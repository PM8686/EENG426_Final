magic
tech sky130l
timestamp 1731220558
<< m2 >>
rect 134 3648 140 3649
rect 110 3645 116 3646
rect 110 3641 111 3645
rect 115 3641 116 3645
rect 134 3644 135 3648
rect 139 3644 140 3648
rect 134 3643 140 3644
rect 214 3648 220 3649
rect 214 3644 215 3648
rect 219 3644 220 3648
rect 214 3643 220 3644
rect 294 3648 300 3649
rect 294 3644 295 3648
rect 299 3644 300 3648
rect 294 3643 300 3644
rect 1830 3645 1836 3646
rect 110 3640 116 3641
rect 1830 3641 1831 3645
rect 1835 3641 1836 3645
rect 1830 3640 1836 3641
rect 110 3628 116 3629
rect 110 3624 111 3628
rect 115 3624 116 3628
rect 110 3623 116 3624
rect 1830 3628 1836 3629
rect 1830 3624 1831 3628
rect 1835 3624 1836 3628
rect 1830 3623 1836 3624
rect 142 3610 148 3611
rect 142 3606 143 3610
rect 147 3606 148 3610
rect 142 3605 148 3606
rect 222 3610 228 3611
rect 222 3606 223 3610
rect 227 3606 228 3610
rect 222 3605 228 3606
rect 302 3610 308 3611
rect 302 3606 303 3610
rect 307 3606 308 3610
rect 302 3605 308 3606
rect 2062 3586 2068 3587
rect 2062 3582 2063 3586
rect 2067 3582 2068 3586
rect 2062 3581 2068 3582
rect 2150 3586 2156 3587
rect 2150 3582 2151 3586
rect 2155 3582 2156 3586
rect 2150 3581 2156 3582
rect 2254 3586 2260 3587
rect 2254 3582 2255 3586
rect 2259 3582 2260 3586
rect 2254 3581 2260 3582
rect 2366 3586 2372 3587
rect 2366 3582 2367 3586
rect 2371 3582 2372 3586
rect 2366 3581 2372 3582
rect 2478 3586 2484 3587
rect 2478 3582 2479 3586
rect 2483 3582 2484 3586
rect 2478 3581 2484 3582
rect 2590 3586 2596 3587
rect 2590 3582 2591 3586
rect 2595 3582 2596 3586
rect 2590 3581 2596 3582
rect 2702 3586 2708 3587
rect 2702 3582 2703 3586
rect 2707 3582 2708 3586
rect 2702 3581 2708 3582
rect 2814 3586 2820 3587
rect 2814 3582 2815 3586
rect 2819 3582 2820 3586
rect 2814 3581 2820 3582
rect 2918 3586 2924 3587
rect 2918 3582 2919 3586
rect 2923 3582 2924 3586
rect 2918 3581 2924 3582
rect 3014 3586 3020 3587
rect 3014 3582 3015 3586
rect 3019 3582 3020 3586
rect 3014 3581 3020 3582
rect 3110 3586 3116 3587
rect 3110 3582 3111 3586
rect 3115 3582 3116 3586
rect 3110 3581 3116 3582
rect 3206 3586 3212 3587
rect 3206 3582 3207 3586
rect 3211 3582 3212 3586
rect 3206 3581 3212 3582
rect 3302 3586 3308 3587
rect 3302 3582 3303 3586
rect 3307 3582 3308 3586
rect 3302 3581 3308 3582
rect 3398 3586 3404 3587
rect 3398 3582 3399 3586
rect 3403 3582 3404 3586
rect 3398 3581 3404 3582
rect 142 3578 148 3579
rect 142 3574 143 3578
rect 147 3574 148 3578
rect 142 3573 148 3574
rect 222 3578 228 3579
rect 222 3574 223 3578
rect 227 3574 228 3578
rect 222 3573 228 3574
rect 342 3578 348 3579
rect 342 3574 343 3578
rect 347 3574 348 3578
rect 342 3573 348 3574
rect 470 3578 476 3579
rect 470 3574 471 3578
rect 475 3574 476 3578
rect 470 3573 476 3574
rect 606 3578 612 3579
rect 606 3574 607 3578
rect 611 3574 612 3578
rect 606 3573 612 3574
rect 742 3578 748 3579
rect 742 3574 743 3578
rect 747 3574 748 3578
rect 742 3573 748 3574
rect 878 3578 884 3579
rect 878 3574 879 3578
rect 883 3574 884 3578
rect 878 3573 884 3574
rect 998 3578 1004 3579
rect 998 3574 999 3578
rect 1003 3574 1004 3578
rect 998 3573 1004 3574
rect 1110 3578 1116 3579
rect 1110 3574 1111 3578
rect 1115 3574 1116 3578
rect 1110 3573 1116 3574
rect 1222 3578 1228 3579
rect 1222 3574 1223 3578
rect 1227 3574 1228 3578
rect 1222 3573 1228 3574
rect 1326 3578 1332 3579
rect 1326 3574 1327 3578
rect 1331 3574 1332 3578
rect 1326 3573 1332 3574
rect 1422 3578 1428 3579
rect 1422 3574 1423 3578
rect 1427 3574 1428 3578
rect 1422 3573 1428 3574
rect 1526 3578 1532 3579
rect 1526 3574 1527 3578
rect 1531 3574 1532 3578
rect 1526 3573 1532 3574
rect 1630 3578 1636 3579
rect 1630 3574 1631 3578
rect 1635 3574 1636 3578
rect 1630 3573 1636 3574
rect 1870 3568 1876 3569
rect 1870 3564 1871 3568
rect 1875 3564 1876 3568
rect 1870 3563 1876 3564
rect 3590 3568 3596 3569
rect 3590 3564 3591 3568
rect 3595 3564 3596 3568
rect 3590 3563 3596 3564
rect 110 3560 116 3561
rect 110 3556 111 3560
rect 115 3556 116 3560
rect 110 3555 116 3556
rect 1830 3560 1836 3561
rect 1830 3556 1831 3560
rect 1835 3556 1836 3560
rect 1830 3555 1836 3556
rect 1870 3551 1876 3552
rect 1870 3547 1871 3551
rect 1875 3547 1876 3551
rect 3590 3551 3596 3552
rect 1870 3546 1876 3547
rect 2054 3548 2060 3549
rect 2054 3544 2055 3548
rect 2059 3544 2060 3548
rect 110 3543 116 3544
rect 110 3539 111 3543
rect 115 3539 116 3543
rect 1830 3543 1836 3544
rect 2054 3543 2060 3544
rect 2142 3548 2148 3549
rect 2142 3544 2143 3548
rect 2147 3544 2148 3548
rect 2142 3543 2148 3544
rect 2246 3548 2252 3549
rect 2246 3544 2247 3548
rect 2251 3544 2252 3548
rect 2246 3543 2252 3544
rect 2358 3548 2364 3549
rect 2358 3544 2359 3548
rect 2363 3544 2364 3548
rect 2358 3543 2364 3544
rect 2470 3548 2476 3549
rect 2470 3544 2471 3548
rect 2475 3544 2476 3548
rect 2470 3543 2476 3544
rect 2582 3548 2588 3549
rect 2582 3544 2583 3548
rect 2587 3544 2588 3548
rect 2582 3543 2588 3544
rect 2694 3548 2700 3549
rect 2694 3544 2695 3548
rect 2699 3544 2700 3548
rect 2694 3543 2700 3544
rect 2806 3548 2812 3549
rect 2806 3544 2807 3548
rect 2811 3544 2812 3548
rect 2806 3543 2812 3544
rect 2910 3548 2916 3549
rect 2910 3544 2911 3548
rect 2915 3544 2916 3548
rect 2910 3543 2916 3544
rect 3006 3548 3012 3549
rect 3006 3544 3007 3548
rect 3011 3544 3012 3548
rect 3006 3543 3012 3544
rect 3102 3548 3108 3549
rect 3102 3544 3103 3548
rect 3107 3544 3108 3548
rect 3102 3543 3108 3544
rect 3198 3548 3204 3549
rect 3198 3544 3199 3548
rect 3203 3544 3204 3548
rect 3198 3543 3204 3544
rect 3294 3548 3300 3549
rect 3294 3544 3295 3548
rect 3299 3544 3300 3548
rect 3294 3543 3300 3544
rect 3390 3548 3396 3549
rect 3390 3544 3391 3548
rect 3395 3544 3396 3548
rect 3590 3547 3591 3551
rect 3595 3547 3596 3551
rect 3590 3546 3596 3547
rect 3390 3543 3396 3544
rect 110 3538 116 3539
rect 134 3540 140 3541
rect 134 3536 135 3540
rect 139 3536 140 3540
rect 134 3535 140 3536
rect 214 3540 220 3541
rect 214 3536 215 3540
rect 219 3536 220 3540
rect 214 3535 220 3536
rect 334 3540 340 3541
rect 334 3536 335 3540
rect 339 3536 340 3540
rect 334 3535 340 3536
rect 462 3540 468 3541
rect 462 3536 463 3540
rect 467 3536 468 3540
rect 462 3535 468 3536
rect 598 3540 604 3541
rect 598 3536 599 3540
rect 603 3536 604 3540
rect 598 3535 604 3536
rect 734 3540 740 3541
rect 734 3536 735 3540
rect 739 3536 740 3540
rect 734 3535 740 3536
rect 870 3540 876 3541
rect 870 3536 871 3540
rect 875 3536 876 3540
rect 870 3535 876 3536
rect 990 3540 996 3541
rect 990 3536 991 3540
rect 995 3536 996 3540
rect 990 3535 996 3536
rect 1102 3540 1108 3541
rect 1102 3536 1103 3540
rect 1107 3536 1108 3540
rect 1102 3535 1108 3536
rect 1214 3540 1220 3541
rect 1214 3536 1215 3540
rect 1219 3536 1220 3540
rect 1214 3535 1220 3536
rect 1318 3540 1324 3541
rect 1318 3536 1319 3540
rect 1323 3536 1324 3540
rect 1318 3535 1324 3536
rect 1414 3540 1420 3541
rect 1414 3536 1415 3540
rect 1419 3536 1420 3540
rect 1414 3535 1420 3536
rect 1518 3540 1524 3541
rect 1518 3536 1519 3540
rect 1523 3536 1524 3540
rect 1518 3535 1524 3536
rect 1622 3540 1628 3541
rect 1622 3536 1623 3540
rect 1627 3536 1628 3540
rect 1830 3539 1831 3543
rect 1835 3539 1836 3543
rect 1830 3538 1836 3539
rect 1622 3535 1628 3536
rect 2086 3504 2092 3505
rect 1870 3501 1876 3502
rect 1870 3497 1871 3501
rect 1875 3497 1876 3501
rect 2086 3500 2087 3504
rect 2091 3500 2092 3504
rect 2086 3499 2092 3500
rect 2166 3504 2172 3505
rect 2166 3500 2167 3504
rect 2171 3500 2172 3504
rect 2166 3499 2172 3500
rect 2262 3504 2268 3505
rect 2262 3500 2263 3504
rect 2267 3500 2268 3504
rect 2262 3499 2268 3500
rect 2366 3504 2372 3505
rect 2366 3500 2367 3504
rect 2371 3500 2372 3504
rect 2366 3499 2372 3500
rect 2486 3504 2492 3505
rect 2486 3500 2487 3504
rect 2491 3500 2492 3504
rect 2486 3499 2492 3500
rect 2614 3504 2620 3505
rect 2614 3500 2615 3504
rect 2619 3500 2620 3504
rect 2614 3499 2620 3500
rect 2742 3504 2748 3505
rect 2742 3500 2743 3504
rect 2747 3500 2748 3504
rect 2742 3499 2748 3500
rect 2870 3504 2876 3505
rect 2870 3500 2871 3504
rect 2875 3500 2876 3504
rect 2870 3499 2876 3500
rect 2990 3504 2996 3505
rect 2990 3500 2991 3504
rect 2995 3500 2996 3504
rect 2990 3499 2996 3500
rect 3118 3504 3124 3505
rect 3118 3500 3119 3504
rect 3123 3500 3124 3504
rect 3118 3499 3124 3500
rect 3246 3504 3252 3505
rect 3246 3500 3247 3504
rect 3251 3500 3252 3504
rect 3246 3499 3252 3500
rect 3374 3504 3380 3505
rect 3374 3500 3375 3504
rect 3379 3500 3380 3504
rect 3374 3499 3380 3500
rect 3590 3501 3596 3502
rect 190 3496 196 3497
rect 110 3493 116 3494
rect 110 3489 111 3493
rect 115 3489 116 3493
rect 190 3492 191 3496
rect 195 3492 196 3496
rect 190 3491 196 3492
rect 326 3496 332 3497
rect 326 3492 327 3496
rect 331 3492 332 3496
rect 326 3491 332 3492
rect 470 3496 476 3497
rect 470 3492 471 3496
rect 475 3492 476 3496
rect 470 3491 476 3492
rect 622 3496 628 3497
rect 622 3492 623 3496
rect 627 3492 628 3496
rect 622 3491 628 3492
rect 774 3496 780 3497
rect 774 3492 775 3496
rect 779 3492 780 3496
rect 774 3491 780 3492
rect 918 3496 924 3497
rect 918 3492 919 3496
rect 923 3492 924 3496
rect 918 3491 924 3492
rect 1054 3496 1060 3497
rect 1054 3492 1055 3496
rect 1059 3492 1060 3496
rect 1054 3491 1060 3492
rect 1182 3496 1188 3497
rect 1182 3492 1183 3496
rect 1187 3492 1188 3496
rect 1182 3491 1188 3492
rect 1310 3496 1316 3497
rect 1310 3492 1311 3496
rect 1315 3492 1316 3496
rect 1310 3491 1316 3492
rect 1438 3496 1444 3497
rect 1438 3492 1439 3496
rect 1443 3492 1444 3496
rect 1438 3491 1444 3492
rect 1566 3496 1572 3497
rect 1870 3496 1876 3497
rect 3590 3497 3591 3501
rect 3595 3497 3596 3501
rect 3590 3496 3596 3497
rect 1566 3492 1567 3496
rect 1571 3492 1572 3496
rect 1566 3491 1572 3492
rect 1830 3493 1836 3494
rect 110 3488 116 3489
rect 1830 3489 1831 3493
rect 1835 3489 1836 3493
rect 1830 3488 1836 3489
rect 1870 3484 1876 3485
rect 1870 3480 1871 3484
rect 1875 3480 1876 3484
rect 1870 3479 1876 3480
rect 3590 3484 3596 3485
rect 3590 3480 3591 3484
rect 3595 3480 3596 3484
rect 3590 3479 3596 3480
rect 110 3476 116 3477
rect 110 3472 111 3476
rect 115 3472 116 3476
rect 110 3471 116 3472
rect 1830 3476 1836 3477
rect 1830 3472 1831 3476
rect 1835 3472 1836 3476
rect 1830 3471 1836 3472
rect 2094 3466 2100 3467
rect 2094 3462 2095 3466
rect 2099 3462 2100 3466
rect 2094 3461 2100 3462
rect 2174 3466 2180 3467
rect 2174 3462 2175 3466
rect 2179 3462 2180 3466
rect 2174 3461 2180 3462
rect 2270 3466 2276 3467
rect 2270 3462 2271 3466
rect 2275 3462 2276 3466
rect 2270 3461 2276 3462
rect 2374 3466 2380 3467
rect 2374 3462 2375 3466
rect 2379 3462 2380 3466
rect 2374 3461 2380 3462
rect 2494 3466 2500 3467
rect 2494 3462 2495 3466
rect 2499 3462 2500 3466
rect 2494 3461 2500 3462
rect 2622 3466 2628 3467
rect 2622 3462 2623 3466
rect 2627 3462 2628 3466
rect 2622 3461 2628 3462
rect 2750 3466 2756 3467
rect 2750 3462 2751 3466
rect 2755 3462 2756 3466
rect 2750 3461 2756 3462
rect 2878 3466 2884 3467
rect 2878 3462 2879 3466
rect 2883 3462 2884 3466
rect 2878 3461 2884 3462
rect 2998 3466 3004 3467
rect 2998 3462 2999 3466
rect 3003 3462 3004 3466
rect 2998 3461 3004 3462
rect 3126 3466 3132 3467
rect 3126 3462 3127 3466
rect 3131 3462 3132 3466
rect 3126 3461 3132 3462
rect 3254 3466 3260 3467
rect 3254 3462 3255 3466
rect 3259 3462 3260 3466
rect 3254 3461 3260 3462
rect 3382 3466 3388 3467
rect 3382 3462 3383 3466
rect 3387 3462 3388 3466
rect 3382 3461 3388 3462
rect 198 3458 204 3459
rect 198 3454 199 3458
rect 203 3454 204 3458
rect 198 3453 204 3454
rect 334 3458 340 3459
rect 334 3454 335 3458
rect 339 3454 340 3458
rect 334 3453 340 3454
rect 478 3458 484 3459
rect 478 3454 479 3458
rect 483 3454 484 3458
rect 478 3453 484 3454
rect 630 3458 636 3459
rect 630 3454 631 3458
rect 635 3454 636 3458
rect 630 3453 636 3454
rect 782 3458 788 3459
rect 782 3454 783 3458
rect 787 3454 788 3458
rect 782 3453 788 3454
rect 926 3458 932 3459
rect 926 3454 927 3458
rect 931 3454 932 3458
rect 926 3453 932 3454
rect 1062 3458 1068 3459
rect 1062 3454 1063 3458
rect 1067 3454 1068 3458
rect 1062 3453 1068 3454
rect 1190 3458 1196 3459
rect 1190 3454 1191 3458
rect 1195 3454 1196 3458
rect 1190 3453 1196 3454
rect 1318 3458 1324 3459
rect 1318 3454 1319 3458
rect 1323 3454 1324 3458
rect 1318 3453 1324 3454
rect 1446 3458 1452 3459
rect 1446 3454 1447 3458
rect 1451 3454 1452 3458
rect 1446 3453 1452 3454
rect 1574 3458 1580 3459
rect 1574 3454 1575 3458
rect 1579 3454 1580 3458
rect 1574 3453 1580 3454
rect 150 3426 156 3427
rect 150 3422 151 3426
rect 155 3422 156 3426
rect 150 3421 156 3422
rect 294 3426 300 3427
rect 294 3422 295 3426
rect 299 3422 300 3426
rect 294 3421 300 3422
rect 454 3426 460 3427
rect 454 3422 455 3426
rect 459 3422 460 3426
rect 454 3421 460 3422
rect 622 3426 628 3427
rect 622 3422 623 3426
rect 627 3422 628 3426
rect 622 3421 628 3422
rect 790 3426 796 3427
rect 790 3422 791 3426
rect 795 3422 796 3426
rect 790 3421 796 3422
rect 958 3426 964 3427
rect 958 3422 959 3426
rect 963 3422 964 3426
rect 958 3421 964 3422
rect 1118 3426 1124 3427
rect 1118 3422 1119 3426
rect 1123 3422 1124 3426
rect 1118 3421 1124 3422
rect 1270 3426 1276 3427
rect 1270 3422 1271 3426
rect 1275 3422 1276 3426
rect 1270 3421 1276 3422
rect 1414 3426 1420 3427
rect 1414 3422 1415 3426
rect 1419 3422 1420 3426
rect 1414 3421 1420 3422
rect 1558 3426 1564 3427
rect 1558 3422 1559 3426
rect 1563 3422 1564 3426
rect 1558 3421 1564 3422
rect 1710 3426 1716 3427
rect 1710 3422 1711 3426
rect 1715 3422 1716 3426
rect 1710 3421 1716 3422
rect 2110 3426 2116 3427
rect 2110 3422 2111 3426
rect 2115 3422 2116 3426
rect 2110 3421 2116 3422
rect 2198 3426 2204 3427
rect 2198 3422 2199 3426
rect 2203 3422 2204 3426
rect 2198 3421 2204 3422
rect 2302 3426 2308 3427
rect 2302 3422 2303 3426
rect 2307 3422 2308 3426
rect 2302 3421 2308 3422
rect 2414 3426 2420 3427
rect 2414 3422 2415 3426
rect 2419 3422 2420 3426
rect 2414 3421 2420 3422
rect 2542 3426 2548 3427
rect 2542 3422 2543 3426
rect 2547 3422 2548 3426
rect 2542 3421 2548 3422
rect 2678 3426 2684 3427
rect 2678 3422 2679 3426
rect 2683 3422 2684 3426
rect 2678 3421 2684 3422
rect 2814 3426 2820 3427
rect 2814 3422 2815 3426
rect 2819 3422 2820 3426
rect 2814 3421 2820 3422
rect 2958 3426 2964 3427
rect 2958 3422 2959 3426
rect 2963 3422 2964 3426
rect 2958 3421 2964 3422
rect 3110 3426 3116 3427
rect 3110 3422 3111 3426
rect 3115 3422 3116 3426
rect 3110 3421 3116 3422
rect 3262 3426 3268 3427
rect 3262 3422 3263 3426
rect 3267 3422 3268 3426
rect 3262 3421 3268 3422
rect 3422 3426 3428 3427
rect 3422 3422 3423 3426
rect 3427 3422 3428 3426
rect 3422 3421 3428 3422
rect 110 3408 116 3409
rect 110 3404 111 3408
rect 115 3404 116 3408
rect 110 3403 116 3404
rect 1830 3408 1836 3409
rect 1830 3404 1831 3408
rect 1835 3404 1836 3408
rect 1830 3403 1836 3404
rect 1870 3408 1876 3409
rect 1870 3404 1871 3408
rect 1875 3404 1876 3408
rect 1870 3403 1876 3404
rect 3590 3408 3596 3409
rect 3590 3404 3591 3408
rect 3595 3404 3596 3408
rect 3590 3403 3596 3404
rect 110 3391 116 3392
rect 110 3387 111 3391
rect 115 3387 116 3391
rect 1830 3391 1836 3392
rect 110 3386 116 3387
rect 142 3388 148 3389
rect 142 3384 143 3388
rect 147 3384 148 3388
rect 142 3383 148 3384
rect 286 3388 292 3389
rect 286 3384 287 3388
rect 291 3384 292 3388
rect 286 3383 292 3384
rect 446 3388 452 3389
rect 446 3384 447 3388
rect 451 3384 452 3388
rect 446 3383 452 3384
rect 614 3388 620 3389
rect 614 3384 615 3388
rect 619 3384 620 3388
rect 614 3383 620 3384
rect 782 3388 788 3389
rect 782 3384 783 3388
rect 787 3384 788 3388
rect 782 3383 788 3384
rect 950 3388 956 3389
rect 950 3384 951 3388
rect 955 3384 956 3388
rect 950 3383 956 3384
rect 1110 3388 1116 3389
rect 1110 3384 1111 3388
rect 1115 3384 1116 3388
rect 1110 3383 1116 3384
rect 1262 3388 1268 3389
rect 1262 3384 1263 3388
rect 1267 3384 1268 3388
rect 1262 3383 1268 3384
rect 1406 3388 1412 3389
rect 1406 3384 1407 3388
rect 1411 3384 1412 3388
rect 1406 3383 1412 3384
rect 1550 3388 1556 3389
rect 1550 3384 1551 3388
rect 1555 3384 1556 3388
rect 1550 3383 1556 3384
rect 1702 3388 1708 3389
rect 1702 3384 1703 3388
rect 1707 3384 1708 3388
rect 1830 3387 1831 3391
rect 1835 3387 1836 3391
rect 1830 3386 1836 3387
rect 1870 3391 1876 3392
rect 1870 3387 1871 3391
rect 1875 3387 1876 3391
rect 3590 3391 3596 3392
rect 1870 3386 1876 3387
rect 2102 3388 2108 3389
rect 1702 3383 1708 3384
rect 2102 3384 2103 3388
rect 2107 3384 2108 3388
rect 2102 3383 2108 3384
rect 2190 3388 2196 3389
rect 2190 3384 2191 3388
rect 2195 3384 2196 3388
rect 2190 3383 2196 3384
rect 2294 3388 2300 3389
rect 2294 3384 2295 3388
rect 2299 3384 2300 3388
rect 2294 3383 2300 3384
rect 2406 3388 2412 3389
rect 2406 3384 2407 3388
rect 2411 3384 2412 3388
rect 2406 3383 2412 3384
rect 2534 3388 2540 3389
rect 2534 3384 2535 3388
rect 2539 3384 2540 3388
rect 2534 3383 2540 3384
rect 2670 3388 2676 3389
rect 2670 3384 2671 3388
rect 2675 3384 2676 3388
rect 2670 3383 2676 3384
rect 2806 3388 2812 3389
rect 2806 3384 2807 3388
rect 2811 3384 2812 3388
rect 2806 3383 2812 3384
rect 2950 3388 2956 3389
rect 2950 3384 2951 3388
rect 2955 3384 2956 3388
rect 2950 3383 2956 3384
rect 3102 3388 3108 3389
rect 3102 3384 3103 3388
rect 3107 3384 3108 3388
rect 3102 3383 3108 3384
rect 3254 3388 3260 3389
rect 3254 3384 3255 3388
rect 3259 3384 3260 3388
rect 3254 3383 3260 3384
rect 3414 3388 3420 3389
rect 3414 3384 3415 3388
rect 3419 3384 3420 3388
rect 3590 3387 3591 3391
rect 3595 3387 3596 3391
rect 3590 3386 3596 3387
rect 3414 3383 3420 3384
rect 206 3344 212 3345
rect 110 3341 116 3342
rect 110 3337 111 3341
rect 115 3337 116 3341
rect 206 3340 207 3344
rect 211 3340 212 3344
rect 206 3339 212 3340
rect 334 3344 340 3345
rect 334 3340 335 3344
rect 339 3340 340 3344
rect 334 3339 340 3340
rect 470 3344 476 3345
rect 470 3340 471 3344
rect 475 3340 476 3344
rect 470 3339 476 3340
rect 622 3344 628 3345
rect 622 3340 623 3344
rect 627 3340 628 3344
rect 622 3339 628 3340
rect 782 3344 788 3345
rect 782 3340 783 3344
rect 787 3340 788 3344
rect 782 3339 788 3340
rect 942 3344 948 3345
rect 942 3340 943 3344
rect 947 3340 948 3344
rect 942 3339 948 3340
rect 1102 3344 1108 3345
rect 1102 3340 1103 3344
rect 1107 3340 1108 3344
rect 1102 3339 1108 3340
rect 1262 3344 1268 3345
rect 1262 3340 1263 3344
rect 1267 3340 1268 3344
rect 1262 3339 1268 3340
rect 1422 3344 1428 3345
rect 1422 3340 1423 3344
rect 1427 3340 1428 3344
rect 1422 3339 1428 3340
rect 1582 3344 1588 3345
rect 1582 3340 1583 3344
rect 1587 3340 1588 3344
rect 1582 3339 1588 3340
rect 1742 3344 1748 3345
rect 1742 3340 1743 3344
rect 1747 3340 1748 3344
rect 1742 3339 1748 3340
rect 1830 3341 1836 3342
rect 110 3336 116 3337
rect 1830 3337 1831 3341
rect 1835 3337 1836 3341
rect 2126 3340 2132 3341
rect 1830 3336 1836 3337
rect 1870 3337 1876 3338
rect 1870 3333 1871 3337
rect 1875 3333 1876 3337
rect 2126 3336 2127 3340
rect 2131 3336 2132 3340
rect 2126 3335 2132 3336
rect 2222 3340 2228 3341
rect 2222 3336 2223 3340
rect 2227 3336 2228 3340
rect 2222 3335 2228 3336
rect 2334 3340 2340 3341
rect 2334 3336 2335 3340
rect 2339 3336 2340 3340
rect 2334 3335 2340 3336
rect 2454 3340 2460 3341
rect 2454 3336 2455 3340
rect 2459 3336 2460 3340
rect 2454 3335 2460 3336
rect 2582 3340 2588 3341
rect 2582 3336 2583 3340
rect 2587 3336 2588 3340
rect 2582 3335 2588 3336
rect 2718 3340 2724 3341
rect 2718 3336 2719 3340
rect 2723 3336 2724 3340
rect 2718 3335 2724 3336
rect 2862 3340 2868 3341
rect 2862 3336 2863 3340
rect 2867 3336 2868 3340
rect 2862 3335 2868 3336
rect 3006 3340 3012 3341
rect 3006 3336 3007 3340
rect 3011 3336 3012 3340
rect 3006 3335 3012 3336
rect 3158 3340 3164 3341
rect 3158 3336 3159 3340
rect 3163 3336 3164 3340
rect 3158 3335 3164 3336
rect 3310 3340 3316 3341
rect 3310 3336 3311 3340
rect 3315 3336 3316 3340
rect 3310 3335 3316 3336
rect 3470 3340 3476 3341
rect 3470 3336 3471 3340
rect 3475 3336 3476 3340
rect 3470 3335 3476 3336
rect 3590 3337 3596 3338
rect 1870 3332 1876 3333
rect 3590 3333 3591 3337
rect 3595 3333 3596 3337
rect 3590 3332 3596 3333
rect 110 3324 116 3325
rect 110 3320 111 3324
rect 115 3320 116 3324
rect 110 3319 116 3320
rect 1830 3324 1836 3325
rect 1830 3320 1831 3324
rect 1835 3320 1836 3324
rect 1830 3319 1836 3320
rect 1870 3320 1876 3321
rect 1870 3316 1871 3320
rect 1875 3316 1876 3320
rect 1870 3315 1876 3316
rect 3590 3320 3596 3321
rect 3590 3316 3591 3320
rect 3595 3316 3596 3320
rect 3590 3315 3596 3316
rect 214 3306 220 3307
rect 214 3302 215 3306
rect 219 3302 220 3306
rect 214 3301 220 3302
rect 342 3306 348 3307
rect 342 3302 343 3306
rect 347 3302 348 3306
rect 342 3301 348 3302
rect 478 3306 484 3307
rect 478 3302 479 3306
rect 483 3302 484 3306
rect 478 3301 484 3302
rect 630 3306 636 3307
rect 630 3302 631 3306
rect 635 3302 636 3306
rect 630 3301 636 3302
rect 790 3306 796 3307
rect 790 3302 791 3306
rect 795 3302 796 3306
rect 790 3301 796 3302
rect 950 3306 956 3307
rect 950 3302 951 3306
rect 955 3302 956 3306
rect 950 3301 956 3302
rect 1110 3306 1116 3307
rect 1110 3302 1111 3306
rect 1115 3302 1116 3306
rect 1110 3301 1116 3302
rect 1270 3306 1276 3307
rect 1270 3302 1271 3306
rect 1275 3302 1276 3306
rect 1270 3301 1276 3302
rect 1430 3306 1436 3307
rect 1430 3302 1431 3306
rect 1435 3302 1436 3306
rect 1430 3301 1436 3302
rect 1590 3306 1596 3307
rect 1590 3302 1591 3306
rect 1595 3302 1596 3306
rect 1590 3301 1596 3302
rect 1750 3306 1756 3307
rect 1750 3302 1751 3306
rect 1755 3302 1756 3306
rect 1750 3301 1756 3302
rect 2134 3302 2140 3303
rect 2134 3298 2135 3302
rect 2139 3298 2140 3302
rect 2134 3297 2140 3298
rect 2230 3302 2236 3303
rect 2230 3298 2231 3302
rect 2235 3298 2236 3302
rect 2230 3297 2236 3298
rect 2342 3302 2348 3303
rect 2342 3298 2343 3302
rect 2347 3298 2348 3302
rect 2342 3297 2348 3298
rect 2462 3302 2468 3303
rect 2462 3298 2463 3302
rect 2467 3298 2468 3302
rect 2462 3297 2468 3298
rect 2590 3302 2596 3303
rect 2590 3298 2591 3302
rect 2595 3298 2596 3302
rect 2590 3297 2596 3298
rect 2726 3302 2732 3303
rect 2726 3298 2727 3302
rect 2731 3298 2732 3302
rect 2726 3297 2732 3298
rect 2870 3302 2876 3303
rect 2870 3298 2871 3302
rect 2875 3298 2876 3302
rect 2870 3297 2876 3298
rect 3014 3302 3020 3303
rect 3014 3298 3015 3302
rect 3019 3298 3020 3302
rect 3014 3297 3020 3298
rect 3166 3302 3172 3303
rect 3166 3298 3167 3302
rect 3171 3298 3172 3302
rect 3166 3297 3172 3298
rect 3318 3302 3324 3303
rect 3318 3298 3319 3302
rect 3323 3298 3324 3302
rect 3318 3297 3324 3298
rect 3478 3302 3484 3303
rect 3478 3298 3479 3302
rect 3483 3298 3484 3302
rect 3478 3297 3484 3298
rect 350 3270 356 3271
rect 350 3266 351 3270
rect 355 3266 356 3270
rect 350 3265 356 3266
rect 454 3270 460 3271
rect 454 3266 455 3270
rect 459 3266 460 3270
rect 454 3265 460 3266
rect 574 3270 580 3271
rect 574 3266 575 3270
rect 579 3266 580 3270
rect 574 3265 580 3266
rect 702 3270 708 3271
rect 702 3266 703 3270
rect 707 3266 708 3270
rect 702 3265 708 3266
rect 838 3270 844 3271
rect 838 3266 839 3270
rect 843 3266 844 3270
rect 838 3265 844 3266
rect 982 3270 988 3271
rect 982 3266 983 3270
rect 987 3266 988 3270
rect 982 3265 988 3266
rect 1118 3270 1124 3271
rect 1118 3266 1119 3270
rect 1123 3266 1124 3270
rect 1118 3265 1124 3266
rect 1254 3270 1260 3271
rect 1254 3266 1255 3270
rect 1259 3266 1260 3270
rect 1254 3265 1260 3266
rect 1382 3270 1388 3271
rect 1382 3266 1383 3270
rect 1387 3266 1388 3270
rect 1382 3265 1388 3266
rect 1510 3270 1516 3271
rect 1510 3266 1511 3270
rect 1515 3266 1516 3270
rect 1510 3265 1516 3266
rect 1638 3270 1644 3271
rect 1638 3266 1639 3270
rect 1643 3266 1644 3270
rect 1638 3265 1644 3266
rect 1750 3270 1756 3271
rect 1750 3266 1751 3270
rect 1755 3266 1756 3270
rect 1750 3265 1756 3266
rect 2134 3258 2140 3259
rect 2134 3254 2135 3258
rect 2139 3254 2140 3258
rect 2134 3253 2140 3254
rect 2278 3258 2284 3259
rect 2278 3254 2279 3258
rect 2283 3254 2284 3258
rect 2278 3253 2284 3254
rect 2414 3258 2420 3259
rect 2414 3254 2415 3258
rect 2419 3254 2420 3258
rect 2414 3253 2420 3254
rect 2550 3258 2556 3259
rect 2550 3254 2551 3258
rect 2555 3254 2556 3258
rect 2550 3253 2556 3254
rect 2686 3258 2692 3259
rect 2686 3254 2687 3258
rect 2691 3254 2692 3258
rect 2686 3253 2692 3254
rect 2822 3258 2828 3259
rect 2822 3254 2823 3258
rect 2827 3254 2828 3258
rect 2822 3253 2828 3254
rect 2958 3258 2964 3259
rect 2958 3254 2959 3258
rect 2963 3254 2964 3258
rect 2958 3253 2964 3254
rect 3094 3258 3100 3259
rect 3094 3254 3095 3258
rect 3099 3254 3100 3258
rect 3094 3253 3100 3254
rect 3230 3258 3236 3259
rect 3230 3254 3231 3258
rect 3235 3254 3236 3258
rect 3230 3253 3236 3254
rect 3374 3258 3380 3259
rect 3374 3254 3375 3258
rect 3379 3254 3380 3258
rect 3374 3253 3380 3254
rect 3510 3258 3516 3259
rect 3510 3254 3511 3258
rect 3515 3254 3516 3258
rect 3510 3253 3516 3254
rect 110 3252 116 3253
rect 110 3248 111 3252
rect 115 3248 116 3252
rect 110 3247 116 3248
rect 1830 3252 1836 3253
rect 1830 3248 1831 3252
rect 1835 3248 1836 3252
rect 1830 3247 1836 3248
rect 1870 3240 1876 3241
rect 1870 3236 1871 3240
rect 1875 3236 1876 3240
rect 110 3235 116 3236
rect 110 3231 111 3235
rect 115 3231 116 3235
rect 1830 3235 1836 3236
rect 1870 3235 1876 3236
rect 3590 3240 3596 3241
rect 3590 3236 3591 3240
rect 3595 3236 3596 3240
rect 3590 3235 3596 3236
rect 110 3230 116 3231
rect 342 3232 348 3233
rect 342 3228 343 3232
rect 347 3228 348 3232
rect 342 3227 348 3228
rect 446 3232 452 3233
rect 446 3228 447 3232
rect 451 3228 452 3232
rect 446 3227 452 3228
rect 566 3232 572 3233
rect 566 3228 567 3232
rect 571 3228 572 3232
rect 566 3227 572 3228
rect 694 3232 700 3233
rect 694 3228 695 3232
rect 699 3228 700 3232
rect 694 3227 700 3228
rect 830 3232 836 3233
rect 830 3228 831 3232
rect 835 3228 836 3232
rect 830 3227 836 3228
rect 974 3232 980 3233
rect 974 3228 975 3232
rect 979 3228 980 3232
rect 974 3227 980 3228
rect 1110 3232 1116 3233
rect 1110 3228 1111 3232
rect 1115 3228 1116 3232
rect 1110 3227 1116 3228
rect 1246 3232 1252 3233
rect 1246 3228 1247 3232
rect 1251 3228 1252 3232
rect 1246 3227 1252 3228
rect 1374 3232 1380 3233
rect 1374 3228 1375 3232
rect 1379 3228 1380 3232
rect 1374 3227 1380 3228
rect 1502 3232 1508 3233
rect 1502 3228 1503 3232
rect 1507 3228 1508 3232
rect 1502 3227 1508 3228
rect 1630 3232 1636 3233
rect 1630 3228 1631 3232
rect 1635 3228 1636 3232
rect 1630 3227 1636 3228
rect 1742 3232 1748 3233
rect 1742 3228 1743 3232
rect 1747 3228 1748 3232
rect 1830 3231 1831 3235
rect 1835 3231 1836 3235
rect 1830 3230 1836 3231
rect 1742 3227 1748 3228
rect 1870 3223 1876 3224
rect 1870 3219 1871 3223
rect 1875 3219 1876 3223
rect 3590 3223 3596 3224
rect 1870 3218 1876 3219
rect 2126 3220 2132 3221
rect 2126 3216 2127 3220
rect 2131 3216 2132 3220
rect 2126 3215 2132 3216
rect 2270 3220 2276 3221
rect 2270 3216 2271 3220
rect 2275 3216 2276 3220
rect 2270 3215 2276 3216
rect 2406 3220 2412 3221
rect 2406 3216 2407 3220
rect 2411 3216 2412 3220
rect 2406 3215 2412 3216
rect 2542 3220 2548 3221
rect 2542 3216 2543 3220
rect 2547 3216 2548 3220
rect 2542 3215 2548 3216
rect 2678 3220 2684 3221
rect 2678 3216 2679 3220
rect 2683 3216 2684 3220
rect 2678 3215 2684 3216
rect 2814 3220 2820 3221
rect 2814 3216 2815 3220
rect 2819 3216 2820 3220
rect 2814 3215 2820 3216
rect 2950 3220 2956 3221
rect 2950 3216 2951 3220
rect 2955 3216 2956 3220
rect 2950 3215 2956 3216
rect 3086 3220 3092 3221
rect 3086 3216 3087 3220
rect 3091 3216 3092 3220
rect 3086 3215 3092 3216
rect 3222 3220 3228 3221
rect 3222 3216 3223 3220
rect 3227 3216 3228 3220
rect 3222 3215 3228 3216
rect 3366 3220 3372 3221
rect 3366 3216 3367 3220
rect 3371 3216 3372 3220
rect 3366 3215 3372 3216
rect 3502 3220 3508 3221
rect 3502 3216 3503 3220
rect 3507 3216 3508 3220
rect 3590 3219 3591 3223
rect 3595 3219 3596 3223
rect 3590 3218 3596 3219
rect 3502 3215 3508 3216
rect 486 3188 492 3189
rect 110 3185 116 3186
rect 110 3181 111 3185
rect 115 3181 116 3185
rect 486 3184 487 3188
rect 491 3184 492 3188
rect 486 3183 492 3184
rect 574 3188 580 3189
rect 574 3184 575 3188
rect 579 3184 580 3188
rect 574 3183 580 3184
rect 662 3188 668 3189
rect 662 3184 663 3188
rect 667 3184 668 3188
rect 662 3183 668 3184
rect 766 3188 772 3189
rect 766 3184 767 3188
rect 771 3184 772 3188
rect 766 3183 772 3184
rect 886 3188 892 3189
rect 886 3184 887 3188
rect 891 3184 892 3188
rect 886 3183 892 3184
rect 1022 3188 1028 3189
rect 1022 3184 1023 3188
rect 1027 3184 1028 3188
rect 1022 3183 1028 3184
rect 1190 3188 1196 3189
rect 1190 3184 1191 3188
rect 1195 3184 1196 3188
rect 1190 3183 1196 3184
rect 1374 3188 1380 3189
rect 1374 3184 1375 3188
rect 1379 3184 1380 3188
rect 1374 3183 1380 3184
rect 1566 3188 1572 3189
rect 1566 3184 1567 3188
rect 1571 3184 1572 3188
rect 1566 3183 1572 3184
rect 1742 3188 1748 3189
rect 1742 3184 1743 3188
rect 1747 3184 1748 3188
rect 1742 3183 1748 3184
rect 1830 3185 1836 3186
rect 110 3180 116 3181
rect 1830 3181 1831 3185
rect 1835 3181 1836 3185
rect 1830 3180 1836 3181
rect 1894 3172 1900 3173
rect 1870 3169 1876 3170
rect 110 3168 116 3169
rect 110 3164 111 3168
rect 115 3164 116 3168
rect 110 3163 116 3164
rect 1830 3168 1836 3169
rect 1830 3164 1831 3168
rect 1835 3164 1836 3168
rect 1870 3165 1871 3169
rect 1875 3165 1876 3169
rect 1894 3168 1895 3172
rect 1899 3168 1900 3172
rect 1894 3167 1900 3168
rect 1990 3172 1996 3173
rect 1990 3168 1991 3172
rect 1995 3168 1996 3172
rect 1990 3167 1996 3168
rect 2118 3172 2124 3173
rect 2118 3168 2119 3172
rect 2123 3168 2124 3172
rect 2118 3167 2124 3168
rect 2246 3172 2252 3173
rect 2246 3168 2247 3172
rect 2251 3168 2252 3172
rect 2246 3167 2252 3168
rect 2382 3172 2388 3173
rect 2382 3168 2383 3172
rect 2387 3168 2388 3172
rect 2382 3167 2388 3168
rect 2510 3172 2516 3173
rect 2510 3168 2511 3172
rect 2515 3168 2516 3172
rect 2510 3167 2516 3168
rect 2638 3172 2644 3173
rect 2638 3168 2639 3172
rect 2643 3168 2644 3172
rect 2638 3167 2644 3168
rect 2766 3172 2772 3173
rect 2766 3168 2767 3172
rect 2771 3168 2772 3172
rect 2766 3167 2772 3168
rect 2894 3172 2900 3173
rect 2894 3168 2895 3172
rect 2899 3168 2900 3172
rect 2894 3167 2900 3168
rect 3030 3172 3036 3173
rect 3030 3168 3031 3172
rect 3035 3168 3036 3172
rect 3030 3167 3036 3168
rect 3174 3172 3180 3173
rect 3174 3168 3175 3172
rect 3179 3168 3180 3172
rect 3174 3167 3180 3168
rect 3326 3172 3332 3173
rect 3326 3168 3327 3172
rect 3331 3168 3332 3172
rect 3326 3167 3332 3168
rect 3486 3172 3492 3173
rect 3486 3168 3487 3172
rect 3491 3168 3492 3172
rect 3486 3167 3492 3168
rect 3590 3169 3596 3170
rect 1870 3164 1876 3165
rect 3590 3165 3591 3169
rect 3595 3165 3596 3169
rect 3590 3164 3596 3165
rect 1830 3163 1836 3164
rect 1870 3152 1876 3153
rect 494 3150 500 3151
rect 494 3146 495 3150
rect 499 3146 500 3150
rect 494 3145 500 3146
rect 582 3150 588 3151
rect 582 3146 583 3150
rect 587 3146 588 3150
rect 582 3145 588 3146
rect 670 3150 676 3151
rect 670 3146 671 3150
rect 675 3146 676 3150
rect 670 3145 676 3146
rect 774 3150 780 3151
rect 774 3146 775 3150
rect 779 3146 780 3150
rect 774 3145 780 3146
rect 894 3150 900 3151
rect 894 3146 895 3150
rect 899 3146 900 3150
rect 894 3145 900 3146
rect 1030 3150 1036 3151
rect 1030 3146 1031 3150
rect 1035 3146 1036 3150
rect 1030 3145 1036 3146
rect 1198 3150 1204 3151
rect 1198 3146 1199 3150
rect 1203 3146 1204 3150
rect 1198 3145 1204 3146
rect 1382 3150 1388 3151
rect 1382 3146 1383 3150
rect 1387 3146 1388 3150
rect 1382 3145 1388 3146
rect 1574 3150 1580 3151
rect 1574 3146 1575 3150
rect 1579 3146 1580 3150
rect 1574 3145 1580 3146
rect 1750 3150 1756 3151
rect 1750 3146 1751 3150
rect 1755 3146 1756 3150
rect 1870 3148 1871 3152
rect 1875 3148 1876 3152
rect 1870 3147 1876 3148
rect 3590 3152 3596 3153
rect 3590 3148 3591 3152
rect 3595 3148 3596 3152
rect 3590 3147 3596 3148
rect 1750 3145 1756 3146
rect 1902 3134 1908 3135
rect 1902 3130 1903 3134
rect 1907 3130 1908 3134
rect 1902 3129 1908 3130
rect 1998 3134 2004 3135
rect 1998 3130 1999 3134
rect 2003 3130 2004 3134
rect 1998 3129 2004 3130
rect 2126 3134 2132 3135
rect 2126 3130 2127 3134
rect 2131 3130 2132 3134
rect 2126 3129 2132 3130
rect 2254 3134 2260 3135
rect 2254 3130 2255 3134
rect 2259 3130 2260 3134
rect 2254 3129 2260 3130
rect 2390 3134 2396 3135
rect 2390 3130 2391 3134
rect 2395 3130 2396 3134
rect 2390 3129 2396 3130
rect 2518 3134 2524 3135
rect 2518 3130 2519 3134
rect 2523 3130 2524 3134
rect 2518 3129 2524 3130
rect 2646 3134 2652 3135
rect 2646 3130 2647 3134
rect 2651 3130 2652 3134
rect 2646 3129 2652 3130
rect 2774 3134 2780 3135
rect 2774 3130 2775 3134
rect 2779 3130 2780 3134
rect 2774 3129 2780 3130
rect 2902 3134 2908 3135
rect 2902 3130 2903 3134
rect 2907 3130 2908 3134
rect 2902 3129 2908 3130
rect 3038 3134 3044 3135
rect 3038 3130 3039 3134
rect 3043 3130 3044 3134
rect 3038 3129 3044 3130
rect 3182 3134 3188 3135
rect 3182 3130 3183 3134
rect 3187 3130 3188 3134
rect 3182 3129 3188 3130
rect 3334 3134 3340 3135
rect 3334 3130 3335 3134
rect 3339 3130 3340 3134
rect 3334 3129 3340 3130
rect 3494 3134 3500 3135
rect 3494 3130 3495 3134
rect 3499 3130 3500 3134
rect 3494 3129 3500 3130
rect 590 3114 596 3115
rect 590 3110 591 3114
rect 595 3110 596 3114
rect 590 3109 596 3110
rect 670 3114 676 3115
rect 670 3110 671 3114
rect 675 3110 676 3114
rect 670 3109 676 3110
rect 758 3114 764 3115
rect 758 3110 759 3114
rect 763 3110 764 3114
rect 758 3109 764 3110
rect 846 3114 852 3115
rect 846 3110 847 3114
rect 851 3110 852 3114
rect 846 3109 852 3110
rect 934 3114 940 3115
rect 934 3110 935 3114
rect 939 3110 940 3114
rect 934 3109 940 3110
rect 1022 3114 1028 3115
rect 1022 3110 1023 3114
rect 1027 3110 1028 3114
rect 1022 3109 1028 3110
rect 1110 3114 1116 3115
rect 1110 3110 1111 3114
rect 1115 3110 1116 3114
rect 1110 3109 1116 3110
rect 1198 3114 1204 3115
rect 1198 3110 1199 3114
rect 1203 3110 1204 3114
rect 1198 3109 1204 3110
rect 1286 3114 1292 3115
rect 1286 3110 1287 3114
rect 1291 3110 1292 3114
rect 1286 3109 1292 3110
rect 1374 3114 1380 3115
rect 1374 3110 1375 3114
rect 1379 3110 1380 3114
rect 1374 3109 1380 3110
rect 110 3096 116 3097
rect 110 3092 111 3096
rect 115 3092 116 3096
rect 110 3091 116 3092
rect 1830 3096 1836 3097
rect 1830 3092 1831 3096
rect 1835 3092 1836 3096
rect 1830 3091 1836 3092
rect 1902 3086 1908 3087
rect 1902 3082 1903 3086
rect 1907 3082 1908 3086
rect 1902 3081 1908 3082
rect 2014 3086 2020 3087
rect 2014 3082 2015 3086
rect 2019 3082 2020 3086
rect 2014 3081 2020 3082
rect 2190 3086 2196 3087
rect 2190 3082 2191 3086
rect 2195 3082 2196 3086
rect 2190 3081 2196 3082
rect 2406 3086 2412 3087
rect 2406 3082 2407 3086
rect 2411 3082 2412 3086
rect 2406 3081 2412 3082
rect 2654 3086 2660 3087
rect 2654 3082 2655 3086
rect 2659 3082 2660 3086
rect 2654 3081 2660 3082
rect 2934 3086 2940 3087
rect 2934 3082 2935 3086
rect 2939 3082 2940 3086
rect 2934 3081 2940 3082
rect 3230 3086 3236 3087
rect 3230 3082 3231 3086
rect 3235 3082 3236 3086
rect 3230 3081 3236 3082
rect 3510 3086 3516 3087
rect 3510 3082 3511 3086
rect 3515 3082 3516 3086
rect 3510 3081 3516 3082
rect 110 3079 116 3080
rect 110 3075 111 3079
rect 115 3075 116 3079
rect 1830 3079 1836 3080
rect 110 3074 116 3075
rect 582 3076 588 3077
rect 582 3072 583 3076
rect 587 3072 588 3076
rect 582 3071 588 3072
rect 662 3076 668 3077
rect 662 3072 663 3076
rect 667 3072 668 3076
rect 662 3071 668 3072
rect 750 3076 756 3077
rect 750 3072 751 3076
rect 755 3072 756 3076
rect 750 3071 756 3072
rect 838 3076 844 3077
rect 838 3072 839 3076
rect 843 3072 844 3076
rect 838 3071 844 3072
rect 926 3076 932 3077
rect 926 3072 927 3076
rect 931 3072 932 3076
rect 926 3071 932 3072
rect 1014 3076 1020 3077
rect 1014 3072 1015 3076
rect 1019 3072 1020 3076
rect 1014 3071 1020 3072
rect 1102 3076 1108 3077
rect 1102 3072 1103 3076
rect 1107 3072 1108 3076
rect 1102 3071 1108 3072
rect 1190 3076 1196 3077
rect 1190 3072 1191 3076
rect 1195 3072 1196 3076
rect 1190 3071 1196 3072
rect 1278 3076 1284 3077
rect 1278 3072 1279 3076
rect 1283 3072 1284 3076
rect 1278 3071 1284 3072
rect 1366 3076 1372 3077
rect 1366 3072 1367 3076
rect 1371 3072 1372 3076
rect 1830 3075 1831 3079
rect 1835 3075 1836 3079
rect 1830 3074 1836 3075
rect 1366 3071 1372 3072
rect 1870 3068 1876 3069
rect 1870 3064 1871 3068
rect 1875 3064 1876 3068
rect 1870 3063 1876 3064
rect 3590 3068 3596 3069
rect 3590 3064 3591 3068
rect 3595 3064 3596 3068
rect 3590 3063 3596 3064
rect 1870 3051 1876 3052
rect 1870 3047 1871 3051
rect 1875 3047 1876 3051
rect 3590 3051 3596 3052
rect 1870 3046 1876 3047
rect 1894 3048 1900 3049
rect 1894 3044 1895 3048
rect 1899 3044 1900 3048
rect 1894 3043 1900 3044
rect 2006 3048 2012 3049
rect 2006 3044 2007 3048
rect 2011 3044 2012 3048
rect 2006 3043 2012 3044
rect 2182 3048 2188 3049
rect 2182 3044 2183 3048
rect 2187 3044 2188 3048
rect 2182 3043 2188 3044
rect 2398 3048 2404 3049
rect 2398 3044 2399 3048
rect 2403 3044 2404 3048
rect 2398 3043 2404 3044
rect 2646 3048 2652 3049
rect 2646 3044 2647 3048
rect 2651 3044 2652 3048
rect 2646 3043 2652 3044
rect 2926 3048 2932 3049
rect 2926 3044 2927 3048
rect 2931 3044 2932 3048
rect 2926 3043 2932 3044
rect 3222 3048 3228 3049
rect 3222 3044 3223 3048
rect 3227 3044 3228 3048
rect 3222 3043 3228 3044
rect 3502 3048 3508 3049
rect 3502 3044 3503 3048
rect 3507 3044 3508 3048
rect 3590 3047 3591 3051
rect 3595 3047 3596 3051
rect 3590 3046 3596 3047
rect 3502 3043 3508 3044
rect 542 3028 548 3029
rect 110 3025 116 3026
rect 110 3021 111 3025
rect 115 3021 116 3025
rect 542 3024 543 3028
rect 547 3024 548 3028
rect 542 3023 548 3024
rect 622 3028 628 3029
rect 622 3024 623 3028
rect 627 3024 628 3028
rect 622 3023 628 3024
rect 710 3028 716 3029
rect 710 3024 711 3028
rect 715 3024 716 3028
rect 710 3023 716 3024
rect 806 3028 812 3029
rect 806 3024 807 3028
rect 811 3024 812 3028
rect 806 3023 812 3024
rect 902 3028 908 3029
rect 902 3024 903 3028
rect 907 3024 908 3028
rect 902 3023 908 3024
rect 998 3028 1004 3029
rect 998 3024 999 3028
rect 1003 3024 1004 3028
rect 998 3023 1004 3024
rect 1086 3028 1092 3029
rect 1086 3024 1087 3028
rect 1091 3024 1092 3028
rect 1086 3023 1092 3024
rect 1182 3028 1188 3029
rect 1182 3024 1183 3028
rect 1187 3024 1188 3028
rect 1182 3023 1188 3024
rect 1278 3028 1284 3029
rect 1278 3024 1279 3028
rect 1283 3024 1284 3028
rect 1278 3023 1284 3024
rect 1374 3028 1380 3029
rect 1374 3024 1375 3028
rect 1379 3024 1380 3028
rect 1374 3023 1380 3024
rect 1470 3028 1476 3029
rect 1470 3024 1471 3028
rect 1475 3024 1476 3028
rect 1470 3023 1476 3024
rect 1830 3025 1836 3026
rect 110 3020 116 3021
rect 1830 3021 1831 3025
rect 1835 3021 1836 3025
rect 1830 3020 1836 3021
rect 110 3008 116 3009
rect 110 3004 111 3008
rect 115 3004 116 3008
rect 110 3003 116 3004
rect 1830 3008 1836 3009
rect 1830 3004 1831 3008
rect 1835 3004 1836 3008
rect 1830 3003 1836 3004
rect 1894 2996 1900 2997
rect 1870 2993 1876 2994
rect 550 2990 556 2991
rect 550 2986 551 2990
rect 555 2986 556 2990
rect 550 2985 556 2986
rect 630 2990 636 2991
rect 630 2986 631 2990
rect 635 2986 636 2990
rect 630 2985 636 2986
rect 718 2990 724 2991
rect 718 2986 719 2990
rect 723 2986 724 2990
rect 718 2985 724 2986
rect 814 2990 820 2991
rect 814 2986 815 2990
rect 819 2986 820 2990
rect 814 2985 820 2986
rect 910 2990 916 2991
rect 910 2986 911 2990
rect 915 2986 916 2990
rect 910 2985 916 2986
rect 1006 2990 1012 2991
rect 1006 2986 1007 2990
rect 1011 2986 1012 2990
rect 1006 2985 1012 2986
rect 1094 2990 1100 2991
rect 1094 2986 1095 2990
rect 1099 2986 1100 2990
rect 1094 2985 1100 2986
rect 1190 2990 1196 2991
rect 1190 2986 1191 2990
rect 1195 2986 1196 2990
rect 1190 2985 1196 2986
rect 1286 2990 1292 2991
rect 1286 2986 1287 2990
rect 1291 2986 1292 2990
rect 1286 2985 1292 2986
rect 1382 2990 1388 2991
rect 1382 2986 1383 2990
rect 1387 2986 1388 2990
rect 1382 2985 1388 2986
rect 1478 2990 1484 2991
rect 1478 2986 1479 2990
rect 1483 2986 1484 2990
rect 1870 2989 1871 2993
rect 1875 2989 1876 2993
rect 1894 2992 1895 2996
rect 1899 2992 1900 2996
rect 1894 2991 1900 2992
rect 2046 2996 2052 2997
rect 2046 2992 2047 2996
rect 2051 2992 2052 2996
rect 2046 2991 2052 2992
rect 2222 2996 2228 2997
rect 2222 2992 2223 2996
rect 2227 2992 2228 2996
rect 2222 2991 2228 2992
rect 2390 2996 2396 2997
rect 2390 2992 2391 2996
rect 2395 2992 2396 2996
rect 2390 2991 2396 2992
rect 2542 2996 2548 2997
rect 2542 2992 2543 2996
rect 2547 2992 2548 2996
rect 2542 2991 2548 2992
rect 2686 2996 2692 2997
rect 2686 2992 2687 2996
rect 2691 2992 2692 2996
rect 2686 2991 2692 2992
rect 2814 2996 2820 2997
rect 2814 2992 2815 2996
rect 2819 2992 2820 2996
rect 2814 2991 2820 2992
rect 2926 2996 2932 2997
rect 2926 2992 2927 2996
rect 2931 2992 2932 2996
rect 2926 2991 2932 2992
rect 3038 2996 3044 2997
rect 3038 2992 3039 2996
rect 3043 2992 3044 2996
rect 3038 2991 3044 2992
rect 3142 2996 3148 2997
rect 3142 2992 3143 2996
rect 3147 2992 3148 2996
rect 3142 2991 3148 2992
rect 3238 2996 3244 2997
rect 3238 2992 3239 2996
rect 3243 2992 3244 2996
rect 3238 2991 3244 2992
rect 3334 2996 3340 2997
rect 3334 2992 3335 2996
rect 3339 2992 3340 2996
rect 3334 2991 3340 2992
rect 3422 2996 3428 2997
rect 3422 2992 3423 2996
rect 3427 2992 3428 2996
rect 3422 2991 3428 2992
rect 3502 2996 3508 2997
rect 3502 2992 3503 2996
rect 3507 2992 3508 2996
rect 3502 2991 3508 2992
rect 3590 2993 3596 2994
rect 1870 2988 1876 2989
rect 3590 2989 3591 2993
rect 3595 2989 3596 2993
rect 3590 2988 3596 2989
rect 1478 2985 1484 2986
rect 1870 2976 1876 2977
rect 1870 2972 1871 2976
rect 1875 2972 1876 2976
rect 1870 2971 1876 2972
rect 3590 2976 3596 2977
rect 3590 2972 3591 2976
rect 3595 2972 3596 2976
rect 3590 2971 3596 2972
rect 470 2958 476 2959
rect 470 2954 471 2958
rect 475 2954 476 2958
rect 470 2953 476 2954
rect 574 2958 580 2959
rect 574 2954 575 2958
rect 579 2954 580 2958
rect 574 2953 580 2954
rect 686 2958 692 2959
rect 686 2954 687 2958
rect 691 2954 692 2958
rect 686 2953 692 2954
rect 806 2958 812 2959
rect 806 2954 807 2958
rect 811 2954 812 2958
rect 806 2953 812 2954
rect 942 2958 948 2959
rect 942 2954 943 2958
rect 947 2954 948 2958
rect 942 2953 948 2954
rect 1086 2958 1092 2959
rect 1086 2954 1087 2958
rect 1091 2954 1092 2958
rect 1086 2953 1092 2954
rect 1246 2958 1252 2959
rect 1246 2954 1247 2958
rect 1251 2954 1252 2958
rect 1246 2953 1252 2954
rect 1414 2958 1420 2959
rect 1414 2954 1415 2958
rect 1419 2954 1420 2958
rect 1414 2953 1420 2954
rect 1590 2958 1596 2959
rect 1590 2954 1591 2958
rect 1595 2954 1596 2958
rect 1590 2953 1596 2954
rect 1750 2958 1756 2959
rect 1750 2954 1751 2958
rect 1755 2954 1756 2958
rect 1750 2953 1756 2954
rect 1902 2958 1908 2959
rect 1902 2954 1903 2958
rect 1907 2954 1908 2958
rect 1902 2953 1908 2954
rect 2054 2958 2060 2959
rect 2054 2954 2055 2958
rect 2059 2954 2060 2958
rect 2054 2953 2060 2954
rect 2230 2958 2236 2959
rect 2230 2954 2231 2958
rect 2235 2954 2236 2958
rect 2230 2953 2236 2954
rect 2398 2958 2404 2959
rect 2398 2954 2399 2958
rect 2403 2954 2404 2958
rect 2398 2953 2404 2954
rect 2550 2958 2556 2959
rect 2550 2954 2551 2958
rect 2555 2954 2556 2958
rect 2550 2953 2556 2954
rect 2694 2958 2700 2959
rect 2694 2954 2695 2958
rect 2699 2954 2700 2958
rect 2694 2953 2700 2954
rect 2822 2958 2828 2959
rect 2822 2954 2823 2958
rect 2827 2954 2828 2958
rect 2822 2953 2828 2954
rect 2934 2958 2940 2959
rect 2934 2954 2935 2958
rect 2939 2954 2940 2958
rect 2934 2953 2940 2954
rect 3046 2958 3052 2959
rect 3046 2954 3047 2958
rect 3051 2954 3052 2958
rect 3046 2953 3052 2954
rect 3150 2958 3156 2959
rect 3150 2954 3151 2958
rect 3155 2954 3156 2958
rect 3150 2953 3156 2954
rect 3246 2958 3252 2959
rect 3246 2954 3247 2958
rect 3251 2954 3252 2958
rect 3246 2953 3252 2954
rect 3342 2958 3348 2959
rect 3342 2954 3343 2958
rect 3347 2954 3348 2958
rect 3342 2953 3348 2954
rect 3430 2958 3436 2959
rect 3430 2954 3431 2958
rect 3435 2954 3436 2958
rect 3430 2953 3436 2954
rect 3510 2958 3516 2959
rect 3510 2954 3511 2958
rect 3515 2954 3516 2958
rect 3510 2953 3516 2954
rect 110 2940 116 2941
rect 110 2936 111 2940
rect 115 2936 116 2940
rect 110 2935 116 2936
rect 1830 2940 1836 2941
rect 1830 2936 1831 2940
rect 1835 2936 1836 2940
rect 1830 2935 1836 2936
rect 1902 2926 1908 2927
rect 110 2923 116 2924
rect 110 2919 111 2923
rect 115 2919 116 2923
rect 1830 2923 1836 2924
rect 110 2918 116 2919
rect 462 2920 468 2921
rect 462 2916 463 2920
rect 467 2916 468 2920
rect 462 2915 468 2916
rect 566 2920 572 2921
rect 566 2916 567 2920
rect 571 2916 572 2920
rect 566 2915 572 2916
rect 678 2920 684 2921
rect 678 2916 679 2920
rect 683 2916 684 2920
rect 678 2915 684 2916
rect 798 2920 804 2921
rect 798 2916 799 2920
rect 803 2916 804 2920
rect 798 2915 804 2916
rect 934 2920 940 2921
rect 934 2916 935 2920
rect 939 2916 940 2920
rect 934 2915 940 2916
rect 1078 2920 1084 2921
rect 1078 2916 1079 2920
rect 1083 2916 1084 2920
rect 1078 2915 1084 2916
rect 1238 2920 1244 2921
rect 1238 2916 1239 2920
rect 1243 2916 1244 2920
rect 1238 2915 1244 2916
rect 1406 2920 1412 2921
rect 1406 2916 1407 2920
rect 1411 2916 1412 2920
rect 1406 2915 1412 2916
rect 1582 2920 1588 2921
rect 1582 2916 1583 2920
rect 1587 2916 1588 2920
rect 1582 2915 1588 2916
rect 1742 2920 1748 2921
rect 1742 2916 1743 2920
rect 1747 2916 1748 2920
rect 1830 2919 1831 2923
rect 1835 2919 1836 2923
rect 1902 2922 1903 2926
rect 1907 2922 1908 2926
rect 1902 2921 1908 2922
rect 2086 2926 2092 2927
rect 2086 2922 2087 2926
rect 2091 2922 2092 2926
rect 2086 2921 2092 2922
rect 2294 2926 2300 2927
rect 2294 2922 2295 2926
rect 2299 2922 2300 2926
rect 2294 2921 2300 2922
rect 2486 2926 2492 2927
rect 2486 2922 2487 2926
rect 2491 2922 2492 2926
rect 2486 2921 2492 2922
rect 2670 2926 2676 2927
rect 2670 2922 2671 2926
rect 2675 2922 2676 2926
rect 2670 2921 2676 2922
rect 2838 2926 2844 2927
rect 2838 2922 2839 2926
rect 2843 2922 2844 2926
rect 2838 2921 2844 2922
rect 2998 2926 3004 2927
rect 2998 2922 2999 2926
rect 3003 2922 3004 2926
rect 2998 2921 3004 2922
rect 3150 2926 3156 2927
rect 3150 2922 3151 2926
rect 3155 2922 3156 2926
rect 3150 2921 3156 2922
rect 3302 2926 3308 2927
rect 3302 2922 3303 2926
rect 3307 2922 3308 2926
rect 3302 2921 3308 2922
rect 3454 2926 3460 2927
rect 3454 2922 3455 2926
rect 3459 2922 3460 2926
rect 3454 2921 3460 2922
rect 1830 2918 1836 2919
rect 1742 2915 1748 2916
rect 1870 2908 1876 2909
rect 1870 2904 1871 2908
rect 1875 2904 1876 2908
rect 1870 2903 1876 2904
rect 3590 2908 3596 2909
rect 3590 2904 3591 2908
rect 3595 2904 3596 2908
rect 3590 2903 3596 2904
rect 1870 2891 1876 2892
rect 1870 2887 1871 2891
rect 1875 2887 1876 2891
rect 3590 2891 3596 2892
rect 1870 2886 1876 2887
rect 1894 2888 1900 2889
rect 1894 2884 1895 2888
rect 1899 2884 1900 2888
rect 1894 2883 1900 2884
rect 2078 2888 2084 2889
rect 2078 2884 2079 2888
rect 2083 2884 2084 2888
rect 2078 2883 2084 2884
rect 2286 2888 2292 2889
rect 2286 2884 2287 2888
rect 2291 2884 2292 2888
rect 2286 2883 2292 2884
rect 2478 2888 2484 2889
rect 2478 2884 2479 2888
rect 2483 2884 2484 2888
rect 2478 2883 2484 2884
rect 2662 2888 2668 2889
rect 2662 2884 2663 2888
rect 2667 2884 2668 2888
rect 2662 2883 2668 2884
rect 2830 2888 2836 2889
rect 2830 2884 2831 2888
rect 2835 2884 2836 2888
rect 2830 2883 2836 2884
rect 2990 2888 2996 2889
rect 2990 2884 2991 2888
rect 2995 2884 2996 2888
rect 2990 2883 2996 2884
rect 3142 2888 3148 2889
rect 3142 2884 3143 2888
rect 3147 2884 3148 2888
rect 3142 2883 3148 2884
rect 3294 2888 3300 2889
rect 3294 2884 3295 2888
rect 3299 2884 3300 2888
rect 3294 2883 3300 2884
rect 3446 2888 3452 2889
rect 3446 2884 3447 2888
rect 3451 2884 3452 2888
rect 3590 2887 3591 2891
rect 3595 2887 3596 2891
rect 3590 2886 3596 2887
rect 3446 2883 3452 2884
rect 310 2876 316 2877
rect 110 2873 116 2874
rect 110 2869 111 2873
rect 115 2869 116 2873
rect 310 2872 311 2876
rect 315 2872 316 2876
rect 310 2871 316 2872
rect 430 2876 436 2877
rect 430 2872 431 2876
rect 435 2872 436 2876
rect 430 2871 436 2872
rect 550 2876 556 2877
rect 550 2872 551 2876
rect 555 2872 556 2876
rect 550 2871 556 2872
rect 678 2876 684 2877
rect 678 2872 679 2876
rect 683 2872 684 2876
rect 678 2871 684 2872
rect 814 2876 820 2877
rect 814 2872 815 2876
rect 819 2872 820 2876
rect 814 2871 820 2872
rect 950 2876 956 2877
rect 950 2872 951 2876
rect 955 2872 956 2876
rect 950 2871 956 2872
rect 1086 2876 1092 2877
rect 1086 2872 1087 2876
rect 1091 2872 1092 2876
rect 1086 2871 1092 2872
rect 1222 2876 1228 2877
rect 1222 2872 1223 2876
rect 1227 2872 1228 2876
rect 1222 2871 1228 2872
rect 1358 2876 1364 2877
rect 1358 2872 1359 2876
rect 1363 2872 1364 2876
rect 1358 2871 1364 2872
rect 1494 2876 1500 2877
rect 1494 2872 1495 2876
rect 1499 2872 1500 2876
rect 1494 2871 1500 2872
rect 1630 2876 1636 2877
rect 1630 2872 1631 2876
rect 1635 2872 1636 2876
rect 1630 2871 1636 2872
rect 1742 2876 1748 2877
rect 1742 2872 1743 2876
rect 1747 2872 1748 2876
rect 1742 2871 1748 2872
rect 1830 2873 1836 2874
rect 110 2868 116 2869
rect 1830 2869 1831 2873
rect 1835 2869 1836 2873
rect 1830 2868 1836 2869
rect 110 2856 116 2857
rect 110 2852 111 2856
rect 115 2852 116 2856
rect 110 2851 116 2852
rect 1830 2856 1836 2857
rect 1830 2852 1831 2856
rect 1835 2852 1836 2856
rect 1830 2851 1836 2852
rect 318 2838 324 2839
rect 318 2834 319 2838
rect 323 2834 324 2838
rect 318 2833 324 2834
rect 438 2838 444 2839
rect 438 2834 439 2838
rect 443 2834 444 2838
rect 438 2833 444 2834
rect 558 2838 564 2839
rect 558 2834 559 2838
rect 563 2834 564 2838
rect 558 2833 564 2834
rect 686 2838 692 2839
rect 686 2834 687 2838
rect 691 2834 692 2838
rect 686 2833 692 2834
rect 822 2838 828 2839
rect 822 2834 823 2838
rect 827 2834 828 2838
rect 822 2833 828 2834
rect 958 2838 964 2839
rect 958 2834 959 2838
rect 963 2834 964 2838
rect 958 2833 964 2834
rect 1094 2838 1100 2839
rect 1094 2834 1095 2838
rect 1099 2834 1100 2838
rect 1094 2833 1100 2834
rect 1230 2838 1236 2839
rect 1230 2834 1231 2838
rect 1235 2834 1236 2838
rect 1230 2833 1236 2834
rect 1366 2838 1372 2839
rect 1366 2834 1367 2838
rect 1371 2834 1372 2838
rect 1366 2833 1372 2834
rect 1502 2838 1508 2839
rect 1502 2834 1503 2838
rect 1507 2834 1508 2838
rect 1502 2833 1508 2834
rect 1638 2838 1644 2839
rect 1638 2834 1639 2838
rect 1643 2834 1644 2838
rect 1638 2833 1644 2834
rect 1750 2838 1756 2839
rect 1750 2834 1751 2838
rect 1755 2834 1756 2838
rect 2134 2836 2140 2837
rect 1750 2833 1756 2834
rect 1870 2833 1876 2834
rect 1870 2829 1871 2833
rect 1875 2829 1876 2833
rect 2134 2832 2135 2836
rect 2139 2832 2140 2836
rect 2134 2831 2140 2832
rect 2262 2836 2268 2837
rect 2262 2832 2263 2836
rect 2267 2832 2268 2836
rect 2262 2831 2268 2832
rect 2390 2836 2396 2837
rect 2390 2832 2391 2836
rect 2395 2832 2396 2836
rect 2390 2831 2396 2832
rect 2518 2836 2524 2837
rect 2518 2832 2519 2836
rect 2523 2832 2524 2836
rect 2518 2831 2524 2832
rect 2646 2836 2652 2837
rect 2646 2832 2647 2836
rect 2651 2832 2652 2836
rect 2646 2831 2652 2832
rect 2766 2836 2772 2837
rect 2766 2832 2767 2836
rect 2771 2832 2772 2836
rect 2766 2831 2772 2832
rect 2886 2836 2892 2837
rect 2886 2832 2887 2836
rect 2891 2832 2892 2836
rect 2886 2831 2892 2832
rect 3006 2836 3012 2837
rect 3006 2832 3007 2836
rect 3011 2832 3012 2836
rect 3006 2831 3012 2832
rect 3134 2836 3140 2837
rect 3134 2832 3135 2836
rect 3139 2832 3140 2836
rect 3134 2831 3140 2832
rect 3590 2833 3596 2834
rect 1870 2828 1876 2829
rect 3590 2829 3591 2833
rect 3595 2829 3596 2833
rect 3590 2828 3596 2829
rect 1870 2816 1876 2817
rect 1870 2812 1871 2816
rect 1875 2812 1876 2816
rect 1870 2811 1876 2812
rect 3590 2816 3596 2817
rect 3590 2812 3591 2816
rect 3595 2812 3596 2816
rect 3590 2811 3596 2812
rect 166 2806 172 2807
rect 166 2802 167 2806
rect 171 2802 172 2806
rect 166 2801 172 2802
rect 302 2806 308 2807
rect 302 2802 303 2806
rect 307 2802 308 2806
rect 302 2801 308 2802
rect 446 2806 452 2807
rect 446 2802 447 2806
rect 451 2802 452 2806
rect 446 2801 452 2802
rect 606 2806 612 2807
rect 606 2802 607 2806
rect 611 2802 612 2806
rect 606 2801 612 2802
rect 782 2806 788 2807
rect 782 2802 783 2806
rect 787 2802 788 2806
rect 782 2801 788 2802
rect 958 2806 964 2807
rect 958 2802 959 2806
rect 963 2802 964 2806
rect 958 2801 964 2802
rect 1142 2806 1148 2807
rect 1142 2802 1143 2806
rect 1147 2802 1148 2806
rect 1142 2801 1148 2802
rect 1334 2806 1340 2807
rect 1334 2802 1335 2806
rect 1339 2802 1340 2806
rect 1334 2801 1340 2802
rect 1534 2806 1540 2807
rect 1534 2802 1535 2806
rect 1539 2802 1540 2806
rect 1534 2801 1540 2802
rect 1734 2806 1740 2807
rect 1734 2802 1735 2806
rect 1739 2802 1740 2806
rect 1734 2801 1740 2802
rect 2142 2798 2148 2799
rect 2142 2794 2143 2798
rect 2147 2794 2148 2798
rect 2142 2793 2148 2794
rect 2270 2798 2276 2799
rect 2270 2794 2271 2798
rect 2275 2794 2276 2798
rect 2270 2793 2276 2794
rect 2398 2798 2404 2799
rect 2398 2794 2399 2798
rect 2403 2794 2404 2798
rect 2398 2793 2404 2794
rect 2526 2798 2532 2799
rect 2526 2794 2527 2798
rect 2531 2794 2532 2798
rect 2526 2793 2532 2794
rect 2654 2798 2660 2799
rect 2654 2794 2655 2798
rect 2659 2794 2660 2798
rect 2654 2793 2660 2794
rect 2774 2798 2780 2799
rect 2774 2794 2775 2798
rect 2779 2794 2780 2798
rect 2774 2793 2780 2794
rect 2894 2798 2900 2799
rect 2894 2794 2895 2798
rect 2899 2794 2900 2798
rect 2894 2793 2900 2794
rect 3014 2798 3020 2799
rect 3014 2794 3015 2798
rect 3019 2794 3020 2798
rect 3014 2793 3020 2794
rect 3142 2798 3148 2799
rect 3142 2794 3143 2798
rect 3147 2794 3148 2798
rect 3142 2793 3148 2794
rect 110 2788 116 2789
rect 110 2784 111 2788
rect 115 2784 116 2788
rect 110 2783 116 2784
rect 1830 2788 1836 2789
rect 1830 2784 1831 2788
rect 1835 2784 1836 2788
rect 1830 2783 1836 2784
rect 110 2771 116 2772
rect 110 2767 111 2771
rect 115 2767 116 2771
rect 1830 2771 1836 2772
rect 110 2766 116 2767
rect 158 2768 164 2769
rect 158 2764 159 2768
rect 163 2764 164 2768
rect 158 2763 164 2764
rect 294 2768 300 2769
rect 294 2764 295 2768
rect 299 2764 300 2768
rect 294 2763 300 2764
rect 438 2768 444 2769
rect 438 2764 439 2768
rect 443 2764 444 2768
rect 438 2763 444 2764
rect 598 2768 604 2769
rect 598 2764 599 2768
rect 603 2764 604 2768
rect 598 2763 604 2764
rect 774 2768 780 2769
rect 774 2764 775 2768
rect 779 2764 780 2768
rect 774 2763 780 2764
rect 950 2768 956 2769
rect 950 2764 951 2768
rect 955 2764 956 2768
rect 950 2763 956 2764
rect 1134 2768 1140 2769
rect 1134 2764 1135 2768
rect 1139 2764 1140 2768
rect 1134 2763 1140 2764
rect 1326 2768 1332 2769
rect 1326 2764 1327 2768
rect 1331 2764 1332 2768
rect 1326 2763 1332 2764
rect 1526 2768 1532 2769
rect 1526 2764 1527 2768
rect 1531 2764 1532 2768
rect 1526 2763 1532 2764
rect 1726 2768 1732 2769
rect 1726 2764 1727 2768
rect 1731 2764 1732 2768
rect 1830 2767 1831 2771
rect 1835 2767 1836 2771
rect 1830 2766 1836 2767
rect 1726 2763 1732 2764
rect 2230 2758 2236 2759
rect 2230 2754 2231 2758
rect 2235 2754 2236 2758
rect 2230 2753 2236 2754
rect 2310 2758 2316 2759
rect 2310 2754 2311 2758
rect 2315 2754 2316 2758
rect 2310 2753 2316 2754
rect 2390 2758 2396 2759
rect 2390 2754 2391 2758
rect 2395 2754 2396 2758
rect 2390 2753 2396 2754
rect 2470 2758 2476 2759
rect 2470 2754 2471 2758
rect 2475 2754 2476 2758
rect 2470 2753 2476 2754
rect 2550 2758 2556 2759
rect 2550 2754 2551 2758
rect 2555 2754 2556 2758
rect 2550 2753 2556 2754
rect 2638 2758 2644 2759
rect 2638 2754 2639 2758
rect 2643 2754 2644 2758
rect 2638 2753 2644 2754
rect 2726 2758 2732 2759
rect 2726 2754 2727 2758
rect 2731 2754 2732 2758
rect 2726 2753 2732 2754
rect 2814 2758 2820 2759
rect 2814 2754 2815 2758
rect 2819 2754 2820 2758
rect 2814 2753 2820 2754
rect 2902 2758 2908 2759
rect 2902 2754 2903 2758
rect 2907 2754 2908 2758
rect 2902 2753 2908 2754
rect 2990 2758 2996 2759
rect 2990 2754 2991 2758
rect 2995 2754 2996 2758
rect 2990 2753 2996 2754
rect 1870 2740 1876 2741
rect 1870 2736 1871 2740
rect 1875 2736 1876 2740
rect 1870 2735 1876 2736
rect 3590 2740 3596 2741
rect 3590 2736 3591 2740
rect 3595 2736 3596 2740
rect 3590 2735 3596 2736
rect 1870 2723 1876 2724
rect 134 2720 140 2721
rect 110 2717 116 2718
rect 110 2713 111 2717
rect 115 2713 116 2717
rect 134 2716 135 2720
rect 139 2716 140 2720
rect 134 2715 140 2716
rect 246 2720 252 2721
rect 246 2716 247 2720
rect 251 2716 252 2720
rect 246 2715 252 2716
rect 390 2720 396 2721
rect 390 2716 391 2720
rect 395 2716 396 2720
rect 390 2715 396 2716
rect 550 2720 556 2721
rect 550 2716 551 2720
rect 555 2716 556 2720
rect 550 2715 556 2716
rect 710 2720 716 2721
rect 710 2716 711 2720
rect 715 2716 716 2720
rect 710 2715 716 2716
rect 878 2720 884 2721
rect 878 2716 879 2720
rect 883 2716 884 2720
rect 878 2715 884 2716
rect 1038 2720 1044 2721
rect 1038 2716 1039 2720
rect 1043 2716 1044 2720
rect 1038 2715 1044 2716
rect 1198 2720 1204 2721
rect 1198 2716 1199 2720
rect 1203 2716 1204 2720
rect 1198 2715 1204 2716
rect 1358 2720 1364 2721
rect 1358 2716 1359 2720
rect 1363 2716 1364 2720
rect 1358 2715 1364 2716
rect 1518 2720 1524 2721
rect 1518 2716 1519 2720
rect 1523 2716 1524 2720
rect 1518 2715 1524 2716
rect 1686 2720 1692 2721
rect 1686 2716 1687 2720
rect 1691 2716 1692 2720
rect 1870 2719 1871 2723
rect 1875 2719 1876 2723
rect 3590 2723 3596 2724
rect 1870 2718 1876 2719
rect 2222 2720 2228 2721
rect 1686 2715 1692 2716
rect 1830 2717 1836 2718
rect 110 2712 116 2713
rect 1830 2713 1831 2717
rect 1835 2713 1836 2717
rect 2222 2716 2223 2720
rect 2227 2716 2228 2720
rect 2222 2715 2228 2716
rect 2302 2720 2308 2721
rect 2302 2716 2303 2720
rect 2307 2716 2308 2720
rect 2302 2715 2308 2716
rect 2382 2720 2388 2721
rect 2382 2716 2383 2720
rect 2387 2716 2388 2720
rect 2382 2715 2388 2716
rect 2462 2720 2468 2721
rect 2462 2716 2463 2720
rect 2467 2716 2468 2720
rect 2462 2715 2468 2716
rect 2542 2720 2548 2721
rect 2542 2716 2543 2720
rect 2547 2716 2548 2720
rect 2542 2715 2548 2716
rect 2630 2720 2636 2721
rect 2630 2716 2631 2720
rect 2635 2716 2636 2720
rect 2630 2715 2636 2716
rect 2718 2720 2724 2721
rect 2718 2716 2719 2720
rect 2723 2716 2724 2720
rect 2718 2715 2724 2716
rect 2806 2720 2812 2721
rect 2806 2716 2807 2720
rect 2811 2716 2812 2720
rect 2806 2715 2812 2716
rect 2894 2720 2900 2721
rect 2894 2716 2895 2720
rect 2899 2716 2900 2720
rect 2894 2715 2900 2716
rect 2982 2720 2988 2721
rect 2982 2716 2983 2720
rect 2987 2716 2988 2720
rect 3590 2719 3591 2723
rect 3595 2719 3596 2723
rect 3590 2718 3596 2719
rect 2982 2715 2988 2716
rect 1830 2712 1836 2713
rect 110 2700 116 2701
rect 110 2696 111 2700
rect 115 2696 116 2700
rect 110 2695 116 2696
rect 1830 2700 1836 2701
rect 1830 2696 1831 2700
rect 1835 2696 1836 2700
rect 1830 2695 1836 2696
rect 142 2682 148 2683
rect 142 2678 143 2682
rect 147 2678 148 2682
rect 142 2677 148 2678
rect 254 2682 260 2683
rect 254 2678 255 2682
rect 259 2678 260 2682
rect 254 2677 260 2678
rect 398 2682 404 2683
rect 398 2678 399 2682
rect 403 2678 404 2682
rect 398 2677 404 2678
rect 558 2682 564 2683
rect 558 2678 559 2682
rect 563 2678 564 2682
rect 558 2677 564 2678
rect 718 2682 724 2683
rect 718 2678 719 2682
rect 723 2678 724 2682
rect 718 2677 724 2678
rect 886 2682 892 2683
rect 886 2678 887 2682
rect 891 2678 892 2682
rect 886 2677 892 2678
rect 1046 2682 1052 2683
rect 1046 2678 1047 2682
rect 1051 2678 1052 2682
rect 1046 2677 1052 2678
rect 1206 2682 1212 2683
rect 1206 2678 1207 2682
rect 1211 2678 1212 2682
rect 1206 2677 1212 2678
rect 1366 2682 1372 2683
rect 1366 2678 1367 2682
rect 1371 2678 1372 2682
rect 1366 2677 1372 2678
rect 1526 2682 1532 2683
rect 1526 2678 1527 2682
rect 1531 2678 1532 2682
rect 1526 2677 1532 2678
rect 1694 2682 1700 2683
rect 1694 2678 1695 2682
rect 1699 2678 1700 2682
rect 1694 2677 1700 2678
rect 2238 2676 2244 2677
rect 1870 2673 1876 2674
rect 1870 2669 1871 2673
rect 1875 2669 1876 2673
rect 2238 2672 2239 2676
rect 2243 2672 2244 2676
rect 2238 2671 2244 2672
rect 2318 2676 2324 2677
rect 2318 2672 2319 2676
rect 2323 2672 2324 2676
rect 2318 2671 2324 2672
rect 2398 2676 2404 2677
rect 2398 2672 2399 2676
rect 2403 2672 2404 2676
rect 2398 2671 2404 2672
rect 2478 2676 2484 2677
rect 2478 2672 2479 2676
rect 2483 2672 2484 2676
rect 2478 2671 2484 2672
rect 2558 2676 2564 2677
rect 2558 2672 2559 2676
rect 2563 2672 2564 2676
rect 2558 2671 2564 2672
rect 2638 2676 2644 2677
rect 2638 2672 2639 2676
rect 2643 2672 2644 2676
rect 2638 2671 2644 2672
rect 2718 2676 2724 2677
rect 2718 2672 2719 2676
rect 2723 2672 2724 2676
rect 2718 2671 2724 2672
rect 2798 2676 2804 2677
rect 2798 2672 2799 2676
rect 2803 2672 2804 2676
rect 2798 2671 2804 2672
rect 2878 2676 2884 2677
rect 2878 2672 2879 2676
rect 2883 2672 2884 2676
rect 2878 2671 2884 2672
rect 2958 2676 2964 2677
rect 2958 2672 2959 2676
rect 2963 2672 2964 2676
rect 2958 2671 2964 2672
rect 3590 2673 3596 2674
rect 1870 2668 1876 2669
rect 3590 2669 3591 2673
rect 3595 2669 3596 2673
rect 3590 2668 3596 2669
rect 1870 2656 1876 2657
rect 1870 2652 1871 2656
rect 1875 2652 1876 2656
rect 1870 2651 1876 2652
rect 3590 2656 3596 2657
rect 3590 2652 3591 2656
rect 3595 2652 3596 2656
rect 3590 2651 3596 2652
rect 142 2650 148 2651
rect 142 2646 143 2650
rect 147 2646 148 2650
rect 142 2645 148 2646
rect 254 2650 260 2651
rect 254 2646 255 2650
rect 259 2646 260 2650
rect 254 2645 260 2646
rect 398 2650 404 2651
rect 398 2646 399 2650
rect 403 2646 404 2650
rect 398 2645 404 2646
rect 550 2650 556 2651
rect 550 2646 551 2650
rect 555 2646 556 2650
rect 550 2645 556 2646
rect 710 2650 716 2651
rect 710 2646 711 2650
rect 715 2646 716 2650
rect 710 2645 716 2646
rect 878 2650 884 2651
rect 878 2646 879 2650
rect 883 2646 884 2650
rect 878 2645 884 2646
rect 1046 2650 1052 2651
rect 1046 2646 1047 2650
rect 1051 2646 1052 2650
rect 1046 2645 1052 2646
rect 1214 2650 1220 2651
rect 1214 2646 1215 2650
rect 1219 2646 1220 2650
rect 1214 2645 1220 2646
rect 1390 2650 1396 2651
rect 1390 2646 1391 2650
rect 1395 2646 1396 2650
rect 1390 2645 1396 2646
rect 1566 2650 1572 2651
rect 1566 2646 1567 2650
rect 1571 2646 1572 2650
rect 1566 2645 1572 2646
rect 2246 2638 2252 2639
rect 2246 2634 2247 2638
rect 2251 2634 2252 2638
rect 2246 2633 2252 2634
rect 2326 2638 2332 2639
rect 2326 2634 2327 2638
rect 2331 2634 2332 2638
rect 2326 2633 2332 2634
rect 2406 2638 2412 2639
rect 2406 2634 2407 2638
rect 2411 2634 2412 2638
rect 2406 2633 2412 2634
rect 2486 2638 2492 2639
rect 2486 2634 2487 2638
rect 2491 2634 2492 2638
rect 2486 2633 2492 2634
rect 2566 2638 2572 2639
rect 2566 2634 2567 2638
rect 2571 2634 2572 2638
rect 2566 2633 2572 2634
rect 2646 2638 2652 2639
rect 2646 2634 2647 2638
rect 2651 2634 2652 2638
rect 2646 2633 2652 2634
rect 2726 2638 2732 2639
rect 2726 2634 2727 2638
rect 2731 2634 2732 2638
rect 2726 2633 2732 2634
rect 2806 2638 2812 2639
rect 2806 2634 2807 2638
rect 2811 2634 2812 2638
rect 2806 2633 2812 2634
rect 2886 2638 2892 2639
rect 2886 2634 2887 2638
rect 2891 2634 2892 2638
rect 2886 2633 2892 2634
rect 2966 2638 2972 2639
rect 2966 2634 2967 2638
rect 2971 2634 2972 2638
rect 2966 2633 2972 2634
rect 110 2632 116 2633
rect 110 2628 111 2632
rect 115 2628 116 2632
rect 110 2627 116 2628
rect 1830 2632 1836 2633
rect 1830 2628 1831 2632
rect 1835 2628 1836 2632
rect 1830 2627 1836 2628
rect 110 2615 116 2616
rect 110 2611 111 2615
rect 115 2611 116 2615
rect 1830 2615 1836 2616
rect 110 2610 116 2611
rect 134 2612 140 2613
rect 134 2608 135 2612
rect 139 2608 140 2612
rect 134 2607 140 2608
rect 246 2612 252 2613
rect 246 2608 247 2612
rect 251 2608 252 2612
rect 246 2607 252 2608
rect 390 2612 396 2613
rect 390 2608 391 2612
rect 395 2608 396 2612
rect 390 2607 396 2608
rect 542 2612 548 2613
rect 542 2608 543 2612
rect 547 2608 548 2612
rect 542 2607 548 2608
rect 702 2612 708 2613
rect 702 2608 703 2612
rect 707 2608 708 2612
rect 702 2607 708 2608
rect 870 2612 876 2613
rect 870 2608 871 2612
rect 875 2608 876 2612
rect 870 2607 876 2608
rect 1038 2612 1044 2613
rect 1038 2608 1039 2612
rect 1043 2608 1044 2612
rect 1038 2607 1044 2608
rect 1206 2612 1212 2613
rect 1206 2608 1207 2612
rect 1211 2608 1212 2612
rect 1206 2607 1212 2608
rect 1382 2612 1388 2613
rect 1382 2608 1383 2612
rect 1387 2608 1388 2612
rect 1382 2607 1388 2608
rect 1558 2612 1564 2613
rect 1558 2608 1559 2612
rect 1563 2608 1564 2612
rect 1830 2611 1831 2615
rect 1835 2611 1836 2615
rect 1830 2610 1836 2611
rect 1558 2607 1564 2608
rect 2190 2598 2196 2599
rect 2190 2594 2191 2598
rect 2195 2594 2196 2598
rect 2190 2593 2196 2594
rect 2270 2598 2276 2599
rect 2270 2594 2271 2598
rect 2275 2594 2276 2598
rect 2270 2593 2276 2594
rect 2350 2598 2356 2599
rect 2350 2594 2351 2598
rect 2355 2594 2356 2598
rect 2350 2593 2356 2594
rect 2430 2598 2436 2599
rect 2430 2594 2431 2598
rect 2435 2594 2436 2598
rect 2430 2593 2436 2594
rect 2510 2598 2516 2599
rect 2510 2594 2511 2598
rect 2515 2594 2516 2598
rect 2510 2593 2516 2594
rect 2590 2598 2596 2599
rect 2590 2594 2591 2598
rect 2595 2594 2596 2598
rect 2590 2593 2596 2594
rect 2670 2598 2676 2599
rect 2670 2594 2671 2598
rect 2675 2594 2676 2598
rect 2670 2593 2676 2594
rect 2750 2598 2756 2599
rect 2750 2594 2751 2598
rect 2755 2594 2756 2598
rect 2750 2593 2756 2594
rect 2830 2598 2836 2599
rect 2830 2594 2831 2598
rect 2835 2594 2836 2598
rect 2830 2593 2836 2594
rect 2910 2598 2916 2599
rect 2910 2594 2911 2598
rect 2915 2594 2916 2598
rect 2910 2593 2916 2594
rect 2990 2598 2996 2599
rect 2990 2594 2991 2598
rect 2995 2594 2996 2598
rect 2990 2593 2996 2594
rect 1870 2580 1876 2581
rect 1870 2576 1871 2580
rect 1875 2576 1876 2580
rect 1870 2575 1876 2576
rect 3590 2580 3596 2581
rect 3590 2576 3591 2580
rect 3595 2576 3596 2580
rect 3590 2575 3596 2576
rect 158 2564 164 2565
rect 110 2561 116 2562
rect 110 2557 111 2561
rect 115 2557 116 2561
rect 158 2560 159 2564
rect 163 2560 164 2564
rect 158 2559 164 2560
rect 278 2564 284 2565
rect 278 2560 279 2564
rect 283 2560 284 2564
rect 278 2559 284 2560
rect 414 2564 420 2565
rect 414 2560 415 2564
rect 419 2560 420 2564
rect 414 2559 420 2560
rect 558 2564 564 2565
rect 558 2560 559 2564
rect 563 2560 564 2564
rect 558 2559 564 2560
rect 702 2564 708 2565
rect 702 2560 703 2564
rect 707 2560 708 2564
rect 702 2559 708 2560
rect 846 2564 852 2565
rect 846 2560 847 2564
rect 851 2560 852 2564
rect 846 2559 852 2560
rect 982 2564 988 2565
rect 982 2560 983 2564
rect 987 2560 988 2564
rect 982 2559 988 2560
rect 1118 2564 1124 2565
rect 1118 2560 1119 2564
rect 1123 2560 1124 2564
rect 1118 2559 1124 2560
rect 1254 2564 1260 2565
rect 1254 2560 1255 2564
rect 1259 2560 1260 2564
rect 1254 2559 1260 2560
rect 1390 2564 1396 2565
rect 1390 2560 1391 2564
rect 1395 2560 1396 2564
rect 1390 2559 1396 2560
rect 1526 2564 1532 2565
rect 1526 2560 1527 2564
rect 1531 2560 1532 2564
rect 1870 2563 1876 2564
rect 1526 2559 1532 2560
rect 1830 2561 1836 2562
rect 110 2556 116 2557
rect 1830 2557 1831 2561
rect 1835 2557 1836 2561
rect 1870 2559 1871 2563
rect 1875 2559 1876 2563
rect 3590 2563 3596 2564
rect 1870 2558 1876 2559
rect 2182 2560 2188 2561
rect 1830 2556 1836 2557
rect 2182 2556 2183 2560
rect 2187 2556 2188 2560
rect 2182 2555 2188 2556
rect 2262 2560 2268 2561
rect 2262 2556 2263 2560
rect 2267 2556 2268 2560
rect 2262 2555 2268 2556
rect 2342 2560 2348 2561
rect 2342 2556 2343 2560
rect 2347 2556 2348 2560
rect 2342 2555 2348 2556
rect 2422 2560 2428 2561
rect 2422 2556 2423 2560
rect 2427 2556 2428 2560
rect 2422 2555 2428 2556
rect 2502 2560 2508 2561
rect 2502 2556 2503 2560
rect 2507 2556 2508 2560
rect 2502 2555 2508 2556
rect 2582 2560 2588 2561
rect 2582 2556 2583 2560
rect 2587 2556 2588 2560
rect 2582 2555 2588 2556
rect 2662 2560 2668 2561
rect 2662 2556 2663 2560
rect 2667 2556 2668 2560
rect 2662 2555 2668 2556
rect 2742 2560 2748 2561
rect 2742 2556 2743 2560
rect 2747 2556 2748 2560
rect 2742 2555 2748 2556
rect 2822 2560 2828 2561
rect 2822 2556 2823 2560
rect 2827 2556 2828 2560
rect 2822 2555 2828 2556
rect 2902 2560 2908 2561
rect 2902 2556 2903 2560
rect 2907 2556 2908 2560
rect 2902 2555 2908 2556
rect 2982 2560 2988 2561
rect 2982 2556 2983 2560
rect 2987 2556 2988 2560
rect 3590 2559 3591 2563
rect 3595 2559 3596 2563
rect 3590 2558 3596 2559
rect 2982 2555 2988 2556
rect 110 2544 116 2545
rect 110 2540 111 2544
rect 115 2540 116 2544
rect 110 2539 116 2540
rect 1830 2544 1836 2545
rect 1830 2540 1831 2544
rect 1835 2540 1836 2544
rect 1830 2539 1836 2540
rect 166 2526 172 2527
rect 166 2522 167 2526
rect 171 2522 172 2526
rect 166 2521 172 2522
rect 286 2526 292 2527
rect 286 2522 287 2526
rect 291 2522 292 2526
rect 286 2521 292 2522
rect 422 2526 428 2527
rect 422 2522 423 2526
rect 427 2522 428 2526
rect 422 2521 428 2522
rect 566 2526 572 2527
rect 566 2522 567 2526
rect 571 2522 572 2526
rect 566 2521 572 2522
rect 710 2526 716 2527
rect 710 2522 711 2526
rect 715 2522 716 2526
rect 710 2521 716 2522
rect 854 2526 860 2527
rect 854 2522 855 2526
rect 859 2522 860 2526
rect 854 2521 860 2522
rect 990 2526 996 2527
rect 990 2522 991 2526
rect 995 2522 996 2526
rect 990 2521 996 2522
rect 1126 2526 1132 2527
rect 1126 2522 1127 2526
rect 1131 2522 1132 2526
rect 1126 2521 1132 2522
rect 1262 2526 1268 2527
rect 1262 2522 1263 2526
rect 1267 2522 1268 2526
rect 1262 2521 1268 2522
rect 1398 2526 1404 2527
rect 1398 2522 1399 2526
rect 1403 2522 1404 2526
rect 1398 2521 1404 2522
rect 1534 2526 1540 2527
rect 1534 2522 1535 2526
rect 1539 2522 1540 2526
rect 1534 2521 1540 2522
rect 2118 2508 2124 2509
rect 1870 2505 1876 2506
rect 1870 2501 1871 2505
rect 1875 2501 1876 2505
rect 2118 2504 2119 2508
rect 2123 2504 2124 2508
rect 2118 2503 2124 2504
rect 2206 2508 2212 2509
rect 2206 2504 2207 2508
rect 2211 2504 2212 2508
rect 2206 2503 2212 2504
rect 2302 2508 2308 2509
rect 2302 2504 2303 2508
rect 2307 2504 2308 2508
rect 2302 2503 2308 2504
rect 2398 2508 2404 2509
rect 2398 2504 2399 2508
rect 2403 2504 2404 2508
rect 2398 2503 2404 2504
rect 2494 2508 2500 2509
rect 2494 2504 2495 2508
rect 2499 2504 2500 2508
rect 2494 2503 2500 2504
rect 2590 2508 2596 2509
rect 2590 2504 2591 2508
rect 2595 2504 2596 2508
rect 2590 2503 2596 2504
rect 2686 2508 2692 2509
rect 2686 2504 2687 2508
rect 2691 2504 2692 2508
rect 2686 2503 2692 2504
rect 2782 2508 2788 2509
rect 2782 2504 2783 2508
rect 2787 2504 2788 2508
rect 2782 2503 2788 2504
rect 2878 2508 2884 2509
rect 2878 2504 2879 2508
rect 2883 2504 2884 2508
rect 2878 2503 2884 2504
rect 2974 2508 2980 2509
rect 2974 2504 2975 2508
rect 2979 2504 2980 2508
rect 2974 2503 2980 2504
rect 3078 2508 3084 2509
rect 3078 2504 3079 2508
rect 3083 2504 3084 2508
rect 3078 2503 3084 2504
rect 3590 2505 3596 2506
rect 1870 2500 1876 2501
rect 3590 2501 3591 2505
rect 3595 2501 3596 2505
rect 3590 2500 3596 2501
rect 334 2490 340 2491
rect 334 2486 335 2490
rect 339 2486 340 2490
rect 334 2485 340 2486
rect 414 2490 420 2491
rect 414 2486 415 2490
rect 419 2486 420 2490
rect 414 2485 420 2486
rect 502 2490 508 2491
rect 502 2486 503 2490
rect 507 2486 508 2490
rect 502 2485 508 2486
rect 598 2490 604 2491
rect 598 2486 599 2490
rect 603 2486 604 2490
rect 598 2485 604 2486
rect 702 2490 708 2491
rect 702 2486 703 2490
rect 707 2486 708 2490
rect 702 2485 708 2486
rect 814 2490 820 2491
rect 814 2486 815 2490
rect 819 2486 820 2490
rect 814 2485 820 2486
rect 934 2490 940 2491
rect 934 2486 935 2490
rect 939 2486 940 2490
rect 934 2485 940 2486
rect 1062 2490 1068 2491
rect 1062 2486 1063 2490
rect 1067 2486 1068 2490
rect 1062 2485 1068 2486
rect 1190 2490 1196 2491
rect 1190 2486 1191 2490
rect 1195 2486 1196 2490
rect 1190 2485 1196 2486
rect 1326 2490 1332 2491
rect 1326 2486 1327 2490
rect 1331 2486 1332 2490
rect 1326 2485 1332 2486
rect 1470 2490 1476 2491
rect 1470 2486 1471 2490
rect 1475 2486 1476 2490
rect 1470 2485 1476 2486
rect 1870 2488 1876 2489
rect 1870 2484 1871 2488
rect 1875 2484 1876 2488
rect 1870 2483 1876 2484
rect 3590 2488 3596 2489
rect 3590 2484 3591 2488
rect 3595 2484 3596 2488
rect 3590 2483 3596 2484
rect 110 2472 116 2473
rect 110 2468 111 2472
rect 115 2468 116 2472
rect 110 2467 116 2468
rect 1830 2472 1836 2473
rect 1830 2468 1831 2472
rect 1835 2468 1836 2472
rect 1830 2467 1836 2468
rect 2126 2470 2132 2471
rect 2126 2466 2127 2470
rect 2131 2466 2132 2470
rect 2126 2465 2132 2466
rect 2214 2470 2220 2471
rect 2214 2466 2215 2470
rect 2219 2466 2220 2470
rect 2214 2465 2220 2466
rect 2310 2470 2316 2471
rect 2310 2466 2311 2470
rect 2315 2466 2316 2470
rect 2310 2465 2316 2466
rect 2406 2470 2412 2471
rect 2406 2466 2407 2470
rect 2411 2466 2412 2470
rect 2406 2465 2412 2466
rect 2502 2470 2508 2471
rect 2502 2466 2503 2470
rect 2507 2466 2508 2470
rect 2502 2465 2508 2466
rect 2598 2470 2604 2471
rect 2598 2466 2599 2470
rect 2603 2466 2604 2470
rect 2598 2465 2604 2466
rect 2694 2470 2700 2471
rect 2694 2466 2695 2470
rect 2699 2466 2700 2470
rect 2694 2465 2700 2466
rect 2790 2470 2796 2471
rect 2790 2466 2791 2470
rect 2795 2466 2796 2470
rect 2790 2465 2796 2466
rect 2886 2470 2892 2471
rect 2886 2466 2887 2470
rect 2891 2466 2892 2470
rect 2886 2465 2892 2466
rect 2982 2470 2988 2471
rect 2982 2466 2983 2470
rect 2987 2466 2988 2470
rect 2982 2465 2988 2466
rect 3086 2470 3092 2471
rect 3086 2466 3087 2470
rect 3091 2466 3092 2470
rect 3086 2465 3092 2466
rect 110 2455 116 2456
rect 110 2451 111 2455
rect 115 2451 116 2455
rect 1830 2455 1836 2456
rect 110 2450 116 2451
rect 326 2452 332 2453
rect 326 2448 327 2452
rect 331 2448 332 2452
rect 326 2447 332 2448
rect 406 2452 412 2453
rect 406 2448 407 2452
rect 411 2448 412 2452
rect 406 2447 412 2448
rect 494 2452 500 2453
rect 494 2448 495 2452
rect 499 2448 500 2452
rect 494 2447 500 2448
rect 590 2452 596 2453
rect 590 2448 591 2452
rect 595 2448 596 2452
rect 590 2447 596 2448
rect 694 2452 700 2453
rect 694 2448 695 2452
rect 699 2448 700 2452
rect 694 2447 700 2448
rect 806 2452 812 2453
rect 806 2448 807 2452
rect 811 2448 812 2452
rect 806 2447 812 2448
rect 926 2452 932 2453
rect 926 2448 927 2452
rect 931 2448 932 2452
rect 926 2447 932 2448
rect 1054 2452 1060 2453
rect 1054 2448 1055 2452
rect 1059 2448 1060 2452
rect 1054 2447 1060 2448
rect 1182 2452 1188 2453
rect 1182 2448 1183 2452
rect 1187 2448 1188 2452
rect 1182 2447 1188 2448
rect 1318 2452 1324 2453
rect 1318 2448 1319 2452
rect 1323 2448 1324 2452
rect 1318 2447 1324 2448
rect 1462 2452 1468 2453
rect 1462 2448 1463 2452
rect 1467 2448 1468 2452
rect 1830 2451 1831 2455
rect 1835 2451 1836 2455
rect 1830 2450 1836 2451
rect 1462 2447 1468 2448
rect 1902 2434 1908 2435
rect 1902 2430 1903 2434
rect 1907 2430 1908 2434
rect 1902 2429 1908 2430
rect 1990 2434 1996 2435
rect 1990 2430 1991 2434
rect 1995 2430 1996 2434
rect 1990 2429 1996 2430
rect 2110 2434 2116 2435
rect 2110 2430 2111 2434
rect 2115 2430 2116 2434
rect 2110 2429 2116 2430
rect 2246 2434 2252 2435
rect 2246 2430 2247 2434
rect 2251 2430 2252 2434
rect 2246 2429 2252 2430
rect 2390 2434 2396 2435
rect 2390 2430 2391 2434
rect 2395 2430 2396 2434
rect 2390 2429 2396 2430
rect 2534 2434 2540 2435
rect 2534 2430 2535 2434
rect 2539 2430 2540 2434
rect 2534 2429 2540 2430
rect 2670 2434 2676 2435
rect 2670 2430 2671 2434
rect 2675 2430 2676 2434
rect 2670 2429 2676 2430
rect 2806 2434 2812 2435
rect 2806 2430 2807 2434
rect 2811 2430 2812 2434
rect 2806 2429 2812 2430
rect 2942 2434 2948 2435
rect 2942 2430 2943 2434
rect 2947 2430 2948 2434
rect 2942 2429 2948 2430
rect 3078 2434 3084 2435
rect 3078 2430 3079 2434
rect 3083 2430 3084 2434
rect 3078 2429 3084 2430
rect 3214 2434 3220 2435
rect 3214 2430 3215 2434
rect 3219 2430 3220 2434
rect 3214 2429 3220 2430
rect 1870 2416 1876 2417
rect 1870 2412 1871 2416
rect 1875 2412 1876 2416
rect 1870 2411 1876 2412
rect 3590 2416 3596 2417
rect 3590 2412 3591 2416
rect 3595 2412 3596 2416
rect 3590 2411 3596 2412
rect 382 2400 388 2401
rect 110 2397 116 2398
rect 110 2393 111 2397
rect 115 2393 116 2397
rect 382 2396 383 2400
rect 387 2396 388 2400
rect 382 2395 388 2396
rect 462 2400 468 2401
rect 462 2396 463 2400
rect 467 2396 468 2400
rect 462 2395 468 2396
rect 542 2400 548 2401
rect 542 2396 543 2400
rect 547 2396 548 2400
rect 542 2395 548 2396
rect 622 2400 628 2401
rect 622 2396 623 2400
rect 627 2396 628 2400
rect 622 2395 628 2396
rect 702 2400 708 2401
rect 702 2396 703 2400
rect 707 2396 708 2400
rect 702 2395 708 2396
rect 782 2400 788 2401
rect 782 2396 783 2400
rect 787 2396 788 2400
rect 782 2395 788 2396
rect 862 2400 868 2401
rect 862 2396 863 2400
rect 867 2396 868 2400
rect 862 2395 868 2396
rect 942 2400 948 2401
rect 942 2396 943 2400
rect 947 2396 948 2400
rect 942 2395 948 2396
rect 1022 2400 1028 2401
rect 1022 2396 1023 2400
rect 1027 2396 1028 2400
rect 1022 2395 1028 2396
rect 1102 2400 1108 2401
rect 1102 2396 1103 2400
rect 1107 2396 1108 2400
rect 1102 2395 1108 2396
rect 1182 2400 1188 2401
rect 1182 2396 1183 2400
rect 1187 2396 1188 2400
rect 1182 2395 1188 2396
rect 1262 2400 1268 2401
rect 1262 2396 1263 2400
rect 1267 2396 1268 2400
rect 1262 2395 1268 2396
rect 1350 2400 1356 2401
rect 1350 2396 1351 2400
rect 1355 2396 1356 2400
rect 1350 2395 1356 2396
rect 1438 2400 1444 2401
rect 1438 2396 1439 2400
rect 1443 2396 1444 2400
rect 1438 2395 1444 2396
rect 1526 2400 1532 2401
rect 1526 2396 1527 2400
rect 1531 2396 1532 2400
rect 1870 2399 1876 2400
rect 1526 2395 1532 2396
rect 1830 2397 1836 2398
rect 110 2392 116 2393
rect 1830 2393 1831 2397
rect 1835 2393 1836 2397
rect 1870 2395 1871 2399
rect 1875 2395 1876 2399
rect 3590 2399 3596 2400
rect 1870 2394 1876 2395
rect 1894 2396 1900 2397
rect 1830 2392 1836 2393
rect 1894 2392 1895 2396
rect 1899 2392 1900 2396
rect 1894 2391 1900 2392
rect 1982 2396 1988 2397
rect 1982 2392 1983 2396
rect 1987 2392 1988 2396
rect 1982 2391 1988 2392
rect 2102 2396 2108 2397
rect 2102 2392 2103 2396
rect 2107 2392 2108 2396
rect 2102 2391 2108 2392
rect 2238 2396 2244 2397
rect 2238 2392 2239 2396
rect 2243 2392 2244 2396
rect 2238 2391 2244 2392
rect 2382 2396 2388 2397
rect 2382 2392 2383 2396
rect 2387 2392 2388 2396
rect 2382 2391 2388 2392
rect 2526 2396 2532 2397
rect 2526 2392 2527 2396
rect 2531 2392 2532 2396
rect 2526 2391 2532 2392
rect 2662 2396 2668 2397
rect 2662 2392 2663 2396
rect 2667 2392 2668 2396
rect 2662 2391 2668 2392
rect 2798 2396 2804 2397
rect 2798 2392 2799 2396
rect 2803 2392 2804 2396
rect 2798 2391 2804 2392
rect 2934 2396 2940 2397
rect 2934 2392 2935 2396
rect 2939 2392 2940 2396
rect 2934 2391 2940 2392
rect 3070 2396 3076 2397
rect 3070 2392 3071 2396
rect 3075 2392 3076 2396
rect 3070 2391 3076 2392
rect 3206 2396 3212 2397
rect 3206 2392 3207 2396
rect 3211 2392 3212 2396
rect 3590 2395 3591 2399
rect 3595 2395 3596 2399
rect 3590 2394 3596 2395
rect 3206 2391 3212 2392
rect 110 2380 116 2381
rect 110 2376 111 2380
rect 115 2376 116 2380
rect 110 2375 116 2376
rect 1830 2380 1836 2381
rect 1830 2376 1831 2380
rect 1835 2376 1836 2380
rect 1830 2375 1836 2376
rect 390 2362 396 2363
rect 390 2358 391 2362
rect 395 2358 396 2362
rect 390 2357 396 2358
rect 470 2362 476 2363
rect 470 2358 471 2362
rect 475 2358 476 2362
rect 470 2357 476 2358
rect 550 2362 556 2363
rect 550 2358 551 2362
rect 555 2358 556 2362
rect 550 2357 556 2358
rect 630 2362 636 2363
rect 630 2358 631 2362
rect 635 2358 636 2362
rect 630 2357 636 2358
rect 710 2362 716 2363
rect 710 2358 711 2362
rect 715 2358 716 2362
rect 710 2357 716 2358
rect 790 2362 796 2363
rect 790 2358 791 2362
rect 795 2358 796 2362
rect 790 2357 796 2358
rect 870 2362 876 2363
rect 870 2358 871 2362
rect 875 2358 876 2362
rect 870 2357 876 2358
rect 950 2362 956 2363
rect 950 2358 951 2362
rect 955 2358 956 2362
rect 950 2357 956 2358
rect 1030 2362 1036 2363
rect 1030 2358 1031 2362
rect 1035 2358 1036 2362
rect 1030 2357 1036 2358
rect 1110 2362 1116 2363
rect 1110 2358 1111 2362
rect 1115 2358 1116 2362
rect 1110 2357 1116 2358
rect 1190 2362 1196 2363
rect 1190 2358 1191 2362
rect 1195 2358 1196 2362
rect 1190 2357 1196 2358
rect 1270 2362 1276 2363
rect 1270 2358 1271 2362
rect 1275 2358 1276 2362
rect 1270 2357 1276 2358
rect 1358 2362 1364 2363
rect 1358 2358 1359 2362
rect 1363 2358 1364 2362
rect 1358 2357 1364 2358
rect 1446 2362 1452 2363
rect 1446 2358 1447 2362
rect 1451 2358 1452 2362
rect 1446 2357 1452 2358
rect 1534 2362 1540 2363
rect 1534 2358 1535 2362
rect 1539 2358 1540 2362
rect 1534 2357 1540 2358
rect 1894 2344 1900 2345
rect 1870 2341 1876 2342
rect 1870 2337 1871 2341
rect 1875 2337 1876 2341
rect 1894 2340 1895 2344
rect 1899 2340 1900 2344
rect 1894 2339 1900 2340
rect 2014 2344 2020 2345
rect 2014 2340 2015 2344
rect 2019 2340 2020 2344
rect 2014 2339 2020 2340
rect 2174 2344 2180 2345
rect 2174 2340 2175 2344
rect 2179 2340 2180 2344
rect 2174 2339 2180 2340
rect 2342 2344 2348 2345
rect 2342 2340 2343 2344
rect 2347 2340 2348 2344
rect 2342 2339 2348 2340
rect 2510 2344 2516 2345
rect 2510 2340 2511 2344
rect 2515 2340 2516 2344
rect 2510 2339 2516 2340
rect 2670 2344 2676 2345
rect 2670 2340 2671 2344
rect 2675 2340 2676 2344
rect 2670 2339 2676 2340
rect 2822 2344 2828 2345
rect 2822 2340 2823 2344
rect 2827 2340 2828 2344
rect 2822 2339 2828 2340
rect 2958 2344 2964 2345
rect 2958 2340 2959 2344
rect 2963 2340 2964 2344
rect 2958 2339 2964 2340
rect 3078 2344 3084 2345
rect 3078 2340 3079 2344
rect 3083 2340 3084 2344
rect 3078 2339 3084 2340
rect 3190 2344 3196 2345
rect 3190 2340 3191 2344
rect 3195 2340 3196 2344
rect 3190 2339 3196 2340
rect 3302 2344 3308 2345
rect 3302 2340 3303 2344
rect 3307 2340 3308 2344
rect 3302 2339 3308 2340
rect 3414 2344 3420 2345
rect 3414 2340 3415 2344
rect 3419 2340 3420 2344
rect 3414 2339 3420 2340
rect 3502 2344 3508 2345
rect 3502 2340 3503 2344
rect 3507 2340 3508 2344
rect 3502 2339 3508 2340
rect 3590 2341 3596 2342
rect 1870 2336 1876 2337
rect 3590 2337 3591 2341
rect 3595 2337 3596 2341
rect 3590 2336 3596 2337
rect 1406 2330 1412 2331
rect 1406 2326 1407 2330
rect 1411 2326 1412 2330
rect 1406 2325 1412 2326
rect 1486 2330 1492 2331
rect 1486 2326 1487 2330
rect 1491 2326 1492 2330
rect 1486 2325 1492 2326
rect 1566 2330 1572 2331
rect 1566 2326 1567 2330
rect 1571 2326 1572 2330
rect 1566 2325 1572 2326
rect 1646 2330 1652 2331
rect 1646 2326 1647 2330
rect 1651 2326 1652 2330
rect 1646 2325 1652 2326
rect 1870 2324 1876 2325
rect 1870 2320 1871 2324
rect 1875 2320 1876 2324
rect 1870 2319 1876 2320
rect 3590 2324 3596 2325
rect 3590 2320 3591 2324
rect 3595 2320 3596 2324
rect 3590 2319 3596 2320
rect 110 2312 116 2313
rect 110 2308 111 2312
rect 115 2308 116 2312
rect 110 2307 116 2308
rect 1830 2312 1836 2313
rect 1830 2308 1831 2312
rect 1835 2308 1836 2312
rect 1830 2307 1836 2308
rect 1902 2306 1908 2307
rect 1902 2302 1903 2306
rect 1907 2302 1908 2306
rect 1902 2301 1908 2302
rect 2022 2306 2028 2307
rect 2022 2302 2023 2306
rect 2027 2302 2028 2306
rect 2022 2301 2028 2302
rect 2182 2306 2188 2307
rect 2182 2302 2183 2306
rect 2187 2302 2188 2306
rect 2182 2301 2188 2302
rect 2350 2306 2356 2307
rect 2350 2302 2351 2306
rect 2355 2302 2356 2306
rect 2350 2301 2356 2302
rect 2518 2306 2524 2307
rect 2518 2302 2519 2306
rect 2523 2302 2524 2306
rect 2518 2301 2524 2302
rect 2678 2306 2684 2307
rect 2678 2302 2679 2306
rect 2683 2302 2684 2306
rect 2678 2301 2684 2302
rect 2830 2306 2836 2307
rect 2830 2302 2831 2306
rect 2835 2302 2836 2306
rect 2830 2301 2836 2302
rect 2966 2306 2972 2307
rect 2966 2302 2967 2306
rect 2971 2302 2972 2306
rect 2966 2301 2972 2302
rect 3086 2306 3092 2307
rect 3086 2302 3087 2306
rect 3091 2302 3092 2306
rect 3086 2301 3092 2302
rect 3198 2306 3204 2307
rect 3198 2302 3199 2306
rect 3203 2302 3204 2306
rect 3198 2301 3204 2302
rect 3310 2306 3316 2307
rect 3310 2302 3311 2306
rect 3315 2302 3316 2306
rect 3310 2301 3316 2302
rect 3422 2306 3428 2307
rect 3422 2302 3423 2306
rect 3427 2302 3428 2306
rect 3422 2301 3428 2302
rect 3510 2306 3516 2307
rect 3510 2302 3511 2306
rect 3515 2302 3516 2306
rect 3510 2301 3516 2302
rect 110 2295 116 2296
rect 110 2291 111 2295
rect 115 2291 116 2295
rect 1830 2295 1836 2296
rect 110 2290 116 2291
rect 1398 2292 1404 2293
rect 1398 2288 1399 2292
rect 1403 2288 1404 2292
rect 1398 2287 1404 2288
rect 1478 2292 1484 2293
rect 1478 2288 1479 2292
rect 1483 2288 1484 2292
rect 1478 2287 1484 2288
rect 1558 2292 1564 2293
rect 1558 2288 1559 2292
rect 1563 2288 1564 2292
rect 1558 2287 1564 2288
rect 1638 2292 1644 2293
rect 1638 2288 1639 2292
rect 1643 2288 1644 2292
rect 1830 2291 1831 2295
rect 1835 2291 1836 2295
rect 1830 2290 1836 2291
rect 1638 2287 1644 2288
rect 1902 2274 1908 2275
rect 1902 2270 1903 2274
rect 1907 2270 1908 2274
rect 1902 2269 1908 2270
rect 2030 2274 2036 2275
rect 2030 2270 2031 2274
rect 2035 2270 2036 2274
rect 2030 2269 2036 2270
rect 2182 2274 2188 2275
rect 2182 2270 2183 2274
rect 2187 2270 2188 2274
rect 2182 2269 2188 2270
rect 2366 2274 2372 2275
rect 2366 2270 2367 2274
rect 2371 2270 2372 2274
rect 2366 2269 2372 2270
rect 2574 2274 2580 2275
rect 2574 2270 2575 2274
rect 2579 2270 2580 2274
rect 2574 2269 2580 2270
rect 2790 2274 2796 2275
rect 2790 2270 2791 2274
rect 2795 2270 2796 2274
rect 2790 2269 2796 2270
rect 3022 2274 3028 2275
rect 3022 2270 3023 2274
rect 3027 2270 3028 2274
rect 3022 2269 3028 2270
rect 3254 2274 3260 2275
rect 3254 2270 3255 2274
rect 3259 2270 3260 2274
rect 3254 2269 3260 2270
rect 3494 2274 3500 2275
rect 3494 2270 3495 2274
rect 3499 2270 3500 2274
rect 3494 2269 3500 2270
rect 1870 2256 1876 2257
rect 1870 2252 1871 2256
rect 1875 2252 1876 2256
rect 1870 2251 1876 2252
rect 3590 2256 3596 2257
rect 3590 2252 3591 2256
rect 3595 2252 3596 2256
rect 3590 2251 3596 2252
rect 134 2240 140 2241
rect 110 2237 116 2238
rect 110 2233 111 2237
rect 115 2233 116 2237
rect 134 2236 135 2240
rect 139 2236 140 2240
rect 134 2235 140 2236
rect 214 2240 220 2241
rect 214 2236 215 2240
rect 219 2236 220 2240
rect 214 2235 220 2236
rect 294 2240 300 2241
rect 294 2236 295 2240
rect 299 2236 300 2240
rect 294 2235 300 2236
rect 382 2240 388 2241
rect 382 2236 383 2240
rect 387 2236 388 2240
rect 382 2235 388 2236
rect 518 2240 524 2241
rect 518 2236 519 2240
rect 523 2236 524 2240
rect 518 2235 524 2236
rect 670 2240 676 2241
rect 670 2236 671 2240
rect 675 2236 676 2240
rect 670 2235 676 2236
rect 830 2240 836 2241
rect 830 2236 831 2240
rect 835 2236 836 2240
rect 830 2235 836 2236
rect 998 2240 1004 2241
rect 998 2236 999 2240
rect 1003 2236 1004 2240
rect 998 2235 1004 2236
rect 1158 2240 1164 2241
rect 1158 2236 1159 2240
rect 1163 2236 1164 2240
rect 1158 2235 1164 2236
rect 1310 2240 1316 2241
rect 1310 2236 1311 2240
rect 1315 2236 1316 2240
rect 1310 2235 1316 2236
rect 1454 2240 1460 2241
rect 1454 2236 1455 2240
rect 1459 2236 1460 2240
rect 1454 2235 1460 2236
rect 1606 2240 1612 2241
rect 1606 2236 1607 2240
rect 1611 2236 1612 2240
rect 1606 2235 1612 2236
rect 1742 2240 1748 2241
rect 1742 2236 1743 2240
rect 1747 2236 1748 2240
rect 1870 2239 1876 2240
rect 1742 2235 1748 2236
rect 1830 2237 1836 2238
rect 110 2232 116 2233
rect 1830 2233 1831 2237
rect 1835 2233 1836 2237
rect 1870 2235 1871 2239
rect 1875 2235 1876 2239
rect 3590 2239 3596 2240
rect 1870 2234 1876 2235
rect 1894 2236 1900 2237
rect 1830 2232 1836 2233
rect 1894 2232 1895 2236
rect 1899 2232 1900 2236
rect 1894 2231 1900 2232
rect 2022 2236 2028 2237
rect 2022 2232 2023 2236
rect 2027 2232 2028 2236
rect 2022 2231 2028 2232
rect 2174 2236 2180 2237
rect 2174 2232 2175 2236
rect 2179 2232 2180 2236
rect 2174 2231 2180 2232
rect 2358 2236 2364 2237
rect 2358 2232 2359 2236
rect 2363 2232 2364 2236
rect 2358 2231 2364 2232
rect 2566 2236 2572 2237
rect 2566 2232 2567 2236
rect 2571 2232 2572 2236
rect 2566 2231 2572 2232
rect 2782 2236 2788 2237
rect 2782 2232 2783 2236
rect 2787 2232 2788 2236
rect 2782 2231 2788 2232
rect 3014 2236 3020 2237
rect 3014 2232 3015 2236
rect 3019 2232 3020 2236
rect 3014 2231 3020 2232
rect 3246 2236 3252 2237
rect 3246 2232 3247 2236
rect 3251 2232 3252 2236
rect 3246 2231 3252 2232
rect 3486 2236 3492 2237
rect 3486 2232 3487 2236
rect 3491 2232 3492 2236
rect 3590 2235 3591 2239
rect 3595 2235 3596 2239
rect 3590 2234 3596 2235
rect 3486 2231 3492 2232
rect 110 2220 116 2221
rect 110 2216 111 2220
rect 115 2216 116 2220
rect 110 2215 116 2216
rect 1830 2220 1836 2221
rect 1830 2216 1831 2220
rect 1835 2216 1836 2220
rect 1830 2215 1836 2216
rect 142 2202 148 2203
rect 142 2198 143 2202
rect 147 2198 148 2202
rect 142 2197 148 2198
rect 222 2202 228 2203
rect 222 2198 223 2202
rect 227 2198 228 2202
rect 222 2197 228 2198
rect 302 2202 308 2203
rect 302 2198 303 2202
rect 307 2198 308 2202
rect 302 2197 308 2198
rect 390 2202 396 2203
rect 390 2198 391 2202
rect 395 2198 396 2202
rect 390 2197 396 2198
rect 526 2202 532 2203
rect 526 2198 527 2202
rect 531 2198 532 2202
rect 526 2197 532 2198
rect 678 2202 684 2203
rect 678 2198 679 2202
rect 683 2198 684 2202
rect 678 2197 684 2198
rect 838 2202 844 2203
rect 838 2198 839 2202
rect 843 2198 844 2202
rect 838 2197 844 2198
rect 1006 2202 1012 2203
rect 1006 2198 1007 2202
rect 1011 2198 1012 2202
rect 1006 2197 1012 2198
rect 1166 2202 1172 2203
rect 1166 2198 1167 2202
rect 1171 2198 1172 2202
rect 1166 2197 1172 2198
rect 1318 2202 1324 2203
rect 1318 2198 1319 2202
rect 1323 2198 1324 2202
rect 1318 2197 1324 2198
rect 1462 2202 1468 2203
rect 1462 2198 1463 2202
rect 1467 2198 1468 2202
rect 1462 2197 1468 2198
rect 1614 2202 1620 2203
rect 1614 2198 1615 2202
rect 1619 2198 1620 2202
rect 1614 2197 1620 2198
rect 1750 2202 1756 2203
rect 1750 2198 1751 2202
rect 1755 2198 1756 2202
rect 1750 2197 1756 2198
rect 2198 2172 2204 2173
rect 1870 2169 1876 2170
rect 190 2166 196 2167
rect 190 2162 191 2166
rect 195 2162 196 2166
rect 190 2161 196 2162
rect 310 2166 316 2167
rect 310 2162 311 2166
rect 315 2162 316 2166
rect 310 2161 316 2162
rect 462 2166 468 2167
rect 462 2162 463 2166
rect 467 2162 468 2166
rect 462 2161 468 2162
rect 638 2166 644 2167
rect 638 2162 639 2166
rect 643 2162 644 2166
rect 638 2161 644 2162
rect 822 2166 828 2167
rect 822 2162 823 2166
rect 827 2162 828 2166
rect 822 2161 828 2162
rect 1014 2166 1020 2167
rect 1014 2162 1015 2166
rect 1019 2162 1020 2166
rect 1014 2161 1020 2162
rect 1198 2166 1204 2167
rect 1198 2162 1199 2166
rect 1203 2162 1204 2166
rect 1198 2161 1204 2162
rect 1390 2166 1396 2167
rect 1390 2162 1391 2166
rect 1395 2162 1396 2166
rect 1390 2161 1396 2162
rect 1582 2166 1588 2167
rect 1582 2162 1583 2166
rect 1587 2162 1588 2166
rect 1582 2161 1588 2162
rect 1750 2166 1756 2167
rect 1750 2162 1751 2166
rect 1755 2162 1756 2166
rect 1870 2165 1871 2169
rect 1875 2165 1876 2169
rect 2198 2168 2199 2172
rect 2203 2168 2204 2172
rect 2198 2167 2204 2168
rect 2294 2172 2300 2173
rect 2294 2168 2295 2172
rect 2299 2168 2300 2172
rect 2294 2167 2300 2168
rect 2398 2172 2404 2173
rect 2398 2168 2399 2172
rect 2403 2168 2404 2172
rect 2398 2167 2404 2168
rect 2518 2172 2524 2173
rect 2518 2168 2519 2172
rect 2523 2168 2524 2172
rect 2518 2167 2524 2168
rect 2638 2172 2644 2173
rect 2638 2168 2639 2172
rect 2643 2168 2644 2172
rect 2638 2167 2644 2168
rect 2758 2172 2764 2173
rect 2758 2168 2759 2172
rect 2763 2168 2764 2172
rect 2758 2167 2764 2168
rect 2878 2172 2884 2173
rect 2878 2168 2879 2172
rect 2883 2168 2884 2172
rect 2878 2167 2884 2168
rect 2990 2172 2996 2173
rect 2990 2168 2991 2172
rect 2995 2168 2996 2172
rect 2990 2167 2996 2168
rect 3094 2172 3100 2173
rect 3094 2168 3095 2172
rect 3099 2168 3100 2172
rect 3094 2167 3100 2168
rect 3198 2172 3204 2173
rect 3198 2168 3199 2172
rect 3203 2168 3204 2172
rect 3198 2167 3204 2168
rect 3302 2172 3308 2173
rect 3302 2168 3303 2172
rect 3307 2168 3308 2172
rect 3302 2167 3308 2168
rect 3406 2172 3412 2173
rect 3406 2168 3407 2172
rect 3411 2168 3412 2172
rect 3406 2167 3412 2168
rect 3502 2172 3508 2173
rect 3502 2168 3503 2172
rect 3507 2168 3508 2172
rect 3502 2167 3508 2168
rect 3590 2169 3596 2170
rect 1870 2164 1876 2165
rect 3590 2165 3591 2169
rect 3595 2165 3596 2169
rect 3590 2164 3596 2165
rect 1750 2161 1756 2162
rect 1870 2152 1876 2153
rect 110 2148 116 2149
rect 110 2144 111 2148
rect 115 2144 116 2148
rect 110 2143 116 2144
rect 1830 2148 1836 2149
rect 1830 2144 1831 2148
rect 1835 2144 1836 2148
rect 1870 2148 1871 2152
rect 1875 2148 1876 2152
rect 1870 2147 1876 2148
rect 3590 2152 3596 2153
rect 3590 2148 3591 2152
rect 3595 2148 3596 2152
rect 3590 2147 3596 2148
rect 1830 2143 1836 2144
rect 2206 2134 2212 2135
rect 110 2131 116 2132
rect 110 2127 111 2131
rect 115 2127 116 2131
rect 1830 2131 1836 2132
rect 110 2126 116 2127
rect 182 2128 188 2129
rect 182 2124 183 2128
rect 187 2124 188 2128
rect 182 2123 188 2124
rect 302 2128 308 2129
rect 302 2124 303 2128
rect 307 2124 308 2128
rect 302 2123 308 2124
rect 454 2128 460 2129
rect 454 2124 455 2128
rect 459 2124 460 2128
rect 454 2123 460 2124
rect 630 2128 636 2129
rect 630 2124 631 2128
rect 635 2124 636 2128
rect 630 2123 636 2124
rect 814 2128 820 2129
rect 814 2124 815 2128
rect 819 2124 820 2128
rect 814 2123 820 2124
rect 1006 2128 1012 2129
rect 1006 2124 1007 2128
rect 1011 2124 1012 2128
rect 1006 2123 1012 2124
rect 1190 2128 1196 2129
rect 1190 2124 1191 2128
rect 1195 2124 1196 2128
rect 1190 2123 1196 2124
rect 1382 2128 1388 2129
rect 1382 2124 1383 2128
rect 1387 2124 1388 2128
rect 1382 2123 1388 2124
rect 1574 2128 1580 2129
rect 1574 2124 1575 2128
rect 1579 2124 1580 2128
rect 1574 2123 1580 2124
rect 1742 2128 1748 2129
rect 1742 2124 1743 2128
rect 1747 2124 1748 2128
rect 1830 2127 1831 2131
rect 1835 2127 1836 2131
rect 2206 2130 2207 2134
rect 2211 2130 2212 2134
rect 2206 2129 2212 2130
rect 2302 2134 2308 2135
rect 2302 2130 2303 2134
rect 2307 2130 2308 2134
rect 2302 2129 2308 2130
rect 2406 2134 2412 2135
rect 2406 2130 2407 2134
rect 2411 2130 2412 2134
rect 2406 2129 2412 2130
rect 2526 2134 2532 2135
rect 2526 2130 2527 2134
rect 2531 2130 2532 2134
rect 2526 2129 2532 2130
rect 2646 2134 2652 2135
rect 2646 2130 2647 2134
rect 2651 2130 2652 2134
rect 2646 2129 2652 2130
rect 2766 2134 2772 2135
rect 2766 2130 2767 2134
rect 2771 2130 2772 2134
rect 2766 2129 2772 2130
rect 2886 2134 2892 2135
rect 2886 2130 2887 2134
rect 2891 2130 2892 2134
rect 2886 2129 2892 2130
rect 2998 2134 3004 2135
rect 2998 2130 2999 2134
rect 3003 2130 3004 2134
rect 2998 2129 3004 2130
rect 3102 2134 3108 2135
rect 3102 2130 3103 2134
rect 3107 2130 3108 2134
rect 3102 2129 3108 2130
rect 3206 2134 3212 2135
rect 3206 2130 3207 2134
rect 3211 2130 3212 2134
rect 3206 2129 3212 2130
rect 3310 2134 3316 2135
rect 3310 2130 3311 2134
rect 3315 2130 3316 2134
rect 3310 2129 3316 2130
rect 3414 2134 3420 2135
rect 3414 2130 3415 2134
rect 3419 2130 3420 2134
rect 3414 2129 3420 2130
rect 3510 2134 3516 2135
rect 3510 2130 3511 2134
rect 3515 2130 3516 2134
rect 3510 2129 3516 2130
rect 1830 2126 1836 2127
rect 1742 2123 1748 2124
rect 2174 2090 2180 2091
rect 2174 2086 2175 2090
rect 2179 2086 2180 2090
rect 2174 2085 2180 2086
rect 2270 2090 2276 2091
rect 2270 2086 2271 2090
rect 2275 2086 2276 2090
rect 2270 2085 2276 2086
rect 2374 2090 2380 2091
rect 2374 2086 2375 2090
rect 2379 2086 2380 2090
rect 2374 2085 2380 2086
rect 2486 2090 2492 2091
rect 2486 2086 2487 2090
rect 2491 2086 2492 2090
rect 2486 2085 2492 2086
rect 2606 2090 2612 2091
rect 2606 2086 2607 2090
rect 2611 2086 2612 2090
rect 2606 2085 2612 2086
rect 2726 2090 2732 2091
rect 2726 2086 2727 2090
rect 2731 2086 2732 2090
rect 2726 2085 2732 2086
rect 2846 2090 2852 2091
rect 2846 2086 2847 2090
rect 2851 2086 2852 2090
rect 2846 2085 2852 2086
rect 2966 2090 2972 2091
rect 2966 2086 2967 2090
rect 2971 2086 2972 2090
rect 2966 2085 2972 2086
rect 3078 2090 3084 2091
rect 3078 2086 3079 2090
rect 3083 2086 3084 2090
rect 3078 2085 3084 2086
rect 3190 2090 3196 2091
rect 3190 2086 3191 2090
rect 3195 2086 3196 2090
rect 3190 2085 3196 2086
rect 3302 2090 3308 2091
rect 3302 2086 3303 2090
rect 3307 2086 3308 2090
rect 3302 2085 3308 2086
rect 3414 2090 3420 2091
rect 3414 2086 3415 2090
rect 3419 2086 3420 2090
rect 3414 2085 3420 2086
rect 3510 2090 3516 2091
rect 3510 2086 3511 2090
rect 3515 2086 3516 2090
rect 3510 2085 3516 2086
rect 214 2080 220 2081
rect 110 2077 116 2078
rect 110 2073 111 2077
rect 115 2073 116 2077
rect 214 2076 215 2080
rect 219 2076 220 2080
rect 214 2075 220 2076
rect 358 2080 364 2081
rect 358 2076 359 2080
rect 363 2076 364 2080
rect 358 2075 364 2076
rect 518 2080 524 2081
rect 518 2076 519 2080
rect 523 2076 524 2080
rect 518 2075 524 2076
rect 702 2080 708 2081
rect 702 2076 703 2080
rect 707 2076 708 2080
rect 702 2075 708 2076
rect 894 2080 900 2081
rect 894 2076 895 2080
rect 899 2076 900 2080
rect 894 2075 900 2076
rect 1102 2080 1108 2081
rect 1102 2076 1103 2080
rect 1107 2076 1108 2080
rect 1102 2075 1108 2076
rect 1310 2080 1316 2081
rect 1310 2076 1311 2080
rect 1315 2076 1316 2080
rect 1310 2075 1316 2076
rect 1526 2080 1532 2081
rect 1526 2076 1527 2080
rect 1531 2076 1532 2080
rect 1526 2075 1532 2076
rect 1742 2080 1748 2081
rect 1742 2076 1743 2080
rect 1747 2076 1748 2080
rect 1742 2075 1748 2076
rect 1830 2077 1836 2078
rect 110 2072 116 2073
rect 1830 2073 1831 2077
rect 1835 2073 1836 2077
rect 1830 2072 1836 2073
rect 1870 2072 1876 2073
rect 1870 2068 1871 2072
rect 1875 2068 1876 2072
rect 1870 2067 1876 2068
rect 3590 2072 3596 2073
rect 3590 2068 3591 2072
rect 3595 2068 3596 2072
rect 3590 2067 3596 2068
rect 110 2060 116 2061
rect 110 2056 111 2060
rect 115 2056 116 2060
rect 110 2055 116 2056
rect 1830 2060 1836 2061
rect 1830 2056 1831 2060
rect 1835 2056 1836 2060
rect 1830 2055 1836 2056
rect 1870 2055 1876 2056
rect 1870 2051 1871 2055
rect 1875 2051 1876 2055
rect 3590 2055 3596 2056
rect 1870 2050 1876 2051
rect 2166 2052 2172 2053
rect 2166 2048 2167 2052
rect 2171 2048 2172 2052
rect 2166 2047 2172 2048
rect 2262 2052 2268 2053
rect 2262 2048 2263 2052
rect 2267 2048 2268 2052
rect 2262 2047 2268 2048
rect 2366 2052 2372 2053
rect 2366 2048 2367 2052
rect 2371 2048 2372 2052
rect 2366 2047 2372 2048
rect 2478 2052 2484 2053
rect 2478 2048 2479 2052
rect 2483 2048 2484 2052
rect 2478 2047 2484 2048
rect 2598 2052 2604 2053
rect 2598 2048 2599 2052
rect 2603 2048 2604 2052
rect 2598 2047 2604 2048
rect 2718 2052 2724 2053
rect 2718 2048 2719 2052
rect 2723 2048 2724 2052
rect 2718 2047 2724 2048
rect 2838 2052 2844 2053
rect 2838 2048 2839 2052
rect 2843 2048 2844 2052
rect 2838 2047 2844 2048
rect 2958 2052 2964 2053
rect 2958 2048 2959 2052
rect 2963 2048 2964 2052
rect 2958 2047 2964 2048
rect 3070 2052 3076 2053
rect 3070 2048 3071 2052
rect 3075 2048 3076 2052
rect 3070 2047 3076 2048
rect 3182 2052 3188 2053
rect 3182 2048 3183 2052
rect 3187 2048 3188 2052
rect 3182 2047 3188 2048
rect 3294 2052 3300 2053
rect 3294 2048 3295 2052
rect 3299 2048 3300 2052
rect 3294 2047 3300 2048
rect 3406 2052 3412 2053
rect 3406 2048 3407 2052
rect 3411 2048 3412 2052
rect 3406 2047 3412 2048
rect 3502 2052 3508 2053
rect 3502 2048 3503 2052
rect 3507 2048 3508 2052
rect 3590 2051 3591 2055
rect 3595 2051 3596 2055
rect 3590 2050 3596 2051
rect 3502 2047 3508 2048
rect 222 2042 228 2043
rect 222 2038 223 2042
rect 227 2038 228 2042
rect 222 2037 228 2038
rect 366 2042 372 2043
rect 366 2038 367 2042
rect 371 2038 372 2042
rect 366 2037 372 2038
rect 526 2042 532 2043
rect 526 2038 527 2042
rect 531 2038 532 2042
rect 526 2037 532 2038
rect 710 2042 716 2043
rect 710 2038 711 2042
rect 715 2038 716 2042
rect 710 2037 716 2038
rect 902 2042 908 2043
rect 902 2038 903 2042
rect 907 2038 908 2042
rect 902 2037 908 2038
rect 1110 2042 1116 2043
rect 1110 2038 1111 2042
rect 1115 2038 1116 2042
rect 1110 2037 1116 2038
rect 1318 2042 1324 2043
rect 1318 2038 1319 2042
rect 1323 2038 1324 2042
rect 1318 2037 1324 2038
rect 1534 2042 1540 2043
rect 1534 2038 1535 2042
rect 1539 2038 1540 2042
rect 1534 2037 1540 2038
rect 1750 2042 1756 2043
rect 1750 2038 1751 2042
rect 1755 2038 1756 2042
rect 1750 2037 1756 2038
rect 142 2010 148 2011
rect 142 2006 143 2010
rect 147 2006 148 2010
rect 142 2005 148 2006
rect 262 2010 268 2011
rect 262 2006 263 2010
rect 267 2006 268 2010
rect 262 2005 268 2006
rect 382 2010 388 2011
rect 382 2006 383 2010
rect 387 2006 388 2010
rect 382 2005 388 2006
rect 494 2010 500 2011
rect 494 2006 495 2010
rect 499 2006 500 2010
rect 494 2005 500 2006
rect 606 2010 612 2011
rect 606 2006 607 2010
rect 611 2006 612 2010
rect 606 2005 612 2006
rect 718 2010 724 2011
rect 718 2006 719 2010
rect 723 2006 724 2010
rect 718 2005 724 2006
rect 822 2010 828 2011
rect 822 2006 823 2010
rect 827 2006 828 2010
rect 822 2005 828 2006
rect 926 2010 932 2011
rect 926 2006 927 2010
rect 931 2006 932 2010
rect 926 2005 932 2006
rect 1022 2010 1028 2011
rect 1022 2006 1023 2010
rect 1027 2006 1028 2010
rect 1022 2005 1028 2006
rect 1110 2010 1116 2011
rect 1110 2006 1111 2010
rect 1115 2006 1116 2010
rect 1110 2005 1116 2006
rect 1206 2010 1212 2011
rect 1206 2006 1207 2010
rect 1211 2006 1212 2010
rect 1206 2005 1212 2006
rect 1294 2010 1300 2011
rect 1294 2006 1295 2010
rect 1299 2006 1300 2010
rect 1294 2005 1300 2006
rect 1390 2010 1396 2011
rect 1390 2006 1391 2010
rect 1395 2006 1396 2010
rect 1390 2005 1396 2006
rect 1486 2010 1492 2011
rect 1486 2006 1487 2010
rect 1491 2006 1492 2010
rect 1486 2005 1492 2006
rect 1582 2010 1588 2011
rect 1582 2006 1583 2010
rect 1587 2006 1588 2010
rect 1582 2005 1588 2006
rect 1670 2010 1676 2011
rect 1670 2006 1671 2010
rect 1675 2006 1676 2010
rect 1670 2005 1676 2006
rect 1750 2010 1756 2011
rect 1750 2006 1751 2010
rect 1755 2006 1756 2010
rect 1750 2005 1756 2006
rect 2070 2004 2076 2005
rect 1870 2001 1876 2002
rect 1870 1997 1871 2001
rect 1875 1997 1876 2001
rect 2070 2000 2071 2004
rect 2075 2000 2076 2004
rect 2070 1999 2076 2000
rect 2206 2004 2212 2005
rect 2206 2000 2207 2004
rect 2211 2000 2212 2004
rect 2206 1999 2212 2000
rect 2358 2004 2364 2005
rect 2358 2000 2359 2004
rect 2363 2000 2364 2004
rect 2358 1999 2364 2000
rect 2518 2004 2524 2005
rect 2518 2000 2519 2004
rect 2523 2000 2524 2004
rect 2518 1999 2524 2000
rect 2678 2004 2684 2005
rect 2678 2000 2679 2004
rect 2683 2000 2684 2004
rect 2678 1999 2684 2000
rect 2846 2004 2852 2005
rect 2846 2000 2847 2004
rect 2851 2000 2852 2004
rect 2846 1999 2852 2000
rect 3014 2004 3020 2005
rect 3014 2000 3015 2004
rect 3019 2000 3020 2004
rect 3014 1999 3020 2000
rect 3182 2004 3188 2005
rect 3182 2000 3183 2004
rect 3187 2000 3188 2004
rect 3182 1999 3188 2000
rect 3350 2004 3356 2005
rect 3350 2000 3351 2004
rect 3355 2000 3356 2004
rect 3350 1999 3356 2000
rect 3502 2004 3508 2005
rect 3502 2000 3503 2004
rect 3507 2000 3508 2004
rect 3502 1999 3508 2000
rect 3590 2001 3596 2002
rect 1870 1996 1876 1997
rect 3590 1997 3591 2001
rect 3595 1997 3596 2001
rect 3590 1996 3596 1997
rect 110 1992 116 1993
rect 110 1988 111 1992
rect 115 1988 116 1992
rect 110 1987 116 1988
rect 1830 1992 1836 1993
rect 1830 1988 1831 1992
rect 1835 1988 1836 1992
rect 1830 1987 1836 1988
rect 1870 1984 1876 1985
rect 1870 1980 1871 1984
rect 1875 1980 1876 1984
rect 1870 1979 1876 1980
rect 3590 1984 3596 1985
rect 3590 1980 3591 1984
rect 3595 1980 3596 1984
rect 3590 1979 3596 1980
rect 110 1975 116 1976
rect 110 1971 111 1975
rect 115 1971 116 1975
rect 1830 1975 1836 1976
rect 110 1970 116 1971
rect 134 1972 140 1973
rect 134 1968 135 1972
rect 139 1968 140 1972
rect 134 1967 140 1968
rect 254 1972 260 1973
rect 254 1968 255 1972
rect 259 1968 260 1972
rect 254 1967 260 1968
rect 374 1972 380 1973
rect 374 1968 375 1972
rect 379 1968 380 1972
rect 374 1967 380 1968
rect 486 1972 492 1973
rect 486 1968 487 1972
rect 491 1968 492 1972
rect 486 1967 492 1968
rect 598 1972 604 1973
rect 598 1968 599 1972
rect 603 1968 604 1972
rect 598 1967 604 1968
rect 710 1972 716 1973
rect 710 1968 711 1972
rect 715 1968 716 1972
rect 710 1967 716 1968
rect 814 1972 820 1973
rect 814 1968 815 1972
rect 819 1968 820 1972
rect 814 1967 820 1968
rect 918 1972 924 1973
rect 918 1968 919 1972
rect 923 1968 924 1972
rect 918 1967 924 1968
rect 1014 1972 1020 1973
rect 1014 1968 1015 1972
rect 1019 1968 1020 1972
rect 1014 1967 1020 1968
rect 1102 1972 1108 1973
rect 1102 1968 1103 1972
rect 1107 1968 1108 1972
rect 1102 1967 1108 1968
rect 1198 1972 1204 1973
rect 1198 1968 1199 1972
rect 1203 1968 1204 1972
rect 1198 1967 1204 1968
rect 1286 1972 1292 1973
rect 1286 1968 1287 1972
rect 1291 1968 1292 1972
rect 1286 1967 1292 1968
rect 1382 1972 1388 1973
rect 1382 1968 1383 1972
rect 1387 1968 1388 1972
rect 1382 1967 1388 1968
rect 1478 1972 1484 1973
rect 1478 1968 1479 1972
rect 1483 1968 1484 1972
rect 1478 1967 1484 1968
rect 1574 1972 1580 1973
rect 1574 1968 1575 1972
rect 1579 1968 1580 1972
rect 1574 1967 1580 1968
rect 1662 1972 1668 1973
rect 1662 1968 1663 1972
rect 1667 1968 1668 1972
rect 1662 1967 1668 1968
rect 1742 1972 1748 1973
rect 1742 1968 1743 1972
rect 1747 1968 1748 1972
rect 1830 1971 1831 1975
rect 1835 1971 1836 1975
rect 1830 1970 1836 1971
rect 1742 1967 1748 1968
rect 2078 1966 2084 1967
rect 2078 1962 2079 1966
rect 2083 1962 2084 1966
rect 2078 1961 2084 1962
rect 2214 1966 2220 1967
rect 2214 1962 2215 1966
rect 2219 1962 2220 1966
rect 2214 1961 2220 1962
rect 2366 1966 2372 1967
rect 2366 1962 2367 1966
rect 2371 1962 2372 1966
rect 2366 1961 2372 1962
rect 2526 1966 2532 1967
rect 2526 1962 2527 1966
rect 2531 1962 2532 1966
rect 2526 1961 2532 1962
rect 2686 1966 2692 1967
rect 2686 1962 2687 1966
rect 2691 1962 2692 1966
rect 2686 1961 2692 1962
rect 2854 1966 2860 1967
rect 2854 1962 2855 1966
rect 2859 1962 2860 1966
rect 2854 1961 2860 1962
rect 3022 1966 3028 1967
rect 3022 1962 3023 1966
rect 3027 1962 3028 1966
rect 3022 1961 3028 1962
rect 3190 1966 3196 1967
rect 3190 1962 3191 1966
rect 3195 1962 3196 1966
rect 3190 1961 3196 1962
rect 3358 1966 3364 1967
rect 3358 1962 3359 1966
rect 3363 1962 3364 1966
rect 3358 1961 3364 1962
rect 3510 1966 3516 1967
rect 3510 1962 3511 1966
rect 3515 1962 3516 1966
rect 3510 1961 3516 1962
rect 1902 1934 1908 1935
rect 1902 1930 1903 1934
rect 1907 1930 1908 1934
rect 1902 1929 1908 1930
rect 2006 1934 2012 1935
rect 2006 1930 2007 1934
rect 2011 1930 2012 1934
rect 2006 1929 2012 1930
rect 2134 1934 2140 1935
rect 2134 1930 2135 1934
rect 2139 1930 2140 1934
rect 2134 1929 2140 1930
rect 2254 1934 2260 1935
rect 2254 1930 2255 1934
rect 2259 1930 2260 1934
rect 2254 1929 2260 1930
rect 2374 1934 2380 1935
rect 2374 1930 2375 1934
rect 2379 1930 2380 1934
rect 2374 1929 2380 1930
rect 2486 1934 2492 1935
rect 2486 1930 2487 1934
rect 2491 1930 2492 1934
rect 2486 1929 2492 1930
rect 2598 1934 2604 1935
rect 2598 1930 2599 1934
rect 2603 1930 2604 1934
rect 2598 1929 2604 1930
rect 2718 1934 2724 1935
rect 2718 1930 2719 1934
rect 2723 1930 2724 1934
rect 2718 1929 2724 1930
rect 2838 1934 2844 1935
rect 2838 1930 2839 1934
rect 2843 1930 2844 1934
rect 2838 1929 2844 1930
rect 166 1920 172 1921
rect 110 1917 116 1918
rect 110 1913 111 1917
rect 115 1913 116 1917
rect 166 1916 167 1920
rect 171 1916 172 1920
rect 166 1915 172 1916
rect 326 1920 332 1921
rect 326 1916 327 1920
rect 331 1916 332 1920
rect 326 1915 332 1916
rect 486 1920 492 1921
rect 486 1916 487 1920
rect 491 1916 492 1920
rect 486 1915 492 1916
rect 646 1920 652 1921
rect 646 1916 647 1920
rect 651 1916 652 1920
rect 646 1915 652 1916
rect 798 1920 804 1921
rect 798 1916 799 1920
rect 803 1916 804 1920
rect 798 1915 804 1916
rect 942 1920 948 1921
rect 942 1916 943 1920
rect 947 1916 948 1920
rect 942 1915 948 1916
rect 1078 1920 1084 1921
rect 1078 1916 1079 1920
rect 1083 1916 1084 1920
rect 1078 1915 1084 1916
rect 1214 1920 1220 1921
rect 1214 1916 1215 1920
rect 1219 1916 1220 1920
rect 1214 1915 1220 1916
rect 1350 1920 1356 1921
rect 1350 1916 1351 1920
rect 1355 1916 1356 1920
rect 1350 1915 1356 1916
rect 1486 1920 1492 1921
rect 1486 1916 1487 1920
rect 1491 1916 1492 1920
rect 1486 1915 1492 1916
rect 1622 1920 1628 1921
rect 1622 1916 1623 1920
rect 1627 1916 1628 1920
rect 1622 1915 1628 1916
rect 1742 1920 1748 1921
rect 1742 1916 1743 1920
rect 1747 1916 1748 1920
rect 1742 1915 1748 1916
rect 1830 1917 1836 1918
rect 110 1912 116 1913
rect 1830 1913 1831 1917
rect 1835 1913 1836 1917
rect 1830 1912 1836 1913
rect 1870 1916 1876 1917
rect 1870 1912 1871 1916
rect 1875 1912 1876 1916
rect 1870 1911 1876 1912
rect 3590 1916 3596 1917
rect 3590 1912 3591 1916
rect 3595 1912 3596 1916
rect 3590 1911 3596 1912
rect 110 1900 116 1901
rect 110 1896 111 1900
rect 115 1896 116 1900
rect 110 1895 116 1896
rect 1830 1900 1836 1901
rect 1830 1896 1831 1900
rect 1835 1896 1836 1900
rect 1830 1895 1836 1896
rect 1870 1899 1876 1900
rect 1870 1895 1871 1899
rect 1875 1895 1876 1899
rect 3590 1899 3596 1900
rect 1870 1894 1876 1895
rect 1894 1896 1900 1897
rect 1894 1892 1895 1896
rect 1899 1892 1900 1896
rect 1894 1891 1900 1892
rect 1998 1896 2004 1897
rect 1998 1892 1999 1896
rect 2003 1892 2004 1896
rect 1998 1891 2004 1892
rect 2126 1896 2132 1897
rect 2126 1892 2127 1896
rect 2131 1892 2132 1896
rect 2126 1891 2132 1892
rect 2246 1896 2252 1897
rect 2246 1892 2247 1896
rect 2251 1892 2252 1896
rect 2246 1891 2252 1892
rect 2366 1896 2372 1897
rect 2366 1892 2367 1896
rect 2371 1892 2372 1896
rect 2366 1891 2372 1892
rect 2478 1896 2484 1897
rect 2478 1892 2479 1896
rect 2483 1892 2484 1896
rect 2478 1891 2484 1892
rect 2590 1896 2596 1897
rect 2590 1892 2591 1896
rect 2595 1892 2596 1896
rect 2590 1891 2596 1892
rect 2710 1896 2716 1897
rect 2710 1892 2711 1896
rect 2715 1892 2716 1896
rect 2710 1891 2716 1892
rect 2830 1896 2836 1897
rect 2830 1892 2831 1896
rect 2835 1892 2836 1896
rect 3590 1895 3591 1899
rect 3595 1895 3596 1899
rect 3590 1894 3596 1895
rect 2830 1891 2836 1892
rect 174 1882 180 1883
rect 174 1878 175 1882
rect 179 1878 180 1882
rect 174 1877 180 1878
rect 334 1882 340 1883
rect 334 1878 335 1882
rect 339 1878 340 1882
rect 334 1877 340 1878
rect 494 1882 500 1883
rect 494 1878 495 1882
rect 499 1878 500 1882
rect 494 1877 500 1878
rect 654 1882 660 1883
rect 654 1878 655 1882
rect 659 1878 660 1882
rect 654 1877 660 1878
rect 806 1882 812 1883
rect 806 1878 807 1882
rect 811 1878 812 1882
rect 806 1877 812 1878
rect 950 1882 956 1883
rect 950 1878 951 1882
rect 955 1878 956 1882
rect 950 1877 956 1878
rect 1086 1882 1092 1883
rect 1086 1878 1087 1882
rect 1091 1878 1092 1882
rect 1086 1877 1092 1878
rect 1222 1882 1228 1883
rect 1222 1878 1223 1882
rect 1227 1878 1228 1882
rect 1222 1877 1228 1878
rect 1358 1882 1364 1883
rect 1358 1878 1359 1882
rect 1363 1878 1364 1882
rect 1358 1877 1364 1878
rect 1494 1882 1500 1883
rect 1494 1878 1495 1882
rect 1499 1878 1500 1882
rect 1494 1877 1500 1878
rect 1630 1882 1636 1883
rect 1630 1878 1631 1882
rect 1635 1878 1636 1882
rect 1630 1877 1636 1878
rect 1750 1882 1756 1883
rect 1750 1878 1751 1882
rect 1755 1878 1756 1882
rect 1750 1877 1756 1878
rect 1894 1852 1900 1853
rect 158 1850 164 1851
rect 158 1846 159 1850
rect 163 1846 164 1850
rect 158 1845 164 1846
rect 302 1850 308 1851
rect 302 1846 303 1850
rect 307 1846 308 1850
rect 302 1845 308 1846
rect 446 1850 452 1851
rect 446 1846 447 1850
rect 451 1846 452 1850
rect 446 1845 452 1846
rect 598 1850 604 1851
rect 598 1846 599 1850
rect 603 1846 604 1850
rect 598 1845 604 1846
rect 750 1850 756 1851
rect 750 1846 751 1850
rect 755 1846 756 1850
rect 750 1845 756 1846
rect 902 1850 908 1851
rect 902 1846 903 1850
rect 907 1846 908 1850
rect 902 1845 908 1846
rect 1054 1850 1060 1851
rect 1054 1846 1055 1850
rect 1059 1846 1060 1850
rect 1054 1845 1060 1846
rect 1206 1850 1212 1851
rect 1206 1846 1207 1850
rect 1211 1846 1212 1850
rect 1206 1845 1212 1846
rect 1350 1850 1356 1851
rect 1350 1846 1351 1850
rect 1355 1846 1356 1850
rect 1350 1845 1356 1846
rect 1486 1850 1492 1851
rect 1486 1846 1487 1850
rect 1491 1846 1492 1850
rect 1486 1845 1492 1846
rect 1630 1850 1636 1851
rect 1630 1846 1631 1850
rect 1635 1846 1636 1850
rect 1630 1845 1636 1846
rect 1750 1850 1756 1851
rect 1750 1846 1751 1850
rect 1755 1846 1756 1850
rect 1750 1845 1756 1846
rect 1870 1849 1876 1850
rect 1870 1845 1871 1849
rect 1875 1845 1876 1849
rect 1894 1848 1895 1852
rect 1899 1848 1900 1852
rect 1894 1847 1900 1848
rect 1990 1852 1996 1853
rect 1990 1848 1991 1852
rect 1995 1848 1996 1852
rect 1990 1847 1996 1848
rect 2118 1852 2124 1853
rect 2118 1848 2119 1852
rect 2123 1848 2124 1852
rect 2118 1847 2124 1848
rect 2246 1852 2252 1853
rect 2246 1848 2247 1852
rect 2251 1848 2252 1852
rect 2246 1847 2252 1848
rect 2382 1852 2388 1853
rect 2382 1848 2383 1852
rect 2387 1848 2388 1852
rect 2382 1847 2388 1848
rect 2518 1852 2524 1853
rect 2518 1848 2519 1852
rect 2523 1848 2524 1852
rect 2518 1847 2524 1848
rect 2654 1852 2660 1853
rect 2654 1848 2655 1852
rect 2659 1848 2660 1852
rect 2654 1847 2660 1848
rect 2806 1852 2812 1853
rect 2806 1848 2807 1852
rect 2811 1848 2812 1852
rect 2806 1847 2812 1848
rect 2974 1852 2980 1853
rect 2974 1848 2975 1852
rect 2979 1848 2980 1852
rect 2974 1847 2980 1848
rect 3150 1852 3156 1853
rect 3150 1848 3151 1852
rect 3155 1848 3156 1852
rect 3150 1847 3156 1848
rect 3334 1852 3340 1853
rect 3334 1848 3335 1852
rect 3339 1848 3340 1852
rect 3334 1847 3340 1848
rect 3502 1852 3508 1853
rect 3502 1848 3503 1852
rect 3507 1848 3508 1852
rect 3502 1847 3508 1848
rect 3590 1849 3596 1850
rect 1870 1844 1876 1845
rect 3590 1845 3591 1849
rect 3595 1845 3596 1849
rect 3590 1844 3596 1845
rect 110 1832 116 1833
rect 110 1828 111 1832
rect 115 1828 116 1832
rect 110 1827 116 1828
rect 1830 1832 1836 1833
rect 1830 1828 1831 1832
rect 1835 1828 1836 1832
rect 1830 1827 1836 1828
rect 1870 1832 1876 1833
rect 1870 1828 1871 1832
rect 1875 1828 1876 1832
rect 1870 1827 1876 1828
rect 3590 1832 3596 1833
rect 3590 1828 3591 1832
rect 3595 1828 3596 1832
rect 3590 1827 3596 1828
rect 110 1815 116 1816
rect 110 1811 111 1815
rect 115 1811 116 1815
rect 1830 1815 1836 1816
rect 110 1810 116 1811
rect 150 1812 156 1813
rect 150 1808 151 1812
rect 155 1808 156 1812
rect 150 1807 156 1808
rect 294 1812 300 1813
rect 294 1808 295 1812
rect 299 1808 300 1812
rect 294 1807 300 1808
rect 438 1812 444 1813
rect 438 1808 439 1812
rect 443 1808 444 1812
rect 438 1807 444 1808
rect 590 1812 596 1813
rect 590 1808 591 1812
rect 595 1808 596 1812
rect 590 1807 596 1808
rect 742 1812 748 1813
rect 742 1808 743 1812
rect 747 1808 748 1812
rect 742 1807 748 1808
rect 894 1812 900 1813
rect 894 1808 895 1812
rect 899 1808 900 1812
rect 894 1807 900 1808
rect 1046 1812 1052 1813
rect 1046 1808 1047 1812
rect 1051 1808 1052 1812
rect 1046 1807 1052 1808
rect 1198 1812 1204 1813
rect 1198 1808 1199 1812
rect 1203 1808 1204 1812
rect 1198 1807 1204 1808
rect 1342 1812 1348 1813
rect 1342 1808 1343 1812
rect 1347 1808 1348 1812
rect 1342 1807 1348 1808
rect 1478 1812 1484 1813
rect 1478 1808 1479 1812
rect 1483 1808 1484 1812
rect 1478 1807 1484 1808
rect 1622 1812 1628 1813
rect 1622 1808 1623 1812
rect 1627 1808 1628 1812
rect 1622 1807 1628 1808
rect 1742 1812 1748 1813
rect 1742 1808 1743 1812
rect 1747 1808 1748 1812
rect 1830 1811 1831 1815
rect 1835 1811 1836 1815
rect 1830 1810 1836 1811
rect 1902 1814 1908 1815
rect 1902 1810 1903 1814
rect 1907 1810 1908 1814
rect 1902 1809 1908 1810
rect 1998 1814 2004 1815
rect 1998 1810 1999 1814
rect 2003 1810 2004 1814
rect 1998 1809 2004 1810
rect 2126 1814 2132 1815
rect 2126 1810 2127 1814
rect 2131 1810 2132 1814
rect 2126 1809 2132 1810
rect 2254 1814 2260 1815
rect 2254 1810 2255 1814
rect 2259 1810 2260 1814
rect 2254 1809 2260 1810
rect 2390 1814 2396 1815
rect 2390 1810 2391 1814
rect 2395 1810 2396 1814
rect 2390 1809 2396 1810
rect 2526 1814 2532 1815
rect 2526 1810 2527 1814
rect 2531 1810 2532 1814
rect 2526 1809 2532 1810
rect 2662 1814 2668 1815
rect 2662 1810 2663 1814
rect 2667 1810 2668 1814
rect 2662 1809 2668 1810
rect 2814 1814 2820 1815
rect 2814 1810 2815 1814
rect 2819 1810 2820 1814
rect 2814 1809 2820 1810
rect 2982 1814 2988 1815
rect 2982 1810 2983 1814
rect 2987 1810 2988 1814
rect 2982 1809 2988 1810
rect 3158 1814 3164 1815
rect 3158 1810 3159 1814
rect 3163 1810 3164 1814
rect 3158 1809 3164 1810
rect 3342 1814 3348 1815
rect 3342 1810 3343 1814
rect 3347 1810 3348 1814
rect 3342 1809 3348 1810
rect 3510 1814 3516 1815
rect 3510 1810 3511 1814
rect 3515 1810 3516 1814
rect 3510 1809 3516 1810
rect 1742 1807 1748 1808
rect 1902 1770 1908 1771
rect 1902 1766 1903 1770
rect 1907 1766 1908 1770
rect 1902 1765 1908 1766
rect 2030 1770 2036 1771
rect 2030 1766 2031 1770
rect 2035 1766 2036 1770
rect 2030 1765 2036 1766
rect 2190 1770 2196 1771
rect 2190 1766 2191 1770
rect 2195 1766 2196 1770
rect 2190 1765 2196 1766
rect 2358 1770 2364 1771
rect 2358 1766 2359 1770
rect 2363 1766 2364 1770
rect 2358 1765 2364 1766
rect 2526 1770 2532 1771
rect 2526 1766 2527 1770
rect 2531 1766 2532 1770
rect 2526 1765 2532 1766
rect 2686 1770 2692 1771
rect 2686 1766 2687 1770
rect 2691 1766 2692 1770
rect 2686 1765 2692 1766
rect 2838 1770 2844 1771
rect 2838 1766 2839 1770
rect 2843 1766 2844 1770
rect 2838 1765 2844 1766
rect 2982 1770 2988 1771
rect 2982 1766 2983 1770
rect 2987 1766 2988 1770
rect 2982 1765 2988 1766
rect 3118 1770 3124 1771
rect 3118 1766 3119 1770
rect 3123 1766 3124 1770
rect 3118 1765 3124 1766
rect 3254 1770 3260 1771
rect 3254 1766 3255 1770
rect 3259 1766 3260 1770
rect 3254 1765 3260 1766
rect 3390 1770 3396 1771
rect 3390 1766 3391 1770
rect 3395 1766 3396 1770
rect 3390 1765 3396 1766
rect 3510 1770 3516 1771
rect 3510 1766 3511 1770
rect 3515 1766 3516 1770
rect 3510 1765 3516 1766
rect 246 1764 252 1765
rect 110 1761 116 1762
rect 110 1757 111 1761
rect 115 1757 116 1761
rect 246 1760 247 1764
rect 251 1760 252 1764
rect 246 1759 252 1760
rect 422 1764 428 1765
rect 422 1760 423 1764
rect 427 1760 428 1764
rect 422 1759 428 1760
rect 590 1764 596 1765
rect 590 1760 591 1764
rect 595 1760 596 1764
rect 590 1759 596 1760
rect 750 1764 756 1765
rect 750 1760 751 1764
rect 755 1760 756 1764
rect 750 1759 756 1760
rect 894 1764 900 1765
rect 894 1760 895 1764
rect 899 1760 900 1764
rect 894 1759 900 1760
rect 1022 1764 1028 1765
rect 1022 1760 1023 1764
rect 1027 1760 1028 1764
rect 1022 1759 1028 1760
rect 1142 1764 1148 1765
rect 1142 1760 1143 1764
rect 1147 1760 1148 1764
rect 1142 1759 1148 1760
rect 1262 1764 1268 1765
rect 1262 1760 1263 1764
rect 1267 1760 1268 1764
rect 1262 1759 1268 1760
rect 1390 1764 1396 1765
rect 1390 1760 1391 1764
rect 1395 1760 1396 1764
rect 1390 1759 1396 1760
rect 1830 1761 1836 1762
rect 110 1756 116 1757
rect 1830 1757 1831 1761
rect 1835 1757 1836 1761
rect 1830 1756 1836 1757
rect 1870 1752 1876 1753
rect 1870 1748 1871 1752
rect 1875 1748 1876 1752
rect 1870 1747 1876 1748
rect 3590 1752 3596 1753
rect 3590 1748 3591 1752
rect 3595 1748 3596 1752
rect 3590 1747 3596 1748
rect 110 1744 116 1745
rect 110 1740 111 1744
rect 115 1740 116 1744
rect 110 1739 116 1740
rect 1830 1744 1836 1745
rect 1830 1740 1831 1744
rect 1835 1740 1836 1744
rect 1830 1739 1836 1740
rect 1870 1735 1876 1736
rect 1870 1731 1871 1735
rect 1875 1731 1876 1735
rect 3590 1735 3596 1736
rect 1870 1730 1876 1731
rect 1894 1732 1900 1733
rect 1894 1728 1895 1732
rect 1899 1728 1900 1732
rect 1894 1727 1900 1728
rect 2022 1732 2028 1733
rect 2022 1728 2023 1732
rect 2027 1728 2028 1732
rect 2022 1727 2028 1728
rect 2182 1732 2188 1733
rect 2182 1728 2183 1732
rect 2187 1728 2188 1732
rect 2182 1727 2188 1728
rect 2350 1732 2356 1733
rect 2350 1728 2351 1732
rect 2355 1728 2356 1732
rect 2350 1727 2356 1728
rect 2518 1732 2524 1733
rect 2518 1728 2519 1732
rect 2523 1728 2524 1732
rect 2518 1727 2524 1728
rect 2678 1732 2684 1733
rect 2678 1728 2679 1732
rect 2683 1728 2684 1732
rect 2678 1727 2684 1728
rect 2830 1732 2836 1733
rect 2830 1728 2831 1732
rect 2835 1728 2836 1732
rect 2830 1727 2836 1728
rect 2974 1732 2980 1733
rect 2974 1728 2975 1732
rect 2979 1728 2980 1732
rect 2974 1727 2980 1728
rect 3110 1732 3116 1733
rect 3110 1728 3111 1732
rect 3115 1728 3116 1732
rect 3110 1727 3116 1728
rect 3246 1732 3252 1733
rect 3246 1728 3247 1732
rect 3251 1728 3252 1732
rect 3246 1727 3252 1728
rect 3382 1732 3388 1733
rect 3382 1728 3383 1732
rect 3387 1728 3388 1732
rect 3382 1727 3388 1728
rect 3502 1732 3508 1733
rect 3502 1728 3503 1732
rect 3507 1728 3508 1732
rect 3590 1731 3591 1735
rect 3595 1731 3596 1735
rect 3590 1730 3596 1731
rect 3502 1727 3508 1728
rect 254 1726 260 1727
rect 254 1722 255 1726
rect 259 1722 260 1726
rect 254 1721 260 1722
rect 430 1726 436 1727
rect 430 1722 431 1726
rect 435 1722 436 1726
rect 430 1721 436 1722
rect 598 1726 604 1727
rect 598 1722 599 1726
rect 603 1722 604 1726
rect 598 1721 604 1722
rect 758 1726 764 1727
rect 758 1722 759 1726
rect 763 1722 764 1726
rect 758 1721 764 1722
rect 902 1726 908 1727
rect 902 1722 903 1726
rect 907 1722 908 1726
rect 902 1721 908 1722
rect 1030 1726 1036 1727
rect 1030 1722 1031 1726
rect 1035 1722 1036 1726
rect 1030 1721 1036 1722
rect 1150 1726 1156 1727
rect 1150 1722 1151 1726
rect 1155 1722 1156 1726
rect 1150 1721 1156 1722
rect 1270 1726 1276 1727
rect 1270 1722 1271 1726
rect 1275 1722 1276 1726
rect 1270 1721 1276 1722
rect 1398 1726 1404 1727
rect 1398 1722 1399 1726
rect 1403 1722 1404 1726
rect 1398 1721 1404 1722
rect 190 1690 196 1691
rect 190 1686 191 1690
rect 195 1686 196 1690
rect 190 1685 196 1686
rect 310 1690 316 1691
rect 310 1686 311 1690
rect 315 1686 316 1690
rect 310 1685 316 1686
rect 446 1690 452 1691
rect 446 1686 447 1690
rect 451 1686 452 1690
rect 446 1685 452 1686
rect 590 1690 596 1691
rect 590 1686 591 1690
rect 595 1686 596 1690
rect 590 1685 596 1686
rect 742 1690 748 1691
rect 742 1686 743 1690
rect 747 1686 748 1690
rect 742 1685 748 1686
rect 894 1690 900 1691
rect 894 1686 895 1690
rect 899 1686 900 1690
rect 894 1685 900 1686
rect 1038 1690 1044 1691
rect 1038 1686 1039 1690
rect 1043 1686 1044 1690
rect 1038 1685 1044 1686
rect 1182 1690 1188 1691
rect 1182 1686 1183 1690
rect 1187 1686 1188 1690
rect 1182 1685 1188 1686
rect 1318 1690 1324 1691
rect 1318 1686 1319 1690
rect 1323 1686 1324 1690
rect 1318 1685 1324 1686
rect 1446 1690 1452 1691
rect 1446 1686 1447 1690
rect 1451 1686 1452 1690
rect 1446 1685 1452 1686
rect 1574 1690 1580 1691
rect 1574 1686 1575 1690
rect 1579 1686 1580 1690
rect 1574 1685 1580 1686
rect 1710 1690 1716 1691
rect 1710 1686 1711 1690
rect 1715 1686 1716 1690
rect 1710 1685 1716 1686
rect 1894 1684 1900 1685
rect 1870 1681 1876 1682
rect 1870 1677 1871 1681
rect 1875 1677 1876 1681
rect 1894 1680 1895 1684
rect 1899 1680 1900 1684
rect 1894 1679 1900 1680
rect 1990 1684 1996 1685
rect 1990 1680 1991 1684
rect 1995 1680 1996 1684
rect 1990 1679 1996 1680
rect 2134 1684 2140 1685
rect 2134 1680 2135 1684
rect 2139 1680 2140 1684
rect 2134 1679 2140 1680
rect 2294 1684 2300 1685
rect 2294 1680 2295 1684
rect 2299 1680 2300 1684
rect 2294 1679 2300 1680
rect 2470 1684 2476 1685
rect 2470 1680 2471 1684
rect 2475 1680 2476 1684
rect 2470 1679 2476 1680
rect 2646 1684 2652 1685
rect 2646 1680 2647 1684
rect 2651 1680 2652 1684
rect 2646 1679 2652 1680
rect 2814 1684 2820 1685
rect 2814 1680 2815 1684
rect 2819 1680 2820 1684
rect 2814 1679 2820 1680
rect 2966 1684 2972 1685
rect 2966 1680 2967 1684
rect 2971 1680 2972 1684
rect 2966 1679 2972 1680
rect 3110 1684 3116 1685
rect 3110 1680 3111 1684
rect 3115 1680 3116 1684
rect 3110 1679 3116 1680
rect 3246 1684 3252 1685
rect 3246 1680 3247 1684
rect 3251 1680 3252 1684
rect 3246 1679 3252 1680
rect 3382 1684 3388 1685
rect 3382 1680 3383 1684
rect 3387 1680 3388 1684
rect 3382 1679 3388 1680
rect 3502 1684 3508 1685
rect 3502 1680 3503 1684
rect 3507 1680 3508 1684
rect 3502 1679 3508 1680
rect 3590 1681 3596 1682
rect 1870 1676 1876 1677
rect 3590 1677 3591 1681
rect 3595 1677 3596 1681
rect 3590 1676 3596 1677
rect 110 1672 116 1673
rect 110 1668 111 1672
rect 115 1668 116 1672
rect 110 1667 116 1668
rect 1830 1672 1836 1673
rect 1830 1668 1831 1672
rect 1835 1668 1836 1672
rect 1830 1667 1836 1668
rect 1870 1664 1876 1665
rect 1870 1660 1871 1664
rect 1875 1660 1876 1664
rect 1870 1659 1876 1660
rect 3590 1664 3596 1665
rect 3590 1660 3591 1664
rect 3595 1660 3596 1664
rect 3590 1659 3596 1660
rect 110 1655 116 1656
rect 110 1651 111 1655
rect 115 1651 116 1655
rect 1830 1655 1836 1656
rect 110 1650 116 1651
rect 182 1652 188 1653
rect 182 1648 183 1652
rect 187 1648 188 1652
rect 182 1647 188 1648
rect 302 1652 308 1653
rect 302 1648 303 1652
rect 307 1648 308 1652
rect 302 1647 308 1648
rect 438 1652 444 1653
rect 438 1648 439 1652
rect 443 1648 444 1652
rect 438 1647 444 1648
rect 582 1652 588 1653
rect 582 1648 583 1652
rect 587 1648 588 1652
rect 582 1647 588 1648
rect 734 1652 740 1653
rect 734 1648 735 1652
rect 739 1648 740 1652
rect 734 1647 740 1648
rect 886 1652 892 1653
rect 886 1648 887 1652
rect 891 1648 892 1652
rect 886 1647 892 1648
rect 1030 1652 1036 1653
rect 1030 1648 1031 1652
rect 1035 1648 1036 1652
rect 1030 1647 1036 1648
rect 1174 1652 1180 1653
rect 1174 1648 1175 1652
rect 1179 1648 1180 1652
rect 1174 1647 1180 1648
rect 1310 1652 1316 1653
rect 1310 1648 1311 1652
rect 1315 1648 1316 1652
rect 1310 1647 1316 1648
rect 1438 1652 1444 1653
rect 1438 1648 1439 1652
rect 1443 1648 1444 1652
rect 1438 1647 1444 1648
rect 1566 1652 1572 1653
rect 1566 1648 1567 1652
rect 1571 1648 1572 1652
rect 1566 1647 1572 1648
rect 1702 1652 1708 1653
rect 1702 1648 1703 1652
rect 1707 1648 1708 1652
rect 1830 1651 1831 1655
rect 1835 1651 1836 1655
rect 1830 1650 1836 1651
rect 1702 1647 1708 1648
rect 1902 1646 1908 1647
rect 1902 1642 1903 1646
rect 1907 1642 1908 1646
rect 1902 1641 1908 1642
rect 1998 1646 2004 1647
rect 1998 1642 1999 1646
rect 2003 1642 2004 1646
rect 1998 1641 2004 1642
rect 2142 1646 2148 1647
rect 2142 1642 2143 1646
rect 2147 1642 2148 1646
rect 2142 1641 2148 1642
rect 2302 1646 2308 1647
rect 2302 1642 2303 1646
rect 2307 1642 2308 1646
rect 2302 1641 2308 1642
rect 2478 1646 2484 1647
rect 2478 1642 2479 1646
rect 2483 1642 2484 1646
rect 2478 1641 2484 1642
rect 2654 1646 2660 1647
rect 2654 1642 2655 1646
rect 2659 1642 2660 1646
rect 2654 1641 2660 1642
rect 2822 1646 2828 1647
rect 2822 1642 2823 1646
rect 2827 1642 2828 1646
rect 2822 1641 2828 1642
rect 2974 1646 2980 1647
rect 2974 1642 2975 1646
rect 2979 1642 2980 1646
rect 2974 1641 2980 1642
rect 3118 1646 3124 1647
rect 3118 1642 3119 1646
rect 3123 1642 3124 1646
rect 3118 1641 3124 1642
rect 3254 1646 3260 1647
rect 3254 1642 3255 1646
rect 3259 1642 3260 1646
rect 3254 1641 3260 1642
rect 3390 1646 3396 1647
rect 3390 1642 3391 1646
rect 3395 1642 3396 1646
rect 3390 1641 3396 1642
rect 3510 1646 3516 1647
rect 3510 1642 3511 1646
rect 3515 1642 3516 1646
rect 3510 1641 3516 1642
rect 1974 1610 1980 1611
rect 1974 1606 1975 1610
rect 1979 1606 1980 1610
rect 1974 1605 1980 1606
rect 2094 1610 2100 1611
rect 2094 1606 2095 1610
rect 2099 1606 2100 1610
rect 2094 1605 2100 1606
rect 2230 1610 2236 1611
rect 2230 1606 2231 1610
rect 2235 1606 2236 1610
rect 2230 1605 2236 1606
rect 2366 1610 2372 1611
rect 2366 1606 2367 1610
rect 2371 1606 2372 1610
rect 2366 1605 2372 1606
rect 2502 1610 2508 1611
rect 2502 1606 2503 1610
rect 2507 1606 2508 1610
rect 2502 1605 2508 1606
rect 2638 1610 2644 1611
rect 2638 1606 2639 1610
rect 2643 1606 2644 1610
rect 2638 1605 2644 1606
rect 2774 1610 2780 1611
rect 2774 1606 2775 1610
rect 2779 1606 2780 1610
rect 2774 1605 2780 1606
rect 2910 1610 2916 1611
rect 2910 1606 2911 1610
rect 2915 1606 2916 1610
rect 2910 1605 2916 1606
rect 3054 1610 3060 1611
rect 3054 1606 3055 1610
rect 3059 1606 3060 1610
rect 3054 1605 3060 1606
rect 3206 1610 3212 1611
rect 3206 1606 3207 1610
rect 3211 1606 3212 1610
rect 3206 1605 3212 1606
rect 3366 1610 3372 1611
rect 3366 1606 3367 1610
rect 3371 1606 3372 1610
rect 3366 1605 3372 1606
rect 3510 1610 3516 1611
rect 3510 1606 3511 1610
rect 3515 1606 3516 1610
rect 3510 1605 3516 1606
rect 166 1600 172 1601
rect 110 1597 116 1598
rect 110 1593 111 1597
rect 115 1593 116 1597
rect 166 1596 167 1600
rect 171 1596 172 1600
rect 166 1595 172 1596
rect 350 1600 356 1601
rect 350 1596 351 1600
rect 355 1596 356 1600
rect 350 1595 356 1596
rect 542 1600 548 1601
rect 542 1596 543 1600
rect 547 1596 548 1600
rect 542 1595 548 1596
rect 726 1600 732 1601
rect 726 1596 727 1600
rect 731 1596 732 1600
rect 726 1595 732 1596
rect 902 1600 908 1601
rect 902 1596 903 1600
rect 907 1596 908 1600
rect 902 1595 908 1596
rect 1070 1600 1076 1601
rect 1070 1596 1071 1600
rect 1075 1596 1076 1600
rect 1070 1595 1076 1596
rect 1222 1600 1228 1601
rect 1222 1596 1223 1600
rect 1227 1596 1228 1600
rect 1222 1595 1228 1596
rect 1358 1600 1364 1601
rect 1358 1596 1359 1600
rect 1363 1596 1364 1600
rect 1358 1595 1364 1596
rect 1494 1600 1500 1601
rect 1494 1596 1495 1600
rect 1499 1596 1500 1600
rect 1494 1595 1500 1596
rect 1622 1600 1628 1601
rect 1622 1596 1623 1600
rect 1627 1596 1628 1600
rect 1622 1595 1628 1596
rect 1742 1600 1748 1601
rect 1742 1596 1743 1600
rect 1747 1596 1748 1600
rect 1742 1595 1748 1596
rect 1830 1597 1836 1598
rect 110 1592 116 1593
rect 1830 1593 1831 1597
rect 1835 1593 1836 1597
rect 1830 1592 1836 1593
rect 1870 1592 1876 1593
rect 1870 1588 1871 1592
rect 1875 1588 1876 1592
rect 1870 1587 1876 1588
rect 3590 1592 3596 1593
rect 3590 1588 3591 1592
rect 3595 1588 3596 1592
rect 3590 1587 3596 1588
rect 110 1580 116 1581
rect 110 1576 111 1580
rect 115 1576 116 1580
rect 110 1575 116 1576
rect 1830 1580 1836 1581
rect 1830 1576 1831 1580
rect 1835 1576 1836 1580
rect 1830 1575 1836 1576
rect 1870 1575 1876 1576
rect 1870 1571 1871 1575
rect 1875 1571 1876 1575
rect 3590 1575 3596 1576
rect 1870 1570 1876 1571
rect 1966 1572 1972 1573
rect 1966 1568 1967 1572
rect 1971 1568 1972 1572
rect 1966 1567 1972 1568
rect 2086 1572 2092 1573
rect 2086 1568 2087 1572
rect 2091 1568 2092 1572
rect 2086 1567 2092 1568
rect 2222 1572 2228 1573
rect 2222 1568 2223 1572
rect 2227 1568 2228 1572
rect 2222 1567 2228 1568
rect 2358 1572 2364 1573
rect 2358 1568 2359 1572
rect 2363 1568 2364 1572
rect 2358 1567 2364 1568
rect 2494 1572 2500 1573
rect 2494 1568 2495 1572
rect 2499 1568 2500 1572
rect 2494 1567 2500 1568
rect 2630 1572 2636 1573
rect 2630 1568 2631 1572
rect 2635 1568 2636 1572
rect 2630 1567 2636 1568
rect 2766 1572 2772 1573
rect 2766 1568 2767 1572
rect 2771 1568 2772 1572
rect 2766 1567 2772 1568
rect 2902 1572 2908 1573
rect 2902 1568 2903 1572
rect 2907 1568 2908 1572
rect 2902 1567 2908 1568
rect 3046 1572 3052 1573
rect 3046 1568 3047 1572
rect 3051 1568 3052 1572
rect 3046 1567 3052 1568
rect 3198 1572 3204 1573
rect 3198 1568 3199 1572
rect 3203 1568 3204 1572
rect 3198 1567 3204 1568
rect 3358 1572 3364 1573
rect 3358 1568 3359 1572
rect 3363 1568 3364 1572
rect 3358 1567 3364 1568
rect 3502 1572 3508 1573
rect 3502 1568 3503 1572
rect 3507 1568 3508 1572
rect 3590 1571 3591 1575
rect 3595 1571 3596 1575
rect 3590 1570 3596 1571
rect 3502 1567 3508 1568
rect 174 1562 180 1563
rect 174 1558 175 1562
rect 179 1558 180 1562
rect 174 1557 180 1558
rect 358 1562 364 1563
rect 358 1558 359 1562
rect 363 1558 364 1562
rect 358 1557 364 1558
rect 550 1562 556 1563
rect 550 1558 551 1562
rect 555 1558 556 1562
rect 550 1557 556 1558
rect 734 1562 740 1563
rect 734 1558 735 1562
rect 739 1558 740 1562
rect 734 1557 740 1558
rect 910 1562 916 1563
rect 910 1558 911 1562
rect 915 1558 916 1562
rect 910 1557 916 1558
rect 1078 1562 1084 1563
rect 1078 1558 1079 1562
rect 1083 1558 1084 1562
rect 1078 1557 1084 1558
rect 1230 1562 1236 1563
rect 1230 1558 1231 1562
rect 1235 1558 1236 1562
rect 1230 1557 1236 1558
rect 1366 1562 1372 1563
rect 1366 1558 1367 1562
rect 1371 1558 1372 1562
rect 1366 1557 1372 1558
rect 1502 1562 1508 1563
rect 1502 1558 1503 1562
rect 1507 1558 1508 1562
rect 1502 1557 1508 1558
rect 1630 1562 1636 1563
rect 1630 1558 1631 1562
rect 1635 1558 1636 1562
rect 1630 1557 1636 1558
rect 1750 1562 1756 1563
rect 1750 1558 1751 1562
rect 1755 1558 1756 1562
rect 1750 1557 1756 1558
rect 142 1526 148 1527
rect 142 1522 143 1526
rect 147 1522 148 1526
rect 142 1521 148 1522
rect 246 1526 252 1527
rect 246 1522 247 1526
rect 251 1522 252 1526
rect 246 1521 252 1522
rect 382 1526 388 1527
rect 382 1522 383 1526
rect 387 1522 388 1526
rect 382 1521 388 1522
rect 526 1526 532 1527
rect 526 1522 527 1526
rect 531 1522 532 1526
rect 526 1521 532 1522
rect 670 1526 676 1527
rect 670 1522 671 1526
rect 675 1522 676 1526
rect 670 1521 676 1522
rect 814 1526 820 1527
rect 814 1522 815 1526
rect 819 1522 820 1526
rect 814 1521 820 1522
rect 950 1526 956 1527
rect 950 1522 951 1526
rect 955 1522 956 1526
rect 950 1521 956 1522
rect 1078 1526 1084 1527
rect 1078 1522 1079 1526
rect 1083 1522 1084 1526
rect 1078 1521 1084 1522
rect 1206 1526 1212 1527
rect 1206 1522 1207 1526
rect 1211 1522 1212 1526
rect 1206 1521 1212 1522
rect 1334 1526 1340 1527
rect 1334 1522 1335 1526
rect 1339 1522 1340 1526
rect 1334 1521 1340 1522
rect 1470 1526 1476 1527
rect 1470 1522 1471 1526
rect 1475 1522 1476 1526
rect 2086 1524 2092 1525
rect 1470 1521 1476 1522
rect 1870 1521 1876 1522
rect 1870 1517 1871 1521
rect 1875 1517 1876 1521
rect 2086 1520 2087 1524
rect 2091 1520 2092 1524
rect 2086 1519 2092 1520
rect 2166 1524 2172 1525
rect 2166 1520 2167 1524
rect 2171 1520 2172 1524
rect 2166 1519 2172 1520
rect 2254 1524 2260 1525
rect 2254 1520 2255 1524
rect 2259 1520 2260 1524
rect 2254 1519 2260 1520
rect 2342 1524 2348 1525
rect 2342 1520 2343 1524
rect 2347 1520 2348 1524
rect 2342 1519 2348 1520
rect 2438 1524 2444 1525
rect 2438 1520 2439 1524
rect 2443 1520 2444 1524
rect 2438 1519 2444 1520
rect 2534 1524 2540 1525
rect 2534 1520 2535 1524
rect 2539 1520 2540 1524
rect 2534 1519 2540 1520
rect 2646 1524 2652 1525
rect 2646 1520 2647 1524
rect 2651 1520 2652 1524
rect 2646 1519 2652 1520
rect 2782 1524 2788 1525
rect 2782 1520 2783 1524
rect 2787 1520 2788 1524
rect 2782 1519 2788 1520
rect 2942 1524 2948 1525
rect 2942 1520 2943 1524
rect 2947 1520 2948 1524
rect 2942 1519 2948 1520
rect 3118 1524 3124 1525
rect 3118 1520 3119 1524
rect 3123 1520 3124 1524
rect 3118 1519 3124 1520
rect 3302 1524 3308 1525
rect 3302 1520 3303 1524
rect 3307 1520 3308 1524
rect 3302 1519 3308 1520
rect 3494 1524 3500 1525
rect 3494 1520 3495 1524
rect 3499 1520 3500 1524
rect 3494 1519 3500 1520
rect 3590 1521 3596 1522
rect 1870 1516 1876 1517
rect 3590 1517 3591 1521
rect 3595 1517 3596 1521
rect 3590 1516 3596 1517
rect 110 1508 116 1509
rect 110 1504 111 1508
rect 115 1504 116 1508
rect 110 1503 116 1504
rect 1830 1508 1836 1509
rect 1830 1504 1831 1508
rect 1835 1504 1836 1508
rect 1830 1503 1836 1504
rect 1870 1504 1876 1505
rect 1870 1500 1871 1504
rect 1875 1500 1876 1504
rect 1870 1499 1876 1500
rect 3590 1504 3596 1505
rect 3590 1500 3591 1504
rect 3595 1500 3596 1504
rect 3590 1499 3596 1500
rect 110 1491 116 1492
rect 110 1487 111 1491
rect 115 1487 116 1491
rect 1830 1491 1836 1492
rect 110 1486 116 1487
rect 134 1488 140 1489
rect 134 1484 135 1488
rect 139 1484 140 1488
rect 134 1483 140 1484
rect 238 1488 244 1489
rect 238 1484 239 1488
rect 243 1484 244 1488
rect 238 1483 244 1484
rect 374 1488 380 1489
rect 374 1484 375 1488
rect 379 1484 380 1488
rect 374 1483 380 1484
rect 518 1488 524 1489
rect 518 1484 519 1488
rect 523 1484 524 1488
rect 518 1483 524 1484
rect 662 1488 668 1489
rect 662 1484 663 1488
rect 667 1484 668 1488
rect 662 1483 668 1484
rect 806 1488 812 1489
rect 806 1484 807 1488
rect 811 1484 812 1488
rect 806 1483 812 1484
rect 942 1488 948 1489
rect 942 1484 943 1488
rect 947 1484 948 1488
rect 942 1483 948 1484
rect 1070 1488 1076 1489
rect 1070 1484 1071 1488
rect 1075 1484 1076 1488
rect 1070 1483 1076 1484
rect 1198 1488 1204 1489
rect 1198 1484 1199 1488
rect 1203 1484 1204 1488
rect 1198 1483 1204 1484
rect 1326 1488 1332 1489
rect 1326 1484 1327 1488
rect 1331 1484 1332 1488
rect 1326 1483 1332 1484
rect 1462 1488 1468 1489
rect 1462 1484 1463 1488
rect 1467 1484 1468 1488
rect 1830 1487 1831 1491
rect 1835 1487 1836 1491
rect 1830 1486 1836 1487
rect 2094 1486 2100 1487
rect 1462 1483 1468 1484
rect 2094 1482 2095 1486
rect 2099 1482 2100 1486
rect 2094 1481 2100 1482
rect 2174 1486 2180 1487
rect 2174 1482 2175 1486
rect 2179 1482 2180 1486
rect 2174 1481 2180 1482
rect 2262 1486 2268 1487
rect 2262 1482 2263 1486
rect 2267 1482 2268 1486
rect 2262 1481 2268 1482
rect 2350 1486 2356 1487
rect 2350 1482 2351 1486
rect 2355 1482 2356 1486
rect 2350 1481 2356 1482
rect 2446 1486 2452 1487
rect 2446 1482 2447 1486
rect 2451 1482 2452 1486
rect 2446 1481 2452 1482
rect 2542 1486 2548 1487
rect 2542 1482 2543 1486
rect 2547 1482 2548 1486
rect 2542 1481 2548 1482
rect 2654 1486 2660 1487
rect 2654 1482 2655 1486
rect 2659 1482 2660 1486
rect 2654 1481 2660 1482
rect 2790 1486 2796 1487
rect 2790 1482 2791 1486
rect 2795 1482 2796 1486
rect 2790 1481 2796 1482
rect 2950 1486 2956 1487
rect 2950 1482 2951 1486
rect 2955 1482 2956 1486
rect 2950 1481 2956 1482
rect 3126 1486 3132 1487
rect 3126 1482 3127 1486
rect 3131 1482 3132 1486
rect 3126 1481 3132 1482
rect 3310 1486 3316 1487
rect 3310 1482 3311 1486
rect 3315 1482 3316 1486
rect 3310 1481 3316 1482
rect 3502 1486 3508 1487
rect 3502 1482 3503 1486
rect 3507 1482 3508 1486
rect 3502 1481 3508 1482
rect 2262 1450 2268 1451
rect 2262 1446 2263 1450
rect 2267 1446 2268 1450
rect 2262 1445 2268 1446
rect 2342 1450 2348 1451
rect 2342 1446 2343 1450
rect 2347 1446 2348 1450
rect 2342 1445 2348 1446
rect 2422 1450 2428 1451
rect 2422 1446 2423 1450
rect 2427 1446 2428 1450
rect 2422 1445 2428 1446
rect 2502 1450 2508 1451
rect 2502 1446 2503 1450
rect 2507 1446 2508 1450
rect 2502 1445 2508 1446
rect 2606 1450 2612 1451
rect 2606 1446 2607 1450
rect 2611 1446 2612 1450
rect 2606 1445 2612 1446
rect 2734 1450 2740 1451
rect 2734 1446 2735 1450
rect 2739 1446 2740 1450
rect 2734 1445 2740 1446
rect 2894 1450 2900 1451
rect 2894 1446 2895 1450
rect 2899 1446 2900 1450
rect 2894 1445 2900 1446
rect 3078 1450 3084 1451
rect 3078 1446 3079 1450
rect 3083 1446 3084 1450
rect 3078 1445 3084 1446
rect 3278 1450 3284 1451
rect 3278 1446 3279 1450
rect 3283 1446 3284 1450
rect 3278 1445 3284 1446
rect 3478 1450 3484 1451
rect 3478 1446 3479 1450
rect 3483 1446 3484 1450
rect 3478 1445 3484 1446
rect 134 1440 140 1441
rect 110 1437 116 1438
rect 110 1433 111 1437
rect 115 1433 116 1437
rect 134 1436 135 1440
rect 139 1436 140 1440
rect 134 1435 140 1436
rect 230 1440 236 1441
rect 230 1436 231 1440
rect 235 1436 236 1440
rect 230 1435 236 1436
rect 358 1440 364 1441
rect 358 1436 359 1440
rect 363 1436 364 1440
rect 358 1435 364 1436
rect 478 1440 484 1441
rect 478 1436 479 1440
rect 483 1436 484 1440
rect 478 1435 484 1436
rect 598 1440 604 1441
rect 598 1436 599 1440
rect 603 1436 604 1440
rect 598 1435 604 1436
rect 718 1440 724 1441
rect 718 1436 719 1440
rect 723 1436 724 1440
rect 718 1435 724 1436
rect 830 1440 836 1441
rect 830 1436 831 1440
rect 835 1436 836 1440
rect 830 1435 836 1436
rect 934 1440 940 1441
rect 934 1436 935 1440
rect 939 1436 940 1440
rect 934 1435 940 1436
rect 1038 1440 1044 1441
rect 1038 1436 1039 1440
rect 1043 1436 1044 1440
rect 1038 1435 1044 1436
rect 1142 1440 1148 1441
rect 1142 1436 1143 1440
rect 1147 1436 1148 1440
rect 1142 1435 1148 1436
rect 1254 1440 1260 1441
rect 1254 1436 1255 1440
rect 1259 1436 1260 1440
rect 1254 1435 1260 1436
rect 1830 1437 1836 1438
rect 110 1432 116 1433
rect 1830 1433 1831 1437
rect 1835 1433 1836 1437
rect 1830 1432 1836 1433
rect 1870 1432 1876 1433
rect 1870 1428 1871 1432
rect 1875 1428 1876 1432
rect 1870 1427 1876 1428
rect 3590 1432 3596 1433
rect 3590 1428 3591 1432
rect 3595 1428 3596 1432
rect 3590 1427 3596 1428
rect 110 1420 116 1421
rect 110 1416 111 1420
rect 115 1416 116 1420
rect 110 1415 116 1416
rect 1830 1420 1836 1421
rect 1830 1416 1831 1420
rect 1835 1416 1836 1420
rect 1830 1415 1836 1416
rect 1870 1415 1876 1416
rect 1870 1411 1871 1415
rect 1875 1411 1876 1415
rect 3590 1415 3596 1416
rect 1870 1410 1876 1411
rect 2254 1412 2260 1413
rect 2254 1408 2255 1412
rect 2259 1408 2260 1412
rect 2254 1407 2260 1408
rect 2334 1412 2340 1413
rect 2334 1408 2335 1412
rect 2339 1408 2340 1412
rect 2334 1407 2340 1408
rect 2414 1412 2420 1413
rect 2414 1408 2415 1412
rect 2419 1408 2420 1412
rect 2414 1407 2420 1408
rect 2494 1412 2500 1413
rect 2494 1408 2495 1412
rect 2499 1408 2500 1412
rect 2494 1407 2500 1408
rect 2598 1412 2604 1413
rect 2598 1408 2599 1412
rect 2603 1408 2604 1412
rect 2598 1407 2604 1408
rect 2726 1412 2732 1413
rect 2726 1408 2727 1412
rect 2731 1408 2732 1412
rect 2726 1407 2732 1408
rect 2886 1412 2892 1413
rect 2886 1408 2887 1412
rect 2891 1408 2892 1412
rect 2886 1407 2892 1408
rect 3070 1412 3076 1413
rect 3070 1408 3071 1412
rect 3075 1408 3076 1412
rect 3070 1407 3076 1408
rect 3270 1412 3276 1413
rect 3270 1408 3271 1412
rect 3275 1408 3276 1412
rect 3270 1407 3276 1408
rect 3470 1412 3476 1413
rect 3470 1408 3471 1412
rect 3475 1408 3476 1412
rect 3590 1411 3591 1415
rect 3595 1411 3596 1415
rect 3590 1410 3596 1411
rect 3470 1407 3476 1408
rect 142 1402 148 1403
rect 142 1398 143 1402
rect 147 1398 148 1402
rect 142 1397 148 1398
rect 238 1402 244 1403
rect 238 1398 239 1402
rect 243 1398 244 1402
rect 238 1397 244 1398
rect 366 1402 372 1403
rect 366 1398 367 1402
rect 371 1398 372 1402
rect 366 1397 372 1398
rect 486 1402 492 1403
rect 486 1398 487 1402
rect 491 1398 492 1402
rect 486 1397 492 1398
rect 606 1402 612 1403
rect 606 1398 607 1402
rect 611 1398 612 1402
rect 606 1397 612 1398
rect 726 1402 732 1403
rect 726 1398 727 1402
rect 731 1398 732 1402
rect 726 1397 732 1398
rect 838 1402 844 1403
rect 838 1398 839 1402
rect 843 1398 844 1402
rect 838 1397 844 1398
rect 942 1402 948 1403
rect 942 1398 943 1402
rect 947 1398 948 1402
rect 942 1397 948 1398
rect 1046 1402 1052 1403
rect 1046 1398 1047 1402
rect 1051 1398 1052 1402
rect 1046 1397 1052 1398
rect 1150 1402 1156 1403
rect 1150 1398 1151 1402
rect 1155 1398 1156 1402
rect 1150 1397 1156 1398
rect 1262 1402 1268 1403
rect 1262 1398 1263 1402
rect 1267 1398 1268 1402
rect 1262 1397 1268 1398
rect 2262 1368 2268 1369
rect 1870 1365 1876 1366
rect 1870 1361 1871 1365
rect 1875 1361 1876 1365
rect 2262 1364 2263 1368
rect 2267 1364 2268 1368
rect 2262 1363 2268 1364
rect 2342 1368 2348 1369
rect 2342 1364 2343 1368
rect 2347 1364 2348 1368
rect 2342 1363 2348 1364
rect 2422 1368 2428 1369
rect 2422 1364 2423 1368
rect 2427 1364 2428 1368
rect 2422 1363 2428 1364
rect 2502 1368 2508 1369
rect 2502 1364 2503 1368
rect 2507 1364 2508 1368
rect 2502 1363 2508 1364
rect 2590 1368 2596 1369
rect 2590 1364 2591 1368
rect 2595 1364 2596 1368
rect 2590 1363 2596 1364
rect 2694 1368 2700 1369
rect 2694 1364 2695 1368
rect 2699 1364 2700 1368
rect 2694 1363 2700 1364
rect 2806 1368 2812 1369
rect 2806 1364 2807 1368
rect 2811 1364 2812 1368
rect 2806 1363 2812 1364
rect 2918 1368 2924 1369
rect 2918 1364 2919 1368
rect 2923 1364 2924 1368
rect 2918 1363 2924 1364
rect 3038 1368 3044 1369
rect 3038 1364 3039 1368
rect 3043 1364 3044 1368
rect 3038 1363 3044 1364
rect 3158 1368 3164 1369
rect 3158 1364 3159 1368
rect 3163 1364 3164 1368
rect 3158 1363 3164 1364
rect 3278 1368 3284 1369
rect 3278 1364 3279 1368
rect 3283 1364 3284 1368
rect 3278 1363 3284 1364
rect 3398 1368 3404 1369
rect 3398 1364 3399 1368
rect 3403 1364 3404 1368
rect 3398 1363 3404 1364
rect 3502 1368 3508 1369
rect 3502 1364 3503 1368
rect 3507 1364 3508 1368
rect 3502 1363 3508 1364
rect 3590 1365 3596 1366
rect 1870 1360 1876 1361
rect 3590 1361 3591 1365
rect 3595 1361 3596 1365
rect 3590 1360 3596 1361
rect 142 1354 148 1355
rect 142 1350 143 1354
rect 147 1350 148 1354
rect 142 1349 148 1350
rect 286 1354 292 1355
rect 286 1350 287 1354
rect 291 1350 292 1354
rect 286 1349 292 1350
rect 430 1354 436 1355
rect 430 1350 431 1354
rect 435 1350 436 1354
rect 430 1349 436 1350
rect 582 1354 588 1355
rect 582 1350 583 1354
rect 587 1350 588 1354
rect 582 1349 588 1350
rect 734 1354 740 1355
rect 734 1350 735 1354
rect 739 1350 740 1354
rect 734 1349 740 1350
rect 878 1354 884 1355
rect 878 1350 879 1354
rect 883 1350 884 1354
rect 878 1349 884 1350
rect 1022 1354 1028 1355
rect 1022 1350 1023 1354
rect 1027 1350 1028 1354
rect 1022 1349 1028 1350
rect 1166 1354 1172 1355
rect 1166 1350 1167 1354
rect 1171 1350 1172 1354
rect 1166 1349 1172 1350
rect 1318 1354 1324 1355
rect 1318 1350 1319 1354
rect 1323 1350 1324 1354
rect 1318 1349 1324 1350
rect 1470 1354 1476 1355
rect 1470 1350 1471 1354
rect 1475 1350 1476 1354
rect 1470 1349 1476 1350
rect 1622 1354 1628 1355
rect 1622 1350 1623 1354
rect 1627 1350 1628 1354
rect 1622 1349 1628 1350
rect 1870 1348 1876 1349
rect 1870 1344 1871 1348
rect 1875 1344 1876 1348
rect 1870 1343 1876 1344
rect 3590 1348 3596 1349
rect 3590 1344 3591 1348
rect 3595 1344 3596 1348
rect 3590 1343 3596 1344
rect 110 1336 116 1337
rect 110 1332 111 1336
rect 115 1332 116 1336
rect 110 1331 116 1332
rect 1830 1336 1836 1337
rect 1830 1332 1831 1336
rect 1835 1332 1836 1336
rect 1830 1331 1836 1332
rect 2270 1330 2276 1331
rect 2270 1326 2271 1330
rect 2275 1326 2276 1330
rect 2270 1325 2276 1326
rect 2350 1330 2356 1331
rect 2350 1326 2351 1330
rect 2355 1326 2356 1330
rect 2350 1325 2356 1326
rect 2430 1330 2436 1331
rect 2430 1326 2431 1330
rect 2435 1326 2436 1330
rect 2430 1325 2436 1326
rect 2510 1330 2516 1331
rect 2510 1326 2511 1330
rect 2515 1326 2516 1330
rect 2510 1325 2516 1326
rect 2598 1330 2604 1331
rect 2598 1326 2599 1330
rect 2603 1326 2604 1330
rect 2598 1325 2604 1326
rect 2702 1330 2708 1331
rect 2702 1326 2703 1330
rect 2707 1326 2708 1330
rect 2702 1325 2708 1326
rect 2814 1330 2820 1331
rect 2814 1326 2815 1330
rect 2819 1326 2820 1330
rect 2814 1325 2820 1326
rect 2926 1330 2932 1331
rect 2926 1326 2927 1330
rect 2931 1326 2932 1330
rect 2926 1325 2932 1326
rect 3046 1330 3052 1331
rect 3046 1326 3047 1330
rect 3051 1326 3052 1330
rect 3046 1325 3052 1326
rect 3166 1330 3172 1331
rect 3166 1326 3167 1330
rect 3171 1326 3172 1330
rect 3166 1325 3172 1326
rect 3286 1330 3292 1331
rect 3286 1326 3287 1330
rect 3291 1326 3292 1330
rect 3286 1325 3292 1326
rect 3406 1330 3412 1331
rect 3406 1326 3407 1330
rect 3411 1326 3412 1330
rect 3406 1325 3412 1326
rect 3510 1330 3516 1331
rect 3510 1326 3511 1330
rect 3515 1326 3516 1330
rect 3510 1325 3516 1326
rect 110 1319 116 1320
rect 110 1315 111 1319
rect 115 1315 116 1319
rect 1830 1319 1836 1320
rect 110 1314 116 1315
rect 134 1316 140 1317
rect 134 1312 135 1316
rect 139 1312 140 1316
rect 134 1311 140 1312
rect 278 1316 284 1317
rect 278 1312 279 1316
rect 283 1312 284 1316
rect 278 1311 284 1312
rect 422 1316 428 1317
rect 422 1312 423 1316
rect 427 1312 428 1316
rect 422 1311 428 1312
rect 574 1316 580 1317
rect 574 1312 575 1316
rect 579 1312 580 1316
rect 574 1311 580 1312
rect 726 1316 732 1317
rect 726 1312 727 1316
rect 731 1312 732 1316
rect 726 1311 732 1312
rect 870 1316 876 1317
rect 870 1312 871 1316
rect 875 1312 876 1316
rect 870 1311 876 1312
rect 1014 1316 1020 1317
rect 1014 1312 1015 1316
rect 1019 1312 1020 1316
rect 1014 1311 1020 1312
rect 1158 1316 1164 1317
rect 1158 1312 1159 1316
rect 1163 1312 1164 1316
rect 1158 1311 1164 1312
rect 1310 1316 1316 1317
rect 1310 1312 1311 1316
rect 1315 1312 1316 1316
rect 1310 1311 1316 1312
rect 1462 1316 1468 1317
rect 1462 1312 1463 1316
rect 1467 1312 1468 1316
rect 1462 1311 1468 1312
rect 1614 1316 1620 1317
rect 1614 1312 1615 1316
rect 1619 1312 1620 1316
rect 1830 1315 1831 1319
rect 1835 1315 1836 1319
rect 1830 1314 1836 1315
rect 1614 1311 1620 1312
rect 2214 1286 2220 1287
rect 2214 1282 2215 1286
rect 2219 1282 2220 1286
rect 2214 1281 2220 1282
rect 2294 1286 2300 1287
rect 2294 1282 2295 1286
rect 2299 1282 2300 1286
rect 2294 1281 2300 1282
rect 2374 1286 2380 1287
rect 2374 1282 2375 1286
rect 2379 1282 2380 1286
rect 2374 1281 2380 1282
rect 2454 1286 2460 1287
rect 2454 1282 2455 1286
rect 2459 1282 2460 1286
rect 2454 1281 2460 1282
rect 2550 1286 2556 1287
rect 2550 1282 2551 1286
rect 2555 1282 2556 1286
rect 2550 1281 2556 1282
rect 2662 1286 2668 1287
rect 2662 1282 2663 1286
rect 2667 1282 2668 1286
rect 2662 1281 2668 1282
rect 2790 1286 2796 1287
rect 2790 1282 2791 1286
rect 2795 1282 2796 1286
rect 2790 1281 2796 1282
rect 2926 1286 2932 1287
rect 2926 1282 2927 1286
rect 2931 1282 2932 1286
rect 2926 1281 2932 1282
rect 3070 1286 3076 1287
rect 3070 1282 3071 1286
rect 3075 1282 3076 1286
rect 3070 1281 3076 1282
rect 3214 1286 3220 1287
rect 3214 1282 3215 1286
rect 3219 1282 3220 1286
rect 3214 1281 3220 1282
rect 3366 1286 3372 1287
rect 3366 1282 3367 1286
rect 3371 1282 3372 1286
rect 3366 1281 3372 1282
rect 3510 1286 3516 1287
rect 3510 1282 3511 1286
rect 3515 1282 3516 1286
rect 3510 1281 3516 1282
rect 134 1268 140 1269
rect 110 1265 116 1266
rect 110 1261 111 1265
rect 115 1261 116 1265
rect 134 1264 135 1268
rect 139 1264 140 1268
rect 134 1263 140 1264
rect 262 1268 268 1269
rect 262 1264 263 1268
rect 267 1264 268 1268
rect 262 1263 268 1264
rect 422 1268 428 1269
rect 422 1264 423 1268
rect 427 1264 428 1268
rect 422 1263 428 1264
rect 590 1268 596 1269
rect 590 1264 591 1268
rect 595 1264 596 1268
rect 590 1263 596 1264
rect 758 1268 764 1269
rect 758 1264 759 1268
rect 763 1264 764 1268
rect 758 1263 764 1264
rect 926 1268 932 1269
rect 926 1264 927 1268
rect 931 1264 932 1268
rect 926 1263 932 1264
rect 1078 1268 1084 1269
rect 1078 1264 1079 1268
rect 1083 1264 1084 1268
rect 1078 1263 1084 1264
rect 1222 1268 1228 1269
rect 1222 1264 1223 1268
rect 1227 1264 1228 1268
rect 1222 1263 1228 1264
rect 1350 1268 1356 1269
rect 1350 1264 1351 1268
rect 1355 1264 1356 1268
rect 1350 1263 1356 1264
rect 1478 1268 1484 1269
rect 1478 1264 1479 1268
rect 1483 1264 1484 1268
rect 1478 1263 1484 1264
rect 1606 1268 1612 1269
rect 1606 1264 1607 1268
rect 1611 1264 1612 1268
rect 1606 1263 1612 1264
rect 1734 1268 1740 1269
rect 1734 1264 1735 1268
rect 1739 1264 1740 1268
rect 1870 1268 1876 1269
rect 1734 1263 1740 1264
rect 1830 1265 1836 1266
rect 110 1260 116 1261
rect 1830 1261 1831 1265
rect 1835 1261 1836 1265
rect 1870 1264 1871 1268
rect 1875 1264 1876 1268
rect 1870 1263 1876 1264
rect 3590 1268 3596 1269
rect 3590 1264 3591 1268
rect 3595 1264 3596 1268
rect 3590 1263 3596 1264
rect 1830 1260 1836 1261
rect 1870 1251 1876 1252
rect 110 1248 116 1249
rect 110 1244 111 1248
rect 115 1244 116 1248
rect 110 1243 116 1244
rect 1830 1248 1836 1249
rect 1830 1244 1831 1248
rect 1835 1244 1836 1248
rect 1870 1247 1871 1251
rect 1875 1247 1876 1251
rect 3590 1251 3596 1252
rect 1870 1246 1876 1247
rect 2206 1248 2212 1249
rect 1830 1243 1836 1244
rect 2206 1244 2207 1248
rect 2211 1244 2212 1248
rect 2206 1243 2212 1244
rect 2286 1248 2292 1249
rect 2286 1244 2287 1248
rect 2291 1244 2292 1248
rect 2286 1243 2292 1244
rect 2366 1248 2372 1249
rect 2366 1244 2367 1248
rect 2371 1244 2372 1248
rect 2366 1243 2372 1244
rect 2446 1248 2452 1249
rect 2446 1244 2447 1248
rect 2451 1244 2452 1248
rect 2446 1243 2452 1244
rect 2542 1248 2548 1249
rect 2542 1244 2543 1248
rect 2547 1244 2548 1248
rect 2542 1243 2548 1244
rect 2654 1248 2660 1249
rect 2654 1244 2655 1248
rect 2659 1244 2660 1248
rect 2654 1243 2660 1244
rect 2782 1248 2788 1249
rect 2782 1244 2783 1248
rect 2787 1244 2788 1248
rect 2782 1243 2788 1244
rect 2918 1248 2924 1249
rect 2918 1244 2919 1248
rect 2923 1244 2924 1248
rect 2918 1243 2924 1244
rect 3062 1248 3068 1249
rect 3062 1244 3063 1248
rect 3067 1244 3068 1248
rect 3062 1243 3068 1244
rect 3206 1248 3212 1249
rect 3206 1244 3207 1248
rect 3211 1244 3212 1248
rect 3206 1243 3212 1244
rect 3358 1248 3364 1249
rect 3358 1244 3359 1248
rect 3363 1244 3364 1248
rect 3358 1243 3364 1244
rect 3502 1248 3508 1249
rect 3502 1244 3503 1248
rect 3507 1244 3508 1248
rect 3590 1247 3591 1251
rect 3595 1247 3596 1251
rect 3590 1246 3596 1247
rect 3502 1243 3508 1244
rect 142 1230 148 1231
rect 142 1226 143 1230
rect 147 1226 148 1230
rect 142 1225 148 1226
rect 270 1230 276 1231
rect 270 1226 271 1230
rect 275 1226 276 1230
rect 270 1225 276 1226
rect 430 1230 436 1231
rect 430 1226 431 1230
rect 435 1226 436 1230
rect 430 1225 436 1226
rect 598 1230 604 1231
rect 598 1226 599 1230
rect 603 1226 604 1230
rect 598 1225 604 1226
rect 766 1230 772 1231
rect 766 1226 767 1230
rect 771 1226 772 1230
rect 766 1225 772 1226
rect 934 1230 940 1231
rect 934 1226 935 1230
rect 939 1226 940 1230
rect 934 1225 940 1226
rect 1086 1230 1092 1231
rect 1086 1226 1087 1230
rect 1091 1226 1092 1230
rect 1086 1225 1092 1226
rect 1230 1230 1236 1231
rect 1230 1226 1231 1230
rect 1235 1226 1236 1230
rect 1230 1225 1236 1226
rect 1358 1230 1364 1231
rect 1358 1226 1359 1230
rect 1363 1226 1364 1230
rect 1358 1225 1364 1226
rect 1486 1230 1492 1231
rect 1486 1226 1487 1230
rect 1491 1226 1492 1230
rect 1486 1225 1492 1226
rect 1614 1230 1620 1231
rect 1614 1226 1615 1230
rect 1619 1226 1620 1230
rect 1614 1225 1620 1226
rect 1742 1230 1748 1231
rect 1742 1226 1743 1230
rect 1747 1226 1748 1230
rect 1742 1225 1748 1226
rect 2110 1200 2116 1201
rect 1870 1197 1876 1198
rect 1870 1193 1871 1197
rect 1875 1193 1876 1197
rect 2110 1196 2111 1200
rect 2115 1196 2116 1200
rect 2110 1195 2116 1196
rect 2206 1200 2212 1201
rect 2206 1196 2207 1200
rect 2211 1196 2212 1200
rect 2206 1195 2212 1196
rect 2302 1200 2308 1201
rect 2302 1196 2303 1200
rect 2307 1196 2308 1200
rect 2302 1195 2308 1196
rect 2406 1200 2412 1201
rect 2406 1196 2407 1200
rect 2411 1196 2412 1200
rect 2406 1195 2412 1196
rect 2526 1200 2532 1201
rect 2526 1196 2527 1200
rect 2531 1196 2532 1200
rect 2526 1195 2532 1196
rect 2646 1200 2652 1201
rect 2646 1196 2647 1200
rect 2651 1196 2652 1200
rect 2646 1195 2652 1196
rect 2774 1200 2780 1201
rect 2774 1196 2775 1200
rect 2779 1196 2780 1200
rect 2774 1195 2780 1196
rect 2910 1200 2916 1201
rect 2910 1196 2911 1200
rect 2915 1196 2916 1200
rect 2910 1195 2916 1196
rect 3054 1200 3060 1201
rect 3054 1196 3055 1200
rect 3059 1196 3060 1200
rect 3054 1195 3060 1196
rect 3198 1200 3204 1201
rect 3198 1196 3199 1200
rect 3203 1196 3204 1200
rect 3198 1195 3204 1196
rect 3342 1200 3348 1201
rect 3342 1196 3343 1200
rect 3347 1196 3348 1200
rect 3342 1195 3348 1196
rect 3494 1200 3500 1201
rect 3494 1196 3495 1200
rect 3499 1196 3500 1200
rect 3494 1195 3500 1196
rect 3590 1197 3596 1198
rect 1870 1192 1876 1193
rect 3590 1193 3591 1197
rect 3595 1193 3596 1197
rect 3590 1192 3596 1193
rect 142 1190 148 1191
rect 142 1186 143 1190
rect 147 1186 148 1190
rect 142 1185 148 1186
rect 310 1190 316 1191
rect 310 1186 311 1190
rect 315 1186 316 1190
rect 310 1185 316 1186
rect 486 1190 492 1191
rect 486 1186 487 1190
rect 491 1186 492 1190
rect 486 1185 492 1186
rect 670 1190 676 1191
rect 670 1186 671 1190
rect 675 1186 676 1190
rect 670 1185 676 1186
rect 846 1190 852 1191
rect 846 1186 847 1190
rect 851 1186 852 1190
rect 846 1185 852 1186
rect 1006 1190 1012 1191
rect 1006 1186 1007 1190
rect 1011 1186 1012 1190
rect 1006 1185 1012 1186
rect 1158 1190 1164 1191
rect 1158 1186 1159 1190
rect 1163 1186 1164 1190
rect 1158 1185 1164 1186
rect 1294 1190 1300 1191
rect 1294 1186 1295 1190
rect 1299 1186 1300 1190
rect 1294 1185 1300 1186
rect 1414 1190 1420 1191
rect 1414 1186 1415 1190
rect 1419 1186 1420 1190
rect 1414 1185 1420 1186
rect 1534 1190 1540 1191
rect 1534 1186 1535 1190
rect 1539 1186 1540 1190
rect 1534 1185 1540 1186
rect 1654 1190 1660 1191
rect 1654 1186 1655 1190
rect 1659 1186 1660 1190
rect 1654 1185 1660 1186
rect 1750 1190 1756 1191
rect 1750 1186 1751 1190
rect 1755 1186 1756 1190
rect 1750 1185 1756 1186
rect 1870 1180 1876 1181
rect 1870 1176 1871 1180
rect 1875 1176 1876 1180
rect 1870 1175 1876 1176
rect 3590 1180 3596 1181
rect 3590 1176 3591 1180
rect 3595 1176 3596 1180
rect 3590 1175 3596 1176
rect 110 1172 116 1173
rect 110 1168 111 1172
rect 115 1168 116 1172
rect 110 1167 116 1168
rect 1830 1172 1836 1173
rect 1830 1168 1831 1172
rect 1835 1168 1836 1172
rect 1830 1167 1836 1168
rect 2118 1162 2124 1163
rect 2118 1158 2119 1162
rect 2123 1158 2124 1162
rect 2118 1157 2124 1158
rect 2214 1162 2220 1163
rect 2214 1158 2215 1162
rect 2219 1158 2220 1162
rect 2214 1157 2220 1158
rect 2310 1162 2316 1163
rect 2310 1158 2311 1162
rect 2315 1158 2316 1162
rect 2310 1157 2316 1158
rect 2414 1162 2420 1163
rect 2414 1158 2415 1162
rect 2419 1158 2420 1162
rect 2414 1157 2420 1158
rect 2534 1162 2540 1163
rect 2534 1158 2535 1162
rect 2539 1158 2540 1162
rect 2534 1157 2540 1158
rect 2654 1162 2660 1163
rect 2654 1158 2655 1162
rect 2659 1158 2660 1162
rect 2654 1157 2660 1158
rect 2782 1162 2788 1163
rect 2782 1158 2783 1162
rect 2787 1158 2788 1162
rect 2782 1157 2788 1158
rect 2918 1162 2924 1163
rect 2918 1158 2919 1162
rect 2923 1158 2924 1162
rect 2918 1157 2924 1158
rect 3062 1162 3068 1163
rect 3062 1158 3063 1162
rect 3067 1158 3068 1162
rect 3062 1157 3068 1158
rect 3206 1162 3212 1163
rect 3206 1158 3207 1162
rect 3211 1158 3212 1162
rect 3206 1157 3212 1158
rect 3350 1162 3356 1163
rect 3350 1158 3351 1162
rect 3355 1158 3356 1162
rect 3350 1157 3356 1158
rect 3502 1162 3508 1163
rect 3502 1158 3503 1162
rect 3507 1158 3508 1162
rect 3502 1157 3508 1158
rect 110 1155 116 1156
rect 110 1151 111 1155
rect 115 1151 116 1155
rect 1830 1155 1836 1156
rect 110 1150 116 1151
rect 134 1152 140 1153
rect 134 1148 135 1152
rect 139 1148 140 1152
rect 134 1147 140 1148
rect 302 1152 308 1153
rect 302 1148 303 1152
rect 307 1148 308 1152
rect 302 1147 308 1148
rect 478 1152 484 1153
rect 478 1148 479 1152
rect 483 1148 484 1152
rect 478 1147 484 1148
rect 662 1152 668 1153
rect 662 1148 663 1152
rect 667 1148 668 1152
rect 662 1147 668 1148
rect 838 1152 844 1153
rect 838 1148 839 1152
rect 843 1148 844 1152
rect 838 1147 844 1148
rect 998 1152 1004 1153
rect 998 1148 999 1152
rect 1003 1148 1004 1152
rect 998 1147 1004 1148
rect 1150 1152 1156 1153
rect 1150 1148 1151 1152
rect 1155 1148 1156 1152
rect 1150 1147 1156 1148
rect 1286 1152 1292 1153
rect 1286 1148 1287 1152
rect 1291 1148 1292 1152
rect 1286 1147 1292 1148
rect 1406 1152 1412 1153
rect 1406 1148 1407 1152
rect 1411 1148 1412 1152
rect 1406 1147 1412 1148
rect 1526 1152 1532 1153
rect 1526 1148 1527 1152
rect 1531 1148 1532 1152
rect 1526 1147 1532 1148
rect 1646 1152 1652 1153
rect 1646 1148 1647 1152
rect 1651 1148 1652 1152
rect 1646 1147 1652 1148
rect 1742 1152 1748 1153
rect 1742 1148 1743 1152
rect 1747 1148 1748 1152
rect 1830 1151 1831 1155
rect 1835 1151 1836 1155
rect 1830 1150 1836 1151
rect 1742 1147 1748 1148
rect 1902 1122 1908 1123
rect 1902 1118 1903 1122
rect 1907 1118 1908 1122
rect 1902 1117 1908 1118
rect 2126 1122 2132 1123
rect 2126 1118 2127 1122
rect 2131 1118 2132 1122
rect 2126 1117 2132 1118
rect 2358 1122 2364 1123
rect 2358 1118 2359 1122
rect 2363 1118 2364 1122
rect 2358 1117 2364 1118
rect 2574 1122 2580 1123
rect 2574 1118 2575 1122
rect 2579 1118 2580 1122
rect 2574 1117 2580 1118
rect 2774 1122 2780 1123
rect 2774 1118 2775 1122
rect 2779 1118 2780 1122
rect 2774 1117 2780 1118
rect 2966 1122 2972 1123
rect 2966 1118 2967 1122
rect 2971 1118 2972 1122
rect 2966 1117 2972 1118
rect 3158 1122 3164 1123
rect 3158 1118 3159 1122
rect 3163 1118 3164 1122
rect 3158 1117 3164 1118
rect 3342 1122 3348 1123
rect 3342 1118 3343 1122
rect 3347 1118 3348 1122
rect 3342 1117 3348 1118
rect 3510 1122 3516 1123
rect 3510 1118 3511 1122
rect 3515 1118 3516 1122
rect 3510 1117 3516 1118
rect 134 1108 140 1109
rect 110 1105 116 1106
rect 110 1101 111 1105
rect 115 1101 116 1105
rect 134 1104 135 1108
rect 139 1104 140 1108
rect 134 1103 140 1104
rect 246 1108 252 1109
rect 246 1104 247 1108
rect 251 1104 252 1108
rect 246 1103 252 1104
rect 382 1108 388 1109
rect 382 1104 383 1108
rect 387 1104 388 1108
rect 382 1103 388 1104
rect 518 1108 524 1109
rect 518 1104 519 1108
rect 523 1104 524 1108
rect 518 1103 524 1104
rect 646 1108 652 1109
rect 646 1104 647 1108
rect 651 1104 652 1108
rect 646 1103 652 1104
rect 774 1108 780 1109
rect 774 1104 775 1108
rect 779 1104 780 1108
rect 774 1103 780 1104
rect 894 1108 900 1109
rect 894 1104 895 1108
rect 899 1104 900 1108
rect 894 1103 900 1104
rect 1014 1108 1020 1109
rect 1014 1104 1015 1108
rect 1019 1104 1020 1108
rect 1014 1103 1020 1104
rect 1134 1108 1140 1109
rect 1134 1104 1135 1108
rect 1139 1104 1140 1108
rect 1134 1103 1140 1104
rect 1254 1108 1260 1109
rect 1254 1104 1255 1108
rect 1259 1104 1260 1108
rect 1254 1103 1260 1104
rect 1374 1108 1380 1109
rect 1374 1104 1375 1108
rect 1379 1104 1380 1108
rect 1374 1103 1380 1104
rect 1502 1108 1508 1109
rect 1502 1104 1503 1108
rect 1507 1104 1508 1108
rect 1502 1103 1508 1104
rect 1630 1108 1636 1109
rect 1630 1104 1631 1108
rect 1635 1104 1636 1108
rect 1630 1103 1636 1104
rect 1742 1108 1748 1109
rect 1742 1104 1743 1108
rect 1747 1104 1748 1108
rect 1742 1103 1748 1104
rect 1830 1105 1836 1106
rect 110 1100 116 1101
rect 1830 1101 1831 1105
rect 1835 1101 1836 1105
rect 1830 1100 1836 1101
rect 1870 1104 1876 1105
rect 1870 1100 1871 1104
rect 1875 1100 1876 1104
rect 1870 1099 1876 1100
rect 3590 1104 3596 1105
rect 3590 1100 3591 1104
rect 3595 1100 3596 1104
rect 3590 1099 3596 1100
rect 110 1088 116 1089
rect 110 1084 111 1088
rect 115 1084 116 1088
rect 110 1083 116 1084
rect 1830 1088 1836 1089
rect 1830 1084 1831 1088
rect 1835 1084 1836 1088
rect 1830 1083 1836 1084
rect 1870 1087 1876 1088
rect 1870 1083 1871 1087
rect 1875 1083 1876 1087
rect 3590 1087 3596 1088
rect 1870 1082 1876 1083
rect 1894 1084 1900 1085
rect 1894 1080 1895 1084
rect 1899 1080 1900 1084
rect 1894 1079 1900 1080
rect 2118 1084 2124 1085
rect 2118 1080 2119 1084
rect 2123 1080 2124 1084
rect 2118 1079 2124 1080
rect 2350 1084 2356 1085
rect 2350 1080 2351 1084
rect 2355 1080 2356 1084
rect 2350 1079 2356 1080
rect 2566 1084 2572 1085
rect 2566 1080 2567 1084
rect 2571 1080 2572 1084
rect 2566 1079 2572 1080
rect 2766 1084 2772 1085
rect 2766 1080 2767 1084
rect 2771 1080 2772 1084
rect 2766 1079 2772 1080
rect 2958 1084 2964 1085
rect 2958 1080 2959 1084
rect 2963 1080 2964 1084
rect 2958 1079 2964 1080
rect 3150 1084 3156 1085
rect 3150 1080 3151 1084
rect 3155 1080 3156 1084
rect 3150 1079 3156 1080
rect 3334 1084 3340 1085
rect 3334 1080 3335 1084
rect 3339 1080 3340 1084
rect 3334 1079 3340 1080
rect 3502 1084 3508 1085
rect 3502 1080 3503 1084
rect 3507 1080 3508 1084
rect 3590 1083 3591 1087
rect 3595 1083 3596 1087
rect 3590 1082 3596 1083
rect 3502 1079 3508 1080
rect 142 1070 148 1071
rect 142 1066 143 1070
rect 147 1066 148 1070
rect 142 1065 148 1066
rect 254 1070 260 1071
rect 254 1066 255 1070
rect 259 1066 260 1070
rect 254 1065 260 1066
rect 390 1070 396 1071
rect 390 1066 391 1070
rect 395 1066 396 1070
rect 390 1065 396 1066
rect 526 1070 532 1071
rect 526 1066 527 1070
rect 531 1066 532 1070
rect 526 1065 532 1066
rect 654 1070 660 1071
rect 654 1066 655 1070
rect 659 1066 660 1070
rect 654 1065 660 1066
rect 782 1070 788 1071
rect 782 1066 783 1070
rect 787 1066 788 1070
rect 782 1065 788 1066
rect 902 1070 908 1071
rect 902 1066 903 1070
rect 907 1066 908 1070
rect 902 1065 908 1066
rect 1022 1070 1028 1071
rect 1022 1066 1023 1070
rect 1027 1066 1028 1070
rect 1022 1065 1028 1066
rect 1142 1070 1148 1071
rect 1142 1066 1143 1070
rect 1147 1066 1148 1070
rect 1142 1065 1148 1066
rect 1262 1070 1268 1071
rect 1262 1066 1263 1070
rect 1267 1066 1268 1070
rect 1262 1065 1268 1066
rect 1382 1070 1388 1071
rect 1382 1066 1383 1070
rect 1387 1066 1388 1070
rect 1382 1065 1388 1066
rect 1510 1070 1516 1071
rect 1510 1066 1511 1070
rect 1515 1066 1516 1070
rect 1510 1065 1516 1066
rect 1638 1070 1644 1071
rect 1638 1066 1639 1070
rect 1643 1066 1644 1070
rect 1638 1065 1644 1066
rect 1750 1070 1756 1071
rect 1750 1066 1751 1070
rect 1755 1066 1756 1070
rect 1750 1065 1756 1066
rect 1894 1040 1900 1041
rect 1870 1037 1876 1038
rect 1870 1033 1871 1037
rect 1875 1033 1876 1037
rect 1894 1036 1895 1040
rect 1899 1036 1900 1040
rect 1894 1035 1900 1036
rect 2014 1040 2020 1041
rect 2014 1036 2015 1040
rect 2019 1036 2020 1040
rect 2014 1035 2020 1036
rect 2166 1040 2172 1041
rect 2166 1036 2167 1040
rect 2171 1036 2172 1040
rect 2166 1035 2172 1036
rect 2326 1040 2332 1041
rect 2326 1036 2327 1040
rect 2331 1036 2332 1040
rect 2326 1035 2332 1036
rect 2486 1040 2492 1041
rect 2486 1036 2487 1040
rect 2491 1036 2492 1040
rect 2486 1035 2492 1036
rect 2638 1040 2644 1041
rect 2638 1036 2639 1040
rect 2643 1036 2644 1040
rect 2638 1035 2644 1036
rect 2790 1040 2796 1041
rect 2790 1036 2791 1040
rect 2795 1036 2796 1040
rect 2790 1035 2796 1036
rect 2934 1040 2940 1041
rect 2934 1036 2935 1040
rect 2939 1036 2940 1040
rect 2934 1035 2940 1036
rect 3078 1040 3084 1041
rect 3078 1036 3079 1040
rect 3083 1036 3084 1040
rect 3078 1035 3084 1036
rect 3222 1040 3228 1041
rect 3222 1036 3223 1040
rect 3227 1036 3228 1040
rect 3222 1035 3228 1036
rect 3374 1040 3380 1041
rect 3374 1036 3375 1040
rect 3379 1036 3380 1040
rect 3374 1035 3380 1036
rect 3502 1040 3508 1041
rect 3502 1036 3503 1040
rect 3507 1036 3508 1040
rect 3502 1035 3508 1036
rect 3590 1037 3596 1038
rect 1870 1032 1876 1033
rect 3590 1033 3591 1037
rect 3595 1033 3596 1037
rect 3590 1032 3596 1033
rect 142 1026 148 1027
rect 142 1022 143 1026
rect 147 1022 148 1026
rect 142 1021 148 1022
rect 238 1026 244 1027
rect 238 1022 239 1026
rect 243 1022 244 1026
rect 238 1021 244 1022
rect 358 1026 364 1027
rect 358 1022 359 1026
rect 363 1022 364 1026
rect 358 1021 364 1022
rect 470 1026 476 1027
rect 470 1022 471 1026
rect 475 1022 476 1026
rect 470 1021 476 1022
rect 574 1026 580 1027
rect 574 1022 575 1026
rect 579 1022 580 1026
rect 574 1021 580 1022
rect 670 1026 676 1027
rect 670 1022 671 1026
rect 675 1022 676 1026
rect 670 1021 676 1022
rect 766 1026 772 1027
rect 766 1022 767 1026
rect 771 1022 772 1026
rect 766 1021 772 1022
rect 854 1026 860 1027
rect 854 1022 855 1026
rect 859 1022 860 1026
rect 854 1021 860 1022
rect 942 1026 948 1027
rect 942 1022 943 1026
rect 947 1022 948 1026
rect 942 1021 948 1022
rect 1030 1026 1036 1027
rect 1030 1022 1031 1026
rect 1035 1022 1036 1026
rect 1030 1021 1036 1022
rect 1126 1026 1132 1027
rect 1126 1022 1127 1026
rect 1131 1022 1132 1026
rect 1126 1021 1132 1022
rect 1222 1026 1228 1027
rect 1222 1022 1223 1026
rect 1227 1022 1228 1026
rect 1222 1021 1228 1022
rect 1870 1020 1876 1021
rect 1870 1016 1871 1020
rect 1875 1016 1876 1020
rect 1870 1015 1876 1016
rect 3590 1020 3596 1021
rect 3590 1016 3591 1020
rect 3595 1016 3596 1020
rect 3590 1015 3596 1016
rect 110 1008 116 1009
rect 110 1004 111 1008
rect 115 1004 116 1008
rect 110 1003 116 1004
rect 1830 1008 1836 1009
rect 1830 1004 1831 1008
rect 1835 1004 1836 1008
rect 1830 1003 1836 1004
rect 1902 1002 1908 1003
rect 1902 998 1903 1002
rect 1907 998 1908 1002
rect 1902 997 1908 998
rect 2022 1002 2028 1003
rect 2022 998 2023 1002
rect 2027 998 2028 1002
rect 2022 997 2028 998
rect 2174 1002 2180 1003
rect 2174 998 2175 1002
rect 2179 998 2180 1002
rect 2174 997 2180 998
rect 2334 1002 2340 1003
rect 2334 998 2335 1002
rect 2339 998 2340 1002
rect 2334 997 2340 998
rect 2494 1002 2500 1003
rect 2494 998 2495 1002
rect 2499 998 2500 1002
rect 2494 997 2500 998
rect 2646 1002 2652 1003
rect 2646 998 2647 1002
rect 2651 998 2652 1002
rect 2646 997 2652 998
rect 2798 1002 2804 1003
rect 2798 998 2799 1002
rect 2803 998 2804 1002
rect 2798 997 2804 998
rect 2942 1002 2948 1003
rect 2942 998 2943 1002
rect 2947 998 2948 1002
rect 2942 997 2948 998
rect 3086 1002 3092 1003
rect 3086 998 3087 1002
rect 3091 998 3092 1002
rect 3086 997 3092 998
rect 3230 1002 3236 1003
rect 3230 998 3231 1002
rect 3235 998 3236 1002
rect 3230 997 3236 998
rect 3382 1002 3388 1003
rect 3382 998 3383 1002
rect 3387 998 3388 1002
rect 3382 997 3388 998
rect 3510 1002 3516 1003
rect 3510 998 3511 1002
rect 3515 998 3516 1002
rect 3510 997 3516 998
rect 110 991 116 992
rect 110 987 111 991
rect 115 987 116 991
rect 1830 991 1836 992
rect 110 986 116 987
rect 134 988 140 989
rect 134 984 135 988
rect 139 984 140 988
rect 134 983 140 984
rect 230 988 236 989
rect 230 984 231 988
rect 235 984 236 988
rect 230 983 236 984
rect 350 988 356 989
rect 350 984 351 988
rect 355 984 356 988
rect 350 983 356 984
rect 462 988 468 989
rect 462 984 463 988
rect 467 984 468 988
rect 462 983 468 984
rect 566 988 572 989
rect 566 984 567 988
rect 571 984 572 988
rect 566 983 572 984
rect 662 988 668 989
rect 662 984 663 988
rect 667 984 668 988
rect 662 983 668 984
rect 758 988 764 989
rect 758 984 759 988
rect 763 984 764 988
rect 758 983 764 984
rect 846 988 852 989
rect 846 984 847 988
rect 851 984 852 988
rect 846 983 852 984
rect 934 988 940 989
rect 934 984 935 988
rect 939 984 940 988
rect 934 983 940 984
rect 1022 988 1028 989
rect 1022 984 1023 988
rect 1027 984 1028 988
rect 1022 983 1028 984
rect 1118 988 1124 989
rect 1118 984 1119 988
rect 1123 984 1124 988
rect 1118 983 1124 984
rect 1214 988 1220 989
rect 1214 984 1215 988
rect 1219 984 1220 988
rect 1830 987 1831 991
rect 1835 987 1836 991
rect 1830 986 1836 987
rect 1214 983 1220 984
rect 1902 966 1908 967
rect 1902 962 1903 966
rect 1907 962 1908 966
rect 1902 961 1908 962
rect 1982 966 1988 967
rect 1982 962 1983 966
rect 1987 962 1988 966
rect 1982 961 1988 962
rect 2078 966 2084 967
rect 2078 962 2079 966
rect 2083 962 2084 966
rect 2078 961 2084 962
rect 2198 966 2204 967
rect 2198 962 2199 966
rect 2203 962 2204 966
rect 2198 961 2204 962
rect 2334 966 2340 967
rect 2334 962 2335 966
rect 2339 962 2340 966
rect 2334 961 2340 962
rect 2478 966 2484 967
rect 2478 962 2479 966
rect 2483 962 2484 966
rect 2478 961 2484 962
rect 2630 966 2636 967
rect 2630 962 2631 966
rect 2635 962 2636 966
rect 2630 961 2636 962
rect 2790 966 2796 967
rect 2790 962 2791 966
rect 2795 962 2796 966
rect 2790 961 2796 962
rect 2966 966 2972 967
rect 2966 962 2967 966
rect 2971 962 2972 966
rect 2966 961 2972 962
rect 3150 966 3156 967
rect 3150 962 3151 966
rect 3155 962 3156 966
rect 3150 961 3156 962
rect 3342 966 3348 967
rect 3342 962 3343 966
rect 3347 962 3348 966
rect 3342 961 3348 962
rect 3510 966 3516 967
rect 3510 962 3511 966
rect 3515 962 3516 966
rect 3510 961 3516 962
rect 1870 948 1876 949
rect 1870 944 1871 948
rect 1875 944 1876 948
rect 1870 943 1876 944
rect 3590 948 3596 949
rect 3590 944 3591 948
rect 3595 944 3596 948
rect 3590 943 3596 944
rect 134 932 140 933
rect 110 929 116 930
rect 110 925 111 929
rect 115 925 116 929
rect 134 928 135 932
rect 139 928 140 932
rect 134 927 140 928
rect 262 932 268 933
rect 262 928 263 932
rect 267 928 268 932
rect 262 927 268 928
rect 414 932 420 933
rect 414 928 415 932
rect 419 928 420 932
rect 414 927 420 928
rect 558 932 564 933
rect 558 928 559 932
rect 563 928 564 932
rect 558 927 564 928
rect 702 932 708 933
rect 702 928 703 932
rect 707 928 708 932
rect 702 927 708 928
rect 838 932 844 933
rect 838 928 839 932
rect 843 928 844 932
rect 838 927 844 928
rect 974 932 980 933
rect 974 928 975 932
rect 979 928 980 932
rect 974 927 980 928
rect 1102 932 1108 933
rect 1102 928 1103 932
rect 1107 928 1108 932
rect 1102 927 1108 928
rect 1222 932 1228 933
rect 1222 928 1223 932
rect 1227 928 1228 932
rect 1222 927 1228 928
rect 1334 932 1340 933
rect 1334 928 1335 932
rect 1339 928 1340 932
rect 1334 927 1340 928
rect 1438 932 1444 933
rect 1438 928 1439 932
rect 1443 928 1444 932
rect 1438 927 1444 928
rect 1542 932 1548 933
rect 1542 928 1543 932
rect 1547 928 1548 932
rect 1542 927 1548 928
rect 1654 932 1660 933
rect 1654 928 1655 932
rect 1659 928 1660 932
rect 1654 927 1660 928
rect 1742 932 1748 933
rect 1742 928 1743 932
rect 1747 928 1748 932
rect 1870 931 1876 932
rect 1742 927 1748 928
rect 1830 929 1836 930
rect 110 924 116 925
rect 1830 925 1831 929
rect 1835 925 1836 929
rect 1870 927 1871 931
rect 1875 927 1876 931
rect 3590 931 3596 932
rect 1870 926 1876 927
rect 1894 928 1900 929
rect 1830 924 1836 925
rect 1894 924 1895 928
rect 1899 924 1900 928
rect 1894 923 1900 924
rect 1974 928 1980 929
rect 1974 924 1975 928
rect 1979 924 1980 928
rect 1974 923 1980 924
rect 2070 928 2076 929
rect 2070 924 2071 928
rect 2075 924 2076 928
rect 2070 923 2076 924
rect 2190 928 2196 929
rect 2190 924 2191 928
rect 2195 924 2196 928
rect 2190 923 2196 924
rect 2326 928 2332 929
rect 2326 924 2327 928
rect 2331 924 2332 928
rect 2326 923 2332 924
rect 2470 928 2476 929
rect 2470 924 2471 928
rect 2475 924 2476 928
rect 2470 923 2476 924
rect 2622 928 2628 929
rect 2622 924 2623 928
rect 2627 924 2628 928
rect 2622 923 2628 924
rect 2782 928 2788 929
rect 2782 924 2783 928
rect 2787 924 2788 928
rect 2782 923 2788 924
rect 2958 928 2964 929
rect 2958 924 2959 928
rect 2963 924 2964 928
rect 2958 923 2964 924
rect 3142 928 3148 929
rect 3142 924 3143 928
rect 3147 924 3148 928
rect 3142 923 3148 924
rect 3334 928 3340 929
rect 3334 924 3335 928
rect 3339 924 3340 928
rect 3334 923 3340 924
rect 3502 928 3508 929
rect 3502 924 3503 928
rect 3507 924 3508 928
rect 3590 927 3591 931
rect 3595 927 3596 931
rect 3590 926 3596 927
rect 3502 923 3508 924
rect 110 912 116 913
rect 110 908 111 912
rect 115 908 116 912
rect 110 907 116 908
rect 1830 912 1836 913
rect 1830 908 1831 912
rect 1835 908 1836 912
rect 1830 907 1836 908
rect 142 894 148 895
rect 142 890 143 894
rect 147 890 148 894
rect 142 889 148 890
rect 270 894 276 895
rect 270 890 271 894
rect 275 890 276 894
rect 270 889 276 890
rect 422 894 428 895
rect 422 890 423 894
rect 427 890 428 894
rect 422 889 428 890
rect 566 894 572 895
rect 566 890 567 894
rect 571 890 572 894
rect 566 889 572 890
rect 710 894 716 895
rect 710 890 711 894
rect 715 890 716 894
rect 710 889 716 890
rect 846 894 852 895
rect 846 890 847 894
rect 851 890 852 894
rect 846 889 852 890
rect 982 894 988 895
rect 982 890 983 894
rect 987 890 988 894
rect 982 889 988 890
rect 1110 894 1116 895
rect 1110 890 1111 894
rect 1115 890 1116 894
rect 1110 889 1116 890
rect 1230 894 1236 895
rect 1230 890 1231 894
rect 1235 890 1236 894
rect 1230 889 1236 890
rect 1342 894 1348 895
rect 1342 890 1343 894
rect 1347 890 1348 894
rect 1342 889 1348 890
rect 1446 894 1452 895
rect 1446 890 1447 894
rect 1451 890 1452 894
rect 1446 889 1452 890
rect 1550 894 1556 895
rect 1550 890 1551 894
rect 1555 890 1556 894
rect 1550 889 1556 890
rect 1662 894 1668 895
rect 1662 890 1663 894
rect 1667 890 1668 894
rect 1662 889 1668 890
rect 1750 894 1756 895
rect 1750 890 1751 894
rect 1755 890 1756 894
rect 1750 889 1756 890
rect 1918 872 1924 873
rect 1870 869 1876 870
rect 1870 865 1871 869
rect 1875 865 1876 869
rect 1918 868 1919 872
rect 1923 868 1924 872
rect 1918 867 1924 868
rect 2094 872 2100 873
rect 2094 868 2095 872
rect 2099 868 2100 872
rect 2094 867 2100 868
rect 2270 872 2276 873
rect 2270 868 2271 872
rect 2275 868 2276 872
rect 2270 867 2276 868
rect 2454 872 2460 873
rect 2454 868 2455 872
rect 2459 868 2460 872
rect 2454 867 2460 868
rect 2654 872 2660 873
rect 2654 868 2655 872
rect 2659 868 2660 872
rect 2654 867 2660 868
rect 2862 872 2868 873
rect 2862 868 2863 872
rect 2867 868 2868 872
rect 2862 867 2868 868
rect 3078 872 3084 873
rect 3078 868 3079 872
rect 3083 868 3084 872
rect 3078 867 3084 868
rect 3302 872 3308 873
rect 3302 868 3303 872
rect 3307 868 3308 872
rect 3302 867 3308 868
rect 3502 872 3508 873
rect 3502 868 3503 872
rect 3507 868 3508 872
rect 3502 867 3508 868
rect 3590 869 3596 870
rect 1870 864 1876 865
rect 3590 865 3591 869
rect 3595 865 3596 869
rect 3590 864 3596 865
rect 142 858 148 859
rect 142 854 143 858
rect 147 854 148 858
rect 142 853 148 854
rect 246 858 252 859
rect 246 854 247 858
rect 251 854 252 858
rect 246 853 252 854
rect 382 858 388 859
rect 382 854 383 858
rect 387 854 388 858
rect 382 853 388 854
rect 518 858 524 859
rect 518 854 519 858
rect 523 854 524 858
rect 518 853 524 854
rect 662 858 668 859
rect 662 854 663 858
rect 667 854 668 858
rect 662 853 668 854
rect 814 858 820 859
rect 814 854 815 858
rect 819 854 820 858
rect 814 853 820 854
rect 958 858 964 859
rect 958 854 959 858
rect 963 854 964 858
rect 958 853 964 854
rect 1102 858 1108 859
rect 1102 854 1103 858
rect 1107 854 1108 858
rect 1102 853 1108 854
rect 1246 858 1252 859
rect 1246 854 1247 858
rect 1251 854 1252 858
rect 1246 853 1252 854
rect 1382 858 1388 859
rect 1382 854 1383 858
rect 1387 854 1388 858
rect 1382 853 1388 854
rect 1510 858 1516 859
rect 1510 854 1511 858
rect 1515 854 1516 858
rect 1510 853 1516 854
rect 1638 858 1644 859
rect 1638 854 1639 858
rect 1643 854 1644 858
rect 1638 853 1644 854
rect 1750 858 1756 859
rect 1750 854 1751 858
rect 1755 854 1756 858
rect 1750 853 1756 854
rect 1870 852 1876 853
rect 1870 848 1871 852
rect 1875 848 1876 852
rect 1870 847 1876 848
rect 3590 852 3596 853
rect 3590 848 3591 852
rect 3595 848 3596 852
rect 3590 847 3596 848
rect 110 840 116 841
rect 110 836 111 840
rect 115 836 116 840
rect 110 835 116 836
rect 1830 840 1836 841
rect 1830 836 1831 840
rect 1835 836 1836 840
rect 1830 835 1836 836
rect 1926 834 1932 835
rect 1926 830 1927 834
rect 1931 830 1932 834
rect 1926 829 1932 830
rect 2102 834 2108 835
rect 2102 830 2103 834
rect 2107 830 2108 834
rect 2102 829 2108 830
rect 2278 834 2284 835
rect 2278 830 2279 834
rect 2283 830 2284 834
rect 2278 829 2284 830
rect 2462 834 2468 835
rect 2462 830 2463 834
rect 2467 830 2468 834
rect 2462 829 2468 830
rect 2662 834 2668 835
rect 2662 830 2663 834
rect 2667 830 2668 834
rect 2662 829 2668 830
rect 2870 834 2876 835
rect 2870 830 2871 834
rect 2875 830 2876 834
rect 2870 829 2876 830
rect 3086 834 3092 835
rect 3086 830 3087 834
rect 3091 830 3092 834
rect 3086 829 3092 830
rect 3310 834 3316 835
rect 3310 830 3311 834
rect 3315 830 3316 834
rect 3310 829 3316 830
rect 3510 834 3516 835
rect 3510 830 3511 834
rect 3515 830 3516 834
rect 3510 829 3516 830
rect 110 823 116 824
rect 110 819 111 823
rect 115 819 116 823
rect 1830 823 1836 824
rect 110 818 116 819
rect 134 820 140 821
rect 134 816 135 820
rect 139 816 140 820
rect 134 815 140 816
rect 238 820 244 821
rect 238 816 239 820
rect 243 816 244 820
rect 238 815 244 816
rect 374 820 380 821
rect 374 816 375 820
rect 379 816 380 820
rect 374 815 380 816
rect 510 820 516 821
rect 510 816 511 820
rect 515 816 516 820
rect 510 815 516 816
rect 654 820 660 821
rect 654 816 655 820
rect 659 816 660 820
rect 654 815 660 816
rect 806 820 812 821
rect 806 816 807 820
rect 811 816 812 820
rect 806 815 812 816
rect 950 820 956 821
rect 950 816 951 820
rect 955 816 956 820
rect 950 815 956 816
rect 1094 820 1100 821
rect 1094 816 1095 820
rect 1099 816 1100 820
rect 1094 815 1100 816
rect 1238 820 1244 821
rect 1238 816 1239 820
rect 1243 816 1244 820
rect 1238 815 1244 816
rect 1374 820 1380 821
rect 1374 816 1375 820
rect 1379 816 1380 820
rect 1374 815 1380 816
rect 1502 820 1508 821
rect 1502 816 1503 820
rect 1507 816 1508 820
rect 1502 815 1508 816
rect 1630 820 1636 821
rect 1630 816 1631 820
rect 1635 816 1636 820
rect 1630 815 1636 816
rect 1742 820 1748 821
rect 1742 816 1743 820
rect 1747 816 1748 820
rect 1830 819 1831 823
rect 1835 819 1836 823
rect 1830 818 1836 819
rect 1742 815 1748 816
rect 1902 802 1908 803
rect 1902 798 1903 802
rect 1907 798 1908 802
rect 1902 797 1908 798
rect 2014 802 2020 803
rect 2014 798 2015 802
rect 2019 798 2020 802
rect 2014 797 2020 798
rect 2166 802 2172 803
rect 2166 798 2167 802
rect 2171 798 2172 802
rect 2166 797 2172 798
rect 2326 802 2332 803
rect 2326 798 2327 802
rect 2331 798 2332 802
rect 2326 797 2332 798
rect 2486 802 2492 803
rect 2486 798 2487 802
rect 2491 798 2492 802
rect 2486 797 2492 798
rect 2646 802 2652 803
rect 2646 798 2647 802
rect 2651 798 2652 802
rect 2646 797 2652 798
rect 2806 802 2812 803
rect 2806 798 2807 802
rect 2811 798 2812 802
rect 2806 797 2812 798
rect 2958 802 2964 803
rect 2958 798 2959 802
rect 2963 798 2964 802
rect 2958 797 2964 798
rect 3102 802 3108 803
rect 3102 798 3103 802
rect 3107 798 3108 802
rect 3102 797 3108 798
rect 3246 802 3252 803
rect 3246 798 3247 802
rect 3251 798 3252 802
rect 3246 797 3252 798
rect 3390 802 3396 803
rect 3390 798 3391 802
rect 3395 798 3396 802
rect 3390 797 3396 798
rect 3510 802 3516 803
rect 3510 798 3511 802
rect 3515 798 3516 802
rect 3510 797 3516 798
rect 1870 784 1876 785
rect 1870 780 1871 784
rect 1875 780 1876 784
rect 1870 779 1876 780
rect 3590 784 3596 785
rect 3590 780 3591 784
rect 3595 780 3596 784
rect 3590 779 3596 780
rect 1870 767 1876 768
rect 134 764 140 765
rect 110 761 116 762
rect 110 757 111 761
rect 115 757 116 761
rect 134 760 135 764
rect 139 760 140 764
rect 134 759 140 760
rect 214 764 220 765
rect 214 760 215 764
rect 219 760 220 764
rect 214 759 220 760
rect 302 764 308 765
rect 302 760 303 764
rect 307 760 308 764
rect 302 759 308 760
rect 414 764 420 765
rect 414 760 415 764
rect 419 760 420 764
rect 414 759 420 760
rect 542 764 548 765
rect 542 760 543 764
rect 547 760 548 764
rect 542 759 548 760
rect 686 764 692 765
rect 686 760 687 764
rect 691 760 692 764
rect 686 759 692 760
rect 838 764 844 765
rect 838 760 839 764
rect 843 760 844 764
rect 838 759 844 760
rect 990 764 996 765
rect 990 760 991 764
rect 995 760 996 764
rect 990 759 996 760
rect 1142 764 1148 765
rect 1142 760 1143 764
rect 1147 760 1148 764
rect 1142 759 1148 760
rect 1294 764 1300 765
rect 1294 760 1295 764
rect 1299 760 1300 764
rect 1294 759 1300 760
rect 1446 764 1452 765
rect 1446 760 1447 764
rect 1451 760 1452 764
rect 1446 759 1452 760
rect 1606 764 1612 765
rect 1606 760 1607 764
rect 1611 760 1612 764
rect 1870 763 1871 767
rect 1875 763 1876 767
rect 3590 767 3596 768
rect 1870 762 1876 763
rect 1894 764 1900 765
rect 1606 759 1612 760
rect 1830 761 1836 762
rect 110 756 116 757
rect 1830 757 1831 761
rect 1835 757 1836 761
rect 1894 760 1895 764
rect 1899 760 1900 764
rect 1894 759 1900 760
rect 2006 764 2012 765
rect 2006 760 2007 764
rect 2011 760 2012 764
rect 2006 759 2012 760
rect 2158 764 2164 765
rect 2158 760 2159 764
rect 2163 760 2164 764
rect 2158 759 2164 760
rect 2318 764 2324 765
rect 2318 760 2319 764
rect 2323 760 2324 764
rect 2318 759 2324 760
rect 2478 764 2484 765
rect 2478 760 2479 764
rect 2483 760 2484 764
rect 2478 759 2484 760
rect 2638 764 2644 765
rect 2638 760 2639 764
rect 2643 760 2644 764
rect 2638 759 2644 760
rect 2798 764 2804 765
rect 2798 760 2799 764
rect 2803 760 2804 764
rect 2798 759 2804 760
rect 2950 764 2956 765
rect 2950 760 2951 764
rect 2955 760 2956 764
rect 2950 759 2956 760
rect 3094 764 3100 765
rect 3094 760 3095 764
rect 3099 760 3100 764
rect 3094 759 3100 760
rect 3238 764 3244 765
rect 3238 760 3239 764
rect 3243 760 3244 764
rect 3238 759 3244 760
rect 3382 764 3388 765
rect 3382 760 3383 764
rect 3387 760 3388 764
rect 3382 759 3388 760
rect 3502 764 3508 765
rect 3502 760 3503 764
rect 3507 760 3508 764
rect 3590 763 3591 767
rect 3595 763 3596 767
rect 3590 762 3596 763
rect 3502 759 3508 760
rect 1830 756 1836 757
rect 110 744 116 745
rect 110 740 111 744
rect 115 740 116 744
rect 110 739 116 740
rect 1830 744 1836 745
rect 1830 740 1831 744
rect 1835 740 1836 744
rect 1830 739 1836 740
rect 142 726 148 727
rect 142 722 143 726
rect 147 722 148 726
rect 142 721 148 722
rect 222 726 228 727
rect 222 722 223 726
rect 227 722 228 726
rect 222 721 228 722
rect 310 726 316 727
rect 310 722 311 726
rect 315 722 316 726
rect 310 721 316 722
rect 422 726 428 727
rect 422 722 423 726
rect 427 722 428 726
rect 422 721 428 722
rect 550 726 556 727
rect 550 722 551 726
rect 555 722 556 726
rect 550 721 556 722
rect 694 726 700 727
rect 694 722 695 726
rect 699 722 700 726
rect 694 721 700 722
rect 846 726 852 727
rect 846 722 847 726
rect 851 722 852 726
rect 846 721 852 722
rect 998 726 1004 727
rect 998 722 999 726
rect 1003 722 1004 726
rect 998 721 1004 722
rect 1150 726 1156 727
rect 1150 722 1151 726
rect 1155 722 1156 726
rect 1150 721 1156 722
rect 1302 726 1308 727
rect 1302 722 1303 726
rect 1307 722 1308 726
rect 1302 721 1308 722
rect 1454 726 1460 727
rect 1454 722 1455 726
rect 1459 722 1460 726
rect 1454 721 1460 722
rect 1614 726 1620 727
rect 1614 722 1615 726
rect 1619 722 1620 726
rect 1614 721 1620 722
rect 1966 720 1972 721
rect 1870 717 1876 718
rect 1870 713 1871 717
rect 1875 713 1876 717
rect 1966 716 1967 720
rect 1971 716 1972 720
rect 1966 715 1972 716
rect 2062 720 2068 721
rect 2062 716 2063 720
rect 2067 716 2068 720
rect 2062 715 2068 716
rect 2174 720 2180 721
rect 2174 716 2175 720
rect 2179 716 2180 720
rect 2174 715 2180 716
rect 2302 720 2308 721
rect 2302 716 2303 720
rect 2307 716 2308 720
rect 2302 715 2308 716
rect 2446 720 2452 721
rect 2446 716 2447 720
rect 2451 716 2452 720
rect 2446 715 2452 716
rect 2598 720 2604 721
rect 2598 716 2599 720
rect 2603 716 2604 720
rect 2598 715 2604 716
rect 2750 720 2756 721
rect 2750 716 2751 720
rect 2755 716 2756 720
rect 2750 715 2756 716
rect 2902 720 2908 721
rect 2902 716 2903 720
rect 2907 716 2908 720
rect 2902 715 2908 716
rect 3054 720 3060 721
rect 3054 716 3055 720
rect 3059 716 3060 720
rect 3054 715 3060 716
rect 3206 720 3212 721
rect 3206 716 3207 720
rect 3211 716 3212 720
rect 3206 715 3212 716
rect 3358 720 3364 721
rect 3358 716 3359 720
rect 3363 716 3364 720
rect 3358 715 3364 716
rect 3502 720 3508 721
rect 3502 716 3503 720
rect 3507 716 3508 720
rect 3502 715 3508 716
rect 3590 717 3596 718
rect 1870 712 1876 713
rect 3590 713 3591 717
rect 3595 713 3596 717
rect 3590 712 3596 713
rect 1870 700 1876 701
rect 1870 696 1871 700
rect 1875 696 1876 700
rect 1870 695 1876 696
rect 3590 700 3596 701
rect 3590 696 3591 700
rect 3595 696 3596 700
rect 3590 695 3596 696
rect 230 686 236 687
rect 230 682 231 686
rect 235 682 236 686
rect 230 681 236 682
rect 318 686 324 687
rect 318 682 319 686
rect 323 682 324 686
rect 318 681 324 682
rect 422 686 428 687
rect 422 682 423 686
rect 427 682 428 686
rect 422 681 428 682
rect 542 686 548 687
rect 542 682 543 686
rect 547 682 548 686
rect 542 681 548 682
rect 678 686 684 687
rect 678 682 679 686
rect 683 682 684 686
rect 678 681 684 682
rect 814 686 820 687
rect 814 682 815 686
rect 819 682 820 686
rect 814 681 820 682
rect 950 686 956 687
rect 950 682 951 686
rect 955 682 956 686
rect 950 681 956 682
rect 1086 686 1092 687
rect 1086 682 1087 686
rect 1091 682 1092 686
rect 1086 681 1092 682
rect 1214 686 1220 687
rect 1214 682 1215 686
rect 1219 682 1220 686
rect 1214 681 1220 682
rect 1334 686 1340 687
rect 1334 682 1335 686
rect 1339 682 1340 686
rect 1334 681 1340 682
rect 1454 686 1460 687
rect 1454 682 1455 686
rect 1459 682 1460 686
rect 1454 681 1460 682
rect 1582 686 1588 687
rect 1582 682 1583 686
rect 1587 682 1588 686
rect 1582 681 1588 682
rect 1974 682 1980 683
rect 1974 678 1975 682
rect 1979 678 1980 682
rect 1974 677 1980 678
rect 2070 682 2076 683
rect 2070 678 2071 682
rect 2075 678 2076 682
rect 2070 677 2076 678
rect 2182 682 2188 683
rect 2182 678 2183 682
rect 2187 678 2188 682
rect 2182 677 2188 678
rect 2310 682 2316 683
rect 2310 678 2311 682
rect 2315 678 2316 682
rect 2310 677 2316 678
rect 2454 682 2460 683
rect 2454 678 2455 682
rect 2459 678 2460 682
rect 2454 677 2460 678
rect 2606 682 2612 683
rect 2606 678 2607 682
rect 2611 678 2612 682
rect 2606 677 2612 678
rect 2758 682 2764 683
rect 2758 678 2759 682
rect 2763 678 2764 682
rect 2758 677 2764 678
rect 2910 682 2916 683
rect 2910 678 2911 682
rect 2915 678 2916 682
rect 2910 677 2916 678
rect 3062 682 3068 683
rect 3062 678 3063 682
rect 3067 678 3068 682
rect 3062 677 3068 678
rect 3214 682 3220 683
rect 3214 678 3215 682
rect 3219 678 3220 682
rect 3214 677 3220 678
rect 3366 682 3372 683
rect 3366 678 3367 682
rect 3371 678 3372 682
rect 3366 677 3372 678
rect 3510 682 3516 683
rect 3510 678 3511 682
rect 3515 678 3516 682
rect 3510 677 3516 678
rect 110 668 116 669
rect 110 664 111 668
rect 115 664 116 668
rect 110 663 116 664
rect 1830 668 1836 669
rect 1830 664 1831 668
rect 1835 664 1836 668
rect 1830 663 1836 664
rect 110 651 116 652
rect 110 647 111 651
rect 115 647 116 651
rect 1830 651 1836 652
rect 110 646 116 647
rect 222 648 228 649
rect 222 644 223 648
rect 227 644 228 648
rect 222 643 228 644
rect 310 648 316 649
rect 310 644 311 648
rect 315 644 316 648
rect 310 643 316 644
rect 414 648 420 649
rect 414 644 415 648
rect 419 644 420 648
rect 414 643 420 644
rect 534 648 540 649
rect 534 644 535 648
rect 539 644 540 648
rect 534 643 540 644
rect 670 648 676 649
rect 670 644 671 648
rect 675 644 676 648
rect 670 643 676 644
rect 806 648 812 649
rect 806 644 807 648
rect 811 644 812 648
rect 806 643 812 644
rect 942 648 948 649
rect 942 644 943 648
rect 947 644 948 648
rect 942 643 948 644
rect 1078 648 1084 649
rect 1078 644 1079 648
rect 1083 644 1084 648
rect 1078 643 1084 644
rect 1206 648 1212 649
rect 1206 644 1207 648
rect 1211 644 1212 648
rect 1206 643 1212 644
rect 1326 648 1332 649
rect 1326 644 1327 648
rect 1331 644 1332 648
rect 1326 643 1332 644
rect 1446 648 1452 649
rect 1446 644 1447 648
rect 1451 644 1452 648
rect 1446 643 1452 644
rect 1574 648 1580 649
rect 1574 644 1575 648
rect 1579 644 1580 648
rect 1830 647 1831 651
rect 1835 647 1836 651
rect 1830 646 1836 647
rect 2174 650 2180 651
rect 2174 646 2175 650
rect 2179 646 2180 650
rect 2174 645 2180 646
rect 2270 650 2276 651
rect 2270 646 2271 650
rect 2275 646 2276 650
rect 2270 645 2276 646
rect 2374 650 2380 651
rect 2374 646 2375 650
rect 2379 646 2380 650
rect 2374 645 2380 646
rect 2486 650 2492 651
rect 2486 646 2487 650
rect 2491 646 2492 650
rect 2486 645 2492 646
rect 2606 650 2612 651
rect 2606 646 2607 650
rect 2611 646 2612 650
rect 2606 645 2612 646
rect 2734 650 2740 651
rect 2734 646 2735 650
rect 2739 646 2740 650
rect 2734 645 2740 646
rect 2862 650 2868 651
rect 2862 646 2863 650
rect 2867 646 2868 650
rect 2862 645 2868 646
rect 2990 650 2996 651
rect 2990 646 2991 650
rect 2995 646 2996 650
rect 2990 645 2996 646
rect 3118 650 3124 651
rect 3118 646 3119 650
rect 3123 646 3124 650
rect 3118 645 3124 646
rect 3246 650 3252 651
rect 3246 646 3247 650
rect 3251 646 3252 650
rect 3246 645 3252 646
rect 3374 650 3380 651
rect 3374 646 3375 650
rect 3379 646 3380 650
rect 3374 645 3380 646
rect 3510 650 3516 651
rect 3510 646 3511 650
rect 3515 646 3516 650
rect 3510 645 3516 646
rect 1574 643 1580 644
rect 1870 632 1876 633
rect 1870 628 1871 632
rect 1875 628 1876 632
rect 1870 627 1876 628
rect 3590 632 3596 633
rect 3590 628 3591 632
rect 3595 628 3596 632
rect 3590 627 3596 628
rect 1870 615 1876 616
rect 1870 611 1871 615
rect 1875 611 1876 615
rect 3590 615 3596 616
rect 1870 610 1876 611
rect 2166 612 2172 613
rect 2166 608 2167 612
rect 2171 608 2172 612
rect 2166 607 2172 608
rect 2262 612 2268 613
rect 2262 608 2263 612
rect 2267 608 2268 612
rect 2262 607 2268 608
rect 2366 612 2372 613
rect 2366 608 2367 612
rect 2371 608 2372 612
rect 2366 607 2372 608
rect 2478 612 2484 613
rect 2478 608 2479 612
rect 2483 608 2484 612
rect 2478 607 2484 608
rect 2598 612 2604 613
rect 2598 608 2599 612
rect 2603 608 2604 612
rect 2598 607 2604 608
rect 2726 612 2732 613
rect 2726 608 2727 612
rect 2731 608 2732 612
rect 2726 607 2732 608
rect 2854 612 2860 613
rect 2854 608 2855 612
rect 2859 608 2860 612
rect 2854 607 2860 608
rect 2982 612 2988 613
rect 2982 608 2983 612
rect 2987 608 2988 612
rect 2982 607 2988 608
rect 3110 612 3116 613
rect 3110 608 3111 612
rect 3115 608 3116 612
rect 3110 607 3116 608
rect 3238 612 3244 613
rect 3238 608 3239 612
rect 3243 608 3244 612
rect 3238 607 3244 608
rect 3366 612 3372 613
rect 3366 608 3367 612
rect 3371 608 3372 612
rect 3366 607 3372 608
rect 3502 612 3508 613
rect 3502 608 3503 612
rect 3507 608 3508 612
rect 3590 611 3591 615
rect 3595 611 3596 615
rect 3590 610 3596 611
rect 3502 607 3508 608
rect 446 596 452 597
rect 110 593 116 594
rect 110 589 111 593
rect 115 589 116 593
rect 446 592 447 596
rect 451 592 452 596
rect 446 591 452 592
rect 526 596 532 597
rect 526 592 527 596
rect 531 592 532 596
rect 526 591 532 592
rect 606 596 612 597
rect 606 592 607 596
rect 611 592 612 596
rect 606 591 612 592
rect 686 596 692 597
rect 686 592 687 596
rect 691 592 692 596
rect 686 591 692 592
rect 774 596 780 597
rect 774 592 775 596
rect 779 592 780 596
rect 774 591 780 592
rect 870 596 876 597
rect 870 592 871 596
rect 875 592 876 596
rect 870 591 876 592
rect 958 596 964 597
rect 958 592 959 596
rect 963 592 964 596
rect 958 591 964 592
rect 1046 596 1052 597
rect 1046 592 1047 596
rect 1051 592 1052 596
rect 1046 591 1052 592
rect 1142 596 1148 597
rect 1142 592 1143 596
rect 1147 592 1148 596
rect 1142 591 1148 592
rect 1238 596 1244 597
rect 1238 592 1239 596
rect 1243 592 1244 596
rect 1238 591 1244 592
rect 1334 596 1340 597
rect 1334 592 1335 596
rect 1339 592 1340 596
rect 1334 591 1340 592
rect 1430 596 1436 597
rect 1430 592 1431 596
rect 1435 592 1436 596
rect 1430 591 1436 592
rect 1830 593 1836 594
rect 110 588 116 589
rect 1830 589 1831 593
rect 1835 589 1836 593
rect 1830 588 1836 589
rect 110 576 116 577
rect 110 572 111 576
rect 115 572 116 576
rect 110 571 116 572
rect 1830 576 1836 577
rect 1830 572 1831 576
rect 1835 572 1836 576
rect 1830 571 1836 572
rect 2262 568 2268 569
rect 1870 565 1876 566
rect 1870 561 1871 565
rect 1875 561 1876 565
rect 2262 564 2263 568
rect 2267 564 2268 568
rect 2262 563 2268 564
rect 2342 568 2348 569
rect 2342 564 2343 568
rect 2347 564 2348 568
rect 2342 563 2348 564
rect 2422 568 2428 569
rect 2422 564 2423 568
rect 2427 564 2428 568
rect 2422 563 2428 564
rect 2502 568 2508 569
rect 2502 564 2503 568
rect 2507 564 2508 568
rect 2502 563 2508 564
rect 2590 568 2596 569
rect 2590 564 2591 568
rect 2595 564 2596 568
rect 2590 563 2596 564
rect 2694 568 2700 569
rect 2694 564 2695 568
rect 2699 564 2700 568
rect 2694 563 2700 564
rect 2814 568 2820 569
rect 2814 564 2815 568
rect 2819 564 2820 568
rect 2814 563 2820 564
rect 2958 568 2964 569
rect 2958 564 2959 568
rect 2963 564 2964 568
rect 2958 563 2964 564
rect 3110 568 3116 569
rect 3110 564 3111 568
rect 3115 564 3116 568
rect 3110 563 3116 564
rect 3278 568 3284 569
rect 3278 564 3279 568
rect 3283 564 3284 568
rect 3278 563 3284 564
rect 3446 568 3452 569
rect 3446 564 3447 568
rect 3451 564 3452 568
rect 3446 563 3452 564
rect 3590 565 3596 566
rect 1870 560 1876 561
rect 3590 561 3591 565
rect 3595 561 3596 565
rect 3590 560 3596 561
rect 454 558 460 559
rect 454 554 455 558
rect 459 554 460 558
rect 454 553 460 554
rect 534 558 540 559
rect 534 554 535 558
rect 539 554 540 558
rect 534 553 540 554
rect 614 558 620 559
rect 614 554 615 558
rect 619 554 620 558
rect 614 553 620 554
rect 694 558 700 559
rect 694 554 695 558
rect 699 554 700 558
rect 694 553 700 554
rect 782 558 788 559
rect 782 554 783 558
rect 787 554 788 558
rect 782 553 788 554
rect 878 558 884 559
rect 878 554 879 558
rect 883 554 884 558
rect 878 553 884 554
rect 966 558 972 559
rect 966 554 967 558
rect 971 554 972 558
rect 966 553 972 554
rect 1054 558 1060 559
rect 1054 554 1055 558
rect 1059 554 1060 558
rect 1054 553 1060 554
rect 1150 558 1156 559
rect 1150 554 1151 558
rect 1155 554 1156 558
rect 1150 553 1156 554
rect 1246 558 1252 559
rect 1246 554 1247 558
rect 1251 554 1252 558
rect 1246 553 1252 554
rect 1342 558 1348 559
rect 1342 554 1343 558
rect 1347 554 1348 558
rect 1342 553 1348 554
rect 1438 558 1444 559
rect 1438 554 1439 558
rect 1443 554 1444 558
rect 1438 553 1444 554
rect 1870 548 1876 549
rect 1870 544 1871 548
rect 1875 544 1876 548
rect 1870 543 1876 544
rect 3590 548 3596 549
rect 3590 544 3591 548
rect 3595 544 3596 548
rect 3590 543 3596 544
rect 2270 530 2276 531
rect 2270 526 2271 530
rect 2275 526 2276 530
rect 2270 525 2276 526
rect 2350 530 2356 531
rect 2350 526 2351 530
rect 2355 526 2356 530
rect 2350 525 2356 526
rect 2430 530 2436 531
rect 2430 526 2431 530
rect 2435 526 2436 530
rect 2430 525 2436 526
rect 2510 530 2516 531
rect 2510 526 2511 530
rect 2515 526 2516 530
rect 2510 525 2516 526
rect 2598 530 2604 531
rect 2598 526 2599 530
rect 2603 526 2604 530
rect 2598 525 2604 526
rect 2702 530 2708 531
rect 2702 526 2703 530
rect 2707 526 2708 530
rect 2702 525 2708 526
rect 2822 530 2828 531
rect 2822 526 2823 530
rect 2827 526 2828 530
rect 2822 525 2828 526
rect 2966 530 2972 531
rect 2966 526 2967 530
rect 2971 526 2972 530
rect 2966 525 2972 526
rect 3118 530 3124 531
rect 3118 526 3119 530
rect 3123 526 3124 530
rect 3118 525 3124 526
rect 3286 530 3292 531
rect 3286 526 3287 530
rect 3291 526 3292 530
rect 3286 525 3292 526
rect 3454 530 3460 531
rect 3454 526 3455 530
rect 3459 526 3460 530
rect 3454 525 3460 526
rect 334 514 340 515
rect 334 510 335 514
rect 339 510 340 514
rect 334 509 340 510
rect 422 514 428 515
rect 422 510 423 514
rect 427 510 428 514
rect 422 509 428 510
rect 510 514 516 515
rect 510 510 511 514
rect 515 510 516 514
rect 510 509 516 510
rect 590 514 596 515
rect 590 510 591 514
rect 595 510 596 514
rect 590 509 596 510
rect 670 514 676 515
rect 670 510 671 514
rect 675 510 676 514
rect 670 509 676 510
rect 750 514 756 515
rect 750 510 751 514
rect 755 510 756 514
rect 750 509 756 510
rect 838 514 844 515
rect 838 510 839 514
rect 843 510 844 514
rect 838 509 844 510
rect 926 514 932 515
rect 926 510 927 514
rect 931 510 932 514
rect 926 509 932 510
rect 1014 514 1020 515
rect 1014 510 1015 514
rect 1019 510 1020 514
rect 1014 509 1020 510
rect 1102 514 1108 515
rect 1102 510 1103 514
rect 1107 510 1108 514
rect 1102 509 1108 510
rect 1190 514 1196 515
rect 1190 510 1191 514
rect 1195 510 1196 514
rect 1190 509 1196 510
rect 1278 514 1284 515
rect 1278 510 1279 514
rect 1283 510 1284 514
rect 1278 509 1284 510
rect 110 496 116 497
rect 110 492 111 496
rect 115 492 116 496
rect 110 491 116 492
rect 1830 496 1836 497
rect 1830 492 1831 496
rect 1835 492 1836 496
rect 1830 491 1836 492
rect 2190 490 2196 491
rect 2190 486 2191 490
rect 2195 486 2196 490
rect 2190 485 2196 486
rect 2286 490 2292 491
rect 2286 486 2287 490
rect 2291 486 2292 490
rect 2286 485 2292 486
rect 2382 490 2388 491
rect 2382 486 2383 490
rect 2387 486 2388 490
rect 2382 485 2388 486
rect 2486 490 2492 491
rect 2486 486 2487 490
rect 2491 486 2492 490
rect 2486 485 2492 486
rect 2582 490 2588 491
rect 2582 486 2583 490
rect 2587 486 2588 490
rect 2582 485 2588 486
rect 2686 490 2692 491
rect 2686 486 2687 490
rect 2691 486 2692 490
rect 2686 485 2692 486
rect 2790 490 2796 491
rect 2790 486 2791 490
rect 2795 486 2796 490
rect 2790 485 2796 486
rect 2910 490 2916 491
rect 2910 486 2911 490
rect 2915 486 2916 490
rect 2910 485 2916 486
rect 3038 490 3044 491
rect 3038 486 3039 490
rect 3043 486 3044 490
rect 3038 485 3044 486
rect 3174 490 3180 491
rect 3174 486 3175 490
rect 3179 486 3180 490
rect 3174 485 3180 486
rect 3318 490 3324 491
rect 3318 486 3319 490
rect 3323 486 3324 490
rect 3318 485 3324 486
rect 3470 490 3476 491
rect 3470 486 3471 490
rect 3475 486 3476 490
rect 3470 485 3476 486
rect 110 479 116 480
rect 110 475 111 479
rect 115 475 116 479
rect 1830 479 1836 480
rect 110 474 116 475
rect 326 476 332 477
rect 326 472 327 476
rect 331 472 332 476
rect 326 471 332 472
rect 414 476 420 477
rect 414 472 415 476
rect 419 472 420 476
rect 414 471 420 472
rect 502 476 508 477
rect 502 472 503 476
rect 507 472 508 476
rect 502 471 508 472
rect 582 476 588 477
rect 582 472 583 476
rect 587 472 588 476
rect 582 471 588 472
rect 662 476 668 477
rect 662 472 663 476
rect 667 472 668 476
rect 662 471 668 472
rect 742 476 748 477
rect 742 472 743 476
rect 747 472 748 476
rect 742 471 748 472
rect 830 476 836 477
rect 830 472 831 476
rect 835 472 836 476
rect 830 471 836 472
rect 918 476 924 477
rect 918 472 919 476
rect 923 472 924 476
rect 918 471 924 472
rect 1006 476 1012 477
rect 1006 472 1007 476
rect 1011 472 1012 476
rect 1006 471 1012 472
rect 1094 476 1100 477
rect 1094 472 1095 476
rect 1099 472 1100 476
rect 1094 471 1100 472
rect 1182 476 1188 477
rect 1182 472 1183 476
rect 1187 472 1188 476
rect 1182 471 1188 472
rect 1270 476 1276 477
rect 1270 472 1271 476
rect 1275 472 1276 476
rect 1830 475 1831 479
rect 1835 475 1836 479
rect 1830 474 1836 475
rect 1270 471 1276 472
rect 1870 472 1876 473
rect 1870 468 1871 472
rect 1875 468 1876 472
rect 1870 467 1876 468
rect 3590 472 3596 473
rect 3590 468 3591 472
rect 3595 468 3596 472
rect 3590 467 3596 468
rect 1870 455 1876 456
rect 1870 451 1871 455
rect 1875 451 1876 455
rect 3590 455 3596 456
rect 1870 450 1876 451
rect 2182 452 2188 453
rect 2182 448 2183 452
rect 2187 448 2188 452
rect 2182 447 2188 448
rect 2278 452 2284 453
rect 2278 448 2279 452
rect 2283 448 2284 452
rect 2278 447 2284 448
rect 2374 452 2380 453
rect 2374 448 2375 452
rect 2379 448 2380 452
rect 2374 447 2380 448
rect 2478 452 2484 453
rect 2478 448 2479 452
rect 2483 448 2484 452
rect 2478 447 2484 448
rect 2574 452 2580 453
rect 2574 448 2575 452
rect 2579 448 2580 452
rect 2574 447 2580 448
rect 2678 452 2684 453
rect 2678 448 2679 452
rect 2683 448 2684 452
rect 2678 447 2684 448
rect 2782 452 2788 453
rect 2782 448 2783 452
rect 2787 448 2788 452
rect 2782 447 2788 448
rect 2902 452 2908 453
rect 2902 448 2903 452
rect 2907 448 2908 452
rect 2902 447 2908 448
rect 3030 452 3036 453
rect 3030 448 3031 452
rect 3035 448 3036 452
rect 3030 447 3036 448
rect 3166 452 3172 453
rect 3166 448 3167 452
rect 3171 448 3172 452
rect 3166 447 3172 448
rect 3310 452 3316 453
rect 3310 448 3311 452
rect 3315 448 3316 452
rect 3310 447 3316 448
rect 3462 452 3468 453
rect 3462 448 3463 452
rect 3467 448 3468 452
rect 3590 451 3591 455
rect 3595 451 3596 455
rect 3590 450 3596 451
rect 3462 447 3468 448
rect 222 424 228 425
rect 110 421 116 422
rect 110 417 111 421
rect 115 417 116 421
rect 222 420 223 424
rect 227 420 228 424
rect 222 419 228 420
rect 334 424 340 425
rect 334 420 335 424
rect 339 420 340 424
rect 334 419 340 420
rect 446 424 452 425
rect 446 420 447 424
rect 451 420 452 424
rect 446 419 452 420
rect 558 424 564 425
rect 558 420 559 424
rect 563 420 564 424
rect 558 419 564 420
rect 662 424 668 425
rect 662 420 663 424
rect 667 420 668 424
rect 662 419 668 420
rect 758 424 764 425
rect 758 420 759 424
rect 763 420 764 424
rect 758 419 764 420
rect 846 424 852 425
rect 846 420 847 424
rect 851 420 852 424
rect 846 419 852 420
rect 934 424 940 425
rect 934 420 935 424
rect 939 420 940 424
rect 934 419 940 420
rect 1022 424 1028 425
rect 1022 420 1023 424
rect 1027 420 1028 424
rect 1022 419 1028 420
rect 1110 424 1116 425
rect 1110 420 1111 424
rect 1115 420 1116 424
rect 1110 419 1116 420
rect 1198 424 1204 425
rect 1198 420 1199 424
rect 1203 420 1204 424
rect 1198 419 1204 420
rect 1294 424 1300 425
rect 1294 420 1295 424
rect 1299 420 1300 424
rect 1294 419 1300 420
rect 1830 421 1836 422
rect 110 416 116 417
rect 1830 417 1831 421
rect 1835 417 1836 421
rect 1830 416 1836 417
rect 110 404 116 405
rect 110 400 111 404
rect 115 400 116 404
rect 110 399 116 400
rect 1830 404 1836 405
rect 1830 400 1831 404
rect 1835 400 1836 404
rect 1974 404 1980 405
rect 1830 399 1836 400
rect 1870 401 1876 402
rect 1870 397 1871 401
rect 1875 397 1876 401
rect 1974 400 1975 404
rect 1979 400 1980 404
rect 1974 399 1980 400
rect 2062 404 2068 405
rect 2062 400 2063 404
rect 2067 400 2068 404
rect 2062 399 2068 400
rect 2158 404 2164 405
rect 2158 400 2159 404
rect 2163 400 2164 404
rect 2158 399 2164 400
rect 2254 404 2260 405
rect 2254 400 2255 404
rect 2259 400 2260 404
rect 2254 399 2260 400
rect 2358 404 2364 405
rect 2358 400 2359 404
rect 2363 400 2364 404
rect 2358 399 2364 400
rect 2470 404 2476 405
rect 2470 400 2471 404
rect 2475 400 2476 404
rect 2470 399 2476 400
rect 2606 404 2612 405
rect 2606 400 2607 404
rect 2611 400 2612 404
rect 2606 399 2612 400
rect 2758 404 2764 405
rect 2758 400 2759 404
rect 2763 400 2764 404
rect 2758 399 2764 400
rect 2926 404 2932 405
rect 2926 400 2927 404
rect 2931 400 2932 404
rect 2926 399 2932 400
rect 3110 404 3116 405
rect 3110 400 3111 404
rect 3115 400 3116 404
rect 3110 399 3116 400
rect 3302 404 3308 405
rect 3302 400 3303 404
rect 3307 400 3308 404
rect 3302 399 3308 400
rect 3494 404 3500 405
rect 3494 400 3495 404
rect 3499 400 3500 404
rect 3494 399 3500 400
rect 3590 401 3596 402
rect 1870 396 1876 397
rect 3590 397 3591 401
rect 3595 397 3596 401
rect 3590 396 3596 397
rect 230 386 236 387
rect 230 382 231 386
rect 235 382 236 386
rect 230 381 236 382
rect 342 386 348 387
rect 342 382 343 386
rect 347 382 348 386
rect 342 381 348 382
rect 454 386 460 387
rect 454 382 455 386
rect 459 382 460 386
rect 454 381 460 382
rect 566 386 572 387
rect 566 382 567 386
rect 571 382 572 386
rect 566 381 572 382
rect 670 386 676 387
rect 670 382 671 386
rect 675 382 676 386
rect 670 381 676 382
rect 766 386 772 387
rect 766 382 767 386
rect 771 382 772 386
rect 766 381 772 382
rect 854 386 860 387
rect 854 382 855 386
rect 859 382 860 386
rect 854 381 860 382
rect 942 386 948 387
rect 942 382 943 386
rect 947 382 948 386
rect 942 381 948 382
rect 1030 386 1036 387
rect 1030 382 1031 386
rect 1035 382 1036 386
rect 1030 381 1036 382
rect 1118 386 1124 387
rect 1118 382 1119 386
rect 1123 382 1124 386
rect 1118 381 1124 382
rect 1206 386 1212 387
rect 1206 382 1207 386
rect 1211 382 1212 386
rect 1206 381 1212 382
rect 1302 386 1308 387
rect 1302 382 1303 386
rect 1307 382 1308 386
rect 1302 381 1308 382
rect 1870 384 1876 385
rect 1870 380 1871 384
rect 1875 380 1876 384
rect 1870 379 1876 380
rect 3590 384 3596 385
rect 3590 380 3591 384
rect 3595 380 3596 384
rect 3590 379 3596 380
rect 1982 366 1988 367
rect 1982 362 1983 366
rect 1987 362 1988 366
rect 1982 361 1988 362
rect 2070 366 2076 367
rect 2070 362 2071 366
rect 2075 362 2076 366
rect 2070 361 2076 362
rect 2166 366 2172 367
rect 2166 362 2167 366
rect 2171 362 2172 366
rect 2166 361 2172 362
rect 2262 366 2268 367
rect 2262 362 2263 366
rect 2267 362 2268 366
rect 2262 361 2268 362
rect 2366 366 2372 367
rect 2366 362 2367 366
rect 2371 362 2372 366
rect 2366 361 2372 362
rect 2478 366 2484 367
rect 2478 362 2479 366
rect 2483 362 2484 366
rect 2478 361 2484 362
rect 2614 366 2620 367
rect 2614 362 2615 366
rect 2619 362 2620 366
rect 2614 361 2620 362
rect 2766 366 2772 367
rect 2766 362 2767 366
rect 2771 362 2772 366
rect 2766 361 2772 362
rect 2934 366 2940 367
rect 2934 362 2935 366
rect 2939 362 2940 366
rect 2934 361 2940 362
rect 3118 366 3124 367
rect 3118 362 3119 366
rect 3123 362 3124 366
rect 3118 361 3124 362
rect 3310 366 3316 367
rect 3310 362 3311 366
rect 3315 362 3316 366
rect 3310 361 3316 362
rect 3502 366 3508 367
rect 3502 362 3503 366
rect 3507 362 3508 366
rect 3502 361 3508 362
rect 142 342 148 343
rect 142 338 143 342
rect 147 338 148 342
rect 142 337 148 338
rect 262 342 268 343
rect 262 338 263 342
rect 267 338 268 342
rect 262 337 268 338
rect 398 342 404 343
rect 398 338 399 342
rect 403 338 404 342
rect 398 337 404 338
rect 534 342 540 343
rect 534 338 535 342
rect 539 338 540 342
rect 534 337 540 338
rect 670 342 676 343
rect 670 338 671 342
rect 675 338 676 342
rect 670 337 676 338
rect 790 342 796 343
rect 790 338 791 342
rect 795 338 796 342
rect 790 337 796 338
rect 910 342 916 343
rect 910 338 911 342
rect 915 338 916 342
rect 910 337 916 338
rect 1022 342 1028 343
rect 1022 338 1023 342
rect 1027 338 1028 342
rect 1022 337 1028 338
rect 1126 342 1132 343
rect 1126 338 1127 342
rect 1131 338 1132 342
rect 1126 337 1132 338
rect 1230 342 1236 343
rect 1230 338 1231 342
rect 1235 338 1236 342
rect 1230 337 1236 338
rect 1334 342 1340 343
rect 1334 338 1335 342
rect 1339 338 1340 342
rect 1334 337 1340 338
rect 1438 342 1444 343
rect 1438 338 1439 342
rect 1443 338 1444 342
rect 1438 337 1444 338
rect 2214 330 2220 331
rect 2214 326 2215 330
rect 2219 326 2220 330
rect 2214 325 2220 326
rect 2294 330 2300 331
rect 2294 326 2295 330
rect 2299 326 2300 330
rect 2294 325 2300 326
rect 2382 330 2388 331
rect 2382 326 2383 330
rect 2387 326 2388 330
rect 2382 325 2388 326
rect 2478 330 2484 331
rect 2478 326 2479 330
rect 2483 326 2484 330
rect 2478 325 2484 326
rect 2590 330 2596 331
rect 2590 326 2591 330
rect 2595 326 2596 330
rect 2590 325 2596 326
rect 2718 330 2724 331
rect 2718 326 2719 330
rect 2723 326 2724 330
rect 2718 325 2724 326
rect 2846 330 2852 331
rect 2846 326 2847 330
rect 2851 326 2852 330
rect 2846 325 2852 326
rect 2982 330 2988 331
rect 2982 326 2983 330
rect 2987 326 2988 330
rect 2982 325 2988 326
rect 3118 330 3124 331
rect 3118 326 3119 330
rect 3123 326 3124 330
rect 3118 325 3124 326
rect 3254 330 3260 331
rect 3254 326 3255 330
rect 3259 326 3260 330
rect 3254 325 3260 326
rect 3390 330 3396 331
rect 3390 326 3391 330
rect 3395 326 3396 330
rect 3390 325 3396 326
rect 3510 330 3516 331
rect 3510 326 3511 330
rect 3515 326 3516 330
rect 3510 325 3516 326
rect 110 324 116 325
rect 110 320 111 324
rect 115 320 116 324
rect 110 319 116 320
rect 1830 324 1836 325
rect 1830 320 1831 324
rect 1835 320 1836 324
rect 1830 319 1836 320
rect 1870 312 1876 313
rect 1870 308 1871 312
rect 1875 308 1876 312
rect 110 307 116 308
rect 110 303 111 307
rect 115 303 116 307
rect 1830 307 1836 308
rect 1870 307 1876 308
rect 3590 312 3596 313
rect 3590 308 3591 312
rect 3595 308 3596 312
rect 3590 307 3596 308
rect 110 302 116 303
rect 134 304 140 305
rect 134 300 135 304
rect 139 300 140 304
rect 134 299 140 300
rect 254 304 260 305
rect 254 300 255 304
rect 259 300 260 304
rect 254 299 260 300
rect 390 304 396 305
rect 390 300 391 304
rect 395 300 396 304
rect 390 299 396 300
rect 526 304 532 305
rect 526 300 527 304
rect 531 300 532 304
rect 526 299 532 300
rect 662 304 668 305
rect 662 300 663 304
rect 667 300 668 304
rect 662 299 668 300
rect 782 304 788 305
rect 782 300 783 304
rect 787 300 788 304
rect 782 299 788 300
rect 902 304 908 305
rect 902 300 903 304
rect 907 300 908 304
rect 902 299 908 300
rect 1014 304 1020 305
rect 1014 300 1015 304
rect 1019 300 1020 304
rect 1014 299 1020 300
rect 1118 304 1124 305
rect 1118 300 1119 304
rect 1123 300 1124 304
rect 1118 299 1124 300
rect 1222 304 1228 305
rect 1222 300 1223 304
rect 1227 300 1228 304
rect 1222 299 1228 300
rect 1326 304 1332 305
rect 1326 300 1327 304
rect 1331 300 1332 304
rect 1326 299 1332 300
rect 1430 304 1436 305
rect 1430 300 1431 304
rect 1435 300 1436 304
rect 1830 303 1831 307
rect 1835 303 1836 307
rect 1830 302 1836 303
rect 1430 299 1436 300
rect 1870 295 1876 296
rect 1870 291 1871 295
rect 1875 291 1876 295
rect 3590 295 3596 296
rect 1870 290 1876 291
rect 2206 292 2212 293
rect 2206 288 2207 292
rect 2211 288 2212 292
rect 2206 287 2212 288
rect 2286 292 2292 293
rect 2286 288 2287 292
rect 2291 288 2292 292
rect 2286 287 2292 288
rect 2374 292 2380 293
rect 2374 288 2375 292
rect 2379 288 2380 292
rect 2374 287 2380 288
rect 2470 292 2476 293
rect 2470 288 2471 292
rect 2475 288 2476 292
rect 2470 287 2476 288
rect 2582 292 2588 293
rect 2582 288 2583 292
rect 2587 288 2588 292
rect 2582 287 2588 288
rect 2710 292 2716 293
rect 2710 288 2711 292
rect 2715 288 2716 292
rect 2710 287 2716 288
rect 2838 292 2844 293
rect 2838 288 2839 292
rect 2843 288 2844 292
rect 2838 287 2844 288
rect 2974 292 2980 293
rect 2974 288 2975 292
rect 2979 288 2980 292
rect 2974 287 2980 288
rect 3110 292 3116 293
rect 3110 288 3111 292
rect 3115 288 3116 292
rect 3110 287 3116 288
rect 3246 292 3252 293
rect 3246 288 3247 292
rect 3251 288 3252 292
rect 3246 287 3252 288
rect 3382 292 3388 293
rect 3382 288 3383 292
rect 3387 288 3388 292
rect 3382 287 3388 288
rect 3502 292 3508 293
rect 3502 288 3503 292
rect 3507 288 3508 292
rect 3590 291 3591 295
rect 3595 291 3596 295
rect 3590 290 3596 291
rect 3502 287 3508 288
rect 134 252 140 253
rect 110 249 116 250
rect 110 245 111 249
rect 115 245 116 249
rect 134 248 135 252
rect 139 248 140 252
rect 134 247 140 248
rect 246 252 252 253
rect 246 248 247 252
rect 251 248 252 252
rect 246 247 252 248
rect 390 252 396 253
rect 390 248 391 252
rect 395 248 396 252
rect 390 247 396 248
rect 542 252 548 253
rect 542 248 543 252
rect 547 248 548 252
rect 542 247 548 248
rect 694 252 700 253
rect 694 248 695 252
rect 699 248 700 252
rect 694 247 700 248
rect 846 252 852 253
rect 846 248 847 252
rect 851 248 852 252
rect 846 247 852 248
rect 990 252 996 253
rect 990 248 991 252
rect 995 248 996 252
rect 990 247 996 248
rect 1118 252 1124 253
rect 1118 248 1119 252
rect 1123 248 1124 252
rect 1118 247 1124 248
rect 1238 252 1244 253
rect 1238 248 1239 252
rect 1243 248 1244 252
rect 1238 247 1244 248
rect 1358 252 1364 253
rect 1358 248 1359 252
rect 1363 248 1364 252
rect 1358 247 1364 248
rect 1478 252 1484 253
rect 1478 248 1479 252
rect 1483 248 1484 252
rect 1478 247 1484 248
rect 1598 252 1604 253
rect 1598 248 1599 252
rect 1603 248 1604 252
rect 1598 247 1604 248
rect 1830 249 1836 250
rect 110 244 116 245
rect 1830 245 1831 249
rect 1835 245 1836 249
rect 1830 244 1836 245
rect 1990 244 1996 245
rect 1870 241 1876 242
rect 1870 237 1871 241
rect 1875 237 1876 241
rect 1990 240 1991 244
rect 1995 240 1996 244
rect 1990 239 1996 240
rect 2118 244 2124 245
rect 2118 240 2119 244
rect 2123 240 2124 244
rect 2118 239 2124 240
rect 2254 244 2260 245
rect 2254 240 2255 244
rect 2259 240 2260 244
rect 2254 239 2260 240
rect 2390 244 2396 245
rect 2390 240 2391 244
rect 2395 240 2396 244
rect 2390 239 2396 240
rect 2534 244 2540 245
rect 2534 240 2535 244
rect 2539 240 2540 244
rect 2534 239 2540 240
rect 2678 244 2684 245
rect 2678 240 2679 244
rect 2683 240 2684 244
rect 2678 239 2684 240
rect 2814 244 2820 245
rect 2814 240 2815 244
rect 2819 240 2820 244
rect 2814 239 2820 240
rect 2950 244 2956 245
rect 2950 240 2951 244
rect 2955 240 2956 244
rect 2950 239 2956 240
rect 3094 244 3100 245
rect 3094 240 3095 244
rect 3099 240 3100 244
rect 3094 239 3100 240
rect 3238 244 3244 245
rect 3238 240 3239 244
rect 3243 240 3244 244
rect 3238 239 3244 240
rect 3382 244 3388 245
rect 3382 240 3383 244
rect 3387 240 3388 244
rect 3382 239 3388 240
rect 3502 244 3508 245
rect 3502 240 3503 244
rect 3507 240 3508 244
rect 3502 239 3508 240
rect 3590 241 3596 242
rect 1870 236 1876 237
rect 3590 237 3591 241
rect 3595 237 3596 241
rect 3590 236 3596 237
rect 110 232 116 233
rect 110 228 111 232
rect 115 228 116 232
rect 110 227 116 228
rect 1830 232 1836 233
rect 1830 228 1831 232
rect 1835 228 1836 232
rect 1830 227 1836 228
rect 1870 224 1876 225
rect 1870 220 1871 224
rect 1875 220 1876 224
rect 1870 219 1876 220
rect 3590 224 3596 225
rect 3590 220 3591 224
rect 3595 220 3596 224
rect 3590 219 3596 220
rect 142 214 148 215
rect 142 210 143 214
rect 147 210 148 214
rect 142 209 148 210
rect 254 214 260 215
rect 254 210 255 214
rect 259 210 260 214
rect 254 209 260 210
rect 398 214 404 215
rect 398 210 399 214
rect 403 210 404 214
rect 398 209 404 210
rect 550 214 556 215
rect 550 210 551 214
rect 555 210 556 214
rect 550 209 556 210
rect 702 214 708 215
rect 702 210 703 214
rect 707 210 708 214
rect 702 209 708 210
rect 854 214 860 215
rect 854 210 855 214
rect 859 210 860 214
rect 854 209 860 210
rect 998 214 1004 215
rect 998 210 999 214
rect 1003 210 1004 214
rect 998 209 1004 210
rect 1126 214 1132 215
rect 1126 210 1127 214
rect 1131 210 1132 214
rect 1126 209 1132 210
rect 1246 214 1252 215
rect 1246 210 1247 214
rect 1251 210 1252 214
rect 1246 209 1252 210
rect 1366 214 1372 215
rect 1366 210 1367 214
rect 1371 210 1372 214
rect 1366 209 1372 210
rect 1486 214 1492 215
rect 1486 210 1487 214
rect 1491 210 1492 214
rect 1486 209 1492 210
rect 1606 214 1612 215
rect 1606 210 1607 214
rect 1611 210 1612 214
rect 1606 209 1612 210
rect 1998 206 2004 207
rect 1998 202 1999 206
rect 2003 202 2004 206
rect 1998 201 2004 202
rect 2126 206 2132 207
rect 2126 202 2127 206
rect 2131 202 2132 206
rect 2126 201 2132 202
rect 2262 206 2268 207
rect 2262 202 2263 206
rect 2267 202 2268 206
rect 2262 201 2268 202
rect 2398 206 2404 207
rect 2398 202 2399 206
rect 2403 202 2404 206
rect 2398 201 2404 202
rect 2542 206 2548 207
rect 2542 202 2543 206
rect 2547 202 2548 206
rect 2542 201 2548 202
rect 2686 206 2692 207
rect 2686 202 2687 206
rect 2691 202 2692 206
rect 2686 201 2692 202
rect 2822 206 2828 207
rect 2822 202 2823 206
rect 2827 202 2828 206
rect 2822 201 2828 202
rect 2958 206 2964 207
rect 2958 202 2959 206
rect 2963 202 2964 206
rect 2958 201 2964 202
rect 3102 206 3108 207
rect 3102 202 3103 206
rect 3107 202 3108 206
rect 3102 201 3108 202
rect 3246 206 3252 207
rect 3246 202 3247 206
rect 3251 202 3252 206
rect 3246 201 3252 202
rect 3390 206 3396 207
rect 3390 202 3391 206
rect 3395 202 3396 206
rect 3390 201 3396 202
rect 3510 206 3516 207
rect 3510 202 3511 206
rect 3515 202 3516 206
rect 3510 201 3516 202
rect 1902 162 1908 163
rect 1902 158 1903 162
rect 1907 158 1908 162
rect 1902 157 1908 158
rect 1982 162 1988 163
rect 1982 158 1983 162
rect 1987 158 1988 162
rect 1982 157 1988 158
rect 2086 162 2092 163
rect 2086 158 2087 162
rect 2091 158 2092 162
rect 2086 157 2092 158
rect 2214 162 2220 163
rect 2214 158 2215 162
rect 2219 158 2220 162
rect 2214 157 2220 158
rect 2350 162 2356 163
rect 2350 158 2351 162
rect 2355 158 2356 162
rect 2350 157 2356 158
rect 2486 162 2492 163
rect 2486 158 2487 162
rect 2491 158 2492 162
rect 2486 157 2492 158
rect 2622 162 2628 163
rect 2622 158 2623 162
rect 2627 158 2628 162
rect 2622 157 2628 158
rect 2742 162 2748 163
rect 2742 158 2743 162
rect 2747 158 2748 162
rect 2742 157 2748 158
rect 2854 162 2860 163
rect 2854 158 2855 162
rect 2859 158 2860 162
rect 2854 157 2860 158
rect 2958 162 2964 163
rect 2958 158 2959 162
rect 2963 158 2964 162
rect 2958 157 2964 158
rect 3062 162 3068 163
rect 3062 158 3063 162
rect 3067 158 3068 162
rect 3062 157 3068 158
rect 3158 162 3164 163
rect 3158 158 3159 162
rect 3163 158 3164 162
rect 3158 157 3164 158
rect 3246 162 3252 163
rect 3246 158 3247 162
rect 3251 158 3252 162
rect 3246 157 3252 158
rect 3342 162 3348 163
rect 3342 158 3343 162
rect 3347 158 3348 162
rect 3342 157 3348 158
rect 3430 162 3436 163
rect 3430 158 3431 162
rect 3435 158 3436 162
rect 3430 157 3436 158
rect 3510 162 3516 163
rect 3510 158 3511 162
rect 3515 158 3516 162
rect 3510 157 3516 158
rect 142 146 148 147
rect 142 142 143 146
rect 147 142 148 146
rect 142 141 148 142
rect 222 146 228 147
rect 222 142 223 146
rect 227 142 228 146
rect 222 141 228 142
rect 302 146 308 147
rect 302 142 303 146
rect 307 142 308 146
rect 302 141 308 142
rect 382 146 388 147
rect 382 142 383 146
rect 387 142 388 146
rect 382 141 388 142
rect 462 146 468 147
rect 462 142 463 146
rect 467 142 468 146
rect 462 141 468 142
rect 542 146 548 147
rect 542 142 543 146
rect 547 142 548 146
rect 542 141 548 142
rect 622 146 628 147
rect 622 142 623 146
rect 627 142 628 146
rect 622 141 628 142
rect 702 146 708 147
rect 702 142 703 146
rect 707 142 708 146
rect 702 141 708 142
rect 782 146 788 147
rect 782 142 783 146
rect 787 142 788 146
rect 782 141 788 142
rect 862 146 868 147
rect 862 142 863 146
rect 867 142 868 146
rect 862 141 868 142
rect 942 146 948 147
rect 942 142 943 146
rect 947 142 948 146
rect 942 141 948 142
rect 1022 146 1028 147
rect 1022 142 1023 146
rect 1027 142 1028 146
rect 1022 141 1028 142
rect 1102 146 1108 147
rect 1102 142 1103 146
rect 1107 142 1108 146
rect 1102 141 1108 142
rect 1182 146 1188 147
rect 1182 142 1183 146
rect 1187 142 1188 146
rect 1182 141 1188 142
rect 1262 146 1268 147
rect 1262 142 1263 146
rect 1267 142 1268 146
rect 1262 141 1268 142
rect 1342 146 1348 147
rect 1342 142 1343 146
rect 1347 142 1348 146
rect 1342 141 1348 142
rect 1422 146 1428 147
rect 1422 142 1423 146
rect 1427 142 1428 146
rect 1422 141 1428 142
rect 1510 146 1516 147
rect 1510 142 1511 146
rect 1515 142 1516 146
rect 1510 141 1516 142
rect 1590 146 1596 147
rect 1590 142 1591 146
rect 1595 142 1596 146
rect 1590 141 1596 142
rect 1670 146 1676 147
rect 1670 142 1671 146
rect 1675 142 1676 146
rect 1670 141 1676 142
rect 1750 146 1756 147
rect 1750 142 1751 146
rect 1755 142 1756 146
rect 1750 141 1756 142
rect 1870 144 1876 145
rect 1870 140 1871 144
rect 1875 140 1876 144
rect 1870 139 1876 140
rect 3590 144 3596 145
rect 3590 140 3591 144
rect 3595 140 3596 144
rect 3590 139 3596 140
rect 110 128 116 129
rect 110 124 111 128
rect 115 124 116 128
rect 110 123 116 124
rect 1830 128 1836 129
rect 1830 124 1831 128
rect 1835 124 1836 128
rect 1830 123 1836 124
rect 1870 127 1876 128
rect 1870 123 1871 127
rect 1875 123 1876 127
rect 3590 127 3596 128
rect 1870 122 1876 123
rect 1894 124 1900 125
rect 1894 120 1895 124
rect 1899 120 1900 124
rect 1894 119 1900 120
rect 1974 124 1980 125
rect 1974 120 1975 124
rect 1979 120 1980 124
rect 1974 119 1980 120
rect 2078 124 2084 125
rect 2078 120 2079 124
rect 2083 120 2084 124
rect 2078 119 2084 120
rect 2206 124 2212 125
rect 2206 120 2207 124
rect 2211 120 2212 124
rect 2206 119 2212 120
rect 2342 124 2348 125
rect 2342 120 2343 124
rect 2347 120 2348 124
rect 2342 119 2348 120
rect 2478 124 2484 125
rect 2478 120 2479 124
rect 2483 120 2484 124
rect 2478 119 2484 120
rect 2614 124 2620 125
rect 2614 120 2615 124
rect 2619 120 2620 124
rect 2614 119 2620 120
rect 2734 124 2740 125
rect 2734 120 2735 124
rect 2739 120 2740 124
rect 2734 119 2740 120
rect 2846 124 2852 125
rect 2846 120 2847 124
rect 2851 120 2852 124
rect 2846 119 2852 120
rect 2950 124 2956 125
rect 2950 120 2951 124
rect 2955 120 2956 124
rect 2950 119 2956 120
rect 3054 124 3060 125
rect 3054 120 3055 124
rect 3059 120 3060 124
rect 3054 119 3060 120
rect 3150 124 3156 125
rect 3150 120 3151 124
rect 3155 120 3156 124
rect 3150 119 3156 120
rect 3238 124 3244 125
rect 3238 120 3239 124
rect 3243 120 3244 124
rect 3238 119 3244 120
rect 3334 124 3340 125
rect 3334 120 3335 124
rect 3339 120 3340 124
rect 3334 119 3340 120
rect 3422 124 3428 125
rect 3422 120 3423 124
rect 3427 120 3428 124
rect 3422 119 3428 120
rect 3502 124 3508 125
rect 3502 120 3503 124
rect 3507 120 3508 124
rect 3590 123 3591 127
rect 3595 123 3596 127
rect 3590 122 3596 123
rect 3502 119 3508 120
rect 110 111 116 112
rect 110 107 111 111
rect 115 107 116 111
rect 1830 111 1836 112
rect 110 106 116 107
rect 134 108 140 109
rect 134 104 135 108
rect 139 104 140 108
rect 134 103 140 104
rect 214 108 220 109
rect 214 104 215 108
rect 219 104 220 108
rect 214 103 220 104
rect 294 108 300 109
rect 294 104 295 108
rect 299 104 300 108
rect 294 103 300 104
rect 374 108 380 109
rect 374 104 375 108
rect 379 104 380 108
rect 374 103 380 104
rect 454 108 460 109
rect 454 104 455 108
rect 459 104 460 108
rect 454 103 460 104
rect 534 108 540 109
rect 534 104 535 108
rect 539 104 540 108
rect 534 103 540 104
rect 614 108 620 109
rect 614 104 615 108
rect 619 104 620 108
rect 614 103 620 104
rect 694 108 700 109
rect 694 104 695 108
rect 699 104 700 108
rect 694 103 700 104
rect 774 108 780 109
rect 774 104 775 108
rect 779 104 780 108
rect 774 103 780 104
rect 854 108 860 109
rect 854 104 855 108
rect 859 104 860 108
rect 854 103 860 104
rect 934 108 940 109
rect 934 104 935 108
rect 939 104 940 108
rect 934 103 940 104
rect 1014 108 1020 109
rect 1014 104 1015 108
rect 1019 104 1020 108
rect 1014 103 1020 104
rect 1094 108 1100 109
rect 1094 104 1095 108
rect 1099 104 1100 108
rect 1094 103 1100 104
rect 1174 108 1180 109
rect 1174 104 1175 108
rect 1179 104 1180 108
rect 1174 103 1180 104
rect 1254 108 1260 109
rect 1254 104 1255 108
rect 1259 104 1260 108
rect 1254 103 1260 104
rect 1334 108 1340 109
rect 1334 104 1335 108
rect 1339 104 1340 108
rect 1334 103 1340 104
rect 1414 108 1420 109
rect 1414 104 1415 108
rect 1419 104 1420 108
rect 1414 103 1420 104
rect 1502 108 1508 109
rect 1502 104 1503 108
rect 1507 104 1508 108
rect 1502 103 1508 104
rect 1582 108 1588 109
rect 1582 104 1583 108
rect 1587 104 1588 108
rect 1582 103 1588 104
rect 1662 108 1668 109
rect 1662 104 1663 108
rect 1667 104 1668 108
rect 1662 103 1668 104
rect 1742 108 1748 109
rect 1742 104 1743 108
rect 1747 104 1748 108
rect 1830 107 1831 111
rect 1835 107 1836 111
rect 1830 106 1836 107
rect 1742 103 1748 104
<< m3c >>
rect 111 3641 115 3645
rect 135 3644 139 3648
rect 215 3644 219 3648
rect 295 3644 299 3648
rect 1831 3641 1835 3645
rect 111 3624 115 3628
rect 1831 3624 1835 3628
rect 143 3606 147 3610
rect 223 3606 227 3610
rect 303 3606 307 3610
rect 2063 3582 2067 3586
rect 2151 3582 2155 3586
rect 2255 3582 2259 3586
rect 2367 3582 2371 3586
rect 2479 3582 2483 3586
rect 2591 3582 2595 3586
rect 2703 3582 2707 3586
rect 2815 3582 2819 3586
rect 2919 3582 2923 3586
rect 3015 3582 3019 3586
rect 3111 3582 3115 3586
rect 3207 3582 3211 3586
rect 3303 3582 3307 3586
rect 3399 3582 3403 3586
rect 143 3574 147 3578
rect 223 3574 227 3578
rect 343 3574 347 3578
rect 471 3574 475 3578
rect 607 3574 611 3578
rect 743 3574 747 3578
rect 879 3574 883 3578
rect 999 3574 1003 3578
rect 1111 3574 1115 3578
rect 1223 3574 1227 3578
rect 1327 3574 1331 3578
rect 1423 3574 1427 3578
rect 1527 3574 1531 3578
rect 1631 3574 1635 3578
rect 1871 3564 1875 3568
rect 3591 3564 3595 3568
rect 111 3556 115 3560
rect 1831 3556 1835 3560
rect 1871 3547 1875 3551
rect 2055 3544 2059 3548
rect 111 3539 115 3543
rect 2143 3544 2147 3548
rect 2247 3544 2251 3548
rect 2359 3544 2363 3548
rect 2471 3544 2475 3548
rect 2583 3544 2587 3548
rect 2695 3544 2699 3548
rect 2807 3544 2811 3548
rect 2911 3544 2915 3548
rect 3007 3544 3011 3548
rect 3103 3544 3107 3548
rect 3199 3544 3203 3548
rect 3295 3544 3299 3548
rect 3391 3544 3395 3548
rect 3591 3547 3595 3551
rect 135 3536 139 3540
rect 215 3536 219 3540
rect 335 3536 339 3540
rect 463 3536 467 3540
rect 599 3536 603 3540
rect 735 3536 739 3540
rect 871 3536 875 3540
rect 991 3536 995 3540
rect 1103 3536 1107 3540
rect 1215 3536 1219 3540
rect 1319 3536 1323 3540
rect 1415 3536 1419 3540
rect 1519 3536 1523 3540
rect 1623 3536 1627 3540
rect 1831 3539 1835 3543
rect 1871 3497 1875 3501
rect 2087 3500 2091 3504
rect 2167 3500 2171 3504
rect 2263 3500 2267 3504
rect 2367 3500 2371 3504
rect 2487 3500 2491 3504
rect 2615 3500 2619 3504
rect 2743 3500 2747 3504
rect 2871 3500 2875 3504
rect 2991 3500 2995 3504
rect 3119 3500 3123 3504
rect 3247 3500 3251 3504
rect 3375 3500 3379 3504
rect 111 3489 115 3493
rect 191 3492 195 3496
rect 327 3492 331 3496
rect 471 3492 475 3496
rect 623 3492 627 3496
rect 775 3492 779 3496
rect 919 3492 923 3496
rect 1055 3492 1059 3496
rect 1183 3492 1187 3496
rect 1311 3492 1315 3496
rect 1439 3492 1443 3496
rect 3591 3497 3595 3501
rect 1567 3492 1571 3496
rect 1831 3489 1835 3493
rect 1871 3480 1875 3484
rect 3591 3480 3595 3484
rect 111 3472 115 3476
rect 1831 3472 1835 3476
rect 2095 3462 2099 3466
rect 2175 3462 2179 3466
rect 2271 3462 2275 3466
rect 2375 3462 2379 3466
rect 2495 3462 2499 3466
rect 2623 3462 2627 3466
rect 2751 3462 2755 3466
rect 2879 3462 2883 3466
rect 2999 3462 3003 3466
rect 3127 3462 3131 3466
rect 3255 3462 3259 3466
rect 3383 3462 3387 3466
rect 199 3454 203 3458
rect 335 3454 339 3458
rect 479 3454 483 3458
rect 631 3454 635 3458
rect 783 3454 787 3458
rect 927 3454 931 3458
rect 1063 3454 1067 3458
rect 1191 3454 1195 3458
rect 1319 3454 1323 3458
rect 1447 3454 1451 3458
rect 1575 3454 1579 3458
rect 151 3422 155 3426
rect 295 3422 299 3426
rect 455 3422 459 3426
rect 623 3422 627 3426
rect 791 3422 795 3426
rect 959 3422 963 3426
rect 1119 3422 1123 3426
rect 1271 3422 1275 3426
rect 1415 3422 1419 3426
rect 1559 3422 1563 3426
rect 1711 3422 1715 3426
rect 2111 3422 2115 3426
rect 2199 3422 2203 3426
rect 2303 3422 2307 3426
rect 2415 3422 2419 3426
rect 2543 3422 2547 3426
rect 2679 3422 2683 3426
rect 2815 3422 2819 3426
rect 2959 3422 2963 3426
rect 3111 3422 3115 3426
rect 3263 3422 3267 3426
rect 3423 3422 3427 3426
rect 111 3404 115 3408
rect 1831 3404 1835 3408
rect 1871 3404 1875 3408
rect 3591 3404 3595 3408
rect 111 3387 115 3391
rect 143 3384 147 3388
rect 287 3384 291 3388
rect 447 3384 451 3388
rect 615 3384 619 3388
rect 783 3384 787 3388
rect 951 3384 955 3388
rect 1111 3384 1115 3388
rect 1263 3384 1267 3388
rect 1407 3384 1411 3388
rect 1551 3384 1555 3388
rect 1703 3384 1707 3388
rect 1831 3387 1835 3391
rect 1871 3387 1875 3391
rect 2103 3384 2107 3388
rect 2191 3384 2195 3388
rect 2295 3384 2299 3388
rect 2407 3384 2411 3388
rect 2535 3384 2539 3388
rect 2671 3384 2675 3388
rect 2807 3384 2811 3388
rect 2951 3384 2955 3388
rect 3103 3384 3107 3388
rect 3255 3384 3259 3388
rect 3415 3384 3419 3388
rect 3591 3387 3595 3391
rect 111 3337 115 3341
rect 207 3340 211 3344
rect 335 3340 339 3344
rect 471 3340 475 3344
rect 623 3340 627 3344
rect 783 3340 787 3344
rect 943 3340 947 3344
rect 1103 3340 1107 3344
rect 1263 3340 1267 3344
rect 1423 3340 1427 3344
rect 1583 3340 1587 3344
rect 1743 3340 1747 3344
rect 1831 3337 1835 3341
rect 1871 3333 1875 3337
rect 2127 3336 2131 3340
rect 2223 3336 2227 3340
rect 2335 3336 2339 3340
rect 2455 3336 2459 3340
rect 2583 3336 2587 3340
rect 2719 3336 2723 3340
rect 2863 3336 2867 3340
rect 3007 3336 3011 3340
rect 3159 3336 3163 3340
rect 3311 3336 3315 3340
rect 3471 3336 3475 3340
rect 3591 3333 3595 3337
rect 111 3320 115 3324
rect 1831 3320 1835 3324
rect 1871 3316 1875 3320
rect 3591 3316 3595 3320
rect 215 3302 219 3306
rect 343 3302 347 3306
rect 479 3302 483 3306
rect 631 3302 635 3306
rect 791 3302 795 3306
rect 951 3302 955 3306
rect 1111 3302 1115 3306
rect 1271 3302 1275 3306
rect 1431 3302 1435 3306
rect 1591 3302 1595 3306
rect 1751 3302 1755 3306
rect 2135 3298 2139 3302
rect 2231 3298 2235 3302
rect 2343 3298 2347 3302
rect 2463 3298 2467 3302
rect 2591 3298 2595 3302
rect 2727 3298 2731 3302
rect 2871 3298 2875 3302
rect 3015 3298 3019 3302
rect 3167 3298 3171 3302
rect 3319 3298 3323 3302
rect 3479 3298 3483 3302
rect 351 3266 355 3270
rect 455 3266 459 3270
rect 575 3266 579 3270
rect 703 3266 707 3270
rect 839 3266 843 3270
rect 983 3266 987 3270
rect 1119 3266 1123 3270
rect 1255 3266 1259 3270
rect 1383 3266 1387 3270
rect 1511 3266 1515 3270
rect 1639 3266 1643 3270
rect 1751 3266 1755 3270
rect 2135 3254 2139 3258
rect 2279 3254 2283 3258
rect 2415 3254 2419 3258
rect 2551 3254 2555 3258
rect 2687 3254 2691 3258
rect 2823 3254 2827 3258
rect 2959 3254 2963 3258
rect 3095 3254 3099 3258
rect 3231 3254 3235 3258
rect 3375 3254 3379 3258
rect 3511 3254 3515 3258
rect 111 3248 115 3252
rect 1831 3248 1835 3252
rect 1871 3236 1875 3240
rect 111 3231 115 3235
rect 3591 3236 3595 3240
rect 343 3228 347 3232
rect 447 3228 451 3232
rect 567 3228 571 3232
rect 695 3228 699 3232
rect 831 3228 835 3232
rect 975 3228 979 3232
rect 1111 3228 1115 3232
rect 1247 3228 1251 3232
rect 1375 3228 1379 3232
rect 1503 3228 1507 3232
rect 1631 3228 1635 3232
rect 1743 3228 1747 3232
rect 1831 3231 1835 3235
rect 1871 3219 1875 3223
rect 2127 3216 2131 3220
rect 2271 3216 2275 3220
rect 2407 3216 2411 3220
rect 2543 3216 2547 3220
rect 2679 3216 2683 3220
rect 2815 3216 2819 3220
rect 2951 3216 2955 3220
rect 3087 3216 3091 3220
rect 3223 3216 3227 3220
rect 3367 3216 3371 3220
rect 3503 3216 3507 3220
rect 3591 3219 3595 3223
rect 111 3181 115 3185
rect 487 3184 491 3188
rect 575 3184 579 3188
rect 663 3184 667 3188
rect 767 3184 771 3188
rect 887 3184 891 3188
rect 1023 3184 1027 3188
rect 1191 3184 1195 3188
rect 1375 3184 1379 3188
rect 1567 3184 1571 3188
rect 1743 3184 1747 3188
rect 1831 3181 1835 3185
rect 111 3164 115 3168
rect 1831 3164 1835 3168
rect 1871 3165 1875 3169
rect 1895 3168 1899 3172
rect 1991 3168 1995 3172
rect 2119 3168 2123 3172
rect 2247 3168 2251 3172
rect 2383 3168 2387 3172
rect 2511 3168 2515 3172
rect 2639 3168 2643 3172
rect 2767 3168 2771 3172
rect 2895 3168 2899 3172
rect 3031 3168 3035 3172
rect 3175 3168 3179 3172
rect 3327 3168 3331 3172
rect 3487 3168 3491 3172
rect 3591 3165 3595 3169
rect 495 3146 499 3150
rect 583 3146 587 3150
rect 671 3146 675 3150
rect 775 3146 779 3150
rect 895 3146 899 3150
rect 1031 3146 1035 3150
rect 1199 3146 1203 3150
rect 1383 3146 1387 3150
rect 1575 3146 1579 3150
rect 1751 3146 1755 3150
rect 1871 3148 1875 3152
rect 3591 3148 3595 3152
rect 1903 3130 1907 3134
rect 1999 3130 2003 3134
rect 2127 3130 2131 3134
rect 2255 3130 2259 3134
rect 2391 3130 2395 3134
rect 2519 3130 2523 3134
rect 2647 3130 2651 3134
rect 2775 3130 2779 3134
rect 2903 3130 2907 3134
rect 3039 3130 3043 3134
rect 3183 3130 3187 3134
rect 3335 3130 3339 3134
rect 3495 3130 3499 3134
rect 591 3110 595 3114
rect 671 3110 675 3114
rect 759 3110 763 3114
rect 847 3110 851 3114
rect 935 3110 939 3114
rect 1023 3110 1027 3114
rect 1111 3110 1115 3114
rect 1199 3110 1203 3114
rect 1287 3110 1291 3114
rect 1375 3110 1379 3114
rect 111 3092 115 3096
rect 1831 3092 1835 3096
rect 1903 3082 1907 3086
rect 2015 3082 2019 3086
rect 2191 3082 2195 3086
rect 2407 3082 2411 3086
rect 2655 3082 2659 3086
rect 2935 3082 2939 3086
rect 3231 3082 3235 3086
rect 3511 3082 3515 3086
rect 111 3075 115 3079
rect 583 3072 587 3076
rect 663 3072 667 3076
rect 751 3072 755 3076
rect 839 3072 843 3076
rect 927 3072 931 3076
rect 1015 3072 1019 3076
rect 1103 3072 1107 3076
rect 1191 3072 1195 3076
rect 1279 3072 1283 3076
rect 1367 3072 1371 3076
rect 1831 3075 1835 3079
rect 1871 3064 1875 3068
rect 3591 3064 3595 3068
rect 1871 3047 1875 3051
rect 1895 3044 1899 3048
rect 2007 3044 2011 3048
rect 2183 3044 2187 3048
rect 2399 3044 2403 3048
rect 2647 3044 2651 3048
rect 2927 3044 2931 3048
rect 3223 3044 3227 3048
rect 3503 3044 3507 3048
rect 3591 3047 3595 3051
rect 111 3021 115 3025
rect 543 3024 547 3028
rect 623 3024 627 3028
rect 711 3024 715 3028
rect 807 3024 811 3028
rect 903 3024 907 3028
rect 999 3024 1003 3028
rect 1087 3024 1091 3028
rect 1183 3024 1187 3028
rect 1279 3024 1283 3028
rect 1375 3024 1379 3028
rect 1471 3024 1475 3028
rect 1831 3021 1835 3025
rect 111 3004 115 3008
rect 1831 3004 1835 3008
rect 551 2986 555 2990
rect 631 2986 635 2990
rect 719 2986 723 2990
rect 815 2986 819 2990
rect 911 2986 915 2990
rect 1007 2986 1011 2990
rect 1095 2986 1099 2990
rect 1191 2986 1195 2990
rect 1287 2986 1291 2990
rect 1383 2986 1387 2990
rect 1479 2986 1483 2990
rect 1871 2989 1875 2993
rect 1895 2992 1899 2996
rect 2047 2992 2051 2996
rect 2223 2992 2227 2996
rect 2391 2992 2395 2996
rect 2543 2992 2547 2996
rect 2687 2992 2691 2996
rect 2815 2992 2819 2996
rect 2927 2992 2931 2996
rect 3039 2992 3043 2996
rect 3143 2992 3147 2996
rect 3239 2992 3243 2996
rect 3335 2992 3339 2996
rect 3423 2992 3427 2996
rect 3503 2992 3507 2996
rect 3591 2989 3595 2993
rect 1871 2972 1875 2976
rect 3591 2972 3595 2976
rect 471 2954 475 2958
rect 575 2954 579 2958
rect 687 2954 691 2958
rect 807 2954 811 2958
rect 943 2954 947 2958
rect 1087 2954 1091 2958
rect 1247 2954 1251 2958
rect 1415 2954 1419 2958
rect 1591 2954 1595 2958
rect 1751 2954 1755 2958
rect 1903 2954 1907 2958
rect 2055 2954 2059 2958
rect 2231 2954 2235 2958
rect 2399 2954 2403 2958
rect 2551 2954 2555 2958
rect 2695 2954 2699 2958
rect 2823 2954 2827 2958
rect 2935 2954 2939 2958
rect 3047 2954 3051 2958
rect 3151 2954 3155 2958
rect 3247 2954 3251 2958
rect 3343 2954 3347 2958
rect 3431 2954 3435 2958
rect 3511 2954 3515 2958
rect 111 2936 115 2940
rect 1831 2936 1835 2940
rect 111 2919 115 2923
rect 463 2916 467 2920
rect 567 2916 571 2920
rect 679 2916 683 2920
rect 799 2916 803 2920
rect 935 2916 939 2920
rect 1079 2916 1083 2920
rect 1239 2916 1243 2920
rect 1407 2916 1411 2920
rect 1583 2916 1587 2920
rect 1743 2916 1747 2920
rect 1831 2919 1835 2923
rect 1903 2922 1907 2926
rect 2087 2922 2091 2926
rect 2295 2922 2299 2926
rect 2487 2922 2491 2926
rect 2671 2922 2675 2926
rect 2839 2922 2843 2926
rect 2999 2922 3003 2926
rect 3151 2922 3155 2926
rect 3303 2922 3307 2926
rect 3455 2922 3459 2926
rect 1871 2904 1875 2908
rect 3591 2904 3595 2908
rect 1871 2887 1875 2891
rect 1895 2884 1899 2888
rect 2079 2884 2083 2888
rect 2287 2884 2291 2888
rect 2479 2884 2483 2888
rect 2663 2884 2667 2888
rect 2831 2884 2835 2888
rect 2991 2884 2995 2888
rect 3143 2884 3147 2888
rect 3295 2884 3299 2888
rect 3447 2884 3451 2888
rect 3591 2887 3595 2891
rect 111 2869 115 2873
rect 311 2872 315 2876
rect 431 2872 435 2876
rect 551 2872 555 2876
rect 679 2872 683 2876
rect 815 2872 819 2876
rect 951 2872 955 2876
rect 1087 2872 1091 2876
rect 1223 2872 1227 2876
rect 1359 2872 1363 2876
rect 1495 2872 1499 2876
rect 1631 2872 1635 2876
rect 1743 2872 1747 2876
rect 1831 2869 1835 2873
rect 111 2852 115 2856
rect 1831 2852 1835 2856
rect 319 2834 323 2838
rect 439 2834 443 2838
rect 559 2834 563 2838
rect 687 2834 691 2838
rect 823 2834 827 2838
rect 959 2834 963 2838
rect 1095 2834 1099 2838
rect 1231 2834 1235 2838
rect 1367 2834 1371 2838
rect 1503 2834 1507 2838
rect 1639 2834 1643 2838
rect 1751 2834 1755 2838
rect 1871 2829 1875 2833
rect 2135 2832 2139 2836
rect 2263 2832 2267 2836
rect 2391 2832 2395 2836
rect 2519 2832 2523 2836
rect 2647 2832 2651 2836
rect 2767 2832 2771 2836
rect 2887 2832 2891 2836
rect 3007 2832 3011 2836
rect 3135 2832 3139 2836
rect 3591 2829 3595 2833
rect 1871 2812 1875 2816
rect 3591 2812 3595 2816
rect 167 2802 171 2806
rect 303 2802 307 2806
rect 447 2802 451 2806
rect 607 2802 611 2806
rect 783 2802 787 2806
rect 959 2802 963 2806
rect 1143 2802 1147 2806
rect 1335 2802 1339 2806
rect 1535 2802 1539 2806
rect 1735 2802 1739 2806
rect 2143 2794 2147 2798
rect 2271 2794 2275 2798
rect 2399 2794 2403 2798
rect 2527 2794 2531 2798
rect 2655 2794 2659 2798
rect 2775 2794 2779 2798
rect 2895 2794 2899 2798
rect 3015 2794 3019 2798
rect 3143 2794 3147 2798
rect 111 2784 115 2788
rect 1831 2784 1835 2788
rect 111 2767 115 2771
rect 159 2764 163 2768
rect 295 2764 299 2768
rect 439 2764 443 2768
rect 599 2764 603 2768
rect 775 2764 779 2768
rect 951 2764 955 2768
rect 1135 2764 1139 2768
rect 1327 2764 1331 2768
rect 1527 2764 1531 2768
rect 1727 2764 1731 2768
rect 1831 2767 1835 2771
rect 2231 2754 2235 2758
rect 2311 2754 2315 2758
rect 2391 2754 2395 2758
rect 2471 2754 2475 2758
rect 2551 2754 2555 2758
rect 2639 2754 2643 2758
rect 2727 2754 2731 2758
rect 2815 2754 2819 2758
rect 2903 2754 2907 2758
rect 2991 2754 2995 2758
rect 1871 2736 1875 2740
rect 3591 2736 3595 2740
rect 111 2713 115 2717
rect 135 2716 139 2720
rect 247 2716 251 2720
rect 391 2716 395 2720
rect 551 2716 555 2720
rect 711 2716 715 2720
rect 879 2716 883 2720
rect 1039 2716 1043 2720
rect 1199 2716 1203 2720
rect 1359 2716 1363 2720
rect 1519 2716 1523 2720
rect 1687 2716 1691 2720
rect 1871 2719 1875 2723
rect 1831 2713 1835 2717
rect 2223 2716 2227 2720
rect 2303 2716 2307 2720
rect 2383 2716 2387 2720
rect 2463 2716 2467 2720
rect 2543 2716 2547 2720
rect 2631 2716 2635 2720
rect 2719 2716 2723 2720
rect 2807 2716 2811 2720
rect 2895 2716 2899 2720
rect 2983 2716 2987 2720
rect 3591 2719 3595 2723
rect 111 2696 115 2700
rect 1831 2696 1835 2700
rect 143 2678 147 2682
rect 255 2678 259 2682
rect 399 2678 403 2682
rect 559 2678 563 2682
rect 719 2678 723 2682
rect 887 2678 891 2682
rect 1047 2678 1051 2682
rect 1207 2678 1211 2682
rect 1367 2678 1371 2682
rect 1527 2678 1531 2682
rect 1695 2678 1699 2682
rect 1871 2669 1875 2673
rect 2239 2672 2243 2676
rect 2319 2672 2323 2676
rect 2399 2672 2403 2676
rect 2479 2672 2483 2676
rect 2559 2672 2563 2676
rect 2639 2672 2643 2676
rect 2719 2672 2723 2676
rect 2799 2672 2803 2676
rect 2879 2672 2883 2676
rect 2959 2672 2963 2676
rect 3591 2669 3595 2673
rect 1871 2652 1875 2656
rect 3591 2652 3595 2656
rect 143 2646 147 2650
rect 255 2646 259 2650
rect 399 2646 403 2650
rect 551 2646 555 2650
rect 711 2646 715 2650
rect 879 2646 883 2650
rect 1047 2646 1051 2650
rect 1215 2646 1219 2650
rect 1391 2646 1395 2650
rect 1567 2646 1571 2650
rect 2247 2634 2251 2638
rect 2327 2634 2331 2638
rect 2407 2634 2411 2638
rect 2487 2634 2491 2638
rect 2567 2634 2571 2638
rect 2647 2634 2651 2638
rect 2727 2634 2731 2638
rect 2807 2634 2811 2638
rect 2887 2634 2891 2638
rect 2967 2634 2971 2638
rect 111 2628 115 2632
rect 1831 2628 1835 2632
rect 111 2611 115 2615
rect 135 2608 139 2612
rect 247 2608 251 2612
rect 391 2608 395 2612
rect 543 2608 547 2612
rect 703 2608 707 2612
rect 871 2608 875 2612
rect 1039 2608 1043 2612
rect 1207 2608 1211 2612
rect 1383 2608 1387 2612
rect 1559 2608 1563 2612
rect 1831 2611 1835 2615
rect 2191 2594 2195 2598
rect 2271 2594 2275 2598
rect 2351 2594 2355 2598
rect 2431 2594 2435 2598
rect 2511 2594 2515 2598
rect 2591 2594 2595 2598
rect 2671 2594 2675 2598
rect 2751 2594 2755 2598
rect 2831 2594 2835 2598
rect 2911 2594 2915 2598
rect 2991 2594 2995 2598
rect 1871 2576 1875 2580
rect 3591 2576 3595 2580
rect 111 2557 115 2561
rect 159 2560 163 2564
rect 279 2560 283 2564
rect 415 2560 419 2564
rect 559 2560 563 2564
rect 703 2560 707 2564
rect 847 2560 851 2564
rect 983 2560 987 2564
rect 1119 2560 1123 2564
rect 1255 2560 1259 2564
rect 1391 2560 1395 2564
rect 1527 2560 1531 2564
rect 1831 2557 1835 2561
rect 1871 2559 1875 2563
rect 2183 2556 2187 2560
rect 2263 2556 2267 2560
rect 2343 2556 2347 2560
rect 2423 2556 2427 2560
rect 2503 2556 2507 2560
rect 2583 2556 2587 2560
rect 2663 2556 2667 2560
rect 2743 2556 2747 2560
rect 2823 2556 2827 2560
rect 2903 2556 2907 2560
rect 2983 2556 2987 2560
rect 3591 2559 3595 2563
rect 111 2540 115 2544
rect 1831 2540 1835 2544
rect 167 2522 171 2526
rect 287 2522 291 2526
rect 423 2522 427 2526
rect 567 2522 571 2526
rect 711 2522 715 2526
rect 855 2522 859 2526
rect 991 2522 995 2526
rect 1127 2522 1131 2526
rect 1263 2522 1267 2526
rect 1399 2522 1403 2526
rect 1535 2522 1539 2526
rect 1871 2501 1875 2505
rect 2119 2504 2123 2508
rect 2207 2504 2211 2508
rect 2303 2504 2307 2508
rect 2399 2504 2403 2508
rect 2495 2504 2499 2508
rect 2591 2504 2595 2508
rect 2687 2504 2691 2508
rect 2783 2504 2787 2508
rect 2879 2504 2883 2508
rect 2975 2504 2979 2508
rect 3079 2504 3083 2508
rect 3591 2501 3595 2505
rect 335 2486 339 2490
rect 415 2486 419 2490
rect 503 2486 507 2490
rect 599 2486 603 2490
rect 703 2486 707 2490
rect 815 2486 819 2490
rect 935 2486 939 2490
rect 1063 2486 1067 2490
rect 1191 2486 1195 2490
rect 1327 2486 1331 2490
rect 1471 2486 1475 2490
rect 1871 2484 1875 2488
rect 3591 2484 3595 2488
rect 111 2468 115 2472
rect 1831 2468 1835 2472
rect 2127 2466 2131 2470
rect 2215 2466 2219 2470
rect 2311 2466 2315 2470
rect 2407 2466 2411 2470
rect 2503 2466 2507 2470
rect 2599 2466 2603 2470
rect 2695 2466 2699 2470
rect 2791 2466 2795 2470
rect 2887 2466 2891 2470
rect 2983 2466 2987 2470
rect 3087 2466 3091 2470
rect 111 2451 115 2455
rect 327 2448 331 2452
rect 407 2448 411 2452
rect 495 2448 499 2452
rect 591 2448 595 2452
rect 695 2448 699 2452
rect 807 2448 811 2452
rect 927 2448 931 2452
rect 1055 2448 1059 2452
rect 1183 2448 1187 2452
rect 1319 2448 1323 2452
rect 1463 2448 1467 2452
rect 1831 2451 1835 2455
rect 1903 2430 1907 2434
rect 1991 2430 1995 2434
rect 2111 2430 2115 2434
rect 2247 2430 2251 2434
rect 2391 2430 2395 2434
rect 2535 2430 2539 2434
rect 2671 2430 2675 2434
rect 2807 2430 2811 2434
rect 2943 2430 2947 2434
rect 3079 2430 3083 2434
rect 3215 2430 3219 2434
rect 1871 2412 1875 2416
rect 3591 2412 3595 2416
rect 111 2393 115 2397
rect 383 2396 387 2400
rect 463 2396 467 2400
rect 543 2396 547 2400
rect 623 2396 627 2400
rect 703 2396 707 2400
rect 783 2396 787 2400
rect 863 2396 867 2400
rect 943 2396 947 2400
rect 1023 2396 1027 2400
rect 1103 2396 1107 2400
rect 1183 2396 1187 2400
rect 1263 2396 1267 2400
rect 1351 2396 1355 2400
rect 1439 2396 1443 2400
rect 1527 2396 1531 2400
rect 1831 2393 1835 2397
rect 1871 2395 1875 2399
rect 1895 2392 1899 2396
rect 1983 2392 1987 2396
rect 2103 2392 2107 2396
rect 2239 2392 2243 2396
rect 2383 2392 2387 2396
rect 2527 2392 2531 2396
rect 2663 2392 2667 2396
rect 2799 2392 2803 2396
rect 2935 2392 2939 2396
rect 3071 2392 3075 2396
rect 3207 2392 3211 2396
rect 3591 2395 3595 2399
rect 111 2376 115 2380
rect 1831 2376 1835 2380
rect 391 2358 395 2362
rect 471 2358 475 2362
rect 551 2358 555 2362
rect 631 2358 635 2362
rect 711 2358 715 2362
rect 791 2358 795 2362
rect 871 2358 875 2362
rect 951 2358 955 2362
rect 1031 2358 1035 2362
rect 1111 2358 1115 2362
rect 1191 2358 1195 2362
rect 1271 2358 1275 2362
rect 1359 2358 1363 2362
rect 1447 2358 1451 2362
rect 1535 2358 1539 2362
rect 1871 2337 1875 2341
rect 1895 2340 1899 2344
rect 2015 2340 2019 2344
rect 2175 2340 2179 2344
rect 2343 2340 2347 2344
rect 2511 2340 2515 2344
rect 2671 2340 2675 2344
rect 2823 2340 2827 2344
rect 2959 2340 2963 2344
rect 3079 2340 3083 2344
rect 3191 2340 3195 2344
rect 3303 2340 3307 2344
rect 3415 2340 3419 2344
rect 3503 2340 3507 2344
rect 3591 2337 3595 2341
rect 1407 2326 1411 2330
rect 1487 2326 1491 2330
rect 1567 2326 1571 2330
rect 1647 2326 1651 2330
rect 1871 2320 1875 2324
rect 3591 2320 3595 2324
rect 111 2308 115 2312
rect 1831 2308 1835 2312
rect 1903 2302 1907 2306
rect 2023 2302 2027 2306
rect 2183 2302 2187 2306
rect 2351 2302 2355 2306
rect 2519 2302 2523 2306
rect 2679 2302 2683 2306
rect 2831 2302 2835 2306
rect 2967 2302 2971 2306
rect 3087 2302 3091 2306
rect 3199 2302 3203 2306
rect 3311 2302 3315 2306
rect 3423 2302 3427 2306
rect 3511 2302 3515 2306
rect 111 2291 115 2295
rect 1399 2288 1403 2292
rect 1479 2288 1483 2292
rect 1559 2288 1563 2292
rect 1639 2288 1643 2292
rect 1831 2291 1835 2295
rect 1903 2270 1907 2274
rect 2031 2270 2035 2274
rect 2183 2270 2187 2274
rect 2367 2270 2371 2274
rect 2575 2270 2579 2274
rect 2791 2270 2795 2274
rect 3023 2270 3027 2274
rect 3255 2270 3259 2274
rect 3495 2270 3499 2274
rect 1871 2252 1875 2256
rect 3591 2252 3595 2256
rect 111 2233 115 2237
rect 135 2236 139 2240
rect 215 2236 219 2240
rect 295 2236 299 2240
rect 383 2236 387 2240
rect 519 2236 523 2240
rect 671 2236 675 2240
rect 831 2236 835 2240
rect 999 2236 1003 2240
rect 1159 2236 1163 2240
rect 1311 2236 1315 2240
rect 1455 2236 1459 2240
rect 1607 2236 1611 2240
rect 1743 2236 1747 2240
rect 1831 2233 1835 2237
rect 1871 2235 1875 2239
rect 1895 2232 1899 2236
rect 2023 2232 2027 2236
rect 2175 2232 2179 2236
rect 2359 2232 2363 2236
rect 2567 2232 2571 2236
rect 2783 2232 2787 2236
rect 3015 2232 3019 2236
rect 3247 2232 3251 2236
rect 3487 2232 3491 2236
rect 3591 2235 3595 2239
rect 111 2216 115 2220
rect 1831 2216 1835 2220
rect 143 2198 147 2202
rect 223 2198 227 2202
rect 303 2198 307 2202
rect 391 2198 395 2202
rect 527 2198 531 2202
rect 679 2198 683 2202
rect 839 2198 843 2202
rect 1007 2198 1011 2202
rect 1167 2198 1171 2202
rect 1319 2198 1323 2202
rect 1463 2198 1467 2202
rect 1615 2198 1619 2202
rect 1751 2198 1755 2202
rect 191 2162 195 2166
rect 311 2162 315 2166
rect 463 2162 467 2166
rect 639 2162 643 2166
rect 823 2162 827 2166
rect 1015 2162 1019 2166
rect 1199 2162 1203 2166
rect 1391 2162 1395 2166
rect 1583 2162 1587 2166
rect 1751 2162 1755 2166
rect 1871 2165 1875 2169
rect 2199 2168 2203 2172
rect 2295 2168 2299 2172
rect 2399 2168 2403 2172
rect 2519 2168 2523 2172
rect 2639 2168 2643 2172
rect 2759 2168 2763 2172
rect 2879 2168 2883 2172
rect 2991 2168 2995 2172
rect 3095 2168 3099 2172
rect 3199 2168 3203 2172
rect 3303 2168 3307 2172
rect 3407 2168 3411 2172
rect 3503 2168 3507 2172
rect 3591 2165 3595 2169
rect 111 2144 115 2148
rect 1831 2144 1835 2148
rect 1871 2148 1875 2152
rect 3591 2148 3595 2152
rect 111 2127 115 2131
rect 183 2124 187 2128
rect 303 2124 307 2128
rect 455 2124 459 2128
rect 631 2124 635 2128
rect 815 2124 819 2128
rect 1007 2124 1011 2128
rect 1191 2124 1195 2128
rect 1383 2124 1387 2128
rect 1575 2124 1579 2128
rect 1743 2124 1747 2128
rect 1831 2127 1835 2131
rect 2207 2130 2211 2134
rect 2303 2130 2307 2134
rect 2407 2130 2411 2134
rect 2527 2130 2531 2134
rect 2647 2130 2651 2134
rect 2767 2130 2771 2134
rect 2887 2130 2891 2134
rect 2999 2130 3003 2134
rect 3103 2130 3107 2134
rect 3207 2130 3211 2134
rect 3311 2130 3315 2134
rect 3415 2130 3419 2134
rect 3511 2130 3515 2134
rect 2175 2086 2179 2090
rect 2271 2086 2275 2090
rect 2375 2086 2379 2090
rect 2487 2086 2491 2090
rect 2607 2086 2611 2090
rect 2727 2086 2731 2090
rect 2847 2086 2851 2090
rect 2967 2086 2971 2090
rect 3079 2086 3083 2090
rect 3191 2086 3195 2090
rect 3303 2086 3307 2090
rect 3415 2086 3419 2090
rect 3511 2086 3515 2090
rect 111 2073 115 2077
rect 215 2076 219 2080
rect 359 2076 363 2080
rect 519 2076 523 2080
rect 703 2076 707 2080
rect 895 2076 899 2080
rect 1103 2076 1107 2080
rect 1311 2076 1315 2080
rect 1527 2076 1531 2080
rect 1743 2076 1747 2080
rect 1831 2073 1835 2077
rect 1871 2068 1875 2072
rect 3591 2068 3595 2072
rect 111 2056 115 2060
rect 1831 2056 1835 2060
rect 1871 2051 1875 2055
rect 2167 2048 2171 2052
rect 2263 2048 2267 2052
rect 2367 2048 2371 2052
rect 2479 2048 2483 2052
rect 2599 2048 2603 2052
rect 2719 2048 2723 2052
rect 2839 2048 2843 2052
rect 2959 2048 2963 2052
rect 3071 2048 3075 2052
rect 3183 2048 3187 2052
rect 3295 2048 3299 2052
rect 3407 2048 3411 2052
rect 3503 2048 3507 2052
rect 3591 2051 3595 2055
rect 223 2038 227 2042
rect 367 2038 371 2042
rect 527 2038 531 2042
rect 711 2038 715 2042
rect 903 2038 907 2042
rect 1111 2038 1115 2042
rect 1319 2038 1323 2042
rect 1535 2038 1539 2042
rect 1751 2038 1755 2042
rect 143 2006 147 2010
rect 263 2006 267 2010
rect 383 2006 387 2010
rect 495 2006 499 2010
rect 607 2006 611 2010
rect 719 2006 723 2010
rect 823 2006 827 2010
rect 927 2006 931 2010
rect 1023 2006 1027 2010
rect 1111 2006 1115 2010
rect 1207 2006 1211 2010
rect 1295 2006 1299 2010
rect 1391 2006 1395 2010
rect 1487 2006 1491 2010
rect 1583 2006 1587 2010
rect 1671 2006 1675 2010
rect 1751 2006 1755 2010
rect 1871 1997 1875 2001
rect 2071 2000 2075 2004
rect 2207 2000 2211 2004
rect 2359 2000 2363 2004
rect 2519 2000 2523 2004
rect 2679 2000 2683 2004
rect 2847 2000 2851 2004
rect 3015 2000 3019 2004
rect 3183 2000 3187 2004
rect 3351 2000 3355 2004
rect 3503 2000 3507 2004
rect 3591 1997 3595 2001
rect 111 1988 115 1992
rect 1831 1988 1835 1992
rect 1871 1980 1875 1984
rect 3591 1980 3595 1984
rect 111 1971 115 1975
rect 135 1968 139 1972
rect 255 1968 259 1972
rect 375 1968 379 1972
rect 487 1968 491 1972
rect 599 1968 603 1972
rect 711 1968 715 1972
rect 815 1968 819 1972
rect 919 1968 923 1972
rect 1015 1968 1019 1972
rect 1103 1968 1107 1972
rect 1199 1968 1203 1972
rect 1287 1968 1291 1972
rect 1383 1968 1387 1972
rect 1479 1968 1483 1972
rect 1575 1968 1579 1972
rect 1663 1968 1667 1972
rect 1743 1968 1747 1972
rect 1831 1971 1835 1975
rect 2079 1962 2083 1966
rect 2215 1962 2219 1966
rect 2367 1962 2371 1966
rect 2527 1962 2531 1966
rect 2687 1962 2691 1966
rect 2855 1962 2859 1966
rect 3023 1962 3027 1966
rect 3191 1962 3195 1966
rect 3359 1962 3363 1966
rect 3511 1962 3515 1966
rect 1903 1930 1907 1934
rect 2007 1930 2011 1934
rect 2135 1930 2139 1934
rect 2255 1930 2259 1934
rect 2375 1930 2379 1934
rect 2487 1930 2491 1934
rect 2599 1930 2603 1934
rect 2719 1930 2723 1934
rect 2839 1930 2843 1934
rect 111 1913 115 1917
rect 167 1916 171 1920
rect 327 1916 331 1920
rect 487 1916 491 1920
rect 647 1916 651 1920
rect 799 1916 803 1920
rect 943 1916 947 1920
rect 1079 1916 1083 1920
rect 1215 1916 1219 1920
rect 1351 1916 1355 1920
rect 1487 1916 1491 1920
rect 1623 1916 1627 1920
rect 1743 1916 1747 1920
rect 1831 1913 1835 1917
rect 1871 1912 1875 1916
rect 3591 1912 3595 1916
rect 111 1896 115 1900
rect 1831 1896 1835 1900
rect 1871 1895 1875 1899
rect 1895 1892 1899 1896
rect 1999 1892 2003 1896
rect 2127 1892 2131 1896
rect 2247 1892 2251 1896
rect 2367 1892 2371 1896
rect 2479 1892 2483 1896
rect 2591 1892 2595 1896
rect 2711 1892 2715 1896
rect 2831 1892 2835 1896
rect 3591 1895 3595 1899
rect 175 1878 179 1882
rect 335 1878 339 1882
rect 495 1878 499 1882
rect 655 1878 659 1882
rect 807 1878 811 1882
rect 951 1878 955 1882
rect 1087 1878 1091 1882
rect 1223 1878 1227 1882
rect 1359 1878 1363 1882
rect 1495 1878 1499 1882
rect 1631 1878 1635 1882
rect 1751 1878 1755 1882
rect 159 1846 163 1850
rect 303 1846 307 1850
rect 447 1846 451 1850
rect 599 1846 603 1850
rect 751 1846 755 1850
rect 903 1846 907 1850
rect 1055 1846 1059 1850
rect 1207 1846 1211 1850
rect 1351 1846 1355 1850
rect 1487 1846 1491 1850
rect 1631 1846 1635 1850
rect 1751 1846 1755 1850
rect 1871 1845 1875 1849
rect 1895 1848 1899 1852
rect 1991 1848 1995 1852
rect 2119 1848 2123 1852
rect 2247 1848 2251 1852
rect 2383 1848 2387 1852
rect 2519 1848 2523 1852
rect 2655 1848 2659 1852
rect 2807 1848 2811 1852
rect 2975 1848 2979 1852
rect 3151 1848 3155 1852
rect 3335 1848 3339 1852
rect 3503 1848 3507 1852
rect 3591 1845 3595 1849
rect 111 1828 115 1832
rect 1831 1828 1835 1832
rect 1871 1828 1875 1832
rect 3591 1828 3595 1832
rect 111 1811 115 1815
rect 151 1808 155 1812
rect 295 1808 299 1812
rect 439 1808 443 1812
rect 591 1808 595 1812
rect 743 1808 747 1812
rect 895 1808 899 1812
rect 1047 1808 1051 1812
rect 1199 1808 1203 1812
rect 1343 1808 1347 1812
rect 1479 1808 1483 1812
rect 1623 1808 1627 1812
rect 1743 1808 1747 1812
rect 1831 1811 1835 1815
rect 1903 1810 1907 1814
rect 1999 1810 2003 1814
rect 2127 1810 2131 1814
rect 2255 1810 2259 1814
rect 2391 1810 2395 1814
rect 2527 1810 2531 1814
rect 2663 1810 2667 1814
rect 2815 1810 2819 1814
rect 2983 1810 2987 1814
rect 3159 1810 3163 1814
rect 3343 1810 3347 1814
rect 3511 1810 3515 1814
rect 1903 1766 1907 1770
rect 2031 1766 2035 1770
rect 2191 1766 2195 1770
rect 2359 1766 2363 1770
rect 2527 1766 2531 1770
rect 2687 1766 2691 1770
rect 2839 1766 2843 1770
rect 2983 1766 2987 1770
rect 3119 1766 3123 1770
rect 3255 1766 3259 1770
rect 3391 1766 3395 1770
rect 3511 1766 3515 1770
rect 111 1757 115 1761
rect 247 1760 251 1764
rect 423 1760 427 1764
rect 591 1760 595 1764
rect 751 1760 755 1764
rect 895 1760 899 1764
rect 1023 1760 1027 1764
rect 1143 1760 1147 1764
rect 1263 1760 1267 1764
rect 1391 1760 1395 1764
rect 1831 1757 1835 1761
rect 1871 1748 1875 1752
rect 3591 1748 3595 1752
rect 111 1740 115 1744
rect 1831 1740 1835 1744
rect 1871 1731 1875 1735
rect 1895 1728 1899 1732
rect 2023 1728 2027 1732
rect 2183 1728 2187 1732
rect 2351 1728 2355 1732
rect 2519 1728 2523 1732
rect 2679 1728 2683 1732
rect 2831 1728 2835 1732
rect 2975 1728 2979 1732
rect 3111 1728 3115 1732
rect 3247 1728 3251 1732
rect 3383 1728 3387 1732
rect 3503 1728 3507 1732
rect 3591 1731 3595 1735
rect 255 1722 259 1726
rect 431 1722 435 1726
rect 599 1722 603 1726
rect 759 1722 763 1726
rect 903 1722 907 1726
rect 1031 1722 1035 1726
rect 1151 1722 1155 1726
rect 1271 1722 1275 1726
rect 1399 1722 1403 1726
rect 191 1686 195 1690
rect 311 1686 315 1690
rect 447 1686 451 1690
rect 591 1686 595 1690
rect 743 1686 747 1690
rect 895 1686 899 1690
rect 1039 1686 1043 1690
rect 1183 1686 1187 1690
rect 1319 1686 1323 1690
rect 1447 1686 1451 1690
rect 1575 1686 1579 1690
rect 1711 1686 1715 1690
rect 1871 1677 1875 1681
rect 1895 1680 1899 1684
rect 1991 1680 1995 1684
rect 2135 1680 2139 1684
rect 2295 1680 2299 1684
rect 2471 1680 2475 1684
rect 2647 1680 2651 1684
rect 2815 1680 2819 1684
rect 2967 1680 2971 1684
rect 3111 1680 3115 1684
rect 3247 1680 3251 1684
rect 3383 1680 3387 1684
rect 3503 1680 3507 1684
rect 3591 1677 3595 1681
rect 111 1668 115 1672
rect 1831 1668 1835 1672
rect 1871 1660 1875 1664
rect 3591 1660 3595 1664
rect 111 1651 115 1655
rect 183 1648 187 1652
rect 303 1648 307 1652
rect 439 1648 443 1652
rect 583 1648 587 1652
rect 735 1648 739 1652
rect 887 1648 891 1652
rect 1031 1648 1035 1652
rect 1175 1648 1179 1652
rect 1311 1648 1315 1652
rect 1439 1648 1443 1652
rect 1567 1648 1571 1652
rect 1703 1648 1707 1652
rect 1831 1651 1835 1655
rect 1903 1642 1907 1646
rect 1999 1642 2003 1646
rect 2143 1642 2147 1646
rect 2303 1642 2307 1646
rect 2479 1642 2483 1646
rect 2655 1642 2659 1646
rect 2823 1642 2827 1646
rect 2975 1642 2979 1646
rect 3119 1642 3123 1646
rect 3255 1642 3259 1646
rect 3391 1642 3395 1646
rect 3511 1642 3515 1646
rect 1975 1606 1979 1610
rect 2095 1606 2099 1610
rect 2231 1606 2235 1610
rect 2367 1606 2371 1610
rect 2503 1606 2507 1610
rect 2639 1606 2643 1610
rect 2775 1606 2779 1610
rect 2911 1606 2915 1610
rect 3055 1606 3059 1610
rect 3207 1606 3211 1610
rect 3367 1606 3371 1610
rect 3511 1606 3515 1610
rect 111 1593 115 1597
rect 167 1596 171 1600
rect 351 1596 355 1600
rect 543 1596 547 1600
rect 727 1596 731 1600
rect 903 1596 907 1600
rect 1071 1596 1075 1600
rect 1223 1596 1227 1600
rect 1359 1596 1363 1600
rect 1495 1596 1499 1600
rect 1623 1596 1627 1600
rect 1743 1596 1747 1600
rect 1831 1593 1835 1597
rect 1871 1588 1875 1592
rect 3591 1588 3595 1592
rect 111 1576 115 1580
rect 1831 1576 1835 1580
rect 1871 1571 1875 1575
rect 1967 1568 1971 1572
rect 2087 1568 2091 1572
rect 2223 1568 2227 1572
rect 2359 1568 2363 1572
rect 2495 1568 2499 1572
rect 2631 1568 2635 1572
rect 2767 1568 2771 1572
rect 2903 1568 2907 1572
rect 3047 1568 3051 1572
rect 3199 1568 3203 1572
rect 3359 1568 3363 1572
rect 3503 1568 3507 1572
rect 3591 1571 3595 1575
rect 175 1558 179 1562
rect 359 1558 363 1562
rect 551 1558 555 1562
rect 735 1558 739 1562
rect 911 1558 915 1562
rect 1079 1558 1083 1562
rect 1231 1558 1235 1562
rect 1367 1558 1371 1562
rect 1503 1558 1507 1562
rect 1631 1558 1635 1562
rect 1751 1558 1755 1562
rect 143 1522 147 1526
rect 247 1522 251 1526
rect 383 1522 387 1526
rect 527 1522 531 1526
rect 671 1522 675 1526
rect 815 1522 819 1526
rect 951 1522 955 1526
rect 1079 1522 1083 1526
rect 1207 1522 1211 1526
rect 1335 1522 1339 1526
rect 1471 1522 1475 1526
rect 1871 1517 1875 1521
rect 2087 1520 2091 1524
rect 2167 1520 2171 1524
rect 2255 1520 2259 1524
rect 2343 1520 2347 1524
rect 2439 1520 2443 1524
rect 2535 1520 2539 1524
rect 2647 1520 2651 1524
rect 2783 1520 2787 1524
rect 2943 1520 2947 1524
rect 3119 1520 3123 1524
rect 3303 1520 3307 1524
rect 3495 1520 3499 1524
rect 3591 1517 3595 1521
rect 111 1504 115 1508
rect 1831 1504 1835 1508
rect 1871 1500 1875 1504
rect 3591 1500 3595 1504
rect 111 1487 115 1491
rect 135 1484 139 1488
rect 239 1484 243 1488
rect 375 1484 379 1488
rect 519 1484 523 1488
rect 663 1484 667 1488
rect 807 1484 811 1488
rect 943 1484 947 1488
rect 1071 1484 1075 1488
rect 1199 1484 1203 1488
rect 1327 1484 1331 1488
rect 1463 1484 1467 1488
rect 1831 1487 1835 1491
rect 2095 1482 2099 1486
rect 2175 1482 2179 1486
rect 2263 1482 2267 1486
rect 2351 1482 2355 1486
rect 2447 1482 2451 1486
rect 2543 1482 2547 1486
rect 2655 1482 2659 1486
rect 2791 1482 2795 1486
rect 2951 1482 2955 1486
rect 3127 1482 3131 1486
rect 3311 1482 3315 1486
rect 3503 1482 3507 1486
rect 2263 1446 2267 1450
rect 2343 1446 2347 1450
rect 2423 1446 2427 1450
rect 2503 1446 2507 1450
rect 2607 1446 2611 1450
rect 2735 1446 2739 1450
rect 2895 1446 2899 1450
rect 3079 1446 3083 1450
rect 3279 1446 3283 1450
rect 3479 1446 3483 1450
rect 111 1433 115 1437
rect 135 1436 139 1440
rect 231 1436 235 1440
rect 359 1436 363 1440
rect 479 1436 483 1440
rect 599 1436 603 1440
rect 719 1436 723 1440
rect 831 1436 835 1440
rect 935 1436 939 1440
rect 1039 1436 1043 1440
rect 1143 1436 1147 1440
rect 1255 1436 1259 1440
rect 1831 1433 1835 1437
rect 1871 1428 1875 1432
rect 3591 1428 3595 1432
rect 111 1416 115 1420
rect 1831 1416 1835 1420
rect 1871 1411 1875 1415
rect 2255 1408 2259 1412
rect 2335 1408 2339 1412
rect 2415 1408 2419 1412
rect 2495 1408 2499 1412
rect 2599 1408 2603 1412
rect 2727 1408 2731 1412
rect 2887 1408 2891 1412
rect 3071 1408 3075 1412
rect 3271 1408 3275 1412
rect 3471 1408 3475 1412
rect 3591 1411 3595 1415
rect 143 1398 147 1402
rect 239 1398 243 1402
rect 367 1398 371 1402
rect 487 1398 491 1402
rect 607 1398 611 1402
rect 727 1398 731 1402
rect 839 1398 843 1402
rect 943 1398 947 1402
rect 1047 1398 1051 1402
rect 1151 1398 1155 1402
rect 1263 1398 1267 1402
rect 1871 1361 1875 1365
rect 2263 1364 2267 1368
rect 2343 1364 2347 1368
rect 2423 1364 2427 1368
rect 2503 1364 2507 1368
rect 2591 1364 2595 1368
rect 2695 1364 2699 1368
rect 2807 1364 2811 1368
rect 2919 1364 2923 1368
rect 3039 1364 3043 1368
rect 3159 1364 3163 1368
rect 3279 1364 3283 1368
rect 3399 1364 3403 1368
rect 3503 1364 3507 1368
rect 3591 1361 3595 1365
rect 143 1350 147 1354
rect 287 1350 291 1354
rect 431 1350 435 1354
rect 583 1350 587 1354
rect 735 1350 739 1354
rect 879 1350 883 1354
rect 1023 1350 1027 1354
rect 1167 1350 1171 1354
rect 1319 1350 1323 1354
rect 1471 1350 1475 1354
rect 1623 1350 1627 1354
rect 1871 1344 1875 1348
rect 3591 1344 3595 1348
rect 111 1332 115 1336
rect 1831 1332 1835 1336
rect 2271 1326 2275 1330
rect 2351 1326 2355 1330
rect 2431 1326 2435 1330
rect 2511 1326 2515 1330
rect 2599 1326 2603 1330
rect 2703 1326 2707 1330
rect 2815 1326 2819 1330
rect 2927 1326 2931 1330
rect 3047 1326 3051 1330
rect 3167 1326 3171 1330
rect 3287 1326 3291 1330
rect 3407 1326 3411 1330
rect 3511 1326 3515 1330
rect 111 1315 115 1319
rect 135 1312 139 1316
rect 279 1312 283 1316
rect 423 1312 427 1316
rect 575 1312 579 1316
rect 727 1312 731 1316
rect 871 1312 875 1316
rect 1015 1312 1019 1316
rect 1159 1312 1163 1316
rect 1311 1312 1315 1316
rect 1463 1312 1467 1316
rect 1615 1312 1619 1316
rect 1831 1315 1835 1319
rect 2215 1282 2219 1286
rect 2295 1282 2299 1286
rect 2375 1282 2379 1286
rect 2455 1282 2459 1286
rect 2551 1282 2555 1286
rect 2663 1282 2667 1286
rect 2791 1282 2795 1286
rect 2927 1282 2931 1286
rect 3071 1282 3075 1286
rect 3215 1282 3219 1286
rect 3367 1282 3371 1286
rect 3511 1282 3515 1286
rect 111 1261 115 1265
rect 135 1264 139 1268
rect 263 1264 267 1268
rect 423 1264 427 1268
rect 591 1264 595 1268
rect 759 1264 763 1268
rect 927 1264 931 1268
rect 1079 1264 1083 1268
rect 1223 1264 1227 1268
rect 1351 1264 1355 1268
rect 1479 1264 1483 1268
rect 1607 1264 1611 1268
rect 1735 1264 1739 1268
rect 1831 1261 1835 1265
rect 1871 1264 1875 1268
rect 3591 1264 3595 1268
rect 111 1244 115 1248
rect 1831 1244 1835 1248
rect 1871 1247 1875 1251
rect 2207 1244 2211 1248
rect 2287 1244 2291 1248
rect 2367 1244 2371 1248
rect 2447 1244 2451 1248
rect 2543 1244 2547 1248
rect 2655 1244 2659 1248
rect 2783 1244 2787 1248
rect 2919 1244 2923 1248
rect 3063 1244 3067 1248
rect 3207 1244 3211 1248
rect 3359 1244 3363 1248
rect 3503 1244 3507 1248
rect 3591 1247 3595 1251
rect 143 1226 147 1230
rect 271 1226 275 1230
rect 431 1226 435 1230
rect 599 1226 603 1230
rect 767 1226 771 1230
rect 935 1226 939 1230
rect 1087 1226 1091 1230
rect 1231 1226 1235 1230
rect 1359 1226 1363 1230
rect 1487 1226 1491 1230
rect 1615 1226 1619 1230
rect 1743 1226 1747 1230
rect 1871 1193 1875 1197
rect 2111 1196 2115 1200
rect 2207 1196 2211 1200
rect 2303 1196 2307 1200
rect 2407 1196 2411 1200
rect 2527 1196 2531 1200
rect 2647 1196 2651 1200
rect 2775 1196 2779 1200
rect 2911 1196 2915 1200
rect 3055 1196 3059 1200
rect 3199 1196 3203 1200
rect 3343 1196 3347 1200
rect 3495 1196 3499 1200
rect 3591 1193 3595 1197
rect 143 1186 147 1190
rect 311 1186 315 1190
rect 487 1186 491 1190
rect 671 1186 675 1190
rect 847 1186 851 1190
rect 1007 1186 1011 1190
rect 1159 1186 1163 1190
rect 1295 1186 1299 1190
rect 1415 1186 1419 1190
rect 1535 1186 1539 1190
rect 1655 1186 1659 1190
rect 1751 1186 1755 1190
rect 1871 1176 1875 1180
rect 3591 1176 3595 1180
rect 111 1168 115 1172
rect 1831 1168 1835 1172
rect 2119 1158 2123 1162
rect 2215 1158 2219 1162
rect 2311 1158 2315 1162
rect 2415 1158 2419 1162
rect 2535 1158 2539 1162
rect 2655 1158 2659 1162
rect 2783 1158 2787 1162
rect 2919 1158 2923 1162
rect 3063 1158 3067 1162
rect 3207 1158 3211 1162
rect 3351 1158 3355 1162
rect 3503 1158 3507 1162
rect 111 1151 115 1155
rect 135 1148 139 1152
rect 303 1148 307 1152
rect 479 1148 483 1152
rect 663 1148 667 1152
rect 839 1148 843 1152
rect 999 1148 1003 1152
rect 1151 1148 1155 1152
rect 1287 1148 1291 1152
rect 1407 1148 1411 1152
rect 1527 1148 1531 1152
rect 1647 1148 1651 1152
rect 1743 1148 1747 1152
rect 1831 1151 1835 1155
rect 1903 1118 1907 1122
rect 2127 1118 2131 1122
rect 2359 1118 2363 1122
rect 2575 1118 2579 1122
rect 2775 1118 2779 1122
rect 2967 1118 2971 1122
rect 3159 1118 3163 1122
rect 3343 1118 3347 1122
rect 3511 1118 3515 1122
rect 111 1101 115 1105
rect 135 1104 139 1108
rect 247 1104 251 1108
rect 383 1104 387 1108
rect 519 1104 523 1108
rect 647 1104 651 1108
rect 775 1104 779 1108
rect 895 1104 899 1108
rect 1015 1104 1019 1108
rect 1135 1104 1139 1108
rect 1255 1104 1259 1108
rect 1375 1104 1379 1108
rect 1503 1104 1507 1108
rect 1631 1104 1635 1108
rect 1743 1104 1747 1108
rect 1831 1101 1835 1105
rect 1871 1100 1875 1104
rect 3591 1100 3595 1104
rect 111 1084 115 1088
rect 1831 1084 1835 1088
rect 1871 1083 1875 1087
rect 1895 1080 1899 1084
rect 2119 1080 2123 1084
rect 2351 1080 2355 1084
rect 2567 1080 2571 1084
rect 2767 1080 2771 1084
rect 2959 1080 2963 1084
rect 3151 1080 3155 1084
rect 3335 1080 3339 1084
rect 3503 1080 3507 1084
rect 3591 1083 3595 1087
rect 143 1066 147 1070
rect 255 1066 259 1070
rect 391 1066 395 1070
rect 527 1066 531 1070
rect 655 1066 659 1070
rect 783 1066 787 1070
rect 903 1066 907 1070
rect 1023 1066 1027 1070
rect 1143 1066 1147 1070
rect 1263 1066 1267 1070
rect 1383 1066 1387 1070
rect 1511 1066 1515 1070
rect 1639 1066 1643 1070
rect 1751 1066 1755 1070
rect 1871 1033 1875 1037
rect 1895 1036 1899 1040
rect 2015 1036 2019 1040
rect 2167 1036 2171 1040
rect 2327 1036 2331 1040
rect 2487 1036 2491 1040
rect 2639 1036 2643 1040
rect 2791 1036 2795 1040
rect 2935 1036 2939 1040
rect 3079 1036 3083 1040
rect 3223 1036 3227 1040
rect 3375 1036 3379 1040
rect 3503 1036 3507 1040
rect 3591 1033 3595 1037
rect 143 1022 147 1026
rect 239 1022 243 1026
rect 359 1022 363 1026
rect 471 1022 475 1026
rect 575 1022 579 1026
rect 671 1022 675 1026
rect 767 1022 771 1026
rect 855 1022 859 1026
rect 943 1022 947 1026
rect 1031 1022 1035 1026
rect 1127 1022 1131 1026
rect 1223 1022 1227 1026
rect 1871 1016 1875 1020
rect 3591 1016 3595 1020
rect 111 1004 115 1008
rect 1831 1004 1835 1008
rect 1903 998 1907 1002
rect 2023 998 2027 1002
rect 2175 998 2179 1002
rect 2335 998 2339 1002
rect 2495 998 2499 1002
rect 2647 998 2651 1002
rect 2799 998 2803 1002
rect 2943 998 2947 1002
rect 3087 998 3091 1002
rect 3231 998 3235 1002
rect 3383 998 3387 1002
rect 3511 998 3515 1002
rect 111 987 115 991
rect 135 984 139 988
rect 231 984 235 988
rect 351 984 355 988
rect 463 984 467 988
rect 567 984 571 988
rect 663 984 667 988
rect 759 984 763 988
rect 847 984 851 988
rect 935 984 939 988
rect 1023 984 1027 988
rect 1119 984 1123 988
rect 1215 984 1219 988
rect 1831 987 1835 991
rect 1903 962 1907 966
rect 1983 962 1987 966
rect 2079 962 2083 966
rect 2199 962 2203 966
rect 2335 962 2339 966
rect 2479 962 2483 966
rect 2631 962 2635 966
rect 2791 962 2795 966
rect 2967 962 2971 966
rect 3151 962 3155 966
rect 3343 962 3347 966
rect 3511 962 3515 966
rect 1871 944 1875 948
rect 3591 944 3595 948
rect 111 925 115 929
rect 135 928 139 932
rect 263 928 267 932
rect 415 928 419 932
rect 559 928 563 932
rect 703 928 707 932
rect 839 928 843 932
rect 975 928 979 932
rect 1103 928 1107 932
rect 1223 928 1227 932
rect 1335 928 1339 932
rect 1439 928 1443 932
rect 1543 928 1547 932
rect 1655 928 1659 932
rect 1743 928 1747 932
rect 1831 925 1835 929
rect 1871 927 1875 931
rect 1895 924 1899 928
rect 1975 924 1979 928
rect 2071 924 2075 928
rect 2191 924 2195 928
rect 2327 924 2331 928
rect 2471 924 2475 928
rect 2623 924 2627 928
rect 2783 924 2787 928
rect 2959 924 2963 928
rect 3143 924 3147 928
rect 3335 924 3339 928
rect 3503 924 3507 928
rect 3591 927 3595 931
rect 111 908 115 912
rect 1831 908 1835 912
rect 143 890 147 894
rect 271 890 275 894
rect 423 890 427 894
rect 567 890 571 894
rect 711 890 715 894
rect 847 890 851 894
rect 983 890 987 894
rect 1111 890 1115 894
rect 1231 890 1235 894
rect 1343 890 1347 894
rect 1447 890 1451 894
rect 1551 890 1555 894
rect 1663 890 1667 894
rect 1751 890 1755 894
rect 1871 865 1875 869
rect 1919 868 1923 872
rect 2095 868 2099 872
rect 2271 868 2275 872
rect 2455 868 2459 872
rect 2655 868 2659 872
rect 2863 868 2867 872
rect 3079 868 3083 872
rect 3303 868 3307 872
rect 3503 868 3507 872
rect 3591 865 3595 869
rect 143 854 147 858
rect 247 854 251 858
rect 383 854 387 858
rect 519 854 523 858
rect 663 854 667 858
rect 815 854 819 858
rect 959 854 963 858
rect 1103 854 1107 858
rect 1247 854 1251 858
rect 1383 854 1387 858
rect 1511 854 1515 858
rect 1639 854 1643 858
rect 1751 854 1755 858
rect 1871 848 1875 852
rect 3591 848 3595 852
rect 111 836 115 840
rect 1831 836 1835 840
rect 1927 830 1931 834
rect 2103 830 2107 834
rect 2279 830 2283 834
rect 2463 830 2467 834
rect 2663 830 2667 834
rect 2871 830 2875 834
rect 3087 830 3091 834
rect 3311 830 3315 834
rect 3511 830 3515 834
rect 111 819 115 823
rect 135 816 139 820
rect 239 816 243 820
rect 375 816 379 820
rect 511 816 515 820
rect 655 816 659 820
rect 807 816 811 820
rect 951 816 955 820
rect 1095 816 1099 820
rect 1239 816 1243 820
rect 1375 816 1379 820
rect 1503 816 1507 820
rect 1631 816 1635 820
rect 1743 816 1747 820
rect 1831 819 1835 823
rect 1903 798 1907 802
rect 2015 798 2019 802
rect 2167 798 2171 802
rect 2327 798 2331 802
rect 2487 798 2491 802
rect 2647 798 2651 802
rect 2807 798 2811 802
rect 2959 798 2963 802
rect 3103 798 3107 802
rect 3247 798 3251 802
rect 3391 798 3395 802
rect 3511 798 3515 802
rect 1871 780 1875 784
rect 3591 780 3595 784
rect 111 757 115 761
rect 135 760 139 764
rect 215 760 219 764
rect 303 760 307 764
rect 415 760 419 764
rect 543 760 547 764
rect 687 760 691 764
rect 839 760 843 764
rect 991 760 995 764
rect 1143 760 1147 764
rect 1295 760 1299 764
rect 1447 760 1451 764
rect 1607 760 1611 764
rect 1871 763 1875 767
rect 1831 757 1835 761
rect 1895 760 1899 764
rect 2007 760 2011 764
rect 2159 760 2163 764
rect 2319 760 2323 764
rect 2479 760 2483 764
rect 2639 760 2643 764
rect 2799 760 2803 764
rect 2951 760 2955 764
rect 3095 760 3099 764
rect 3239 760 3243 764
rect 3383 760 3387 764
rect 3503 760 3507 764
rect 3591 763 3595 767
rect 111 740 115 744
rect 1831 740 1835 744
rect 143 722 147 726
rect 223 722 227 726
rect 311 722 315 726
rect 423 722 427 726
rect 551 722 555 726
rect 695 722 699 726
rect 847 722 851 726
rect 999 722 1003 726
rect 1151 722 1155 726
rect 1303 722 1307 726
rect 1455 722 1459 726
rect 1615 722 1619 726
rect 1871 713 1875 717
rect 1967 716 1971 720
rect 2063 716 2067 720
rect 2175 716 2179 720
rect 2303 716 2307 720
rect 2447 716 2451 720
rect 2599 716 2603 720
rect 2751 716 2755 720
rect 2903 716 2907 720
rect 3055 716 3059 720
rect 3207 716 3211 720
rect 3359 716 3363 720
rect 3503 716 3507 720
rect 3591 713 3595 717
rect 1871 696 1875 700
rect 3591 696 3595 700
rect 231 682 235 686
rect 319 682 323 686
rect 423 682 427 686
rect 543 682 547 686
rect 679 682 683 686
rect 815 682 819 686
rect 951 682 955 686
rect 1087 682 1091 686
rect 1215 682 1219 686
rect 1335 682 1339 686
rect 1455 682 1459 686
rect 1583 682 1587 686
rect 1975 678 1979 682
rect 2071 678 2075 682
rect 2183 678 2187 682
rect 2311 678 2315 682
rect 2455 678 2459 682
rect 2607 678 2611 682
rect 2759 678 2763 682
rect 2911 678 2915 682
rect 3063 678 3067 682
rect 3215 678 3219 682
rect 3367 678 3371 682
rect 3511 678 3515 682
rect 111 664 115 668
rect 1831 664 1835 668
rect 111 647 115 651
rect 223 644 227 648
rect 311 644 315 648
rect 415 644 419 648
rect 535 644 539 648
rect 671 644 675 648
rect 807 644 811 648
rect 943 644 947 648
rect 1079 644 1083 648
rect 1207 644 1211 648
rect 1327 644 1331 648
rect 1447 644 1451 648
rect 1575 644 1579 648
rect 1831 647 1835 651
rect 2175 646 2179 650
rect 2271 646 2275 650
rect 2375 646 2379 650
rect 2487 646 2491 650
rect 2607 646 2611 650
rect 2735 646 2739 650
rect 2863 646 2867 650
rect 2991 646 2995 650
rect 3119 646 3123 650
rect 3247 646 3251 650
rect 3375 646 3379 650
rect 3511 646 3515 650
rect 1871 628 1875 632
rect 3591 628 3595 632
rect 1871 611 1875 615
rect 2167 608 2171 612
rect 2263 608 2267 612
rect 2367 608 2371 612
rect 2479 608 2483 612
rect 2599 608 2603 612
rect 2727 608 2731 612
rect 2855 608 2859 612
rect 2983 608 2987 612
rect 3111 608 3115 612
rect 3239 608 3243 612
rect 3367 608 3371 612
rect 3503 608 3507 612
rect 3591 611 3595 615
rect 111 589 115 593
rect 447 592 451 596
rect 527 592 531 596
rect 607 592 611 596
rect 687 592 691 596
rect 775 592 779 596
rect 871 592 875 596
rect 959 592 963 596
rect 1047 592 1051 596
rect 1143 592 1147 596
rect 1239 592 1243 596
rect 1335 592 1339 596
rect 1431 592 1435 596
rect 1831 589 1835 593
rect 111 572 115 576
rect 1831 572 1835 576
rect 1871 561 1875 565
rect 2263 564 2267 568
rect 2343 564 2347 568
rect 2423 564 2427 568
rect 2503 564 2507 568
rect 2591 564 2595 568
rect 2695 564 2699 568
rect 2815 564 2819 568
rect 2959 564 2963 568
rect 3111 564 3115 568
rect 3279 564 3283 568
rect 3447 564 3451 568
rect 3591 561 3595 565
rect 455 554 459 558
rect 535 554 539 558
rect 615 554 619 558
rect 695 554 699 558
rect 783 554 787 558
rect 879 554 883 558
rect 967 554 971 558
rect 1055 554 1059 558
rect 1151 554 1155 558
rect 1247 554 1251 558
rect 1343 554 1347 558
rect 1439 554 1443 558
rect 1871 544 1875 548
rect 3591 544 3595 548
rect 2271 526 2275 530
rect 2351 526 2355 530
rect 2431 526 2435 530
rect 2511 526 2515 530
rect 2599 526 2603 530
rect 2703 526 2707 530
rect 2823 526 2827 530
rect 2967 526 2971 530
rect 3119 526 3123 530
rect 3287 526 3291 530
rect 3455 526 3459 530
rect 335 510 339 514
rect 423 510 427 514
rect 511 510 515 514
rect 591 510 595 514
rect 671 510 675 514
rect 751 510 755 514
rect 839 510 843 514
rect 927 510 931 514
rect 1015 510 1019 514
rect 1103 510 1107 514
rect 1191 510 1195 514
rect 1279 510 1283 514
rect 111 492 115 496
rect 1831 492 1835 496
rect 2191 486 2195 490
rect 2287 486 2291 490
rect 2383 486 2387 490
rect 2487 486 2491 490
rect 2583 486 2587 490
rect 2687 486 2691 490
rect 2791 486 2795 490
rect 2911 486 2915 490
rect 3039 486 3043 490
rect 3175 486 3179 490
rect 3319 486 3323 490
rect 3471 486 3475 490
rect 111 475 115 479
rect 327 472 331 476
rect 415 472 419 476
rect 503 472 507 476
rect 583 472 587 476
rect 663 472 667 476
rect 743 472 747 476
rect 831 472 835 476
rect 919 472 923 476
rect 1007 472 1011 476
rect 1095 472 1099 476
rect 1183 472 1187 476
rect 1271 472 1275 476
rect 1831 475 1835 479
rect 1871 468 1875 472
rect 3591 468 3595 472
rect 1871 451 1875 455
rect 2183 448 2187 452
rect 2279 448 2283 452
rect 2375 448 2379 452
rect 2479 448 2483 452
rect 2575 448 2579 452
rect 2679 448 2683 452
rect 2783 448 2787 452
rect 2903 448 2907 452
rect 3031 448 3035 452
rect 3167 448 3171 452
rect 3311 448 3315 452
rect 3463 448 3467 452
rect 3591 451 3595 455
rect 111 417 115 421
rect 223 420 227 424
rect 335 420 339 424
rect 447 420 451 424
rect 559 420 563 424
rect 663 420 667 424
rect 759 420 763 424
rect 847 420 851 424
rect 935 420 939 424
rect 1023 420 1027 424
rect 1111 420 1115 424
rect 1199 420 1203 424
rect 1295 420 1299 424
rect 1831 417 1835 421
rect 111 400 115 404
rect 1831 400 1835 404
rect 1871 397 1875 401
rect 1975 400 1979 404
rect 2063 400 2067 404
rect 2159 400 2163 404
rect 2255 400 2259 404
rect 2359 400 2363 404
rect 2471 400 2475 404
rect 2607 400 2611 404
rect 2759 400 2763 404
rect 2927 400 2931 404
rect 3111 400 3115 404
rect 3303 400 3307 404
rect 3495 400 3499 404
rect 3591 397 3595 401
rect 231 382 235 386
rect 343 382 347 386
rect 455 382 459 386
rect 567 382 571 386
rect 671 382 675 386
rect 767 382 771 386
rect 855 382 859 386
rect 943 382 947 386
rect 1031 382 1035 386
rect 1119 382 1123 386
rect 1207 382 1211 386
rect 1303 382 1307 386
rect 1871 380 1875 384
rect 3591 380 3595 384
rect 1983 362 1987 366
rect 2071 362 2075 366
rect 2167 362 2171 366
rect 2263 362 2267 366
rect 2367 362 2371 366
rect 2479 362 2483 366
rect 2615 362 2619 366
rect 2767 362 2771 366
rect 2935 362 2939 366
rect 3119 362 3123 366
rect 3311 362 3315 366
rect 3503 362 3507 366
rect 143 338 147 342
rect 263 338 267 342
rect 399 338 403 342
rect 535 338 539 342
rect 671 338 675 342
rect 791 338 795 342
rect 911 338 915 342
rect 1023 338 1027 342
rect 1127 338 1131 342
rect 1231 338 1235 342
rect 1335 338 1339 342
rect 1439 338 1443 342
rect 2215 326 2219 330
rect 2295 326 2299 330
rect 2383 326 2387 330
rect 2479 326 2483 330
rect 2591 326 2595 330
rect 2719 326 2723 330
rect 2847 326 2851 330
rect 2983 326 2987 330
rect 3119 326 3123 330
rect 3255 326 3259 330
rect 3391 326 3395 330
rect 3511 326 3515 330
rect 111 320 115 324
rect 1831 320 1835 324
rect 1871 308 1875 312
rect 111 303 115 307
rect 3591 308 3595 312
rect 135 300 139 304
rect 255 300 259 304
rect 391 300 395 304
rect 527 300 531 304
rect 663 300 667 304
rect 783 300 787 304
rect 903 300 907 304
rect 1015 300 1019 304
rect 1119 300 1123 304
rect 1223 300 1227 304
rect 1327 300 1331 304
rect 1431 300 1435 304
rect 1831 303 1835 307
rect 1871 291 1875 295
rect 2207 288 2211 292
rect 2287 288 2291 292
rect 2375 288 2379 292
rect 2471 288 2475 292
rect 2583 288 2587 292
rect 2711 288 2715 292
rect 2839 288 2843 292
rect 2975 288 2979 292
rect 3111 288 3115 292
rect 3247 288 3251 292
rect 3383 288 3387 292
rect 3503 288 3507 292
rect 3591 291 3595 295
rect 111 245 115 249
rect 135 248 139 252
rect 247 248 251 252
rect 391 248 395 252
rect 543 248 547 252
rect 695 248 699 252
rect 847 248 851 252
rect 991 248 995 252
rect 1119 248 1123 252
rect 1239 248 1243 252
rect 1359 248 1363 252
rect 1479 248 1483 252
rect 1599 248 1603 252
rect 1831 245 1835 249
rect 1871 237 1875 241
rect 1991 240 1995 244
rect 2119 240 2123 244
rect 2255 240 2259 244
rect 2391 240 2395 244
rect 2535 240 2539 244
rect 2679 240 2683 244
rect 2815 240 2819 244
rect 2951 240 2955 244
rect 3095 240 3099 244
rect 3239 240 3243 244
rect 3383 240 3387 244
rect 3503 240 3507 244
rect 3591 237 3595 241
rect 111 228 115 232
rect 1831 228 1835 232
rect 1871 220 1875 224
rect 3591 220 3595 224
rect 143 210 147 214
rect 255 210 259 214
rect 399 210 403 214
rect 551 210 555 214
rect 703 210 707 214
rect 855 210 859 214
rect 999 210 1003 214
rect 1127 210 1131 214
rect 1247 210 1251 214
rect 1367 210 1371 214
rect 1487 210 1491 214
rect 1607 210 1611 214
rect 1999 202 2003 206
rect 2127 202 2131 206
rect 2263 202 2267 206
rect 2399 202 2403 206
rect 2543 202 2547 206
rect 2687 202 2691 206
rect 2823 202 2827 206
rect 2959 202 2963 206
rect 3103 202 3107 206
rect 3247 202 3251 206
rect 3391 202 3395 206
rect 3511 202 3515 206
rect 1903 158 1907 162
rect 1983 158 1987 162
rect 2087 158 2091 162
rect 2215 158 2219 162
rect 2351 158 2355 162
rect 2487 158 2491 162
rect 2623 158 2627 162
rect 2743 158 2747 162
rect 2855 158 2859 162
rect 2959 158 2963 162
rect 3063 158 3067 162
rect 3159 158 3163 162
rect 3247 158 3251 162
rect 3343 158 3347 162
rect 3431 158 3435 162
rect 3511 158 3515 162
rect 143 142 147 146
rect 223 142 227 146
rect 303 142 307 146
rect 383 142 387 146
rect 463 142 467 146
rect 543 142 547 146
rect 623 142 627 146
rect 703 142 707 146
rect 783 142 787 146
rect 863 142 867 146
rect 943 142 947 146
rect 1023 142 1027 146
rect 1103 142 1107 146
rect 1183 142 1187 146
rect 1263 142 1267 146
rect 1343 142 1347 146
rect 1423 142 1427 146
rect 1511 142 1515 146
rect 1591 142 1595 146
rect 1671 142 1675 146
rect 1751 142 1755 146
rect 1871 140 1875 144
rect 3591 140 3595 144
rect 111 124 115 128
rect 1831 124 1835 128
rect 1871 123 1875 127
rect 1895 120 1899 124
rect 1975 120 1979 124
rect 2079 120 2083 124
rect 2207 120 2211 124
rect 2343 120 2347 124
rect 2479 120 2483 124
rect 2615 120 2619 124
rect 2735 120 2739 124
rect 2847 120 2851 124
rect 2951 120 2955 124
rect 3055 120 3059 124
rect 3151 120 3155 124
rect 3239 120 3243 124
rect 3335 120 3339 124
rect 3423 120 3427 124
rect 3503 120 3507 124
rect 3591 123 3595 127
rect 111 107 115 111
rect 135 104 139 108
rect 215 104 219 108
rect 295 104 299 108
rect 375 104 379 108
rect 455 104 459 108
rect 535 104 539 108
rect 615 104 619 108
rect 695 104 699 108
rect 775 104 779 108
rect 855 104 859 108
rect 935 104 939 108
rect 1015 104 1019 108
rect 1095 104 1099 108
rect 1175 104 1179 108
rect 1255 104 1259 108
rect 1335 104 1339 108
rect 1415 104 1419 108
rect 1503 104 1507 108
rect 1583 104 1587 108
rect 1663 104 1667 108
rect 1743 104 1747 108
rect 1831 107 1835 111
<< m3 >>
rect 111 3670 115 3671
rect 111 3665 115 3666
rect 135 3670 139 3671
rect 135 3665 139 3666
rect 215 3670 219 3671
rect 215 3665 219 3666
rect 295 3670 299 3671
rect 295 3665 299 3666
rect 1831 3670 1835 3671
rect 1831 3665 1835 3666
rect 112 3646 114 3665
rect 136 3649 138 3665
rect 216 3649 218 3665
rect 296 3649 298 3665
rect 134 3648 140 3649
rect 110 3645 116 3646
rect 110 3641 111 3645
rect 115 3641 116 3645
rect 134 3644 135 3648
rect 139 3644 140 3648
rect 134 3643 140 3644
rect 214 3648 220 3649
rect 214 3644 215 3648
rect 219 3644 220 3648
rect 214 3643 220 3644
rect 294 3648 300 3649
rect 294 3644 295 3648
rect 299 3644 300 3648
rect 1832 3646 1834 3665
rect 294 3643 300 3644
rect 1830 3645 1836 3646
rect 110 3640 116 3641
rect 1830 3641 1831 3645
rect 1835 3641 1836 3645
rect 1830 3640 1836 3641
rect 110 3628 116 3629
rect 110 3624 111 3628
rect 115 3624 116 3628
rect 110 3623 116 3624
rect 1830 3628 1836 3629
rect 1830 3624 1831 3628
rect 1835 3624 1836 3628
rect 1830 3623 1836 3624
rect 112 3595 114 3623
rect 142 3610 148 3611
rect 142 3606 143 3610
rect 147 3606 148 3610
rect 142 3605 148 3606
rect 222 3610 228 3611
rect 222 3606 223 3610
rect 227 3606 228 3610
rect 222 3605 228 3606
rect 302 3610 308 3611
rect 302 3606 303 3610
rect 307 3606 308 3610
rect 302 3605 308 3606
rect 144 3595 146 3605
rect 224 3595 226 3605
rect 304 3595 306 3605
rect 1832 3595 1834 3623
rect 1871 3602 1875 3603
rect 1871 3597 1875 3598
rect 2063 3602 2067 3603
rect 2063 3597 2067 3598
rect 2151 3602 2155 3603
rect 2151 3597 2155 3598
rect 2255 3602 2259 3603
rect 2255 3597 2259 3598
rect 2367 3602 2371 3603
rect 2367 3597 2371 3598
rect 2479 3602 2483 3603
rect 2479 3597 2483 3598
rect 2591 3602 2595 3603
rect 2591 3597 2595 3598
rect 2703 3602 2707 3603
rect 2703 3597 2707 3598
rect 2815 3602 2819 3603
rect 2815 3597 2819 3598
rect 2919 3602 2923 3603
rect 2919 3597 2923 3598
rect 3015 3602 3019 3603
rect 3015 3597 3019 3598
rect 3111 3602 3115 3603
rect 3111 3597 3115 3598
rect 3207 3602 3211 3603
rect 3207 3597 3211 3598
rect 3303 3602 3307 3603
rect 3303 3597 3307 3598
rect 3399 3602 3403 3603
rect 3399 3597 3403 3598
rect 3591 3602 3595 3603
rect 3591 3597 3595 3598
rect 111 3594 115 3595
rect 111 3589 115 3590
rect 143 3594 147 3595
rect 143 3589 147 3590
rect 223 3594 227 3595
rect 223 3589 227 3590
rect 303 3594 307 3595
rect 303 3589 307 3590
rect 343 3594 347 3595
rect 343 3589 347 3590
rect 471 3594 475 3595
rect 471 3589 475 3590
rect 607 3594 611 3595
rect 607 3589 611 3590
rect 743 3594 747 3595
rect 743 3589 747 3590
rect 879 3594 883 3595
rect 879 3589 883 3590
rect 999 3594 1003 3595
rect 999 3589 1003 3590
rect 1111 3594 1115 3595
rect 1111 3589 1115 3590
rect 1223 3594 1227 3595
rect 1223 3589 1227 3590
rect 1327 3594 1331 3595
rect 1327 3589 1331 3590
rect 1423 3594 1427 3595
rect 1423 3589 1427 3590
rect 1527 3594 1531 3595
rect 1527 3589 1531 3590
rect 1631 3594 1635 3595
rect 1631 3589 1635 3590
rect 1831 3594 1835 3595
rect 1831 3589 1835 3590
rect 112 3561 114 3589
rect 144 3579 146 3589
rect 224 3579 226 3589
rect 344 3579 346 3589
rect 472 3579 474 3589
rect 608 3579 610 3589
rect 744 3579 746 3589
rect 880 3579 882 3589
rect 1000 3579 1002 3589
rect 1112 3579 1114 3589
rect 1224 3579 1226 3589
rect 1328 3579 1330 3589
rect 1424 3579 1426 3589
rect 1528 3579 1530 3589
rect 1632 3579 1634 3589
rect 142 3578 148 3579
rect 142 3574 143 3578
rect 147 3574 148 3578
rect 142 3573 148 3574
rect 222 3578 228 3579
rect 222 3574 223 3578
rect 227 3574 228 3578
rect 222 3573 228 3574
rect 342 3578 348 3579
rect 342 3574 343 3578
rect 347 3574 348 3578
rect 342 3573 348 3574
rect 470 3578 476 3579
rect 470 3574 471 3578
rect 475 3574 476 3578
rect 470 3573 476 3574
rect 606 3578 612 3579
rect 606 3574 607 3578
rect 611 3574 612 3578
rect 606 3573 612 3574
rect 742 3578 748 3579
rect 742 3574 743 3578
rect 747 3574 748 3578
rect 742 3573 748 3574
rect 878 3578 884 3579
rect 878 3574 879 3578
rect 883 3574 884 3578
rect 878 3573 884 3574
rect 998 3578 1004 3579
rect 998 3574 999 3578
rect 1003 3574 1004 3578
rect 998 3573 1004 3574
rect 1110 3578 1116 3579
rect 1110 3574 1111 3578
rect 1115 3574 1116 3578
rect 1110 3573 1116 3574
rect 1222 3578 1228 3579
rect 1222 3574 1223 3578
rect 1227 3574 1228 3578
rect 1222 3573 1228 3574
rect 1326 3578 1332 3579
rect 1326 3574 1327 3578
rect 1331 3574 1332 3578
rect 1326 3573 1332 3574
rect 1422 3578 1428 3579
rect 1422 3574 1423 3578
rect 1427 3574 1428 3578
rect 1422 3573 1428 3574
rect 1526 3578 1532 3579
rect 1526 3574 1527 3578
rect 1531 3574 1532 3578
rect 1526 3573 1532 3574
rect 1630 3578 1636 3579
rect 1630 3574 1631 3578
rect 1635 3574 1636 3578
rect 1630 3573 1636 3574
rect 1832 3561 1834 3589
rect 1872 3569 1874 3597
rect 2064 3587 2066 3597
rect 2152 3587 2154 3597
rect 2256 3587 2258 3597
rect 2368 3587 2370 3597
rect 2480 3587 2482 3597
rect 2592 3587 2594 3597
rect 2704 3587 2706 3597
rect 2816 3587 2818 3597
rect 2920 3587 2922 3597
rect 3016 3587 3018 3597
rect 3112 3587 3114 3597
rect 3208 3587 3210 3597
rect 3304 3587 3306 3597
rect 3400 3587 3402 3597
rect 2062 3586 2068 3587
rect 2062 3582 2063 3586
rect 2067 3582 2068 3586
rect 2062 3581 2068 3582
rect 2150 3586 2156 3587
rect 2150 3582 2151 3586
rect 2155 3582 2156 3586
rect 2150 3581 2156 3582
rect 2254 3586 2260 3587
rect 2254 3582 2255 3586
rect 2259 3582 2260 3586
rect 2254 3581 2260 3582
rect 2366 3586 2372 3587
rect 2366 3582 2367 3586
rect 2371 3582 2372 3586
rect 2366 3581 2372 3582
rect 2478 3586 2484 3587
rect 2478 3582 2479 3586
rect 2483 3582 2484 3586
rect 2478 3581 2484 3582
rect 2590 3586 2596 3587
rect 2590 3582 2591 3586
rect 2595 3582 2596 3586
rect 2590 3581 2596 3582
rect 2702 3586 2708 3587
rect 2702 3582 2703 3586
rect 2707 3582 2708 3586
rect 2702 3581 2708 3582
rect 2814 3586 2820 3587
rect 2814 3582 2815 3586
rect 2819 3582 2820 3586
rect 2814 3581 2820 3582
rect 2918 3586 2924 3587
rect 2918 3582 2919 3586
rect 2923 3582 2924 3586
rect 2918 3581 2924 3582
rect 3014 3586 3020 3587
rect 3014 3582 3015 3586
rect 3019 3582 3020 3586
rect 3014 3581 3020 3582
rect 3110 3586 3116 3587
rect 3110 3582 3111 3586
rect 3115 3582 3116 3586
rect 3110 3581 3116 3582
rect 3206 3586 3212 3587
rect 3206 3582 3207 3586
rect 3211 3582 3212 3586
rect 3206 3581 3212 3582
rect 3302 3586 3308 3587
rect 3302 3582 3303 3586
rect 3307 3582 3308 3586
rect 3302 3581 3308 3582
rect 3398 3586 3404 3587
rect 3398 3582 3399 3586
rect 3403 3582 3404 3586
rect 3398 3581 3404 3582
rect 3592 3569 3594 3597
rect 1870 3568 1876 3569
rect 1870 3564 1871 3568
rect 1875 3564 1876 3568
rect 1870 3563 1876 3564
rect 3590 3568 3596 3569
rect 3590 3564 3591 3568
rect 3595 3564 3596 3568
rect 3590 3563 3596 3564
rect 110 3560 116 3561
rect 110 3556 111 3560
rect 115 3556 116 3560
rect 110 3555 116 3556
rect 1830 3560 1836 3561
rect 1830 3556 1831 3560
rect 1835 3556 1836 3560
rect 1830 3555 1836 3556
rect 1870 3551 1876 3552
rect 1870 3547 1871 3551
rect 1875 3547 1876 3551
rect 3590 3551 3596 3552
rect 1870 3546 1876 3547
rect 2054 3548 2060 3549
rect 110 3543 116 3544
rect 110 3539 111 3543
rect 115 3539 116 3543
rect 1830 3543 1836 3544
rect 110 3538 116 3539
rect 134 3540 140 3541
rect 112 3519 114 3538
rect 134 3536 135 3540
rect 139 3536 140 3540
rect 134 3535 140 3536
rect 214 3540 220 3541
rect 214 3536 215 3540
rect 219 3536 220 3540
rect 214 3535 220 3536
rect 334 3540 340 3541
rect 334 3536 335 3540
rect 339 3536 340 3540
rect 334 3535 340 3536
rect 462 3540 468 3541
rect 462 3536 463 3540
rect 467 3536 468 3540
rect 462 3535 468 3536
rect 598 3540 604 3541
rect 598 3536 599 3540
rect 603 3536 604 3540
rect 598 3535 604 3536
rect 734 3540 740 3541
rect 734 3536 735 3540
rect 739 3536 740 3540
rect 734 3535 740 3536
rect 870 3540 876 3541
rect 870 3536 871 3540
rect 875 3536 876 3540
rect 870 3535 876 3536
rect 990 3540 996 3541
rect 990 3536 991 3540
rect 995 3536 996 3540
rect 990 3535 996 3536
rect 1102 3540 1108 3541
rect 1102 3536 1103 3540
rect 1107 3536 1108 3540
rect 1102 3535 1108 3536
rect 1214 3540 1220 3541
rect 1214 3536 1215 3540
rect 1219 3536 1220 3540
rect 1214 3535 1220 3536
rect 1318 3540 1324 3541
rect 1318 3536 1319 3540
rect 1323 3536 1324 3540
rect 1318 3535 1324 3536
rect 1414 3540 1420 3541
rect 1414 3536 1415 3540
rect 1419 3536 1420 3540
rect 1414 3535 1420 3536
rect 1518 3540 1524 3541
rect 1518 3536 1519 3540
rect 1523 3536 1524 3540
rect 1518 3535 1524 3536
rect 1622 3540 1628 3541
rect 1622 3536 1623 3540
rect 1627 3536 1628 3540
rect 1830 3539 1831 3543
rect 1835 3539 1836 3543
rect 1830 3538 1836 3539
rect 1622 3535 1628 3536
rect 136 3519 138 3535
rect 216 3519 218 3535
rect 336 3519 338 3535
rect 464 3519 466 3535
rect 600 3519 602 3535
rect 736 3519 738 3535
rect 872 3519 874 3535
rect 992 3519 994 3535
rect 1104 3519 1106 3535
rect 1216 3519 1218 3535
rect 1320 3519 1322 3535
rect 1416 3519 1418 3535
rect 1520 3519 1522 3535
rect 1624 3519 1626 3535
rect 1832 3519 1834 3538
rect 1872 3527 1874 3546
rect 2054 3544 2055 3548
rect 2059 3544 2060 3548
rect 2054 3543 2060 3544
rect 2142 3548 2148 3549
rect 2142 3544 2143 3548
rect 2147 3544 2148 3548
rect 2142 3543 2148 3544
rect 2246 3548 2252 3549
rect 2246 3544 2247 3548
rect 2251 3544 2252 3548
rect 2246 3543 2252 3544
rect 2358 3548 2364 3549
rect 2358 3544 2359 3548
rect 2363 3544 2364 3548
rect 2358 3543 2364 3544
rect 2470 3548 2476 3549
rect 2470 3544 2471 3548
rect 2475 3544 2476 3548
rect 2470 3543 2476 3544
rect 2582 3548 2588 3549
rect 2582 3544 2583 3548
rect 2587 3544 2588 3548
rect 2582 3543 2588 3544
rect 2694 3548 2700 3549
rect 2694 3544 2695 3548
rect 2699 3544 2700 3548
rect 2694 3543 2700 3544
rect 2806 3548 2812 3549
rect 2806 3544 2807 3548
rect 2811 3544 2812 3548
rect 2806 3543 2812 3544
rect 2910 3548 2916 3549
rect 2910 3544 2911 3548
rect 2915 3544 2916 3548
rect 2910 3543 2916 3544
rect 3006 3548 3012 3549
rect 3006 3544 3007 3548
rect 3011 3544 3012 3548
rect 3006 3543 3012 3544
rect 3102 3548 3108 3549
rect 3102 3544 3103 3548
rect 3107 3544 3108 3548
rect 3102 3543 3108 3544
rect 3198 3548 3204 3549
rect 3198 3544 3199 3548
rect 3203 3544 3204 3548
rect 3198 3543 3204 3544
rect 3294 3548 3300 3549
rect 3294 3544 3295 3548
rect 3299 3544 3300 3548
rect 3294 3543 3300 3544
rect 3390 3548 3396 3549
rect 3390 3544 3391 3548
rect 3395 3544 3396 3548
rect 3590 3547 3591 3551
rect 3595 3547 3596 3551
rect 3590 3546 3596 3547
rect 3390 3543 3396 3544
rect 2056 3527 2058 3543
rect 2144 3527 2146 3543
rect 2248 3527 2250 3543
rect 2360 3527 2362 3543
rect 2472 3527 2474 3543
rect 2584 3527 2586 3543
rect 2696 3527 2698 3543
rect 2808 3527 2810 3543
rect 2912 3527 2914 3543
rect 3008 3527 3010 3543
rect 3104 3527 3106 3543
rect 3200 3527 3202 3543
rect 3296 3527 3298 3543
rect 3392 3527 3394 3543
rect 3592 3527 3594 3546
rect 1871 3526 1875 3527
rect 1871 3521 1875 3522
rect 2055 3526 2059 3527
rect 2055 3521 2059 3522
rect 2087 3526 2091 3527
rect 2087 3521 2091 3522
rect 2143 3526 2147 3527
rect 2143 3521 2147 3522
rect 2167 3526 2171 3527
rect 2167 3521 2171 3522
rect 2247 3526 2251 3527
rect 2247 3521 2251 3522
rect 2263 3526 2267 3527
rect 2263 3521 2267 3522
rect 2359 3526 2363 3527
rect 2359 3521 2363 3522
rect 2367 3526 2371 3527
rect 2367 3521 2371 3522
rect 2471 3526 2475 3527
rect 2471 3521 2475 3522
rect 2487 3526 2491 3527
rect 2487 3521 2491 3522
rect 2583 3526 2587 3527
rect 2583 3521 2587 3522
rect 2615 3526 2619 3527
rect 2615 3521 2619 3522
rect 2695 3526 2699 3527
rect 2695 3521 2699 3522
rect 2743 3526 2747 3527
rect 2743 3521 2747 3522
rect 2807 3526 2811 3527
rect 2807 3521 2811 3522
rect 2871 3526 2875 3527
rect 2871 3521 2875 3522
rect 2911 3526 2915 3527
rect 2911 3521 2915 3522
rect 2991 3526 2995 3527
rect 2991 3521 2995 3522
rect 3007 3526 3011 3527
rect 3007 3521 3011 3522
rect 3103 3526 3107 3527
rect 3103 3521 3107 3522
rect 3119 3526 3123 3527
rect 3119 3521 3123 3522
rect 3199 3526 3203 3527
rect 3199 3521 3203 3522
rect 3247 3526 3251 3527
rect 3247 3521 3251 3522
rect 3295 3526 3299 3527
rect 3295 3521 3299 3522
rect 3375 3526 3379 3527
rect 3375 3521 3379 3522
rect 3391 3526 3395 3527
rect 3391 3521 3395 3522
rect 3591 3526 3595 3527
rect 3591 3521 3595 3522
rect 111 3518 115 3519
rect 111 3513 115 3514
rect 135 3518 139 3519
rect 135 3513 139 3514
rect 191 3518 195 3519
rect 191 3513 195 3514
rect 215 3518 219 3519
rect 215 3513 219 3514
rect 327 3518 331 3519
rect 327 3513 331 3514
rect 335 3518 339 3519
rect 335 3513 339 3514
rect 463 3518 467 3519
rect 463 3513 467 3514
rect 471 3518 475 3519
rect 471 3513 475 3514
rect 599 3518 603 3519
rect 599 3513 603 3514
rect 623 3518 627 3519
rect 623 3513 627 3514
rect 735 3518 739 3519
rect 735 3513 739 3514
rect 775 3518 779 3519
rect 775 3513 779 3514
rect 871 3518 875 3519
rect 871 3513 875 3514
rect 919 3518 923 3519
rect 919 3513 923 3514
rect 991 3518 995 3519
rect 991 3513 995 3514
rect 1055 3518 1059 3519
rect 1055 3513 1059 3514
rect 1103 3518 1107 3519
rect 1103 3513 1107 3514
rect 1183 3518 1187 3519
rect 1183 3513 1187 3514
rect 1215 3518 1219 3519
rect 1215 3513 1219 3514
rect 1311 3518 1315 3519
rect 1311 3513 1315 3514
rect 1319 3518 1323 3519
rect 1319 3513 1323 3514
rect 1415 3518 1419 3519
rect 1415 3513 1419 3514
rect 1439 3518 1443 3519
rect 1439 3513 1443 3514
rect 1519 3518 1523 3519
rect 1519 3513 1523 3514
rect 1567 3518 1571 3519
rect 1567 3513 1571 3514
rect 1623 3518 1627 3519
rect 1623 3513 1627 3514
rect 1831 3518 1835 3519
rect 1831 3513 1835 3514
rect 112 3494 114 3513
rect 192 3497 194 3513
rect 328 3497 330 3513
rect 472 3497 474 3513
rect 624 3497 626 3513
rect 776 3497 778 3513
rect 920 3497 922 3513
rect 1056 3497 1058 3513
rect 1184 3497 1186 3513
rect 1312 3497 1314 3513
rect 1440 3497 1442 3513
rect 1568 3497 1570 3513
rect 190 3496 196 3497
rect 110 3493 116 3494
rect 110 3489 111 3493
rect 115 3489 116 3493
rect 190 3492 191 3496
rect 195 3492 196 3496
rect 190 3491 196 3492
rect 326 3496 332 3497
rect 326 3492 327 3496
rect 331 3492 332 3496
rect 326 3491 332 3492
rect 470 3496 476 3497
rect 470 3492 471 3496
rect 475 3492 476 3496
rect 470 3491 476 3492
rect 622 3496 628 3497
rect 622 3492 623 3496
rect 627 3492 628 3496
rect 622 3491 628 3492
rect 774 3496 780 3497
rect 774 3492 775 3496
rect 779 3492 780 3496
rect 774 3491 780 3492
rect 918 3496 924 3497
rect 918 3492 919 3496
rect 923 3492 924 3496
rect 918 3491 924 3492
rect 1054 3496 1060 3497
rect 1054 3492 1055 3496
rect 1059 3492 1060 3496
rect 1054 3491 1060 3492
rect 1182 3496 1188 3497
rect 1182 3492 1183 3496
rect 1187 3492 1188 3496
rect 1182 3491 1188 3492
rect 1310 3496 1316 3497
rect 1310 3492 1311 3496
rect 1315 3492 1316 3496
rect 1310 3491 1316 3492
rect 1438 3496 1444 3497
rect 1438 3492 1439 3496
rect 1443 3492 1444 3496
rect 1438 3491 1444 3492
rect 1566 3496 1572 3497
rect 1566 3492 1567 3496
rect 1571 3492 1572 3496
rect 1832 3494 1834 3513
rect 1872 3502 1874 3521
rect 2088 3505 2090 3521
rect 2168 3505 2170 3521
rect 2264 3505 2266 3521
rect 2368 3505 2370 3521
rect 2488 3505 2490 3521
rect 2616 3505 2618 3521
rect 2744 3505 2746 3521
rect 2872 3505 2874 3521
rect 2992 3505 2994 3521
rect 3120 3505 3122 3521
rect 3248 3505 3250 3521
rect 3376 3505 3378 3521
rect 2086 3504 2092 3505
rect 1870 3501 1876 3502
rect 1870 3497 1871 3501
rect 1875 3497 1876 3501
rect 2086 3500 2087 3504
rect 2091 3500 2092 3504
rect 2086 3499 2092 3500
rect 2166 3504 2172 3505
rect 2166 3500 2167 3504
rect 2171 3500 2172 3504
rect 2166 3499 2172 3500
rect 2262 3504 2268 3505
rect 2262 3500 2263 3504
rect 2267 3500 2268 3504
rect 2262 3499 2268 3500
rect 2366 3504 2372 3505
rect 2366 3500 2367 3504
rect 2371 3500 2372 3504
rect 2366 3499 2372 3500
rect 2486 3504 2492 3505
rect 2486 3500 2487 3504
rect 2491 3500 2492 3504
rect 2486 3499 2492 3500
rect 2614 3504 2620 3505
rect 2614 3500 2615 3504
rect 2619 3500 2620 3504
rect 2614 3499 2620 3500
rect 2742 3504 2748 3505
rect 2742 3500 2743 3504
rect 2747 3500 2748 3504
rect 2742 3499 2748 3500
rect 2870 3504 2876 3505
rect 2870 3500 2871 3504
rect 2875 3500 2876 3504
rect 2870 3499 2876 3500
rect 2990 3504 2996 3505
rect 2990 3500 2991 3504
rect 2995 3500 2996 3504
rect 2990 3499 2996 3500
rect 3118 3504 3124 3505
rect 3118 3500 3119 3504
rect 3123 3500 3124 3504
rect 3118 3499 3124 3500
rect 3246 3504 3252 3505
rect 3246 3500 3247 3504
rect 3251 3500 3252 3504
rect 3246 3499 3252 3500
rect 3374 3504 3380 3505
rect 3374 3500 3375 3504
rect 3379 3500 3380 3504
rect 3592 3502 3594 3521
rect 3374 3499 3380 3500
rect 3590 3501 3596 3502
rect 1870 3496 1876 3497
rect 3590 3497 3591 3501
rect 3595 3497 3596 3501
rect 3590 3496 3596 3497
rect 1566 3491 1572 3492
rect 1830 3493 1836 3494
rect 110 3488 116 3489
rect 1830 3489 1831 3493
rect 1835 3489 1836 3493
rect 1830 3488 1836 3489
rect 1870 3484 1876 3485
rect 1870 3480 1871 3484
rect 1875 3480 1876 3484
rect 1870 3479 1876 3480
rect 3590 3484 3596 3485
rect 3590 3480 3591 3484
rect 3595 3480 3596 3484
rect 3590 3479 3596 3480
rect 110 3476 116 3477
rect 110 3472 111 3476
rect 115 3472 116 3476
rect 110 3471 116 3472
rect 1830 3476 1836 3477
rect 1830 3472 1831 3476
rect 1835 3472 1836 3476
rect 1830 3471 1836 3472
rect 112 3443 114 3471
rect 198 3458 204 3459
rect 198 3454 199 3458
rect 203 3454 204 3458
rect 198 3453 204 3454
rect 334 3458 340 3459
rect 334 3454 335 3458
rect 339 3454 340 3458
rect 334 3453 340 3454
rect 478 3458 484 3459
rect 478 3454 479 3458
rect 483 3454 484 3458
rect 478 3453 484 3454
rect 630 3458 636 3459
rect 630 3454 631 3458
rect 635 3454 636 3458
rect 630 3453 636 3454
rect 782 3458 788 3459
rect 782 3454 783 3458
rect 787 3454 788 3458
rect 782 3453 788 3454
rect 926 3458 932 3459
rect 926 3454 927 3458
rect 931 3454 932 3458
rect 926 3453 932 3454
rect 1062 3458 1068 3459
rect 1062 3454 1063 3458
rect 1067 3454 1068 3458
rect 1062 3453 1068 3454
rect 1190 3458 1196 3459
rect 1190 3454 1191 3458
rect 1195 3454 1196 3458
rect 1190 3453 1196 3454
rect 1318 3458 1324 3459
rect 1318 3454 1319 3458
rect 1323 3454 1324 3458
rect 1318 3453 1324 3454
rect 1446 3458 1452 3459
rect 1446 3454 1447 3458
rect 1451 3454 1452 3458
rect 1446 3453 1452 3454
rect 1574 3458 1580 3459
rect 1574 3454 1575 3458
rect 1579 3454 1580 3458
rect 1574 3453 1580 3454
rect 200 3443 202 3453
rect 336 3443 338 3453
rect 480 3443 482 3453
rect 632 3443 634 3453
rect 784 3443 786 3453
rect 928 3443 930 3453
rect 1064 3443 1066 3453
rect 1192 3443 1194 3453
rect 1320 3443 1322 3453
rect 1448 3443 1450 3453
rect 1576 3443 1578 3453
rect 1832 3443 1834 3471
rect 1872 3443 1874 3479
rect 2094 3466 2100 3467
rect 2094 3462 2095 3466
rect 2099 3462 2100 3466
rect 2094 3461 2100 3462
rect 2174 3466 2180 3467
rect 2174 3462 2175 3466
rect 2179 3462 2180 3466
rect 2174 3461 2180 3462
rect 2270 3466 2276 3467
rect 2270 3462 2271 3466
rect 2275 3462 2276 3466
rect 2270 3461 2276 3462
rect 2374 3466 2380 3467
rect 2374 3462 2375 3466
rect 2379 3462 2380 3466
rect 2374 3461 2380 3462
rect 2494 3466 2500 3467
rect 2494 3462 2495 3466
rect 2499 3462 2500 3466
rect 2494 3461 2500 3462
rect 2622 3466 2628 3467
rect 2622 3462 2623 3466
rect 2627 3462 2628 3466
rect 2622 3461 2628 3462
rect 2750 3466 2756 3467
rect 2750 3462 2751 3466
rect 2755 3462 2756 3466
rect 2750 3461 2756 3462
rect 2878 3466 2884 3467
rect 2878 3462 2879 3466
rect 2883 3462 2884 3466
rect 2878 3461 2884 3462
rect 2998 3466 3004 3467
rect 2998 3462 2999 3466
rect 3003 3462 3004 3466
rect 2998 3461 3004 3462
rect 3126 3466 3132 3467
rect 3126 3462 3127 3466
rect 3131 3462 3132 3466
rect 3126 3461 3132 3462
rect 3254 3466 3260 3467
rect 3254 3462 3255 3466
rect 3259 3462 3260 3466
rect 3254 3461 3260 3462
rect 3382 3466 3388 3467
rect 3382 3462 3383 3466
rect 3387 3462 3388 3466
rect 3382 3461 3388 3462
rect 2096 3443 2098 3461
rect 2176 3443 2178 3461
rect 2272 3443 2274 3461
rect 2376 3443 2378 3461
rect 2496 3443 2498 3461
rect 2624 3443 2626 3461
rect 2752 3443 2754 3461
rect 2880 3443 2882 3461
rect 3000 3443 3002 3461
rect 3128 3443 3130 3461
rect 3256 3443 3258 3461
rect 3384 3443 3386 3461
rect 3592 3443 3594 3479
rect 111 3442 115 3443
rect 111 3437 115 3438
rect 151 3442 155 3443
rect 151 3437 155 3438
rect 199 3442 203 3443
rect 199 3437 203 3438
rect 295 3442 299 3443
rect 295 3437 299 3438
rect 335 3442 339 3443
rect 335 3437 339 3438
rect 455 3442 459 3443
rect 455 3437 459 3438
rect 479 3442 483 3443
rect 479 3437 483 3438
rect 623 3442 627 3443
rect 623 3437 627 3438
rect 631 3442 635 3443
rect 631 3437 635 3438
rect 783 3442 787 3443
rect 783 3437 787 3438
rect 791 3442 795 3443
rect 791 3437 795 3438
rect 927 3442 931 3443
rect 927 3437 931 3438
rect 959 3442 963 3443
rect 959 3437 963 3438
rect 1063 3442 1067 3443
rect 1063 3437 1067 3438
rect 1119 3442 1123 3443
rect 1119 3437 1123 3438
rect 1191 3442 1195 3443
rect 1191 3437 1195 3438
rect 1271 3442 1275 3443
rect 1271 3437 1275 3438
rect 1319 3442 1323 3443
rect 1319 3437 1323 3438
rect 1415 3442 1419 3443
rect 1415 3437 1419 3438
rect 1447 3442 1451 3443
rect 1447 3437 1451 3438
rect 1559 3442 1563 3443
rect 1559 3437 1563 3438
rect 1575 3442 1579 3443
rect 1575 3437 1579 3438
rect 1711 3442 1715 3443
rect 1711 3437 1715 3438
rect 1831 3442 1835 3443
rect 1831 3437 1835 3438
rect 1871 3442 1875 3443
rect 1871 3437 1875 3438
rect 2095 3442 2099 3443
rect 2095 3437 2099 3438
rect 2111 3442 2115 3443
rect 2111 3437 2115 3438
rect 2175 3442 2179 3443
rect 2175 3437 2179 3438
rect 2199 3442 2203 3443
rect 2199 3437 2203 3438
rect 2271 3442 2275 3443
rect 2271 3437 2275 3438
rect 2303 3442 2307 3443
rect 2303 3437 2307 3438
rect 2375 3442 2379 3443
rect 2375 3437 2379 3438
rect 2415 3442 2419 3443
rect 2415 3437 2419 3438
rect 2495 3442 2499 3443
rect 2495 3437 2499 3438
rect 2543 3442 2547 3443
rect 2543 3437 2547 3438
rect 2623 3442 2627 3443
rect 2623 3437 2627 3438
rect 2679 3442 2683 3443
rect 2679 3437 2683 3438
rect 2751 3442 2755 3443
rect 2751 3437 2755 3438
rect 2815 3442 2819 3443
rect 2815 3437 2819 3438
rect 2879 3442 2883 3443
rect 2879 3437 2883 3438
rect 2959 3442 2963 3443
rect 2959 3437 2963 3438
rect 2999 3442 3003 3443
rect 2999 3437 3003 3438
rect 3111 3442 3115 3443
rect 3111 3437 3115 3438
rect 3127 3442 3131 3443
rect 3127 3437 3131 3438
rect 3255 3442 3259 3443
rect 3255 3437 3259 3438
rect 3263 3442 3267 3443
rect 3263 3437 3267 3438
rect 3383 3442 3387 3443
rect 3383 3437 3387 3438
rect 3423 3442 3427 3443
rect 3423 3437 3427 3438
rect 3591 3442 3595 3443
rect 3591 3437 3595 3438
rect 112 3409 114 3437
rect 152 3427 154 3437
rect 296 3427 298 3437
rect 456 3427 458 3437
rect 624 3427 626 3437
rect 792 3427 794 3437
rect 960 3427 962 3437
rect 1120 3427 1122 3437
rect 1272 3427 1274 3437
rect 1416 3427 1418 3437
rect 1560 3427 1562 3437
rect 1712 3427 1714 3437
rect 150 3426 156 3427
rect 150 3422 151 3426
rect 155 3422 156 3426
rect 150 3421 156 3422
rect 294 3426 300 3427
rect 294 3422 295 3426
rect 299 3422 300 3426
rect 294 3421 300 3422
rect 454 3426 460 3427
rect 454 3422 455 3426
rect 459 3422 460 3426
rect 454 3421 460 3422
rect 622 3426 628 3427
rect 622 3422 623 3426
rect 627 3422 628 3426
rect 622 3421 628 3422
rect 790 3426 796 3427
rect 790 3422 791 3426
rect 795 3422 796 3426
rect 790 3421 796 3422
rect 958 3426 964 3427
rect 958 3422 959 3426
rect 963 3422 964 3426
rect 958 3421 964 3422
rect 1118 3426 1124 3427
rect 1118 3422 1119 3426
rect 1123 3422 1124 3426
rect 1118 3421 1124 3422
rect 1270 3426 1276 3427
rect 1270 3422 1271 3426
rect 1275 3422 1276 3426
rect 1270 3421 1276 3422
rect 1414 3426 1420 3427
rect 1414 3422 1415 3426
rect 1419 3422 1420 3426
rect 1414 3421 1420 3422
rect 1558 3426 1564 3427
rect 1558 3422 1559 3426
rect 1563 3422 1564 3426
rect 1558 3421 1564 3422
rect 1710 3426 1716 3427
rect 1710 3422 1711 3426
rect 1715 3422 1716 3426
rect 1710 3421 1716 3422
rect 1832 3409 1834 3437
rect 1872 3409 1874 3437
rect 2112 3427 2114 3437
rect 2200 3427 2202 3437
rect 2304 3427 2306 3437
rect 2416 3427 2418 3437
rect 2544 3427 2546 3437
rect 2680 3427 2682 3437
rect 2816 3427 2818 3437
rect 2960 3427 2962 3437
rect 3112 3427 3114 3437
rect 3264 3427 3266 3437
rect 3424 3427 3426 3437
rect 2110 3426 2116 3427
rect 2110 3422 2111 3426
rect 2115 3422 2116 3426
rect 2110 3421 2116 3422
rect 2198 3426 2204 3427
rect 2198 3422 2199 3426
rect 2203 3422 2204 3426
rect 2198 3421 2204 3422
rect 2302 3426 2308 3427
rect 2302 3422 2303 3426
rect 2307 3422 2308 3426
rect 2302 3421 2308 3422
rect 2414 3426 2420 3427
rect 2414 3422 2415 3426
rect 2419 3422 2420 3426
rect 2414 3421 2420 3422
rect 2542 3426 2548 3427
rect 2542 3422 2543 3426
rect 2547 3422 2548 3426
rect 2542 3421 2548 3422
rect 2678 3426 2684 3427
rect 2678 3422 2679 3426
rect 2683 3422 2684 3426
rect 2678 3421 2684 3422
rect 2814 3426 2820 3427
rect 2814 3422 2815 3426
rect 2819 3422 2820 3426
rect 2814 3421 2820 3422
rect 2958 3426 2964 3427
rect 2958 3422 2959 3426
rect 2963 3422 2964 3426
rect 2958 3421 2964 3422
rect 3110 3426 3116 3427
rect 3110 3422 3111 3426
rect 3115 3422 3116 3426
rect 3110 3421 3116 3422
rect 3262 3426 3268 3427
rect 3262 3422 3263 3426
rect 3267 3422 3268 3426
rect 3262 3421 3268 3422
rect 3422 3426 3428 3427
rect 3422 3422 3423 3426
rect 3427 3422 3428 3426
rect 3422 3421 3428 3422
rect 3592 3409 3594 3437
rect 110 3408 116 3409
rect 110 3404 111 3408
rect 115 3404 116 3408
rect 110 3403 116 3404
rect 1830 3408 1836 3409
rect 1830 3404 1831 3408
rect 1835 3404 1836 3408
rect 1830 3403 1836 3404
rect 1870 3408 1876 3409
rect 1870 3404 1871 3408
rect 1875 3404 1876 3408
rect 1870 3403 1876 3404
rect 3590 3408 3596 3409
rect 3590 3404 3591 3408
rect 3595 3404 3596 3408
rect 3590 3403 3596 3404
rect 110 3391 116 3392
rect 110 3387 111 3391
rect 115 3387 116 3391
rect 1830 3391 1836 3392
rect 110 3386 116 3387
rect 142 3388 148 3389
rect 112 3367 114 3386
rect 142 3384 143 3388
rect 147 3384 148 3388
rect 142 3383 148 3384
rect 286 3388 292 3389
rect 286 3384 287 3388
rect 291 3384 292 3388
rect 286 3383 292 3384
rect 446 3388 452 3389
rect 446 3384 447 3388
rect 451 3384 452 3388
rect 446 3383 452 3384
rect 614 3388 620 3389
rect 614 3384 615 3388
rect 619 3384 620 3388
rect 614 3383 620 3384
rect 782 3388 788 3389
rect 782 3384 783 3388
rect 787 3384 788 3388
rect 782 3383 788 3384
rect 950 3388 956 3389
rect 950 3384 951 3388
rect 955 3384 956 3388
rect 950 3383 956 3384
rect 1110 3388 1116 3389
rect 1110 3384 1111 3388
rect 1115 3384 1116 3388
rect 1110 3383 1116 3384
rect 1262 3388 1268 3389
rect 1262 3384 1263 3388
rect 1267 3384 1268 3388
rect 1262 3383 1268 3384
rect 1406 3388 1412 3389
rect 1406 3384 1407 3388
rect 1411 3384 1412 3388
rect 1406 3383 1412 3384
rect 1550 3388 1556 3389
rect 1550 3384 1551 3388
rect 1555 3384 1556 3388
rect 1550 3383 1556 3384
rect 1702 3388 1708 3389
rect 1702 3384 1703 3388
rect 1707 3384 1708 3388
rect 1830 3387 1831 3391
rect 1835 3387 1836 3391
rect 1830 3386 1836 3387
rect 1870 3391 1876 3392
rect 1870 3387 1871 3391
rect 1875 3387 1876 3391
rect 3590 3391 3596 3392
rect 1870 3386 1876 3387
rect 2102 3388 2108 3389
rect 1702 3383 1708 3384
rect 144 3367 146 3383
rect 288 3367 290 3383
rect 448 3367 450 3383
rect 616 3367 618 3383
rect 784 3367 786 3383
rect 952 3367 954 3383
rect 1112 3367 1114 3383
rect 1264 3367 1266 3383
rect 1408 3367 1410 3383
rect 1552 3367 1554 3383
rect 1704 3367 1706 3383
rect 1832 3367 1834 3386
rect 111 3366 115 3367
rect 111 3361 115 3362
rect 143 3366 147 3367
rect 143 3361 147 3362
rect 207 3366 211 3367
rect 207 3361 211 3362
rect 287 3366 291 3367
rect 287 3361 291 3362
rect 335 3366 339 3367
rect 335 3361 339 3362
rect 447 3366 451 3367
rect 447 3361 451 3362
rect 471 3366 475 3367
rect 471 3361 475 3362
rect 615 3366 619 3367
rect 615 3361 619 3362
rect 623 3366 627 3367
rect 623 3361 627 3362
rect 783 3366 787 3367
rect 783 3361 787 3362
rect 943 3366 947 3367
rect 943 3361 947 3362
rect 951 3366 955 3367
rect 951 3361 955 3362
rect 1103 3366 1107 3367
rect 1103 3361 1107 3362
rect 1111 3366 1115 3367
rect 1111 3361 1115 3362
rect 1263 3366 1267 3367
rect 1263 3361 1267 3362
rect 1407 3366 1411 3367
rect 1407 3361 1411 3362
rect 1423 3366 1427 3367
rect 1423 3361 1427 3362
rect 1551 3366 1555 3367
rect 1551 3361 1555 3362
rect 1583 3366 1587 3367
rect 1583 3361 1587 3362
rect 1703 3366 1707 3367
rect 1703 3361 1707 3362
rect 1743 3366 1747 3367
rect 1743 3361 1747 3362
rect 1831 3366 1835 3367
rect 1872 3363 1874 3386
rect 2102 3384 2103 3388
rect 2107 3384 2108 3388
rect 2102 3383 2108 3384
rect 2190 3388 2196 3389
rect 2190 3384 2191 3388
rect 2195 3384 2196 3388
rect 2190 3383 2196 3384
rect 2294 3388 2300 3389
rect 2294 3384 2295 3388
rect 2299 3384 2300 3388
rect 2294 3383 2300 3384
rect 2406 3388 2412 3389
rect 2406 3384 2407 3388
rect 2411 3384 2412 3388
rect 2406 3383 2412 3384
rect 2534 3388 2540 3389
rect 2534 3384 2535 3388
rect 2539 3384 2540 3388
rect 2534 3383 2540 3384
rect 2670 3388 2676 3389
rect 2670 3384 2671 3388
rect 2675 3384 2676 3388
rect 2670 3383 2676 3384
rect 2806 3388 2812 3389
rect 2806 3384 2807 3388
rect 2811 3384 2812 3388
rect 2806 3383 2812 3384
rect 2950 3388 2956 3389
rect 2950 3384 2951 3388
rect 2955 3384 2956 3388
rect 2950 3383 2956 3384
rect 3102 3388 3108 3389
rect 3102 3384 3103 3388
rect 3107 3384 3108 3388
rect 3102 3383 3108 3384
rect 3254 3388 3260 3389
rect 3254 3384 3255 3388
rect 3259 3384 3260 3388
rect 3254 3383 3260 3384
rect 3414 3388 3420 3389
rect 3414 3384 3415 3388
rect 3419 3384 3420 3388
rect 3590 3387 3591 3391
rect 3595 3387 3596 3391
rect 3590 3386 3596 3387
rect 3414 3383 3420 3384
rect 2104 3363 2106 3383
rect 2192 3363 2194 3383
rect 2296 3363 2298 3383
rect 2408 3363 2410 3383
rect 2536 3363 2538 3383
rect 2672 3363 2674 3383
rect 2808 3363 2810 3383
rect 2952 3363 2954 3383
rect 3104 3363 3106 3383
rect 3256 3363 3258 3383
rect 3416 3363 3418 3383
rect 3592 3363 3594 3386
rect 1831 3361 1835 3362
rect 1871 3362 1875 3363
rect 112 3342 114 3361
rect 208 3345 210 3361
rect 336 3345 338 3361
rect 472 3345 474 3361
rect 624 3345 626 3361
rect 784 3345 786 3361
rect 944 3345 946 3361
rect 1104 3345 1106 3361
rect 1264 3345 1266 3361
rect 1424 3345 1426 3361
rect 1584 3345 1586 3361
rect 1744 3345 1746 3361
rect 206 3344 212 3345
rect 110 3341 116 3342
rect 110 3337 111 3341
rect 115 3337 116 3341
rect 206 3340 207 3344
rect 211 3340 212 3344
rect 206 3339 212 3340
rect 334 3344 340 3345
rect 334 3340 335 3344
rect 339 3340 340 3344
rect 334 3339 340 3340
rect 470 3344 476 3345
rect 470 3340 471 3344
rect 475 3340 476 3344
rect 470 3339 476 3340
rect 622 3344 628 3345
rect 622 3340 623 3344
rect 627 3340 628 3344
rect 622 3339 628 3340
rect 782 3344 788 3345
rect 782 3340 783 3344
rect 787 3340 788 3344
rect 782 3339 788 3340
rect 942 3344 948 3345
rect 942 3340 943 3344
rect 947 3340 948 3344
rect 942 3339 948 3340
rect 1102 3344 1108 3345
rect 1102 3340 1103 3344
rect 1107 3340 1108 3344
rect 1102 3339 1108 3340
rect 1262 3344 1268 3345
rect 1262 3340 1263 3344
rect 1267 3340 1268 3344
rect 1262 3339 1268 3340
rect 1422 3344 1428 3345
rect 1422 3340 1423 3344
rect 1427 3340 1428 3344
rect 1422 3339 1428 3340
rect 1582 3344 1588 3345
rect 1582 3340 1583 3344
rect 1587 3340 1588 3344
rect 1582 3339 1588 3340
rect 1742 3344 1748 3345
rect 1742 3340 1743 3344
rect 1747 3340 1748 3344
rect 1832 3342 1834 3361
rect 1871 3357 1875 3358
rect 2103 3362 2107 3363
rect 2103 3357 2107 3358
rect 2127 3362 2131 3363
rect 2127 3357 2131 3358
rect 2191 3362 2195 3363
rect 2191 3357 2195 3358
rect 2223 3362 2227 3363
rect 2223 3357 2227 3358
rect 2295 3362 2299 3363
rect 2295 3357 2299 3358
rect 2335 3362 2339 3363
rect 2335 3357 2339 3358
rect 2407 3362 2411 3363
rect 2407 3357 2411 3358
rect 2455 3362 2459 3363
rect 2455 3357 2459 3358
rect 2535 3362 2539 3363
rect 2535 3357 2539 3358
rect 2583 3362 2587 3363
rect 2583 3357 2587 3358
rect 2671 3362 2675 3363
rect 2671 3357 2675 3358
rect 2719 3362 2723 3363
rect 2719 3357 2723 3358
rect 2807 3362 2811 3363
rect 2807 3357 2811 3358
rect 2863 3362 2867 3363
rect 2863 3357 2867 3358
rect 2951 3362 2955 3363
rect 2951 3357 2955 3358
rect 3007 3362 3011 3363
rect 3007 3357 3011 3358
rect 3103 3362 3107 3363
rect 3103 3357 3107 3358
rect 3159 3362 3163 3363
rect 3159 3357 3163 3358
rect 3255 3362 3259 3363
rect 3255 3357 3259 3358
rect 3311 3362 3315 3363
rect 3311 3357 3315 3358
rect 3415 3362 3419 3363
rect 3415 3357 3419 3358
rect 3471 3362 3475 3363
rect 3471 3357 3475 3358
rect 3591 3362 3595 3363
rect 3591 3357 3595 3358
rect 1742 3339 1748 3340
rect 1830 3341 1836 3342
rect 110 3336 116 3337
rect 1830 3337 1831 3341
rect 1835 3337 1836 3341
rect 1872 3338 1874 3357
rect 2128 3341 2130 3357
rect 2224 3341 2226 3357
rect 2336 3341 2338 3357
rect 2456 3341 2458 3357
rect 2584 3341 2586 3357
rect 2720 3341 2722 3357
rect 2864 3341 2866 3357
rect 3008 3341 3010 3357
rect 3160 3341 3162 3357
rect 3312 3341 3314 3357
rect 3472 3341 3474 3357
rect 2126 3340 2132 3341
rect 1830 3336 1836 3337
rect 1870 3337 1876 3338
rect 1870 3333 1871 3337
rect 1875 3333 1876 3337
rect 2126 3336 2127 3340
rect 2131 3336 2132 3340
rect 2126 3335 2132 3336
rect 2222 3340 2228 3341
rect 2222 3336 2223 3340
rect 2227 3336 2228 3340
rect 2222 3335 2228 3336
rect 2334 3340 2340 3341
rect 2334 3336 2335 3340
rect 2339 3336 2340 3340
rect 2334 3335 2340 3336
rect 2454 3340 2460 3341
rect 2454 3336 2455 3340
rect 2459 3336 2460 3340
rect 2454 3335 2460 3336
rect 2582 3340 2588 3341
rect 2582 3336 2583 3340
rect 2587 3336 2588 3340
rect 2582 3335 2588 3336
rect 2718 3340 2724 3341
rect 2718 3336 2719 3340
rect 2723 3336 2724 3340
rect 2718 3335 2724 3336
rect 2862 3340 2868 3341
rect 2862 3336 2863 3340
rect 2867 3336 2868 3340
rect 2862 3335 2868 3336
rect 3006 3340 3012 3341
rect 3006 3336 3007 3340
rect 3011 3336 3012 3340
rect 3006 3335 3012 3336
rect 3158 3340 3164 3341
rect 3158 3336 3159 3340
rect 3163 3336 3164 3340
rect 3158 3335 3164 3336
rect 3310 3340 3316 3341
rect 3310 3336 3311 3340
rect 3315 3336 3316 3340
rect 3310 3335 3316 3336
rect 3470 3340 3476 3341
rect 3470 3336 3471 3340
rect 3475 3336 3476 3340
rect 3592 3338 3594 3357
rect 3470 3335 3476 3336
rect 3590 3337 3596 3338
rect 1870 3332 1876 3333
rect 3590 3333 3591 3337
rect 3595 3333 3596 3337
rect 3590 3332 3596 3333
rect 110 3324 116 3325
rect 110 3320 111 3324
rect 115 3320 116 3324
rect 110 3319 116 3320
rect 1830 3324 1836 3325
rect 1830 3320 1831 3324
rect 1835 3320 1836 3324
rect 1830 3319 1836 3320
rect 1870 3320 1876 3321
rect 112 3287 114 3319
rect 214 3306 220 3307
rect 214 3302 215 3306
rect 219 3302 220 3306
rect 214 3301 220 3302
rect 342 3306 348 3307
rect 342 3302 343 3306
rect 347 3302 348 3306
rect 342 3301 348 3302
rect 478 3306 484 3307
rect 478 3302 479 3306
rect 483 3302 484 3306
rect 478 3301 484 3302
rect 630 3306 636 3307
rect 630 3302 631 3306
rect 635 3302 636 3306
rect 630 3301 636 3302
rect 790 3306 796 3307
rect 790 3302 791 3306
rect 795 3302 796 3306
rect 790 3301 796 3302
rect 950 3306 956 3307
rect 950 3302 951 3306
rect 955 3302 956 3306
rect 950 3301 956 3302
rect 1110 3306 1116 3307
rect 1110 3302 1111 3306
rect 1115 3302 1116 3306
rect 1110 3301 1116 3302
rect 1270 3306 1276 3307
rect 1270 3302 1271 3306
rect 1275 3302 1276 3306
rect 1270 3301 1276 3302
rect 1430 3306 1436 3307
rect 1430 3302 1431 3306
rect 1435 3302 1436 3306
rect 1430 3301 1436 3302
rect 1590 3306 1596 3307
rect 1590 3302 1591 3306
rect 1595 3302 1596 3306
rect 1590 3301 1596 3302
rect 1750 3306 1756 3307
rect 1750 3302 1751 3306
rect 1755 3302 1756 3306
rect 1750 3301 1756 3302
rect 216 3287 218 3301
rect 344 3287 346 3301
rect 480 3287 482 3301
rect 632 3287 634 3301
rect 792 3287 794 3301
rect 952 3287 954 3301
rect 1112 3287 1114 3301
rect 1272 3287 1274 3301
rect 1432 3287 1434 3301
rect 1592 3287 1594 3301
rect 1752 3287 1754 3301
rect 1832 3287 1834 3319
rect 1870 3316 1871 3320
rect 1875 3316 1876 3320
rect 1870 3315 1876 3316
rect 3590 3320 3596 3321
rect 3590 3316 3591 3320
rect 3595 3316 3596 3320
rect 3590 3315 3596 3316
rect 111 3286 115 3287
rect 111 3281 115 3282
rect 215 3286 219 3287
rect 215 3281 219 3282
rect 343 3286 347 3287
rect 343 3281 347 3282
rect 351 3286 355 3287
rect 351 3281 355 3282
rect 455 3286 459 3287
rect 455 3281 459 3282
rect 479 3286 483 3287
rect 479 3281 483 3282
rect 575 3286 579 3287
rect 575 3281 579 3282
rect 631 3286 635 3287
rect 631 3281 635 3282
rect 703 3286 707 3287
rect 703 3281 707 3282
rect 791 3286 795 3287
rect 791 3281 795 3282
rect 839 3286 843 3287
rect 839 3281 843 3282
rect 951 3286 955 3287
rect 951 3281 955 3282
rect 983 3286 987 3287
rect 983 3281 987 3282
rect 1111 3286 1115 3287
rect 1111 3281 1115 3282
rect 1119 3286 1123 3287
rect 1119 3281 1123 3282
rect 1255 3286 1259 3287
rect 1255 3281 1259 3282
rect 1271 3286 1275 3287
rect 1271 3281 1275 3282
rect 1383 3286 1387 3287
rect 1383 3281 1387 3282
rect 1431 3286 1435 3287
rect 1431 3281 1435 3282
rect 1511 3286 1515 3287
rect 1511 3281 1515 3282
rect 1591 3286 1595 3287
rect 1591 3281 1595 3282
rect 1639 3286 1643 3287
rect 1639 3281 1643 3282
rect 1751 3286 1755 3287
rect 1751 3281 1755 3282
rect 1831 3286 1835 3287
rect 1831 3281 1835 3282
rect 112 3253 114 3281
rect 352 3271 354 3281
rect 456 3271 458 3281
rect 576 3271 578 3281
rect 704 3271 706 3281
rect 840 3271 842 3281
rect 984 3271 986 3281
rect 1120 3271 1122 3281
rect 1256 3271 1258 3281
rect 1384 3271 1386 3281
rect 1512 3271 1514 3281
rect 1640 3271 1642 3281
rect 1752 3271 1754 3281
rect 350 3270 356 3271
rect 350 3266 351 3270
rect 355 3266 356 3270
rect 350 3265 356 3266
rect 454 3270 460 3271
rect 454 3266 455 3270
rect 459 3266 460 3270
rect 454 3265 460 3266
rect 574 3270 580 3271
rect 574 3266 575 3270
rect 579 3266 580 3270
rect 574 3265 580 3266
rect 702 3270 708 3271
rect 702 3266 703 3270
rect 707 3266 708 3270
rect 702 3265 708 3266
rect 838 3270 844 3271
rect 838 3266 839 3270
rect 843 3266 844 3270
rect 838 3265 844 3266
rect 982 3270 988 3271
rect 982 3266 983 3270
rect 987 3266 988 3270
rect 982 3265 988 3266
rect 1118 3270 1124 3271
rect 1118 3266 1119 3270
rect 1123 3266 1124 3270
rect 1118 3265 1124 3266
rect 1254 3270 1260 3271
rect 1254 3266 1255 3270
rect 1259 3266 1260 3270
rect 1254 3265 1260 3266
rect 1382 3270 1388 3271
rect 1382 3266 1383 3270
rect 1387 3266 1388 3270
rect 1382 3265 1388 3266
rect 1510 3270 1516 3271
rect 1510 3266 1511 3270
rect 1515 3266 1516 3270
rect 1510 3265 1516 3266
rect 1638 3270 1644 3271
rect 1638 3266 1639 3270
rect 1643 3266 1644 3270
rect 1638 3265 1644 3266
rect 1750 3270 1756 3271
rect 1750 3266 1751 3270
rect 1755 3266 1756 3270
rect 1750 3265 1756 3266
rect 1832 3253 1834 3281
rect 1872 3275 1874 3315
rect 2134 3302 2140 3303
rect 2134 3298 2135 3302
rect 2139 3298 2140 3302
rect 2134 3297 2140 3298
rect 2230 3302 2236 3303
rect 2230 3298 2231 3302
rect 2235 3298 2236 3302
rect 2230 3297 2236 3298
rect 2342 3302 2348 3303
rect 2342 3298 2343 3302
rect 2347 3298 2348 3302
rect 2342 3297 2348 3298
rect 2462 3302 2468 3303
rect 2462 3298 2463 3302
rect 2467 3298 2468 3302
rect 2462 3297 2468 3298
rect 2590 3302 2596 3303
rect 2590 3298 2591 3302
rect 2595 3298 2596 3302
rect 2590 3297 2596 3298
rect 2726 3302 2732 3303
rect 2726 3298 2727 3302
rect 2731 3298 2732 3302
rect 2726 3297 2732 3298
rect 2870 3302 2876 3303
rect 2870 3298 2871 3302
rect 2875 3298 2876 3302
rect 2870 3297 2876 3298
rect 3014 3302 3020 3303
rect 3014 3298 3015 3302
rect 3019 3298 3020 3302
rect 3014 3297 3020 3298
rect 3166 3302 3172 3303
rect 3166 3298 3167 3302
rect 3171 3298 3172 3302
rect 3166 3297 3172 3298
rect 3318 3302 3324 3303
rect 3318 3298 3319 3302
rect 3323 3298 3324 3302
rect 3318 3297 3324 3298
rect 3478 3302 3484 3303
rect 3478 3298 3479 3302
rect 3483 3298 3484 3302
rect 3478 3297 3484 3298
rect 2136 3275 2138 3297
rect 2232 3275 2234 3297
rect 2344 3275 2346 3297
rect 2464 3275 2466 3297
rect 2592 3275 2594 3297
rect 2728 3275 2730 3297
rect 2872 3275 2874 3297
rect 3016 3275 3018 3297
rect 3168 3275 3170 3297
rect 3320 3275 3322 3297
rect 3480 3275 3482 3297
rect 3592 3275 3594 3315
rect 1871 3274 1875 3275
rect 1871 3269 1875 3270
rect 2135 3274 2139 3275
rect 2135 3269 2139 3270
rect 2231 3274 2235 3275
rect 2231 3269 2235 3270
rect 2279 3274 2283 3275
rect 2279 3269 2283 3270
rect 2343 3274 2347 3275
rect 2343 3269 2347 3270
rect 2415 3274 2419 3275
rect 2415 3269 2419 3270
rect 2463 3274 2467 3275
rect 2463 3269 2467 3270
rect 2551 3274 2555 3275
rect 2551 3269 2555 3270
rect 2591 3274 2595 3275
rect 2591 3269 2595 3270
rect 2687 3274 2691 3275
rect 2687 3269 2691 3270
rect 2727 3274 2731 3275
rect 2727 3269 2731 3270
rect 2823 3274 2827 3275
rect 2823 3269 2827 3270
rect 2871 3274 2875 3275
rect 2871 3269 2875 3270
rect 2959 3274 2963 3275
rect 2959 3269 2963 3270
rect 3015 3274 3019 3275
rect 3015 3269 3019 3270
rect 3095 3274 3099 3275
rect 3095 3269 3099 3270
rect 3167 3274 3171 3275
rect 3167 3269 3171 3270
rect 3231 3274 3235 3275
rect 3231 3269 3235 3270
rect 3319 3274 3323 3275
rect 3319 3269 3323 3270
rect 3375 3274 3379 3275
rect 3375 3269 3379 3270
rect 3479 3274 3483 3275
rect 3479 3269 3483 3270
rect 3511 3274 3515 3275
rect 3511 3269 3515 3270
rect 3591 3274 3595 3275
rect 3591 3269 3595 3270
rect 110 3252 116 3253
rect 110 3248 111 3252
rect 115 3248 116 3252
rect 110 3247 116 3248
rect 1830 3252 1836 3253
rect 1830 3248 1831 3252
rect 1835 3248 1836 3252
rect 1830 3247 1836 3248
rect 1872 3241 1874 3269
rect 2136 3259 2138 3269
rect 2280 3259 2282 3269
rect 2416 3259 2418 3269
rect 2552 3259 2554 3269
rect 2688 3259 2690 3269
rect 2824 3259 2826 3269
rect 2960 3259 2962 3269
rect 3096 3259 3098 3269
rect 3232 3259 3234 3269
rect 3376 3259 3378 3269
rect 3512 3259 3514 3269
rect 2134 3258 2140 3259
rect 2134 3254 2135 3258
rect 2139 3254 2140 3258
rect 2134 3253 2140 3254
rect 2278 3258 2284 3259
rect 2278 3254 2279 3258
rect 2283 3254 2284 3258
rect 2278 3253 2284 3254
rect 2414 3258 2420 3259
rect 2414 3254 2415 3258
rect 2419 3254 2420 3258
rect 2414 3253 2420 3254
rect 2550 3258 2556 3259
rect 2550 3254 2551 3258
rect 2555 3254 2556 3258
rect 2550 3253 2556 3254
rect 2686 3258 2692 3259
rect 2686 3254 2687 3258
rect 2691 3254 2692 3258
rect 2686 3253 2692 3254
rect 2822 3258 2828 3259
rect 2822 3254 2823 3258
rect 2827 3254 2828 3258
rect 2822 3253 2828 3254
rect 2958 3258 2964 3259
rect 2958 3254 2959 3258
rect 2963 3254 2964 3258
rect 2958 3253 2964 3254
rect 3094 3258 3100 3259
rect 3094 3254 3095 3258
rect 3099 3254 3100 3258
rect 3094 3253 3100 3254
rect 3230 3258 3236 3259
rect 3230 3254 3231 3258
rect 3235 3254 3236 3258
rect 3230 3253 3236 3254
rect 3374 3258 3380 3259
rect 3374 3254 3375 3258
rect 3379 3254 3380 3258
rect 3374 3253 3380 3254
rect 3510 3258 3516 3259
rect 3510 3254 3511 3258
rect 3515 3254 3516 3258
rect 3510 3253 3516 3254
rect 3592 3241 3594 3269
rect 1870 3240 1876 3241
rect 1870 3236 1871 3240
rect 1875 3236 1876 3240
rect 110 3235 116 3236
rect 110 3231 111 3235
rect 115 3231 116 3235
rect 1830 3235 1836 3236
rect 1870 3235 1876 3236
rect 3590 3240 3596 3241
rect 3590 3236 3591 3240
rect 3595 3236 3596 3240
rect 3590 3235 3596 3236
rect 110 3230 116 3231
rect 342 3232 348 3233
rect 112 3211 114 3230
rect 342 3228 343 3232
rect 347 3228 348 3232
rect 342 3227 348 3228
rect 446 3232 452 3233
rect 446 3228 447 3232
rect 451 3228 452 3232
rect 446 3227 452 3228
rect 566 3232 572 3233
rect 566 3228 567 3232
rect 571 3228 572 3232
rect 566 3227 572 3228
rect 694 3232 700 3233
rect 694 3228 695 3232
rect 699 3228 700 3232
rect 694 3227 700 3228
rect 830 3232 836 3233
rect 830 3228 831 3232
rect 835 3228 836 3232
rect 830 3227 836 3228
rect 974 3232 980 3233
rect 974 3228 975 3232
rect 979 3228 980 3232
rect 974 3227 980 3228
rect 1110 3232 1116 3233
rect 1110 3228 1111 3232
rect 1115 3228 1116 3232
rect 1110 3227 1116 3228
rect 1246 3232 1252 3233
rect 1246 3228 1247 3232
rect 1251 3228 1252 3232
rect 1246 3227 1252 3228
rect 1374 3232 1380 3233
rect 1374 3228 1375 3232
rect 1379 3228 1380 3232
rect 1374 3227 1380 3228
rect 1502 3232 1508 3233
rect 1502 3228 1503 3232
rect 1507 3228 1508 3232
rect 1502 3227 1508 3228
rect 1630 3232 1636 3233
rect 1630 3228 1631 3232
rect 1635 3228 1636 3232
rect 1630 3227 1636 3228
rect 1742 3232 1748 3233
rect 1742 3228 1743 3232
rect 1747 3228 1748 3232
rect 1830 3231 1831 3235
rect 1835 3231 1836 3235
rect 1830 3230 1836 3231
rect 1742 3227 1748 3228
rect 344 3211 346 3227
rect 448 3211 450 3227
rect 568 3211 570 3227
rect 696 3211 698 3227
rect 832 3211 834 3227
rect 976 3211 978 3227
rect 1112 3211 1114 3227
rect 1248 3211 1250 3227
rect 1376 3211 1378 3227
rect 1504 3211 1506 3227
rect 1632 3211 1634 3227
rect 1744 3211 1746 3227
rect 1832 3211 1834 3230
rect 1870 3223 1876 3224
rect 1870 3219 1871 3223
rect 1875 3219 1876 3223
rect 3590 3223 3596 3224
rect 1870 3218 1876 3219
rect 2126 3220 2132 3221
rect 111 3210 115 3211
rect 111 3205 115 3206
rect 343 3210 347 3211
rect 343 3205 347 3206
rect 447 3210 451 3211
rect 447 3205 451 3206
rect 487 3210 491 3211
rect 487 3205 491 3206
rect 567 3210 571 3211
rect 567 3205 571 3206
rect 575 3210 579 3211
rect 575 3205 579 3206
rect 663 3210 667 3211
rect 663 3205 667 3206
rect 695 3210 699 3211
rect 695 3205 699 3206
rect 767 3210 771 3211
rect 767 3205 771 3206
rect 831 3210 835 3211
rect 831 3205 835 3206
rect 887 3210 891 3211
rect 887 3205 891 3206
rect 975 3210 979 3211
rect 975 3205 979 3206
rect 1023 3210 1027 3211
rect 1023 3205 1027 3206
rect 1111 3210 1115 3211
rect 1111 3205 1115 3206
rect 1191 3210 1195 3211
rect 1191 3205 1195 3206
rect 1247 3210 1251 3211
rect 1247 3205 1251 3206
rect 1375 3210 1379 3211
rect 1375 3205 1379 3206
rect 1503 3210 1507 3211
rect 1503 3205 1507 3206
rect 1567 3210 1571 3211
rect 1567 3205 1571 3206
rect 1631 3210 1635 3211
rect 1631 3205 1635 3206
rect 1743 3210 1747 3211
rect 1743 3205 1747 3206
rect 1831 3210 1835 3211
rect 1831 3205 1835 3206
rect 112 3186 114 3205
rect 488 3189 490 3205
rect 576 3189 578 3205
rect 664 3189 666 3205
rect 768 3189 770 3205
rect 888 3189 890 3205
rect 1024 3189 1026 3205
rect 1192 3189 1194 3205
rect 1376 3189 1378 3205
rect 1568 3189 1570 3205
rect 1744 3189 1746 3205
rect 486 3188 492 3189
rect 110 3185 116 3186
rect 110 3181 111 3185
rect 115 3181 116 3185
rect 486 3184 487 3188
rect 491 3184 492 3188
rect 486 3183 492 3184
rect 574 3188 580 3189
rect 574 3184 575 3188
rect 579 3184 580 3188
rect 574 3183 580 3184
rect 662 3188 668 3189
rect 662 3184 663 3188
rect 667 3184 668 3188
rect 662 3183 668 3184
rect 766 3188 772 3189
rect 766 3184 767 3188
rect 771 3184 772 3188
rect 766 3183 772 3184
rect 886 3188 892 3189
rect 886 3184 887 3188
rect 891 3184 892 3188
rect 886 3183 892 3184
rect 1022 3188 1028 3189
rect 1022 3184 1023 3188
rect 1027 3184 1028 3188
rect 1022 3183 1028 3184
rect 1190 3188 1196 3189
rect 1190 3184 1191 3188
rect 1195 3184 1196 3188
rect 1190 3183 1196 3184
rect 1374 3188 1380 3189
rect 1374 3184 1375 3188
rect 1379 3184 1380 3188
rect 1374 3183 1380 3184
rect 1566 3188 1572 3189
rect 1566 3184 1567 3188
rect 1571 3184 1572 3188
rect 1566 3183 1572 3184
rect 1742 3188 1748 3189
rect 1742 3184 1743 3188
rect 1747 3184 1748 3188
rect 1832 3186 1834 3205
rect 1872 3195 1874 3218
rect 2126 3216 2127 3220
rect 2131 3216 2132 3220
rect 2126 3215 2132 3216
rect 2270 3220 2276 3221
rect 2270 3216 2271 3220
rect 2275 3216 2276 3220
rect 2270 3215 2276 3216
rect 2406 3220 2412 3221
rect 2406 3216 2407 3220
rect 2411 3216 2412 3220
rect 2406 3215 2412 3216
rect 2542 3220 2548 3221
rect 2542 3216 2543 3220
rect 2547 3216 2548 3220
rect 2542 3215 2548 3216
rect 2678 3220 2684 3221
rect 2678 3216 2679 3220
rect 2683 3216 2684 3220
rect 2678 3215 2684 3216
rect 2814 3220 2820 3221
rect 2814 3216 2815 3220
rect 2819 3216 2820 3220
rect 2814 3215 2820 3216
rect 2950 3220 2956 3221
rect 2950 3216 2951 3220
rect 2955 3216 2956 3220
rect 2950 3215 2956 3216
rect 3086 3220 3092 3221
rect 3086 3216 3087 3220
rect 3091 3216 3092 3220
rect 3086 3215 3092 3216
rect 3222 3220 3228 3221
rect 3222 3216 3223 3220
rect 3227 3216 3228 3220
rect 3222 3215 3228 3216
rect 3366 3220 3372 3221
rect 3366 3216 3367 3220
rect 3371 3216 3372 3220
rect 3366 3215 3372 3216
rect 3502 3220 3508 3221
rect 3502 3216 3503 3220
rect 3507 3216 3508 3220
rect 3590 3219 3591 3223
rect 3595 3219 3596 3223
rect 3590 3218 3596 3219
rect 3502 3215 3508 3216
rect 2128 3195 2130 3215
rect 2272 3195 2274 3215
rect 2408 3195 2410 3215
rect 2544 3195 2546 3215
rect 2680 3195 2682 3215
rect 2816 3195 2818 3215
rect 2952 3195 2954 3215
rect 3088 3195 3090 3215
rect 3224 3195 3226 3215
rect 3368 3195 3370 3215
rect 3504 3195 3506 3215
rect 3592 3195 3594 3218
rect 1871 3194 1875 3195
rect 1871 3189 1875 3190
rect 1895 3194 1899 3195
rect 1895 3189 1899 3190
rect 1991 3194 1995 3195
rect 1991 3189 1995 3190
rect 2119 3194 2123 3195
rect 2119 3189 2123 3190
rect 2127 3194 2131 3195
rect 2127 3189 2131 3190
rect 2247 3194 2251 3195
rect 2247 3189 2251 3190
rect 2271 3194 2275 3195
rect 2271 3189 2275 3190
rect 2383 3194 2387 3195
rect 2383 3189 2387 3190
rect 2407 3194 2411 3195
rect 2407 3189 2411 3190
rect 2511 3194 2515 3195
rect 2511 3189 2515 3190
rect 2543 3194 2547 3195
rect 2543 3189 2547 3190
rect 2639 3194 2643 3195
rect 2639 3189 2643 3190
rect 2679 3194 2683 3195
rect 2679 3189 2683 3190
rect 2767 3194 2771 3195
rect 2767 3189 2771 3190
rect 2815 3194 2819 3195
rect 2815 3189 2819 3190
rect 2895 3194 2899 3195
rect 2895 3189 2899 3190
rect 2951 3194 2955 3195
rect 2951 3189 2955 3190
rect 3031 3194 3035 3195
rect 3031 3189 3035 3190
rect 3087 3194 3091 3195
rect 3087 3189 3091 3190
rect 3175 3194 3179 3195
rect 3175 3189 3179 3190
rect 3223 3194 3227 3195
rect 3223 3189 3227 3190
rect 3327 3194 3331 3195
rect 3327 3189 3331 3190
rect 3367 3194 3371 3195
rect 3367 3189 3371 3190
rect 3487 3194 3491 3195
rect 3487 3189 3491 3190
rect 3503 3194 3507 3195
rect 3503 3189 3507 3190
rect 3591 3194 3595 3195
rect 3591 3189 3595 3190
rect 1742 3183 1748 3184
rect 1830 3185 1836 3186
rect 110 3180 116 3181
rect 1830 3181 1831 3185
rect 1835 3181 1836 3185
rect 1830 3180 1836 3181
rect 1872 3170 1874 3189
rect 1896 3173 1898 3189
rect 1992 3173 1994 3189
rect 2120 3173 2122 3189
rect 2248 3173 2250 3189
rect 2384 3173 2386 3189
rect 2512 3173 2514 3189
rect 2640 3173 2642 3189
rect 2768 3173 2770 3189
rect 2896 3173 2898 3189
rect 3032 3173 3034 3189
rect 3176 3173 3178 3189
rect 3328 3173 3330 3189
rect 3488 3173 3490 3189
rect 1894 3172 1900 3173
rect 1870 3169 1876 3170
rect 110 3168 116 3169
rect 110 3164 111 3168
rect 115 3164 116 3168
rect 110 3163 116 3164
rect 1830 3168 1836 3169
rect 1830 3164 1831 3168
rect 1835 3164 1836 3168
rect 1870 3165 1871 3169
rect 1875 3165 1876 3169
rect 1894 3168 1895 3172
rect 1899 3168 1900 3172
rect 1894 3167 1900 3168
rect 1990 3172 1996 3173
rect 1990 3168 1991 3172
rect 1995 3168 1996 3172
rect 1990 3167 1996 3168
rect 2118 3172 2124 3173
rect 2118 3168 2119 3172
rect 2123 3168 2124 3172
rect 2118 3167 2124 3168
rect 2246 3172 2252 3173
rect 2246 3168 2247 3172
rect 2251 3168 2252 3172
rect 2246 3167 2252 3168
rect 2382 3172 2388 3173
rect 2382 3168 2383 3172
rect 2387 3168 2388 3172
rect 2382 3167 2388 3168
rect 2510 3172 2516 3173
rect 2510 3168 2511 3172
rect 2515 3168 2516 3172
rect 2510 3167 2516 3168
rect 2638 3172 2644 3173
rect 2638 3168 2639 3172
rect 2643 3168 2644 3172
rect 2638 3167 2644 3168
rect 2766 3172 2772 3173
rect 2766 3168 2767 3172
rect 2771 3168 2772 3172
rect 2766 3167 2772 3168
rect 2894 3172 2900 3173
rect 2894 3168 2895 3172
rect 2899 3168 2900 3172
rect 2894 3167 2900 3168
rect 3030 3172 3036 3173
rect 3030 3168 3031 3172
rect 3035 3168 3036 3172
rect 3030 3167 3036 3168
rect 3174 3172 3180 3173
rect 3174 3168 3175 3172
rect 3179 3168 3180 3172
rect 3174 3167 3180 3168
rect 3326 3172 3332 3173
rect 3326 3168 3327 3172
rect 3331 3168 3332 3172
rect 3326 3167 3332 3168
rect 3486 3172 3492 3173
rect 3486 3168 3487 3172
rect 3491 3168 3492 3172
rect 3592 3170 3594 3189
rect 3486 3167 3492 3168
rect 3590 3169 3596 3170
rect 1870 3164 1876 3165
rect 3590 3165 3591 3169
rect 3595 3165 3596 3169
rect 3590 3164 3596 3165
rect 1830 3163 1836 3164
rect 112 3131 114 3163
rect 494 3150 500 3151
rect 494 3146 495 3150
rect 499 3146 500 3150
rect 494 3145 500 3146
rect 582 3150 588 3151
rect 582 3146 583 3150
rect 587 3146 588 3150
rect 582 3145 588 3146
rect 670 3150 676 3151
rect 670 3146 671 3150
rect 675 3146 676 3150
rect 670 3145 676 3146
rect 774 3150 780 3151
rect 774 3146 775 3150
rect 779 3146 780 3150
rect 774 3145 780 3146
rect 894 3150 900 3151
rect 894 3146 895 3150
rect 899 3146 900 3150
rect 894 3145 900 3146
rect 1030 3150 1036 3151
rect 1030 3146 1031 3150
rect 1035 3146 1036 3150
rect 1030 3145 1036 3146
rect 1198 3150 1204 3151
rect 1198 3146 1199 3150
rect 1203 3146 1204 3150
rect 1198 3145 1204 3146
rect 1382 3150 1388 3151
rect 1382 3146 1383 3150
rect 1387 3146 1388 3150
rect 1382 3145 1388 3146
rect 1574 3150 1580 3151
rect 1574 3146 1575 3150
rect 1579 3146 1580 3150
rect 1574 3145 1580 3146
rect 1750 3150 1756 3151
rect 1750 3146 1751 3150
rect 1755 3146 1756 3150
rect 1750 3145 1756 3146
rect 496 3131 498 3145
rect 584 3131 586 3145
rect 672 3131 674 3145
rect 776 3131 778 3145
rect 896 3131 898 3145
rect 1032 3131 1034 3145
rect 1200 3131 1202 3145
rect 1384 3131 1386 3145
rect 1576 3131 1578 3145
rect 1752 3131 1754 3145
rect 1832 3131 1834 3163
rect 1870 3152 1876 3153
rect 1870 3148 1871 3152
rect 1875 3148 1876 3152
rect 1870 3147 1876 3148
rect 3590 3152 3596 3153
rect 3590 3148 3591 3152
rect 3595 3148 3596 3152
rect 3590 3147 3596 3148
rect 111 3130 115 3131
rect 111 3125 115 3126
rect 495 3130 499 3131
rect 495 3125 499 3126
rect 583 3130 587 3131
rect 583 3125 587 3126
rect 591 3130 595 3131
rect 591 3125 595 3126
rect 671 3130 675 3131
rect 671 3125 675 3126
rect 759 3130 763 3131
rect 759 3125 763 3126
rect 775 3130 779 3131
rect 775 3125 779 3126
rect 847 3130 851 3131
rect 847 3125 851 3126
rect 895 3130 899 3131
rect 895 3125 899 3126
rect 935 3130 939 3131
rect 935 3125 939 3126
rect 1023 3130 1027 3131
rect 1023 3125 1027 3126
rect 1031 3130 1035 3131
rect 1031 3125 1035 3126
rect 1111 3130 1115 3131
rect 1111 3125 1115 3126
rect 1199 3130 1203 3131
rect 1199 3125 1203 3126
rect 1287 3130 1291 3131
rect 1287 3125 1291 3126
rect 1375 3130 1379 3131
rect 1375 3125 1379 3126
rect 1383 3130 1387 3131
rect 1383 3125 1387 3126
rect 1575 3130 1579 3131
rect 1575 3125 1579 3126
rect 1751 3130 1755 3131
rect 1751 3125 1755 3126
rect 1831 3130 1835 3131
rect 1831 3125 1835 3126
rect 112 3097 114 3125
rect 592 3115 594 3125
rect 672 3115 674 3125
rect 760 3115 762 3125
rect 848 3115 850 3125
rect 936 3115 938 3125
rect 1024 3115 1026 3125
rect 1112 3115 1114 3125
rect 1200 3115 1202 3125
rect 1288 3115 1290 3125
rect 1376 3115 1378 3125
rect 590 3114 596 3115
rect 590 3110 591 3114
rect 595 3110 596 3114
rect 590 3109 596 3110
rect 670 3114 676 3115
rect 670 3110 671 3114
rect 675 3110 676 3114
rect 670 3109 676 3110
rect 758 3114 764 3115
rect 758 3110 759 3114
rect 763 3110 764 3114
rect 758 3109 764 3110
rect 846 3114 852 3115
rect 846 3110 847 3114
rect 851 3110 852 3114
rect 846 3109 852 3110
rect 934 3114 940 3115
rect 934 3110 935 3114
rect 939 3110 940 3114
rect 934 3109 940 3110
rect 1022 3114 1028 3115
rect 1022 3110 1023 3114
rect 1027 3110 1028 3114
rect 1022 3109 1028 3110
rect 1110 3114 1116 3115
rect 1110 3110 1111 3114
rect 1115 3110 1116 3114
rect 1110 3109 1116 3110
rect 1198 3114 1204 3115
rect 1198 3110 1199 3114
rect 1203 3110 1204 3114
rect 1198 3109 1204 3110
rect 1286 3114 1292 3115
rect 1286 3110 1287 3114
rect 1291 3110 1292 3114
rect 1286 3109 1292 3110
rect 1374 3114 1380 3115
rect 1374 3110 1375 3114
rect 1379 3110 1380 3114
rect 1374 3109 1380 3110
rect 1832 3097 1834 3125
rect 1872 3103 1874 3147
rect 1902 3134 1908 3135
rect 1902 3130 1903 3134
rect 1907 3130 1908 3134
rect 1902 3129 1908 3130
rect 1998 3134 2004 3135
rect 1998 3130 1999 3134
rect 2003 3130 2004 3134
rect 1998 3129 2004 3130
rect 2126 3134 2132 3135
rect 2126 3130 2127 3134
rect 2131 3130 2132 3134
rect 2126 3129 2132 3130
rect 2254 3134 2260 3135
rect 2254 3130 2255 3134
rect 2259 3130 2260 3134
rect 2254 3129 2260 3130
rect 2390 3134 2396 3135
rect 2390 3130 2391 3134
rect 2395 3130 2396 3134
rect 2390 3129 2396 3130
rect 2518 3134 2524 3135
rect 2518 3130 2519 3134
rect 2523 3130 2524 3134
rect 2518 3129 2524 3130
rect 2646 3134 2652 3135
rect 2646 3130 2647 3134
rect 2651 3130 2652 3134
rect 2646 3129 2652 3130
rect 2774 3134 2780 3135
rect 2774 3130 2775 3134
rect 2779 3130 2780 3134
rect 2774 3129 2780 3130
rect 2902 3134 2908 3135
rect 2902 3130 2903 3134
rect 2907 3130 2908 3134
rect 2902 3129 2908 3130
rect 3038 3134 3044 3135
rect 3038 3130 3039 3134
rect 3043 3130 3044 3134
rect 3038 3129 3044 3130
rect 3182 3134 3188 3135
rect 3182 3130 3183 3134
rect 3187 3130 3188 3134
rect 3182 3129 3188 3130
rect 3334 3134 3340 3135
rect 3334 3130 3335 3134
rect 3339 3130 3340 3134
rect 3334 3129 3340 3130
rect 3494 3134 3500 3135
rect 3494 3130 3495 3134
rect 3499 3130 3500 3134
rect 3494 3129 3500 3130
rect 1904 3103 1906 3129
rect 2000 3103 2002 3129
rect 2128 3103 2130 3129
rect 2256 3103 2258 3129
rect 2392 3103 2394 3129
rect 2520 3103 2522 3129
rect 2648 3103 2650 3129
rect 2776 3103 2778 3129
rect 2904 3103 2906 3129
rect 3040 3103 3042 3129
rect 3184 3103 3186 3129
rect 3336 3103 3338 3129
rect 3496 3103 3498 3129
rect 3592 3103 3594 3147
rect 1871 3102 1875 3103
rect 1871 3097 1875 3098
rect 1903 3102 1907 3103
rect 1903 3097 1907 3098
rect 1999 3102 2003 3103
rect 1999 3097 2003 3098
rect 2015 3102 2019 3103
rect 2015 3097 2019 3098
rect 2127 3102 2131 3103
rect 2127 3097 2131 3098
rect 2191 3102 2195 3103
rect 2191 3097 2195 3098
rect 2255 3102 2259 3103
rect 2255 3097 2259 3098
rect 2391 3102 2395 3103
rect 2391 3097 2395 3098
rect 2407 3102 2411 3103
rect 2407 3097 2411 3098
rect 2519 3102 2523 3103
rect 2519 3097 2523 3098
rect 2647 3102 2651 3103
rect 2647 3097 2651 3098
rect 2655 3102 2659 3103
rect 2655 3097 2659 3098
rect 2775 3102 2779 3103
rect 2775 3097 2779 3098
rect 2903 3102 2907 3103
rect 2903 3097 2907 3098
rect 2935 3102 2939 3103
rect 2935 3097 2939 3098
rect 3039 3102 3043 3103
rect 3039 3097 3043 3098
rect 3183 3102 3187 3103
rect 3183 3097 3187 3098
rect 3231 3102 3235 3103
rect 3231 3097 3235 3098
rect 3335 3102 3339 3103
rect 3335 3097 3339 3098
rect 3495 3102 3499 3103
rect 3495 3097 3499 3098
rect 3511 3102 3515 3103
rect 3511 3097 3515 3098
rect 3591 3102 3595 3103
rect 3591 3097 3595 3098
rect 110 3096 116 3097
rect 110 3092 111 3096
rect 115 3092 116 3096
rect 110 3091 116 3092
rect 1830 3096 1836 3097
rect 1830 3092 1831 3096
rect 1835 3092 1836 3096
rect 1830 3091 1836 3092
rect 110 3079 116 3080
rect 110 3075 111 3079
rect 115 3075 116 3079
rect 1830 3079 1836 3080
rect 110 3074 116 3075
rect 582 3076 588 3077
rect 112 3051 114 3074
rect 582 3072 583 3076
rect 587 3072 588 3076
rect 582 3071 588 3072
rect 662 3076 668 3077
rect 662 3072 663 3076
rect 667 3072 668 3076
rect 662 3071 668 3072
rect 750 3076 756 3077
rect 750 3072 751 3076
rect 755 3072 756 3076
rect 750 3071 756 3072
rect 838 3076 844 3077
rect 838 3072 839 3076
rect 843 3072 844 3076
rect 838 3071 844 3072
rect 926 3076 932 3077
rect 926 3072 927 3076
rect 931 3072 932 3076
rect 926 3071 932 3072
rect 1014 3076 1020 3077
rect 1014 3072 1015 3076
rect 1019 3072 1020 3076
rect 1014 3071 1020 3072
rect 1102 3076 1108 3077
rect 1102 3072 1103 3076
rect 1107 3072 1108 3076
rect 1102 3071 1108 3072
rect 1190 3076 1196 3077
rect 1190 3072 1191 3076
rect 1195 3072 1196 3076
rect 1190 3071 1196 3072
rect 1278 3076 1284 3077
rect 1278 3072 1279 3076
rect 1283 3072 1284 3076
rect 1278 3071 1284 3072
rect 1366 3076 1372 3077
rect 1366 3072 1367 3076
rect 1371 3072 1372 3076
rect 1830 3075 1831 3079
rect 1835 3075 1836 3079
rect 1830 3074 1836 3075
rect 1366 3071 1372 3072
rect 584 3051 586 3071
rect 664 3051 666 3071
rect 752 3051 754 3071
rect 840 3051 842 3071
rect 928 3051 930 3071
rect 1016 3051 1018 3071
rect 1104 3051 1106 3071
rect 1192 3051 1194 3071
rect 1280 3051 1282 3071
rect 1368 3051 1370 3071
rect 1832 3051 1834 3074
rect 1872 3069 1874 3097
rect 1904 3087 1906 3097
rect 2016 3087 2018 3097
rect 2192 3087 2194 3097
rect 2408 3087 2410 3097
rect 2656 3087 2658 3097
rect 2936 3087 2938 3097
rect 3232 3087 3234 3097
rect 3512 3087 3514 3097
rect 1902 3086 1908 3087
rect 1902 3082 1903 3086
rect 1907 3082 1908 3086
rect 1902 3081 1908 3082
rect 2014 3086 2020 3087
rect 2014 3082 2015 3086
rect 2019 3082 2020 3086
rect 2014 3081 2020 3082
rect 2190 3086 2196 3087
rect 2190 3082 2191 3086
rect 2195 3082 2196 3086
rect 2190 3081 2196 3082
rect 2406 3086 2412 3087
rect 2406 3082 2407 3086
rect 2411 3082 2412 3086
rect 2406 3081 2412 3082
rect 2654 3086 2660 3087
rect 2654 3082 2655 3086
rect 2659 3082 2660 3086
rect 2654 3081 2660 3082
rect 2934 3086 2940 3087
rect 2934 3082 2935 3086
rect 2939 3082 2940 3086
rect 2934 3081 2940 3082
rect 3230 3086 3236 3087
rect 3230 3082 3231 3086
rect 3235 3082 3236 3086
rect 3230 3081 3236 3082
rect 3510 3086 3516 3087
rect 3510 3082 3511 3086
rect 3515 3082 3516 3086
rect 3510 3081 3516 3082
rect 3592 3069 3594 3097
rect 1870 3068 1876 3069
rect 1870 3064 1871 3068
rect 1875 3064 1876 3068
rect 1870 3063 1876 3064
rect 3590 3068 3596 3069
rect 3590 3064 3591 3068
rect 3595 3064 3596 3068
rect 3590 3063 3596 3064
rect 1870 3051 1876 3052
rect 111 3050 115 3051
rect 111 3045 115 3046
rect 543 3050 547 3051
rect 543 3045 547 3046
rect 583 3050 587 3051
rect 583 3045 587 3046
rect 623 3050 627 3051
rect 623 3045 627 3046
rect 663 3050 667 3051
rect 663 3045 667 3046
rect 711 3050 715 3051
rect 711 3045 715 3046
rect 751 3050 755 3051
rect 751 3045 755 3046
rect 807 3050 811 3051
rect 807 3045 811 3046
rect 839 3050 843 3051
rect 839 3045 843 3046
rect 903 3050 907 3051
rect 903 3045 907 3046
rect 927 3050 931 3051
rect 927 3045 931 3046
rect 999 3050 1003 3051
rect 999 3045 1003 3046
rect 1015 3050 1019 3051
rect 1015 3045 1019 3046
rect 1087 3050 1091 3051
rect 1087 3045 1091 3046
rect 1103 3050 1107 3051
rect 1103 3045 1107 3046
rect 1183 3050 1187 3051
rect 1183 3045 1187 3046
rect 1191 3050 1195 3051
rect 1191 3045 1195 3046
rect 1279 3050 1283 3051
rect 1279 3045 1283 3046
rect 1367 3050 1371 3051
rect 1367 3045 1371 3046
rect 1375 3050 1379 3051
rect 1375 3045 1379 3046
rect 1471 3050 1475 3051
rect 1471 3045 1475 3046
rect 1831 3050 1835 3051
rect 1870 3047 1871 3051
rect 1875 3047 1876 3051
rect 3590 3051 3596 3052
rect 1870 3046 1876 3047
rect 1894 3048 1900 3049
rect 1831 3045 1835 3046
rect 112 3026 114 3045
rect 544 3029 546 3045
rect 624 3029 626 3045
rect 712 3029 714 3045
rect 808 3029 810 3045
rect 904 3029 906 3045
rect 1000 3029 1002 3045
rect 1088 3029 1090 3045
rect 1184 3029 1186 3045
rect 1280 3029 1282 3045
rect 1376 3029 1378 3045
rect 1472 3029 1474 3045
rect 542 3028 548 3029
rect 110 3025 116 3026
rect 110 3021 111 3025
rect 115 3021 116 3025
rect 542 3024 543 3028
rect 547 3024 548 3028
rect 542 3023 548 3024
rect 622 3028 628 3029
rect 622 3024 623 3028
rect 627 3024 628 3028
rect 622 3023 628 3024
rect 710 3028 716 3029
rect 710 3024 711 3028
rect 715 3024 716 3028
rect 710 3023 716 3024
rect 806 3028 812 3029
rect 806 3024 807 3028
rect 811 3024 812 3028
rect 806 3023 812 3024
rect 902 3028 908 3029
rect 902 3024 903 3028
rect 907 3024 908 3028
rect 902 3023 908 3024
rect 998 3028 1004 3029
rect 998 3024 999 3028
rect 1003 3024 1004 3028
rect 998 3023 1004 3024
rect 1086 3028 1092 3029
rect 1086 3024 1087 3028
rect 1091 3024 1092 3028
rect 1086 3023 1092 3024
rect 1182 3028 1188 3029
rect 1182 3024 1183 3028
rect 1187 3024 1188 3028
rect 1182 3023 1188 3024
rect 1278 3028 1284 3029
rect 1278 3024 1279 3028
rect 1283 3024 1284 3028
rect 1278 3023 1284 3024
rect 1374 3028 1380 3029
rect 1374 3024 1375 3028
rect 1379 3024 1380 3028
rect 1374 3023 1380 3024
rect 1470 3028 1476 3029
rect 1470 3024 1471 3028
rect 1475 3024 1476 3028
rect 1832 3026 1834 3045
rect 1470 3023 1476 3024
rect 1830 3025 1836 3026
rect 110 3020 116 3021
rect 1830 3021 1831 3025
rect 1835 3021 1836 3025
rect 1830 3020 1836 3021
rect 1872 3019 1874 3046
rect 1894 3044 1895 3048
rect 1899 3044 1900 3048
rect 1894 3043 1900 3044
rect 2006 3048 2012 3049
rect 2006 3044 2007 3048
rect 2011 3044 2012 3048
rect 2006 3043 2012 3044
rect 2182 3048 2188 3049
rect 2182 3044 2183 3048
rect 2187 3044 2188 3048
rect 2182 3043 2188 3044
rect 2398 3048 2404 3049
rect 2398 3044 2399 3048
rect 2403 3044 2404 3048
rect 2398 3043 2404 3044
rect 2646 3048 2652 3049
rect 2646 3044 2647 3048
rect 2651 3044 2652 3048
rect 2646 3043 2652 3044
rect 2926 3048 2932 3049
rect 2926 3044 2927 3048
rect 2931 3044 2932 3048
rect 2926 3043 2932 3044
rect 3222 3048 3228 3049
rect 3222 3044 3223 3048
rect 3227 3044 3228 3048
rect 3222 3043 3228 3044
rect 3502 3048 3508 3049
rect 3502 3044 3503 3048
rect 3507 3044 3508 3048
rect 3590 3047 3591 3051
rect 3595 3047 3596 3051
rect 3590 3046 3596 3047
rect 3502 3043 3508 3044
rect 1896 3019 1898 3043
rect 2008 3019 2010 3043
rect 2184 3019 2186 3043
rect 2400 3019 2402 3043
rect 2648 3019 2650 3043
rect 2928 3019 2930 3043
rect 3224 3019 3226 3043
rect 3504 3019 3506 3043
rect 3592 3019 3594 3046
rect 1871 3018 1875 3019
rect 1871 3013 1875 3014
rect 1895 3018 1899 3019
rect 1895 3013 1899 3014
rect 2007 3018 2011 3019
rect 2007 3013 2011 3014
rect 2047 3018 2051 3019
rect 2047 3013 2051 3014
rect 2183 3018 2187 3019
rect 2183 3013 2187 3014
rect 2223 3018 2227 3019
rect 2223 3013 2227 3014
rect 2391 3018 2395 3019
rect 2391 3013 2395 3014
rect 2399 3018 2403 3019
rect 2399 3013 2403 3014
rect 2543 3018 2547 3019
rect 2543 3013 2547 3014
rect 2647 3018 2651 3019
rect 2647 3013 2651 3014
rect 2687 3018 2691 3019
rect 2687 3013 2691 3014
rect 2815 3018 2819 3019
rect 2815 3013 2819 3014
rect 2927 3018 2931 3019
rect 2927 3013 2931 3014
rect 3039 3018 3043 3019
rect 3039 3013 3043 3014
rect 3143 3018 3147 3019
rect 3143 3013 3147 3014
rect 3223 3018 3227 3019
rect 3223 3013 3227 3014
rect 3239 3018 3243 3019
rect 3239 3013 3243 3014
rect 3335 3018 3339 3019
rect 3335 3013 3339 3014
rect 3423 3018 3427 3019
rect 3423 3013 3427 3014
rect 3503 3018 3507 3019
rect 3503 3013 3507 3014
rect 3591 3018 3595 3019
rect 3591 3013 3595 3014
rect 110 3008 116 3009
rect 110 3004 111 3008
rect 115 3004 116 3008
rect 110 3003 116 3004
rect 1830 3008 1836 3009
rect 1830 3004 1831 3008
rect 1835 3004 1836 3008
rect 1830 3003 1836 3004
rect 112 2975 114 3003
rect 550 2990 556 2991
rect 550 2986 551 2990
rect 555 2986 556 2990
rect 550 2985 556 2986
rect 630 2990 636 2991
rect 630 2986 631 2990
rect 635 2986 636 2990
rect 630 2985 636 2986
rect 718 2990 724 2991
rect 718 2986 719 2990
rect 723 2986 724 2990
rect 718 2985 724 2986
rect 814 2990 820 2991
rect 814 2986 815 2990
rect 819 2986 820 2990
rect 814 2985 820 2986
rect 910 2990 916 2991
rect 910 2986 911 2990
rect 915 2986 916 2990
rect 910 2985 916 2986
rect 1006 2990 1012 2991
rect 1006 2986 1007 2990
rect 1011 2986 1012 2990
rect 1006 2985 1012 2986
rect 1094 2990 1100 2991
rect 1094 2986 1095 2990
rect 1099 2986 1100 2990
rect 1094 2985 1100 2986
rect 1190 2990 1196 2991
rect 1190 2986 1191 2990
rect 1195 2986 1196 2990
rect 1190 2985 1196 2986
rect 1286 2990 1292 2991
rect 1286 2986 1287 2990
rect 1291 2986 1292 2990
rect 1286 2985 1292 2986
rect 1382 2990 1388 2991
rect 1382 2986 1383 2990
rect 1387 2986 1388 2990
rect 1382 2985 1388 2986
rect 1478 2990 1484 2991
rect 1478 2986 1479 2990
rect 1483 2986 1484 2990
rect 1478 2985 1484 2986
rect 552 2975 554 2985
rect 632 2975 634 2985
rect 720 2975 722 2985
rect 816 2975 818 2985
rect 912 2975 914 2985
rect 1008 2975 1010 2985
rect 1096 2975 1098 2985
rect 1192 2975 1194 2985
rect 1288 2975 1290 2985
rect 1384 2975 1386 2985
rect 1480 2975 1482 2985
rect 1832 2975 1834 3003
rect 1872 2994 1874 3013
rect 1896 2997 1898 3013
rect 2048 2997 2050 3013
rect 2224 2997 2226 3013
rect 2392 2997 2394 3013
rect 2544 2997 2546 3013
rect 2688 2997 2690 3013
rect 2816 2997 2818 3013
rect 2928 2997 2930 3013
rect 3040 2997 3042 3013
rect 3144 2997 3146 3013
rect 3240 2997 3242 3013
rect 3336 2997 3338 3013
rect 3424 2997 3426 3013
rect 3504 2997 3506 3013
rect 1894 2996 1900 2997
rect 1870 2993 1876 2994
rect 1870 2989 1871 2993
rect 1875 2989 1876 2993
rect 1894 2992 1895 2996
rect 1899 2992 1900 2996
rect 1894 2991 1900 2992
rect 2046 2996 2052 2997
rect 2046 2992 2047 2996
rect 2051 2992 2052 2996
rect 2046 2991 2052 2992
rect 2222 2996 2228 2997
rect 2222 2992 2223 2996
rect 2227 2992 2228 2996
rect 2222 2991 2228 2992
rect 2390 2996 2396 2997
rect 2390 2992 2391 2996
rect 2395 2992 2396 2996
rect 2390 2991 2396 2992
rect 2542 2996 2548 2997
rect 2542 2992 2543 2996
rect 2547 2992 2548 2996
rect 2542 2991 2548 2992
rect 2686 2996 2692 2997
rect 2686 2992 2687 2996
rect 2691 2992 2692 2996
rect 2686 2991 2692 2992
rect 2814 2996 2820 2997
rect 2814 2992 2815 2996
rect 2819 2992 2820 2996
rect 2814 2991 2820 2992
rect 2926 2996 2932 2997
rect 2926 2992 2927 2996
rect 2931 2992 2932 2996
rect 2926 2991 2932 2992
rect 3038 2996 3044 2997
rect 3038 2992 3039 2996
rect 3043 2992 3044 2996
rect 3038 2991 3044 2992
rect 3142 2996 3148 2997
rect 3142 2992 3143 2996
rect 3147 2992 3148 2996
rect 3142 2991 3148 2992
rect 3238 2996 3244 2997
rect 3238 2992 3239 2996
rect 3243 2992 3244 2996
rect 3238 2991 3244 2992
rect 3334 2996 3340 2997
rect 3334 2992 3335 2996
rect 3339 2992 3340 2996
rect 3334 2991 3340 2992
rect 3422 2996 3428 2997
rect 3422 2992 3423 2996
rect 3427 2992 3428 2996
rect 3422 2991 3428 2992
rect 3502 2996 3508 2997
rect 3502 2992 3503 2996
rect 3507 2992 3508 2996
rect 3592 2994 3594 3013
rect 3502 2991 3508 2992
rect 3590 2993 3596 2994
rect 1870 2988 1876 2989
rect 3590 2989 3591 2993
rect 3595 2989 3596 2993
rect 3590 2988 3596 2989
rect 1870 2976 1876 2977
rect 111 2974 115 2975
rect 111 2969 115 2970
rect 471 2974 475 2975
rect 471 2969 475 2970
rect 551 2974 555 2975
rect 551 2969 555 2970
rect 575 2974 579 2975
rect 575 2969 579 2970
rect 631 2974 635 2975
rect 631 2969 635 2970
rect 687 2974 691 2975
rect 687 2969 691 2970
rect 719 2974 723 2975
rect 719 2969 723 2970
rect 807 2974 811 2975
rect 807 2969 811 2970
rect 815 2974 819 2975
rect 815 2969 819 2970
rect 911 2974 915 2975
rect 911 2969 915 2970
rect 943 2974 947 2975
rect 943 2969 947 2970
rect 1007 2974 1011 2975
rect 1007 2969 1011 2970
rect 1087 2974 1091 2975
rect 1087 2969 1091 2970
rect 1095 2974 1099 2975
rect 1095 2969 1099 2970
rect 1191 2974 1195 2975
rect 1191 2969 1195 2970
rect 1247 2974 1251 2975
rect 1247 2969 1251 2970
rect 1287 2974 1291 2975
rect 1287 2969 1291 2970
rect 1383 2974 1387 2975
rect 1383 2969 1387 2970
rect 1415 2974 1419 2975
rect 1415 2969 1419 2970
rect 1479 2974 1483 2975
rect 1479 2969 1483 2970
rect 1591 2974 1595 2975
rect 1591 2969 1595 2970
rect 1751 2974 1755 2975
rect 1751 2969 1755 2970
rect 1831 2974 1835 2975
rect 1870 2972 1871 2976
rect 1875 2972 1876 2976
rect 1870 2971 1876 2972
rect 3590 2976 3596 2977
rect 3590 2972 3591 2976
rect 3595 2972 3596 2976
rect 3590 2971 3596 2972
rect 1831 2969 1835 2970
rect 112 2941 114 2969
rect 472 2959 474 2969
rect 576 2959 578 2969
rect 688 2959 690 2969
rect 808 2959 810 2969
rect 944 2959 946 2969
rect 1088 2959 1090 2969
rect 1248 2959 1250 2969
rect 1416 2959 1418 2969
rect 1592 2959 1594 2969
rect 1752 2959 1754 2969
rect 470 2958 476 2959
rect 470 2954 471 2958
rect 475 2954 476 2958
rect 470 2953 476 2954
rect 574 2958 580 2959
rect 574 2954 575 2958
rect 579 2954 580 2958
rect 574 2953 580 2954
rect 686 2958 692 2959
rect 686 2954 687 2958
rect 691 2954 692 2958
rect 686 2953 692 2954
rect 806 2958 812 2959
rect 806 2954 807 2958
rect 811 2954 812 2958
rect 806 2953 812 2954
rect 942 2958 948 2959
rect 942 2954 943 2958
rect 947 2954 948 2958
rect 942 2953 948 2954
rect 1086 2958 1092 2959
rect 1086 2954 1087 2958
rect 1091 2954 1092 2958
rect 1086 2953 1092 2954
rect 1246 2958 1252 2959
rect 1246 2954 1247 2958
rect 1251 2954 1252 2958
rect 1246 2953 1252 2954
rect 1414 2958 1420 2959
rect 1414 2954 1415 2958
rect 1419 2954 1420 2958
rect 1414 2953 1420 2954
rect 1590 2958 1596 2959
rect 1590 2954 1591 2958
rect 1595 2954 1596 2958
rect 1590 2953 1596 2954
rect 1750 2958 1756 2959
rect 1750 2954 1751 2958
rect 1755 2954 1756 2958
rect 1750 2953 1756 2954
rect 1832 2941 1834 2969
rect 1872 2943 1874 2971
rect 1902 2958 1908 2959
rect 1902 2954 1903 2958
rect 1907 2954 1908 2958
rect 1902 2953 1908 2954
rect 2054 2958 2060 2959
rect 2054 2954 2055 2958
rect 2059 2954 2060 2958
rect 2054 2953 2060 2954
rect 2230 2958 2236 2959
rect 2230 2954 2231 2958
rect 2235 2954 2236 2958
rect 2230 2953 2236 2954
rect 2398 2958 2404 2959
rect 2398 2954 2399 2958
rect 2403 2954 2404 2958
rect 2398 2953 2404 2954
rect 2550 2958 2556 2959
rect 2550 2954 2551 2958
rect 2555 2954 2556 2958
rect 2550 2953 2556 2954
rect 2694 2958 2700 2959
rect 2694 2954 2695 2958
rect 2699 2954 2700 2958
rect 2694 2953 2700 2954
rect 2822 2958 2828 2959
rect 2822 2954 2823 2958
rect 2827 2954 2828 2958
rect 2822 2953 2828 2954
rect 2934 2958 2940 2959
rect 2934 2954 2935 2958
rect 2939 2954 2940 2958
rect 2934 2953 2940 2954
rect 3046 2958 3052 2959
rect 3046 2954 3047 2958
rect 3051 2954 3052 2958
rect 3046 2953 3052 2954
rect 3150 2958 3156 2959
rect 3150 2954 3151 2958
rect 3155 2954 3156 2958
rect 3150 2953 3156 2954
rect 3246 2958 3252 2959
rect 3246 2954 3247 2958
rect 3251 2954 3252 2958
rect 3246 2953 3252 2954
rect 3342 2958 3348 2959
rect 3342 2954 3343 2958
rect 3347 2954 3348 2958
rect 3342 2953 3348 2954
rect 3430 2958 3436 2959
rect 3430 2954 3431 2958
rect 3435 2954 3436 2958
rect 3430 2953 3436 2954
rect 3510 2958 3516 2959
rect 3510 2954 3511 2958
rect 3515 2954 3516 2958
rect 3510 2953 3516 2954
rect 1904 2943 1906 2953
rect 2056 2943 2058 2953
rect 2232 2943 2234 2953
rect 2400 2943 2402 2953
rect 2552 2943 2554 2953
rect 2696 2943 2698 2953
rect 2824 2943 2826 2953
rect 2936 2943 2938 2953
rect 3048 2943 3050 2953
rect 3152 2943 3154 2953
rect 3248 2943 3250 2953
rect 3344 2943 3346 2953
rect 3432 2943 3434 2953
rect 3512 2943 3514 2953
rect 3592 2943 3594 2971
rect 1871 2942 1875 2943
rect 110 2940 116 2941
rect 110 2936 111 2940
rect 115 2936 116 2940
rect 110 2935 116 2936
rect 1830 2940 1836 2941
rect 1830 2936 1831 2940
rect 1835 2936 1836 2940
rect 1871 2937 1875 2938
rect 1903 2942 1907 2943
rect 1903 2937 1907 2938
rect 2055 2942 2059 2943
rect 2055 2937 2059 2938
rect 2087 2942 2091 2943
rect 2087 2937 2091 2938
rect 2231 2942 2235 2943
rect 2231 2937 2235 2938
rect 2295 2942 2299 2943
rect 2295 2937 2299 2938
rect 2399 2942 2403 2943
rect 2399 2937 2403 2938
rect 2487 2942 2491 2943
rect 2487 2937 2491 2938
rect 2551 2942 2555 2943
rect 2551 2937 2555 2938
rect 2671 2942 2675 2943
rect 2671 2937 2675 2938
rect 2695 2942 2699 2943
rect 2695 2937 2699 2938
rect 2823 2942 2827 2943
rect 2823 2937 2827 2938
rect 2839 2942 2843 2943
rect 2839 2937 2843 2938
rect 2935 2942 2939 2943
rect 2935 2937 2939 2938
rect 2999 2942 3003 2943
rect 2999 2937 3003 2938
rect 3047 2942 3051 2943
rect 3047 2937 3051 2938
rect 3151 2942 3155 2943
rect 3151 2937 3155 2938
rect 3247 2942 3251 2943
rect 3247 2937 3251 2938
rect 3303 2942 3307 2943
rect 3303 2937 3307 2938
rect 3343 2942 3347 2943
rect 3343 2937 3347 2938
rect 3431 2942 3435 2943
rect 3431 2937 3435 2938
rect 3455 2942 3459 2943
rect 3455 2937 3459 2938
rect 3511 2942 3515 2943
rect 3511 2937 3515 2938
rect 3591 2942 3595 2943
rect 3591 2937 3595 2938
rect 1830 2935 1836 2936
rect 110 2923 116 2924
rect 110 2919 111 2923
rect 115 2919 116 2923
rect 1830 2923 1836 2924
rect 110 2918 116 2919
rect 462 2920 468 2921
rect 112 2899 114 2918
rect 462 2916 463 2920
rect 467 2916 468 2920
rect 462 2915 468 2916
rect 566 2920 572 2921
rect 566 2916 567 2920
rect 571 2916 572 2920
rect 566 2915 572 2916
rect 678 2920 684 2921
rect 678 2916 679 2920
rect 683 2916 684 2920
rect 678 2915 684 2916
rect 798 2920 804 2921
rect 798 2916 799 2920
rect 803 2916 804 2920
rect 798 2915 804 2916
rect 934 2920 940 2921
rect 934 2916 935 2920
rect 939 2916 940 2920
rect 934 2915 940 2916
rect 1078 2920 1084 2921
rect 1078 2916 1079 2920
rect 1083 2916 1084 2920
rect 1078 2915 1084 2916
rect 1238 2920 1244 2921
rect 1238 2916 1239 2920
rect 1243 2916 1244 2920
rect 1238 2915 1244 2916
rect 1406 2920 1412 2921
rect 1406 2916 1407 2920
rect 1411 2916 1412 2920
rect 1406 2915 1412 2916
rect 1582 2920 1588 2921
rect 1582 2916 1583 2920
rect 1587 2916 1588 2920
rect 1582 2915 1588 2916
rect 1742 2920 1748 2921
rect 1742 2916 1743 2920
rect 1747 2916 1748 2920
rect 1830 2919 1831 2923
rect 1835 2919 1836 2923
rect 1830 2918 1836 2919
rect 1742 2915 1748 2916
rect 464 2899 466 2915
rect 568 2899 570 2915
rect 680 2899 682 2915
rect 800 2899 802 2915
rect 936 2899 938 2915
rect 1080 2899 1082 2915
rect 1240 2899 1242 2915
rect 1408 2899 1410 2915
rect 1584 2899 1586 2915
rect 1744 2899 1746 2915
rect 1832 2899 1834 2918
rect 1872 2909 1874 2937
rect 1904 2927 1906 2937
rect 2088 2927 2090 2937
rect 2296 2927 2298 2937
rect 2488 2927 2490 2937
rect 2672 2927 2674 2937
rect 2840 2927 2842 2937
rect 3000 2927 3002 2937
rect 3152 2927 3154 2937
rect 3304 2927 3306 2937
rect 3456 2927 3458 2937
rect 1902 2926 1908 2927
rect 1902 2922 1903 2926
rect 1907 2922 1908 2926
rect 1902 2921 1908 2922
rect 2086 2926 2092 2927
rect 2086 2922 2087 2926
rect 2091 2922 2092 2926
rect 2086 2921 2092 2922
rect 2294 2926 2300 2927
rect 2294 2922 2295 2926
rect 2299 2922 2300 2926
rect 2294 2921 2300 2922
rect 2486 2926 2492 2927
rect 2486 2922 2487 2926
rect 2491 2922 2492 2926
rect 2486 2921 2492 2922
rect 2670 2926 2676 2927
rect 2670 2922 2671 2926
rect 2675 2922 2676 2926
rect 2670 2921 2676 2922
rect 2838 2926 2844 2927
rect 2838 2922 2839 2926
rect 2843 2922 2844 2926
rect 2838 2921 2844 2922
rect 2998 2926 3004 2927
rect 2998 2922 2999 2926
rect 3003 2922 3004 2926
rect 2998 2921 3004 2922
rect 3150 2926 3156 2927
rect 3150 2922 3151 2926
rect 3155 2922 3156 2926
rect 3150 2921 3156 2922
rect 3302 2926 3308 2927
rect 3302 2922 3303 2926
rect 3307 2922 3308 2926
rect 3302 2921 3308 2922
rect 3454 2926 3460 2927
rect 3454 2922 3455 2926
rect 3459 2922 3460 2926
rect 3454 2921 3460 2922
rect 3592 2909 3594 2937
rect 1870 2908 1876 2909
rect 1870 2904 1871 2908
rect 1875 2904 1876 2908
rect 1870 2903 1876 2904
rect 3590 2908 3596 2909
rect 3590 2904 3591 2908
rect 3595 2904 3596 2908
rect 3590 2903 3596 2904
rect 111 2898 115 2899
rect 111 2893 115 2894
rect 311 2898 315 2899
rect 311 2893 315 2894
rect 431 2898 435 2899
rect 431 2893 435 2894
rect 463 2898 467 2899
rect 463 2893 467 2894
rect 551 2898 555 2899
rect 551 2893 555 2894
rect 567 2898 571 2899
rect 567 2893 571 2894
rect 679 2898 683 2899
rect 679 2893 683 2894
rect 799 2898 803 2899
rect 799 2893 803 2894
rect 815 2898 819 2899
rect 815 2893 819 2894
rect 935 2898 939 2899
rect 935 2893 939 2894
rect 951 2898 955 2899
rect 951 2893 955 2894
rect 1079 2898 1083 2899
rect 1079 2893 1083 2894
rect 1087 2898 1091 2899
rect 1087 2893 1091 2894
rect 1223 2898 1227 2899
rect 1223 2893 1227 2894
rect 1239 2898 1243 2899
rect 1239 2893 1243 2894
rect 1359 2898 1363 2899
rect 1359 2893 1363 2894
rect 1407 2898 1411 2899
rect 1407 2893 1411 2894
rect 1495 2898 1499 2899
rect 1495 2893 1499 2894
rect 1583 2898 1587 2899
rect 1583 2893 1587 2894
rect 1631 2898 1635 2899
rect 1631 2893 1635 2894
rect 1743 2898 1747 2899
rect 1743 2893 1747 2894
rect 1831 2898 1835 2899
rect 1831 2893 1835 2894
rect 112 2874 114 2893
rect 312 2877 314 2893
rect 432 2877 434 2893
rect 552 2877 554 2893
rect 680 2877 682 2893
rect 816 2877 818 2893
rect 952 2877 954 2893
rect 1088 2877 1090 2893
rect 1224 2877 1226 2893
rect 1360 2877 1362 2893
rect 1496 2877 1498 2893
rect 1632 2877 1634 2893
rect 1744 2877 1746 2893
rect 310 2876 316 2877
rect 110 2873 116 2874
rect 110 2869 111 2873
rect 115 2869 116 2873
rect 310 2872 311 2876
rect 315 2872 316 2876
rect 310 2871 316 2872
rect 430 2876 436 2877
rect 430 2872 431 2876
rect 435 2872 436 2876
rect 430 2871 436 2872
rect 550 2876 556 2877
rect 550 2872 551 2876
rect 555 2872 556 2876
rect 550 2871 556 2872
rect 678 2876 684 2877
rect 678 2872 679 2876
rect 683 2872 684 2876
rect 678 2871 684 2872
rect 814 2876 820 2877
rect 814 2872 815 2876
rect 819 2872 820 2876
rect 814 2871 820 2872
rect 950 2876 956 2877
rect 950 2872 951 2876
rect 955 2872 956 2876
rect 950 2871 956 2872
rect 1086 2876 1092 2877
rect 1086 2872 1087 2876
rect 1091 2872 1092 2876
rect 1086 2871 1092 2872
rect 1222 2876 1228 2877
rect 1222 2872 1223 2876
rect 1227 2872 1228 2876
rect 1222 2871 1228 2872
rect 1358 2876 1364 2877
rect 1358 2872 1359 2876
rect 1363 2872 1364 2876
rect 1358 2871 1364 2872
rect 1494 2876 1500 2877
rect 1494 2872 1495 2876
rect 1499 2872 1500 2876
rect 1494 2871 1500 2872
rect 1630 2876 1636 2877
rect 1630 2872 1631 2876
rect 1635 2872 1636 2876
rect 1630 2871 1636 2872
rect 1742 2876 1748 2877
rect 1742 2872 1743 2876
rect 1747 2872 1748 2876
rect 1832 2874 1834 2893
rect 1870 2891 1876 2892
rect 1870 2887 1871 2891
rect 1875 2887 1876 2891
rect 3590 2891 3596 2892
rect 1870 2886 1876 2887
rect 1894 2888 1900 2889
rect 1742 2871 1748 2872
rect 1830 2873 1836 2874
rect 110 2868 116 2869
rect 1830 2869 1831 2873
rect 1835 2869 1836 2873
rect 1830 2868 1836 2869
rect 1872 2859 1874 2886
rect 1894 2884 1895 2888
rect 1899 2884 1900 2888
rect 1894 2883 1900 2884
rect 2078 2888 2084 2889
rect 2078 2884 2079 2888
rect 2083 2884 2084 2888
rect 2078 2883 2084 2884
rect 2286 2888 2292 2889
rect 2286 2884 2287 2888
rect 2291 2884 2292 2888
rect 2286 2883 2292 2884
rect 2478 2888 2484 2889
rect 2478 2884 2479 2888
rect 2483 2884 2484 2888
rect 2478 2883 2484 2884
rect 2662 2888 2668 2889
rect 2662 2884 2663 2888
rect 2667 2884 2668 2888
rect 2662 2883 2668 2884
rect 2830 2888 2836 2889
rect 2830 2884 2831 2888
rect 2835 2884 2836 2888
rect 2830 2883 2836 2884
rect 2990 2888 2996 2889
rect 2990 2884 2991 2888
rect 2995 2884 2996 2888
rect 2990 2883 2996 2884
rect 3142 2888 3148 2889
rect 3142 2884 3143 2888
rect 3147 2884 3148 2888
rect 3142 2883 3148 2884
rect 3294 2888 3300 2889
rect 3294 2884 3295 2888
rect 3299 2884 3300 2888
rect 3294 2883 3300 2884
rect 3446 2888 3452 2889
rect 3446 2884 3447 2888
rect 3451 2884 3452 2888
rect 3590 2887 3591 2891
rect 3595 2887 3596 2891
rect 3590 2886 3596 2887
rect 3446 2883 3452 2884
rect 1896 2859 1898 2883
rect 2080 2859 2082 2883
rect 2288 2859 2290 2883
rect 2480 2859 2482 2883
rect 2664 2859 2666 2883
rect 2832 2859 2834 2883
rect 2992 2859 2994 2883
rect 3144 2859 3146 2883
rect 3296 2859 3298 2883
rect 3448 2859 3450 2883
rect 3592 2859 3594 2886
rect 1871 2858 1875 2859
rect 110 2856 116 2857
rect 110 2852 111 2856
rect 115 2852 116 2856
rect 110 2851 116 2852
rect 1830 2856 1836 2857
rect 1830 2852 1831 2856
rect 1835 2852 1836 2856
rect 1871 2853 1875 2854
rect 1895 2858 1899 2859
rect 1895 2853 1899 2854
rect 2079 2858 2083 2859
rect 2079 2853 2083 2854
rect 2135 2858 2139 2859
rect 2135 2853 2139 2854
rect 2263 2858 2267 2859
rect 2263 2853 2267 2854
rect 2287 2858 2291 2859
rect 2287 2853 2291 2854
rect 2391 2858 2395 2859
rect 2391 2853 2395 2854
rect 2479 2858 2483 2859
rect 2479 2853 2483 2854
rect 2519 2858 2523 2859
rect 2519 2853 2523 2854
rect 2647 2858 2651 2859
rect 2647 2853 2651 2854
rect 2663 2858 2667 2859
rect 2663 2853 2667 2854
rect 2767 2858 2771 2859
rect 2767 2853 2771 2854
rect 2831 2858 2835 2859
rect 2831 2853 2835 2854
rect 2887 2858 2891 2859
rect 2887 2853 2891 2854
rect 2991 2858 2995 2859
rect 2991 2853 2995 2854
rect 3007 2858 3011 2859
rect 3007 2853 3011 2854
rect 3135 2858 3139 2859
rect 3135 2853 3139 2854
rect 3143 2858 3147 2859
rect 3143 2853 3147 2854
rect 3295 2858 3299 2859
rect 3295 2853 3299 2854
rect 3447 2858 3451 2859
rect 3447 2853 3451 2854
rect 3591 2858 3595 2859
rect 3591 2853 3595 2854
rect 1830 2851 1836 2852
rect 112 2823 114 2851
rect 318 2838 324 2839
rect 318 2834 319 2838
rect 323 2834 324 2838
rect 318 2833 324 2834
rect 438 2838 444 2839
rect 438 2834 439 2838
rect 443 2834 444 2838
rect 438 2833 444 2834
rect 558 2838 564 2839
rect 558 2834 559 2838
rect 563 2834 564 2838
rect 558 2833 564 2834
rect 686 2838 692 2839
rect 686 2834 687 2838
rect 691 2834 692 2838
rect 686 2833 692 2834
rect 822 2838 828 2839
rect 822 2834 823 2838
rect 827 2834 828 2838
rect 822 2833 828 2834
rect 958 2838 964 2839
rect 958 2834 959 2838
rect 963 2834 964 2838
rect 958 2833 964 2834
rect 1094 2838 1100 2839
rect 1094 2834 1095 2838
rect 1099 2834 1100 2838
rect 1094 2833 1100 2834
rect 1230 2838 1236 2839
rect 1230 2834 1231 2838
rect 1235 2834 1236 2838
rect 1230 2833 1236 2834
rect 1366 2838 1372 2839
rect 1366 2834 1367 2838
rect 1371 2834 1372 2838
rect 1366 2833 1372 2834
rect 1502 2838 1508 2839
rect 1502 2834 1503 2838
rect 1507 2834 1508 2838
rect 1502 2833 1508 2834
rect 1638 2838 1644 2839
rect 1638 2834 1639 2838
rect 1643 2834 1644 2838
rect 1638 2833 1644 2834
rect 1750 2838 1756 2839
rect 1750 2834 1751 2838
rect 1755 2834 1756 2838
rect 1750 2833 1756 2834
rect 320 2823 322 2833
rect 440 2823 442 2833
rect 560 2823 562 2833
rect 688 2823 690 2833
rect 824 2823 826 2833
rect 960 2823 962 2833
rect 1096 2823 1098 2833
rect 1232 2823 1234 2833
rect 1368 2823 1370 2833
rect 1504 2823 1506 2833
rect 1640 2823 1642 2833
rect 1752 2823 1754 2833
rect 1832 2823 1834 2851
rect 1872 2834 1874 2853
rect 2136 2837 2138 2853
rect 2264 2837 2266 2853
rect 2392 2837 2394 2853
rect 2520 2837 2522 2853
rect 2648 2837 2650 2853
rect 2768 2837 2770 2853
rect 2888 2837 2890 2853
rect 3008 2837 3010 2853
rect 3136 2837 3138 2853
rect 2134 2836 2140 2837
rect 1870 2833 1876 2834
rect 1870 2829 1871 2833
rect 1875 2829 1876 2833
rect 2134 2832 2135 2836
rect 2139 2832 2140 2836
rect 2134 2831 2140 2832
rect 2262 2836 2268 2837
rect 2262 2832 2263 2836
rect 2267 2832 2268 2836
rect 2262 2831 2268 2832
rect 2390 2836 2396 2837
rect 2390 2832 2391 2836
rect 2395 2832 2396 2836
rect 2390 2831 2396 2832
rect 2518 2836 2524 2837
rect 2518 2832 2519 2836
rect 2523 2832 2524 2836
rect 2518 2831 2524 2832
rect 2646 2836 2652 2837
rect 2646 2832 2647 2836
rect 2651 2832 2652 2836
rect 2646 2831 2652 2832
rect 2766 2836 2772 2837
rect 2766 2832 2767 2836
rect 2771 2832 2772 2836
rect 2766 2831 2772 2832
rect 2886 2836 2892 2837
rect 2886 2832 2887 2836
rect 2891 2832 2892 2836
rect 2886 2831 2892 2832
rect 3006 2836 3012 2837
rect 3006 2832 3007 2836
rect 3011 2832 3012 2836
rect 3006 2831 3012 2832
rect 3134 2836 3140 2837
rect 3134 2832 3135 2836
rect 3139 2832 3140 2836
rect 3592 2834 3594 2853
rect 3134 2831 3140 2832
rect 3590 2833 3596 2834
rect 1870 2828 1876 2829
rect 3590 2829 3591 2833
rect 3595 2829 3596 2833
rect 3590 2828 3596 2829
rect 111 2822 115 2823
rect 111 2817 115 2818
rect 167 2822 171 2823
rect 167 2817 171 2818
rect 303 2822 307 2823
rect 303 2817 307 2818
rect 319 2822 323 2823
rect 319 2817 323 2818
rect 439 2822 443 2823
rect 439 2817 443 2818
rect 447 2822 451 2823
rect 447 2817 451 2818
rect 559 2822 563 2823
rect 559 2817 563 2818
rect 607 2822 611 2823
rect 607 2817 611 2818
rect 687 2822 691 2823
rect 687 2817 691 2818
rect 783 2822 787 2823
rect 783 2817 787 2818
rect 823 2822 827 2823
rect 823 2817 827 2818
rect 959 2822 963 2823
rect 959 2817 963 2818
rect 1095 2822 1099 2823
rect 1095 2817 1099 2818
rect 1143 2822 1147 2823
rect 1143 2817 1147 2818
rect 1231 2822 1235 2823
rect 1231 2817 1235 2818
rect 1335 2822 1339 2823
rect 1335 2817 1339 2818
rect 1367 2822 1371 2823
rect 1367 2817 1371 2818
rect 1503 2822 1507 2823
rect 1503 2817 1507 2818
rect 1535 2822 1539 2823
rect 1535 2817 1539 2818
rect 1639 2822 1643 2823
rect 1639 2817 1643 2818
rect 1735 2822 1739 2823
rect 1735 2817 1739 2818
rect 1751 2822 1755 2823
rect 1751 2817 1755 2818
rect 1831 2822 1835 2823
rect 1831 2817 1835 2818
rect 112 2789 114 2817
rect 168 2807 170 2817
rect 304 2807 306 2817
rect 448 2807 450 2817
rect 608 2807 610 2817
rect 784 2807 786 2817
rect 960 2807 962 2817
rect 1144 2807 1146 2817
rect 1336 2807 1338 2817
rect 1536 2807 1538 2817
rect 1736 2807 1738 2817
rect 166 2806 172 2807
rect 166 2802 167 2806
rect 171 2802 172 2806
rect 166 2801 172 2802
rect 302 2806 308 2807
rect 302 2802 303 2806
rect 307 2802 308 2806
rect 302 2801 308 2802
rect 446 2806 452 2807
rect 446 2802 447 2806
rect 451 2802 452 2806
rect 446 2801 452 2802
rect 606 2806 612 2807
rect 606 2802 607 2806
rect 611 2802 612 2806
rect 606 2801 612 2802
rect 782 2806 788 2807
rect 782 2802 783 2806
rect 787 2802 788 2806
rect 782 2801 788 2802
rect 958 2806 964 2807
rect 958 2802 959 2806
rect 963 2802 964 2806
rect 958 2801 964 2802
rect 1142 2806 1148 2807
rect 1142 2802 1143 2806
rect 1147 2802 1148 2806
rect 1142 2801 1148 2802
rect 1334 2806 1340 2807
rect 1334 2802 1335 2806
rect 1339 2802 1340 2806
rect 1334 2801 1340 2802
rect 1534 2806 1540 2807
rect 1534 2802 1535 2806
rect 1539 2802 1540 2806
rect 1534 2801 1540 2802
rect 1734 2806 1740 2807
rect 1734 2802 1735 2806
rect 1739 2802 1740 2806
rect 1734 2801 1740 2802
rect 1832 2789 1834 2817
rect 1870 2816 1876 2817
rect 1870 2812 1871 2816
rect 1875 2812 1876 2816
rect 1870 2811 1876 2812
rect 3590 2816 3596 2817
rect 3590 2812 3591 2816
rect 3595 2812 3596 2816
rect 3590 2811 3596 2812
rect 110 2788 116 2789
rect 110 2784 111 2788
rect 115 2784 116 2788
rect 110 2783 116 2784
rect 1830 2788 1836 2789
rect 1830 2784 1831 2788
rect 1835 2784 1836 2788
rect 1830 2783 1836 2784
rect 1872 2775 1874 2811
rect 2142 2798 2148 2799
rect 2142 2794 2143 2798
rect 2147 2794 2148 2798
rect 2142 2793 2148 2794
rect 2270 2798 2276 2799
rect 2270 2794 2271 2798
rect 2275 2794 2276 2798
rect 2270 2793 2276 2794
rect 2398 2798 2404 2799
rect 2398 2794 2399 2798
rect 2403 2794 2404 2798
rect 2398 2793 2404 2794
rect 2526 2798 2532 2799
rect 2526 2794 2527 2798
rect 2531 2794 2532 2798
rect 2526 2793 2532 2794
rect 2654 2798 2660 2799
rect 2654 2794 2655 2798
rect 2659 2794 2660 2798
rect 2654 2793 2660 2794
rect 2774 2798 2780 2799
rect 2774 2794 2775 2798
rect 2779 2794 2780 2798
rect 2774 2793 2780 2794
rect 2894 2798 2900 2799
rect 2894 2794 2895 2798
rect 2899 2794 2900 2798
rect 2894 2793 2900 2794
rect 3014 2798 3020 2799
rect 3014 2794 3015 2798
rect 3019 2794 3020 2798
rect 3014 2793 3020 2794
rect 3142 2798 3148 2799
rect 3142 2794 3143 2798
rect 3147 2794 3148 2798
rect 3142 2793 3148 2794
rect 2144 2775 2146 2793
rect 2272 2775 2274 2793
rect 2400 2775 2402 2793
rect 2528 2775 2530 2793
rect 2656 2775 2658 2793
rect 2776 2775 2778 2793
rect 2896 2775 2898 2793
rect 3016 2775 3018 2793
rect 3144 2775 3146 2793
rect 3592 2775 3594 2811
rect 1871 2774 1875 2775
rect 110 2771 116 2772
rect 110 2767 111 2771
rect 115 2767 116 2771
rect 1830 2771 1836 2772
rect 110 2766 116 2767
rect 158 2768 164 2769
rect 112 2743 114 2766
rect 158 2764 159 2768
rect 163 2764 164 2768
rect 158 2763 164 2764
rect 294 2768 300 2769
rect 294 2764 295 2768
rect 299 2764 300 2768
rect 294 2763 300 2764
rect 438 2768 444 2769
rect 438 2764 439 2768
rect 443 2764 444 2768
rect 438 2763 444 2764
rect 598 2768 604 2769
rect 598 2764 599 2768
rect 603 2764 604 2768
rect 598 2763 604 2764
rect 774 2768 780 2769
rect 774 2764 775 2768
rect 779 2764 780 2768
rect 774 2763 780 2764
rect 950 2768 956 2769
rect 950 2764 951 2768
rect 955 2764 956 2768
rect 950 2763 956 2764
rect 1134 2768 1140 2769
rect 1134 2764 1135 2768
rect 1139 2764 1140 2768
rect 1134 2763 1140 2764
rect 1326 2768 1332 2769
rect 1326 2764 1327 2768
rect 1331 2764 1332 2768
rect 1326 2763 1332 2764
rect 1526 2768 1532 2769
rect 1526 2764 1527 2768
rect 1531 2764 1532 2768
rect 1526 2763 1532 2764
rect 1726 2768 1732 2769
rect 1726 2764 1727 2768
rect 1731 2764 1732 2768
rect 1830 2767 1831 2771
rect 1835 2767 1836 2771
rect 1871 2769 1875 2770
rect 2143 2774 2147 2775
rect 2143 2769 2147 2770
rect 2231 2774 2235 2775
rect 2231 2769 2235 2770
rect 2271 2774 2275 2775
rect 2271 2769 2275 2770
rect 2311 2774 2315 2775
rect 2311 2769 2315 2770
rect 2391 2774 2395 2775
rect 2391 2769 2395 2770
rect 2399 2774 2403 2775
rect 2399 2769 2403 2770
rect 2471 2774 2475 2775
rect 2471 2769 2475 2770
rect 2527 2774 2531 2775
rect 2527 2769 2531 2770
rect 2551 2774 2555 2775
rect 2551 2769 2555 2770
rect 2639 2774 2643 2775
rect 2639 2769 2643 2770
rect 2655 2774 2659 2775
rect 2655 2769 2659 2770
rect 2727 2774 2731 2775
rect 2727 2769 2731 2770
rect 2775 2774 2779 2775
rect 2775 2769 2779 2770
rect 2815 2774 2819 2775
rect 2815 2769 2819 2770
rect 2895 2774 2899 2775
rect 2895 2769 2899 2770
rect 2903 2774 2907 2775
rect 2903 2769 2907 2770
rect 2991 2774 2995 2775
rect 2991 2769 2995 2770
rect 3015 2774 3019 2775
rect 3015 2769 3019 2770
rect 3143 2774 3147 2775
rect 3143 2769 3147 2770
rect 3591 2774 3595 2775
rect 3591 2769 3595 2770
rect 1830 2766 1836 2767
rect 1726 2763 1732 2764
rect 160 2743 162 2763
rect 296 2743 298 2763
rect 440 2743 442 2763
rect 600 2743 602 2763
rect 776 2743 778 2763
rect 952 2743 954 2763
rect 1136 2743 1138 2763
rect 1328 2743 1330 2763
rect 1528 2743 1530 2763
rect 1728 2743 1730 2763
rect 1832 2743 1834 2766
rect 111 2742 115 2743
rect 111 2737 115 2738
rect 135 2742 139 2743
rect 135 2737 139 2738
rect 159 2742 163 2743
rect 159 2737 163 2738
rect 247 2742 251 2743
rect 247 2737 251 2738
rect 295 2742 299 2743
rect 295 2737 299 2738
rect 391 2742 395 2743
rect 391 2737 395 2738
rect 439 2742 443 2743
rect 439 2737 443 2738
rect 551 2742 555 2743
rect 551 2737 555 2738
rect 599 2742 603 2743
rect 599 2737 603 2738
rect 711 2742 715 2743
rect 711 2737 715 2738
rect 775 2742 779 2743
rect 775 2737 779 2738
rect 879 2742 883 2743
rect 879 2737 883 2738
rect 951 2742 955 2743
rect 951 2737 955 2738
rect 1039 2742 1043 2743
rect 1039 2737 1043 2738
rect 1135 2742 1139 2743
rect 1135 2737 1139 2738
rect 1199 2742 1203 2743
rect 1199 2737 1203 2738
rect 1327 2742 1331 2743
rect 1327 2737 1331 2738
rect 1359 2742 1363 2743
rect 1359 2737 1363 2738
rect 1519 2742 1523 2743
rect 1519 2737 1523 2738
rect 1527 2742 1531 2743
rect 1527 2737 1531 2738
rect 1687 2742 1691 2743
rect 1687 2737 1691 2738
rect 1727 2742 1731 2743
rect 1727 2737 1731 2738
rect 1831 2742 1835 2743
rect 1872 2741 1874 2769
rect 2232 2759 2234 2769
rect 2312 2759 2314 2769
rect 2392 2759 2394 2769
rect 2472 2759 2474 2769
rect 2552 2759 2554 2769
rect 2640 2759 2642 2769
rect 2728 2759 2730 2769
rect 2816 2759 2818 2769
rect 2904 2759 2906 2769
rect 2992 2759 2994 2769
rect 2230 2758 2236 2759
rect 2230 2754 2231 2758
rect 2235 2754 2236 2758
rect 2230 2753 2236 2754
rect 2310 2758 2316 2759
rect 2310 2754 2311 2758
rect 2315 2754 2316 2758
rect 2310 2753 2316 2754
rect 2390 2758 2396 2759
rect 2390 2754 2391 2758
rect 2395 2754 2396 2758
rect 2390 2753 2396 2754
rect 2470 2758 2476 2759
rect 2470 2754 2471 2758
rect 2475 2754 2476 2758
rect 2470 2753 2476 2754
rect 2550 2758 2556 2759
rect 2550 2754 2551 2758
rect 2555 2754 2556 2758
rect 2550 2753 2556 2754
rect 2638 2758 2644 2759
rect 2638 2754 2639 2758
rect 2643 2754 2644 2758
rect 2638 2753 2644 2754
rect 2726 2758 2732 2759
rect 2726 2754 2727 2758
rect 2731 2754 2732 2758
rect 2726 2753 2732 2754
rect 2814 2758 2820 2759
rect 2814 2754 2815 2758
rect 2819 2754 2820 2758
rect 2814 2753 2820 2754
rect 2902 2758 2908 2759
rect 2902 2754 2903 2758
rect 2907 2754 2908 2758
rect 2902 2753 2908 2754
rect 2990 2758 2996 2759
rect 2990 2754 2991 2758
rect 2995 2754 2996 2758
rect 2990 2753 2996 2754
rect 3592 2741 3594 2769
rect 1831 2737 1835 2738
rect 1870 2740 1876 2741
rect 112 2718 114 2737
rect 136 2721 138 2737
rect 248 2721 250 2737
rect 392 2721 394 2737
rect 552 2721 554 2737
rect 712 2721 714 2737
rect 880 2721 882 2737
rect 1040 2721 1042 2737
rect 1200 2721 1202 2737
rect 1360 2721 1362 2737
rect 1520 2721 1522 2737
rect 1688 2721 1690 2737
rect 134 2720 140 2721
rect 110 2717 116 2718
rect 110 2713 111 2717
rect 115 2713 116 2717
rect 134 2716 135 2720
rect 139 2716 140 2720
rect 134 2715 140 2716
rect 246 2720 252 2721
rect 246 2716 247 2720
rect 251 2716 252 2720
rect 246 2715 252 2716
rect 390 2720 396 2721
rect 390 2716 391 2720
rect 395 2716 396 2720
rect 390 2715 396 2716
rect 550 2720 556 2721
rect 550 2716 551 2720
rect 555 2716 556 2720
rect 550 2715 556 2716
rect 710 2720 716 2721
rect 710 2716 711 2720
rect 715 2716 716 2720
rect 710 2715 716 2716
rect 878 2720 884 2721
rect 878 2716 879 2720
rect 883 2716 884 2720
rect 878 2715 884 2716
rect 1038 2720 1044 2721
rect 1038 2716 1039 2720
rect 1043 2716 1044 2720
rect 1038 2715 1044 2716
rect 1198 2720 1204 2721
rect 1198 2716 1199 2720
rect 1203 2716 1204 2720
rect 1198 2715 1204 2716
rect 1358 2720 1364 2721
rect 1358 2716 1359 2720
rect 1363 2716 1364 2720
rect 1358 2715 1364 2716
rect 1518 2720 1524 2721
rect 1518 2716 1519 2720
rect 1523 2716 1524 2720
rect 1518 2715 1524 2716
rect 1686 2720 1692 2721
rect 1686 2716 1687 2720
rect 1691 2716 1692 2720
rect 1832 2718 1834 2737
rect 1870 2736 1871 2740
rect 1875 2736 1876 2740
rect 1870 2735 1876 2736
rect 3590 2740 3596 2741
rect 3590 2736 3591 2740
rect 3595 2736 3596 2740
rect 3590 2735 3596 2736
rect 1870 2723 1876 2724
rect 1870 2719 1871 2723
rect 1875 2719 1876 2723
rect 3590 2723 3596 2724
rect 1870 2718 1876 2719
rect 2222 2720 2228 2721
rect 1686 2715 1692 2716
rect 1830 2717 1836 2718
rect 110 2712 116 2713
rect 1830 2713 1831 2717
rect 1835 2713 1836 2717
rect 1830 2712 1836 2713
rect 110 2700 116 2701
rect 110 2696 111 2700
rect 115 2696 116 2700
rect 110 2695 116 2696
rect 1830 2700 1836 2701
rect 1830 2696 1831 2700
rect 1835 2696 1836 2700
rect 1872 2699 1874 2718
rect 2222 2716 2223 2720
rect 2227 2716 2228 2720
rect 2222 2715 2228 2716
rect 2302 2720 2308 2721
rect 2302 2716 2303 2720
rect 2307 2716 2308 2720
rect 2302 2715 2308 2716
rect 2382 2720 2388 2721
rect 2382 2716 2383 2720
rect 2387 2716 2388 2720
rect 2382 2715 2388 2716
rect 2462 2720 2468 2721
rect 2462 2716 2463 2720
rect 2467 2716 2468 2720
rect 2462 2715 2468 2716
rect 2542 2720 2548 2721
rect 2542 2716 2543 2720
rect 2547 2716 2548 2720
rect 2542 2715 2548 2716
rect 2630 2720 2636 2721
rect 2630 2716 2631 2720
rect 2635 2716 2636 2720
rect 2630 2715 2636 2716
rect 2718 2720 2724 2721
rect 2718 2716 2719 2720
rect 2723 2716 2724 2720
rect 2718 2715 2724 2716
rect 2806 2720 2812 2721
rect 2806 2716 2807 2720
rect 2811 2716 2812 2720
rect 2806 2715 2812 2716
rect 2894 2720 2900 2721
rect 2894 2716 2895 2720
rect 2899 2716 2900 2720
rect 2894 2715 2900 2716
rect 2982 2720 2988 2721
rect 2982 2716 2983 2720
rect 2987 2716 2988 2720
rect 3590 2719 3591 2723
rect 3595 2719 3596 2723
rect 3590 2718 3596 2719
rect 2982 2715 2988 2716
rect 2224 2699 2226 2715
rect 2304 2699 2306 2715
rect 2384 2699 2386 2715
rect 2464 2699 2466 2715
rect 2544 2699 2546 2715
rect 2632 2699 2634 2715
rect 2720 2699 2722 2715
rect 2808 2699 2810 2715
rect 2896 2699 2898 2715
rect 2984 2699 2986 2715
rect 3592 2699 3594 2718
rect 1830 2695 1836 2696
rect 1871 2698 1875 2699
rect 112 2667 114 2695
rect 142 2682 148 2683
rect 142 2678 143 2682
rect 147 2678 148 2682
rect 142 2677 148 2678
rect 254 2682 260 2683
rect 254 2678 255 2682
rect 259 2678 260 2682
rect 254 2677 260 2678
rect 398 2682 404 2683
rect 398 2678 399 2682
rect 403 2678 404 2682
rect 398 2677 404 2678
rect 558 2682 564 2683
rect 558 2678 559 2682
rect 563 2678 564 2682
rect 558 2677 564 2678
rect 718 2682 724 2683
rect 718 2678 719 2682
rect 723 2678 724 2682
rect 718 2677 724 2678
rect 886 2682 892 2683
rect 886 2678 887 2682
rect 891 2678 892 2682
rect 886 2677 892 2678
rect 1046 2682 1052 2683
rect 1046 2678 1047 2682
rect 1051 2678 1052 2682
rect 1046 2677 1052 2678
rect 1206 2682 1212 2683
rect 1206 2678 1207 2682
rect 1211 2678 1212 2682
rect 1206 2677 1212 2678
rect 1366 2682 1372 2683
rect 1366 2678 1367 2682
rect 1371 2678 1372 2682
rect 1366 2677 1372 2678
rect 1526 2682 1532 2683
rect 1526 2678 1527 2682
rect 1531 2678 1532 2682
rect 1526 2677 1532 2678
rect 1694 2682 1700 2683
rect 1694 2678 1695 2682
rect 1699 2678 1700 2682
rect 1694 2677 1700 2678
rect 144 2667 146 2677
rect 256 2667 258 2677
rect 400 2667 402 2677
rect 560 2667 562 2677
rect 720 2667 722 2677
rect 888 2667 890 2677
rect 1048 2667 1050 2677
rect 1208 2667 1210 2677
rect 1368 2667 1370 2677
rect 1528 2667 1530 2677
rect 1696 2667 1698 2677
rect 1832 2667 1834 2695
rect 1871 2693 1875 2694
rect 2223 2698 2227 2699
rect 2223 2693 2227 2694
rect 2239 2698 2243 2699
rect 2239 2693 2243 2694
rect 2303 2698 2307 2699
rect 2303 2693 2307 2694
rect 2319 2698 2323 2699
rect 2319 2693 2323 2694
rect 2383 2698 2387 2699
rect 2383 2693 2387 2694
rect 2399 2698 2403 2699
rect 2399 2693 2403 2694
rect 2463 2698 2467 2699
rect 2463 2693 2467 2694
rect 2479 2698 2483 2699
rect 2479 2693 2483 2694
rect 2543 2698 2547 2699
rect 2543 2693 2547 2694
rect 2559 2698 2563 2699
rect 2559 2693 2563 2694
rect 2631 2698 2635 2699
rect 2631 2693 2635 2694
rect 2639 2698 2643 2699
rect 2639 2693 2643 2694
rect 2719 2698 2723 2699
rect 2719 2693 2723 2694
rect 2799 2698 2803 2699
rect 2799 2693 2803 2694
rect 2807 2698 2811 2699
rect 2807 2693 2811 2694
rect 2879 2698 2883 2699
rect 2879 2693 2883 2694
rect 2895 2698 2899 2699
rect 2895 2693 2899 2694
rect 2959 2698 2963 2699
rect 2959 2693 2963 2694
rect 2983 2698 2987 2699
rect 2983 2693 2987 2694
rect 3591 2698 3595 2699
rect 3591 2693 3595 2694
rect 1872 2674 1874 2693
rect 2240 2677 2242 2693
rect 2320 2677 2322 2693
rect 2400 2677 2402 2693
rect 2480 2677 2482 2693
rect 2560 2677 2562 2693
rect 2640 2677 2642 2693
rect 2720 2677 2722 2693
rect 2800 2677 2802 2693
rect 2880 2677 2882 2693
rect 2960 2677 2962 2693
rect 2238 2676 2244 2677
rect 1870 2673 1876 2674
rect 1870 2669 1871 2673
rect 1875 2669 1876 2673
rect 2238 2672 2239 2676
rect 2243 2672 2244 2676
rect 2238 2671 2244 2672
rect 2318 2676 2324 2677
rect 2318 2672 2319 2676
rect 2323 2672 2324 2676
rect 2318 2671 2324 2672
rect 2398 2676 2404 2677
rect 2398 2672 2399 2676
rect 2403 2672 2404 2676
rect 2398 2671 2404 2672
rect 2478 2676 2484 2677
rect 2478 2672 2479 2676
rect 2483 2672 2484 2676
rect 2478 2671 2484 2672
rect 2558 2676 2564 2677
rect 2558 2672 2559 2676
rect 2563 2672 2564 2676
rect 2558 2671 2564 2672
rect 2638 2676 2644 2677
rect 2638 2672 2639 2676
rect 2643 2672 2644 2676
rect 2638 2671 2644 2672
rect 2718 2676 2724 2677
rect 2718 2672 2719 2676
rect 2723 2672 2724 2676
rect 2718 2671 2724 2672
rect 2798 2676 2804 2677
rect 2798 2672 2799 2676
rect 2803 2672 2804 2676
rect 2798 2671 2804 2672
rect 2878 2676 2884 2677
rect 2878 2672 2879 2676
rect 2883 2672 2884 2676
rect 2878 2671 2884 2672
rect 2958 2676 2964 2677
rect 2958 2672 2959 2676
rect 2963 2672 2964 2676
rect 3592 2674 3594 2693
rect 2958 2671 2964 2672
rect 3590 2673 3596 2674
rect 1870 2668 1876 2669
rect 3590 2669 3591 2673
rect 3595 2669 3596 2673
rect 3590 2668 3596 2669
rect 111 2666 115 2667
rect 111 2661 115 2662
rect 143 2666 147 2667
rect 143 2661 147 2662
rect 255 2666 259 2667
rect 255 2661 259 2662
rect 399 2666 403 2667
rect 399 2661 403 2662
rect 551 2666 555 2667
rect 551 2661 555 2662
rect 559 2666 563 2667
rect 559 2661 563 2662
rect 711 2666 715 2667
rect 711 2661 715 2662
rect 719 2666 723 2667
rect 719 2661 723 2662
rect 879 2666 883 2667
rect 879 2661 883 2662
rect 887 2666 891 2667
rect 887 2661 891 2662
rect 1047 2666 1051 2667
rect 1047 2661 1051 2662
rect 1207 2666 1211 2667
rect 1207 2661 1211 2662
rect 1215 2666 1219 2667
rect 1215 2661 1219 2662
rect 1367 2666 1371 2667
rect 1367 2661 1371 2662
rect 1391 2666 1395 2667
rect 1391 2661 1395 2662
rect 1527 2666 1531 2667
rect 1527 2661 1531 2662
rect 1567 2666 1571 2667
rect 1567 2661 1571 2662
rect 1695 2666 1699 2667
rect 1695 2661 1699 2662
rect 1831 2666 1835 2667
rect 1831 2661 1835 2662
rect 112 2633 114 2661
rect 144 2651 146 2661
rect 256 2651 258 2661
rect 400 2651 402 2661
rect 552 2651 554 2661
rect 712 2651 714 2661
rect 880 2651 882 2661
rect 1048 2651 1050 2661
rect 1216 2651 1218 2661
rect 1392 2651 1394 2661
rect 1568 2651 1570 2661
rect 142 2650 148 2651
rect 142 2646 143 2650
rect 147 2646 148 2650
rect 142 2645 148 2646
rect 254 2650 260 2651
rect 254 2646 255 2650
rect 259 2646 260 2650
rect 254 2645 260 2646
rect 398 2650 404 2651
rect 398 2646 399 2650
rect 403 2646 404 2650
rect 398 2645 404 2646
rect 550 2650 556 2651
rect 550 2646 551 2650
rect 555 2646 556 2650
rect 550 2645 556 2646
rect 710 2650 716 2651
rect 710 2646 711 2650
rect 715 2646 716 2650
rect 710 2645 716 2646
rect 878 2650 884 2651
rect 878 2646 879 2650
rect 883 2646 884 2650
rect 878 2645 884 2646
rect 1046 2650 1052 2651
rect 1046 2646 1047 2650
rect 1051 2646 1052 2650
rect 1046 2645 1052 2646
rect 1214 2650 1220 2651
rect 1214 2646 1215 2650
rect 1219 2646 1220 2650
rect 1214 2645 1220 2646
rect 1390 2650 1396 2651
rect 1390 2646 1391 2650
rect 1395 2646 1396 2650
rect 1390 2645 1396 2646
rect 1566 2650 1572 2651
rect 1566 2646 1567 2650
rect 1571 2646 1572 2650
rect 1566 2645 1572 2646
rect 1832 2633 1834 2661
rect 1870 2656 1876 2657
rect 1870 2652 1871 2656
rect 1875 2652 1876 2656
rect 1870 2651 1876 2652
rect 3590 2656 3596 2657
rect 3590 2652 3591 2656
rect 3595 2652 3596 2656
rect 3590 2651 3596 2652
rect 110 2632 116 2633
rect 110 2628 111 2632
rect 115 2628 116 2632
rect 110 2627 116 2628
rect 1830 2632 1836 2633
rect 1830 2628 1831 2632
rect 1835 2628 1836 2632
rect 1830 2627 1836 2628
rect 110 2615 116 2616
rect 110 2611 111 2615
rect 115 2611 116 2615
rect 1830 2615 1836 2616
rect 1872 2615 1874 2651
rect 2246 2638 2252 2639
rect 2246 2634 2247 2638
rect 2251 2634 2252 2638
rect 2246 2633 2252 2634
rect 2326 2638 2332 2639
rect 2326 2634 2327 2638
rect 2331 2634 2332 2638
rect 2326 2633 2332 2634
rect 2406 2638 2412 2639
rect 2406 2634 2407 2638
rect 2411 2634 2412 2638
rect 2406 2633 2412 2634
rect 2486 2638 2492 2639
rect 2486 2634 2487 2638
rect 2491 2634 2492 2638
rect 2486 2633 2492 2634
rect 2566 2638 2572 2639
rect 2566 2634 2567 2638
rect 2571 2634 2572 2638
rect 2566 2633 2572 2634
rect 2646 2638 2652 2639
rect 2646 2634 2647 2638
rect 2651 2634 2652 2638
rect 2646 2633 2652 2634
rect 2726 2638 2732 2639
rect 2726 2634 2727 2638
rect 2731 2634 2732 2638
rect 2726 2633 2732 2634
rect 2806 2638 2812 2639
rect 2806 2634 2807 2638
rect 2811 2634 2812 2638
rect 2806 2633 2812 2634
rect 2886 2638 2892 2639
rect 2886 2634 2887 2638
rect 2891 2634 2892 2638
rect 2886 2633 2892 2634
rect 2966 2638 2972 2639
rect 2966 2634 2967 2638
rect 2971 2634 2972 2638
rect 2966 2633 2972 2634
rect 2248 2615 2250 2633
rect 2328 2615 2330 2633
rect 2408 2615 2410 2633
rect 2488 2615 2490 2633
rect 2568 2615 2570 2633
rect 2648 2615 2650 2633
rect 2728 2615 2730 2633
rect 2808 2615 2810 2633
rect 2888 2615 2890 2633
rect 2968 2615 2970 2633
rect 3592 2615 3594 2651
rect 110 2610 116 2611
rect 134 2612 140 2613
rect 112 2587 114 2610
rect 134 2608 135 2612
rect 139 2608 140 2612
rect 134 2607 140 2608
rect 246 2612 252 2613
rect 246 2608 247 2612
rect 251 2608 252 2612
rect 246 2607 252 2608
rect 390 2612 396 2613
rect 390 2608 391 2612
rect 395 2608 396 2612
rect 390 2607 396 2608
rect 542 2612 548 2613
rect 542 2608 543 2612
rect 547 2608 548 2612
rect 542 2607 548 2608
rect 702 2612 708 2613
rect 702 2608 703 2612
rect 707 2608 708 2612
rect 702 2607 708 2608
rect 870 2612 876 2613
rect 870 2608 871 2612
rect 875 2608 876 2612
rect 870 2607 876 2608
rect 1038 2612 1044 2613
rect 1038 2608 1039 2612
rect 1043 2608 1044 2612
rect 1038 2607 1044 2608
rect 1206 2612 1212 2613
rect 1206 2608 1207 2612
rect 1211 2608 1212 2612
rect 1206 2607 1212 2608
rect 1382 2612 1388 2613
rect 1382 2608 1383 2612
rect 1387 2608 1388 2612
rect 1382 2607 1388 2608
rect 1558 2612 1564 2613
rect 1558 2608 1559 2612
rect 1563 2608 1564 2612
rect 1830 2611 1831 2615
rect 1835 2611 1836 2615
rect 1830 2610 1836 2611
rect 1871 2614 1875 2615
rect 1558 2607 1564 2608
rect 136 2587 138 2607
rect 248 2587 250 2607
rect 392 2587 394 2607
rect 544 2587 546 2607
rect 704 2587 706 2607
rect 872 2587 874 2607
rect 1040 2587 1042 2607
rect 1208 2587 1210 2607
rect 1384 2587 1386 2607
rect 1560 2587 1562 2607
rect 1832 2587 1834 2610
rect 1871 2609 1875 2610
rect 2191 2614 2195 2615
rect 2191 2609 2195 2610
rect 2247 2614 2251 2615
rect 2247 2609 2251 2610
rect 2271 2614 2275 2615
rect 2271 2609 2275 2610
rect 2327 2614 2331 2615
rect 2327 2609 2331 2610
rect 2351 2614 2355 2615
rect 2351 2609 2355 2610
rect 2407 2614 2411 2615
rect 2407 2609 2411 2610
rect 2431 2614 2435 2615
rect 2431 2609 2435 2610
rect 2487 2614 2491 2615
rect 2487 2609 2491 2610
rect 2511 2614 2515 2615
rect 2511 2609 2515 2610
rect 2567 2614 2571 2615
rect 2567 2609 2571 2610
rect 2591 2614 2595 2615
rect 2591 2609 2595 2610
rect 2647 2614 2651 2615
rect 2647 2609 2651 2610
rect 2671 2614 2675 2615
rect 2671 2609 2675 2610
rect 2727 2614 2731 2615
rect 2727 2609 2731 2610
rect 2751 2614 2755 2615
rect 2751 2609 2755 2610
rect 2807 2614 2811 2615
rect 2807 2609 2811 2610
rect 2831 2614 2835 2615
rect 2831 2609 2835 2610
rect 2887 2614 2891 2615
rect 2887 2609 2891 2610
rect 2911 2614 2915 2615
rect 2911 2609 2915 2610
rect 2967 2614 2971 2615
rect 2967 2609 2971 2610
rect 2991 2614 2995 2615
rect 2991 2609 2995 2610
rect 3591 2614 3595 2615
rect 3591 2609 3595 2610
rect 111 2586 115 2587
rect 111 2581 115 2582
rect 135 2586 139 2587
rect 135 2581 139 2582
rect 159 2586 163 2587
rect 159 2581 163 2582
rect 247 2586 251 2587
rect 247 2581 251 2582
rect 279 2586 283 2587
rect 279 2581 283 2582
rect 391 2586 395 2587
rect 391 2581 395 2582
rect 415 2586 419 2587
rect 415 2581 419 2582
rect 543 2586 547 2587
rect 543 2581 547 2582
rect 559 2586 563 2587
rect 559 2581 563 2582
rect 703 2586 707 2587
rect 703 2581 707 2582
rect 847 2586 851 2587
rect 847 2581 851 2582
rect 871 2586 875 2587
rect 871 2581 875 2582
rect 983 2586 987 2587
rect 983 2581 987 2582
rect 1039 2586 1043 2587
rect 1039 2581 1043 2582
rect 1119 2586 1123 2587
rect 1119 2581 1123 2582
rect 1207 2586 1211 2587
rect 1207 2581 1211 2582
rect 1255 2586 1259 2587
rect 1255 2581 1259 2582
rect 1383 2586 1387 2587
rect 1383 2581 1387 2582
rect 1391 2586 1395 2587
rect 1391 2581 1395 2582
rect 1527 2586 1531 2587
rect 1527 2581 1531 2582
rect 1559 2586 1563 2587
rect 1559 2581 1563 2582
rect 1831 2586 1835 2587
rect 1831 2581 1835 2582
rect 1872 2581 1874 2609
rect 2192 2599 2194 2609
rect 2272 2599 2274 2609
rect 2352 2599 2354 2609
rect 2432 2599 2434 2609
rect 2512 2599 2514 2609
rect 2592 2599 2594 2609
rect 2672 2599 2674 2609
rect 2752 2599 2754 2609
rect 2832 2599 2834 2609
rect 2912 2599 2914 2609
rect 2992 2599 2994 2609
rect 2190 2598 2196 2599
rect 2190 2594 2191 2598
rect 2195 2594 2196 2598
rect 2190 2593 2196 2594
rect 2270 2598 2276 2599
rect 2270 2594 2271 2598
rect 2275 2594 2276 2598
rect 2270 2593 2276 2594
rect 2350 2598 2356 2599
rect 2350 2594 2351 2598
rect 2355 2594 2356 2598
rect 2350 2593 2356 2594
rect 2430 2598 2436 2599
rect 2430 2594 2431 2598
rect 2435 2594 2436 2598
rect 2430 2593 2436 2594
rect 2510 2598 2516 2599
rect 2510 2594 2511 2598
rect 2515 2594 2516 2598
rect 2510 2593 2516 2594
rect 2590 2598 2596 2599
rect 2590 2594 2591 2598
rect 2595 2594 2596 2598
rect 2590 2593 2596 2594
rect 2670 2598 2676 2599
rect 2670 2594 2671 2598
rect 2675 2594 2676 2598
rect 2670 2593 2676 2594
rect 2750 2598 2756 2599
rect 2750 2594 2751 2598
rect 2755 2594 2756 2598
rect 2750 2593 2756 2594
rect 2830 2598 2836 2599
rect 2830 2594 2831 2598
rect 2835 2594 2836 2598
rect 2830 2593 2836 2594
rect 2910 2598 2916 2599
rect 2910 2594 2911 2598
rect 2915 2594 2916 2598
rect 2910 2593 2916 2594
rect 2990 2598 2996 2599
rect 2990 2594 2991 2598
rect 2995 2594 2996 2598
rect 2990 2593 2996 2594
rect 3592 2581 3594 2609
rect 112 2562 114 2581
rect 160 2565 162 2581
rect 280 2565 282 2581
rect 416 2565 418 2581
rect 560 2565 562 2581
rect 704 2565 706 2581
rect 848 2565 850 2581
rect 984 2565 986 2581
rect 1120 2565 1122 2581
rect 1256 2565 1258 2581
rect 1392 2565 1394 2581
rect 1528 2565 1530 2581
rect 158 2564 164 2565
rect 110 2561 116 2562
rect 110 2557 111 2561
rect 115 2557 116 2561
rect 158 2560 159 2564
rect 163 2560 164 2564
rect 158 2559 164 2560
rect 278 2564 284 2565
rect 278 2560 279 2564
rect 283 2560 284 2564
rect 278 2559 284 2560
rect 414 2564 420 2565
rect 414 2560 415 2564
rect 419 2560 420 2564
rect 414 2559 420 2560
rect 558 2564 564 2565
rect 558 2560 559 2564
rect 563 2560 564 2564
rect 558 2559 564 2560
rect 702 2564 708 2565
rect 702 2560 703 2564
rect 707 2560 708 2564
rect 702 2559 708 2560
rect 846 2564 852 2565
rect 846 2560 847 2564
rect 851 2560 852 2564
rect 846 2559 852 2560
rect 982 2564 988 2565
rect 982 2560 983 2564
rect 987 2560 988 2564
rect 982 2559 988 2560
rect 1118 2564 1124 2565
rect 1118 2560 1119 2564
rect 1123 2560 1124 2564
rect 1118 2559 1124 2560
rect 1254 2564 1260 2565
rect 1254 2560 1255 2564
rect 1259 2560 1260 2564
rect 1254 2559 1260 2560
rect 1390 2564 1396 2565
rect 1390 2560 1391 2564
rect 1395 2560 1396 2564
rect 1390 2559 1396 2560
rect 1526 2564 1532 2565
rect 1526 2560 1527 2564
rect 1531 2560 1532 2564
rect 1832 2562 1834 2581
rect 1870 2580 1876 2581
rect 1870 2576 1871 2580
rect 1875 2576 1876 2580
rect 1870 2575 1876 2576
rect 3590 2580 3596 2581
rect 3590 2576 3591 2580
rect 3595 2576 3596 2580
rect 3590 2575 3596 2576
rect 1870 2563 1876 2564
rect 1526 2559 1532 2560
rect 1830 2561 1836 2562
rect 110 2556 116 2557
rect 1830 2557 1831 2561
rect 1835 2557 1836 2561
rect 1870 2559 1871 2563
rect 1875 2559 1876 2563
rect 3590 2563 3596 2564
rect 1870 2558 1876 2559
rect 2182 2560 2188 2561
rect 1830 2556 1836 2557
rect 110 2544 116 2545
rect 110 2540 111 2544
rect 115 2540 116 2544
rect 110 2539 116 2540
rect 1830 2544 1836 2545
rect 1830 2540 1831 2544
rect 1835 2540 1836 2544
rect 1830 2539 1836 2540
rect 112 2507 114 2539
rect 166 2526 172 2527
rect 166 2522 167 2526
rect 171 2522 172 2526
rect 166 2521 172 2522
rect 286 2526 292 2527
rect 286 2522 287 2526
rect 291 2522 292 2526
rect 286 2521 292 2522
rect 422 2526 428 2527
rect 422 2522 423 2526
rect 427 2522 428 2526
rect 422 2521 428 2522
rect 566 2526 572 2527
rect 566 2522 567 2526
rect 571 2522 572 2526
rect 566 2521 572 2522
rect 710 2526 716 2527
rect 710 2522 711 2526
rect 715 2522 716 2526
rect 710 2521 716 2522
rect 854 2526 860 2527
rect 854 2522 855 2526
rect 859 2522 860 2526
rect 854 2521 860 2522
rect 990 2526 996 2527
rect 990 2522 991 2526
rect 995 2522 996 2526
rect 990 2521 996 2522
rect 1126 2526 1132 2527
rect 1126 2522 1127 2526
rect 1131 2522 1132 2526
rect 1126 2521 1132 2522
rect 1262 2526 1268 2527
rect 1262 2522 1263 2526
rect 1267 2522 1268 2526
rect 1262 2521 1268 2522
rect 1398 2526 1404 2527
rect 1398 2522 1399 2526
rect 1403 2522 1404 2526
rect 1398 2521 1404 2522
rect 1534 2526 1540 2527
rect 1534 2522 1535 2526
rect 1539 2522 1540 2526
rect 1534 2521 1540 2522
rect 168 2507 170 2521
rect 288 2507 290 2521
rect 424 2507 426 2521
rect 568 2507 570 2521
rect 712 2507 714 2521
rect 856 2507 858 2521
rect 992 2507 994 2521
rect 1128 2507 1130 2521
rect 1264 2507 1266 2521
rect 1400 2507 1402 2521
rect 1536 2507 1538 2521
rect 1832 2507 1834 2539
rect 1872 2531 1874 2558
rect 2182 2556 2183 2560
rect 2187 2556 2188 2560
rect 2182 2555 2188 2556
rect 2262 2560 2268 2561
rect 2262 2556 2263 2560
rect 2267 2556 2268 2560
rect 2262 2555 2268 2556
rect 2342 2560 2348 2561
rect 2342 2556 2343 2560
rect 2347 2556 2348 2560
rect 2342 2555 2348 2556
rect 2422 2560 2428 2561
rect 2422 2556 2423 2560
rect 2427 2556 2428 2560
rect 2422 2555 2428 2556
rect 2502 2560 2508 2561
rect 2502 2556 2503 2560
rect 2507 2556 2508 2560
rect 2502 2555 2508 2556
rect 2582 2560 2588 2561
rect 2582 2556 2583 2560
rect 2587 2556 2588 2560
rect 2582 2555 2588 2556
rect 2662 2560 2668 2561
rect 2662 2556 2663 2560
rect 2667 2556 2668 2560
rect 2662 2555 2668 2556
rect 2742 2560 2748 2561
rect 2742 2556 2743 2560
rect 2747 2556 2748 2560
rect 2742 2555 2748 2556
rect 2822 2560 2828 2561
rect 2822 2556 2823 2560
rect 2827 2556 2828 2560
rect 2822 2555 2828 2556
rect 2902 2560 2908 2561
rect 2902 2556 2903 2560
rect 2907 2556 2908 2560
rect 2902 2555 2908 2556
rect 2982 2560 2988 2561
rect 2982 2556 2983 2560
rect 2987 2556 2988 2560
rect 3590 2559 3591 2563
rect 3595 2559 3596 2563
rect 3590 2558 3596 2559
rect 2982 2555 2988 2556
rect 2184 2531 2186 2555
rect 2264 2531 2266 2555
rect 2344 2531 2346 2555
rect 2424 2531 2426 2555
rect 2504 2531 2506 2555
rect 2584 2531 2586 2555
rect 2664 2531 2666 2555
rect 2744 2531 2746 2555
rect 2824 2531 2826 2555
rect 2904 2531 2906 2555
rect 2984 2531 2986 2555
rect 3592 2531 3594 2558
rect 1871 2530 1875 2531
rect 1871 2525 1875 2526
rect 2119 2530 2123 2531
rect 2119 2525 2123 2526
rect 2183 2530 2187 2531
rect 2183 2525 2187 2526
rect 2207 2530 2211 2531
rect 2207 2525 2211 2526
rect 2263 2530 2267 2531
rect 2263 2525 2267 2526
rect 2303 2530 2307 2531
rect 2303 2525 2307 2526
rect 2343 2530 2347 2531
rect 2343 2525 2347 2526
rect 2399 2530 2403 2531
rect 2399 2525 2403 2526
rect 2423 2530 2427 2531
rect 2423 2525 2427 2526
rect 2495 2530 2499 2531
rect 2495 2525 2499 2526
rect 2503 2530 2507 2531
rect 2503 2525 2507 2526
rect 2583 2530 2587 2531
rect 2583 2525 2587 2526
rect 2591 2530 2595 2531
rect 2591 2525 2595 2526
rect 2663 2530 2667 2531
rect 2663 2525 2667 2526
rect 2687 2530 2691 2531
rect 2687 2525 2691 2526
rect 2743 2530 2747 2531
rect 2743 2525 2747 2526
rect 2783 2530 2787 2531
rect 2783 2525 2787 2526
rect 2823 2530 2827 2531
rect 2823 2525 2827 2526
rect 2879 2530 2883 2531
rect 2879 2525 2883 2526
rect 2903 2530 2907 2531
rect 2903 2525 2907 2526
rect 2975 2530 2979 2531
rect 2975 2525 2979 2526
rect 2983 2530 2987 2531
rect 2983 2525 2987 2526
rect 3079 2530 3083 2531
rect 3079 2525 3083 2526
rect 3591 2530 3595 2531
rect 3591 2525 3595 2526
rect 111 2506 115 2507
rect 111 2501 115 2502
rect 167 2506 171 2507
rect 167 2501 171 2502
rect 287 2506 291 2507
rect 287 2501 291 2502
rect 335 2506 339 2507
rect 335 2501 339 2502
rect 415 2506 419 2507
rect 415 2501 419 2502
rect 423 2506 427 2507
rect 423 2501 427 2502
rect 503 2506 507 2507
rect 503 2501 507 2502
rect 567 2506 571 2507
rect 567 2501 571 2502
rect 599 2506 603 2507
rect 599 2501 603 2502
rect 703 2506 707 2507
rect 703 2501 707 2502
rect 711 2506 715 2507
rect 711 2501 715 2502
rect 815 2506 819 2507
rect 815 2501 819 2502
rect 855 2506 859 2507
rect 855 2501 859 2502
rect 935 2506 939 2507
rect 935 2501 939 2502
rect 991 2506 995 2507
rect 991 2501 995 2502
rect 1063 2506 1067 2507
rect 1063 2501 1067 2502
rect 1127 2506 1131 2507
rect 1127 2501 1131 2502
rect 1191 2506 1195 2507
rect 1191 2501 1195 2502
rect 1263 2506 1267 2507
rect 1263 2501 1267 2502
rect 1327 2506 1331 2507
rect 1327 2501 1331 2502
rect 1399 2506 1403 2507
rect 1399 2501 1403 2502
rect 1471 2506 1475 2507
rect 1471 2501 1475 2502
rect 1535 2506 1539 2507
rect 1535 2501 1539 2502
rect 1831 2506 1835 2507
rect 1872 2506 1874 2525
rect 2120 2509 2122 2525
rect 2208 2509 2210 2525
rect 2304 2509 2306 2525
rect 2400 2509 2402 2525
rect 2496 2509 2498 2525
rect 2592 2509 2594 2525
rect 2688 2509 2690 2525
rect 2784 2509 2786 2525
rect 2880 2509 2882 2525
rect 2976 2509 2978 2525
rect 3080 2509 3082 2525
rect 2118 2508 2124 2509
rect 1831 2501 1835 2502
rect 1870 2505 1876 2506
rect 1870 2501 1871 2505
rect 1875 2501 1876 2505
rect 2118 2504 2119 2508
rect 2123 2504 2124 2508
rect 2118 2503 2124 2504
rect 2206 2508 2212 2509
rect 2206 2504 2207 2508
rect 2211 2504 2212 2508
rect 2206 2503 2212 2504
rect 2302 2508 2308 2509
rect 2302 2504 2303 2508
rect 2307 2504 2308 2508
rect 2302 2503 2308 2504
rect 2398 2508 2404 2509
rect 2398 2504 2399 2508
rect 2403 2504 2404 2508
rect 2398 2503 2404 2504
rect 2494 2508 2500 2509
rect 2494 2504 2495 2508
rect 2499 2504 2500 2508
rect 2494 2503 2500 2504
rect 2590 2508 2596 2509
rect 2590 2504 2591 2508
rect 2595 2504 2596 2508
rect 2590 2503 2596 2504
rect 2686 2508 2692 2509
rect 2686 2504 2687 2508
rect 2691 2504 2692 2508
rect 2686 2503 2692 2504
rect 2782 2508 2788 2509
rect 2782 2504 2783 2508
rect 2787 2504 2788 2508
rect 2782 2503 2788 2504
rect 2878 2508 2884 2509
rect 2878 2504 2879 2508
rect 2883 2504 2884 2508
rect 2878 2503 2884 2504
rect 2974 2508 2980 2509
rect 2974 2504 2975 2508
rect 2979 2504 2980 2508
rect 2974 2503 2980 2504
rect 3078 2508 3084 2509
rect 3078 2504 3079 2508
rect 3083 2504 3084 2508
rect 3592 2506 3594 2525
rect 3078 2503 3084 2504
rect 3590 2505 3596 2506
rect 112 2473 114 2501
rect 336 2491 338 2501
rect 416 2491 418 2501
rect 504 2491 506 2501
rect 600 2491 602 2501
rect 704 2491 706 2501
rect 816 2491 818 2501
rect 936 2491 938 2501
rect 1064 2491 1066 2501
rect 1192 2491 1194 2501
rect 1328 2491 1330 2501
rect 1472 2491 1474 2501
rect 334 2490 340 2491
rect 334 2486 335 2490
rect 339 2486 340 2490
rect 334 2485 340 2486
rect 414 2490 420 2491
rect 414 2486 415 2490
rect 419 2486 420 2490
rect 414 2485 420 2486
rect 502 2490 508 2491
rect 502 2486 503 2490
rect 507 2486 508 2490
rect 502 2485 508 2486
rect 598 2490 604 2491
rect 598 2486 599 2490
rect 603 2486 604 2490
rect 598 2485 604 2486
rect 702 2490 708 2491
rect 702 2486 703 2490
rect 707 2486 708 2490
rect 702 2485 708 2486
rect 814 2490 820 2491
rect 814 2486 815 2490
rect 819 2486 820 2490
rect 814 2485 820 2486
rect 934 2490 940 2491
rect 934 2486 935 2490
rect 939 2486 940 2490
rect 934 2485 940 2486
rect 1062 2490 1068 2491
rect 1062 2486 1063 2490
rect 1067 2486 1068 2490
rect 1062 2485 1068 2486
rect 1190 2490 1196 2491
rect 1190 2486 1191 2490
rect 1195 2486 1196 2490
rect 1190 2485 1196 2486
rect 1326 2490 1332 2491
rect 1326 2486 1327 2490
rect 1331 2486 1332 2490
rect 1326 2485 1332 2486
rect 1470 2490 1476 2491
rect 1470 2486 1471 2490
rect 1475 2486 1476 2490
rect 1470 2485 1476 2486
rect 1832 2473 1834 2501
rect 1870 2500 1876 2501
rect 3590 2501 3591 2505
rect 3595 2501 3596 2505
rect 3590 2500 3596 2501
rect 1870 2488 1876 2489
rect 1870 2484 1871 2488
rect 1875 2484 1876 2488
rect 1870 2483 1876 2484
rect 3590 2488 3596 2489
rect 3590 2484 3591 2488
rect 3595 2484 3596 2488
rect 3590 2483 3596 2484
rect 110 2472 116 2473
rect 110 2468 111 2472
rect 115 2468 116 2472
rect 110 2467 116 2468
rect 1830 2472 1836 2473
rect 1830 2468 1831 2472
rect 1835 2468 1836 2472
rect 1830 2467 1836 2468
rect 110 2455 116 2456
rect 110 2451 111 2455
rect 115 2451 116 2455
rect 1830 2455 1836 2456
rect 110 2450 116 2451
rect 326 2452 332 2453
rect 112 2423 114 2450
rect 326 2448 327 2452
rect 331 2448 332 2452
rect 326 2447 332 2448
rect 406 2452 412 2453
rect 406 2448 407 2452
rect 411 2448 412 2452
rect 406 2447 412 2448
rect 494 2452 500 2453
rect 494 2448 495 2452
rect 499 2448 500 2452
rect 494 2447 500 2448
rect 590 2452 596 2453
rect 590 2448 591 2452
rect 595 2448 596 2452
rect 590 2447 596 2448
rect 694 2452 700 2453
rect 694 2448 695 2452
rect 699 2448 700 2452
rect 694 2447 700 2448
rect 806 2452 812 2453
rect 806 2448 807 2452
rect 811 2448 812 2452
rect 806 2447 812 2448
rect 926 2452 932 2453
rect 926 2448 927 2452
rect 931 2448 932 2452
rect 926 2447 932 2448
rect 1054 2452 1060 2453
rect 1054 2448 1055 2452
rect 1059 2448 1060 2452
rect 1054 2447 1060 2448
rect 1182 2452 1188 2453
rect 1182 2448 1183 2452
rect 1187 2448 1188 2452
rect 1182 2447 1188 2448
rect 1318 2452 1324 2453
rect 1318 2448 1319 2452
rect 1323 2448 1324 2452
rect 1318 2447 1324 2448
rect 1462 2452 1468 2453
rect 1462 2448 1463 2452
rect 1467 2448 1468 2452
rect 1830 2451 1831 2455
rect 1835 2451 1836 2455
rect 1872 2451 1874 2483
rect 2126 2470 2132 2471
rect 2126 2466 2127 2470
rect 2131 2466 2132 2470
rect 2126 2465 2132 2466
rect 2214 2470 2220 2471
rect 2214 2466 2215 2470
rect 2219 2466 2220 2470
rect 2214 2465 2220 2466
rect 2310 2470 2316 2471
rect 2310 2466 2311 2470
rect 2315 2466 2316 2470
rect 2310 2465 2316 2466
rect 2406 2470 2412 2471
rect 2406 2466 2407 2470
rect 2411 2466 2412 2470
rect 2406 2465 2412 2466
rect 2502 2470 2508 2471
rect 2502 2466 2503 2470
rect 2507 2466 2508 2470
rect 2502 2465 2508 2466
rect 2598 2470 2604 2471
rect 2598 2466 2599 2470
rect 2603 2466 2604 2470
rect 2598 2465 2604 2466
rect 2694 2470 2700 2471
rect 2694 2466 2695 2470
rect 2699 2466 2700 2470
rect 2694 2465 2700 2466
rect 2790 2470 2796 2471
rect 2790 2466 2791 2470
rect 2795 2466 2796 2470
rect 2790 2465 2796 2466
rect 2886 2470 2892 2471
rect 2886 2466 2887 2470
rect 2891 2466 2892 2470
rect 2886 2465 2892 2466
rect 2982 2470 2988 2471
rect 2982 2466 2983 2470
rect 2987 2466 2988 2470
rect 2982 2465 2988 2466
rect 3086 2470 3092 2471
rect 3086 2466 3087 2470
rect 3091 2466 3092 2470
rect 3086 2465 3092 2466
rect 2128 2451 2130 2465
rect 2216 2451 2218 2465
rect 2312 2451 2314 2465
rect 2408 2451 2410 2465
rect 2504 2451 2506 2465
rect 2600 2451 2602 2465
rect 2696 2451 2698 2465
rect 2792 2451 2794 2465
rect 2888 2451 2890 2465
rect 2984 2451 2986 2465
rect 3088 2451 3090 2465
rect 3592 2451 3594 2483
rect 1830 2450 1836 2451
rect 1871 2450 1875 2451
rect 1462 2447 1468 2448
rect 328 2423 330 2447
rect 408 2423 410 2447
rect 496 2423 498 2447
rect 592 2423 594 2447
rect 696 2423 698 2447
rect 808 2423 810 2447
rect 928 2423 930 2447
rect 1056 2423 1058 2447
rect 1184 2423 1186 2447
rect 1320 2423 1322 2447
rect 1464 2423 1466 2447
rect 1832 2423 1834 2450
rect 1871 2445 1875 2446
rect 1903 2450 1907 2451
rect 1903 2445 1907 2446
rect 1991 2450 1995 2451
rect 1991 2445 1995 2446
rect 2111 2450 2115 2451
rect 2111 2445 2115 2446
rect 2127 2450 2131 2451
rect 2127 2445 2131 2446
rect 2215 2450 2219 2451
rect 2215 2445 2219 2446
rect 2247 2450 2251 2451
rect 2247 2445 2251 2446
rect 2311 2450 2315 2451
rect 2311 2445 2315 2446
rect 2391 2450 2395 2451
rect 2391 2445 2395 2446
rect 2407 2450 2411 2451
rect 2407 2445 2411 2446
rect 2503 2450 2507 2451
rect 2503 2445 2507 2446
rect 2535 2450 2539 2451
rect 2535 2445 2539 2446
rect 2599 2450 2603 2451
rect 2599 2445 2603 2446
rect 2671 2450 2675 2451
rect 2671 2445 2675 2446
rect 2695 2450 2699 2451
rect 2695 2445 2699 2446
rect 2791 2450 2795 2451
rect 2791 2445 2795 2446
rect 2807 2450 2811 2451
rect 2807 2445 2811 2446
rect 2887 2450 2891 2451
rect 2887 2445 2891 2446
rect 2943 2450 2947 2451
rect 2943 2445 2947 2446
rect 2983 2450 2987 2451
rect 2983 2445 2987 2446
rect 3079 2450 3083 2451
rect 3079 2445 3083 2446
rect 3087 2450 3091 2451
rect 3087 2445 3091 2446
rect 3215 2450 3219 2451
rect 3215 2445 3219 2446
rect 3591 2450 3595 2451
rect 3591 2445 3595 2446
rect 111 2422 115 2423
rect 111 2417 115 2418
rect 327 2422 331 2423
rect 327 2417 331 2418
rect 383 2422 387 2423
rect 383 2417 387 2418
rect 407 2422 411 2423
rect 407 2417 411 2418
rect 463 2422 467 2423
rect 463 2417 467 2418
rect 495 2422 499 2423
rect 495 2417 499 2418
rect 543 2422 547 2423
rect 543 2417 547 2418
rect 591 2422 595 2423
rect 591 2417 595 2418
rect 623 2422 627 2423
rect 623 2417 627 2418
rect 695 2422 699 2423
rect 695 2417 699 2418
rect 703 2422 707 2423
rect 703 2417 707 2418
rect 783 2422 787 2423
rect 783 2417 787 2418
rect 807 2422 811 2423
rect 807 2417 811 2418
rect 863 2422 867 2423
rect 863 2417 867 2418
rect 927 2422 931 2423
rect 927 2417 931 2418
rect 943 2422 947 2423
rect 943 2417 947 2418
rect 1023 2422 1027 2423
rect 1023 2417 1027 2418
rect 1055 2422 1059 2423
rect 1055 2417 1059 2418
rect 1103 2422 1107 2423
rect 1103 2417 1107 2418
rect 1183 2422 1187 2423
rect 1183 2417 1187 2418
rect 1263 2422 1267 2423
rect 1263 2417 1267 2418
rect 1319 2422 1323 2423
rect 1319 2417 1323 2418
rect 1351 2422 1355 2423
rect 1351 2417 1355 2418
rect 1439 2422 1443 2423
rect 1439 2417 1443 2418
rect 1463 2422 1467 2423
rect 1463 2417 1467 2418
rect 1527 2422 1531 2423
rect 1527 2417 1531 2418
rect 1831 2422 1835 2423
rect 1831 2417 1835 2418
rect 1872 2417 1874 2445
rect 1904 2435 1906 2445
rect 1992 2435 1994 2445
rect 2112 2435 2114 2445
rect 2248 2435 2250 2445
rect 2392 2435 2394 2445
rect 2536 2435 2538 2445
rect 2672 2435 2674 2445
rect 2808 2435 2810 2445
rect 2944 2435 2946 2445
rect 3080 2435 3082 2445
rect 3216 2435 3218 2445
rect 1902 2434 1908 2435
rect 1902 2430 1903 2434
rect 1907 2430 1908 2434
rect 1902 2429 1908 2430
rect 1990 2434 1996 2435
rect 1990 2430 1991 2434
rect 1995 2430 1996 2434
rect 1990 2429 1996 2430
rect 2110 2434 2116 2435
rect 2110 2430 2111 2434
rect 2115 2430 2116 2434
rect 2110 2429 2116 2430
rect 2246 2434 2252 2435
rect 2246 2430 2247 2434
rect 2251 2430 2252 2434
rect 2246 2429 2252 2430
rect 2390 2434 2396 2435
rect 2390 2430 2391 2434
rect 2395 2430 2396 2434
rect 2390 2429 2396 2430
rect 2534 2434 2540 2435
rect 2534 2430 2535 2434
rect 2539 2430 2540 2434
rect 2534 2429 2540 2430
rect 2670 2434 2676 2435
rect 2670 2430 2671 2434
rect 2675 2430 2676 2434
rect 2670 2429 2676 2430
rect 2806 2434 2812 2435
rect 2806 2430 2807 2434
rect 2811 2430 2812 2434
rect 2806 2429 2812 2430
rect 2942 2434 2948 2435
rect 2942 2430 2943 2434
rect 2947 2430 2948 2434
rect 2942 2429 2948 2430
rect 3078 2434 3084 2435
rect 3078 2430 3079 2434
rect 3083 2430 3084 2434
rect 3078 2429 3084 2430
rect 3214 2434 3220 2435
rect 3214 2430 3215 2434
rect 3219 2430 3220 2434
rect 3214 2429 3220 2430
rect 3592 2417 3594 2445
rect 112 2398 114 2417
rect 384 2401 386 2417
rect 464 2401 466 2417
rect 544 2401 546 2417
rect 624 2401 626 2417
rect 704 2401 706 2417
rect 784 2401 786 2417
rect 864 2401 866 2417
rect 944 2401 946 2417
rect 1024 2401 1026 2417
rect 1104 2401 1106 2417
rect 1184 2401 1186 2417
rect 1264 2401 1266 2417
rect 1352 2401 1354 2417
rect 1440 2401 1442 2417
rect 1528 2401 1530 2417
rect 382 2400 388 2401
rect 110 2397 116 2398
rect 110 2393 111 2397
rect 115 2393 116 2397
rect 382 2396 383 2400
rect 387 2396 388 2400
rect 382 2395 388 2396
rect 462 2400 468 2401
rect 462 2396 463 2400
rect 467 2396 468 2400
rect 462 2395 468 2396
rect 542 2400 548 2401
rect 542 2396 543 2400
rect 547 2396 548 2400
rect 542 2395 548 2396
rect 622 2400 628 2401
rect 622 2396 623 2400
rect 627 2396 628 2400
rect 622 2395 628 2396
rect 702 2400 708 2401
rect 702 2396 703 2400
rect 707 2396 708 2400
rect 702 2395 708 2396
rect 782 2400 788 2401
rect 782 2396 783 2400
rect 787 2396 788 2400
rect 782 2395 788 2396
rect 862 2400 868 2401
rect 862 2396 863 2400
rect 867 2396 868 2400
rect 862 2395 868 2396
rect 942 2400 948 2401
rect 942 2396 943 2400
rect 947 2396 948 2400
rect 942 2395 948 2396
rect 1022 2400 1028 2401
rect 1022 2396 1023 2400
rect 1027 2396 1028 2400
rect 1022 2395 1028 2396
rect 1102 2400 1108 2401
rect 1102 2396 1103 2400
rect 1107 2396 1108 2400
rect 1102 2395 1108 2396
rect 1182 2400 1188 2401
rect 1182 2396 1183 2400
rect 1187 2396 1188 2400
rect 1182 2395 1188 2396
rect 1262 2400 1268 2401
rect 1262 2396 1263 2400
rect 1267 2396 1268 2400
rect 1262 2395 1268 2396
rect 1350 2400 1356 2401
rect 1350 2396 1351 2400
rect 1355 2396 1356 2400
rect 1350 2395 1356 2396
rect 1438 2400 1444 2401
rect 1438 2396 1439 2400
rect 1443 2396 1444 2400
rect 1438 2395 1444 2396
rect 1526 2400 1532 2401
rect 1526 2396 1527 2400
rect 1531 2396 1532 2400
rect 1832 2398 1834 2417
rect 1870 2416 1876 2417
rect 1870 2412 1871 2416
rect 1875 2412 1876 2416
rect 1870 2411 1876 2412
rect 3590 2416 3596 2417
rect 3590 2412 3591 2416
rect 3595 2412 3596 2416
rect 3590 2411 3596 2412
rect 1870 2399 1876 2400
rect 1526 2395 1532 2396
rect 1830 2397 1836 2398
rect 110 2392 116 2393
rect 1830 2393 1831 2397
rect 1835 2393 1836 2397
rect 1870 2395 1871 2399
rect 1875 2395 1876 2399
rect 3590 2399 3596 2400
rect 1870 2394 1876 2395
rect 1894 2396 1900 2397
rect 1830 2392 1836 2393
rect 110 2380 116 2381
rect 110 2376 111 2380
rect 115 2376 116 2380
rect 110 2375 116 2376
rect 1830 2380 1836 2381
rect 1830 2376 1831 2380
rect 1835 2376 1836 2380
rect 1830 2375 1836 2376
rect 112 2347 114 2375
rect 390 2362 396 2363
rect 390 2358 391 2362
rect 395 2358 396 2362
rect 390 2357 396 2358
rect 470 2362 476 2363
rect 470 2358 471 2362
rect 475 2358 476 2362
rect 470 2357 476 2358
rect 550 2362 556 2363
rect 550 2358 551 2362
rect 555 2358 556 2362
rect 550 2357 556 2358
rect 630 2362 636 2363
rect 630 2358 631 2362
rect 635 2358 636 2362
rect 630 2357 636 2358
rect 710 2362 716 2363
rect 710 2358 711 2362
rect 715 2358 716 2362
rect 710 2357 716 2358
rect 790 2362 796 2363
rect 790 2358 791 2362
rect 795 2358 796 2362
rect 790 2357 796 2358
rect 870 2362 876 2363
rect 870 2358 871 2362
rect 875 2358 876 2362
rect 870 2357 876 2358
rect 950 2362 956 2363
rect 950 2358 951 2362
rect 955 2358 956 2362
rect 950 2357 956 2358
rect 1030 2362 1036 2363
rect 1030 2358 1031 2362
rect 1035 2358 1036 2362
rect 1030 2357 1036 2358
rect 1110 2362 1116 2363
rect 1110 2358 1111 2362
rect 1115 2358 1116 2362
rect 1110 2357 1116 2358
rect 1190 2362 1196 2363
rect 1190 2358 1191 2362
rect 1195 2358 1196 2362
rect 1190 2357 1196 2358
rect 1270 2362 1276 2363
rect 1270 2358 1271 2362
rect 1275 2358 1276 2362
rect 1270 2357 1276 2358
rect 1358 2362 1364 2363
rect 1358 2358 1359 2362
rect 1363 2358 1364 2362
rect 1358 2357 1364 2358
rect 1446 2362 1452 2363
rect 1446 2358 1447 2362
rect 1451 2358 1452 2362
rect 1446 2357 1452 2358
rect 1534 2362 1540 2363
rect 1534 2358 1535 2362
rect 1539 2358 1540 2362
rect 1534 2357 1540 2358
rect 392 2347 394 2357
rect 472 2347 474 2357
rect 552 2347 554 2357
rect 632 2347 634 2357
rect 712 2347 714 2357
rect 792 2347 794 2357
rect 872 2347 874 2357
rect 952 2347 954 2357
rect 1032 2347 1034 2357
rect 1112 2347 1114 2357
rect 1192 2347 1194 2357
rect 1272 2347 1274 2357
rect 1360 2347 1362 2357
rect 1448 2347 1450 2357
rect 1536 2347 1538 2357
rect 1832 2347 1834 2375
rect 1872 2367 1874 2394
rect 1894 2392 1895 2396
rect 1899 2392 1900 2396
rect 1894 2391 1900 2392
rect 1982 2396 1988 2397
rect 1982 2392 1983 2396
rect 1987 2392 1988 2396
rect 1982 2391 1988 2392
rect 2102 2396 2108 2397
rect 2102 2392 2103 2396
rect 2107 2392 2108 2396
rect 2102 2391 2108 2392
rect 2238 2396 2244 2397
rect 2238 2392 2239 2396
rect 2243 2392 2244 2396
rect 2238 2391 2244 2392
rect 2382 2396 2388 2397
rect 2382 2392 2383 2396
rect 2387 2392 2388 2396
rect 2382 2391 2388 2392
rect 2526 2396 2532 2397
rect 2526 2392 2527 2396
rect 2531 2392 2532 2396
rect 2526 2391 2532 2392
rect 2662 2396 2668 2397
rect 2662 2392 2663 2396
rect 2667 2392 2668 2396
rect 2662 2391 2668 2392
rect 2798 2396 2804 2397
rect 2798 2392 2799 2396
rect 2803 2392 2804 2396
rect 2798 2391 2804 2392
rect 2934 2396 2940 2397
rect 2934 2392 2935 2396
rect 2939 2392 2940 2396
rect 2934 2391 2940 2392
rect 3070 2396 3076 2397
rect 3070 2392 3071 2396
rect 3075 2392 3076 2396
rect 3070 2391 3076 2392
rect 3206 2396 3212 2397
rect 3206 2392 3207 2396
rect 3211 2392 3212 2396
rect 3590 2395 3591 2399
rect 3595 2395 3596 2399
rect 3590 2394 3596 2395
rect 3206 2391 3212 2392
rect 1896 2367 1898 2391
rect 1984 2367 1986 2391
rect 2104 2367 2106 2391
rect 2240 2367 2242 2391
rect 2384 2367 2386 2391
rect 2528 2367 2530 2391
rect 2664 2367 2666 2391
rect 2800 2367 2802 2391
rect 2936 2367 2938 2391
rect 3072 2367 3074 2391
rect 3208 2367 3210 2391
rect 3592 2367 3594 2394
rect 1871 2366 1875 2367
rect 1871 2361 1875 2362
rect 1895 2366 1899 2367
rect 1895 2361 1899 2362
rect 1983 2366 1987 2367
rect 1983 2361 1987 2362
rect 2015 2366 2019 2367
rect 2015 2361 2019 2362
rect 2103 2366 2107 2367
rect 2103 2361 2107 2362
rect 2175 2366 2179 2367
rect 2175 2361 2179 2362
rect 2239 2366 2243 2367
rect 2239 2361 2243 2362
rect 2343 2366 2347 2367
rect 2343 2361 2347 2362
rect 2383 2366 2387 2367
rect 2383 2361 2387 2362
rect 2511 2366 2515 2367
rect 2511 2361 2515 2362
rect 2527 2366 2531 2367
rect 2527 2361 2531 2362
rect 2663 2366 2667 2367
rect 2663 2361 2667 2362
rect 2671 2366 2675 2367
rect 2671 2361 2675 2362
rect 2799 2366 2803 2367
rect 2799 2361 2803 2362
rect 2823 2366 2827 2367
rect 2823 2361 2827 2362
rect 2935 2366 2939 2367
rect 2935 2361 2939 2362
rect 2959 2366 2963 2367
rect 2959 2361 2963 2362
rect 3071 2366 3075 2367
rect 3071 2361 3075 2362
rect 3079 2366 3083 2367
rect 3079 2361 3083 2362
rect 3191 2366 3195 2367
rect 3191 2361 3195 2362
rect 3207 2366 3211 2367
rect 3207 2361 3211 2362
rect 3303 2366 3307 2367
rect 3303 2361 3307 2362
rect 3415 2366 3419 2367
rect 3415 2361 3419 2362
rect 3503 2366 3507 2367
rect 3503 2361 3507 2362
rect 3591 2366 3595 2367
rect 3591 2361 3595 2362
rect 111 2346 115 2347
rect 111 2341 115 2342
rect 391 2346 395 2347
rect 391 2341 395 2342
rect 471 2346 475 2347
rect 471 2341 475 2342
rect 551 2346 555 2347
rect 551 2341 555 2342
rect 631 2346 635 2347
rect 631 2341 635 2342
rect 711 2346 715 2347
rect 711 2341 715 2342
rect 791 2346 795 2347
rect 791 2341 795 2342
rect 871 2346 875 2347
rect 871 2341 875 2342
rect 951 2346 955 2347
rect 951 2341 955 2342
rect 1031 2346 1035 2347
rect 1031 2341 1035 2342
rect 1111 2346 1115 2347
rect 1111 2341 1115 2342
rect 1191 2346 1195 2347
rect 1191 2341 1195 2342
rect 1271 2346 1275 2347
rect 1271 2341 1275 2342
rect 1359 2346 1363 2347
rect 1359 2341 1363 2342
rect 1407 2346 1411 2347
rect 1407 2341 1411 2342
rect 1447 2346 1451 2347
rect 1447 2341 1451 2342
rect 1487 2346 1491 2347
rect 1487 2341 1491 2342
rect 1535 2346 1539 2347
rect 1535 2341 1539 2342
rect 1567 2346 1571 2347
rect 1567 2341 1571 2342
rect 1647 2346 1651 2347
rect 1647 2341 1651 2342
rect 1831 2346 1835 2347
rect 1872 2342 1874 2361
rect 1896 2345 1898 2361
rect 2016 2345 2018 2361
rect 2176 2345 2178 2361
rect 2344 2345 2346 2361
rect 2512 2345 2514 2361
rect 2672 2345 2674 2361
rect 2824 2345 2826 2361
rect 2960 2345 2962 2361
rect 3080 2345 3082 2361
rect 3192 2345 3194 2361
rect 3304 2345 3306 2361
rect 3416 2345 3418 2361
rect 3504 2345 3506 2361
rect 1894 2344 1900 2345
rect 1831 2341 1835 2342
rect 1870 2341 1876 2342
rect 112 2313 114 2341
rect 1408 2331 1410 2341
rect 1488 2331 1490 2341
rect 1568 2331 1570 2341
rect 1648 2331 1650 2341
rect 1406 2330 1412 2331
rect 1406 2326 1407 2330
rect 1411 2326 1412 2330
rect 1406 2325 1412 2326
rect 1486 2330 1492 2331
rect 1486 2326 1487 2330
rect 1491 2326 1492 2330
rect 1486 2325 1492 2326
rect 1566 2330 1572 2331
rect 1566 2326 1567 2330
rect 1571 2326 1572 2330
rect 1566 2325 1572 2326
rect 1646 2330 1652 2331
rect 1646 2326 1647 2330
rect 1651 2326 1652 2330
rect 1646 2325 1652 2326
rect 1832 2313 1834 2341
rect 1870 2337 1871 2341
rect 1875 2337 1876 2341
rect 1894 2340 1895 2344
rect 1899 2340 1900 2344
rect 1894 2339 1900 2340
rect 2014 2344 2020 2345
rect 2014 2340 2015 2344
rect 2019 2340 2020 2344
rect 2014 2339 2020 2340
rect 2174 2344 2180 2345
rect 2174 2340 2175 2344
rect 2179 2340 2180 2344
rect 2174 2339 2180 2340
rect 2342 2344 2348 2345
rect 2342 2340 2343 2344
rect 2347 2340 2348 2344
rect 2342 2339 2348 2340
rect 2510 2344 2516 2345
rect 2510 2340 2511 2344
rect 2515 2340 2516 2344
rect 2510 2339 2516 2340
rect 2670 2344 2676 2345
rect 2670 2340 2671 2344
rect 2675 2340 2676 2344
rect 2670 2339 2676 2340
rect 2822 2344 2828 2345
rect 2822 2340 2823 2344
rect 2827 2340 2828 2344
rect 2822 2339 2828 2340
rect 2958 2344 2964 2345
rect 2958 2340 2959 2344
rect 2963 2340 2964 2344
rect 2958 2339 2964 2340
rect 3078 2344 3084 2345
rect 3078 2340 3079 2344
rect 3083 2340 3084 2344
rect 3078 2339 3084 2340
rect 3190 2344 3196 2345
rect 3190 2340 3191 2344
rect 3195 2340 3196 2344
rect 3190 2339 3196 2340
rect 3302 2344 3308 2345
rect 3302 2340 3303 2344
rect 3307 2340 3308 2344
rect 3302 2339 3308 2340
rect 3414 2344 3420 2345
rect 3414 2340 3415 2344
rect 3419 2340 3420 2344
rect 3414 2339 3420 2340
rect 3502 2344 3508 2345
rect 3502 2340 3503 2344
rect 3507 2340 3508 2344
rect 3592 2342 3594 2361
rect 3502 2339 3508 2340
rect 3590 2341 3596 2342
rect 1870 2336 1876 2337
rect 3590 2337 3591 2341
rect 3595 2337 3596 2341
rect 3590 2336 3596 2337
rect 1870 2324 1876 2325
rect 1870 2320 1871 2324
rect 1875 2320 1876 2324
rect 1870 2319 1876 2320
rect 3590 2324 3596 2325
rect 3590 2320 3591 2324
rect 3595 2320 3596 2324
rect 3590 2319 3596 2320
rect 110 2312 116 2313
rect 110 2308 111 2312
rect 115 2308 116 2312
rect 110 2307 116 2308
rect 1830 2312 1836 2313
rect 1830 2308 1831 2312
rect 1835 2308 1836 2312
rect 1830 2307 1836 2308
rect 110 2295 116 2296
rect 110 2291 111 2295
rect 115 2291 116 2295
rect 1830 2295 1836 2296
rect 110 2290 116 2291
rect 1398 2292 1404 2293
rect 112 2263 114 2290
rect 1398 2288 1399 2292
rect 1403 2288 1404 2292
rect 1398 2287 1404 2288
rect 1478 2292 1484 2293
rect 1478 2288 1479 2292
rect 1483 2288 1484 2292
rect 1478 2287 1484 2288
rect 1558 2292 1564 2293
rect 1558 2288 1559 2292
rect 1563 2288 1564 2292
rect 1558 2287 1564 2288
rect 1638 2292 1644 2293
rect 1638 2288 1639 2292
rect 1643 2288 1644 2292
rect 1830 2291 1831 2295
rect 1835 2291 1836 2295
rect 1872 2291 1874 2319
rect 1902 2306 1908 2307
rect 1902 2302 1903 2306
rect 1907 2302 1908 2306
rect 1902 2301 1908 2302
rect 2022 2306 2028 2307
rect 2022 2302 2023 2306
rect 2027 2302 2028 2306
rect 2022 2301 2028 2302
rect 2182 2306 2188 2307
rect 2182 2302 2183 2306
rect 2187 2302 2188 2306
rect 2182 2301 2188 2302
rect 2350 2306 2356 2307
rect 2350 2302 2351 2306
rect 2355 2302 2356 2306
rect 2350 2301 2356 2302
rect 2518 2306 2524 2307
rect 2518 2302 2519 2306
rect 2523 2302 2524 2306
rect 2518 2301 2524 2302
rect 2678 2306 2684 2307
rect 2678 2302 2679 2306
rect 2683 2302 2684 2306
rect 2678 2301 2684 2302
rect 2830 2306 2836 2307
rect 2830 2302 2831 2306
rect 2835 2302 2836 2306
rect 2830 2301 2836 2302
rect 2966 2306 2972 2307
rect 2966 2302 2967 2306
rect 2971 2302 2972 2306
rect 2966 2301 2972 2302
rect 3086 2306 3092 2307
rect 3086 2302 3087 2306
rect 3091 2302 3092 2306
rect 3086 2301 3092 2302
rect 3198 2306 3204 2307
rect 3198 2302 3199 2306
rect 3203 2302 3204 2306
rect 3198 2301 3204 2302
rect 3310 2306 3316 2307
rect 3310 2302 3311 2306
rect 3315 2302 3316 2306
rect 3310 2301 3316 2302
rect 3422 2306 3428 2307
rect 3422 2302 3423 2306
rect 3427 2302 3428 2306
rect 3422 2301 3428 2302
rect 3510 2306 3516 2307
rect 3510 2302 3511 2306
rect 3515 2302 3516 2306
rect 3510 2301 3516 2302
rect 1904 2291 1906 2301
rect 2024 2291 2026 2301
rect 2184 2291 2186 2301
rect 2352 2291 2354 2301
rect 2520 2291 2522 2301
rect 2680 2291 2682 2301
rect 2832 2291 2834 2301
rect 2968 2291 2970 2301
rect 3088 2291 3090 2301
rect 3200 2291 3202 2301
rect 3312 2291 3314 2301
rect 3424 2291 3426 2301
rect 3512 2291 3514 2301
rect 3592 2291 3594 2319
rect 1830 2290 1836 2291
rect 1871 2290 1875 2291
rect 1638 2287 1644 2288
rect 1400 2263 1402 2287
rect 1480 2263 1482 2287
rect 1560 2263 1562 2287
rect 1640 2263 1642 2287
rect 1832 2263 1834 2290
rect 1871 2285 1875 2286
rect 1903 2290 1907 2291
rect 1903 2285 1907 2286
rect 2023 2290 2027 2291
rect 2023 2285 2027 2286
rect 2031 2290 2035 2291
rect 2031 2285 2035 2286
rect 2183 2290 2187 2291
rect 2183 2285 2187 2286
rect 2351 2290 2355 2291
rect 2351 2285 2355 2286
rect 2367 2290 2371 2291
rect 2367 2285 2371 2286
rect 2519 2290 2523 2291
rect 2519 2285 2523 2286
rect 2575 2290 2579 2291
rect 2575 2285 2579 2286
rect 2679 2290 2683 2291
rect 2679 2285 2683 2286
rect 2791 2290 2795 2291
rect 2791 2285 2795 2286
rect 2831 2290 2835 2291
rect 2831 2285 2835 2286
rect 2967 2290 2971 2291
rect 2967 2285 2971 2286
rect 3023 2290 3027 2291
rect 3023 2285 3027 2286
rect 3087 2290 3091 2291
rect 3087 2285 3091 2286
rect 3199 2290 3203 2291
rect 3199 2285 3203 2286
rect 3255 2290 3259 2291
rect 3255 2285 3259 2286
rect 3311 2290 3315 2291
rect 3311 2285 3315 2286
rect 3423 2290 3427 2291
rect 3423 2285 3427 2286
rect 3495 2290 3499 2291
rect 3495 2285 3499 2286
rect 3511 2290 3515 2291
rect 3511 2285 3515 2286
rect 3591 2290 3595 2291
rect 3591 2285 3595 2286
rect 111 2262 115 2263
rect 111 2257 115 2258
rect 135 2262 139 2263
rect 135 2257 139 2258
rect 215 2262 219 2263
rect 215 2257 219 2258
rect 295 2262 299 2263
rect 295 2257 299 2258
rect 383 2262 387 2263
rect 383 2257 387 2258
rect 519 2262 523 2263
rect 519 2257 523 2258
rect 671 2262 675 2263
rect 671 2257 675 2258
rect 831 2262 835 2263
rect 831 2257 835 2258
rect 999 2262 1003 2263
rect 999 2257 1003 2258
rect 1159 2262 1163 2263
rect 1159 2257 1163 2258
rect 1311 2262 1315 2263
rect 1311 2257 1315 2258
rect 1399 2262 1403 2263
rect 1399 2257 1403 2258
rect 1455 2262 1459 2263
rect 1455 2257 1459 2258
rect 1479 2262 1483 2263
rect 1479 2257 1483 2258
rect 1559 2262 1563 2263
rect 1559 2257 1563 2258
rect 1607 2262 1611 2263
rect 1607 2257 1611 2258
rect 1639 2262 1643 2263
rect 1639 2257 1643 2258
rect 1743 2262 1747 2263
rect 1743 2257 1747 2258
rect 1831 2262 1835 2263
rect 1831 2257 1835 2258
rect 1872 2257 1874 2285
rect 1904 2275 1906 2285
rect 2032 2275 2034 2285
rect 2184 2275 2186 2285
rect 2368 2275 2370 2285
rect 2576 2275 2578 2285
rect 2792 2275 2794 2285
rect 3024 2275 3026 2285
rect 3256 2275 3258 2285
rect 3496 2275 3498 2285
rect 1902 2274 1908 2275
rect 1902 2270 1903 2274
rect 1907 2270 1908 2274
rect 1902 2269 1908 2270
rect 2030 2274 2036 2275
rect 2030 2270 2031 2274
rect 2035 2270 2036 2274
rect 2030 2269 2036 2270
rect 2182 2274 2188 2275
rect 2182 2270 2183 2274
rect 2187 2270 2188 2274
rect 2182 2269 2188 2270
rect 2366 2274 2372 2275
rect 2366 2270 2367 2274
rect 2371 2270 2372 2274
rect 2366 2269 2372 2270
rect 2574 2274 2580 2275
rect 2574 2270 2575 2274
rect 2579 2270 2580 2274
rect 2574 2269 2580 2270
rect 2790 2274 2796 2275
rect 2790 2270 2791 2274
rect 2795 2270 2796 2274
rect 2790 2269 2796 2270
rect 3022 2274 3028 2275
rect 3022 2270 3023 2274
rect 3027 2270 3028 2274
rect 3022 2269 3028 2270
rect 3254 2274 3260 2275
rect 3254 2270 3255 2274
rect 3259 2270 3260 2274
rect 3254 2269 3260 2270
rect 3494 2274 3500 2275
rect 3494 2270 3495 2274
rect 3499 2270 3500 2274
rect 3494 2269 3500 2270
rect 3592 2257 3594 2285
rect 112 2238 114 2257
rect 136 2241 138 2257
rect 216 2241 218 2257
rect 296 2241 298 2257
rect 384 2241 386 2257
rect 520 2241 522 2257
rect 672 2241 674 2257
rect 832 2241 834 2257
rect 1000 2241 1002 2257
rect 1160 2241 1162 2257
rect 1312 2241 1314 2257
rect 1456 2241 1458 2257
rect 1608 2241 1610 2257
rect 1744 2241 1746 2257
rect 134 2240 140 2241
rect 110 2237 116 2238
rect 110 2233 111 2237
rect 115 2233 116 2237
rect 134 2236 135 2240
rect 139 2236 140 2240
rect 134 2235 140 2236
rect 214 2240 220 2241
rect 214 2236 215 2240
rect 219 2236 220 2240
rect 214 2235 220 2236
rect 294 2240 300 2241
rect 294 2236 295 2240
rect 299 2236 300 2240
rect 294 2235 300 2236
rect 382 2240 388 2241
rect 382 2236 383 2240
rect 387 2236 388 2240
rect 382 2235 388 2236
rect 518 2240 524 2241
rect 518 2236 519 2240
rect 523 2236 524 2240
rect 518 2235 524 2236
rect 670 2240 676 2241
rect 670 2236 671 2240
rect 675 2236 676 2240
rect 670 2235 676 2236
rect 830 2240 836 2241
rect 830 2236 831 2240
rect 835 2236 836 2240
rect 830 2235 836 2236
rect 998 2240 1004 2241
rect 998 2236 999 2240
rect 1003 2236 1004 2240
rect 998 2235 1004 2236
rect 1158 2240 1164 2241
rect 1158 2236 1159 2240
rect 1163 2236 1164 2240
rect 1158 2235 1164 2236
rect 1310 2240 1316 2241
rect 1310 2236 1311 2240
rect 1315 2236 1316 2240
rect 1310 2235 1316 2236
rect 1454 2240 1460 2241
rect 1454 2236 1455 2240
rect 1459 2236 1460 2240
rect 1454 2235 1460 2236
rect 1606 2240 1612 2241
rect 1606 2236 1607 2240
rect 1611 2236 1612 2240
rect 1606 2235 1612 2236
rect 1742 2240 1748 2241
rect 1742 2236 1743 2240
rect 1747 2236 1748 2240
rect 1832 2238 1834 2257
rect 1870 2256 1876 2257
rect 1870 2252 1871 2256
rect 1875 2252 1876 2256
rect 1870 2251 1876 2252
rect 3590 2256 3596 2257
rect 3590 2252 3591 2256
rect 3595 2252 3596 2256
rect 3590 2251 3596 2252
rect 1870 2239 1876 2240
rect 1742 2235 1748 2236
rect 1830 2237 1836 2238
rect 110 2232 116 2233
rect 1830 2233 1831 2237
rect 1835 2233 1836 2237
rect 1870 2235 1871 2239
rect 1875 2235 1876 2239
rect 3590 2239 3596 2240
rect 1870 2234 1876 2235
rect 1894 2236 1900 2237
rect 1830 2232 1836 2233
rect 110 2220 116 2221
rect 110 2216 111 2220
rect 115 2216 116 2220
rect 110 2215 116 2216
rect 1830 2220 1836 2221
rect 1830 2216 1831 2220
rect 1835 2216 1836 2220
rect 1830 2215 1836 2216
rect 112 2183 114 2215
rect 142 2202 148 2203
rect 142 2198 143 2202
rect 147 2198 148 2202
rect 142 2197 148 2198
rect 222 2202 228 2203
rect 222 2198 223 2202
rect 227 2198 228 2202
rect 222 2197 228 2198
rect 302 2202 308 2203
rect 302 2198 303 2202
rect 307 2198 308 2202
rect 302 2197 308 2198
rect 390 2202 396 2203
rect 390 2198 391 2202
rect 395 2198 396 2202
rect 390 2197 396 2198
rect 526 2202 532 2203
rect 526 2198 527 2202
rect 531 2198 532 2202
rect 526 2197 532 2198
rect 678 2202 684 2203
rect 678 2198 679 2202
rect 683 2198 684 2202
rect 678 2197 684 2198
rect 838 2202 844 2203
rect 838 2198 839 2202
rect 843 2198 844 2202
rect 838 2197 844 2198
rect 1006 2202 1012 2203
rect 1006 2198 1007 2202
rect 1011 2198 1012 2202
rect 1006 2197 1012 2198
rect 1166 2202 1172 2203
rect 1166 2198 1167 2202
rect 1171 2198 1172 2202
rect 1166 2197 1172 2198
rect 1318 2202 1324 2203
rect 1318 2198 1319 2202
rect 1323 2198 1324 2202
rect 1318 2197 1324 2198
rect 1462 2202 1468 2203
rect 1462 2198 1463 2202
rect 1467 2198 1468 2202
rect 1462 2197 1468 2198
rect 1614 2202 1620 2203
rect 1614 2198 1615 2202
rect 1619 2198 1620 2202
rect 1614 2197 1620 2198
rect 1750 2202 1756 2203
rect 1750 2198 1751 2202
rect 1755 2198 1756 2202
rect 1750 2197 1756 2198
rect 144 2183 146 2197
rect 224 2183 226 2197
rect 304 2183 306 2197
rect 392 2183 394 2197
rect 528 2183 530 2197
rect 680 2183 682 2197
rect 840 2183 842 2197
rect 1008 2183 1010 2197
rect 1168 2183 1170 2197
rect 1320 2183 1322 2197
rect 1464 2183 1466 2197
rect 1616 2183 1618 2197
rect 1752 2183 1754 2197
rect 1832 2183 1834 2215
rect 1872 2195 1874 2234
rect 1894 2232 1895 2236
rect 1899 2232 1900 2236
rect 1894 2231 1900 2232
rect 2022 2236 2028 2237
rect 2022 2232 2023 2236
rect 2027 2232 2028 2236
rect 2022 2231 2028 2232
rect 2174 2236 2180 2237
rect 2174 2232 2175 2236
rect 2179 2232 2180 2236
rect 2174 2231 2180 2232
rect 2358 2236 2364 2237
rect 2358 2232 2359 2236
rect 2363 2232 2364 2236
rect 2358 2231 2364 2232
rect 2566 2236 2572 2237
rect 2566 2232 2567 2236
rect 2571 2232 2572 2236
rect 2566 2231 2572 2232
rect 2782 2236 2788 2237
rect 2782 2232 2783 2236
rect 2787 2232 2788 2236
rect 2782 2231 2788 2232
rect 3014 2236 3020 2237
rect 3014 2232 3015 2236
rect 3019 2232 3020 2236
rect 3014 2231 3020 2232
rect 3246 2236 3252 2237
rect 3246 2232 3247 2236
rect 3251 2232 3252 2236
rect 3246 2231 3252 2232
rect 3486 2236 3492 2237
rect 3486 2232 3487 2236
rect 3491 2232 3492 2236
rect 3590 2235 3591 2239
rect 3595 2235 3596 2239
rect 3590 2234 3596 2235
rect 3486 2231 3492 2232
rect 1896 2195 1898 2231
rect 2024 2195 2026 2231
rect 2176 2195 2178 2231
rect 2360 2195 2362 2231
rect 2568 2195 2570 2231
rect 2784 2195 2786 2231
rect 3016 2195 3018 2231
rect 3248 2195 3250 2231
rect 3488 2195 3490 2231
rect 3592 2195 3594 2234
rect 1871 2194 1875 2195
rect 1871 2189 1875 2190
rect 1895 2194 1899 2195
rect 1895 2189 1899 2190
rect 2023 2194 2027 2195
rect 2023 2189 2027 2190
rect 2175 2194 2179 2195
rect 2175 2189 2179 2190
rect 2199 2194 2203 2195
rect 2199 2189 2203 2190
rect 2295 2194 2299 2195
rect 2295 2189 2299 2190
rect 2359 2194 2363 2195
rect 2359 2189 2363 2190
rect 2399 2194 2403 2195
rect 2399 2189 2403 2190
rect 2519 2194 2523 2195
rect 2519 2189 2523 2190
rect 2567 2194 2571 2195
rect 2567 2189 2571 2190
rect 2639 2194 2643 2195
rect 2639 2189 2643 2190
rect 2759 2194 2763 2195
rect 2759 2189 2763 2190
rect 2783 2194 2787 2195
rect 2783 2189 2787 2190
rect 2879 2194 2883 2195
rect 2879 2189 2883 2190
rect 2991 2194 2995 2195
rect 2991 2189 2995 2190
rect 3015 2194 3019 2195
rect 3015 2189 3019 2190
rect 3095 2194 3099 2195
rect 3095 2189 3099 2190
rect 3199 2194 3203 2195
rect 3199 2189 3203 2190
rect 3247 2194 3251 2195
rect 3247 2189 3251 2190
rect 3303 2194 3307 2195
rect 3303 2189 3307 2190
rect 3407 2194 3411 2195
rect 3407 2189 3411 2190
rect 3487 2194 3491 2195
rect 3487 2189 3491 2190
rect 3503 2194 3507 2195
rect 3503 2189 3507 2190
rect 3591 2194 3595 2195
rect 3591 2189 3595 2190
rect 111 2182 115 2183
rect 111 2177 115 2178
rect 143 2182 147 2183
rect 143 2177 147 2178
rect 191 2182 195 2183
rect 191 2177 195 2178
rect 223 2182 227 2183
rect 223 2177 227 2178
rect 303 2182 307 2183
rect 303 2177 307 2178
rect 311 2182 315 2183
rect 311 2177 315 2178
rect 391 2182 395 2183
rect 391 2177 395 2178
rect 463 2182 467 2183
rect 463 2177 467 2178
rect 527 2182 531 2183
rect 527 2177 531 2178
rect 639 2182 643 2183
rect 639 2177 643 2178
rect 679 2182 683 2183
rect 679 2177 683 2178
rect 823 2182 827 2183
rect 823 2177 827 2178
rect 839 2182 843 2183
rect 839 2177 843 2178
rect 1007 2182 1011 2183
rect 1007 2177 1011 2178
rect 1015 2182 1019 2183
rect 1015 2177 1019 2178
rect 1167 2182 1171 2183
rect 1167 2177 1171 2178
rect 1199 2182 1203 2183
rect 1199 2177 1203 2178
rect 1319 2182 1323 2183
rect 1319 2177 1323 2178
rect 1391 2182 1395 2183
rect 1391 2177 1395 2178
rect 1463 2182 1467 2183
rect 1463 2177 1467 2178
rect 1583 2182 1587 2183
rect 1583 2177 1587 2178
rect 1615 2182 1619 2183
rect 1615 2177 1619 2178
rect 1751 2182 1755 2183
rect 1751 2177 1755 2178
rect 1831 2182 1835 2183
rect 1831 2177 1835 2178
rect 112 2149 114 2177
rect 192 2167 194 2177
rect 312 2167 314 2177
rect 464 2167 466 2177
rect 640 2167 642 2177
rect 824 2167 826 2177
rect 1016 2167 1018 2177
rect 1200 2167 1202 2177
rect 1392 2167 1394 2177
rect 1584 2167 1586 2177
rect 1752 2167 1754 2177
rect 190 2166 196 2167
rect 190 2162 191 2166
rect 195 2162 196 2166
rect 190 2161 196 2162
rect 310 2166 316 2167
rect 310 2162 311 2166
rect 315 2162 316 2166
rect 310 2161 316 2162
rect 462 2166 468 2167
rect 462 2162 463 2166
rect 467 2162 468 2166
rect 462 2161 468 2162
rect 638 2166 644 2167
rect 638 2162 639 2166
rect 643 2162 644 2166
rect 638 2161 644 2162
rect 822 2166 828 2167
rect 822 2162 823 2166
rect 827 2162 828 2166
rect 822 2161 828 2162
rect 1014 2166 1020 2167
rect 1014 2162 1015 2166
rect 1019 2162 1020 2166
rect 1014 2161 1020 2162
rect 1198 2166 1204 2167
rect 1198 2162 1199 2166
rect 1203 2162 1204 2166
rect 1198 2161 1204 2162
rect 1390 2166 1396 2167
rect 1390 2162 1391 2166
rect 1395 2162 1396 2166
rect 1390 2161 1396 2162
rect 1582 2166 1588 2167
rect 1582 2162 1583 2166
rect 1587 2162 1588 2166
rect 1582 2161 1588 2162
rect 1750 2166 1756 2167
rect 1750 2162 1751 2166
rect 1755 2162 1756 2166
rect 1750 2161 1756 2162
rect 1832 2149 1834 2177
rect 1872 2170 1874 2189
rect 2200 2173 2202 2189
rect 2296 2173 2298 2189
rect 2400 2173 2402 2189
rect 2520 2173 2522 2189
rect 2640 2173 2642 2189
rect 2760 2173 2762 2189
rect 2880 2173 2882 2189
rect 2992 2173 2994 2189
rect 3096 2173 3098 2189
rect 3200 2173 3202 2189
rect 3304 2173 3306 2189
rect 3408 2173 3410 2189
rect 3504 2173 3506 2189
rect 2198 2172 2204 2173
rect 1870 2169 1876 2170
rect 1870 2165 1871 2169
rect 1875 2165 1876 2169
rect 2198 2168 2199 2172
rect 2203 2168 2204 2172
rect 2198 2167 2204 2168
rect 2294 2172 2300 2173
rect 2294 2168 2295 2172
rect 2299 2168 2300 2172
rect 2294 2167 2300 2168
rect 2398 2172 2404 2173
rect 2398 2168 2399 2172
rect 2403 2168 2404 2172
rect 2398 2167 2404 2168
rect 2518 2172 2524 2173
rect 2518 2168 2519 2172
rect 2523 2168 2524 2172
rect 2518 2167 2524 2168
rect 2638 2172 2644 2173
rect 2638 2168 2639 2172
rect 2643 2168 2644 2172
rect 2638 2167 2644 2168
rect 2758 2172 2764 2173
rect 2758 2168 2759 2172
rect 2763 2168 2764 2172
rect 2758 2167 2764 2168
rect 2878 2172 2884 2173
rect 2878 2168 2879 2172
rect 2883 2168 2884 2172
rect 2878 2167 2884 2168
rect 2990 2172 2996 2173
rect 2990 2168 2991 2172
rect 2995 2168 2996 2172
rect 2990 2167 2996 2168
rect 3094 2172 3100 2173
rect 3094 2168 3095 2172
rect 3099 2168 3100 2172
rect 3094 2167 3100 2168
rect 3198 2172 3204 2173
rect 3198 2168 3199 2172
rect 3203 2168 3204 2172
rect 3198 2167 3204 2168
rect 3302 2172 3308 2173
rect 3302 2168 3303 2172
rect 3307 2168 3308 2172
rect 3302 2167 3308 2168
rect 3406 2172 3412 2173
rect 3406 2168 3407 2172
rect 3411 2168 3412 2172
rect 3406 2167 3412 2168
rect 3502 2172 3508 2173
rect 3502 2168 3503 2172
rect 3507 2168 3508 2172
rect 3592 2170 3594 2189
rect 3502 2167 3508 2168
rect 3590 2169 3596 2170
rect 1870 2164 1876 2165
rect 3590 2165 3591 2169
rect 3595 2165 3596 2169
rect 3590 2164 3596 2165
rect 1870 2152 1876 2153
rect 110 2148 116 2149
rect 110 2144 111 2148
rect 115 2144 116 2148
rect 110 2143 116 2144
rect 1830 2148 1836 2149
rect 1830 2144 1831 2148
rect 1835 2144 1836 2148
rect 1870 2148 1871 2152
rect 1875 2148 1876 2152
rect 1870 2147 1876 2148
rect 3590 2152 3596 2153
rect 3590 2148 3591 2152
rect 3595 2148 3596 2152
rect 3590 2147 3596 2148
rect 1830 2143 1836 2144
rect 110 2131 116 2132
rect 110 2127 111 2131
rect 115 2127 116 2131
rect 1830 2131 1836 2132
rect 110 2126 116 2127
rect 182 2128 188 2129
rect 112 2103 114 2126
rect 182 2124 183 2128
rect 187 2124 188 2128
rect 182 2123 188 2124
rect 302 2128 308 2129
rect 302 2124 303 2128
rect 307 2124 308 2128
rect 302 2123 308 2124
rect 454 2128 460 2129
rect 454 2124 455 2128
rect 459 2124 460 2128
rect 454 2123 460 2124
rect 630 2128 636 2129
rect 630 2124 631 2128
rect 635 2124 636 2128
rect 630 2123 636 2124
rect 814 2128 820 2129
rect 814 2124 815 2128
rect 819 2124 820 2128
rect 814 2123 820 2124
rect 1006 2128 1012 2129
rect 1006 2124 1007 2128
rect 1011 2124 1012 2128
rect 1006 2123 1012 2124
rect 1190 2128 1196 2129
rect 1190 2124 1191 2128
rect 1195 2124 1196 2128
rect 1190 2123 1196 2124
rect 1382 2128 1388 2129
rect 1382 2124 1383 2128
rect 1387 2124 1388 2128
rect 1382 2123 1388 2124
rect 1574 2128 1580 2129
rect 1574 2124 1575 2128
rect 1579 2124 1580 2128
rect 1574 2123 1580 2124
rect 1742 2128 1748 2129
rect 1742 2124 1743 2128
rect 1747 2124 1748 2128
rect 1830 2127 1831 2131
rect 1835 2127 1836 2131
rect 1830 2126 1836 2127
rect 1742 2123 1748 2124
rect 184 2103 186 2123
rect 304 2103 306 2123
rect 456 2103 458 2123
rect 632 2103 634 2123
rect 816 2103 818 2123
rect 1008 2103 1010 2123
rect 1192 2103 1194 2123
rect 1384 2103 1386 2123
rect 1576 2103 1578 2123
rect 1744 2103 1746 2123
rect 1832 2103 1834 2126
rect 1872 2107 1874 2147
rect 2206 2134 2212 2135
rect 2206 2130 2207 2134
rect 2211 2130 2212 2134
rect 2206 2129 2212 2130
rect 2302 2134 2308 2135
rect 2302 2130 2303 2134
rect 2307 2130 2308 2134
rect 2302 2129 2308 2130
rect 2406 2134 2412 2135
rect 2406 2130 2407 2134
rect 2411 2130 2412 2134
rect 2406 2129 2412 2130
rect 2526 2134 2532 2135
rect 2526 2130 2527 2134
rect 2531 2130 2532 2134
rect 2526 2129 2532 2130
rect 2646 2134 2652 2135
rect 2646 2130 2647 2134
rect 2651 2130 2652 2134
rect 2646 2129 2652 2130
rect 2766 2134 2772 2135
rect 2766 2130 2767 2134
rect 2771 2130 2772 2134
rect 2766 2129 2772 2130
rect 2886 2134 2892 2135
rect 2886 2130 2887 2134
rect 2891 2130 2892 2134
rect 2886 2129 2892 2130
rect 2998 2134 3004 2135
rect 2998 2130 2999 2134
rect 3003 2130 3004 2134
rect 2998 2129 3004 2130
rect 3102 2134 3108 2135
rect 3102 2130 3103 2134
rect 3107 2130 3108 2134
rect 3102 2129 3108 2130
rect 3206 2134 3212 2135
rect 3206 2130 3207 2134
rect 3211 2130 3212 2134
rect 3206 2129 3212 2130
rect 3310 2134 3316 2135
rect 3310 2130 3311 2134
rect 3315 2130 3316 2134
rect 3310 2129 3316 2130
rect 3414 2134 3420 2135
rect 3414 2130 3415 2134
rect 3419 2130 3420 2134
rect 3414 2129 3420 2130
rect 3510 2134 3516 2135
rect 3510 2130 3511 2134
rect 3515 2130 3516 2134
rect 3510 2129 3516 2130
rect 2208 2107 2210 2129
rect 2304 2107 2306 2129
rect 2408 2107 2410 2129
rect 2528 2107 2530 2129
rect 2648 2107 2650 2129
rect 2768 2107 2770 2129
rect 2888 2107 2890 2129
rect 3000 2107 3002 2129
rect 3104 2107 3106 2129
rect 3208 2107 3210 2129
rect 3312 2107 3314 2129
rect 3416 2107 3418 2129
rect 3512 2107 3514 2129
rect 3592 2107 3594 2147
rect 1871 2106 1875 2107
rect 111 2102 115 2103
rect 111 2097 115 2098
rect 183 2102 187 2103
rect 183 2097 187 2098
rect 215 2102 219 2103
rect 215 2097 219 2098
rect 303 2102 307 2103
rect 303 2097 307 2098
rect 359 2102 363 2103
rect 359 2097 363 2098
rect 455 2102 459 2103
rect 455 2097 459 2098
rect 519 2102 523 2103
rect 519 2097 523 2098
rect 631 2102 635 2103
rect 631 2097 635 2098
rect 703 2102 707 2103
rect 703 2097 707 2098
rect 815 2102 819 2103
rect 815 2097 819 2098
rect 895 2102 899 2103
rect 895 2097 899 2098
rect 1007 2102 1011 2103
rect 1007 2097 1011 2098
rect 1103 2102 1107 2103
rect 1103 2097 1107 2098
rect 1191 2102 1195 2103
rect 1191 2097 1195 2098
rect 1311 2102 1315 2103
rect 1311 2097 1315 2098
rect 1383 2102 1387 2103
rect 1383 2097 1387 2098
rect 1527 2102 1531 2103
rect 1527 2097 1531 2098
rect 1575 2102 1579 2103
rect 1575 2097 1579 2098
rect 1743 2102 1747 2103
rect 1743 2097 1747 2098
rect 1831 2102 1835 2103
rect 1871 2101 1875 2102
rect 2175 2106 2179 2107
rect 2175 2101 2179 2102
rect 2207 2106 2211 2107
rect 2207 2101 2211 2102
rect 2271 2106 2275 2107
rect 2271 2101 2275 2102
rect 2303 2106 2307 2107
rect 2303 2101 2307 2102
rect 2375 2106 2379 2107
rect 2375 2101 2379 2102
rect 2407 2106 2411 2107
rect 2407 2101 2411 2102
rect 2487 2106 2491 2107
rect 2487 2101 2491 2102
rect 2527 2106 2531 2107
rect 2527 2101 2531 2102
rect 2607 2106 2611 2107
rect 2607 2101 2611 2102
rect 2647 2106 2651 2107
rect 2647 2101 2651 2102
rect 2727 2106 2731 2107
rect 2727 2101 2731 2102
rect 2767 2106 2771 2107
rect 2767 2101 2771 2102
rect 2847 2106 2851 2107
rect 2847 2101 2851 2102
rect 2887 2106 2891 2107
rect 2887 2101 2891 2102
rect 2967 2106 2971 2107
rect 2967 2101 2971 2102
rect 2999 2106 3003 2107
rect 2999 2101 3003 2102
rect 3079 2106 3083 2107
rect 3079 2101 3083 2102
rect 3103 2106 3107 2107
rect 3103 2101 3107 2102
rect 3191 2106 3195 2107
rect 3191 2101 3195 2102
rect 3207 2106 3211 2107
rect 3207 2101 3211 2102
rect 3303 2106 3307 2107
rect 3303 2101 3307 2102
rect 3311 2106 3315 2107
rect 3311 2101 3315 2102
rect 3415 2106 3419 2107
rect 3415 2101 3419 2102
rect 3511 2106 3515 2107
rect 3511 2101 3515 2102
rect 3591 2106 3595 2107
rect 3591 2101 3595 2102
rect 1831 2097 1835 2098
rect 112 2078 114 2097
rect 216 2081 218 2097
rect 360 2081 362 2097
rect 520 2081 522 2097
rect 704 2081 706 2097
rect 896 2081 898 2097
rect 1104 2081 1106 2097
rect 1312 2081 1314 2097
rect 1528 2081 1530 2097
rect 1744 2081 1746 2097
rect 214 2080 220 2081
rect 110 2077 116 2078
rect 110 2073 111 2077
rect 115 2073 116 2077
rect 214 2076 215 2080
rect 219 2076 220 2080
rect 214 2075 220 2076
rect 358 2080 364 2081
rect 358 2076 359 2080
rect 363 2076 364 2080
rect 358 2075 364 2076
rect 518 2080 524 2081
rect 518 2076 519 2080
rect 523 2076 524 2080
rect 518 2075 524 2076
rect 702 2080 708 2081
rect 702 2076 703 2080
rect 707 2076 708 2080
rect 702 2075 708 2076
rect 894 2080 900 2081
rect 894 2076 895 2080
rect 899 2076 900 2080
rect 894 2075 900 2076
rect 1102 2080 1108 2081
rect 1102 2076 1103 2080
rect 1107 2076 1108 2080
rect 1102 2075 1108 2076
rect 1310 2080 1316 2081
rect 1310 2076 1311 2080
rect 1315 2076 1316 2080
rect 1310 2075 1316 2076
rect 1526 2080 1532 2081
rect 1526 2076 1527 2080
rect 1531 2076 1532 2080
rect 1526 2075 1532 2076
rect 1742 2080 1748 2081
rect 1742 2076 1743 2080
rect 1747 2076 1748 2080
rect 1832 2078 1834 2097
rect 1742 2075 1748 2076
rect 1830 2077 1836 2078
rect 110 2072 116 2073
rect 1830 2073 1831 2077
rect 1835 2073 1836 2077
rect 1872 2073 1874 2101
rect 2176 2091 2178 2101
rect 2272 2091 2274 2101
rect 2376 2091 2378 2101
rect 2488 2091 2490 2101
rect 2608 2091 2610 2101
rect 2728 2091 2730 2101
rect 2848 2091 2850 2101
rect 2968 2091 2970 2101
rect 3080 2091 3082 2101
rect 3192 2091 3194 2101
rect 3304 2091 3306 2101
rect 3416 2091 3418 2101
rect 3512 2091 3514 2101
rect 2174 2090 2180 2091
rect 2174 2086 2175 2090
rect 2179 2086 2180 2090
rect 2174 2085 2180 2086
rect 2270 2090 2276 2091
rect 2270 2086 2271 2090
rect 2275 2086 2276 2090
rect 2270 2085 2276 2086
rect 2374 2090 2380 2091
rect 2374 2086 2375 2090
rect 2379 2086 2380 2090
rect 2374 2085 2380 2086
rect 2486 2090 2492 2091
rect 2486 2086 2487 2090
rect 2491 2086 2492 2090
rect 2486 2085 2492 2086
rect 2606 2090 2612 2091
rect 2606 2086 2607 2090
rect 2611 2086 2612 2090
rect 2606 2085 2612 2086
rect 2726 2090 2732 2091
rect 2726 2086 2727 2090
rect 2731 2086 2732 2090
rect 2726 2085 2732 2086
rect 2846 2090 2852 2091
rect 2846 2086 2847 2090
rect 2851 2086 2852 2090
rect 2846 2085 2852 2086
rect 2966 2090 2972 2091
rect 2966 2086 2967 2090
rect 2971 2086 2972 2090
rect 2966 2085 2972 2086
rect 3078 2090 3084 2091
rect 3078 2086 3079 2090
rect 3083 2086 3084 2090
rect 3078 2085 3084 2086
rect 3190 2090 3196 2091
rect 3190 2086 3191 2090
rect 3195 2086 3196 2090
rect 3190 2085 3196 2086
rect 3302 2090 3308 2091
rect 3302 2086 3303 2090
rect 3307 2086 3308 2090
rect 3302 2085 3308 2086
rect 3414 2090 3420 2091
rect 3414 2086 3415 2090
rect 3419 2086 3420 2090
rect 3414 2085 3420 2086
rect 3510 2090 3516 2091
rect 3510 2086 3511 2090
rect 3515 2086 3516 2090
rect 3510 2085 3516 2086
rect 3592 2073 3594 2101
rect 1830 2072 1836 2073
rect 1870 2072 1876 2073
rect 1870 2068 1871 2072
rect 1875 2068 1876 2072
rect 1870 2067 1876 2068
rect 3590 2072 3596 2073
rect 3590 2068 3591 2072
rect 3595 2068 3596 2072
rect 3590 2067 3596 2068
rect 110 2060 116 2061
rect 110 2056 111 2060
rect 115 2056 116 2060
rect 110 2055 116 2056
rect 1830 2060 1836 2061
rect 1830 2056 1831 2060
rect 1835 2056 1836 2060
rect 1830 2055 1836 2056
rect 1870 2055 1876 2056
rect 112 2027 114 2055
rect 222 2042 228 2043
rect 222 2038 223 2042
rect 227 2038 228 2042
rect 222 2037 228 2038
rect 366 2042 372 2043
rect 366 2038 367 2042
rect 371 2038 372 2042
rect 366 2037 372 2038
rect 526 2042 532 2043
rect 526 2038 527 2042
rect 531 2038 532 2042
rect 526 2037 532 2038
rect 710 2042 716 2043
rect 710 2038 711 2042
rect 715 2038 716 2042
rect 710 2037 716 2038
rect 902 2042 908 2043
rect 902 2038 903 2042
rect 907 2038 908 2042
rect 902 2037 908 2038
rect 1110 2042 1116 2043
rect 1110 2038 1111 2042
rect 1115 2038 1116 2042
rect 1110 2037 1116 2038
rect 1318 2042 1324 2043
rect 1318 2038 1319 2042
rect 1323 2038 1324 2042
rect 1318 2037 1324 2038
rect 1534 2042 1540 2043
rect 1534 2038 1535 2042
rect 1539 2038 1540 2042
rect 1534 2037 1540 2038
rect 1750 2042 1756 2043
rect 1750 2038 1751 2042
rect 1755 2038 1756 2042
rect 1750 2037 1756 2038
rect 224 2027 226 2037
rect 368 2027 370 2037
rect 528 2027 530 2037
rect 712 2027 714 2037
rect 904 2027 906 2037
rect 1112 2027 1114 2037
rect 1320 2027 1322 2037
rect 1536 2027 1538 2037
rect 1752 2027 1754 2037
rect 1832 2027 1834 2055
rect 1870 2051 1871 2055
rect 1875 2051 1876 2055
rect 3590 2055 3596 2056
rect 1870 2050 1876 2051
rect 2166 2052 2172 2053
rect 1872 2027 1874 2050
rect 2166 2048 2167 2052
rect 2171 2048 2172 2052
rect 2166 2047 2172 2048
rect 2262 2052 2268 2053
rect 2262 2048 2263 2052
rect 2267 2048 2268 2052
rect 2262 2047 2268 2048
rect 2366 2052 2372 2053
rect 2366 2048 2367 2052
rect 2371 2048 2372 2052
rect 2366 2047 2372 2048
rect 2478 2052 2484 2053
rect 2478 2048 2479 2052
rect 2483 2048 2484 2052
rect 2478 2047 2484 2048
rect 2598 2052 2604 2053
rect 2598 2048 2599 2052
rect 2603 2048 2604 2052
rect 2598 2047 2604 2048
rect 2718 2052 2724 2053
rect 2718 2048 2719 2052
rect 2723 2048 2724 2052
rect 2718 2047 2724 2048
rect 2838 2052 2844 2053
rect 2838 2048 2839 2052
rect 2843 2048 2844 2052
rect 2838 2047 2844 2048
rect 2958 2052 2964 2053
rect 2958 2048 2959 2052
rect 2963 2048 2964 2052
rect 2958 2047 2964 2048
rect 3070 2052 3076 2053
rect 3070 2048 3071 2052
rect 3075 2048 3076 2052
rect 3070 2047 3076 2048
rect 3182 2052 3188 2053
rect 3182 2048 3183 2052
rect 3187 2048 3188 2052
rect 3182 2047 3188 2048
rect 3294 2052 3300 2053
rect 3294 2048 3295 2052
rect 3299 2048 3300 2052
rect 3294 2047 3300 2048
rect 3406 2052 3412 2053
rect 3406 2048 3407 2052
rect 3411 2048 3412 2052
rect 3406 2047 3412 2048
rect 3502 2052 3508 2053
rect 3502 2048 3503 2052
rect 3507 2048 3508 2052
rect 3590 2051 3591 2055
rect 3595 2051 3596 2055
rect 3590 2050 3596 2051
rect 3502 2047 3508 2048
rect 2168 2027 2170 2047
rect 2264 2027 2266 2047
rect 2368 2027 2370 2047
rect 2480 2027 2482 2047
rect 2600 2027 2602 2047
rect 2720 2027 2722 2047
rect 2840 2027 2842 2047
rect 2960 2027 2962 2047
rect 3072 2027 3074 2047
rect 3184 2027 3186 2047
rect 3296 2027 3298 2047
rect 3408 2027 3410 2047
rect 3504 2027 3506 2047
rect 3592 2027 3594 2050
rect 111 2026 115 2027
rect 111 2021 115 2022
rect 143 2026 147 2027
rect 143 2021 147 2022
rect 223 2026 227 2027
rect 223 2021 227 2022
rect 263 2026 267 2027
rect 263 2021 267 2022
rect 367 2026 371 2027
rect 367 2021 371 2022
rect 383 2026 387 2027
rect 383 2021 387 2022
rect 495 2026 499 2027
rect 495 2021 499 2022
rect 527 2026 531 2027
rect 527 2021 531 2022
rect 607 2026 611 2027
rect 607 2021 611 2022
rect 711 2026 715 2027
rect 711 2021 715 2022
rect 719 2026 723 2027
rect 719 2021 723 2022
rect 823 2026 827 2027
rect 823 2021 827 2022
rect 903 2026 907 2027
rect 903 2021 907 2022
rect 927 2026 931 2027
rect 927 2021 931 2022
rect 1023 2026 1027 2027
rect 1023 2021 1027 2022
rect 1111 2026 1115 2027
rect 1111 2021 1115 2022
rect 1207 2026 1211 2027
rect 1207 2021 1211 2022
rect 1295 2026 1299 2027
rect 1295 2021 1299 2022
rect 1319 2026 1323 2027
rect 1319 2021 1323 2022
rect 1391 2026 1395 2027
rect 1391 2021 1395 2022
rect 1487 2026 1491 2027
rect 1487 2021 1491 2022
rect 1535 2026 1539 2027
rect 1535 2021 1539 2022
rect 1583 2026 1587 2027
rect 1583 2021 1587 2022
rect 1671 2026 1675 2027
rect 1671 2021 1675 2022
rect 1751 2026 1755 2027
rect 1751 2021 1755 2022
rect 1831 2026 1835 2027
rect 1831 2021 1835 2022
rect 1871 2026 1875 2027
rect 1871 2021 1875 2022
rect 2071 2026 2075 2027
rect 2071 2021 2075 2022
rect 2167 2026 2171 2027
rect 2167 2021 2171 2022
rect 2207 2026 2211 2027
rect 2207 2021 2211 2022
rect 2263 2026 2267 2027
rect 2263 2021 2267 2022
rect 2359 2026 2363 2027
rect 2359 2021 2363 2022
rect 2367 2026 2371 2027
rect 2367 2021 2371 2022
rect 2479 2026 2483 2027
rect 2479 2021 2483 2022
rect 2519 2026 2523 2027
rect 2519 2021 2523 2022
rect 2599 2026 2603 2027
rect 2599 2021 2603 2022
rect 2679 2026 2683 2027
rect 2679 2021 2683 2022
rect 2719 2026 2723 2027
rect 2719 2021 2723 2022
rect 2839 2026 2843 2027
rect 2839 2021 2843 2022
rect 2847 2026 2851 2027
rect 2847 2021 2851 2022
rect 2959 2026 2963 2027
rect 2959 2021 2963 2022
rect 3015 2026 3019 2027
rect 3015 2021 3019 2022
rect 3071 2026 3075 2027
rect 3071 2021 3075 2022
rect 3183 2026 3187 2027
rect 3183 2021 3187 2022
rect 3295 2026 3299 2027
rect 3295 2021 3299 2022
rect 3351 2026 3355 2027
rect 3351 2021 3355 2022
rect 3407 2026 3411 2027
rect 3407 2021 3411 2022
rect 3503 2026 3507 2027
rect 3503 2021 3507 2022
rect 3591 2026 3595 2027
rect 3591 2021 3595 2022
rect 112 1993 114 2021
rect 144 2011 146 2021
rect 264 2011 266 2021
rect 384 2011 386 2021
rect 496 2011 498 2021
rect 608 2011 610 2021
rect 720 2011 722 2021
rect 824 2011 826 2021
rect 928 2011 930 2021
rect 1024 2011 1026 2021
rect 1112 2011 1114 2021
rect 1208 2011 1210 2021
rect 1296 2011 1298 2021
rect 1392 2011 1394 2021
rect 1488 2011 1490 2021
rect 1584 2011 1586 2021
rect 1672 2011 1674 2021
rect 1752 2011 1754 2021
rect 142 2010 148 2011
rect 142 2006 143 2010
rect 147 2006 148 2010
rect 142 2005 148 2006
rect 262 2010 268 2011
rect 262 2006 263 2010
rect 267 2006 268 2010
rect 262 2005 268 2006
rect 382 2010 388 2011
rect 382 2006 383 2010
rect 387 2006 388 2010
rect 382 2005 388 2006
rect 494 2010 500 2011
rect 494 2006 495 2010
rect 499 2006 500 2010
rect 494 2005 500 2006
rect 606 2010 612 2011
rect 606 2006 607 2010
rect 611 2006 612 2010
rect 606 2005 612 2006
rect 718 2010 724 2011
rect 718 2006 719 2010
rect 723 2006 724 2010
rect 718 2005 724 2006
rect 822 2010 828 2011
rect 822 2006 823 2010
rect 827 2006 828 2010
rect 822 2005 828 2006
rect 926 2010 932 2011
rect 926 2006 927 2010
rect 931 2006 932 2010
rect 926 2005 932 2006
rect 1022 2010 1028 2011
rect 1022 2006 1023 2010
rect 1027 2006 1028 2010
rect 1022 2005 1028 2006
rect 1110 2010 1116 2011
rect 1110 2006 1111 2010
rect 1115 2006 1116 2010
rect 1110 2005 1116 2006
rect 1206 2010 1212 2011
rect 1206 2006 1207 2010
rect 1211 2006 1212 2010
rect 1206 2005 1212 2006
rect 1294 2010 1300 2011
rect 1294 2006 1295 2010
rect 1299 2006 1300 2010
rect 1294 2005 1300 2006
rect 1390 2010 1396 2011
rect 1390 2006 1391 2010
rect 1395 2006 1396 2010
rect 1390 2005 1396 2006
rect 1486 2010 1492 2011
rect 1486 2006 1487 2010
rect 1491 2006 1492 2010
rect 1486 2005 1492 2006
rect 1582 2010 1588 2011
rect 1582 2006 1583 2010
rect 1587 2006 1588 2010
rect 1582 2005 1588 2006
rect 1670 2010 1676 2011
rect 1670 2006 1671 2010
rect 1675 2006 1676 2010
rect 1670 2005 1676 2006
rect 1750 2010 1756 2011
rect 1750 2006 1751 2010
rect 1755 2006 1756 2010
rect 1750 2005 1756 2006
rect 1832 1993 1834 2021
rect 1872 2002 1874 2021
rect 2072 2005 2074 2021
rect 2208 2005 2210 2021
rect 2360 2005 2362 2021
rect 2520 2005 2522 2021
rect 2680 2005 2682 2021
rect 2848 2005 2850 2021
rect 3016 2005 3018 2021
rect 3184 2005 3186 2021
rect 3352 2005 3354 2021
rect 3504 2005 3506 2021
rect 2070 2004 2076 2005
rect 1870 2001 1876 2002
rect 1870 1997 1871 2001
rect 1875 1997 1876 2001
rect 2070 2000 2071 2004
rect 2075 2000 2076 2004
rect 2070 1999 2076 2000
rect 2206 2004 2212 2005
rect 2206 2000 2207 2004
rect 2211 2000 2212 2004
rect 2206 1999 2212 2000
rect 2358 2004 2364 2005
rect 2358 2000 2359 2004
rect 2363 2000 2364 2004
rect 2358 1999 2364 2000
rect 2518 2004 2524 2005
rect 2518 2000 2519 2004
rect 2523 2000 2524 2004
rect 2518 1999 2524 2000
rect 2678 2004 2684 2005
rect 2678 2000 2679 2004
rect 2683 2000 2684 2004
rect 2678 1999 2684 2000
rect 2846 2004 2852 2005
rect 2846 2000 2847 2004
rect 2851 2000 2852 2004
rect 2846 1999 2852 2000
rect 3014 2004 3020 2005
rect 3014 2000 3015 2004
rect 3019 2000 3020 2004
rect 3014 1999 3020 2000
rect 3182 2004 3188 2005
rect 3182 2000 3183 2004
rect 3187 2000 3188 2004
rect 3182 1999 3188 2000
rect 3350 2004 3356 2005
rect 3350 2000 3351 2004
rect 3355 2000 3356 2004
rect 3350 1999 3356 2000
rect 3502 2004 3508 2005
rect 3502 2000 3503 2004
rect 3507 2000 3508 2004
rect 3592 2002 3594 2021
rect 3502 1999 3508 2000
rect 3590 2001 3596 2002
rect 1870 1996 1876 1997
rect 3590 1997 3591 2001
rect 3595 1997 3596 2001
rect 3590 1996 3596 1997
rect 110 1992 116 1993
rect 110 1988 111 1992
rect 115 1988 116 1992
rect 110 1987 116 1988
rect 1830 1992 1836 1993
rect 1830 1988 1831 1992
rect 1835 1988 1836 1992
rect 1830 1987 1836 1988
rect 1870 1984 1876 1985
rect 1870 1980 1871 1984
rect 1875 1980 1876 1984
rect 1870 1979 1876 1980
rect 3590 1984 3596 1985
rect 3590 1980 3591 1984
rect 3595 1980 3596 1984
rect 3590 1979 3596 1980
rect 110 1975 116 1976
rect 110 1971 111 1975
rect 115 1971 116 1975
rect 1830 1975 1836 1976
rect 110 1970 116 1971
rect 134 1972 140 1973
rect 112 1943 114 1970
rect 134 1968 135 1972
rect 139 1968 140 1972
rect 134 1967 140 1968
rect 254 1972 260 1973
rect 254 1968 255 1972
rect 259 1968 260 1972
rect 254 1967 260 1968
rect 374 1972 380 1973
rect 374 1968 375 1972
rect 379 1968 380 1972
rect 374 1967 380 1968
rect 486 1972 492 1973
rect 486 1968 487 1972
rect 491 1968 492 1972
rect 486 1967 492 1968
rect 598 1972 604 1973
rect 598 1968 599 1972
rect 603 1968 604 1972
rect 598 1967 604 1968
rect 710 1972 716 1973
rect 710 1968 711 1972
rect 715 1968 716 1972
rect 710 1967 716 1968
rect 814 1972 820 1973
rect 814 1968 815 1972
rect 819 1968 820 1972
rect 814 1967 820 1968
rect 918 1972 924 1973
rect 918 1968 919 1972
rect 923 1968 924 1972
rect 918 1967 924 1968
rect 1014 1972 1020 1973
rect 1014 1968 1015 1972
rect 1019 1968 1020 1972
rect 1014 1967 1020 1968
rect 1102 1972 1108 1973
rect 1102 1968 1103 1972
rect 1107 1968 1108 1972
rect 1102 1967 1108 1968
rect 1198 1972 1204 1973
rect 1198 1968 1199 1972
rect 1203 1968 1204 1972
rect 1198 1967 1204 1968
rect 1286 1972 1292 1973
rect 1286 1968 1287 1972
rect 1291 1968 1292 1972
rect 1286 1967 1292 1968
rect 1382 1972 1388 1973
rect 1382 1968 1383 1972
rect 1387 1968 1388 1972
rect 1382 1967 1388 1968
rect 1478 1972 1484 1973
rect 1478 1968 1479 1972
rect 1483 1968 1484 1972
rect 1478 1967 1484 1968
rect 1574 1972 1580 1973
rect 1574 1968 1575 1972
rect 1579 1968 1580 1972
rect 1574 1967 1580 1968
rect 1662 1972 1668 1973
rect 1662 1968 1663 1972
rect 1667 1968 1668 1972
rect 1662 1967 1668 1968
rect 1742 1972 1748 1973
rect 1742 1968 1743 1972
rect 1747 1968 1748 1972
rect 1830 1971 1831 1975
rect 1835 1971 1836 1975
rect 1830 1970 1836 1971
rect 1742 1967 1748 1968
rect 136 1943 138 1967
rect 256 1943 258 1967
rect 376 1943 378 1967
rect 488 1943 490 1967
rect 600 1943 602 1967
rect 712 1943 714 1967
rect 816 1943 818 1967
rect 920 1943 922 1967
rect 1016 1943 1018 1967
rect 1104 1943 1106 1967
rect 1200 1943 1202 1967
rect 1288 1943 1290 1967
rect 1384 1943 1386 1967
rect 1480 1943 1482 1967
rect 1576 1943 1578 1967
rect 1664 1943 1666 1967
rect 1744 1943 1746 1967
rect 1832 1943 1834 1970
rect 1872 1951 1874 1979
rect 2078 1966 2084 1967
rect 2078 1962 2079 1966
rect 2083 1962 2084 1966
rect 2078 1961 2084 1962
rect 2214 1966 2220 1967
rect 2214 1962 2215 1966
rect 2219 1962 2220 1966
rect 2214 1961 2220 1962
rect 2366 1966 2372 1967
rect 2366 1962 2367 1966
rect 2371 1962 2372 1966
rect 2366 1961 2372 1962
rect 2526 1966 2532 1967
rect 2526 1962 2527 1966
rect 2531 1962 2532 1966
rect 2526 1961 2532 1962
rect 2686 1966 2692 1967
rect 2686 1962 2687 1966
rect 2691 1962 2692 1966
rect 2686 1961 2692 1962
rect 2854 1966 2860 1967
rect 2854 1962 2855 1966
rect 2859 1962 2860 1966
rect 2854 1961 2860 1962
rect 3022 1966 3028 1967
rect 3022 1962 3023 1966
rect 3027 1962 3028 1966
rect 3022 1961 3028 1962
rect 3190 1966 3196 1967
rect 3190 1962 3191 1966
rect 3195 1962 3196 1966
rect 3190 1961 3196 1962
rect 3358 1966 3364 1967
rect 3358 1962 3359 1966
rect 3363 1962 3364 1966
rect 3358 1961 3364 1962
rect 3510 1966 3516 1967
rect 3510 1962 3511 1966
rect 3515 1962 3516 1966
rect 3510 1961 3516 1962
rect 2080 1951 2082 1961
rect 2216 1951 2218 1961
rect 2368 1951 2370 1961
rect 2528 1951 2530 1961
rect 2688 1951 2690 1961
rect 2856 1951 2858 1961
rect 3024 1951 3026 1961
rect 3192 1951 3194 1961
rect 3360 1951 3362 1961
rect 3512 1951 3514 1961
rect 3592 1951 3594 1979
rect 1871 1950 1875 1951
rect 1871 1945 1875 1946
rect 1903 1950 1907 1951
rect 1903 1945 1907 1946
rect 2007 1950 2011 1951
rect 2007 1945 2011 1946
rect 2079 1950 2083 1951
rect 2079 1945 2083 1946
rect 2135 1950 2139 1951
rect 2135 1945 2139 1946
rect 2215 1950 2219 1951
rect 2215 1945 2219 1946
rect 2255 1950 2259 1951
rect 2255 1945 2259 1946
rect 2367 1950 2371 1951
rect 2367 1945 2371 1946
rect 2375 1950 2379 1951
rect 2375 1945 2379 1946
rect 2487 1950 2491 1951
rect 2487 1945 2491 1946
rect 2527 1950 2531 1951
rect 2527 1945 2531 1946
rect 2599 1950 2603 1951
rect 2599 1945 2603 1946
rect 2687 1950 2691 1951
rect 2687 1945 2691 1946
rect 2719 1950 2723 1951
rect 2719 1945 2723 1946
rect 2839 1950 2843 1951
rect 2839 1945 2843 1946
rect 2855 1950 2859 1951
rect 2855 1945 2859 1946
rect 3023 1950 3027 1951
rect 3023 1945 3027 1946
rect 3191 1950 3195 1951
rect 3191 1945 3195 1946
rect 3359 1950 3363 1951
rect 3359 1945 3363 1946
rect 3511 1950 3515 1951
rect 3511 1945 3515 1946
rect 3591 1950 3595 1951
rect 3591 1945 3595 1946
rect 111 1942 115 1943
rect 111 1937 115 1938
rect 135 1942 139 1943
rect 135 1937 139 1938
rect 167 1942 171 1943
rect 167 1937 171 1938
rect 255 1942 259 1943
rect 255 1937 259 1938
rect 327 1942 331 1943
rect 327 1937 331 1938
rect 375 1942 379 1943
rect 375 1937 379 1938
rect 487 1942 491 1943
rect 487 1937 491 1938
rect 599 1942 603 1943
rect 599 1937 603 1938
rect 647 1942 651 1943
rect 647 1937 651 1938
rect 711 1942 715 1943
rect 711 1937 715 1938
rect 799 1942 803 1943
rect 799 1937 803 1938
rect 815 1942 819 1943
rect 815 1937 819 1938
rect 919 1942 923 1943
rect 919 1937 923 1938
rect 943 1942 947 1943
rect 943 1937 947 1938
rect 1015 1942 1019 1943
rect 1015 1937 1019 1938
rect 1079 1942 1083 1943
rect 1079 1937 1083 1938
rect 1103 1942 1107 1943
rect 1103 1937 1107 1938
rect 1199 1942 1203 1943
rect 1199 1937 1203 1938
rect 1215 1942 1219 1943
rect 1215 1937 1219 1938
rect 1287 1942 1291 1943
rect 1287 1937 1291 1938
rect 1351 1942 1355 1943
rect 1351 1937 1355 1938
rect 1383 1942 1387 1943
rect 1383 1937 1387 1938
rect 1479 1942 1483 1943
rect 1479 1937 1483 1938
rect 1487 1942 1491 1943
rect 1487 1937 1491 1938
rect 1575 1942 1579 1943
rect 1575 1937 1579 1938
rect 1623 1942 1627 1943
rect 1623 1937 1627 1938
rect 1663 1942 1667 1943
rect 1663 1937 1667 1938
rect 1743 1942 1747 1943
rect 1743 1937 1747 1938
rect 1831 1942 1835 1943
rect 1831 1937 1835 1938
rect 112 1918 114 1937
rect 168 1921 170 1937
rect 328 1921 330 1937
rect 488 1921 490 1937
rect 648 1921 650 1937
rect 800 1921 802 1937
rect 944 1921 946 1937
rect 1080 1921 1082 1937
rect 1216 1921 1218 1937
rect 1352 1921 1354 1937
rect 1488 1921 1490 1937
rect 1624 1921 1626 1937
rect 1744 1921 1746 1937
rect 166 1920 172 1921
rect 110 1917 116 1918
rect 110 1913 111 1917
rect 115 1913 116 1917
rect 166 1916 167 1920
rect 171 1916 172 1920
rect 166 1915 172 1916
rect 326 1920 332 1921
rect 326 1916 327 1920
rect 331 1916 332 1920
rect 326 1915 332 1916
rect 486 1920 492 1921
rect 486 1916 487 1920
rect 491 1916 492 1920
rect 486 1915 492 1916
rect 646 1920 652 1921
rect 646 1916 647 1920
rect 651 1916 652 1920
rect 646 1915 652 1916
rect 798 1920 804 1921
rect 798 1916 799 1920
rect 803 1916 804 1920
rect 798 1915 804 1916
rect 942 1920 948 1921
rect 942 1916 943 1920
rect 947 1916 948 1920
rect 942 1915 948 1916
rect 1078 1920 1084 1921
rect 1078 1916 1079 1920
rect 1083 1916 1084 1920
rect 1078 1915 1084 1916
rect 1214 1920 1220 1921
rect 1214 1916 1215 1920
rect 1219 1916 1220 1920
rect 1214 1915 1220 1916
rect 1350 1920 1356 1921
rect 1350 1916 1351 1920
rect 1355 1916 1356 1920
rect 1350 1915 1356 1916
rect 1486 1920 1492 1921
rect 1486 1916 1487 1920
rect 1491 1916 1492 1920
rect 1486 1915 1492 1916
rect 1622 1920 1628 1921
rect 1622 1916 1623 1920
rect 1627 1916 1628 1920
rect 1622 1915 1628 1916
rect 1742 1920 1748 1921
rect 1742 1916 1743 1920
rect 1747 1916 1748 1920
rect 1832 1918 1834 1937
rect 1742 1915 1748 1916
rect 1830 1917 1836 1918
rect 1872 1917 1874 1945
rect 1904 1935 1906 1945
rect 2008 1935 2010 1945
rect 2136 1935 2138 1945
rect 2256 1935 2258 1945
rect 2376 1935 2378 1945
rect 2488 1935 2490 1945
rect 2600 1935 2602 1945
rect 2720 1935 2722 1945
rect 2840 1935 2842 1945
rect 1902 1934 1908 1935
rect 1902 1930 1903 1934
rect 1907 1930 1908 1934
rect 1902 1929 1908 1930
rect 2006 1934 2012 1935
rect 2006 1930 2007 1934
rect 2011 1930 2012 1934
rect 2006 1929 2012 1930
rect 2134 1934 2140 1935
rect 2134 1930 2135 1934
rect 2139 1930 2140 1934
rect 2134 1929 2140 1930
rect 2254 1934 2260 1935
rect 2254 1930 2255 1934
rect 2259 1930 2260 1934
rect 2254 1929 2260 1930
rect 2374 1934 2380 1935
rect 2374 1930 2375 1934
rect 2379 1930 2380 1934
rect 2374 1929 2380 1930
rect 2486 1934 2492 1935
rect 2486 1930 2487 1934
rect 2491 1930 2492 1934
rect 2486 1929 2492 1930
rect 2598 1934 2604 1935
rect 2598 1930 2599 1934
rect 2603 1930 2604 1934
rect 2598 1929 2604 1930
rect 2718 1934 2724 1935
rect 2718 1930 2719 1934
rect 2723 1930 2724 1934
rect 2718 1929 2724 1930
rect 2838 1934 2844 1935
rect 2838 1930 2839 1934
rect 2843 1930 2844 1934
rect 2838 1929 2844 1930
rect 3592 1917 3594 1945
rect 110 1912 116 1913
rect 1830 1913 1831 1917
rect 1835 1913 1836 1917
rect 1830 1912 1836 1913
rect 1870 1916 1876 1917
rect 1870 1912 1871 1916
rect 1875 1912 1876 1916
rect 1870 1911 1876 1912
rect 3590 1916 3596 1917
rect 3590 1912 3591 1916
rect 3595 1912 3596 1916
rect 3590 1911 3596 1912
rect 110 1900 116 1901
rect 110 1896 111 1900
rect 115 1896 116 1900
rect 110 1895 116 1896
rect 1830 1900 1836 1901
rect 1830 1896 1831 1900
rect 1835 1896 1836 1900
rect 1830 1895 1836 1896
rect 1870 1899 1876 1900
rect 1870 1895 1871 1899
rect 1875 1895 1876 1899
rect 3590 1899 3596 1900
rect 112 1867 114 1895
rect 174 1882 180 1883
rect 174 1878 175 1882
rect 179 1878 180 1882
rect 174 1877 180 1878
rect 334 1882 340 1883
rect 334 1878 335 1882
rect 339 1878 340 1882
rect 334 1877 340 1878
rect 494 1882 500 1883
rect 494 1878 495 1882
rect 499 1878 500 1882
rect 494 1877 500 1878
rect 654 1882 660 1883
rect 654 1878 655 1882
rect 659 1878 660 1882
rect 654 1877 660 1878
rect 806 1882 812 1883
rect 806 1878 807 1882
rect 811 1878 812 1882
rect 806 1877 812 1878
rect 950 1882 956 1883
rect 950 1878 951 1882
rect 955 1878 956 1882
rect 950 1877 956 1878
rect 1086 1882 1092 1883
rect 1086 1878 1087 1882
rect 1091 1878 1092 1882
rect 1086 1877 1092 1878
rect 1222 1882 1228 1883
rect 1222 1878 1223 1882
rect 1227 1878 1228 1882
rect 1222 1877 1228 1878
rect 1358 1882 1364 1883
rect 1358 1878 1359 1882
rect 1363 1878 1364 1882
rect 1358 1877 1364 1878
rect 1494 1882 1500 1883
rect 1494 1878 1495 1882
rect 1499 1878 1500 1882
rect 1494 1877 1500 1878
rect 1630 1882 1636 1883
rect 1630 1878 1631 1882
rect 1635 1878 1636 1882
rect 1630 1877 1636 1878
rect 1750 1882 1756 1883
rect 1750 1878 1751 1882
rect 1755 1878 1756 1882
rect 1750 1877 1756 1878
rect 176 1867 178 1877
rect 336 1867 338 1877
rect 496 1867 498 1877
rect 656 1867 658 1877
rect 808 1867 810 1877
rect 952 1867 954 1877
rect 1088 1867 1090 1877
rect 1224 1867 1226 1877
rect 1360 1867 1362 1877
rect 1496 1867 1498 1877
rect 1632 1867 1634 1877
rect 1752 1867 1754 1877
rect 1832 1867 1834 1895
rect 1870 1894 1876 1895
rect 1894 1896 1900 1897
rect 1872 1875 1874 1894
rect 1894 1892 1895 1896
rect 1899 1892 1900 1896
rect 1894 1891 1900 1892
rect 1998 1896 2004 1897
rect 1998 1892 1999 1896
rect 2003 1892 2004 1896
rect 1998 1891 2004 1892
rect 2126 1896 2132 1897
rect 2126 1892 2127 1896
rect 2131 1892 2132 1896
rect 2126 1891 2132 1892
rect 2246 1896 2252 1897
rect 2246 1892 2247 1896
rect 2251 1892 2252 1896
rect 2246 1891 2252 1892
rect 2366 1896 2372 1897
rect 2366 1892 2367 1896
rect 2371 1892 2372 1896
rect 2366 1891 2372 1892
rect 2478 1896 2484 1897
rect 2478 1892 2479 1896
rect 2483 1892 2484 1896
rect 2478 1891 2484 1892
rect 2590 1896 2596 1897
rect 2590 1892 2591 1896
rect 2595 1892 2596 1896
rect 2590 1891 2596 1892
rect 2710 1896 2716 1897
rect 2710 1892 2711 1896
rect 2715 1892 2716 1896
rect 2710 1891 2716 1892
rect 2830 1896 2836 1897
rect 2830 1892 2831 1896
rect 2835 1892 2836 1896
rect 3590 1895 3591 1899
rect 3595 1895 3596 1899
rect 3590 1894 3596 1895
rect 2830 1891 2836 1892
rect 1896 1875 1898 1891
rect 2000 1875 2002 1891
rect 2128 1875 2130 1891
rect 2248 1875 2250 1891
rect 2368 1875 2370 1891
rect 2480 1875 2482 1891
rect 2592 1875 2594 1891
rect 2712 1875 2714 1891
rect 2832 1875 2834 1891
rect 3592 1875 3594 1894
rect 1871 1874 1875 1875
rect 1871 1869 1875 1870
rect 1895 1874 1899 1875
rect 1895 1869 1899 1870
rect 1991 1874 1995 1875
rect 1991 1869 1995 1870
rect 1999 1874 2003 1875
rect 1999 1869 2003 1870
rect 2119 1874 2123 1875
rect 2119 1869 2123 1870
rect 2127 1874 2131 1875
rect 2127 1869 2131 1870
rect 2247 1874 2251 1875
rect 2247 1869 2251 1870
rect 2367 1874 2371 1875
rect 2367 1869 2371 1870
rect 2383 1874 2387 1875
rect 2383 1869 2387 1870
rect 2479 1874 2483 1875
rect 2479 1869 2483 1870
rect 2519 1874 2523 1875
rect 2519 1869 2523 1870
rect 2591 1874 2595 1875
rect 2591 1869 2595 1870
rect 2655 1874 2659 1875
rect 2655 1869 2659 1870
rect 2711 1874 2715 1875
rect 2711 1869 2715 1870
rect 2807 1874 2811 1875
rect 2807 1869 2811 1870
rect 2831 1874 2835 1875
rect 2831 1869 2835 1870
rect 2975 1874 2979 1875
rect 2975 1869 2979 1870
rect 3151 1874 3155 1875
rect 3151 1869 3155 1870
rect 3335 1874 3339 1875
rect 3335 1869 3339 1870
rect 3503 1874 3507 1875
rect 3503 1869 3507 1870
rect 3591 1874 3595 1875
rect 3591 1869 3595 1870
rect 111 1866 115 1867
rect 111 1861 115 1862
rect 159 1866 163 1867
rect 159 1861 163 1862
rect 175 1866 179 1867
rect 175 1861 179 1862
rect 303 1866 307 1867
rect 303 1861 307 1862
rect 335 1866 339 1867
rect 335 1861 339 1862
rect 447 1866 451 1867
rect 447 1861 451 1862
rect 495 1866 499 1867
rect 495 1861 499 1862
rect 599 1866 603 1867
rect 599 1861 603 1862
rect 655 1866 659 1867
rect 655 1861 659 1862
rect 751 1866 755 1867
rect 751 1861 755 1862
rect 807 1866 811 1867
rect 807 1861 811 1862
rect 903 1866 907 1867
rect 903 1861 907 1862
rect 951 1866 955 1867
rect 951 1861 955 1862
rect 1055 1866 1059 1867
rect 1055 1861 1059 1862
rect 1087 1866 1091 1867
rect 1087 1861 1091 1862
rect 1207 1866 1211 1867
rect 1207 1861 1211 1862
rect 1223 1866 1227 1867
rect 1223 1861 1227 1862
rect 1351 1866 1355 1867
rect 1351 1861 1355 1862
rect 1359 1866 1363 1867
rect 1359 1861 1363 1862
rect 1487 1866 1491 1867
rect 1487 1861 1491 1862
rect 1495 1866 1499 1867
rect 1495 1861 1499 1862
rect 1631 1866 1635 1867
rect 1631 1861 1635 1862
rect 1751 1866 1755 1867
rect 1751 1861 1755 1862
rect 1831 1866 1835 1867
rect 1831 1861 1835 1862
rect 112 1833 114 1861
rect 160 1851 162 1861
rect 304 1851 306 1861
rect 448 1851 450 1861
rect 600 1851 602 1861
rect 752 1851 754 1861
rect 904 1851 906 1861
rect 1056 1851 1058 1861
rect 1208 1851 1210 1861
rect 1352 1851 1354 1861
rect 1488 1851 1490 1861
rect 1632 1851 1634 1861
rect 1752 1851 1754 1861
rect 158 1850 164 1851
rect 158 1846 159 1850
rect 163 1846 164 1850
rect 158 1845 164 1846
rect 302 1850 308 1851
rect 302 1846 303 1850
rect 307 1846 308 1850
rect 302 1845 308 1846
rect 446 1850 452 1851
rect 446 1846 447 1850
rect 451 1846 452 1850
rect 446 1845 452 1846
rect 598 1850 604 1851
rect 598 1846 599 1850
rect 603 1846 604 1850
rect 598 1845 604 1846
rect 750 1850 756 1851
rect 750 1846 751 1850
rect 755 1846 756 1850
rect 750 1845 756 1846
rect 902 1850 908 1851
rect 902 1846 903 1850
rect 907 1846 908 1850
rect 902 1845 908 1846
rect 1054 1850 1060 1851
rect 1054 1846 1055 1850
rect 1059 1846 1060 1850
rect 1054 1845 1060 1846
rect 1206 1850 1212 1851
rect 1206 1846 1207 1850
rect 1211 1846 1212 1850
rect 1206 1845 1212 1846
rect 1350 1850 1356 1851
rect 1350 1846 1351 1850
rect 1355 1846 1356 1850
rect 1350 1845 1356 1846
rect 1486 1850 1492 1851
rect 1486 1846 1487 1850
rect 1491 1846 1492 1850
rect 1486 1845 1492 1846
rect 1630 1850 1636 1851
rect 1630 1846 1631 1850
rect 1635 1846 1636 1850
rect 1630 1845 1636 1846
rect 1750 1850 1756 1851
rect 1750 1846 1751 1850
rect 1755 1846 1756 1850
rect 1750 1845 1756 1846
rect 1832 1833 1834 1861
rect 1872 1850 1874 1869
rect 1896 1853 1898 1869
rect 1992 1853 1994 1869
rect 2120 1853 2122 1869
rect 2248 1853 2250 1869
rect 2384 1853 2386 1869
rect 2520 1853 2522 1869
rect 2656 1853 2658 1869
rect 2808 1853 2810 1869
rect 2976 1853 2978 1869
rect 3152 1853 3154 1869
rect 3336 1853 3338 1869
rect 3504 1853 3506 1869
rect 1894 1852 1900 1853
rect 1870 1849 1876 1850
rect 1870 1845 1871 1849
rect 1875 1845 1876 1849
rect 1894 1848 1895 1852
rect 1899 1848 1900 1852
rect 1894 1847 1900 1848
rect 1990 1852 1996 1853
rect 1990 1848 1991 1852
rect 1995 1848 1996 1852
rect 1990 1847 1996 1848
rect 2118 1852 2124 1853
rect 2118 1848 2119 1852
rect 2123 1848 2124 1852
rect 2118 1847 2124 1848
rect 2246 1852 2252 1853
rect 2246 1848 2247 1852
rect 2251 1848 2252 1852
rect 2246 1847 2252 1848
rect 2382 1852 2388 1853
rect 2382 1848 2383 1852
rect 2387 1848 2388 1852
rect 2382 1847 2388 1848
rect 2518 1852 2524 1853
rect 2518 1848 2519 1852
rect 2523 1848 2524 1852
rect 2518 1847 2524 1848
rect 2654 1852 2660 1853
rect 2654 1848 2655 1852
rect 2659 1848 2660 1852
rect 2654 1847 2660 1848
rect 2806 1852 2812 1853
rect 2806 1848 2807 1852
rect 2811 1848 2812 1852
rect 2806 1847 2812 1848
rect 2974 1852 2980 1853
rect 2974 1848 2975 1852
rect 2979 1848 2980 1852
rect 2974 1847 2980 1848
rect 3150 1852 3156 1853
rect 3150 1848 3151 1852
rect 3155 1848 3156 1852
rect 3150 1847 3156 1848
rect 3334 1852 3340 1853
rect 3334 1848 3335 1852
rect 3339 1848 3340 1852
rect 3334 1847 3340 1848
rect 3502 1852 3508 1853
rect 3502 1848 3503 1852
rect 3507 1848 3508 1852
rect 3592 1850 3594 1869
rect 3502 1847 3508 1848
rect 3590 1849 3596 1850
rect 1870 1844 1876 1845
rect 3590 1845 3591 1849
rect 3595 1845 3596 1849
rect 3590 1844 3596 1845
rect 110 1832 116 1833
rect 110 1828 111 1832
rect 115 1828 116 1832
rect 110 1827 116 1828
rect 1830 1832 1836 1833
rect 1830 1828 1831 1832
rect 1835 1828 1836 1832
rect 1830 1827 1836 1828
rect 1870 1832 1876 1833
rect 1870 1828 1871 1832
rect 1875 1828 1876 1832
rect 1870 1827 1876 1828
rect 3590 1832 3596 1833
rect 3590 1828 3591 1832
rect 3595 1828 3596 1832
rect 3590 1827 3596 1828
rect 110 1815 116 1816
rect 110 1811 111 1815
rect 115 1811 116 1815
rect 1830 1815 1836 1816
rect 110 1810 116 1811
rect 150 1812 156 1813
rect 112 1787 114 1810
rect 150 1808 151 1812
rect 155 1808 156 1812
rect 150 1807 156 1808
rect 294 1812 300 1813
rect 294 1808 295 1812
rect 299 1808 300 1812
rect 294 1807 300 1808
rect 438 1812 444 1813
rect 438 1808 439 1812
rect 443 1808 444 1812
rect 438 1807 444 1808
rect 590 1812 596 1813
rect 590 1808 591 1812
rect 595 1808 596 1812
rect 590 1807 596 1808
rect 742 1812 748 1813
rect 742 1808 743 1812
rect 747 1808 748 1812
rect 742 1807 748 1808
rect 894 1812 900 1813
rect 894 1808 895 1812
rect 899 1808 900 1812
rect 894 1807 900 1808
rect 1046 1812 1052 1813
rect 1046 1808 1047 1812
rect 1051 1808 1052 1812
rect 1046 1807 1052 1808
rect 1198 1812 1204 1813
rect 1198 1808 1199 1812
rect 1203 1808 1204 1812
rect 1198 1807 1204 1808
rect 1342 1812 1348 1813
rect 1342 1808 1343 1812
rect 1347 1808 1348 1812
rect 1342 1807 1348 1808
rect 1478 1812 1484 1813
rect 1478 1808 1479 1812
rect 1483 1808 1484 1812
rect 1478 1807 1484 1808
rect 1622 1812 1628 1813
rect 1622 1808 1623 1812
rect 1627 1808 1628 1812
rect 1622 1807 1628 1808
rect 1742 1812 1748 1813
rect 1742 1808 1743 1812
rect 1747 1808 1748 1812
rect 1830 1811 1831 1815
rect 1835 1811 1836 1815
rect 1830 1810 1836 1811
rect 1742 1807 1748 1808
rect 152 1787 154 1807
rect 296 1787 298 1807
rect 440 1787 442 1807
rect 592 1787 594 1807
rect 744 1787 746 1807
rect 896 1787 898 1807
rect 1048 1787 1050 1807
rect 1200 1787 1202 1807
rect 1344 1787 1346 1807
rect 1480 1787 1482 1807
rect 1624 1787 1626 1807
rect 1744 1787 1746 1807
rect 1832 1787 1834 1810
rect 1872 1787 1874 1827
rect 1902 1814 1908 1815
rect 1902 1810 1903 1814
rect 1907 1810 1908 1814
rect 1902 1809 1908 1810
rect 1998 1814 2004 1815
rect 1998 1810 1999 1814
rect 2003 1810 2004 1814
rect 1998 1809 2004 1810
rect 2126 1814 2132 1815
rect 2126 1810 2127 1814
rect 2131 1810 2132 1814
rect 2126 1809 2132 1810
rect 2254 1814 2260 1815
rect 2254 1810 2255 1814
rect 2259 1810 2260 1814
rect 2254 1809 2260 1810
rect 2390 1814 2396 1815
rect 2390 1810 2391 1814
rect 2395 1810 2396 1814
rect 2390 1809 2396 1810
rect 2526 1814 2532 1815
rect 2526 1810 2527 1814
rect 2531 1810 2532 1814
rect 2526 1809 2532 1810
rect 2662 1814 2668 1815
rect 2662 1810 2663 1814
rect 2667 1810 2668 1814
rect 2662 1809 2668 1810
rect 2814 1814 2820 1815
rect 2814 1810 2815 1814
rect 2819 1810 2820 1814
rect 2814 1809 2820 1810
rect 2982 1814 2988 1815
rect 2982 1810 2983 1814
rect 2987 1810 2988 1814
rect 2982 1809 2988 1810
rect 3158 1814 3164 1815
rect 3158 1810 3159 1814
rect 3163 1810 3164 1814
rect 3158 1809 3164 1810
rect 3342 1814 3348 1815
rect 3342 1810 3343 1814
rect 3347 1810 3348 1814
rect 3342 1809 3348 1810
rect 3510 1814 3516 1815
rect 3510 1810 3511 1814
rect 3515 1810 3516 1814
rect 3510 1809 3516 1810
rect 1904 1787 1906 1809
rect 2000 1787 2002 1809
rect 2128 1787 2130 1809
rect 2256 1787 2258 1809
rect 2392 1787 2394 1809
rect 2528 1787 2530 1809
rect 2664 1787 2666 1809
rect 2816 1787 2818 1809
rect 2984 1787 2986 1809
rect 3160 1787 3162 1809
rect 3344 1787 3346 1809
rect 3512 1787 3514 1809
rect 3592 1787 3594 1827
rect 111 1786 115 1787
rect 111 1781 115 1782
rect 151 1786 155 1787
rect 151 1781 155 1782
rect 247 1786 251 1787
rect 247 1781 251 1782
rect 295 1786 299 1787
rect 295 1781 299 1782
rect 423 1786 427 1787
rect 423 1781 427 1782
rect 439 1786 443 1787
rect 439 1781 443 1782
rect 591 1786 595 1787
rect 591 1781 595 1782
rect 743 1786 747 1787
rect 743 1781 747 1782
rect 751 1786 755 1787
rect 751 1781 755 1782
rect 895 1786 899 1787
rect 895 1781 899 1782
rect 1023 1786 1027 1787
rect 1023 1781 1027 1782
rect 1047 1786 1051 1787
rect 1047 1781 1051 1782
rect 1143 1786 1147 1787
rect 1143 1781 1147 1782
rect 1199 1786 1203 1787
rect 1199 1781 1203 1782
rect 1263 1786 1267 1787
rect 1263 1781 1267 1782
rect 1343 1786 1347 1787
rect 1343 1781 1347 1782
rect 1391 1786 1395 1787
rect 1391 1781 1395 1782
rect 1479 1786 1483 1787
rect 1479 1781 1483 1782
rect 1623 1786 1627 1787
rect 1623 1781 1627 1782
rect 1743 1786 1747 1787
rect 1743 1781 1747 1782
rect 1831 1786 1835 1787
rect 1831 1781 1835 1782
rect 1871 1786 1875 1787
rect 1871 1781 1875 1782
rect 1903 1786 1907 1787
rect 1903 1781 1907 1782
rect 1999 1786 2003 1787
rect 1999 1781 2003 1782
rect 2031 1786 2035 1787
rect 2031 1781 2035 1782
rect 2127 1786 2131 1787
rect 2127 1781 2131 1782
rect 2191 1786 2195 1787
rect 2191 1781 2195 1782
rect 2255 1786 2259 1787
rect 2255 1781 2259 1782
rect 2359 1786 2363 1787
rect 2359 1781 2363 1782
rect 2391 1786 2395 1787
rect 2391 1781 2395 1782
rect 2527 1786 2531 1787
rect 2527 1781 2531 1782
rect 2663 1786 2667 1787
rect 2663 1781 2667 1782
rect 2687 1786 2691 1787
rect 2687 1781 2691 1782
rect 2815 1786 2819 1787
rect 2815 1781 2819 1782
rect 2839 1786 2843 1787
rect 2839 1781 2843 1782
rect 2983 1786 2987 1787
rect 2983 1781 2987 1782
rect 3119 1786 3123 1787
rect 3119 1781 3123 1782
rect 3159 1786 3163 1787
rect 3159 1781 3163 1782
rect 3255 1786 3259 1787
rect 3255 1781 3259 1782
rect 3343 1786 3347 1787
rect 3343 1781 3347 1782
rect 3391 1786 3395 1787
rect 3391 1781 3395 1782
rect 3511 1786 3515 1787
rect 3511 1781 3515 1782
rect 3591 1786 3595 1787
rect 3591 1781 3595 1782
rect 112 1762 114 1781
rect 248 1765 250 1781
rect 424 1765 426 1781
rect 592 1765 594 1781
rect 752 1765 754 1781
rect 896 1765 898 1781
rect 1024 1765 1026 1781
rect 1144 1765 1146 1781
rect 1264 1765 1266 1781
rect 1392 1765 1394 1781
rect 246 1764 252 1765
rect 110 1761 116 1762
rect 110 1757 111 1761
rect 115 1757 116 1761
rect 246 1760 247 1764
rect 251 1760 252 1764
rect 246 1759 252 1760
rect 422 1764 428 1765
rect 422 1760 423 1764
rect 427 1760 428 1764
rect 422 1759 428 1760
rect 590 1764 596 1765
rect 590 1760 591 1764
rect 595 1760 596 1764
rect 590 1759 596 1760
rect 750 1764 756 1765
rect 750 1760 751 1764
rect 755 1760 756 1764
rect 750 1759 756 1760
rect 894 1764 900 1765
rect 894 1760 895 1764
rect 899 1760 900 1764
rect 894 1759 900 1760
rect 1022 1764 1028 1765
rect 1022 1760 1023 1764
rect 1027 1760 1028 1764
rect 1022 1759 1028 1760
rect 1142 1764 1148 1765
rect 1142 1760 1143 1764
rect 1147 1760 1148 1764
rect 1142 1759 1148 1760
rect 1262 1764 1268 1765
rect 1262 1760 1263 1764
rect 1267 1760 1268 1764
rect 1262 1759 1268 1760
rect 1390 1764 1396 1765
rect 1390 1760 1391 1764
rect 1395 1760 1396 1764
rect 1832 1762 1834 1781
rect 1390 1759 1396 1760
rect 1830 1761 1836 1762
rect 110 1756 116 1757
rect 1830 1757 1831 1761
rect 1835 1757 1836 1761
rect 1830 1756 1836 1757
rect 1872 1753 1874 1781
rect 1904 1771 1906 1781
rect 2032 1771 2034 1781
rect 2192 1771 2194 1781
rect 2360 1771 2362 1781
rect 2528 1771 2530 1781
rect 2688 1771 2690 1781
rect 2840 1771 2842 1781
rect 2984 1771 2986 1781
rect 3120 1771 3122 1781
rect 3256 1771 3258 1781
rect 3392 1771 3394 1781
rect 3512 1771 3514 1781
rect 1902 1770 1908 1771
rect 1902 1766 1903 1770
rect 1907 1766 1908 1770
rect 1902 1765 1908 1766
rect 2030 1770 2036 1771
rect 2030 1766 2031 1770
rect 2035 1766 2036 1770
rect 2030 1765 2036 1766
rect 2190 1770 2196 1771
rect 2190 1766 2191 1770
rect 2195 1766 2196 1770
rect 2190 1765 2196 1766
rect 2358 1770 2364 1771
rect 2358 1766 2359 1770
rect 2363 1766 2364 1770
rect 2358 1765 2364 1766
rect 2526 1770 2532 1771
rect 2526 1766 2527 1770
rect 2531 1766 2532 1770
rect 2526 1765 2532 1766
rect 2686 1770 2692 1771
rect 2686 1766 2687 1770
rect 2691 1766 2692 1770
rect 2686 1765 2692 1766
rect 2838 1770 2844 1771
rect 2838 1766 2839 1770
rect 2843 1766 2844 1770
rect 2838 1765 2844 1766
rect 2982 1770 2988 1771
rect 2982 1766 2983 1770
rect 2987 1766 2988 1770
rect 2982 1765 2988 1766
rect 3118 1770 3124 1771
rect 3118 1766 3119 1770
rect 3123 1766 3124 1770
rect 3118 1765 3124 1766
rect 3254 1770 3260 1771
rect 3254 1766 3255 1770
rect 3259 1766 3260 1770
rect 3254 1765 3260 1766
rect 3390 1770 3396 1771
rect 3390 1766 3391 1770
rect 3395 1766 3396 1770
rect 3390 1765 3396 1766
rect 3510 1770 3516 1771
rect 3510 1766 3511 1770
rect 3515 1766 3516 1770
rect 3510 1765 3516 1766
rect 3592 1753 3594 1781
rect 1870 1752 1876 1753
rect 1870 1748 1871 1752
rect 1875 1748 1876 1752
rect 1870 1747 1876 1748
rect 3590 1752 3596 1753
rect 3590 1748 3591 1752
rect 3595 1748 3596 1752
rect 3590 1747 3596 1748
rect 110 1744 116 1745
rect 110 1740 111 1744
rect 115 1740 116 1744
rect 110 1739 116 1740
rect 1830 1744 1836 1745
rect 1830 1740 1831 1744
rect 1835 1740 1836 1744
rect 1830 1739 1836 1740
rect 112 1707 114 1739
rect 254 1726 260 1727
rect 254 1722 255 1726
rect 259 1722 260 1726
rect 254 1721 260 1722
rect 430 1726 436 1727
rect 430 1722 431 1726
rect 435 1722 436 1726
rect 430 1721 436 1722
rect 598 1726 604 1727
rect 598 1722 599 1726
rect 603 1722 604 1726
rect 598 1721 604 1722
rect 758 1726 764 1727
rect 758 1722 759 1726
rect 763 1722 764 1726
rect 758 1721 764 1722
rect 902 1726 908 1727
rect 902 1722 903 1726
rect 907 1722 908 1726
rect 902 1721 908 1722
rect 1030 1726 1036 1727
rect 1030 1722 1031 1726
rect 1035 1722 1036 1726
rect 1030 1721 1036 1722
rect 1150 1726 1156 1727
rect 1150 1722 1151 1726
rect 1155 1722 1156 1726
rect 1150 1721 1156 1722
rect 1270 1726 1276 1727
rect 1270 1722 1271 1726
rect 1275 1722 1276 1726
rect 1270 1721 1276 1722
rect 1398 1726 1404 1727
rect 1398 1722 1399 1726
rect 1403 1722 1404 1726
rect 1398 1721 1404 1722
rect 256 1707 258 1721
rect 432 1707 434 1721
rect 600 1707 602 1721
rect 760 1707 762 1721
rect 904 1707 906 1721
rect 1032 1707 1034 1721
rect 1152 1707 1154 1721
rect 1272 1707 1274 1721
rect 1400 1707 1402 1721
rect 1832 1707 1834 1739
rect 1870 1735 1876 1736
rect 1870 1731 1871 1735
rect 1875 1731 1876 1735
rect 3590 1735 3596 1736
rect 1870 1730 1876 1731
rect 1894 1732 1900 1733
rect 1872 1707 1874 1730
rect 1894 1728 1895 1732
rect 1899 1728 1900 1732
rect 1894 1727 1900 1728
rect 2022 1732 2028 1733
rect 2022 1728 2023 1732
rect 2027 1728 2028 1732
rect 2022 1727 2028 1728
rect 2182 1732 2188 1733
rect 2182 1728 2183 1732
rect 2187 1728 2188 1732
rect 2182 1727 2188 1728
rect 2350 1732 2356 1733
rect 2350 1728 2351 1732
rect 2355 1728 2356 1732
rect 2350 1727 2356 1728
rect 2518 1732 2524 1733
rect 2518 1728 2519 1732
rect 2523 1728 2524 1732
rect 2518 1727 2524 1728
rect 2678 1732 2684 1733
rect 2678 1728 2679 1732
rect 2683 1728 2684 1732
rect 2678 1727 2684 1728
rect 2830 1732 2836 1733
rect 2830 1728 2831 1732
rect 2835 1728 2836 1732
rect 2830 1727 2836 1728
rect 2974 1732 2980 1733
rect 2974 1728 2975 1732
rect 2979 1728 2980 1732
rect 2974 1727 2980 1728
rect 3110 1732 3116 1733
rect 3110 1728 3111 1732
rect 3115 1728 3116 1732
rect 3110 1727 3116 1728
rect 3246 1732 3252 1733
rect 3246 1728 3247 1732
rect 3251 1728 3252 1732
rect 3246 1727 3252 1728
rect 3382 1732 3388 1733
rect 3382 1728 3383 1732
rect 3387 1728 3388 1732
rect 3382 1727 3388 1728
rect 3502 1732 3508 1733
rect 3502 1728 3503 1732
rect 3507 1728 3508 1732
rect 3590 1731 3591 1735
rect 3595 1731 3596 1735
rect 3590 1730 3596 1731
rect 3502 1727 3508 1728
rect 1896 1707 1898 1727
rect 2024 1707 2026 1727
rect 2184 1707 2186 1727
rect 2352 1707 2354 1727
rect 2520 1707 2522 1727
rect 2680 1707 2682 1727
rect 2832 1707 2834 1727
rect 2976 1707 2978 1727
rect 3112 1707 3114 1727
rect 3248 1707 3250 1727
rect 3384 1707 3386 1727
rect 3504 1707 3506 1727
rect 3592 1707 3594 1730
rect 111 1706 115 1707
rect 111 1701 115 1702
rect 191 1706 195 1707
rect 191 1701 195 1702
rect 255 1706 259 1707
rect 255 1701 259 1702
rect 311 1706 315 1707
rect 311 1701 315 1702
rect 431 1706 435 1707
rect 431 1701 435 1702
rect 447 1706 451 1707
rect 447 1701 451 1702
rect 591 1706 595 1707
rect 591 1701 595 1702
rect 599 1706 603 1707
rect 599 1701 603 1702
rect 743 1706 747 1707
rect 743 1701 747 1702
rect 759 1706 763 1707
rect 759 1701 763 1702
rect 895 1706 899 1707
rect 895 1701 899 1702
rect 903 1706 907 1707
rect 903 1701 907 1702
rect 1031 1706 1035 1707
rect 1031 1701 1035 1702
rect 1039 1706 1043 1707
rect 1039 1701 1043 1702
rect 1151 1706 1155 1707
rect 1151 1701 1155 1702
rect 1183 1706 1187 1707
rect 1183 1701 1187 1702
rect 1271 1706 1275 1707
rect 1271 1701 1275 1702
rect 1319 1706 1323 1707
rect 1319 1701 1323 1702
rect 1399 1706 1403 1707
rect 1399 1701 1403 1702
rect 1447 1706 1451 1707
rect 1447 1701 1451 1702
rect 1575 1706 1579 1707
rect 1575 1701 1579 1702
rect 1711 1706 1715 1707
rect 1711 1701 1715 1702
rect 1831 1706 1835 1707
rect 1831 1701 1835 1702
rect 1871 1706 1875 1707
rect 1871 1701 1875 1702
rect 1895 1706 1899 1707
rect 1895 1701 1899 1702
rect 1991 1706 1995 1707
rect 1991 1701 1995 1702
rect 2023 1706 2027 1707
rect 2023 1701 2027 1702
rect 2135 1706 2139 1707
rect 2135 1701 2139 1702
rect 2183 1706 2187 1707
rect 2183 1701 2187 1702
rect 2295 1706 2299 1707
rect 2295 1701 2299 1702
rect 2351 1706 2355 1707
rect 2351 1701 2355 1702
rect 2471 1706 2475 1707
rect 2471 1701 2475 1702
rect 2519 1706 2523 1707
rect 2519 1701 2523 1702
rect 2647 1706 2651 1707
rect 2647 1701 2651 1702
rect 2679 1706 2683 1707
rect 2679 1701 2683 1702
rect 2815 1706 2819 1707
rect 2815 1701 2819 1702
rect 2831 1706 2835 1707
rect 2831 1701 2835 1702
rect 2967 1706 2971 1707
rect 2967 1701 2971 1702
rect 2975 1706 2979 1707
rect 2975 1701 2979 1702
rect 3111 1706 3115 1707
rect 3111 1701 3115 1702
rect 3247 1706 3251 1707
rect 3247 1701 3251 1702
rect 3383 1706 3387 1707
rect 3383 1701 3387 1702
rect 3503 1706 3507 1707
rect 3503 1701 3507 1702
rect 3591 1706 3595 1707
rect 3591 1701 3595 1702
rect 112 1673 114 1701
rect 192 1691 194 1701
rect 312 1691 314 1701
rect 448 1691 450 1701
rect 592 1691 594 1701
rect 744 1691 746 1701
rect 896 1691 898 1701
rect 1040 1691 1042 1701
rect 1184 1691 1186 1701
rect 1320 1691 1322 1701
rect 1448 1691 1450 1701
rect 1576 1691 1578 1701
rect 1712 1691 1714 1701
rect 190 1690 196 1691
rect 190 1686 191 1690
rect 195 1686 196 1690
rect 190 1685 196 1686
rect 310 1690 316 1691
rect 310 1686 311 1690
rect 315 1686 316 1690
rect 310 1685 316 1686
rect 446 1690 452 1691
rect 446 1686 447 1690
rect 451 1686 452 1690
rect 446 1685 452 1686
rect 590 1690 596 1691
rect 590 1686 591 1690
rect 595 1686 596 1690
rect 590 1685 596 1686
rect 742 1690 748 1691
rect 742 1686 743 1690
rect 747 1686 748 1690
rect 742 1685 748 1686
rect 894 1690 900 1691
rect 894 1686 895 1690
rect 899 1686 900 1690
rect 894 1685 900 1686
rect 1038 1690 1044 1691
rect 1038 1686 1039 1690
rect 1043 1686 1044 1690
rect 1038 1685 1044 1686
rect 1182 1690 1188 1691
rect 1182 1686 1183 1690
rect 1187 1686 1188 1690
rect 1182 1685 1188 1686
rect 1318 1690 1324 1691
rect 1318 1686 1319 1690
rect 1323 1686 1324 1690
rect 1318 1685 1324 1686
rect 1446 1690 1452 1691
rect 1446 1686 1447 1690
rect 1451 1686 1452 1690
rect 1446 1685 1452 1686
rect 1574 1690 1580 1691
rect 1574 1686 1575 1690
rect 1579 1686 1580 1690
rect 1574 1685 1580 1686
rect 1710 1690 1716 1691
rect 1710 1686 1711 1690
rect 1715 1686 1716 1690
rect 1710 1685 1716 1686
rect 1832 1673 1834 1701
rect 1872 1682 1874 1701
rect 1896 1685 1898 1701
rect 1992 1685 1994 1701
rect 2136 1685 2138 1701
rect 2296 1685 2298 1701
rect 2472 1685 2474 1701
rect 2648 1685 2650 1701
rect 2816 1685 2818 1701
rect 2968 1685 2970 1701
rect 3112 1685 3114 1701
rect 3248 1685 3250 1701
rect 3384 1685 3386 1701
rect 3504 1685 3506 1701
rect 1894 1684 1900 1685
rect 1870 1681 1876 1682
rect 1870 1677 1871 1681
rect 1875 1677 1876 1681
rect 1894 1680 1895 1684
rect 1899 1680 1900 1684
rect 1894 1679 1900 1680
rect 1990 1684 1996 1685
rect 1990 1680 1991 1684
rect 1995 1680 1996 1684
rect 1990 1679 1996 1680
rect 2134 1684 2140 1685
rect 2134 1680 2135 1684
rect 2139 1680 2140 1684
rect 2134 1679 2140 1680
rect 2294 1684 2300 1685
rect 2294 1680 2295 1684
rect 2299 1680 2300 1684
rect 2294 1679 2300 1680
rect 2470 1684 2476 1685
rect 2470 1680 2471 1684
rect 2475 1680 2476 1684
rect 2470 1679 2476 1680
rect 2646 1684 2652 1685
rect 2646 1680 2647 1684
rect 2651 1680 2652 1684
rect 2646 1679 2652 1680
rect 2814 1684 2820 1685
rect 2814 1680 2815 1684
rect 2819 1680 2820 1684
rect 2814 1679 2820 1680
rect 2966 1684 2972 1685
rect 2966 1680 2967 1684
rect 2971 1680 2972 1684
rect 2966 1679 2972 1680
rect 3110 1684 3116 1685
rect 3110 1680 3111 1684
rect 3115 1680 3116 1684
rect 3110 1679 3116 1680
rect 3246 1684 3252 1685
rect 3246 1680 3247 1684
rect 3251 1680 3252 1684
rect 3246 1679 3252 1680
rect 3382 1684 3388 1685
rect 3382 1680 3383 1684
rect 3387 1680 3388 1684
rect 3382 1679 3388 1680
rect 3502 1684 3508 1685
rect 3502 1680 3503 1684
rect 3507 1680 3508 1684
rect 3592 1682 3594 1701
rect 3502 1679 3508 1680
rect 3590 1681 3596 1682
rect 1870 1676 1876 1677
rect 3590 1677 3591 1681
rect 3595 1677 3596 1681
rect 3590 1676 3596 1677
rect 110 1672 116 1673
rect 110 1668 111 1672
rect 115 1668 116 1672
rect 110 1667 116 1668
rect 1830 1672 1836 1673
rect 1830 1668 1831 1672
rect 1835 1668 1836 1672
rect 1830 1667 1836 1668
rect 1870 1664 1876 1665
rect 1870 1660 1871 1664
rect 1875 1660 1876 1664
rect 1870 1659 1876 1660
rect 3590 1664 3596 1665
rect 3590 1660 3591 1664
rect 3595 1660 3596 1664
rect 3590 1659 3596 1660
rect 110 1655 116 1656
rect 110 1651 111 1655
rect 115 1651 116 1655
rect 1830 1655 1836 1656
rect 110 1650 116 1651
rect 182 1652 188 1653
rect 112 1623 114 1650
rect 182 1648 183 1652
rect 187 1648 188 1652
rect 182 1647 188 1648
rect 302 1652 308 1653
rect 302 1648 303 1652
rect 307 1648 308 1652
rect 302 1647 308 1648
rect 438 1652 444 1653
rect 438 1648 439 1652
rect 443 1648 444 1652
rect 438 1647 444 1648
rect 582 1652 588 1653
rect 582 1648 583 1652
rect 587 1648 588 1652
rect 582 1647 588 1648
rect 734 1652 740 1653
rect 734 1648 735 1652
rect 739 1648 740 1652
rect 734 1647 740 1648
rect 886 1652 892 1653
rect 886 1648 887 1652
rect 891 1648 892 1652
rect 886 1647 892 1648
rect 1030 1652 1036 1653
rect 1030 1648 1031 1652
rect 1035 1648 1036 1652
rect 1030 1647 1036 1648
rect 1174 1652 1180 1653
rect 1174 1648 1175 1652
rect 1179 1648 1180 1652
rect 1174 1647 1180 1648
rect 1310 1652 1316 1653
rect 1310 1648 1311 1652
rect 1315 1648 1316 1652
rect 1310 1647 1316 1648
rect 1438 1652 1444 1653
rect 1438 1648 1439 1652
rect 1443 1648 1444 1652
rect 1438 1647 1444 1648
rect 1566 1652 1572 1653
rect 1566 1648 1567 1652
rect 1571 1648 1572 1652
rect 1566 1647 1572 1648
rect 1702 1652 1708 1653
rect 1702 1648 1703 1652
rect 1707 1648 1708 1652
rect 1830 1651 1831 1655
rect 1835 1651 1836 1655
rect 1830 1650 1836 1651
rect 1702 1647 1708 1648
rect 184 1623 186 1647
rect 304 1623 306 1647
rect 440 1623 442 1647
rect 584 1623 586 1647
rect 736 1623 738 1647
rect 888 1623 890 1647
rect 1032 1623 1034 1647
rect 1176 1623 1178 1647
rect 1312 1623 1314 1647
rect 1440 1623 1442 1647
rect 1568 1623 1570 1647
rect 1704 1623 1706 1647
rect 1832 1623 1834 1650
rect 1872 1627 1874 1659
rect 1902 1646 1908 1647
rect 1902 1642 1903 1646
rect 1907 1642 1908 1646
rect 1902 1641 1908 1642
rect 1998 1646 2004 1647
rect 1998 1642 1999 1646
rect 2003 1642 2004 1646
rect 1998 1641 2004 1642
rect 2142 1646 2148 1647
rect 2142 1642 2143 1646
rect 2147 1642 2148 1646
rect 2142 1641 2148 1642
rect 2302 1646 2308 1647
rect 2302 1642 2303 1646
rect 2307 1642 2308 1646
rect 2302 1641 2308 1642
rect 2478 1646 2484 1647
rect 2478 1642 2479 1646
rect 2483 1642 2484 1646
rect 2478 1641 2484 1642
rect 2654 1646 2660 1647
rect 2654 1642 2655 1646
rect 2659 1642 2660 1646
rect 2654 1641 2660 1642
rect 2822 1646 2828 1647
rect 2822 1642 2823 1646
rect 2827 1642 2828 1646
rect 2822 1641 2828 1642
rect 2974 1646 2980 1647
rect 2974 1642 2975 1646
rect 2979 1642 2980 1646
rect 2974 1641 2980 1642
rect 3118 1646 3124 1647
rect 3118 1642 3119 1646
rect 3123 1642 3124 1646
rect 3118 1641 3124 1642
rect 3254 1646 3260 1647
rect 3254 1642 3255 1646
rect 3259 1642 3260 1646
rect 3254 1641 3260 1642
rect 3390 1646 3396 1647
rect 3390 1642 3391 1646
rect 3395 1642 3396 1646
rect 3390 1641 3396 1642
rect 3510 1646 3516 1647
rect 3510 1642 3511 1646
rect 3515 1642 3516 1646
rect 3510 1641 3516 1642
rect 1904 1627 1906 1641
rect 2000 1627 2002 1641
rect 2144 1627 2146 1641
rect 2304 1627 2306 1641
rect 2480 1627 2482 1641
rect 2656 1627 2658 1641
rect 2824 1627 2826 1641
rect 2976 1627 2978 1641
rect 3120 1627 3122 1641
rect 3256 1627 3258 1641
rect 3392 1627 3394 1641
rect 3512 1627 3514 1641
rect 3592 1627 3594 1659
rect 1871 1626 1875 1627
rect 111 1622 115 1623
rect 111 1617 115 1618
rect 167 1622 171 1623
rect 167 1617 171 1618
rect 183 1622 187 1623
rect 183 1617 187 1618
rect 303 1622 307 1623
rect 303 1617 307 1618
rect 351 1622 355 1623
rect 351 1617 355 1618
rect 439 1622 443 1623
rect 439 1617 443 1618
rect 543 1622 547 1623
rect 543 1617 547 1618
rect 583 1622 587 1623
rect 583 1617 587 1618
rect 727 1622 731 1623
rect 727 1617 731 1618
rect 735 1622 739 1623
rect 735 1617 739 1618
rect 887 1622 891 1623
rect 887 1617 891 1618
rect 903 1622 907 1623
rect 903 1617 907 1618
rect 1031 1622 1035 1623
rect 1031 1617 1035 1618
rect 1071 1622 1075 1623
rect 1071 1617 1075 1618
rect 1175 1622 1179 1623
rect 1175 1617 1179 1618
rect 1223 1622 1227 1623
rect 1223 1617 1227 1618
rect 1311 1622 1315 1623
rect 1311 1617 1315 1618
rect 1359 1622 1363 1623
rect 1359 1617 1363 1618
rect 1439 1622 1443 1623
rect 1439 1617 1443 1618
rect 1495 1622 1499 1623
rect 1495 1617 1499 1618
rect 1567 1622 1571 1623
rect 1567 1617 1571 1618
rect 1623 1622 1627 1623
rect 1623 1617 1627 1618
rect 1703 1622 1707 1623
rect 1703 1617 1707 1618
rect 1743 1622 1747 1623
rect 1743 1617 1747 1618
rect 1831 1622 1835 1623
rect 1871 1621 1875 1622
rect 1903 1626 1907 1627
rect 1903 1621 1907 1622
rect 1975 1626 1979 1627
rect 1975 1621 1979 1622
rect 1999 1626 2003 1627
rect 1999 1621 2003 1622
rect 2095 1626 2099 1627
rect 2095 1621 2099 1622
rect 2143 1626 2147 1627
rect 2143 1621 2147 1622
rect 2231 1626 2235 1627
rect 2231 1621 2235 1622
rect 2303 1626 2307 1627
rect 2303 1621 2307 1622
rect 2367 1626 2371 1627
rect 2367 1621 2371 1622
rect 2479 1626 2483 1627
rect 2479 1621 2483 1622
rect 2503 1626 2507 1627
rect 2503 1621 2507 1622
rect 2639 1626 2643 1627
rect 2639 1621 2643 1622
rect 2655 1626 2659 1627
rect 2655 1621 2659 1622
rect 2775 1626 2779 1627
rect 2775 1621 2779 1622
rect 2823 1626 2827 1627
rect 2823 1621 2827 1622
rect 2911 1626 2915 1627
rect 2911 1621 2915 1622
rect 2975 1626 2979 1627
rect 2975 1621 2979 1622
rect 3055 1626 3059 1627
rect 3055 1621 3059 1622
rect 3119 1626 3123 1627
rect 3119 1621 3123 1622
rect 3207 1626 3211 1627
rect 3207 1621 3211 1622
rect 3255 1626 3259 1627
rect 3255 1621 3259 1622
rect 3367 1626 3371 1627
rect 3367 1621 3371 1622
rect 3391 1626 3395 1627
rect 3391 1621 3395 1622
rect 3511 1626 3515 1627
rect 3511 1621 3515 1622
rect 3591 1626 3595 1627
rect 3591 1621 3595 1622
rect 1831 1617 1835 1618
rect 112 1598 114 1617
rect 168 1601 170 1617
rect 352 1601 354 1617
rect 544 1601 546 1617
rect 728 1601 730 1617
rect 904 1601 906 1617
rect 1072 1601 1074 1617
rect 1224 1601 1226 1617
rect 1360 1601 1362 1617
rect 1496 1601 1498 1617
rect 1624 1601 1626 1617
rect 1744 1601 1746 1617
rect 166 1600 172 1601
rect 110 1597 116 1598
rect 110 1593 111 1597
rect 115 1593 116 1597
rect 166 1596 167 1600
rect 171 1596 172 1600
rect 166 1595 172 1596
rect 350 1600 356 1601
rect 350 1596 351 1600
rect 355 1596 356 1600
rect 350 1595 356 1596
rect 542 1600 548 1601
rect 542 1596 543 1600
rect 547 1596 548 1600
rect 542 1595 548 1596
rect 726 1600 732 1601
rect 726 1596 727 1600
rect 731 1596 732 1600
rect 726 1595 732 1596
rect 902 1600 908 1601
rect 902 1596 903 1600
rect 907 1596 908 1600
rect 902 1595 908 1596
rect 1070 1600 1076 1601
rect 1070 1596 1071 1600
rect 1075 1596 1076 1600
rect 1070 1595 1076 1596
rect 1222 1600 1228 1601
rect 1222 1596 1223 1600
rect 1227 1596 1228 1600
rect 1222 1595 1228 1596
rect 1358 1600 1364 1601
rect 1358 1596 1359 1600
rect 1363 1596 1364 1600
rect 1358 1595 1364 1596
rect 1494 1600 1500 1601
rect 1494 1596 1495 1600
rect 1499 1596 1500 1600
rect 1494 1595 1500 1596
rect 1622 1600 1628 1601
rect 1622 1596 1623 1600
rect 1627 1596 1628 1600
rect 1622 1595 1628 1596
rect 1742 1600 1748 1601
rect 1742 1596 1743 1600
rect 1747 1596 1748 1600
rect 1832 1598 1834 1617
rect 1742 1595 1748 1596
rect 1830 1597 1836 1598
rect 110 1592 116 1593
rect 1830 1593 1831 1597
rect 1835 1593 1836 1597
rect 1872 1593 1874 1621
rect 1976 1611 1978 1621
rect 2096 1611 2098 1621
rect 2232 1611 2234 1621
rect 2368 1611 2370 1621
rect 2504 1611 2506 1621
rect 2640 1611 2642 1621
rect 2776 1611 2778 1621
rect 2912 1611 2914 1621
rect 3056 1611 3058 1621
rect 3208 1611 3210 1621
rect 3368 1611 3370 1621
rect 3512 1611 3514 1621
rect 1974 1610 1980 1611
rect 1974 1606 1975 1610
rect 1979 1606 1980 1610
rect 1974 1605 1980 1606
rect 2094 1610 2100 1611
rect 2094 1606 2095 1610
rect 2099 1606 2100 1610
rect 2094 1605 2100 1606
rect 2230 1610 2236 1611
rect 2230 1606 2231 1610
rect 2235 1606 2236 1610
rect 2230 1605 2236 1606
rect 2366 1610 2372 1611
rect 2366 1606 2367 1610
rect 2371 1606 2372 1610
rect 2366 1605 2372 1606
rect 2502 1610 2508 1611
rect 2502 1606 2503 1610
rect 2507 1606 2508 1610
rect 2502 1605 2508 1606
rect 2638 1610 2644 1611
rect 2638 1606 2639 1610
rect 2643 1606 2644 1610
rect 2638 1605 2644 1606
rect 2774 1610 2780 1611
rect 2774 1606 2775 1610
rect 2779 1606 2780 1610
rect 2774 1605 2780 1606
rect 2910 1610 2916 1611
rect 2910 1606 2911 1610
rect 2915 1606 2916 1610
rect 2910 1605 2916 1606
rect 3054 1610 3060 1611
rect 3054 1606 3055 1610
rect 3059 1606 3060 1610
rect 3054 1605 3060 1606
rect 3206 1610 3212 1611
rect 3206 1606 3207 1610
rect 3211 1606 3212 1610
rect 3206 1605 3212 1606
rect 3366 1610 3372 1611
rect 3366 1606 3367 1610
rect 3371 1606 3372 1610
rect 3366 1605 3372 1606
rect 3510 1610 3516 1611
rect 3510 1606 3511 1610
rect 3515 1606 3516 1610
rect 3510 1605 3516 1606
rect 3592 1593 3594 1621
rect 1830 1592 1836 1593
rect 1870 1592 1876 1593
rect 1870 1588 1871 1592
rect 1875 1588 1876 1592
rect 1870 1587 1876 1588
rect 3590 1592 3596 1593
rect 3590 1588 3591 1592
rect 3595 1588 3596 1592
rect 3590 1587 3596 1588
rect 110 1580 116 1581
rect 110 1576 111 1580
rect 115 1576 116 1580
rect 110 1575 116 1576
rect 1830 1580 1836 1581
rect 1830 1576 1831 1580
rect 1835 1576 1836 1580
rect 1830 1575 1836 1576
rect 1870 1575 1876 1576
rect 112 1543 114 1575
rect 174 1562 180 1563
rect 174 1558 175 1562
rect 179 1558 180 1562
rect 174 1557 180 1558
rect 358 1562 364 1563
rect 358 1558 359 1562
rect 363 1558 364 1562
rect 358 1557 364 1558
rect 550 1562 556 1563
rect 550 1558 551 1562
rect 555 1558 556 1562
rect 550 1557 556 1558
rect 734 1562 740 1563
rect 734 1558 735 1562
rect 739 1558 740 1562
rect 734 1557 740 1558
rect 910 1562 916 1563
rect 910 1558 911 1562
rect 915 1558 916 1562
rect 910 1557 916 1558
rect 1078 1562 1084 1563
rect 1078 1558 1079 1562
rect 1083 1558 1084 1562
rect 1078 1557 1084 1558
rect 1230 1562 1236 1563
rect 1230 1558 1231 1562
rect 1235 1558 1236 1562
rect 1230 1557 1236 1558
rect 1366 1562 1372 1563
rect 1366 1558 1367 1562
rect 1371 1558 1372 1562
rect 1366 1557 1372 1558
rect 1502 1562 1508 1563
rect 1502 1558 1503 1562
rect 1507 1558 1508 1562
rect 1502 1557 1508 1558
rect 1630 1562 1636 1563
rect 1630 1558 1631 1562
rect 1635 1558 1636 1562
rect 1630 1557 1636 1558
rect 1750 1562 1756 1563
rect 1750 1558 1751 1562
rect 1755 1558 1756 1562
rect 1750 1557 1756 1558
rect 176 1543 178 1557
rect 360 1543 362 1557
rect 552 1543 554 1557
rect 736 1543 738 1557
rect 912 1543 914 1557
rect 1080 1543 1082 1557
rect 1232 1543 1234 1557
rect 1368 1543 1370 1557
rect 1504 1543 1506 1557
rect 1632 1543 1634 1557
rect 1752 1543 1754 1557
rect 1832 1543 1834 1575
rect 1870 1571 1871 1575
rect 1875 1571 1876 1575
rect 3590 1575 3596 1576
rect 1870 1570 1876 1571
rect 1966 1572 1972 1573
rect 1872 1547 1874 1570
rect 1966 1568 1967 1572
rect 1971 1568 1972 1572
rect 1966 1567 1972 1568
rect 2086 1572 2092 1573
rect 2086 1568 2087 1572
rect 2091 1568 2092 1572
rect 2086 1567 2092 1568
rect 2222 1572 2228 1573
rect 2222 1568 2223 1572
rect 2227 1568 2228 1572
rect 2222 1567 2228 1568
rect 2358 1572 2364 1573
rect 2358 1568 2359 1572
rect 2363 1568 2364 1572
rect 2358 1567 2364 1568
rect 2494 1572 2500 1573
rect 2494 1568 2495 1572
rect 2499 1568 2500 1572
rect 2494 1567 2500 1568
rect 2630 1572 2636 1573
rect 2630 1568 2631 1572
rect 2635 1568 2636 1572
rect 2630 1567 2636 1568
rect 2766 1572 2772 1573
rect 2766 1568 2767 1572
rect 2771 1568 2772 1572
rect 2766 1567 2772 1568
rect 2902 1572 2908 1573
rect 2902 1568 2903 1572
rect 2907 1568 2908 1572
rect 2902 1567 2908 1568
rect 3046 1572 3052 1573
rect 3046 1568 3047 1572
rect 3051 1568 3052 1572
rect 3046 1567 3052 1568
rect 3198 1572 3204 1573
rect 3198 1568 3199 1572
rect 3203 1568 3204 1572
rect 3198 1567 3204 1568
rect 3358 1572 3364 1573
rect 3358 1568 3359 1572
rect 3363 1568 3364 1572
rect 3358 1567 3364 1568
rect 3502 1572 3508 1573
rect 3502 1568 3503 1572
rect 3507 1568 3508 1572
rect 3590 1571 3591 1575
rect 3595 1571 3596 1575
rect 3590 1570 3596 1571
rect 3502 1567 3508 1568
rect 1968 1547 1970 1567
rect 2088 1547 2090 1567
rect 2224 1547 2226 1567
rect 2360 1547 2362 1567
rect 2496 1547 2498 1567
rect 2632 1547 2634 1567
rect 2768 1547 2770 1567
rect 2904 1547 2906 1567
rect 3048 1547 3050 1567
rect 3200 1547 3202 1567
rect 3360 1547 3362 1567
rect 3504 1547 3506 1567
rect 3592 1547 3594 1570
rect 1871 1546 1875 1547
rect 111 1542 115 1543
rect 111 1537 115 1538
rect 143 1542 147 1543
rect 143 1537 147 1538
rect 175 1542 179 1543
rect 175 1537 179 1538
rect 247 1542 251 1543
rect 247 1537 251 1538
rect 359 1542 363 1543
rect 359 1537 363 1538
rect 383 1542 387 1543
rect 383 1537 387 1538
rect 527 1542 531 1543
rect 527 1537 531 1538
rect 551 1542 555 1543
rect 551 1537 555 1538
rect 671 1542 675 1543
rect 671 1537 675 1538
rect 735 1542 739 1543
rect 735 1537 739 1538
rect 815 1542 819 1543
rect 815 1537 819 1538
rect 911 1542 915 1543
rect 911 1537 915 1538
rect 951 1542 955 1543
rect 951 1537 955 1538
rect 1079 1542 1083 1543
rect 1079 1537 1083 1538
rect 1207 1542 1211 1543
rect 1207 1537 1211 1538
rect 1231 1542 1235 1543
rect 1231 1537 1235 1538
rect 1335 1542 1339 1543
rect 1335 1537 1339 1538
rect 1367 1542 1371 1543
rect 1367 1537 1371 1538
rect 1471 1542 1475 1543
rect 1471 1537 1475 1538
rect 1503 1542 1507 1543
rect 1503 1537 1507 1538
rect 1631 1542 1635 1543
rect 1631 1537 1635 1538
rect 1751 1542 1755 1543
rect 1751 1537 1755 1538
rect 1831 1542 1835 1543
rect 1871 1541 1875 1542
rect 1967 1546 1971 1547
rect 1967 1541 1971 1542
rect 2087 1546 2091 1547
rect 2087 1541 2091 1542
rect 2167 1546 2171 1547
rect 2167 1541 2171 1542
rect 2223 1546 2227 1547
rect 2223 1541 2227 1542
rect 2255 1546 2259 1547
rect 2255 1541 2259 1542
rect 2343 1546 2347 1547
rect 2343 1541 2347 1542
rect 2359 1546 2363 1547
rect 2359 1541 2363 1542
rect 2439 1546 2443 1547
rect 2439 1541 2443 1542
rect 2495 1546 2499 1547
rect 2495 1541 2499 1542
rect 2535 1546 2539 1547
rect 2535 1541 2539 1542
rect 2631 1546 2635 1547
rect 2631 1541 2635 1542
rect 2647 1546 2651 1547
rect 2647 1541 2651 1542
rect 2767 1546 2771 1547
rect 2767 1541 2771 1542
rect 2783 1546 2787 1547
rect 2783 1541 2787 1542
rect 2903 1546 2907 1547
rect 2903 1541 2907 1542
rect 2943 1546 2947 1547
rect 2943 1541 2947 1542
rect 3047 1546 3051 1547
rect 3047 1541 3051 1542
rect 3119 1546 3123 1547
rect 3119 1541 3123 1542
rect 3199 1546 3203 1547
rect 3199 1541 3203 1542
rect 3303 1546 3307 1547
rect 3303 1541 3307 1542
rect 3359 1546 3363 1547
rect 3359 1541 3363 1542
rect 3495 1546 3499 1547
rect 3495 1541 3499 1542
rect 3503 1546 3507 1547
rect 3503 1541 3507 1542
rect 3591 1546 3595 1547
rect 3591 1541 3595 1542
rect 1831 1537 1835 1538
rect 112 1509 114 1537
rect 144 1527 146 1537
rect 248 1527 250 1537
rect 384 1527 386 1537
rect 528 1527 530 1537
rect 672 1527 674 1537
rect 816 1527 818 1537
rect 952 1527 954 1537
rect 1080 1527 1082 1537
rect 1208 1527 1210 1537
rect 1336 1527 1338 1537
rect 1472 1527 1474 1537
rect 142 1526 148 1527
rect 142 1522 143 1526
rect 147 1522 148 1526
rect 142 1521 148 1522
rect 246 1526 252 1527
rect 246 1522 247 1526
rect 251 1522 252 1526
rect 246 1521 252 1522
rect 382 1526 388 1527
rect 382 1522 383 1526
rect 387 1522 388 1526
rect 382 1521 388 1522
rect 526 1526 532 1527
rect 526 1522 527 1526
rect 531 1522 532 1526
rect 526 1521 532 1522
rect 670 1526 676 1527
rect 670 1522 671 1526
rect 675 1522 676 1526
rect 670 1521 676 1522
rect 814 1526 820 1527
rect 814 1522 815 1526
rect 819 1522 820 1526
rect 814 1521 820 1522
rect 950 1526 956 1527
rect 950 1522 951 1526
rect 955 1522 956 1526
rect 950 1521 956 1522
rect 1078 1526 1084 1527
rect 1078 1522 1079 1526
rect 1083 1522 1084 1526
rect 1078 1521 1084 1522
rect 1206 1526 1212 1527
rect 1206 1522 1207 1526
rect 1211 1522 1212 1526
rect 1206 1521 1212 1522
rect 1334 1526 1340 1527
rect 1334 1522 1335 1526
rect 1339 1522 1340 1526
rect 1334 1521 1340 1522
rect 1470 1526 1476 1527
rect 1470 1522 1471 1526
rect 1475 1522 1476 1526
rect 1470 1521 1476 1522
rect 1832 1509 1834 1537
rect 1872 1522 1874 1541
rect 2088 1525 2090 1541
rect 2168 1525 2170 1541
rect 2256 1525 2258 1541
rect 2344 1525 2346 1541
rect 2440 1525 2442 1541
rect 2536 1525 2538 1541
rect 2648 1525 2650 1541
rect 2784 1525 2786 1541
rect 2944 1525 2946 1541
rect 3120 1525 3122 1541
rect 3304 1525 3306 1541
rect 3496 1525 3498 1541
rect 2086 1524 2092 1525
rect 1870 1521 1876 1522
rect 1870 1517 1871 1521
rect 1875 1517 1876 1521
rect 2086 1520 2087 1524
rect 2091 1520 2092 1524
rect 2086 1519 2092 1520
rect 2166 1524 2172 1525
rect 2166 1520 2167 1524
rect 2171 1520 2172 1524
rect 2166 1519 2172 1520
rect 2254 1524 2260 1525
rect 2254 1520 2255 1524
rect 2259 1520 2260 1524
rect 2254 1519 2260 1520
rect 2342 1524 2348 1525
rect 2342 1520 2343 1524
rect 2347 1520 2348 1524
rect 2342 1519 2348 1520
rect 2438 1524 2444 1525
rect 2438 1520 2439 1524
rect 2443 1520 2444 1524
rect 2438 1519 2444 1520
rect 2534 1524 2540 1525
rect 2534 1520 2535 1524
rect 2539 1520 2540 1524
rect 2534 1519 2540 1520
rect 2646 1524 2652 1525
rect 2646 1520 2647 1524
rect 2651 1520 2652 1524
rect 2646 1519 2652 1520
rect 2782 1524 2788 1525
rect 2782 1520 2783 1524
rect 2787 1520 2788 1524
rect 2782 1519 2788 1520
rect 2942 1524 2948 1525
rect 2942 1520 2943 1524
rect 2947 1520 2948 1524
rect 2942 1519 2948 1520
rect 3118 1524 3124 1525
rect 3118 1520 3119 1524
rect 3123 1520 3124 1524
rect 3118 1519 3124 1520
rect 3302 1524 3308 1525
rect 3302 1520 3303 1524
rect 3307 1520 3308 1524
rect 3302 1519 3308 1520
rect 3494 1524 3500 1525
rect 3494 1520 3495 1524
rect 3499 1520 3500 1524
rect 3592 1522 3594 1541
rect 3494 1519 3500 1520
rect 3590 1521 3596 1522
rect 1870 1516 1876 1517
rect 3590 1517 3591 1521
rect 3595 1517 3596 1521
rect 3590 1516 3596 1517
rect 110 1508 116 1509
rect 110 1504 111 1508
rect 115 1504 116 1508
rect 110 1503 116 1504
rect 1830 1508 1836 1509
rect 1830 1504 1831 1508
rect 1835 1504 1836 1508
rect 1830 1503 1836 1504
rect 1870 1504 1876 1505
rect 1870 1500 1871 1504
rect 1875 1500 1876 1504
rect 1870 1499 1876 1500
rect 3590 1504 3596 1505
rect 3590 1500 3591 1504
rect 3595 1500 3596 1504
rect 3590 1499 3596 1500
rect 110 1491 116 1492
rect 110 1487 111 1491
rect 115 1487 116 1491
rect 1830 1491 1836 1492
rect 110 1486 116 1487
rect 134 1488 140 1489
rect 112 1463 114 1486
rect 134 1484 135 1488
rect 139 1484 140 1488
rect 134 1483 140 1484
rect 238 1488 244 1489
rect 238 1484 239 1488
rect 243 1484 244 1488
rect 238 1483 244 1484
rect 374 1488 380 1489
rect 374 1484 375 1488
rect 379 1484 380 1488
rect 374 1483 380 1484
rect 518 1488 524 1489
rect 518 1484 519 1488
rect 523 1484 524 1488
rect 518 1483 524 1484
rect 662 1488 668 1489
rect 662 1484 663 1488
rect 667 1484 668 1488
rect 662 1483 668 1484
rect 806 1488 812 1489
rect 806 1484 807 1488
rect 811 1484 812 1488
rect 806 1483 812 1484
rect 942 1488 948 1489
rect 942 1484 943 1488
rect 947 1484 948 1488
rect 942 1483 948 1484
rect 1070 1488 1076 1489
rect 1070 1484 1071 1488
rect 1075 1484 1076 1488
rect 1070 1483 1076 1484
rect 1198 1488 1204 1489
rect 1198 1484 1199 1488
rect 1203 1484 1204 1488
rect 1198 1483 1204 1484
rect 1326 1488 1332 1489
rect 1326 1484 1327 1488
rect 1331 1484 1332 1488
rect 1326 1483 1332 1484
rect 1462 1488 1468 1489
rect 1462 1484 1463 1488
rect 1467 1484 1468 1488
rect 1830 1487 1831 1491
rect 1835 1487 1836 1491
rect 1830 1486 1836 1487
rect 1462 1483 1468 1484
rect 136 1463 138 1483
rect 240 1463 242 1483
rect 376 1463 378 1483
rect 520 1463 522 1483
rect 664 1463 666 1483
rect 808 1463 810 1483
rect 944 1463 946 1483
rect 1072 1463 1074 1483
rect 1200 1463 1202 1483
rect 1328 1463 1330 1483
rect 1464 1463 1466 1483
rect 1832 1463 1834 1486
rect 1872 1467 1874 1499
rect 2094 1486 2100 1487
rect 2094 1482 2095 1486
rect 2099 1482 2100 1486
rect 2094 1481 2100 1482
rect 2174 1486 2180 1487
rect 2174 1482 2175 1486
rect 2179 1482 2180 1486
rect 2174 1481 2180 1482
rect 2262 1486 2268 1487
rect 2262 1482 2263 1486
rect 2267 1482 2268 1486
rect 2262 1481 2268 1482
rect 2350 1486 2356 1487
rect 2350 1482 2351 1486
rect 2355 1482 2356 1486
rect 2350 1481 2356 1482
rect 2446 1486 2452 1487
rect 2446 1482 2447 1486
rect 2451 1482 2452 1486
rect 2446 1481 2452 1482
rect 2542 1486 2548 1487
rect 2542 1482 2543 1486
rect 2547 1482 2548 1486
rect 2542 1481 2548 1482
rect 2654 1486 2660 1487
rect 2654 1482 2655 1486
rect 2659 1482 2660 1486
rect 2654 1481 2660 1482
rect 2790 1486 2796 1487
rect 2790 1482 2791 1486
rect 2795 1482 2796 1486
rect 2790 1481 2796 1482
rect 2950 1486 2956 1487
rect 2950 1482 2951 1486
rect 2955 1482 2956 1486
rect 2950 1481 2956 1482
rect 3126 1486 3132 1487
rect 3126 1482 3127 1486
rect 3131 1482 3132 1486
rect 3126 1481 3132 1482
rect 3310 1486 3316 1487
rect 3310 1482 3311 1486
rect 3315 1482 3316 1486
rect 3310 1481 3316 1482
rect 3502 1486 3508 1487
rect 3502 1482 3503 1486
rect 3507 1482 3508 1486
rect 3502 1481 3508 1482
rect 2096 1467 2098 1481
rect 2176 1467 2178 1481
rect 2264 1467 2266 1481
rect 2352 1467 2354 1481
rect 2448 1467 2450 1481
rect 2544 1467 2546 1481
rect 2656 1467 2658 1481
rect 2792 1467 2794 1481
rect 2952 1467 2954 1481
rect 3128 1467 3130 1481
rect 3312 1467 3314 1481
rect 3504 1467 3506 1481
rect 3592 1467 3594 1499
rect 1871 1466 1875 1467
rect 111 1462 115 1463
rect 111 1457 115 1458
rect 135 1462 139 1463
rect 135 1457 139 1458
rect 231 1462 235 1463
rect 231 1457 235 1458
rect 239 1462 243 1463
rect 239 1457 243 1458
rect 359 1462 363 1463
rect 359 1457 363 1458
rect 375 1462 379 1463
rect 375 1457 379 1458
rect 479 1462 483 1463
rect 479 1457 483 1458
rect 519 1462 523 1463
rect 519 1457 523 1458
rect 599 1462 603 1463
rect 599 1457 603 1458
rect 663 1462 667 1463
rect 663 1457 667 1458
rect 719 1462 723 1463
rect 719 1457 723 1458
rect 807 1462 811 1463
rect 807 1457 811 1458
rect 831 1462 835 1463
rect 831 1457 835 1458
rect 935 1462 939 1463
rect 935 1457 939 1458
rect 943 1462 947 1463
rect 943 1457 947 1458
rect 1039 1462 1043 1463
rect 1039 1457 1043 1458
rect 1071 1462 1075 1463
rect 1071 1457 1075 1458
rect 1143 1462 1147 1463
rect 1143 1457 1147 1458
rect 1199 1462 1203 1463
rect 1199 1457 1203 1458
rect 1255 1462 1259 1463
rect 1255 1457 1259 1458
rect 1327 1462 1331 1463
rect 1327 1457 1331 1458
rect 1463 1462 1467 1463
rect 1463 1457 1467 1458
rect 1831 1462 1835 1463
rect 1871 1461 1875 1462
rect 2095 1466 2099 1467
rect 2095 1461 2099 1462
rect 2175 1466 2179 1467
rect 2175 1461 2179 1462
rect 2263 1466 2267 1467
rect 2263 1461 2267 1462
rect 2343 1466 2347 1467
rect 2343 1461 2347 1462
rect 2351 1466 2355 1467
rect 2351 1461 2355 1462
rect 2423 1466 2427 1467
rect 2423 1461 2427 1462
rect 2447 1466 2451 1467
rect 2447 1461 2451 1462
rect 2503 1466 2507 1467
rect 2503 1461 2507 1462
rect 2543 1466 2547 1467
rect 2543 1461 2547 1462
rect 2607 1466 2611 1467
rect 2607 1461 2611 1462
rect 2655 1466 2659 1467
rect 2655 1461 2659 1462
rect 2735 1466 2739 1467
rect 2735 1461 2739 1462
rect 2791 1466 2795 1467
rect 2791 1461 2795 1462
rect 2895 1466 2899 1467
rect 2895 1461 2899 1462
rect 2951 1466 2955 1467
rect 2951 1461 2955 1462
rect 3079 1466 3083 1467
rect 3079 1461 3083 1462
rect 3127 1466 3131 1467
rect 3127 1461 3131 1462
rect 3279 1466 3283 1467
rect 3279 1461 3283 1462
rect 3311 1466 3315 1467
rect 3311 1461 3315 1462
rect 3479 1466 3483 1467
rect 3479 1461 3483 1462
rect 3503 1466 3507 1467
rect 3503 1461 3507 1462
rect 3591 1466 3595 1467
rect 3591 1461 3595 1462
rect 1831 1457 1835 1458
rect 112 1438 114 1457
rect 136 1441 138 1457
rect 232 1441 234 1457
rect 360 1441 362 1457
rect 480 1441 482 1457
rect 600 1441 602 1457
rect 720 1441 722 1457
rect 832 1441 834 1457
rect 936 1441 938 1457
rect 1040 1441 1042 1457
rect 1144 1441 1146 1457
rect 1256 1441 1258 1457
rect 134 1440 140 1441
rect 110 1437 116 1438
rect 110 1433 111 1437
rect 115 1433 116 1437
rect 134 1436 135 1440
rect 139 1436 140 1440
rect 134 1435 140 1436
rect 230 1440 236 1441
rect 230 1436 231 1440
rect 235 1436 236 1440
rect 230 1435 236 1436
rect 358 1440 364 1441
rect 358 1436 359 1440
rect 363 1436 364 1440
rect 358 1435 364 1436
rect 478 1440 484 1441
rect 478 1436 479 1440
rect 483 1436 484 1440
rect 478 1435 484 1436
rect 598 1440 604 1441
rect 598 1436 599 1440
rect 603 1436 604 1440
rect 598 1435 604 1436
rect 718 1440 724 1441
rect 718 1436 719 1440
rect 723 1436 724 1440
rect 718 1435 724 1436
rect 830 1440 836 1441
rect 830 1436 831 1440
rect 835 1436 836 1440
rect 830 1435 836 1436
rect 934 1440 940 1441
rect 934 1436 935 1440
rect 939 1436 940 1440
rect 934 1435 940 1436
rect 1038 1440 1044 1441
rect 1038 1436 1039 1440
rect 1043 1436 1044 1440
rect 1038 1435 1044 1436
rect 1142 1440 1148 1441
rect 1142 1436 1143 1440
rect 1147 1436 1148 1440
rect 1142 1435 1148 1436
rect 1254 1440 1260 1441
rect 1254 1436 1255 1440
rect 1259 1436 1260 1440
rect 1832 1438 1834 1457
rect 1254 1435 1260 1436
rect 1830 1437 1836 1438
rect 110 1432 116 1433
rect 1830 1433 1831 1437
rect 1835 1433 1836 1437
rect 1872 1433 1874 1461
rect 2264 1451 2266 1461
rect 2344 1451 2346 1461
rect 2424 1451 2426 1461
rect 2504 1451 2506 1461
rect 2608 1451 2610 1461
rect 2736 1451 2738 1461
rect 2896 1451 2898 1461
rect 3080 1451 3082 1461
rect 3280 1451 3282 1461
rect 3480 1451 3482 1461
rect 2262 1450 2268 1451
rect 2262 1446 2263 1450
rect 2267 1446 2268 1450
rect 2262 1445 2268 1446
rect 2342 1450 2348 1451
rect 2342 1446 2343 1450
rect 2347 1446 2348 1450
rect 2342 1445 2348 1446
rect 2422 1450 2428 1451
rect 2422 1446 2423 1450
rect 2427 1446 2428 1450
rect 2422 1445 2428 1446
rect 2502 1450 2508 1451
rect 2502 1446 2503 1450
rect 2507 1446 2508 1450
rect 2502 1445 2508 1446
rect 2606 1450 2612 1451
rect 2606 1446 2607 1450
rect 2611 1446 2612 1450
rect 2606 1445 2612 1446
rect 2734 1450 2740 1451
rect 2734 1446 2735 1450
rect 2739 1446 2740 1450
rect 2734 1445 2740 1446
rect 2894 1450 2900 1451
rect 2894 1446 2895 1450
rect 2899 1446 2900 1450
rect 2894 1445 2900 1446
rect 3078 1450 3084 1451
rect 3078 1446 3079 1450
rect 3083 1446 3084 1450
rect 3078 1445 3084 1446
rect 3278 1450 3284 1451
rect 3278 1446 3279 1450
rect 3283 1446 3284 1450
rect 3278 1445 3284 1446
rect 3478 1450 3484 1451
rect 3478 1446 3479 1450
rect 3483 1446 3484 1450
rect 3478 1445 3484 1446
rect 3592 1433 3594 1461
rect 1830 1432 1836 1433
rect 1870 1432 1876 1433
rect 1870 1428 1871 1432
rect 1875 1428 1876 1432
rect 1870 1427 1876 1428
rect 3590 1432 3596 1433
rect 3590 1428 3591 1432
rect 3595 1428 3596 1432
rect 3590 1427 3596 1428
rect 110 1420 116 1421
rect 110 1416 111 1420
rect 115 1416 116 1420
rect 110 1415 116 1416
rect 1830 1420 1836 1421
rect 1830 1416 1831 1420
rect 1835 1416 1836 1420
rect 1830 1415 1836 1416
rect 1870 1415 1876 1416
rect 112 1371 114 1415
rect 142 1402 148 1403
rect 142 1398 143 1402
rect 147 1398 148 1402
rect 142 1397 148 1398
rect 238 1402 244 1403
rect 238 1398 239 1402
rect 243 1398 244 1402
rect 238 1397 244 1398
rect 366 1402 372 1403
rect 366 1398 367 1402
rect 371 1398 372 1402
rect 366 1397 372 1398
rect 486 1402 492 1403
rect 486 1398 487 1402
rect 491 1398 492 1402
rect 486 1397 492 1398
rect 606 1402 612 1403
rect 606 1398 607 1402
rect 611 1398 612 1402
rect 606 1397 612 1398
rect 726 1402 732 1403
rect 726 1398 727 1402
rect 731 1398 732 1402
rect 726 1397 732 1398
rect 838 1402 844 1403
rect 838 1398 839 1402
rect 843 1398 844 1402
rect 838 1397 844 1398
rect 942 1402 948 1403
rect 942 1398 943 1402
rect 947 1398 948 1402
rect 942 1397 948 1398
rect 1046 1402 1052 1403
rect 1046 1398 1047 1402
rect 1051 1398 1052 1402
rect 1046 1397 1052 1398
rect 1150 1402 1156 1403
rect 1150 1398 1151 1402
rect 1155 1398 1156 1402
rect 1150 1397 1156 1398
rect 1262 1402 1268 1403
rect 1262 1398 1263 1402
rect 1267 1398 1268 1402
rect 1262 1397 1268 1398
rect 144 1371 146 1397
rect 240 1371 242 1397
rect 368 1371 370 1397
rect 488 1371 490 1397
rect 608 1371 610 1397
rect 728 1371 730 1397
rect 840 1371 842 1397
rect 944 1371 946 1397
rect 1048 1371 1050 1397
rect 1152 1371 1154 1397
rect 1264 1371 1266 1397
rect 1832 1371 1834 1415
rect 1870 1411 1871 1415
rect 1875 1411 1876 1415
rect 3590 1415 3596 1416
rect 1870 1410 1876 1411
rect 2254 1412 2260 1413
rect 1872 1391 1874 1410
rect 2254 1408 2255 1412
rect 2259 1408 2260 1412
rect 2254 1407 2260 1408
rect 2334 1412 2340 1413
rect 2334 1408 2335 1412
rect 2339 1408 2340 1412
rect 2334 1407 2340 1408
rect 2414 1412 2420 1413
rect 2414 1408 2415 1412
rect 2419 1408 2420 1412
rect 2414 1407 2420 1408
rect 2494 1412 2500 1413
rect 2494 1408 2495 1412
rect 2499 1408 2500 1412
rect 2494 1407 2500 1408
rect 2598 1412 2604 1413
rect 2598 1408 2599 1412
rect 2603 1408 2604 1412
rect 2598 1407 2604 1408
rect 2726 1412 2732 1413
rect 2726 1408 2727 1412
rect 2731 1408 2732 1412
rect 2726 1407 2732 1408
rect 2886 1412 2892 1413
rect 2886 1408 2887 1412
rect 2891 1408 2892 1412
rect 2886 1407 2892 1408
rect 3070 1412 3076 1413
rect 3070 1408 3071 1412
rect 3075 1408 3076 1412
rect 3070 1407 3076 1408
rect 3270 1412 3276 1413
rect 3270 1408 3271 1412
rect 3275 1408 3276 1412
rect 3270 1407 3276 1408
rect 3470 1412 3476 1413
rect 3470 1408 3471 1412
rect 3475 1408 3476 1412
rect 3590 1411 3591 1415
rect 3595 1411 3596 1415
rect 3590 1410 3596 1411
rect 3470 1407 3476 1408
rect 2256 1391 2258 1407
rect 2336 1391 2338 1407
rect 2416 1391 2418 1407
rect 2496 1391 2498 1407
rect 2600 1391 2602 1407
rect 2728 1391 2730 1407
rect 2888 1391 2890 1407
rect 3072 1391 3074 1407
rect 3272 1391 3274 1407
rect 3472 1391 3474 1407
rect 3592 1391 3594 1410
rect 1871 1390 1875 1391
rect 1871 1385 1875 1386
rect 2255 1390 2259 1391
rect 2255 1385 2259 1386
rect 2263 1390 2267 1391
rect 2263 1385 2267 1386
rect 2335 1390 2339 1391
rect 2335 1385 2339 1386
rect 2343 1390 2347 1391
rect 2343 1385 2347 1386
rect 2415 1390 2419 1391
rect 2415 1385 2419 1386
rect 2423 1390 2427 1391
rect 2423 1385 2427 1386
rect 2495 1390 2499 1391
rect 2495 1385 2499 1386
rect 2503 1390 2507 1391
rect 2503 1385 2507 1386
rect 2591 1390 2595 1391
rect 2591 1385 2595 1386
rect 2599 1390 2603 1391
rect 2599 1385 2603 1386
rect 2695 1390 2699 1391
rect 2695 1385 2699 1386
rect 2727 1390 2731 1391
rect 2727 1385 2731 1386
rect 2807 1390 2811 1391
rect 2807 1385 2811 1386
rect 2887 1390 2891 1391
rect 2887 1385 2891 1386
rect 2919 1390 2923 1391
rect 2919 1385 2923 1386
rect 3039 1390 3043 1391
rect 3039 1385 3043 1386
rect 3071 1390 3075 1391
rect 3071 1385 3075 1386
rect 3159 1390 3163 1391
rect 3159 1385 3163 1386
rect 3271 1390 3275 1391
rect 3271 1385 3275 1386
rect 3279 1390 3283 1391
rect 3279 1385 3283 1386
rect 3399 1390 3403 1391
rect 3399 1385 3403 1386
rect 3471 1390 3475 1391
rect 3471 1385 3475 1386
rect 3503 1390 3507 1391
rect 3503 1385 3507 1386
rect 3591 1390 3595 1391
rect 3591 1385 3595 1386
rect 111 1370 115 1371
rect 111 1365 115 1366
rect 143 1370 147 1371
rect 143 1365 147 1366
rect 239 1370 243 1371
rect 239 1365 243 1366
rect 287 1370 291 1371
rect 287 1365 291 1366
rect 367 1370 371 1371
rect 367 1365 371 1366
rect 431 1370 435 1371
rect 431 1365 435 1366
rect 487 1370 491 1371
rect 487 1365 491 1366
rect 583 1370 587 1371
rect 583 1365 587 1366
rect 607 1370 611 1371
rect 607 1365 611 1366
rect 727 1370 731 1371
rect 727 1365 731 1366
rect 735 1370 739 1371
rect 735 1365 739 1366
rect 839 1370 843 1371
rect 839 1365 843 1366
rect 879 1370 883 1371
rect 879 1365 883 1366
rect 943 1370 947 1371
rect 943 1365 947 1366
rect 1023 1370 1027 1371
rect 1023 1365 1027 1366
rect 1047 1370 1051 1371
rect 1047 1365 1051 1366
rect 1151 1370 1155 1371
rect 1151 1365 1155 1366
rect 1167 1370 1171 1371
rect 1167 1365 1171 1366
rect 1263 1370 1267 1371
rect 1263 1365 1267 1366
rect 1319 1370 1323 1371
rect 1319 1365 1323 1366
rect 1471 1370 1475 1371
rect 1471 1365 1475 1366
rect 1623 1370 1627 1371
rect 1623 1365 1627 1366
rect 1831 1370 1835 1371
rect 1872 1366 1874 1385
rect 2264 1369 2266 1385
rect 2344 1369 2346 1385
rect 2424 1369 2426 1385
rect 2504 1369 2506 1385
rect 2592 1369 2594 1385
rect 2696 1369 2698 1385
rect 2808 1369 2810 1385
rect 2920 1369 2922 1385
rect 3040 1369 3042 1385
rect 3160 1369 3162 1385
rect 3280 1369 3282 1385
rect 3400 1369 3402 1385
rect 3504 1369 3506 1385
rect 2262 1368 2268 1369
rect 1831 1365 1835 1366
rect 1870 1365 1876 1366
rect 112 1337 114 1365
rect 144 1355 146 1365
rect 288 1355 290 1365
rect 432 1355 434 1365
rect 584 1355 586 1365
rect 736 1355 738 1365
rect 880 1355 882 1365
rect 1024 1355 1026 1365
rect 1168 1355 1170 1365
rect 1320 1355 1322 1365
rect 1472 1355 1474 1365
rect 1624 1355 1626 1365
rect 142 1354 148 1355
rect 142 1350 143 1354
rect 147 1350 148 1354
rect 142 1349 148 1350
rect 286 1354 292 1355
rect 286 1350 287 1354
rect 291 1350 292 1354
rect 286 1349 292 1350
rect 430 1354 436 1355
rect 430 1350 431 1354
rect 435 1350 436 1354
rect 430 1349 436 1350
rect 582 1354 588 1355
rect 582 1350 583 1354
rect 587 1350 588 1354
rect 582 1349 588 1350
rect 734 1354 740 1355
rect 734 1350 735 1354
rect 739 1350 740 1354
rect 734 1349 740 1350
rect 878 1354 884 1355
rect 878 1350 879 1354
rect 883 1350 884 1354
rect 878 1349 884 1350
rect 1022 1354 1028 1355
rect 1022 1350 1023 1354
rect 1027 1350 1028 1354
rect 1022 1349 1028 1350
rect 1166 1354 1172 1355
rect 1166 1350 1167 1354
rect 1171 1350 1172 1354
rect 1166 1349 1172 1350
rect 1318 1354 1324 1355
rect 1318 1350 1319 1354
rect 1323 1350 1324 1354
rect 1318 1349 1324 1350
rect 1470 1354 1476 1355
rect 1470 1350 1471 1354
rect 1475 1350 1476 1354
rect 1470 1349 1476 1350
rect 1622 1354 1628 1355
rect 1622 1350 1623 1354
rect 1627 1350 1628 1354
rect 1622 1349 1628 1350
rect 1832 1337 1834 1365
rect 1870 1361 1871 1365
rect 1875 1361 1876 1365
rect 2262 1364 2263 1368
rect 2267 1364 2268 1368
rect 2262 1363 2268 1364
rect 2342 1368 2348 1369
rect 2342 1364 2343 1368
rect 2347 1364 2348 1368
rect 2342 1363 2348 1364
rect 2422 1368 2428 1369
rect 2422 1364 2423 1368
rect 2427 1364 2428 1368
rect 2422 1363 2428 1364
rect 2502 1368 2508 1369
rect 2502 1364 2503 1368
rect 2507 1364 2508 1368
rect 2502 1363 2508 1364
rect 2590 1368 2596 1369
rect 2590 1364 2591 1368
rect 2595 1364 2596 1368
rect 2590 1363 2596 1364
rect 2694 1368 2700 1369
rect 2694 1364 2695 1368
rect 2699 1364 2700 1368
rect 2694 1363 2700 1364
rect 2806 1368 2812 1369
rect 2806 1364 2807 1368
rect 2811 1364 2812 1368
rect 2806 1363 2812 1364
rect 2918 1368 2924 1369
rect 2918 1364 2919 1368
rect 2923 1364 2924 1368
rect 2918 1363 2924 1364
rect 3038 1368 3044 1369
rect 3038 1364 3039 1368
rect 3043 1364 3044 1368
rect 3038 1363 3044 1364
rect 3158 1368 3164 1369
rect 3158 1364 3159 1368
rect 3163 1364 3164 1368
rect 3158 1363 3164 1364
rect 3278 1368 3284 1369
rect 3278 1364 3279 1368
rect 3283 1364 3284 1368
rect 3278 1363 3284 1364
rect 3398 1368 3404 1369
rect 3398 1364 3399 1368
rect 3403 1364 3404 1368
rect 3398 1363 3404 1364
rect 3502 1368 3508 1369
rect 3502 1364 3503 1368
rect 3507 1364 3508 1368
rect 3592 1366 3594 1385
rect 3502 1363 3508 1364
rect 3590 1365 3596 1366
rect 1870 1360 1876 1361
rect 3590 1361 3591 1365
rect 3595 1361 3596 1365
rect 3590 1360 3596 1361
rect 1870 1348 1876 1349
rect 1870 1344 1871 1348
rect 1875 1344 1876 1348
rect 1870 1343 1876 1344
rect 3590 1348 3596 1349
rect 3590 1344 3591 1348
rect 3595 1344 3596 1348
rect 3590 1343 3596 1344
rect 110 1336 116 1337
rect 110 1332 111 1336
rect 115 1332 116 1336
rect 110 1331 116 1332
rect 1830 1336 1836 1337
rect 1830 1332 1831 1336
rect 1835 1332 1836 1336
rect 1830 1331 1836 1332
rect 110 1319 116 1320
rect 110 1315 111 1319
rect 115 1315 116 1319
rect 1830 1319 1836 1320
rect 110 1314 116 1315
rect 134 1316 140 1317
rect 112 1291 114 1314
rect 134 1312 135 1316
rect 139 1312 140 1316
rect 134 1311 140 1312
rect 278 1316 284 1317
rect 278 1312 279 1316
rect 283 1312 284 1316
rect 278 1311 284 1312
rect 422 1316 428 1317
rect 422 1312 423 1316
rect 427 1312 428 1316
rect 422 1311 428 1312
rect 574 1316 580 1317
rect 574 1312 575 1316
rect 579 1312 580 1316
rect 574 1311 580 1312
rect 726 1316 732 1317
rect 726 1312 727 1316
rect 731 1312 732 1316
rect 726 1311 732 1312
rect 870 1316 876 1317
rect 870 1312 871 1316
rect 875 1312 876 1316
rect 870 1311 876 1312
rect 1014 1316 1020 1317
rect 1014 1312 1015 1316
rect 1019 1312 1020 1316
rect 1014 1311 1020 1312
rect 1158 1316 1164 1317
rect 1158 1312 1159 1316
rect 1163 1312 1164 1316
rect 1158 1311 1164 1312
rect 1310 1316 1316 1317
rect 1310 1312 1311 1316
rect 1315 1312 1316 1316
rect 1310 1311 1316 1312
rect 1462 1316 1468 1317
rect 1462 1312 1463 1316
rect 1467 1312 1468 1316
rect 1462 1311 1468 1312
rect 1614 1316 1620 1317
rect 1614 1312 1615 1316
rect 1619 1312 1620 1316
rect 1830 1315 1831 1319
rect 1835 1315 1836 1319
rect 1830 1314 1836 1315
rect 1614 1311 1620 1312
rect 136 1291 138 1311
rect 280 1291 282 1311
rect 424 1291 426 1311
rect 576 1291 578 1311
rect 728 1291 730 1311
rect 872 1291 874 1311
rect 1016 1291 1018 1311
rect 1160 1291 1162 1311
rect 1312 1291 1314 1311
rect 1464 1291 1466 1311
rect 1616 1291 1618 1311
rect 1832 1291 1834 1314
rect 1872 1303 1874 1343
rect 2270 1330 2276 1331
rect 2270 1326 2271 1330
rect 2275 1326 2276 1330
rect 2270 1325 2276 1326
rect 2350 1330 2356 1331
rect 2350 1326 2351 1330
rect 2355 1326 2356 1330
rect 2350 1325 2356 1326
rect 2430 1330 2436 1331
rect 2430 1326 2431 1330
rect 2435 1326 2436 1330
rect 2430 1325 2436 1326
rect 2510 1330 2516 1331
rect 2510 1326 2511 1330
rect 2515 1326 2516 1330
rect 2510 1325 2516 1326
rect 2598 1330 2604 1331
rect 2598 1326 2599 1330
rect 2603 1326 2604 1330
rect 2598 1325 2604 1326
rect 2702 1330 2708 1331
rect 2702 1326 2703 1330
rect 2707 1326 2708 1330
rect 2702 1325 2708 1326
rect 2814 1330 2820 1331
rect 2814 1326 2815 1330
rect 2819 1326 2820 1330
rect 2814 1325 2820 1326
rect 2926 1330 2932 1331
rect 2926 1326 2927 1330
rect 2931 1326 2932 1330
rect 2926 1325 2932 1326
rect 3046 1330 3052 1331
rect 3046 1326 3047 1330
rect 3051 1326 3052 1330
rect 3046 1325 3052 1326
rect 3166 1330 3172 1331
rect 3166 1326 3167 1330
rect 3171 1326 3172 1330
rect 3166 1325 3172 1326
rect 3286 1330 3292 1331
rect 3286 1326 3287 1330
rect 3291 1326 3292 1330
rect 3286 1325 3292 1326
rect 3406 1330 3412 1331
rect 3406 1326 3407 1330
rect 3411 1326 3412 1330
rect 3406 1325 3412 1326
rect 3510 1330 3516 1331
rect 3510 1326 3511 1330
rect 3515 1326 3516 1330
rect 3510 1325 3516 1326
rect 2272 1303 2274 1325
rect 2352 1303 2354 1325
rect 2432 1303 2434 1325
rect 2512 1303 2514 1325
rect 2600 1303 2602 1325
rect 2704 1303 2706 1325
rect 2816 1303 2818 1325
rect 2928 1303 2930 1325
rect 3048 1303 3050 1325
rect 3168 1303 3170 1325
rect 3288 1303 3290 1325
rect 3408 1303 3410 1325
rect 3512 1303 3514 1325
rect 3592 1303 3594 1343
rect 1871 1302 1875 1303
rect 1871 1297 1875 1298
rect 2215 1302 2219 1303
rect 2215 1297 2219 1298
rect 2271 1302 2275 1303
rect 2271 1297 2275 1298
rect 2295 1302 2299 1303
rect 2295 1297 2299 1298
rect 2351 1302 2355 1303
rect 2351 1297 2355 1298
rect 2375 1302 2379 1303
rect 2375 1297 2379 1298
rect 2431 1302 2435 1303
rect 2431 1297 2435 1298
rect 2455 1302 2459 1303
rect 2455 1297 2459 1298
rect 2511 1302 2515 1303
rect 2511 1297 2515 1298
rect 2551 1302 2555 1303
rect 2551 1297 2555 1298
rect 2599 1302 2603 1303
rect 2599 1297 2603 1298
rect 2663 1302 2667 1303
rect 2663 1297 2667 1298
rect 2703 1302 2707 1303
rect 2703 1297 2707 1298
rect 2791 1302 2795 1303
rect 2791 1297 2795 1298
rect 2815 1302 2819 1303
rect 2815 1297 2819 1298
rect 2927 1302 2931 1303
rect 2927 1297 2931 1298
rect 3047 1302 3051 1303
rect 3047 1297 3051 1298
rect 3071 1302 3075 1303
rect 3071 1297 3075 1298
rect 3167 1302 3171 1303
rect 3167 1297 3171 1298
rect 3215 1302 3219 1303
rect 3215 1297 3219 1298
rect 3287 1302 3291 1303
rect 3287 1297 3291 1298
rect 3367 1302 3371 1303
rect 3367 1297 3371 1298
rect 3407 1302 3411 1303
rect 3407 1297 3411 1298
rect 3511 1302 3515 1303
rect 3511 1297 3515 1298
rect 3591 1302 3595 1303
rect 3591 1297 3595 1298
rect 111 1290 115 1291
rect 111 1285 115 1286
rect 135 1290 139 1291
rect 135 1285 139 1286
rect 263 1290 267 1291
rect 263 1285 267 1286
rect 279 1290 283 1291
rect 279 1285 283 1286
rect 423 1290 427 1291
rect 423 1285 427 1286
rect 575 1290 579 1291
rect 575 1285 579 1286
rect 591 1290 595 1291
rect 591 1285 595 1286
rect 727 1290 731 1291
rect 727 1285 731 1286
rect 759 1290 763 1291
rect 759 1285 763 1286
rect 871 1290 875 1291
rect 871 1285 875 1286
rect 927 1290 931 1291
rect 927 1285 931 1286
rect 1015 1290 1019 1291
rect 1015 1285 1019 1286
rect 1079 1290 1083 1291
rect 1079 1285 1083 1286
rect 1159 1290 1163 1291
rect 1159 1285 1163 1286
rect 1223 1290 1227 1291
rect 1223 1285 1227 1286
rect 1311 1290 1315 1291
rect 1311 1285 1315 1286
rect 1351 1290 1355 1291
rect 1351 1285 1355 1286
rect 1463 1290 1467 1291
rect 1463 1285 1467 1286
rect 1479 1290 1483 1291
rect 1479 1285 1483 1286
rect 1607 1290 1611 1291
rect 1607 1285 1611 1286
rect 1615 1290 1619 1291
rect 1615 1285 1619 1286
rect 1735 1290 1739 1291
rect 1735 1285 1739 1286
rect 1831 1290 1835 1291
rect 1831 1285 1835 1286
rect 112 1266 114 1285
rect 136 1269 138 1285
rect 264 1269 266 1285
rect 424 1269 426 1285
rect 592 1269 594 1285
rect 760 1269 762 1285
rect 928 1269 930 1285
rect 1080 1269 1082 1285
rect 1224 1269 1226 1285
rect 1352 1269 1354 1285
rect 1480 1269 1482 1285
rect 1608 1269 1610 1285
rect 1736 1269 1738 1285
rect 134 1268 140 1269
rect 110 1265 116 1266
rect 110 1261 111 1265
rect 115 1261 116 1265
rect 134 1264 135 1268
rect 139 1264 140 1268
rect 134 1263 140 1264
rect 262 1268 268 1269
rect 262 1264 263 1268
rect 267 1264 268 1268
rect 262 1263 268 1264
rect 422 1268 428 1269
rect 422 1264 423 1268
rect 427 1264 428 1268
rect 422 1263 428 1264
rect 590 1268 596 1269
rect 590 1264 591 1268
rect 595 1264 596 1268
rect 590 1263 596 1264
rect 758 1268 764 1269
rect 758 1264 759 1268
rect 763 1264 764 1268
rect 758 1263 764 1264
rect 926 1268 932 1269
rect 926 1264 927 1268
rect 931 1264 932 1268
rect 926 1263 932 1264
rect 1078 1268 1084 1269
rect 1078 1264 1079 1268
rect 1083 1264 1084 1268
rect 1078 1263 1084 1264
rect 1222 1268 1228 1269
rect 1222 1264 1223 1268
rect 1227 1264 1228 1268
rect 1222 1263 1228 1264
rect 1350 1268 1356 1269
rect 1350 1264 1351 1268
rect 1355 1264 1356 1268
rect 1350 1263 1356 1264
rect 1478 1268 1484 1269
rect 1478 1264 1479 1268
rect 1483 1264 1484 1268
rect 1478 1263 1484 1264
rect 1606 1268 1612 1269
rect 1606 1264 1607 1268
rect 1611 1264 1612 1268
rect 1606 1263 1612 1264
rect 1734 1268 1740 1269
rect 1734 1264 1735 1268
rect 1739 1264 1740 1268
rect 1832 1266 1834 1285
rect 1872 1269 1874 1297
rect 2216 1287 2218 1297
rect 2296 1287 2298 1297
rect 2376 1287 2378 1297
rect 2456 1287 2458 1297
rect 2552 1287 2554 1297
rect 2664 1287 2666 1297
rect 2792 1287 2794 1297
rect 2928 1287 2930 1297
rect 3072 1287 3074 1297
rect 3216 1287 3218 1297
rect 3368 1287 3370 1297
rect 3512 1287 3514 1297
rect 2214 1286 2220 1287
rect 2214 1282 2215 1286
rect 2219 1282 2220 1286
rect 2214 1281 2220 1282
rect 2294 1286 2300 1287
rect 2294 1282 2295 1286
rect 2299 1282 2300 1286
rect 2294 1281 2300 1282
rect 2374 1286 2380 1287
rect 2374 1282 2375 1286
rect 2379 1282 2380 1286
rect 2374 1281 2380 1282
rect 2454 1286 2460 1287
rect 2454 1282 2455 1286
rect 2459 1282 2460 1286
rect 2454 1281 2460 1282
rect 2550 1286 2556 1287
rect 2550 1282 2551 1286
rect 2555 1282 2556 1286
rect 2550 1281 2556 1282
rect 2662 1286 2668 1287
rect 2662 1282 2663 1286
rect 2667 1282 2668 1286
rect 2662 1281 2668 1282
rect 2790 1286 2796 1287
rect 2790 1282 2791 1286
rect 2795 1282 2796 1286
rect 2790 1281 2796 1282
rect 2926 1286 2932 1287
rect 2926 1282 2927 1286
rect 2931 1282 2932 1286
rect 2926 1281 2932 1282
rect 3070 1286 3076 1287
rect 3070 1282 3071 1286
rect 3075 1282 3076 1286
rect 3070 1281 3076 1282
rect 3214 1286 3220 1287
rect 3214 1282 3215 1286
rect 3219 1282 3220 1286
rect 3214 1281 3220 1282
rect 3366 1286 3372 1287
rect 3366 1282 3367 1286
rect 3371 1282 3372 1286
rect 3366 1281 3372 1282
rect 3510 1286 3516 1287
rect 3510 1282 3511 1286
rect 3515 1282 3516 1286
rect 3510 1281 3516 1282
rect 3592 1269 3594 1297
rect 1870 1268 1876 1269
rect 1734 1263 1740 1264
rect 1830 1265 1836 1266
rect 110 1260 116 1261
rect 1830 1261 1831 1265
rect 1835 1261 1836 1265
rect 1870 1264 1871 1268
rect 1875 1264 1876 1268
rect 1870 1263 1876 1264
rect 3590 1268 3596 1269
rect 3590 1264 3591 1268
rect 3595 1264 3596 1268
rect 3590 1263 3596 1264
rect 1830 1260 1836 1261
rect 1870 1251 1876 1252
rect 110 1248 116 1249
rect 110 1244 111 1248
rect 115 1244 116 1248
rect 110 1243 116 1244
rect 1830 1248 1836 1249
rect 1830 1244 1831 1248
rect 1835 1244 1836 1248
rect 1870 1247 1871 1251
rect 1875 1247 1876 1251
rect 3590 1251 3596 1252
rect 1870 1246 1876 1247
rect 2206 1248 2212 1249
rect 1830 1243 1836 1244
rect 112 1207 114 1243
rect 142 1230 148 1231
rect 142 1226 143 1230
rect 147 1226 148 1230
rect 142 1225 148 1226
rect 270 1230 276 1231
rect 270 1226 271 1230
rect 275 1226 276 1230
rect 270 1225 276 1226
rect 430 1230 436 1231
rect 430 1226 431 1230
rect 435 1226 436 1230
rect 430 1225 436 1226
rect 598 1230 604 1231
rect 598 1226 599 1230
rect 603 1226 604 1230
rect 598 1225 604 1226
rect 766 1230 772 1231
rect 766 1226 767 1230
rect 771 1226 772 1230
rect 766 1225 772 1226
rect 934 1230 940 1231
rect 934 1226 935 1230
rect 939 1226 940 1230
rect 934 1225 940 1226
rect 1086 1230 1092 1231
rect 1086 1226 1087 1230
rect 1091 1226 1092 1230
rect 1086 1225 1092 1226
rect 1230 1230 1236 1231
rect 1230 1226 1231 1230
rect 1235 1226 1236 1230
rect 1230 1225 1236 1226
rect 1358 1230 1364 1231
rect 1358 1226 1359 1230
rect 1363 1226 1364 1230
rect 1358 1225 1364 1226
rect 1486 1230 1492 1231
rect 1486 1226 1487 1230
rect 1491 1226 1492 1230
rect 1486 1225 1492 1226
rect 1614 1230 1620 1231
rect 1614 1226 1615 1230
rect 1619 1226 1620 1230
rect 1614 1225 1620 1226
rect 1742 1230 1748 1231
rect 1742 1226 1743 1230
rect 1747 1226 1748 1230
rect 1742 1225 1748 1226
rect 144 1207 146 1225
rect 272 1207 274 1225
rect 432 1207 434 1225
rect 600 1207 602 1225
rect 768 1207 770 1225
rect 936 1207 938 1225
rect 1088 1207 1090 1225
rect 1232 1207 1234 1225
rect 1360 1207 1362 1225
rect 1488 1207 1490 1225
rect 1616 1207 1618 1225
rect 1744 1207 1746 1225
rect 1832 1207 1834 1243
rect 1872 1223 1874 1246
rect 2206 1244 2207 1248
rect 2211 1244 2212 1248
rect 2206 1243 2212 1244
rect 2286 1248 2292 1249
rect 2286 1244 2287 1248
rect 2291 1244 2292 1248
rect 2286 1243 2292 1244
rect 2366 1248 2372 1249
rect 2366 1244 2367 1248
rect 2371 1244 2372 1248
rect 2366 1243 2372 1244
rect 2446 1248 2452 1249
rect 2446 1244 2447 1248
rect 2451 1244 2452 1248
rect 2446 1243 2452 1244
rect 2542 1248 2548 1249
rect 2542 1244 2543 1248
rect 2547 1244 2548 1248
rect 2542 1243 2548 1244
rect 2654 1248 2660 1249
rect 2654 1244 2655 1248
rect 2659 1244 2660 1248
rect 2654 1243 2660 1244
rect 2782 1248 2788 1249
rect 2782 1244 2783 1248
rect 2787 1244 2788 1248
rect 2782 1243 2788 1244
rect 2918 1248 2924 1249
rect 2918 1244 2919 1248
rect 2923 1244 2924 1248
rect 2918 1243 2924 1244
rect 3062 1248 3068 1249
rect 3062 1244 3063 1248
rect 3067 1244 3068 1248
rect 3062 1243 3068 1244
rect 3206 1248 3212 1249
rect 3206 1244 3207 1248
rect 3211 1244 3212 1248
rect 3206 1243 3212 1244
rect 3358 1248 3364 1249
rect 3358 1244 3359 1248
rect 3363 1244 3364 1248
rect 3358 1243 3364 1244
rect 3502 1248 3508 1249
rect 3502 1244 3503 1248
rect 3507 1244 3508 1248
rect 3590 1247 3591 1251
rect 3595 1247 3596 1251
rect 3590 1246 3596 1247
rect 3502 1243 3508 1244
rect 2208 1223 2210 1243
rect 2288 1223 2290 1243
rect 2368 1223 2370 1243
rect 2448 1223 2450 1243
rect 2544 1223 2546 1243
rect 2656 1223 2658 1243
rect 2784 1223 2786 1243
rect 2920 1223 2922 1243
rect 3064 1223 3066 1243
rect 3208 1223 3210 1243
rect 3360 1223 3362 1243
rect 3504 1223 3506 1243
rect 3592 1223 3594 1246
rect 1871 1222 1875 1223
rect 1871 1217 1875 1218
rect 2111 1222 2115 1223
rect 2111 1217 2115 1218
rect 2207 1222 2211 1223
rect 2207 1217 2211 1218
rect 2287 1222 2291 1223
rect 2287 1217 2291 1218
rect 2303 1222 2307 1223
rect 2303 1217 2307 1218
rect 2367 1222 2371 1223
rect 2367 1217 2371 1218
rect 2407 1222 2411 1223
rect 2407 1217 2411 1218
rect 2447 1222 2451 1223
rect 2447 1217 2451 1218
rect 2527 1222 2531 1223
rect 2527 1217 2531 1218
rect 2543 1222 2547 1223
rect 2543 1217 2547 1218
rect 2647 1222 2651 1223
rect 2647 1217 2651 1218
rect 2655 1222 2659 1223
rect 2655 1217 2659 1218
rect 2775 1222 2779 1223
rect 2775 1217 2779 1218
rect 2783 1222 2787 1223
rect 2783 1217 2787 1218
rect 2911 1222 2915 1223
rect 2911 1217 2915 1218
rect 2919 1222 2923 1223
rect 2919 1217 2923 1218
rect 3055 1222 3059 1223
rect 3055 1217 3059 1218
rect 3063 1222 3067 1223
rect 3063 1217 3067 1218
rect 3199 1222 3203 1223
rect 3199 1217 3203 1218
rect 3207 1222 3211 1223
rect 3207 1217 3211 1218
rect 3343 1222 3347 1223
rect 3343 1217 3347 1218
rect 3359 1222 3363 1223
rect 3359 1217 3363 1218
rect 3495 1222 3499 1223
rect 3495 1217 3499 1218
rect 3503 1222 3507 1223
rect 3503 1217 3507 1218
rect 3591 1222 3595 1223
rect 3591 1217 3595 1218
rect 111 1206 115 1207
rect 111 1201 115 1202
rect 143 1206 147 1207
rect 143 1201 147 1202
rect 271 1206 275 1207
rect 271 1201 275 1202
rect 311 1206 315 1207
rect 311 1201 315 1202
rect 431 1206 435 1207
rect 431 1201 435 1202
rect 487 1206 491 1207
rect 487 1201 491 1202
rect 599 1206 603 1207
rect 599 1201 603 1202
rect 671 1206 675 1207
rect 671 1201 675 1202
rect 767 1206 771 1207
rect 767 1201 771 1202
rect 847 1206 851 1207
rect 847 1201 851 1202
rect 935 1206 939 1207
rect 935 1201 939 1202
rect 1007 1206 1011 1207
rect 1007 1201 1011 1202
rect 1087 1206 1091 1207
rect 1087 1201 1091 1202
rect 1159 1206 1163 1207
rect 1159 1201 1163 1202
rect 1231 1206 1235 1207
rect 1231 1201 1235 1202
rect 1295 1206 1299 1207
rect 1295 1201 1299 1202
rect 1359 1206 1363 1207
rect 1359 1201 1363 1202
rect 1415 1206 1419 1207
rect 1415 1201 1419 1202
rect 1487 1206 1491 1207
rect 1487 1201 1491 1202
rect 1535 1206 1539 1207
rect 1535 1201 1539 1202
rect 1615 1206 1619 1207
rect 1615 1201 1619 1202
rect 1655 1206 1659 1207
rect 1655 1201 1659 1202
rect 1743 1206 1747 1207
rect 1743 1201 1747 1202
rect 1751 1206 1755 1207
rect 1751 1201 1755 1202
rect 1831 1206 1835 1207
rect 1831 1201 1835 1202
rect 112 1173 114 1201
rect 144 1191 146 1201
rect 312 1191 314 1201
rect 488 1191 490 1201
rect 672 1191 674 1201
rect 848 1191 850 1201
rect 1008 1191 1010 1201
rect 1160 1191 1162 1201
rect 1296 1191 1298 1201
rect 1416 1191 1418 1201
rect 1536 1191 1538 1201
rect 1656 1191 1658 1201
rect 1752 1191 1754 1201
rect 142 1190 148 1191
rect 142 1186 143 1190
rect 147 1186 148 1190
rect 142 1185 148 1186
rect 310 1190 316 1191
rect 310 1186 311 1190
rect 315 1186 316 1190
rect 310 1185 316 1186
rect 486 1190 492 1191
rect 486 1186 487 1190
rect 491 1186 492 1190
rect 486 1185 492 1186
rect 670 1190 676 1191
rect 670 1186 671 1190
rect 675 1186 676 1190
rect 670 1185 676 1186
rect 846 1190 852 1191
rect 846 1186 847 1190
rect 851 1186 852 1190
rect 846 1185 852 1186
rect 1006 1190 1012 1191
rect 1006 1186 1007 1190
rect 1011 1186 1012 1190
rect 1006 1185 1012 1186
rect 1158 1190 1164 1191
rect 1158 1186 1159 1190
rect 1163 1186 1164 1190
rect 1158 1185 1164 1186
rect 1294 1190 1300 1191
rect 1294 1186 1295 1190
rect 1299 1186 1300 1190
rect 1294 1185 1300 1186
rect 1414 1190 1420 1191
rect 1414 1186 1415 1190
rect 1419 1186 1420 1190
rect 1414 1185 1420 1186
rect 1534 1190 1540 1191
rect 1534 1186 1535 1190
rect 1539 1186 1540 1190
rect 1534 1185 1540 1186
rect 1654 1190 1660 1191
rect 1654 1186 1655 1190
rect 1659 1186 1660 1190
rect 1654 1185 1660 1186
rect 1750 1190 1756 1191
rect 1750 1186 1751 1190
rect 1755 1186 1756 1190
rect 1750 1185 1756 1186
rect 1832 1173 1834 1201
rect 1872 1198 1874 1217
rect 2112 1201 2114 1217
rect 2208 1201 2210 1217
rect 2304 1201 2306 1217
rect 2408 1201 2410 1217
rect 2528 1201 2530 1217
rect 2648 1201 2650 1217
rect 2776 1201 2778 1217
rect 2912 1201 2914 1217
rect 3056 1201 3058 1217
rect 3200 1201 3202 1217
rect 3344 1201 3346 1217
rect 3496 1201 3498 1217
rect 2110 1200 2116 1201
rect 1870 1197 1876 1198
rect 1870 1193 1871 1197
rect 1875 1193 1876 1197
rect 2110 1196 2111 1200
rect 2115 1196 2116 1200
rect 2110 1195 2116 1196
rect 2206 1200 2212 1201
rect 2206 1196 2207 1200
rect 2211 1196 2212 1200
rect 2206 1195 2212 1196
rect 2302 1200 2308 1201
rect 2302 1196 2303 1200
rect 2307 1196 2308 1200
rect 2302 1195 2308 1196
rect 2406 1200 2412 1201
rect 2406 1196 2407 1200
rect 2411 1196 2412 1200
rect 2406 1195 2412 1196
rect 2526 1200 2532 1201
rect 2526 1196 2527 1200
rect 2531 1196 2532 1200
rect 2526 1195 2532 1196
rect 2646 1200 2652 1201
rect 2646 1196 2647 1200
rect 2651 1196 2652 1200
rect 2646 1195 2652 1196
rect 2774 1200 2780 1201
rect 2774 1196 2775 1200
rect 2779 1196 2780 1200
rect 2774 1195 2780 1196
rect 2910 1200 2916 1201
rect 2910 1196 2911 1200
rect 2915 1196 2916 1200
rect 2910 1195 2916 1196
rect 3054 1200 3060 1201
rect 3054 1196 3055 1200
rect 3059 1196 3060 1200
rect 3054 1195 3060 1196
rect 3198 1200 3204 1201
rect 3198 1196 3199 1200
rect 3203 1196 3204 1200
rect 3198 1195 3204 1196
rect 3342 1200 3348 1201
rect 3342 1196 3343 1200
rect 3347 1196 3348 1200
rect 3342 1195 3348 1196
rect 3494 1200 3500 1201
rect 3494 1196 3495 1200
rect 3499 1196 3500 1200
rect 3592 1198 3594 1217
rect 3494 1195 3500 1196
rect 3590 1197 3596 1198
rect 1870 1192 1876 1193
rect 3590 1193 3591 1197
rect 3595 1193 3596 1197
rect 3590 1192 3596 1193
rect 1870 1180 1876 1181
rect 1870 1176 1871 1180
rect 1875 1176 1876 1180
rect 1870 1175 1876 1176
rect 3590 1180 3596 1181
rect 3590 1176 3591 1180
rect 3595 1176 3596 1180
rect 3590 1175 3596 1176
rect 110 1172 116 1173
rect 110 1168 111 1172
rect 115 1168 116 1172
rect 110 1167 116 1168
rect 1830 1172 1836 1173
rect 1830 1168 1831 1172
rect 1835 1168 1836 1172
rect 1830 1167 1836 1168
rect 110 1155 116 1156
rect 110 1151 111 1155
rect 115 1151 116 1155
rect 1830 1155 1836 1156
rect 110 1150 116 1151
rect 134 1152 140 1153
rect 112 1131 114 1150
rect 134 1148 135 1152
rect 139 1148 140 1152
rect 134 1147 140 1148
rect 302 1152 308 1153
rect 302 1148 303 1152
rect 307 1148 308 1152
rect 302 1147 308 1148
rect 478 1152 484 1153
rect 478 1148 479 1152
rect 483 1148 484 1152
rect 478 1147 484 1148
rect 662 1152 668 1153
rect 662 1148 663 1152
rect 667 1148 668 1152
rect 662 1147 668 1148
rect 838 1152 844 1153
rect 838 1148 839 1152
rect 843 1148 844 1152
rect 838 1147 844 1148
rect 998 1152 1004 1153
rect 998 1148 999 1152
rect 1003 1148 1004 1152
rect 998 1147 1004 1148
rect 1150 1152 1156 1153
rect 1150 1148 1151 1152
rect 1155 1148 1156 1152
rect 1150 1147 1156 1148
rect 1286 1152 1292 1153
rect 1286 1148 1287 1152
rect 1291 1148 1292 1152
rect 1286 1147 1292 1148
rect 1406 1152 1412 1153
rect 1406 1148 1407 1152
rect 1411 1148 1412 1152
rect 1406 1147 1412 1148
rect 1526 1152 1532 1153
rect 1526 1148 1527 1152
rect 1531 1148 1532 1152
rect 1526 1147 1532 1148
rect 1646 1152 1652 1153
rect 1646 1148 1647 1152
rect 1651 1148 1652 1152
rect 1646 1147 1652 1148
rect 1742 1152 1748 1153
rect 1742 1148 1743 1152
rect 1747 1148 1748 1152
rect 1830 1151 1831 1155
rect 1835 1151 1836 1155
rect 1830 1150 1836 1151
rect 1742 1147 1748 1148
rect 136 1131 138 1147
rect 304 1131 306 1147
rect 480 1131 482 1147
rect 664 1131 666 1147
rect 840 1131 842 1147
rect 1000 1131 1002 1147
rect 1152 1131 1154 1147
rect 1288 1131 1290 1147
rect 1408 1131 1410 1147
rect 1528 1131 1530 1147
rect 1648 1131 1650 1147
rect 1744 1131 1746 1147
rect 1832 1131 1834 1150
rect 1872 1139 1874 1175
rect 2118 1162 2124 1163
rect 2118 1158 2119 1162
rect 2123 1158 2124 1162
rect 2118 1157 2124 1158
rect 2214 1162 2220 1163
rect 2214 1158 2215 1162
rect 2219 1158 2220 1162
rect 2214 1157 2220 1158
rect 2310 1162 2316 1163
rect 2310 1158 2311 1162
rect 2315 1158 2316 1162
rect 2310 1157 2316 1158
rect 2414 1162 2420 1163
rect 2414 1158 2415 1162
rect 2419 1158 2420 1162
rect 2414 1157 2420 1158
rect 2534 1162 2540 1163
rect 2534 1158 2535 1162
rect 2539 1158 2540 1162
rect 2534 1157 2540 1158
rect 2654 1162 2660 1163
rect 2654 1158 2655 1162
rect 2659 1158 2660 1162
rect 2654 1157 2660 1158
rect 2782 1162 2788 1163
rect 2782 1158 2783 1162
rect 2787 1158 2788 1162
rect 2782 1157 2788 1158
rect 2918 1162 2924 1163
rect 2918 1158 2919 1162
rect 2923 1158 2924 1162
rect 2918 1157 2924 1158
rect 3062 1162 3068 1163
rect 3062 1158 3063 1162
rect 3067 1158 3068 1162
rect 3062 1157 3068 1158
rect 3206 1162 3212 1163
rect 3206 1158 3207 1162
rect 3211 1158 3212 1162
rect 3206 1157 3212 1158
rect 3350 1162 3356 1163
rect 3350 1158 3351 1162
rect 3355 1158 3356 1162
rect 3350 1157 3356 1158
rect 3502 1162 3508 1163
rect 3502 1158 3503 1162
rect 3507 1158 3508 1162
rect 3502 1157 3508 1158
rect 2120 1139 2122 1157
rect 2216 1139 2218 1157
rect 2312 1139 2314 1157
rect 2416 1139 2418 1157
rect 2536 1139 2538 1157
rect 2656 1139 2658 1157
rect 2784 1139 2786 1157
rect 2920 1139 2922 1157
rect 3064 1139 3066 1157
rect 3208 1139 3210 1157
rect 3352 1139 3354 1157
rect 3504 1139 3506 1157
rect 3592 1139 3594 1175
rect 1871 1138 1875 1139
rect 1871 1133 1875 1134
rect 1903 1138 1907 1139
rect 1903 1133 1907 1134
rect 2119 1138 2123 1139
rect 2119 1133 2123 1134
rect 2127 1138 2131 1139
rect 2127 1133 2131 1134
rect 2215 1138 2219 1139
rect 2215 1133 2219 1134
rect 2311 1138 2315 1139
rect 2311 1133 2315 1134
rect 2359 1138 2363 1139
rect 2359 1133 2363 1134
rect 2415 1138 2419 1139
rect 2415 1133 2419 1134
rect 2535 1138 2539 1139
rect 2535 1133 2539 1134
rect 2575 1138 2579 1139
rect 2575 1133 2579 1134
rect 2655 1138 2659 1139
rect 2655 1133 2659 1134
rect 2775 1138 2779 1139
rect 2775 1133 2779 1134
rect 2783 1138 2787 1139
rect 2783 1133 2787 1134
rect 2919 1138 2923 1139
rect 2919 1133 2923 1134
rect 2967 1138 2971 1139
rect 2967 1133 2971 1134
rect 3063 1138 3067 1139
rect 3063 1133 3067 1134
rect 3159 1138 3163 1139
rect 3159 1133 3163 1134
rect 3207 1138 3211 1139
rect 3207 1133 3211 1134
rect 3343 1138 3347 1139
rect 3343 1133 3347 1134
rect 3351 1138 3355 1139
rect 3351 1133 3355 1134
rect 3503 1138 3507 1139
rect 3503 1133 3507 1134
rect 3511 1138 3515 1139
rect 3511 1133 3515 1134
rect 3591 1138 3595 1139
rect 3591 1133 3595 1134
rect 111 1130 115 1131
rect 111 1125 115 1126
rect 135 1130 139 1131
rect 135 1125 139 1126
rect 247 1130 251 1131
rect 247 1125 251 1126
rect 303 1130 307 1131
rect 303 1125 307 1126
rect 383 1130 387 1131
rect 383 1125 387 1126
rect 479 1130 483 1131
rect 479 1125 483 1126
rect 519 1130 523 1131
rect 519 1125 523 1126
rect 647 1130 651 1131
rect 647 1125 651 1126
rect 663 1130 667 1131
rect 663 1125 667 1126
rect 775 1130 779 1131
rect 775 1125 779 1126
rect 839 1130 843 1131
rect 839 1125 843 1126
rect 895 1130 899 1131
rect 895 1125 899 1126
rect 999 1130 1003 1131
rect 999 1125 1003 1126
rect 1015 1130 1019 1131
rect 1015 1125 1019 1126
rect 1135 1130 1139 1131
rect 1135 1125 1139 1126
rect 1151 1130 1155 1131
rect 1151 1125 1155 1126
rect 1255 1130 1259 1131
rect 1255 1125 1259 1126
rect 1287 1130 1291 1131
rect 1287 1125 1291 1126
rect 1375 1130 1379 1131
rect 1375 1125 1379 1126
rect 1407 1130 1411 1131
rect 1407 1125 1411 1126
rect 1503 1130 1507 1131
rect 1503 1125 1507 1126
rect 1527 1130 1531 1131
rect 1527 1125 1531 1126
rect 1631 1130 1635 1131
rect 1631 1125 1635 1126
rect 1647 1130 1651 1131
rect 1647 1125 1651 1126
rect 1743 1130 1747 1131
rect 1743 1125 1747 1126
rect 1831 1130 1835 1131
rect 1831 1125 1835 1126
rect 112 1106 114 1125
rect 136 1109 138 1125
rect 248 1109 250 1125
rect 384 1109 386 1125
rect 520 1109 522 1125
rect 648 1109 650 1125
rect 776 1109 778 1125
rect 896 1109 898 1125
rect 1016 1109 1018 1125
rect 1136 1109 1138 1125
rect 1256 1109 1258 1125
rect 1376 1109 1378 1125
rect 1504 1109 1506 1125
rect 1632 1109 1634 1125
rect 1744 1109 1746 1125
rect 134 1108 140 1109
rect 110 1105 116 1106
rect 110 1101 111 1105
rect 115 1101 116 1105
rect 134 1104 135 1108
rect 139 1104 140 1108
rect 134 1103 140 1104
rect 246 1108 252 1109
rect 246 1104 247 1108
rect 251 1104 252 1108
rect 246 1103 252 1104
rect 382 1108 388 1109
rect 382 1104 383 1108
rect 387 1104 388 1108
rect 382 1103 388 1104
rect 518 1108 524 1109
rect 518 1104 519 1108
rect 523 1104 524 1108
rect 518 1103 524 1104
rect 646 1108 652 1109
rect 646 1104 647 1108
rect 651 1104 652 1108
rect 646 1103 652 1104
rect 774 1108 780 1109
rect 774 1104 775 1108
rect 779 1104 780 1108
rect 774 1103 780 1104
rect 894 1108 900 1109
rect 894 1104 895 1108
rect 899 1104 900 1108
rect 894 1103 900 1104
rect 1014 1108 1020 1109
rect 1014 1104 1015 1108
rect 1019 1104 1020 1108
rect 1014 1103 1020 1104
rect 1134 1108 1140 1109
rect 1134 1104 1135 1108
rect 1139 1104 1140 1108
rect 1134 1103 1140 1104
rect 1254 1108 1260 1109
rect 1254 1104 1255 1108
rect 1259 1104 1260 1108
rect 1254 1103 1260 1104
rect 1374 1108 1380 1109
rect 1374 1104 1375 1108
rect 1379 1104 1380 1108
rect 1374 1103 1380 1104
rect 1502 1108 1508 1109
rect 1502 1104 1503 1108
rect 1507 1104 1508 1108
rect 1502 1103 1508 1104
rect 1630 1108 1636 1109
rect 1630 1104 1631 1108
rect 1635 1104 1636 1108
rect 1630 1103 1636 1104
rect 1742 1108 1748 1109
rect 1742 1104 1743 1108
rect 1747 1104 1748 1108
rect 1832 1106 1834 1125
rect 1742 1103 1748 1104
rect 1830 1105 1836 1106
rect 1872 1105 1874 1133
rect 1904 1123 1906 1133
rect 2128 1123 2130 1133
rect 2360 1123 2362 1133
rect 2576 1123 2578 1133
rect 2776 1123 2778 1133
rect 2968 1123 2970 1133
rect 3160 1123 3162 1133
rect 3344 1123 3346 1133
rect 3512 1123 3514 1133
rect 1902 1122 1908 1123
rect 1902 1118 1903 1122
rect 1907 1118 1908 1122
rect 1902 1117 1908 1118
rect 2126 1122 2132 1123
rect 2126 1118 2127 1122
rect 2131 1118 2132 1122
rect 2126 1117 2132 1118
rect 2358 1122 2364 1123
rect 2358 1118 2359 1122
rect 2363 1118 2364 1122
rect 2358 1117 2364 1118
rect 2574 1122 2580 1123
rect 2574 1118 2575 1122
rect 2579 1118 2580 1122
rect 2574 1117 2580 1118
rect 2774 1122 2780 1123
rect 2774 1118 2775 1122
rect 2779 1118 2780 1122
rect 2774 1117 2780 1118
rect 2966 1122 2972 1123
rect 2966 1118 2967 1122
rect 2971 1118 2972 1122
rect 2966 1117 2972 1118
rect 3158 1122 3164 1123
rect 3158 1118 3159 1122
rect 3163 1118 3164 1122
rect 3158 1117 3164 1118
rect 3342 1122 3348 1123
rect 3342 1118 3343 1122
rect 3347 1118 3348 1122
rect 3342 1117 3348 1118
rect 3510 1122 3516 1123
rect 3510 1118 3511 1122
rect 3515 1118 3516 1122
rect 3510 1117 3516 1118
rect 3592 1105 3594 1133
rect 110 1100 116 1101
rect 1830 1101 1831 1105
rect 1835 1101 1836 1105
rect 1830 1100 1836 1101
rect 1870 1104 1876 1105
rect 1870 1100 1871 1104
rect 1875 1100 1876 1104
rect 1870 1099 1876 1100
rect 3590 1104 3596 1105
rect 3590 1100 3591 1104
rect 3595 1100 3596 1104
rect 3590 1099 3596 1100
rect 110 1088 116 1089
rect 110 1084 111 1088
rect 115 1084 116 1088
rect 110 1083 116 1084
rect 1830 1088 1836 1089
rect 1830 1084 1831 1088
rect 1835 1084 1836 1088
rect 1830 1083 1836 1084
rect 1870 1087 1876 1088
rect 1870 1083 1871 1087
rect 1875 1083 1876 1087
rect 3590 1087 3596 1088
rect 112 1043 114 1083
rect 142 1070 148 1071
rect 142 1066 143 1070
rect 147 1066 148 1070
rect 142 1065 148 1066
rect 254 1070 260 1071
rect 254 1066 255 1070
rect 259 1066 260 1070
rect 254 1065 260 1066
rect 390 1070 396 1071
rect 390 1066 391 1070
rect 395 1066 396 1070
rect 390 1065 396 1066
rect 526 1070 532 1071
rect 526 1066 527 1070
rect 531 1066 532 1070
rect 526 1065 532 1066
rect 654 1070 660 1071
rect 654 1066 655 1070
rect 659 1066 660 1070
rect 654 1065 660 1066
rect 782 1070 788 1071
rect 782 1066 783 1070
rect 787 1066 788 1070
rect 782 1065 788 1066
rect 902 1070 908 1071
rect 902 1066 903 1070
rect 907 1066 908 1070
rect 902 1065 908 1066
rect 1022 1070 1028 1071
rect 1022 1066 1023 1070
rect 1027 1066 1028 1070
rect 1022 1065 1028 1066
rect 1142 1070 1148 1071
rect 1142 1066 1143 1070
rect 1147 1066 1148 1070
rect 1142 1065 1148 1066
rect 1262 1070 1268 1071
rect 1262 1066 1263 1070
rect 1267 1066 1268 1070
rect 1262 1065 1268 1066
rect 1382 1070 1388 1071
rect 1382 1066 1383 1070
rect 1387 1066 1388 1070
rect 1382 1065 1388 1066
rect 1510 1070 1516 1071
rect 1510 1066 1511 1070
rect 1515 1066 1516 1070
rect 1510 1065 1516 1066
rect 1638 1070 1644 1071
rect 1638 1066 1639 1070
rect 1643 1066 1644 1070
rect 1638 1065 1644 1066
rect 1750 1070 1756 1071
rect 1750 1066 1751 1070
rect 1755 1066 1756 1070
rect 1750 1065 1756 1066
rect 144 1043 146 1065
rect 256 1043 258 1065
rect 392 1043 394 1065
rect 528 1043 530 1065
rect 656 1043 658 1065
rect 784 1043 786 1065
rect 904 1043 906 1065
rect 1024 1043 1026 1065
rect 1144 1043 1146 1065
rect 1264 1043 1266 1065
rect 1384 1043 1386 1065
rect 1512 1043 1514 1065
rect 1640 1043 1642 1065
rect 1752 1043 1754 1065
rect 1832 1043 1834 1083
rect 1870 1082 1876 1083
rect 1894 1084 1900 1085
rect 1872 1063 1874 1082
rect 1894 1080 1895 1084
rect 1899 1080 1900 1084
rect 1894 1079 1900 1080
rect 2118 1084 2124 1085
rect 2118 1080 2119 1084
rect 2123 1080 2124 1084
rect 2118 1079 2124 1080
rect 2350 1084 2356 1085
rect 2350 1080 2351 1084
rect 2355 1080 2356 1084
rect 2350 1079 2356 1080
rect 2566 1084 2572 1085
rect 2566 1080 2567 1084
rect 2571 1080 2572 1084
rect 2566 1079 2572 1080
rect 2766 1084 2772 1085
rect 2766 1080 2767 1084
rect 2771 1080 2772 1084
rect 2766 1079 2772 1080
rect 2958 1084 2964 1085
rect 2958 1080 2959 1084
rect 2963 1080 2964 1084
rect 2958 1079 2964 1080
rect 3150 1084 3156 1085
rect 3150 1080 3151 1084
rect 3155 1080 3156 1084
rect 3150 1079 3156 1080
rect 3334 1084 3340 1085
rect 3334 1080 3335 1084
rect 3339 1080 3340 1084
rect 3334 1079 3340 1080
rect 3502 1084 3508 1085
rect 3502 1080 3503 1084
rect 3507 1080 3508 1084
rect 3590 1083 3591 1087
rect 3595 1083 3596 1087
rect 3590 1082 3596 1083
rect 3502 1079 3508 1080
rect 1896 1063 1898 1079
rect 2120 1063 2122 1079
rect 2352 1063 2354 1079
rect 2568 1063 2570 1079
rect 2768 1063 2770 1079
rect 2960 1063 2962 1079
rect 3152 1063 3154 1079
rect 3336 1063 3338 1079
rect 3504 1063 3506 1079
rect 3592 1063 3594 1082
rect 1871 1062 1875 1063
rect 1871 1057 1875 1058
rect 1895 1062 1899 1063
rect 1895 1057 1899 1058
rect 2015 1062 2019 1063
rect 2015 1057 2019 1058
rect 2119 1062 2123 1063
rect 2119 1057 2123 1058
rect 2167 1062 2171 1063
rect 2167 1057 2171 1058
rect 2327 1062 2331 1063
rect 2327 1057 2331 1058
rect 2351 1062 2355 1063
rect 2351 1057 2355 1058
rect 2487 1062 2491 1063
rect 2487 1057 2491 1058
rect 2567 1062 2571 1063
rect 2567 1057 2571 1058
rect 2639 1062 2643 1063
rect 2639 1057 2643 1058
rect 2767 1062 2771 1063
rect 2767 1057 2771 1058
rect 2791 1062 2795 1063
rect 2791 1057 2795 1058
rect 2935 1062 2939 1063
rect 2935 1057 2939 1058
rect 2959 1062 2963 1063
rect 2959 1057 2963 1058
rect 3079 1062 3083 1063
rect 3079 1057 3083 1058
rect 3151 1062 3155 1063
rect 3151 1057 3155 1058
rect 3223 1062 3227 1063
rect 3223 1057 3227 1058
rect 3335 1062 3339 1063
rect 3335 1057 3339 1058
rect 3375 1062 3379 1063
rect 3375 1057 3379 1058
rect 3503 1062 3507 1063
rect 3503 1057 3507 1058
rect 3591 1062 3595 1063
rect 3591 1057 3595 1058
rect 111 1042 115 1043
rect 111 1037 115 1038
rect 143 1042 147 1043
rect 143 1037 147 1038
rect 239 1042 243 1043
rect 239 1037 243 1038
rect 255 1042 259 1043
rect 255 1037 259 1038
rect 359 1042 363 1043
rect 359 1037 363 1038
rect 391 1042 395 1043
rect 391 1037 395 1038
rect 471 1042 475 1043
rect 471 1037 475 1038
rect 527 1042 531 1043
rect 527 1037 531 1038
rect 575 1042 579 1043
rect 575 1037 579 1038
rect 655 1042 659 1043
rect 655 1037 659 1038
rect 671 1042 675 1043
rect 671 1037 675 1038
rect 767 1042 771 1043
rect 767 1037 771 1038
rect 783 1042 787 1043
rect 783 1037 787 1038
rect 855 1042 859 1043
rect 855 1037 859 1038
rect 903 1042 907 1043
rect 903 1037 907 1038
rect 943 1042 947 1043
rect 943 1037 947 1038
rect 1023 1042 1027 1043
rect 1023 1037 1027 1038
rect 1031 1042 1035 1043
rect 1031 1037 1035 1038
rect 1127 1042 1131 1043
rect 1127 1037 1131 1038
rect 1143 1042 1147 1043
rect 1143 1037 1147 1038
rect 1223 1042 1227 1043
rect 1223 1037 1227 1038
rect 1263 1042 1267 1043
rect 1263 1037 1267 1038
rect 1383 1042 1387 1043
rect 1383 1037 1387 1038
rect 1511 1042 1515 1043
rect 1511 1037 1515 1038
rect 1639 1042 1643 1043
rect 1639 1037 1643 1038
rect 1751 1042 1755 1043
rect 1751 1037 1755 1038
rect 1831 1042 1835 1043
rect 1872 1038 1874 1057
rect 1896 1041 1898 1057
rect 2016 1041 2018 1057
rect 2168 1041 2170 1057
rect 2328 1041 2330 1057
rect 2488 1041 2490 1057
rect 2640 1041 2642 1057
rect 2792 1041 2794 1057
rect 2936 1041 2938 1057
rect 3080 1041 3082 1057
rect 3224 1041 3226 1057
rect 3376 1041 3378 1057
rect 3504 1041 3506 1057
rect 1894 1040 1900 1041
rect 1831 1037 1835 1038
rect 1870 1037 1876 1038
rect 112 1009 114 1037
rect 144 1027 146 1037
rect 240 1027 242 1037
rect 360 1027 362 1037
rect 472 1027 474 1037
rect 576 1027 578 1037
rect 672 1027 674 1037
rect 768 1027 770 1037
rect 856 1027 858 1037
rect 944 1027 946 1037
rect 1032 1027 1034 1037
rect 1128 1027 1130 1037
rect 1224 1027 1226 1037
rect 142 1026 148 1027
rect 142 1022 143 1026
rect 147 1022 148 1026
rect 142 1021 148 1022
rect 238 1026 244 1027
rect 238 1022 239 1026
rect 243 1022 244 1026
rect 238 1021 244 1022
rect 358 1026 364 1027
rect 358 1022 359 1026
rect 363 1022 364 1026
rect 358 1021 364 1022
rect 470 1026 476 1027
rect 470 1022 471 1026
rect 475 1022 476 1026
rect 470 1021 476 1022
rect 574 1026 580 1027
rect 574 1022 575 1026
rect 579 1022 580 1026
rect 574 1021 580 1022
rect 670 1026 676 1027
rect 670 1022 671 1026
rect 675 1022 676 1026
rect 670 1021 676 1022
rect 766 1026 772 1027
rect 766 1022 767 1026
rect 771 1022 772 1026
rect 766 1021 772 1022
rect 854 1026 860 1027
rect 854 1022 855 1026
rect 859 1022 860 1026
rect 854 1021 860 1022
rect 942 1026 948 1027
rect 942 1022 943 1026
rect 947 1022 948 1026
rect 942 1021 948 1022
rect 1030 1026 1036 1027
rect 1030 1022 1031 1026
rect 1035 1022 1036 1026
rect 1030 1021 1036 1022
rect 1126 1026 1132 1027
rect 1126 1022 1127 1026
rect 1131 1022 1132 1026
rect 1126 1021 1132 1022
rect 1222 1026 1228 1027
rect 1222 1022 1223 1026
rect 1227 1022 1228 1026
rect 1222 1021 1228 1022
rect 1832 1009 1834 1037
rect 1870 1033 1871 1037
rect 1875 1033 1876 1037
rect 1894 1036 1895 1040
rect 1899 1036 1900 1040
rect 1894 1035 1900 1036
rect 2014 1040 2020 1041
rect 2014 1036 2015 1040
rect 2019 1036 2020 1040
rect 2014 1035 2020 1036
rect 2166 1040 2172 1041
rect 2166 1036 2167 1040
rect 2171 1036 2172 1040
rect 2166 1035 2172 1036
rect 2326 1040 2332 1041
rect 2326 1036 2327 1040
rect 2331 1036 2332 1040
rect 2326 1035 2332 1036
rect 2486 1040 2492 1041
rect 2486 1036 2487 1040
rect 2491 1036 2492 1040
rect 2486 1035 2492 1036
rect 2638 1040 2644 1041
rect 2638 1036 2639 1040
rect 2643 1036 2644 1040
rect 2638 1035 2644 1036
rect 2790 1040 2796 1041
rect 2790 1036 2791 1040
rect 2795 1036 2796 1040
rect 2790 1035 2796 1036
rect 2934 1040 2940 1041
rect 2934 1036 2935 1040
rect 2939 1036 2940 1040
rect 2934 1035 2940 1036
rect 3078 1040 3084 1041
rect 3078 1036 3079 1040
rect 3083 1036 3084 1040
rect 3078 1035 3084 1036
rect 3222 1040 3228 1041
rect 3222 1036 3223 1040
rect 3227 1036 3228 1040
rect 3222 1035 3228 1036
rect 3374 1040 3380 1041
rect 3374 1036 3375 1040
rect 3379 1036 3380 1040
rect 3374 1035 3380 1036
rect 3502 1040 3508 1041
rect 3502 1036 3503 1040
rect 3507 1036 3508 1040
rect 3592 1038 3594 1057
rect 3502 1035 3508 1036
rect 3590 1037 3596 1038
rect 1870 1032 1876 1033
rect 3590 1033 3591 1037
rect 3595 1033 3596 1037
rect 3590 1032 3596 1033
rect 1870 1020 1876 1021
rect 1870 1016 1871 1020
rect 1875 1016 1876 1020
rect 1870 1015 1876 1016
rect 3590 1020 3596 1021
rect 3590 1016 3591 1020
rect 3595 1016 3596 1020
rect 3590 1015 3596 1016
rect 110 1008 116 1009
rect 110 1004 111 1008
rect 115 1004 116 1008
rect 110 1003 116 1004
rect 1830 1008 1836 1009
rect 1830 1004 1831 1008
rect 1835 1004 1836 1008
rect 1830 1003 1836 1004
rect 110 991 116 992
rect 110 987 111 991
rect 115 987 116 991
rect 1830 991 1836 992
rect 110 986 116 987
rect 134 988 140 989
rect 112 955 114 986
rect 134 984 135 988
rect 139 984 140 988
rect 134 983 140 984
rect 230 988 236 989
rect 230 984 231 988
rect 235 984 236 988
rect 230 983 236 984
rect 350 988 356 989
rect 350 984 351 988
rect 355 984 356 988
rect 350 983 356 984
rect 462 988 468 989
rect 462 984 463 988
rect 467 984 468 988
rect 462 983 468 984
rect 566 988 572 989
rect 566 984 567 988
rect 571 984 572 988
rect 566 983 572 984
rect 662 988 668 989
rect 662 984 663 988
rect 667 984 668 988
rect 662 983 668 984
rect 758 988 764 989
rect 758 984 759 988
rect 763 984 764 988
rect 758 983 764 984
rect 846 988 852 989
rect 846 984 847 988
rect 851 984 852 988
rect 846 983 852 984
rect 934 988 940 989
rect 934 984 935 988
rect 939 984 940 988
rect 934 983 940 984
rect 1022 988 1028 989
rect 1022 984 1023 988
rect 1027 984 1028 988
rect 1022 983 1028 984
rect 1118 988 1124 989
rect 1118 984 1119 988
rect 1123 984 1124 988
rect 1118 983 1124 984
rect 1214 988 1220 989
rect 1214 984 1215 988
rect 1219 984 1220 988
rect 1830 987 1831 991
rect 1835 987 1836 991
rect 1830 986 1836 987
rect 1214 983 1220 984
rect 136 955 138 983
rect 232 955 234 983
rect 352 955 354 983
rect 464 955 466 983
rect 568 955 570 983
rect 664 955 666 983
rect 760 955 762 983
rect 848 955 850 983
rect 936 955 938 983
rect 1024 955 1026 983
rect 1120 955 1122 983
rect 1216 955 1218 983
rect 1832 955 1834 986
rect 1872 983 1874 1015
rect 1902 1002 1908 1003
rect 1902 998 1903 1002
rect 1907 998 1908 1002
rect 1902 997 1908 998
rect 2022 1002 2028 1003
rect 2022 998 2023 1002
rect 2027 998 2028 1002
rect 2022 997 2028 998
rect 2174 1002 2180 1003
rect 2174 998 2175 1002
rect 2179 998 2180 1002
rect 2174 997 2180 998
rect 2334 1002 2340 1003
rect 2334 998 2335 1002
rect 2339 998 2340 1002
rect 2334 997 2340 998
rect 2494 1002 2500 1003
rect 2494 998 2495 1002
rect 2499 998 2500 1002
rect 2494 997 2500 998
rect 2646 1002 2652 1003
rect 2646 998 2647 1002
rect 2651 998 2652 1002
rect 2646 997 2652 998
rect 2798 1002 2804 1003
rect 2798 998 2799 1002
rect 2803 998 2804 1002
rect 2798 997 2804 998
rect 2942 1002 2948 1003
rect 2942 998 2943 1002
rect 2947 998 2948 1002
rect 2942 997 2948 998
rect 3086 1002 3092 1003
rect 3086 998 3087 1002
rect 3091 998 3092 1002
rect 3086 997 3092 998
rect 3230 1002 3236 1003
rect 3230 998 3231 1002
rect 3235 998 3236 1002
rect 3230 997 3236 998
rect 3382 1002 3388 1003
rect 3382 998 3383 1002
rect 3387 998 3388 1002
rect 3382 997 3388 998
rect 3510 1002 3516 1003
rect 3510 998 3511 1002
rect 3515 998 3516 1002
rect 3510 997 3516 998
rect 1904 983 1906 997
rect 2024 983 2026 997
rect 2176 983 2178 997
rect 2336 983 2338 997
rect 2496 983 2498 997
rect 2648 983 2650 997
rect 2800 983 2802 997
rect 2944 983 2946 997
rect 3088 983 3090 997
rect 3232 983 3234 997
rect 3384 983 3386 997
rect 3512 983 3514 997
rect 3592 983 3594 1015
rect 1871 982 1875 983
rect 1871 977 1875 978
rect 1903 982 1907 983
rect 1903 977 1907 978
rect 1983 982 1987 983
rect 1983 977 1987 978
rect 2023 982 2027 983
rect 2023 977 2027 978
rect 2079 982 2083 983
rect 2079 977 2083 978
rect 2175 982 2179 983
rect 2175 977 2179 978
rect 2199 982 2203 983
rect 2199 977 2203 978
rect 2335 982 2339 983
rect 2335 977 2339 978
rect 2479 982 2483 983
rect 2479 977 2483 978
rect 2495 982 2499 983
rect 2495 977 2499 978
rect 2631 982 2635 983
rect 2631 977 2635 978
rect 2647 982 2651 983
rect 2647 977 2651 978
rect 2791 982 2795 983
rect 2791 977 2795 978
rect 2799 982 2803 983
rect 2799 977 2803 978
rect 2943 982 2947 983
rect 2943 977 2947 978
rect 2967 982 2971 983
rect 2967 977 2971 978
rect 3087 982 3091 983
rect 3087 977 3091 978
rect 3151 982 3155 983
rect 3151 977 3155 978
rect 3231 982 3235 983
rect 3231 977 3235 978
rect 3343 982 3347 983
rect 3343 977 3347 978
rect 3383 982 3387 983
rect 3383 977 3387 978
rect 3511 982 3515 983
rect 3511 977 3515 978
rect 3591 982 3595 983
rect 3591 977 3595 978
rect 111 954 115 955
rect 111 949 115 950
rect 135 954 139 955
rect 135 949 139 950
rect 231 954 235 955
rect 231 949 235 950
rect 263 954 267 955
rect 263 949 267 950
rect 351 954 355 955
rect 351 949 355 950
rect 415 954 419 955
rect 415 949 419 950
rect 463 954 467 955
rect 463 949 467 950
rect 559 954 563 955
rect 559 949 563 950
rect 567 954 571 955
rect 567 949 571 950
rect 663 954 667 955
rect 663 949 667 950
rect 703 954 707 955
rect 703 949 707 950
rect 759 954 763 955
rect 759 949 763 950
rect 839 954 843 955
rect 839 949 843 950
rect 847 954 851 955
rect 847 949 851 950
rect 935 954 939 955
rect 935 949 939 950
rect 975 954 979 955
rect 975 949 979 950
rect 1023 954 1027 955
rect 1023 949 1027 950
rect 1103 954 1107 955
rect 1103 949 1107 950
rect 1119 954 1123 955
rect 1119 949 1123 950
rect 1215 954 1219 955
rect 1215 949 1219 950
rect 1223 954 1227 955
rect 1223 949 1227 950
rect 1335 954 1339 955
rect 1335 949 1339 950
rect 1439 954 1443 955
rect 1439 949 1443 950
rect 1543 954 1547 955
rect 1543 949 1547 950
rect 1655 954 1659 955
rect 1655 949 1659 950
rect 1743 954 1747 955
rect 1743 949 1747 950
rect 1831 954 1835 955
rect 1831 949 1835 950
rect 1872 949 1874 977
rect 1904 967 1906 977
rect 1984 967 1986 977
rect 2080 967 2082 977
rect 2200 967 2202 977
rect 2336 967 2338 977
rect 2480 967 2482 977
rect 2632 967 2634 977
rect 2792 967 2794 977
rect 2968 967 2970 977
rect 3152 967 3154 977
rect 3344 967 3346 977
rect 3512 967 3514 977
rect 1902 966 1908 967
rect 1902 962 1903 966
rect 1907 962 1908 966
rect 1902 961 1908 962
rect 1982 966 1988 967
rect 1982 962 1983 966
rect 1987 962 1988 966
rect 1982 961 1988 962
rect 2078 966 2084 967
rect 2078 962 2079 966
rect 2083 962 2084 966
rect 2078 961 2084 962
rect 2198 966 2204 967
rect 2198 962 2199 966
rect 2203 962 2204 966
rect 2198 961 2204 962
rect 2334 966 2340 967
rect 2334 962 2335 966
rect 2339 962 2340 966
rect 2334 961 2340 962
rect 2478 966 2484 967
rect 2478 962 2479 966
rect 2483 962 2484 966
rect 2478 961 2484 962
rect 2630 966 2636 967
rect 2630 962 2631 966
rect 2635 962 2636 966
rect 2630 961 2636 962
rect 2790 966 2796 967
rect 2790 962 2791 966
rect 2795 962 2796 966
rect 2790 961 2796 962
rect 2966 966 2972 967
rect 2966 962 2967 966
rect 2971 962 2972 966
rect 2966 961 2972 962
rect 3150 966 3156 967
rect 3150 962 3151 966
rect 3155 962 3156 966
rect 3150 961 3156 962
rect 3342 966 3348 967
rect 3342 962 3343 966
rect 3347 962 3348 966
rect 3342 961 3348 962
rect 3510 966 3516 967
rect 3510 962 3511 966
rect 3515 962 3516 966
rect 3510 961 3516 962
rect 3592 949 3594 977
rect 112 930 114 949
rect 136 933 138 949
rect 264 933 266 949
rect 416 933 418 949
rect 560 933 562 949
rect 704 933 706 949
rect 840 933 842 949
rect 976 933 978 949
rect 1104 933 1106 949
rect 1224 933 1226 949
rect 1336 933 1338 949
rect 1440 933 1442 949
rect 1544 933 1546 949
rect 1656 933 1658 949
rect 1744 933 1746 949
rect 134 932 140 933
rect 110 929 116 930
rect 110 925 111 929
rect 115 925 116 929
rect 134 928 135 932
rect 139 928 140 932
rect 134 927 140 928
rect 262 932 268 933
rect 262 928 263 932
rect 267 928 268 932
rect 262 927 268 928
rect 414 932 420 933
rect 414 928 415 932
rect 419 928 420 932
rect 414 927 420 928
rect 558 932 564 933
rect 558 928 559 932
rect 563 928 564 932
rect 558 927 564 928
rect 702 932 708 933
rect 702 928 703 932
rect 707 928 708 932
rect 702 927 708 928
rect 838 932 844 933
rect 838 928 839 932
rect 843 928 844 932
rect 838 927 844 928
rect 974 932 980 933
rect 974 928 975 932
rect 979 928 980 932
rect 974 927 980 928
rect 1102 932 1108 933
rect 1102 928 1103 932
rect 1107 928 1108 932
rect 1102 927 1108 928
rect 1222 932 1228 933
rect 1222 928 1223 932
rect 1227 928 1228 932
rect 1222 927 1228 928
rect 1334 932 1340 933
rect 1334 928 1335 932
rect 1339 928 1340 932
rect 1334 927 1340 928
rect 1438 932 1444 933
rect 1438 928 1439 932
rect 1443 928 1444 932
rect 1438 927 1444 928
rect 1542 932 1548 933
rect 1542 928 1543 932
rect 1547 928 1548 932
rect 1542 927 1548 928
rect 1654 932 1660 933
rect 1654 928 1655 932
rect 1659 928 1660 932
rect 1654 927 1660 928
rect 1742 932 1748 933
rect 1742 928 1743 932
rect 1747 928 1748 932
rect 1832 930 1834 949
rect 1870 948 1876 949
rect 1870 944 1871 948
rect 1875 944 1876 948
rect 1870 943 1876 944
rect 3590 948 3596 949
rect 3590 944 3591 948
rect 3595 944 3596 948
rect 3590 943 3596 944
rect 1870 931 1876 932
rect 1742 927 1748 928
rect 1830 929 1836 930
rect 110 924 116 925
rect 1830 925 1831 929
rect 1835 925 1836 929
rect 1870 927 1871 931
rect 1875 927 1876 931
rect 3590 931 3596 932
rect 1870 926 1876 927
rect 1894 928 1900 929
rect 1830 924 1836 925
rect 110 912 116 913
rect 110 908 111 912
rect 115 908 116 912
rect 110 907 116 908
rect 1830 912 1836 913
rect 1830 908 1831 912
rect 1835 908 1836 912
rect 1830 907 1836 908
rect 112 875 114 907
rect 142 894 148 895
rect 142 890 143 894
rect 147 890 148 894
rect 142 889 148 890
rect 270 894 276 895
rect 270 890 271 894
rect 275 890 276 894
rect 270 889 276 890
rect 422 894 428 895
rect 422 890 423 894
rect 427 890 428 894
rect 422 889 428 890
rect 566 894 572 895
rect 566 890 567 894
rect 571 890 572 894
rect 566 889 572 890
rect 710 894 716 895
rect 710 890 711 894
rect 715 890 716 894
rect 710 889 716 890
rect 846 894 852 895
rect 846 890 847 894
rect 851 890 852 894
rect 846 889 852 890
rect 982 894 988 895
rect 982 890 983 894
rect 987 890 988 894
rect 982 889 988 890
rect 1110 894 1116 895
rect 1110 890 1111 894
rect 1115 890 1116 894
rect 1110 889 1116 890
rect 1230 894 1236 895
rect 1230 890 1231 894
rect 1235 890 1236 894
rect 1230 889 1236 890
rect 1342 894 1348 895
rect 1342 890 1343 894
rect 1347 890 1348 894
rect 1342 889 1348 890
rect 1446 894 1452 895
rect 1446 890 1447 894
rect 1451 890 1452 894
rect 1446 889 1452 890
rect 1550 894 1556 895
rect 1550 890 1551 894
rect 1555 890 1556 894
rect 1550 889 1556 890
rect 1662 894 1668 895
rect 1662 890 1663 894
rect 1667 890 1668 894
rect 1662 889 1668 890
rect 1750 894 1756 895
rect 1750 890 1751 894
rect 1755 890 1756 894
rect 1750 889 1756 890
rect 144 875 146 889
rect 272 875 274 889
rect 424 875 426 889
rect 568 875 570 889
rect 712 875 714 889
rect 848 875 850 889
rect 984 875 986 889
rect 1112 875 1114 889
rect 1232 875 1234 889
rect 1344 875 1346 889
rect 1448 875 1450 889
rect 1552 875 1554 889
rect 1664 875 1666 889
rect 1752 875 1754 889
rect 1832 875 1834 907
rect 1872 895 1874 926
rect 1894 924 1895 928
rect 1899 924 1900 928
rect 1894 923 1900 924
rect 1974 928 1980 929
rect 1974 924 1975 928
rect 1979 924 1980 928
rect 1974 923 1980 924
rect 2070 928 2076 929
rect 2070 924 2071 928
rect 2075 924 2076 928
rect 2070 923 2076 924
rect 2190 928 2196 929
rect 2190 924 2191 928
rect 2195 924 2196 928
rect 2190 923 2196 924
rect 2326 928 2332 929
rect 2326 924 2327 928
rect 2331 924 2332 928
rect 2326 923 2332 924
rect 2470 928 2476 929
rect 2470 924 2471 928
rect 2475 924 2476 928
rect 2470 923 2476 924
rect 2622 928 2628 929
rect 2622 924 2623 928
rect 2627 924 2628 928
rect 2622 923 2628 924
rect 2782 928 2788 929
rect 2782 924 2783 928
rect 2787 924 2788 928
rect 2782 923 2788 924
rect 2958 928 2964 929
rect 2958 924 2959 928
rect 2963 924 2964 928
rect 2958 923 2964 924
rect 3142 928 3148 929
rect 3142 924 3143 928
rect 3147 924 3148 928
rect 3142 923 3148 924
rect 3334 928 3340 929
rect 3334 924 3335 928
rect 3339 924 3340 928
rect 3334 923 3340 924
rect 3502 928 3508 929
rect 3502 924 3503 928
rect 3507 924 3508 928
rect 3590 927 3591 931
rect 3595 927 3596 931
rect 3590 926 3596 927
rect 3502 923 3508 924
rect 1896 895 1898 923
rect 1976 895 1978 923
rect 2072 895 2074 923
rect 2192 895 2194 923
rect 2328 895 2330 923
rect 2472 895 2474 923
rect 2624 895 2626 923
rect 2784 895 2786 923
rect 2960 895 2962 923
rect 3144 895 3146 923
rect 3336 895 3338 923
rect 3504 895 3506 923
rect 3592 895 3594 926
rect 1871 894 1875 895
rect 1871 889 1875 890
rect 1895 894 1899 895
rect 1895 889 1899 890
rect 1919 894 1923 895
rect 1919 889 1923 890
rect 1975 894 1979 895
rect 1975 889 1979 890
rect 2071 894 2075 895
rect 2071 889 2075 890
rect 2095 894 2099 895
rect 2095 889 2099 890
rect 2191 894 2195 895
rect 2191 889 2195 890
rect 2271 894 2275 895
rect 2271 889 2275 890
rect 2327 894 2331 895
rect 2327 889 2331 890
rect 2455 894 2459 895
rect 2455 889 2459 890
rect 2471 894 2475 895
rect 2471 889 2475 890
rect 2623 894 2627 895
rect 2623 889 2627 890
rect 2655 894 2659 895
rect 2655 889 2659 890
rect 2783 894 2787 895
rect 2783 889 2787 890
rect 2863 894 2867 895
rect 2863 889 2867 890
rect 2959 894 2963 895
rect 2959 889 2963 890
rect 3079 894 3083 895
rect 3079 889 3083 890
rect 3143 894 3147 895
rect 3143 889 3147 890
rect 3303 894 3307 895
rect 3303 889 3307 890
rect 3335 894 3339 895
rect 3335 889 3339 890
rect 3503 894 3507 895
rect 3503 889 3507 890
rect 3591 894 3595 895
rect 3591 889 3595 890
rect 111 874 115 875
rect 111 869 115 870
rect 143 874 147 875
rect 143 869 147 870
rect 247 874 251 875
rect 247 869 251 870
rect 271 874 275 875
rect 271 869 275 870
rect 383 874 387 875
rect 383 869 387 870
rect 423 874 427 875
rect 423 869 427 870
rect 519 874 523 875
rect 519 869 523 870
rect 567 874 571 875
rect 567 869 571 870
rect 663 874 667 875
rect 663 869 667 870
rect 711 874 715 875
rect 711 869 715 870
rect 815 874 819 875
rect 815 869 819 870
rect 847 874 851 875
rect 847 869 851 870
rect 959 874 963 875
rect 959 869 963 870
rect 983 874 987 875
rect 983 869 987 870
rect 1103 874 1107 875
rect 1103 869 1107 870
rect 1111 874 1115 875
rect 1111 869 1115 870
rect 1231 874 1235 875
rect 1231 869 1235 870
rect 1247 874 1251 875
rect 1247 869 1251 870
rect 1343 874 1347 875
rect 1343 869 1347 870
rect 1383 874 1387 875
rect 1383 869 1387 870
rect 1447 874 1451 875
rect 1447 869 1451 870
rect 1511 874 1515 875
rect 1511 869 1515 870
rect 1551 874 1555 875
rect 1551 869 1555 870
rect 1639 874 1643 875
rect 1639 869 1643 870
rect 1663 874 1667 875
rect 1663 869 1667 870
rect 1751 874 1755 875
rect 1751 869 1755 870
rect 1831 874 1835 875
rect 1872 870 1874 889
rect 1920 873 1922 889
rect 2096 873 2098 889
rect 2272 873 2274 889
rect 2456 873 2458 889
rect 2656 873 2658 889
rect 2864 873 2866 889
rect 3080 873 3082 889
rect 3304 873 3306 889
rect 3504 873 3506 889
rect 1918 872 1924 873
rect 1831 869 1835 870
rect 1870 869 1876 870
rect 112 841 114 869
rect 144 859 146 869
rect 248 859 250 869
rect 384 859 386 869
rect 520 859 522 869
rect 664 859 666 869
rect 816 859 818 869
rect 960 859 962 869
rect 1104 859 1106 869
rect 1248 859 1250 869
rect 1384 859 1386 869
rect 1512 859 1514 869
rect 1640 859 1642 869
rect 1752 859 1754 869
rect 142 858 148 859
rect 142 854 143 858
rect 147 854 148 858
rect 142 853 148 854
rect 246 858 252 859
rect 246 854 247 858
rect 251 854 252 858
rect 246 853 252 854
rect 382 858 388 859
rect 382 854 383 858
rect 387 854 388 858
rect 382 853 388 854
rect 518 858 524 859
rect 518 854 519 858
rect 523 854 524 858
rect 518 853 524 854
rect 662 858 668 859
rect 662 854 663 858
rect 667 854 668 858
rect 662 853 668 854
rect 814 858 820 859
rect 814 854 815 858
rect 819 854 820 858
rect 814 853 820 854
rect 958 858 964 859
rect 958 854 959 858
rect 963 854 964 858
rect 958 853 964 854
rect 1102 858 1108 859
rect 1102 854 1103 858
rect 1107 854 1108 858
rect 1102 853 1108 854
rect 1246 858 1252 859
rect 1246 854 1247 858
rect 1251 854 1252 858
rect 1246 853 1252 854
rect 1382 858 1388 859
rect 1382 854 1383 858
rect 1387 854 1388 858
rect 1382 853 1388 854
rect 1510 858 1516 859
rect 1510 854 1511 858
rect 1515 854 1516 858
rect 1510 853 1516 854
rect 1638 858 1644 859
rect 1638 854 1639 858
rect 1643 854 1644 858
rect 1638 853 1644 854
rect 1750 858 1756 859
rect 1750 854 1751 858
rect 1755 854 1756 858
rect 1750 853 1756 854
rect 1832 841 1834 869
rect 1870 865 1871 869
rect 1875 865 1876 869
rect 1918 868 1919 872
rect 1923 868 1924 872
rect 1918 867 1924 868
rect 2094 872 2100 873
rect 2094 868 2095 872
rect 2099 868 2100 872
rect 2094 867 2100 868
rect 2270 872 2276 873
rect 2270 868 2271 872
rect 2275 868 2276 872
rect 2270 867 2276 868
rect 2454 872 2460 873
rect 2454 868 2455 872
rect 2459 868 2460 872
rect 2454 867 2460 868
rect 2654 872 2660 873
rect 2654 868 2655 872
rect 2659 868 2660 872
rect 2654 867 2660 868
rect 2862 872 2868 873
rect 2862 868 2863 872
rect 2867 868 2868 872
rect 2862 867 2868 868
rect 3078 872 3084 873
rect 3078 868 3079 872
rect 3083 868 3084 872
rect 3078 867 3084 868
rect 3302 872 3308 873
rect 3302 868 3303 872
rect 3307 868 3308 872
rect 3302 867 3308 868
rect 3502 872 3508 873
rect 3502 868 3503 872
rect 3507 868 3508 872
rect 3592 870 3594 889
rect 3502 867 3508 868
rect 3590 869 3596 870
rect 1870 864 1876 865
rect 3590 865 3591 869
rect 3595 865 3596 869
rect 3590 864 3596 865
rect 1870 852 1876 853
rect 1870 848 1871 852
rect 1875 848 1876 852
rect 1870 847 1876 848
rect 3590 852 3596 853
rect 3590 848 3591 852
rect 3595 848 3596 852
rect 3590 847 3596 848
rect 110 840 116 841
rect 110 836 111 840
rect 115 836 116 840
rect 110 835 116 836
rect 1830 840 1836 841
rect 1830 836 1831 840
rect 1835 836 1836 840
rect 1830 835 1836 836
rect 110 823 116 824
rect 110 819 111 823
rect 115 819 116 823
rect 1830 823 1836 824
rect 110 818 116 819
rect 134 820 140 821
rect 112 787 114 818
rect 134 816 135 820
rect 139 816 140 820
rect 134 815 140 816
rect 238 820 244 821
rect 238 816 239 820
rect 243 816 244 820
rect 238 815 244 816
rect 374 820 380 821
rect 374 816 375 820
rect 379 816 380 820
rect 374 815 380 816
rect 510 820 516 821
rect 510 816 511 820
rect 515 816 516 820
rect 510 815 516 816
rect 654 820 660 821
rect 654 816 655 820
rect 659 816 660 820
rect 654 815 660 816
rect 806 820 812 821
rect 806 816 807 820
rect 811 816 812 820
rect 806 815 812 816
rect 950 820 956 821
rect 950 816 951 820
rect 955 816 956 820
rect 950 815 956 816
rect 1094 820 1100 821
rect 1094 816 1095 820
rect 1099 816 1100 820
rect 1094 815 1100 816
rect 1238 820 1244 821
rect 1238 816 1239 820
rect 1243 816 1244 820
rect 1238 815 1244 816
rect 1374 820 1380 821
rect 1374 816 1375 820
rect 1379 816 1380 820
rect 1374 815 1380 816
rect 1502 820 1508 821
rect 1502 816 1503 820
rect 1507 816 1508 820
rect 1502 815 1508 816
rect 1630 820 1636 821
rect 1630 816 1631 820
rect 1635 816 1636 820
rect 1630 815 1636 816
rect 1742 820 1748 821
rect 1742 816 1743 820
rect 1747 816 1748 820
rect 1830 819 1831 823
rect 1835 819 1836 823
rect 1872 819 1874 847
rect 1926 834 1932 835
rect 1926 830 1927 834
rect 1931 830 1932 834
rect 1926 829 1932 830
rect 2102 834 2108 835
rect 2102 830 2103 834
rect 2107 830 2108 834
rect 2102 829 2108 830
rect 2278 834 2284 835
rect 2278 830 2279 834
rect 2283 830 2284 834
rect 2278 829 2284 830
rect 2462 834 2468 835
rect 2462 830 2463 834
rect 2467 830 2468 834
rect 2462 829 2468 830
rect 2662 834 2668 835
rect 2662 830 2663 834
rect 2667 830 2668 834
rect 2662 829 2668 830
rect 2870 834 2876 835
rect 2870 830 2871 834
rect 2875 830 2876 834
rect 2870 829 2876 830
rect 3086 834 3092 835
rect 3086 830 3087 834
rect 3091 830 3092 834
rect 3086 829 3092 830
rect 3310 834 3316 835
rect 3310 830 3311 834
rect 3315 830 3316 834
rect 3310 829 3316 830
rect 3510 834 3516 835
rect 3510 830 3511 834
rect 3515 830 3516 834
rect 3510 829 3516 830
rect 1928 819 1930 829
rect 2104 819 2106 829
rect 2280 819 2282 829
rect 2464 819 2466 829
rect 2664 819 2666 829
rect 2872 819 2874 829
rect 3088 819 3090 829
rect 3312 819 3314 829
rect 3512 819 3514 829
rect 3592 819 3594 847
rect 1830 818 1836 819
rect 1871 818 1875 819
rect 1742 815 1748 816
rect 136 787 138 815
rect 240 787 242 815
rect 376 787 378 815
rect 512 787 514 815
rect 656 787 658 815
rect 808 787 810 815
rect 952 787 954 815
rect 1096 787 1098 815
rect 1240 787 1242 815
rect 1376 787 1378 815
rect 1504 787 1506 815
rect 1632 787 1634 815
rect 1744 787 1746 815
rect 1832 787 1834 818
rect 1871 813 1875 814
rect 1903 818 1907 819
rect 1903 813 1907 814
rect 1927 818 1931 819
rect 1927 813 1931 814
rect 2015 818 2019 819
rect 2015 813 2019 814
rect 2103 818 2107 819
rect 2103 813 2107 814
rect 2167 818 2171 819
rect 2167 813 2171 814
rect 2279 818 2283 819
rect 2279 813 2283 814
rect 2327 818 2331 819
rect 2327 813 2331 814
rect 2463 818 2467 819
rect 2463 813 2467 814
rect 2487 818 2491 819
rect 2487 813 2491 814
rect 2647 818 2651 819
rect 2647 813 2651 814
rect 2663 818 2667 819
rect 2663 813 2667 814
rect 2807 818 2811 819
rect 2807 813 2811 814
rect 2871 818 2875 819
rect 2871 813 2875 814
rect 2959 818 2963 819
rect 2959 813 2963 814
rect 3087 818 3091 819
rect 3087 813 3091 814
rect 3103 818 3107 819
rect 3103 813 3107 814
rect 3247 818 3251 819
rect 3247 813 3251 814
rect 3311 818 3315 819
rect 3311 813 3315 814
rect 3391 818 3395 819
rect 3391 813 3395 814
rect 3511 818 3515 819
rect 3511 813 3515 814
rect 3591 818 3595 819
rect 3591 813 3595 814
rect 111 786 115 787
rect 111 781 115 782
rect 135 786 139 787
rect 135 781 139 782
rect 215 786 219 787
rect 215 781 219 782
rect 239 786 243 787
rect 239 781 243 782
rect 303 786 307 787
rect 303 781 307 782
rect 375 786 379 787
rect 375 781 379 782
rect 415 786 419 787
rect 415 781 419 782
rect 511 786 515 787
rect 511 781 515 782
rect 543 786 547 787
rect 543 781 547 782
rect 655 786 659 787
rect 655 781 659 782
rect 687 786 691 787
rect 687 781 691 782
rect 807 786 811 787
rect 807 781 811 782
rect 839 786 843 787
rect 839 781 843 782
rect 951 786 955 787
rect 951 781 955 782
rect 991 786 995 787
rect 991 781 995 782
rect 1095 786 1099 787
rect 1095 781 1099 782
rect 1143 786 1147 787
rect 1143 781 1147 782
rect 1239 786 1243 787
rect 1239 781 1243 782
rect 1295 786 1299 787
rect 1295 781 1299 782
rect 1375 786 1379 787
rect 1375 781 1379 782
rect 1447 786 1451 787
rect 1447 781 1451 782
rect 1503 786 1507 787
rect 1503 781 1507 782
rect 1607 786 1611 787
rect 1607 781 1611 782
rect 1631 786 1635 787
rect 1631 781 1635 782
rect 1743 786 1747 787
rect 1743 781 1747 782
rect 1831 786 1835 787
rect 1872 785 1874 813
rect 1904 803 1906 813
rect 2016 803 2018 813
rect 2168 803 2170 813
rect 2328 803 2330 813
rect 2488 803 2490 813
rect 2648 803 2650 813
rect 2808 803 2810 813
rect 2960 803 2962 813
rect 3104 803 3106 813
rect 3248 803 3250 813
rect 3392 803 3394 813
rect 3512 803 3514 813
rect 1902 802 1908 803
rect 1902 798 1903 802
rect 1907 798 1908 802
rect 1902 797 1908 798
rect 2014 802 2020 803
rect 2014 798 2015 802
rect 2019 798 2020 802
rect 2014 797 2020 798
rect 2166 802 2172 803
rect 2166 798 2167 802
rect 2171 798 2172 802
rect 2166 797 2172 798
rect 2326 802 2332 803
rect 2326 798 2327 802
rect 2331 798 2332 802
rect 2326 797 2332 798
rect 2486 802 2492 803
rect 2486 798 2487 802
rect 2491 798 2492 802
rect 2486 797 2492 798
rect 2646 802 2652 803
rect 2646 798 2647 802
rect 2651 798 2652 802
rect 2646 797 2652 798
rect 2806 802 2812 803
rect 2806 798 2807 802
rect 2811 798 2812 802
rect 2806 797 2812 798
rect 2958 802 2964 803
rect 2958 798 2959 802
rect 2963 798 2964 802
rect 2958 797 2964 798
rect 3102 802 3108 803
rect 3102 798 3103 802
rect 3107 798 3108 802
rect 3102 797 3108 798
rect 3246 802 3252 803
rect 3246 798 3247 802
rect 3251 798 3252 802
rect 3246 797 3252 798
rect 3390 802 3396 803
rect 3390 798 3391 802
rect 3395 798 3396 802
rect 3390 797 3396 798
rect 3510 802 3516 803
rect 3510 798 3511 802
rect 3515 798 3516 802
rect 3510 797 3516 798
rect 3592 785 3594 813
rect 1831 781 1835 782
rect 1870 784 1876 785
rect 112 762 114 781
rect 136 765 138 781
rect 216 765 218 781
rect 304 765 306 781
rect 416 765 418 781
rect 544 765 546 781
rect 688 765 690 781
rect 840 765 842 781
rect 992 765 994 781
rect 1144 765 1146 781
rect 1296 765 1298 781
rect 1448 765 1450 781
rect 1608 765 1610 781
rect 134 764 140 765
rect 110 761 116 762
rect 110 757 111 761
rect 115 757 116 761
rect 134 760 135 764
rect 139 760 140 764
rect 134 759 140 760
rect 214 764 220 765
rect 214 760 215 764
rect 219 760 220 764
rect 214 759 220 760
rect 302 764 308 765
rect 302 760 303 764
rect 307 760 308 764
rect 302 759 308 760
rect 414 764 420 765
rect 414 760 415 764
rect 419 760 420 764
rect 414 759 420 760
rect 542 764 548 765
rect 542 760 543 764
rect 547 760 548 764
rect 542 759 548 760
rect 686 764 692 765
rect 686 760 687 764
rect 691 760 692 764
rect 686 759 692 760
rect 838 764 844 765
rect 838 760 839 764
rect 843 760 844 764
rect 838 759 844 760
rect 990 764 996 765
rect 990 760 991 764
rect 995 760 996 764
rect 990 759 996 760
rect 1142 764 1148 765
rect 1142 760 1143 764
rect 1147 760 1148 764
rect 1142 759 1148 760
rect 1294 764 1300 765
rect 1294 760 1295 764
rect 1299 760 1300 764
rect 1294 759 1300 760
rect 1446 764 1452 765
rect 1446 760 1447 764
rect 1451 760 1452 764
rect 1446 759 1452 760
rect 1606 764 1612 765
rect 1606 760 1607 764
rect 1611 760 1612 764
rect 1832 762 1834 781
rect 1870 780 1871 784
rect 1875 780 1876 784
rect 1870 779 1876 780
rect 3590 784 3596 785
rect 3590 780 3591 784
rect 3595 780 3596 784
rect 3590 779 3596 780
rect 1870 767 1876 768
rect 1870 763 1871 767
rect 1875 763 1876 767
rect 3590 767 3596 768
rect 1870 762 1876 763
rect 1894 764 1900 765
rect 1606 759 1612 760
rect 1830 761 1836 762
rect 110 756 116 757
rect 1830 757 1831 761
rect 1835 757 1836 761
rect 1830 756 1836 757
rect 110 744 116 745
rect 110 740 111 744
rect 115 740 116 744
rect 110 739 116 740
rect 1830 744 1836 745
rect 1830 740 1831 744
rect 1835 740 1836 744
rect 1872 743 1874 762
rect 1894 760 1895 764
rect 1899 760 1900 764
rect 1894 759 1900 760
rect 2006 764 2012 765
rect 2006 760 2007 764
rect 2011 760 2012 764
rect 2006 759 2012 760
rect 2158 764 2164 765
rect 2158 760 2159 764
rect 2163 760 2164 764
rect 2158 759 2164 760
rect 2318 764 2324 765
rect 2318 760 2319 764
rect 2323 760 2324 764
rect 2318 759 2324 760
rect 2478 764 2484 765
rect 2478 760 2479 764
rect 2483 760 2484 764
rect 2478 759 2484 760
rect 2638 764 2644 765
rect 2638 760 2639 764
rect 2643 760 2644 764
rect 2638 759 2644 760
rect 2798 764 2804 765
rect 2798 760 2799 764
rect 2803 760 2804 764
rect 2798 759 2804 760
rect 2950 764 2956 765
rect 2950 760 2951 764
rect 2955 760 2956 764
rect 2950 759 2956 760
rect 3094 764 3100 765
rect 3094 760 3095 764
rect 3099 760 3100 764
rect 3094 759 3100 760
rect 3238 764 3244 765
rect 3238 760 3239 764
rect 3243 760 3244 764
rect 3238 759 3244 760
rect 3382 764 3388 765
rect 3382 760 3383 764
rect 3387 760 3388 764
rect 3382 759 3388 760
rect 3502 764 3508 765
rect 3502 760 3503 764
rect 3507 760 3508 764
rect 3590 763 3591 767
rect 3595 763 3596 767
rect 3590 762 3596 763
rect 3502 759 3508 760
rect 1896 743 1898 759
rect 2008 743 2010 759
rect 2160 743 2162 759
rect 2320 743 2322 759
rect 2480 743 2482 759
rect 2640 743 2642 759
rect 2800 743 2802 759
rect 2952 743 2954 759
rect 3096 743 3098 759
rect 3240 743 3242 759
rect 3384 743 3386 759
rect 3504 743 3506 759
rect 3592 743 3594 762
rect 1830 739 1836 740
rect 1871 742 1875 743
rect 112 703 114 739
rect 142 726 148 727
rect 142 722 143 726
rect 147 722 148 726
rect 142 721 148 722
rect 222 726 228 727
rect 222 722 223 726
rect 227 722 228 726
rect 222 721 228 722
rect 310 726 316 727
rect 310 722 311 726
rect 315 722 316 726
rect 310 721 316 722
rect 422 726 428 727
rect 422 722 423 726
rect 427 722 428 726
rect 422 721 428 722
rect 550 726 556 727
rect 550 722 551 726
rect 555 722 556 726
rect 550 721 556 722
rect 694 726 700 727
rect 694 722 695 726
rect 699 722 700 726
rect 694 721 700 722
rect 846 726 852 727
rect 846 722 847 726
rect 851 722 852 726
rect 846 721 852 722
rect 998 726 1004 727
rect 998 722 999 726
rect 1003 722 1004 726
rect 998 721 1004 722
rect 1150 726 1156 727
rect 1150 722 1151 726
rect 1155 722 1156 726
rect 1150 721 1156 722
rect 1302 726 1308 727
rect 1302 722 1303 726
rect 1307 722 1308 726
rect 1302 721 1308 722
rect 1454 726 1460 727
rect 1454 722 1455 726
rect 1459 722 1460 726
rect 1454 721 1460 722
rect 1614 726 1620 727
rect 1614 722 1615 726
rect 1619 722 1620 726
rect 1614 721 1620 722
rect 144 703 146 721
rect 224 703 226 721
rect 312 703 314 721
rect 424 703 426 721
rect 552 703 554 721
rect 696 703 698 721
rect 848 703 850 721
rect 1000 703 1002 721
rect 1152 703 1154 721
rect 1304 703 1306 721
rect 1456 703 1458 721
rect 1616 703 1618 721
rect 1832 703 1834 739
rect 1871 737 1875 738
rect 1895 742 1899 743
rect 1895 737 1899 738
rect 1967 742 1971 743
rect 1967 737 1971 738
rect 2007 742 2011 743
rect 2007 737 2011 738
rect 2063 742 2067 743
rect 2063 737 2067 738
rect 2159 742 2163 743
rect 2159 737 2163 738
rect 2175 742 2179 743
rect 2175 737 2179 738
rect 2303 742 2307 743
rect 2303 737 2307 738
rect 2319 742 2323 743
rect 2319 737 2323 738
rect 2447 742 2451 743
rect 2447 737 2451 738
rect 2479 742 2483 743
rect 2479 737 2483 738
rect 2599 742 2603 743
rect 2599 737 2603 738
rect 2639 742 2643 743
rect 2639 737 2643 738
rect 2751 742 2755 743
rect 2751 737 2755 738
rect 2799 742 2803 743
rect 2799 737 2803 738
rect 2903 742 2907 743
rect 2903 737 2907 738
rect 2951 742 2955 743
rect 2951 737 2955 738
rect 3055 742 3059 743
rect 3055 737 3059 738
rect 3095 742 3099 743
rect 3095 737 3099 738
rect 3207 742 3211 743
rect 3207 737 3211 738
rect 3239 742 3243 743
rect 3239 737 3243 738
rect 3359 742 3363 743
rect 3359 737 3363 738
rect 3383 742 3387 743
rect 3383 737 3387 738
rect 3503 742 3507 743
rect 3503 737 3507 738
rect 3591 742 3595 743
rect 3591 737 3595 738
rect 1872 718 1874 737
rect 1968 721 1970 737
rect 2064 721 2066 737
rect 2176 721 2178 737
rect 2304 721 2306 737
rect 2448 721 2450 737
rect 2600 721 2602 737
rect 2752 721 2754 737
rect 2904 721 2906 737
rect 3056 721 3058 737
rect 3208 721 3210 737
rect 3360 721 3362 737
rect 3504 721 3506 737
rect 1966 720 1972 721
rect 1870 717 1876 718
rect 1870 713 1871 717
rect 1875 713 1876 717
rect 1966 716 1967 720
rect 1971 716 1972 720
rect 1966 715 1972 716
rect 2062 720 2068 721
rect 2062 716 2063 720
rect 2067 716 2068 720
rect 2062 715 2068 716
rect 2174 720 2180 721
rect 2174 716 2175 720
rect 2179 716 2180 720
rect 2174 715 2180 716
rect 2302 720 2308 721
rect 2302 716 2303 720
rect 2307 716 2308 720
rect 2302 715 2308 716
rect 2446 720 2452 721
rect 2446 716 2447 720
rect 2451 716 2452 720
rect 2446 715 2452 716
rect 2598 720 2604 721
rect 2598 716 2599 720
rect 2603 716 2604 720
rect 2598 715 2604 716
rect 2750 720 2756 721
rect 2750 716 2751 720
rect 2755 716 2756 720
rect 2750 715 2756 716
rect 2902 720 2908 721
rect 2902 716 2903 720
rect 2907 716 2908 720
rect 2902 715 2908 716
rect 3054 720 3060 721
rect 3054 716 3055 720
rect 3059 716 3060 720
rect 3054 715 3060 716
rect 3206 720 3212 721
rect 3206 716 3207 720
rect 3211 716 3212 720
rect 3206 715 3212 716
rect 3358 720 3364 721
rect 3358 716 3359 720
rect 3363 716 3364 720
rect 3358 715 3364 716
rect 3502 720 3508 721
rect 3502 716 3503 720
rect 3507 716 3508 720
rect 3592 718 3594 737
rect 3502 715 3508 716
rect 3590 717 3596 718
rect 1870 712 1876 713
rect 3590 713 3591 717
rect 3595 713 3596 717
rect 3590 712 3596 713
rect 111 702 115 703
rect 111 697 115 698
rect 143 702 147 703
rect 143 697 147 698
rect 223 702 227 703
rect 223 697 227 698
rect 231 702 235 703
rect 231 697 235 698
rect 311 702 315 703
rect 311 697 315 698
rect 319 702 323 703
rect 319 697 323 698
rect 423 702 427 703
rect 423 697 427 698
rect 543 702 547 703
rect 543 697 547 698
rect 551 702 555 703
rect 551 697 555 698
rect 679 702 683 703
rect 679 697 683 698
rect 695 702 699 703
rect 695 697 699 698
rect 815 702 819 703
rect 815 697 819 698
rect 847 702 851 703
rect 847 697 851 698
rect 951 702 955 703
rect 951 697 955 698
rect 999 702 1003 703
rect 999 697 1003 698
rect 1087 702 1091 703
rect 1087 697 1091 698
rect 1151 702 1155 703
rect 1151 697 1155 698
rect 1215 702 1219 703
rect 1215 697 1219 698
rect 1303 702 1307 703
rect 1303 697 1307 698
rect 1335 702 1339 703
rect 1335 697 1339 698
rect 1455 702 1459 703
rect 1455 697 1459 698
rect 1583 702 1587 703
rect 1583 697 1587 698
rect 1615 702 1619 703
rect 1615 697 1619 698
rect 1831 702 1835 703
rect 1831 697 1835 698
rect 1870 700 1876 701
rect 112 669 114 697
rect 232 687 234 697
rect 320 687 322 697
rect 424 687 426 697
rect 544 687 546 697
rect 680 687 682 697
rect 816 687 818 697
rect 952 687 954 697
rect 1088 687 1090 697
rect 1216 687 1218 697
rect 1336 687 1338 697
rect 1456 687 1458 697
rect 1584 687 1586 697
rect 230 686 236 687
rect 230 682 231 686
rect 235 682 236 686
rect 230 681 236 682
rect 318 686 324 687
rect 318 682 319 686
rect 323 682 324 686
rect 318 681 324 682
rect 422 686 428 687
rect 422 682 423 686
rect 427 682 428 686
rect 422 681 428 682
rect 542 686 548 687
rect 542 682 543 686
rect 547 682 548 686
rect 542 681 548 682
rect 678 686 684 687
rect 678 682 679 686
rect 683 682 684 686
rect 678 681 684 682
rect 814 686 820 687
rect 814 682 815 686
rect 819 682 820 686
rect 814 681 820 682
rect 950 686 956 687
rect 950 682 951 686
rect 955 682 956 686
rect 950 681 956 682
rect 1086 686 1092 687
rect 1086 682 1087 686
rect 1091 682 1092 686
rect 1086 681 1092 682
rect 1214 686 1220 687
rect 1214 682 1215 686
rect 1219 682 1220 686
rect 1214 681 1220 682
rect 1334 686 1340 687
rect 1334 682 1335 686
rect 1339 682 1340 686
rect 1334 681 1340 682
rect 1454 686 1460 687
rect 1454 682 1455 686
rect 1459 682 1460 686
rect 1454 681 1460 682
rect 1582 686 1588 687
rect 1582 682 1583 686
rect 1587 682 1588 686
rect 1582 681 1588 682
rect 1832 669 1834 697
rect 1870 696 1871 700
rect 1875 696 1876 700
rect 1870 695 1876 696
rect 3590 700 3596 701
rect 3590 696 3591 700
rect 3595 696 3596 700
rect 3590 695 3596 696
rect 110 668 116 669
rect 110 664 111 668
rect 115 664 116 668
rect 110 663 116 664
rect 1830 668 1836 669
rect 1830 664 1831 668
rect 1835 664 1836 668
rect 1872 667 1874 695
rect 1974 682 1980 683
rect 1974 678 1975 682
rect 1979 678 1980 682
rect 1974 677 1980 678
rect 2070 682 2076 683
rect 2070 678 2071 682
rect 2075 678 2076 682
rect 2070 677 2076 678
rect 2182 682 2188 683
rect 2182 678 2183 682
rect 2187 678 2188 682
rect 2182 677 2188 678
rect 2310 682 2316 683
rect 2310 678 2311 682
rect 2315 678 2316 682
rect 2310 677 2316 678
rect 2454 682 2460 683
rect 2454 678 2455 682
rect 2459 678 2460 682
rect 2454 677 2460 678
rect 2606 682 2612 683
rect 2606 678 2607 682
rect 2611 678 2612 682
rect 2606 677 2612 678
rect 2758 682 2764 683
rect 2758 678 2759 682
rect 2763 678 2764 682
rect 2758 677 2764 678
rect 2910 682 2916 683
rect 2910 678 2911 682
rect 2915 678 2916 682
rect 2910 677 2916 678
rect 3062 682 3068 683
rect 3062 678 3063 682
rect 3067 678 3068 682
rect 3062 677 3068 678
rect 3214 682 3220 683
rect 3214 678 3215 682
rect 3219 678 3220 682
rect 3214 677 3220 678
rect 3366 682 3372 683
rect 3366 678 3367 682
rect 3371 678 3372 682
rect 3366 677 3372 678
rect 3510 682 3516 683
rect 3510 678 3511 682
rect 3515 678 3516 682
rect 3510 677 3516 678
rect 1976 667 1978 677
rect 2072 667 2074 677
rect 2184 667 2186 677
rect 2312 667 2314 677
rect 2456 667 2458 677
rect 2608 667 2610 677
rect 2760 667 2762 677
rect 2912 667 2914 677
rect 3064 667 3066 677
rect 3216 667 3218 677
rect 3368 667 3370 677
rect 3512 667 3514 677
rect 3592 667 3594 695
rect 1830 663 1836 664
rect 1871 666 1875 667
rect 1871 661 1875 662
rect 1975 666 1979 667
rect 1975 661 1979 662
rect 2071 666 2075 667
rect 2071 661 2075 662
rect 2175 666 2179 667
rect 2175 661 2179 662
rect 2183 666 2187 667
rect 2183 661 2187 662
rect 2271 666 2275 667
rect 2271 661 2275 662
rect 2311 666 2315 667
rect 2311 661 2315 662
rect 2375 666 2379 667
rect 2375 661 2379 662
rect 2455 666 2459 667
rect 2455 661 2459 662
rect 2487 666 2491 667
rect 2487 661 2491 662
rect 2607 666 2611 667
rect 2607 661 2611 662
rect 2735 666 2739 667
rect 2735 661 2739 662
rect 2759 666 2763 667
rect 2759 661 2763 662
rect 2863 666 2867 667
rect 2863 661 2867 662
rect 2911 666 2915 667
rect 2911 661 2915 662
rect 2991 666 2995 667
rect 2991 661 2995 662
rect 3063 666 3067 667
rect 3063 661 3067 662
rect 3119 666 3123 667
rect 3119 661 3123 662
rect 3215 666 3219 667
rect 3215 661 3219 662
rect 3247 666 3251 667
rect 3247 661 3251 662
rect 3367 666 3371 667
rect 3367 661 3371 662
rect 3375 666 3379 667
rect 3375 661 3379 662
rect 3511 666 3515 667
rect 3511 661 3515 662
rect 3591 666 3595 667
rect 3591 661 3595 662
rect 110 651 116 652
rect 110 647 111 651
rect 115 647 116 651
rect 1830 651 1836 652
rect 110 646 116 647
rect 222 648 228 649
rect 112 619 114 646
rect 222 644 223 648
rect 227 644 228 648
rect 222 643 228 644
rect 310 648 316 649
rect 310 644 311 648
rect 315 644 316 648
rect 310 643 316 644
rect 414 648 420 649
rect 414 644 415 648
rect 419 644 420 648
rect 414 643 420 644
rect 534 648 540 649
rect 534 644 535 648
rect 539 644 540 648
rect 534 643 540 644
rect 670 648 676 649
rect 670 644 671 648
rect 675 644 676 648
rect 670 643 676 644
rect 806 648 812 649
rect 806 644 807 648
rect 811 644 812 648
rect 806 643 812 644
rect 942 648 948 649
rect 942 644 943 648
rect 947 644 948 648
rect 942 643 948 644
rect 1078 648 1084 649
rect 1078 644 1079 648
rect 1083 644 1084 648
rect 1078 643 1084 644
rect 1206 648 1212 649
rect 1206 644 1207 648
rect 1211 644 1212 648
rect 1206 643 1212 644
rect 1326 648 1332 649
rect 1326 644 1327 648
rect 1331 644 1332 648
rect 1326 643 1332 644
rect 1446 648 1452 649
rect 1446 644 1447 648
rect 1451 644 1452 648
rect 1446 643 1452 644
rect 1574 648 1580 649
rect 1574 644 1575 648
rect 1579 644 1580 648
rect 1830 647 1831 651
rect 1835 647 1836 651
rect 1830 646 1836 647
rect 1574 643 1580 644
rect 224 619 226 643
rect 312 619 314 643
rect 416 619 418 643
rect 536 619 538 643
rect 672 619 674 643
rect 808 619 810 643
rect 944 619 946 643
rect 1080 619 1082 643
rect 1208 619 1210 643
rect 1328 619 1330 643
rect 1448 619 1450 643
rect 1576 619 1578 643
rect 1832 619 1834 646
rect 1872 633 1874 661
rect 2176 651 2178 661
rect 2272 651 2274 661
rect 2376 651 2378 661
rect 2488 651 2490 661
rect 2608 651 2610 661
rect 2736 651 2738 661
rect 2864 651 2866 661
rect 2992 651 2994 661
rect 3120 651 3122 661
rect 3248 651 3250 661
rect 3376 651 3378 661
rect 3512 651 3514 661
rect 2174 650 2180 651
rect 2174 646 2175 650
rect 2179 646 2180 650
rect 2174 645 2180 646
rect 2270 650 2276 651
rect 2270 646 2271 650
rect 2275 646 2276 650
rect 2270 645 2276 646
rect 2374 650 2380 651
rect 2374 646 2375 650
rect 2379 646 2380 650
rect 2374 645 2380 646
rect 2486 650 2492 651
rect 2486 646 2487 650
rect 2491 646 2492 650
rect 2486 645 2492 646
rect 2606 650 2612 651
rect 2606 646 2607 650
rect 2611 646 2612 650
rect 2606 645 2612 646
rect 2734 650 2740 651
rect 2734 646 2735 650
rect 2739 646 2740 650
rect 2734 645 2740 646
rect 2862 650 2868 651
rect 2862 646 2863 650
rect 2867 646 2868 650
rect 2862 645 2868 646
rect 2990 650 2996 651
rect 2990 646 2991 650
rect 2995 646 2996 650
rect 2990 645 2996 646
rect 3118 650 3124 651
rect 3118 646 3119 650
rect 3123 646 3124 650
rect 3118 645 3124 646
rect 3246 650 3252 651
rect 3246 646 3247 650
rect 3251 646 3252 650
rect 3246 645 3252 646
rect 3374 650 3380 651
rect 3374 646 3375 650
rect 3379 646 3380 650
rect 3374 645 3380 646
rect 3510 650 3516 651
rect 3510 646 3511 650
rect 3515 646 3516 650
rect 3510 645 3516 646
rect 3592 633 3594 661
rect 1870 632 1876 633
rect 1870 628 1871 632
rect 1875 628 1876 632
rect 1870 627 1876 628
rect 3590 632 3596 633
rect 3590 628 3591 632
rect 3595 628 3596 632
rect 3590 627 3596 628
rect 111 618 115 619
rect 111 613 115 614
rect 223 618 227 619
rect 223 613 227 614
rect 311 618 315 619
rect 311 613 315 614
rect 415 618 419 619
rect 415 613 419 614
rect 447 618 451 619
rect 447 613 451 614
rect 527 618 531 619
rect 527 613 531 614
rect 535 618 539 619
rect 535 613 539 614
rect 607 618 611 619
rect 607 613 611 614
rect 671 618 675 619
rect 671 613 675 614
rect 687 618 691 619
rect 687 613 691 614
rect 775 618 779 619
rect 775 613 779 614
rect 807 618 811 619
rect 807 613 811 614
rect 871 618 875 619
rect 871 613 875 614
rect 943 618 947 619
rect 943 613 947 614
rect 959 618 963 619
rect 959 613 963 614
rect 1047 618 1051 619
rect 1047 613 1051 614
rect 1079 618 1083 619
rect 1079 613 1083 614
rect 1143 618 1147 619
rect 1143 613 1147 614
rect 1207 618 1211 619
rect 1207 613 1211 614
rect 1239 618 1243 619
rect 1239 613 1243 614
rect 1327 618 1331 619
rect 1327 613 1331 614
rect 1335 618 1339 619
rect 1335 613 1339 614
rect 1431 618 1435 619
rect 1431 613 1435 614
rect 1447 618 1451 619
rect 1447 613 1451 614
rect 1575 618 1579 619
rect 1575 613 1579 614
rect 1831 618 1835 619
rect 1831 613 1835 614
rect 1870 615 1876 616
rect 112 594 114 613
rect 448 597 450 613
rect 528 597 530 613
rect 608 597 610 613
rect 688 597 690 613
rect 776 597 778 613
rect 872 597 874 613
rect 960 597 962 613
rect 1048 597 1050 613
rect 1144 597 1146 613
rect 1240 597 1242 613
rect 1336 597 1338 613
rect 1432 597 1434 613
rect 446 596 452 597
rect 110 593 116 594
rect 110 589 111 593
rect 115 589 116 593
rect 446 592 447 596
rect 451 592 452 596
rect 446 591 452 592
rect 526 596 532 597
rect 526 592 527 596
rect 531 592 532 596
rect 526 591 532 592
rect 606 596 612 597
rect 606 592 607 596
rect 611 592 612 596
rect 606 591 612 592
rect 686 596 692 597
rect 686 592 687 596
rect 691 592 692 596
rect 686 591 692 592
rect 774 596 780 597
rect 774 592 775 596
rect 779 592 780 596
rect 774 591 780 592
rect 870 596 876 597
rect 870 592 871 596
rect 875 592 876 596
rect 870 591 876 592
rect 958 596 964 597
rect 958 592 959 596
rect 963 592 964 596
rect 958 591 964 592
rect 1046 596 1052 597
rect 1046 592 1047 596
rect 1051 592 1052 596
rect 1046 591 1052 592
rect 1142 596 1148 597
rect 1142 592 1143 596
rect 1147 592 1148 596
rect 1142 591 1148 592
rect 1238 596 1244 597
rect 1238 592 1239 596
rect 1243 592 1244 596
rect 1238 591 1244 592
rect 1334 596 1340 597
rect 1334 592 1335 596
rect 1339 592 1340 596
rect 1334 591 1340 592
rect 1430 596 1436 597
rect 1430 592 1431 596
rect 1435 592 1436 596
rect 1832 594 1834 613
rect 1870 611 1871 615
rect 1875 611 1876 615
rect 3590 615 3596 616
rect 1870 610 1876 611
rect 2166 612 2172 613
rect 1430 591 1436 592
rect 1830 593 1836 594
rect 110 588 116 589
rect 1830 589 1831 593
rect 1835 589 1836 593
rect 1872 591 1874 610
rect 2166 608 2167 612
rect 2171 608 2172 612
rect 2166 607 2172 608
rect 2262 612 2268 613
rect 2262 608 2263 612
rect 2267 608 2268 612
rect 2262 607 2268 608
rect 2366 612 2372 613
rect 2366 608 2367 612
rect 2371 608 2372 612
rect 2366 607 2372 608
rect 2478 612 2484 613
rect 2478 608 2479 612
rect 2483 608 2484 612
rect 2478 607 2484 608
rect 2598 612 2604 613
rect 2598 608 2599 612
rect 2603 608 2604 612
rect 2598 607 2604 608
rect 2726 612 2732 613
rect 2726 608 2727 612
rect 2731 608 2732 612
rect 2726 607 2732 608
rect 2854 612 2860 613
rect 2854 608 2855 612
rect 2859 608 2860 612
rect 2854 607 2860 608
rect 2982 612 2988 613
rect 2982 608 2983 612
rect 2987 608 2988 612
rect 2982 607 2988 608
rect 3110 612 3116 613
rect 3110 608 3111 612
rect 3115 608 3116 612
rect 3110 607 3116 608
rect 3238 612 3244 613
rect 3238 608 3239 612
rect 3243 608 3244 612
rect 3238 607 3244 608
rect 3366 612 3372 613
rect 3366 608 3367 612
rect 3371 608 3372 612
rect 3366 607 3372 608
rect 3502 612 3508 613
rect 3502 608 3503 612
rect 3507 608 3508 612
rect 3590 611 3591 615
rect 3595 611 3596 615
rect 3590 610 3596 611
rect 3502 607 3508 608
rect 2168 591 2170 607
rect 2264 591 2266 607
rect 2368 591 2370 607
rect 2480 591 2482 607
rect 2600 591 2602 607
rect 2728 591 2730 607
rect 2856 591 2858 607
rect 2984 591 2986 607
rect 3112 591 3114 607
rect 3240 591 3242 607
rect 3368 591 3370 607
rect 3504 591 3506 607
rect 3592 591 3594 610
rect 1830 588 1836 589
rect 1871 590 1875 591
rect 1871 585 1875 586
rect 2167 590 2171 591
rect 2167 585 2171 586
rect 2263 590 2267 591
rect 2263 585 2267 586
rect 2343 590 2347 591
rect 2343 585 2347 586
rect 2367 590 2371 591
rect 2367 585 2371 586
rect 2423 590 2427 591
rect 2423 585 2427 586
rect 2479 590 2483 591
rect 2479 585 2483 586
rect 2503 590 2507 591
rect 2503 585 2507 586
rect 2591 590 2595 591
rect 2591 585 2595 586
rect 2599 590 2603 591
rect 2599 585 2603 586
rect 2695 590 2699 591
rect 2695 585 2699 586
rect 2727 590 2731 591
rect 2727 585 2731 586
rect 2815 590 2819 591
rect 2815 585 2819 586
rect 2855 590 2859 591
rect 2855 585 2859 586
rect 2959 590 2963 591
rect 2959 585 2963 586
rect 2983 590 2987 591
rect 2983 585 2987 586
rect 3111 590 3115 591
rect 3111 585 3115 586
rect 3239 590 3243 591
rect 3239 585 3243 586
rect 3279 590 3283 591
rect 3279 585 3283 586
rect 3367 590 3371 591
rect 3367 585 3371 586
rect 3447 590 3451 591
rect 3447 585 3451 586
rect 3503 590 3507 591
rect 3503 585 3507 586
rect 3591 590 3595 591
rect 3591 585 3595 586
rect 110 576 116 577
rect 110 572 111 576
rect 115 572 116 576
rect 110 571 116 572
rect 1830 576 1836 577
rect 1830 572 1831 576
rect 1835 572 1836 576
rect 1830 571 1836 572
rect 112 531 114 571
rect 454 558 460 559
rect 454 554 455 558
rect 459 554 460 558
rect 454 553 460 554
rect 534 558 540 559
rect 534 554 535 558
rect 539 554 540 558
rect 534 553 540 554
rect 614 558 620 559
rect 614 554 615 558
rect 619 554 620 558
rect 614 553 620 554
rect 694 558 700 559
rect 694 554 695 558
rect 699 554 700 558
rect 694 553 700 554
rect 782 558 788 559
rect 782 554 783 558
rect 787 554 788 558
rect 782 553 788 554
rect 878 558 884 559
rect 878 554 879 558
rect 883 554 884 558
rect 878 553 884 554
rect 966 558 972 559
rect 966 554 967 558
rect 971 554 972 558
rect 966 553 972 554
rect 1054 558 1060 559
rect 1054 554 1055 558
rect 1059 554 1060 558
rect 1054 553 1060 554
rect 1150 558 1156 559
rect 1150 554 1151 558
rect 1155 554 1156 558
rect 1150 553 1156 554
rect 1246 558 1252 559
rect 1246 554 1247 558
rect 1251 554 1252 558
rect 1246 553 1252 554
rect 1342 558 1348 559
rect 1342 554 1343 558
rect 1347 554 1348 558
rect 1342 553 1348 554
rect 1438 558 1444 559
rect 1438 554 1439 558
rect 1443 554 1444 558
rect 1438 553 1444 554
rect 456 531 458 553
rect 536 531 538 553
rect 616 531 618 553
rect 696 531 698 553
rect 784 531 786 553
rect 880 531 882 553
rect 968 531 970 553
rect 1056 531 1058 553
rect 1152 531 1154 553
rect 1248 531 1250 553
rect 1344 531 1346 553
rect 1440 531 1442 553
rect 1832 531 1834 571
rect 1872 566 1874 585
rect 2264 569 2266 585
rect 2344 569 2346 585
rect 2424 569 2426 585
rect 2504 569 2506 585
rect 2592 569 2594 585
rect 2696 569 2698 585
rect 2816 569 2818 585
rect 2960 569 2962 585
rect 3112 569 3114 585
rect 3280 569 3282 585
rect 3448 569 3450 585
rect 2262 568 2268 569
rect 1870 565 1876 566
rect 1870 561 1871 565
rect 1875 561 1876 565
rect 2262 564 2263 568
rect 2267 564 2268 568
rect 2262 563 2268 564
rect 2342 568 2348 569
rect 2342 564 2343 568
rect 2347 564 2348 568
rect 2342 563 2348 564
rect 2422 568 2428 569
rect 2422 564 2423 568
rect 2427 564 2428 568
rect 2422 563 2428 564
rect 2502 568 2508 569
rect 2502 564 2503 568
rect 2507 564 2508 568
rect 2502 563 2508 564
rect 2590 568 2596 569
rect 2590 564 2591 568
rect 2595 564 2596 568
rect 2590 563 2596 564
rect 2694 568 2700 569
rect 2694 564 2695 568
rect 2699 564 2700 568
rect 2694 563 2700 564
rect 2814 568 2820 569
rect 2814 564 2815 568
rect 2819 564 2820 568
rect 2814 563 2820 564
rect 2958 568 2964 569
rect 2958 564 2959 568
rect 2963 564 2964 568
rect 2958 563 2964 564
rect 3110 568 3116 569
rect 3110 564 3111 568
rect 3115 564 3116 568
rect 3110 563 3116 564
rect 3278 568 3284 569
rect 3278 564 3279 568
rect 3283 564 3284 568
rect 3278 563 3284 564
rect 3446 568 3452 569
rect 3446 564 3447 568
rect 3451 564 3452 568
rect 3592 566 3594 585
rect 3446 563 3452 564
rect 3590 565 3596 566
rect 1870 560 1876 561
rect 3590 561 3591 565
rect 3595 561 3596 565
rect 3590 560 3596 561
rect 1870 548 1876 549
rect 1870 544 1871 548
rect 1875 544 1876 548
rect 1870 543 1876 544
rect 3590 548 3596 549
rect 3590 544 3591 548
rect 3595 544 3596 548
rect 3590 543 3596 544
rect 111 530 115 531
rect 111 525 115 526
rect 335 530 339 531
rect 335 525 339 526
rect 423 530 427 531
rect 423 525 427 526
rect 455 530 459 531
rect 455 525 459 526
rect 511 530 515 531
rect 511 525 515 526
rect 535 530 539 531
rect 535 525 539 526
rect 591 530 595 531
rect 591 525 595 526
rect 615 530 619 531
rect 615 525 619 526
rect 671 530 675 531
rect 671 525 675 526
rect 695 530 699 531
rect 695 525 699 526
rect 751 530 755 531
rect 751 525 755 526
rect 783 530 787 531
rect 783 525 787 526
rect 839 530 843 531
rect 839 525 843 526
rect 879 530 883 531
rect 879 525 883 526
rect 927 530 931 531
rect 927 525 931 526
rect 967 530 971 531
rect 967 525 971 526
rect 1015 530 1019 531
rect 1015 525 1019 526
rect 1055 530 1059 531
rect 1055 525 1059 526
rect 1103 530 1107 531
rect 1103 525 1107 526
rect 1151 530 1155 531
rect 1151 525 1155 526
rect 1191 530 1195 531
rect 1191 525 1195 526
rect 1247 530 1251 531
rect 1247 525 1251 526
rect 1279 530 1283 531
rect 1279 525 1283 526
rect 1343 530 1347 531
rect 1343 525 1347 526
rect 1439 530 1443 531
rect 1439 525 1443 526
rect 1831 530 1835 531
rect 1831 525 1835 526
rect 112 497 114 525
rect 336 515 338 525
rect 424 515 426 525
rect 512 515 514 525
rect 592 515 594 525
rect 672 515 674 525
rect 752 515 754 525
rect 840 515 842 525
rect 928 515 930 525
rect 1016 515 1018 525
rect 1104 515 1106 525
rect 1192 515 1194 525
rect 1280 515 1282 525
rect 334 514 340 515
rect 334 510 335 514
rect 339 510 340 514
rect 334 509 340 510
rect 422 514 428 515
rect 422 510 423 514
rect 427 510 428 514
rect 422 509 428 510
rect 510 514 516 515
rect 510 510 511 514
rect 515 510 516 514
rect 510 509 516 510
rect 590 514 596 515
rect 590 510 591 514
rect 595 510 596 514
rect 590 509 596 510
rect 670 514 676 515
rect 670 510 671 514
rect 675 510 676 514
rect 670 509 676 510
rect 750 514 756 515
rect 750 510 751 514
rect 755 510 756 514
rect 750 509 756 510
rect 838 514 844 515
rect 838 510 839 514
rect 843 510 844 514
rect 838 509 844 510
rect 926 514 932 515
rect 926 510 927 514
rect 931 510 932 514
rect 926 509 932 510
rect 1014 514 1020 515
rect 1014 510 1015 514
rect 1019 510 1020 514
rect 1014 509 1020 510
rect 1102 514 1108 515
rect 1102 510 1103 514
rect 1107 510 1108 514
rect 1102 509 1108 510
rect 1190 514 1196 515
rect 1190 510 1191 514
rect 1195 510 1196 514
rect 1190 509 1196 510
rect 1278 514 1284 515
rect 1278 510 1279 514
rect 1283 510 1284 514
rect 1278 509 1284 510
rect 1832 497 1834 525
rect 1872 507 1874 543
rect 2270 530 2276 531
rect 2270 526 2271 530
rect 2275 526 2276 530
rect 2270 525 2276 526
rect 2350 530 2356 531
rect 2350 526 2351 530
rect 2355 526 2356 530
rect 2350 525 2356 526
rect 2430 530 2436 531
rect 2430 526 2431 530
rect 2435 526 2436 530
rect 2430 525 2436 526
rect 2510 530 2516 531
rect 2510 526 2511 530
rect 2515 526 2516 530
rect 2510 525 2516 526
rect 2598 530 2604 531
rect 2598 526 2599 530
rect 2603 526 2604 530
rect 2598 525 2604 526
rect 2702 530 2708 531
rect 2702 526 2703 530
rect 2707 526 2708 530
rect 2702 525 2708 526
rect 2822 530 2828 531
rect 2822 526 2823 530
rect 2827 526 2828 530
rect 2822 525 2828 526
rect 2966 530 2972 531
rect 2966 526 2967 530
rect 2971 526 2972 530
rect 2966 525 2972 526
rect 3118 530 3124 531
rect 3118 526 3119 530
rect 3123 526 3124 530
rect 3118 525 3124 526
rect 3286 530 3292 531
rect 3286 526 3287 530
rect 3291 526 3292 530
rect 3286 525 3292 526
rect 3454 530 3460 531
rect 3454 526 3455 530
rect 3459 526 3460 530
rect 3454 525 3460 526
rect 2272 507 2274 525
rect 2352 507 2354 525
rect 2432 507 2434 525
rect 2512 507 2514 525
rect 2600 507 2602 525
rect 2704 507 2706 525
rect 2824 507 2826 525
rect 2968 507 2970 525
rect 3120 507 3122 525
rect 3288 507 3290 525
rect 3456 507 3458 525
rect 3592 507 3594 543
rect 1871 506 1875 507
rect 1871 501 1875 502
rect 2191 506 2195 507
rect 2191 501 2195 502
rect 2271 506 2275 507
rect 2271 501 2275 502
rect 2287 506 2291 507
rect 2287 501 2291 502
rect 2351 506 2355 507
rect 2351 501 2355 502
rect 2383 506 2387 507
rect 2383 501 2387 502
rect 2431 506 2435 507
rect 2431 501 2435 502
rect 2487 506 2491 507
rect 2487 501 2491 502
rect 2511 506 2515 507
rect 2511 501 2515 502
rect 2583 506 2587 507
rect 2583 501 2587 502
rect 2599 506 2603 507
rect 2599 501 2603 502
rect 2687 506 2691 507
rect 2687 501 2691 502
rect 2703 506 2707 507
rect 2703 501 2707 502
rect 2791 506 2795 507
rect 2791 501 2795 502
rect 2823 506 2827 507
rect 2823 501 2827 502
rect 2911 506 2915 507
rect 2911 501 2915 502
rect 2967 506 2971 507
rect 2967 501 2971 502
rect 3039 506 3043 507
rect 3039 501 3043 502
rect 3119 506 3123 507
rect 3119 501 3123 502
rect 3175 506 3179 507
rect 3175 501 3179 502
rect 3287 506 3291 507
rect 3287 501 3291 502
rect 3319 506 3323 507
rect 3319 501 3323 502
rect 3455 506 3459 507
rect 3455 501 3459 502
rect 3471 506 3475 507
rect 3471 501 3475 502
rect 3591 506 3595 507
rect 3591 501 3595 502
rect 110 496 116 497
rect 110 492 111 496
rect 115 492 116 496
rect 110 491 116 492
rect 1830 496 1836 497
rect 1830 492 1831 496
rect 1835 492 1836 496
rect 1830 491 1836 492
rect 110 479 116 480
rect 110 475 111 479
rect 115 475 116 479
rect 1830 479 1836 480
rect 110 474 116 475
rect 326 476 332 477
rect 112 447 114 474
rect 326 472 327 476
rect 331 472 332 476
rect 326 471 332 472
rect 414 476 420 477
rect 414 472 415 476
rect 419 472 420 476
rect 414 471 420 472
rect 502 476 508 477
rect 502 472 503 476
rect 507 472 508 476
rect 502 471 508 472
rect 582 476 588 477
rect 582 472 583 476
rect 587 472 588 476
rect 582 471 588 472
rect 662 476 668 477
rect 662 472 663 476
rect 667 472 668 476
rect 662 471 668 472
rect 742 476 748 477
rect 742 472 743 476
rect 747 472 748 476
rect 742 471 748 472
rect 830 476 836 477
rect 830 472 831 476
rect 835 472 836 476
rect 830 471 836 472
rect 918 476 924 477
rect 918 472 919 476
rect 923 472 924 476
rect 918 471 924 472
rect 1006 476 1012 477
rect 1006 472 1007 476
rect 1011 472 1012 476
rect 1006 471 1012 472
rect 1094 476 1100 477
rect 1094 472 1095 476
rect 1099 472 1100 476
rect 1094 471 1100 472
rect 1182 476 1188 477
rect 1182 472 1183 476
rect 1187 472 1188 476
rect 1182 471 1188 472
rect 1270 476 1276 477
rect 1270 472 1271 476
rect 1275 472 1276 476
rect 1830 475 1831 479
rect 1835 475 1836 479
rect 1830 474 1836 475
rect 1270 471 1276 472
rect 328 447 330 471
rect 416 447 418 471
rect 504 447 506 471
rect 584 447 586 471
rect 664 447 666 471
rect 744 447 746 471
rect 832 447 834 471
rect 920 447 922 471
rect 1008 447 1010 471
rect 1096 447 1098 471
rect 1184 447 1186 471
rect 1272 447 1274 471
rect 1832 447 1834 474
rect 1872 473 1874 501
rect 2192 491 2194 501
rect 2288 491 2290 501
rect 2384 491 2386 501
rect 2488 491 2490 501
rect 2584 491 2586 501
rect 2688 491 2690 501
rect 2792 491 2794 501
rect 2912 491 2914 501
rect 3040 491 3042 501
rect 3176 491 3178 501
rect 3320 491 3322 501
rect 3472 491 3474 501
rect 2190 490 2196 491
rect 2190 486 2191 490
rect 2195 486 2196 490
rect 2190 485 2196 486
rect 2286 490 2292 491
rect 2286 486 2287 490
rect 2291 486 2292 490
rect 2286 485 2292 486
rect 2382 490 2388 491
rect 2382 486 2383 490
rect 2387 486 2388 490
rect 2382 485 2388 486
rect 2486 490 2492 491
rect 2486 486 2487 490
rect 2491 486 2492 490
rect 2486 485 2492 486
rect 2582 490 2588 491
rect 2582 486 2583 490
rect 2587 486 2588 490
rect 2582 485 2588 486
rect 2686 490 2692 491
rect 2686 486 2687 490
rect 2691 486 2692 490
rect 2686 485 2692 486
rect 2790 490 2796 491
rect 2790 486 2791 490
rect 2795 486 2796 490
rect 2790 485 2796 486
rect 2910 490 2916 491
rect 2910 486 2911 490
rect 2915 486 2916 490
rect 2910 485 2916 486
rect 3038 490 3044 491
rect 3038 486 3039 490
rect 3043 486 3044 490
rect 3038 485 3044 486
rect 3174 490 3180 491
rect 3174 486 3175 490
rect 3179 486 3180 490
rect 3174 485 3180 486
rect 3318 490 3324 491
rect 3318 486 3319 490
rect 3323 486 3324 490
rect 3318 485 3324 486
rect 3470 490 3476 491
rect 3470 486 3471 490
rect 3475 486 3476 490
rect 3470 485 3476 486
rect 3592 473 3594 501
rect 1870 472 1876 473
rect 1870 468 1871 472
rect 1875 468 1876 472
rect 1870 467 1876 468
rect 3590 472 3596 473
rect 3590 468 3591 472
rect 3595 468 3596 472
rect 3590 467 3596 468
rect 1870 455 1876 456
rect 1870 451 1871 455
rect 1875 451 1876 455
rect 3590 455 3596 456
rect 1870 450 1876 451
rect 2182 452 2188 453
rect 111 446 115 447
rect 111 441 115 442
rect 223 446 227 447
rect 223 441 227 442
rect 327 446 331 447
rect 327 441 331 442
rect 335 446 339 447
rect 335 441 339 442
rect 415 446 419 447
rect 415 441 419 442
rect 447 446 451 447
rect 447 441 451 442
rect 503 446 507 447
rect 503 441 507 442
rect 559 446 563 447
rect 559 441 563 442
rect 583 446 587 447
rect 583 441 587 442
rect 663 446 667 447
rect 663 441 667 442
rect 743 446 747 447
rect 743 441 747 442
rect 759 446 763 447
rect 759 441 763 442
rect 831 446 835 447
rect 831 441 835 442
rect 847 446 851 447
rect 847 441 851 442
rect 919 446 923 447
rect 919 441 923 442
rect 935 446 939 447
rect 935 441 939 442
rect 1007 446 1011 447
rect 1007 441 1011 442
rect 1023 446 1027 447
rect 1023 441 1027 442
rect 1095 446 1099 447
rect 1095 441 1099 442
rect 1111 446 1115 447
rect 1111 441 1115 442
rect 1183 446 1187 447
rect 1183 441 1187 442
rect 1199 446 1203 447
rect 1199 441 1203 442
rect 1271 446 1275 447
rect 1271 441 1275 442
rect 1295 446 1299 447
rect 1295 441 1299 442
rect 1831 446 1835 447
rect 1831 441 1835 442
rect 112 422 114 441
rect 224 425 226 441
rect 336 425 338 441
rect 448 425 450 441
rect 560 425 562 441
rect 664 425 666 441
rect 760 425 762 441
rect 848 425 850 441
rect 936 425 938 441
rect 1024 425 1026 441
rect 1112 425 1114 441
rect 1200 425 1202 441
rect 1296 425 1298 441
rect 222 424 228 425
rect 110 421 116 422
rect 110 417 111 421
rect 115 417 116 421
rect 222 420 223 424
rect 227 420 228 424
rect 222 419 228 420
rect 334 424 340 425
rect 334 420 335 424
rect 339 420 340 424
rect 334 419 340 420
rect 446 424 452 425
rect 446 420 447 424
rect 451 420 452 424
rect 446 419 452 420
rect 558 424 564 425
rect 558 420 559 424
rect 563 420 564 424
rect 558 419 564 420
rect 662 424 668 425
rect 662 420 663 424
rect 667 420 668 424
rect 662 419 668 420
rect 758 424 764 425
rect 758 420 759 424
rect 763 420 764 424
rect 758 419 764 420
rect 846 424 852 425
rect 846 420 847 424
rect 851 420 852 424
rect 846 419 852 420
rect 934 424 940 425
rect 934 420 935 424
rect 939 420 940 424
rect 934 419 940 420
rect 1022 424 1028 425
rect 1022 420 1023 424
rect 1027 420 1028 424
rect 1022 419 1028 420
rect 1110 424 1116 425
rect 1110 420 1111 424
rect 1115 420 1116 424
rect 1110 419 1116 420
rect 1198 424 1204 425
rect 1198 420 1199 424
rect 1203 420 1204 424
rect 1198 419 1204 420
rect 1294 424 1300 425
rect 1294 420 1295 424
rect 1299 420 1300 424
rect 1832 422 1834 441
rect 1872 427 1874 450
rect 2182 448 2183 452
rect 2187 448 2188 452
rect 2182 447 2188 448
rect 2278 452 2284 453
rect 2278 448 2279 452
rect 2283 448 2284 452
rect 2278 447 2284 448
rect 2374 452 2380 453
rect 2374 448 2375 452
rect 2379 448 2380 452
rect 2374 447 2380 448
rect 2478 452 2484 453
rect 2478 448 2479 452
rect 2483 448 2484 452
rect 2478 447 2484 448
rect 2574 452 2580 453
rect 2574 448 2575 452
rect 2579 448 2580 452
rect 2574 447 2580 448
rect 2678 452 2684 453
rect 2678 448 2679 452
rect 2683 448 2684 452
rect 2678 447 2684 448
rect 2782 452 2788 453
rect 2782 448 2783 452
rect 2787 448 2788 452
rect 2782 447 2788 448
rect 2902 452 2908 453
rect 2902 448 2903 452
rect 2907 448 2908 452
rect 2902 447 2908 448
rect 3030 452 3036 453
rect 3030 448 3031 452
rect 3035 448 3036 452
rect 3030 447 3036 448
rect 3166 452 3172 453
rect 3166 448 3167 452
rect 3171 448 3172 452
rect 3166 447 3172 448
rect 3310 452 3316 453
rect 3310 448 3311 452
rect 3315 448 3316 452
rect 3310 447 3316 448
rect 3462 452 3468 453
rect 3462 448 3463 452
rect 3467 448 3468 452
rect 3590 451 3591 455
rect 3595 451 3596 455
rect 3590 450 3596 451
rect 3462 447 3468 448
rect 2184 427 2186 447
rect 2280 427 2282 447
rect 2376 427 2378 447
rect 2480 427 2482 447
rect 2576 427 2578 447
rect 2680 427 2682 447
rect 2784 427 2786 447
rect 2904 427 2906 447
rect 3032 427 3034 447
rect 3168 427 3170 447
rect 3312 427 3314 447
rect 3464 427 3466 447
rect 3592 427 3594 450
rect 1871 426 1875 427
rect 1294 419 1300 420
rect 1830 421 1836 422
rect 1871 421 1875 422
rect 1975 426 1979 427
rect 1975 421 1979 422
rect 2063 426 2067 427
rect 2063 421 2067 422
rect 2159 426 2163 427
rect 2159 421 2163 422
rect 2183 426 2187 427
rect 2183 421 2187 422
rect 2255 426 2259 427
rect 2255 421 2259 422
rect 2279 426 2283 427
rect 2279 421 2283 422
rect 2359 426 2363 427
rect 2359 421 2363 422
rect 2375 426 2379 427
rect 2375 421 2379 422
rect 2471 426 2475 427
rect 2471 421 2475 422
rect 2479 426 2483 427
rect 2479 421 2483 422
rect 2575 426 2579 427
rect 2575 421 2579 422
rect 2607 426 2611 427
rect 2607 421 2611 422
rect 2679 426 2683 427
rect 2679 421 2683 422
rect 2759 426 2763 427
rect 2759 421 2763 422
rect 2783 426 2787 427
rect 2783 421 2787 422
rect 2903 426 2907 427
rect 2903 421 2907 422
rect 2927 426 2931 427
rect 2927 421 2931 422
rect 3031 426 3035 427
rect 3031 421 3035 422
rect 3111 426 3115 427
rect 3111 421 3115 422
rect 3167 426 3171 427
rect 3167 421 3171 422
rect 3303 426 3307 427
rect 3303 421 3307 422
rect 3311 426 3315 427
rect 3311 421 3315 422
rect 3463 426 3467 427
rect 3463 421 3467 422
rect 3495 426 3499 427
rect 3495 421 3499 422
rect 3591 426 3595 427
rect 3591 421 3595 422
rect 110 416 116 417
rect 1830 417 1831 421
rect 1835 417 1836 421
rect 1830 416 1836 417
rect 110 404 116 405
rect 110 400 111 404
rect 115 400 116 404
rect 110 399 116 400
rect 1830 404 1836 405
rect 1830 400 1831 404
rect 1835 400 1836 404
rect 1872 402 1874 421
rect 1976 405 1978 421
rect 2064 405 2066 421
rect 2160 405 2162 421
rect 2256 405 2258 421
rect 2360 405 2362 421
rect 2472 405 2474 421
rect 2608 405 2610 421
rect 2760 405 2762 421
rect 2928 405 2930 421
rect 3112 405 3114 421
rect 3304 405 3306 421
rect 3496 405 3498 421
rect 1974 404 1980 405
rect 1830 399 1836 400
rect 1870 401 1876 402
rect 112 359 114 399
rect 230 386 236 387
rect 230 382 231 386
rect 235 382 236 386
rect 230 381 236 382
rect 342 386 348 387
rect 342 382 343 386
rect 347 382 348 386
rect 342 381 348 382
rect 454 386 460 387
rect 454 382 455 386
rect 459 382 460 386
rect 454 381 460 382
rect 566 386 572 387
rect 566 382 567 386
rect 571 382 572 386
rect 566 381 572 382
rect 670 386 676 387
rect 670 382 671 386
rect 675 382 676 386
rect 670 381 676 382
rect 766 386 772 387
rect 766 382 767 386
rect 771 382 772 386
rect 766 381 772 382
rect 854 386 860 387
rect 854 382 855 386
rect 859 382 860 386
rect 854 381 860 382
rect 942 386 948 387
rect 942 382 943 386
rect 947 382 948 386
rect 942 381 948 382
rect 1030 386 1036 387
rect 1030 382 1031 386
rect 1035 382 1036 386
rect 1030 381 1036 382
rect 1118 386 1124 387
rect 1118 382 1119 386
rect 1123 382 1124 386
rect 1118 381 1124 382
rect 1206 386 1212 387
rect 1206 382 1207 386
rect 1211 382 1212 386
rect 1206 381 1212 382
rect 1302 386 1308 387
rect 1302 382 1303 386
rect 1307 382 1308 386
rect 1302 381 1308 382
rect 232 359 234 381
rect 344 359 346 381
rect 456 359 458 381
rect 568 359 570 381
rect 672 359 674 381
rect 768 359 770 381
rect 856 359 858 381
rect 944 359 946 381
rect 1032 359 1034 381
rect 1120 359 1122 381
rect 1208 359 1210 381
rect 1304 359 1306 381
rect 1832 359 1834 399
rect 1870 397 1871 401
rect 1875 397 1876 401
rect 1974 400 1975 404
rect 1979 400 1980 404
rect 1974 399 1980 400
rect 2062 404 2068 405
rect 2062 400 2063 404
rect 2067 400 2068 404
rect 2062 399 2068 400
rect 2158 404 2164 405
rect 2158 400 2159 404
rect 2163 400 2164 404
rect 2158 399 2164 400
rect 2254 404 2260 405
rect 2254 400 2255 404
rect 2259 400 2260 404
rect 2254 399 2260 400
rect 2358 404 2364 405
rect 2358 400 2359 404
rect 2363 400 2364 404
rect 2358 399 2364 400
rect 2470 404 2476 405
rect 2470 400 2471 404
rect 2475 400 2476 404
rect 2470 399 2476 400
rect 2606 404 2612 405
rect 2606 400 2607 404
rect 2611 400 2612 404
rect 2606 399 2612 400
rect 2758 404 2764 405
rect 2758 400 2759 404
rect 2763 400 2764 404
rect 2758 399 2764 400
rect 2926 404 2932 405
rect 2926 400 2927 404
rect 2931 400 2932 404
rect 2926 399 2932 400
rect 3110 404 3116 405
rect 3110 400 3111 404
rect 3115 400 3116 404
rect 3110 399 3116 400
rect 3302 404 3308 405
rect 3302 400 3303 404
rect 3307 400 3308 404
rect 3302 399 3308 400
rect 3494 404 3500 405
rect 3494 400 3495 404
rect 3499 400 3500 404
rect 3592 402 3594 421
rect 3494 399 3500 400
rect 3590 401 3596 402
rect 1870 396 1876 397
rect 3590 397 3591 401
rect 3595 397 3596 401
rect 3590 396 3596 397
rect 1870 384 1876 385
rect 1870 380 1871 384
rect 1875 380 1876 384
rect 1870 379 1876 380
rect 3590 384 3596 385
rect 3590 380 3591 384
rect 3595 380 3596 384
rect 3590 379 3596 380
rect 111 358 115 359
rect 111 353 115 354
rect 143 358 147 359
rect 143 353 147 354
rect 231 358 235 359
rect 231 353 235 354
rect 263 358 267 359
rect 263 353 267 354
rect 343 358 347 359
rect 343 353 347 354
rect 399 358 403 359
rect 399 353 403 354
rect 455 358 459 359
rect 455 353 459 354
rect 535 358 539 359
rect 535 353 539 354
rect 567 358 571 359
rect 567 353 571 354
rect 671 358 675 359
rect 671 353 675 354
rect 767 358 771 359
rect 767 353 771 354
rect 791 358 795 359
rect 791 353 795 354
rect 855 358 859 359
rect 855 353 859 354
rect 911 358 915 359
rect 911 353 915 354
rect 943 358 947 359
rect 943 353 947 354
rect 1023 358 1027 359
rect 1023 353 1027 354
rect 1031 358 1035 359
rect 1031 353 1035 354
rect 1119 358 1123 359
rect 1119 353 1123 354
rect 1127 358 1131 359
rect 1127 353 1131 354
rect 1207 358 1211 359
rect 1207 353 1211 354
rect 1231 358 1235 359
rect 1231 353 1235 354
rect 1303 358 1307 359
rect 1303 353 1307 354
rect 1335 358 1339 359
rect 1335 353 1339 354
rect 1439 358 1443 359
rect 1439 353 1443 354
rect 1831 358 1835 359
rect 1831 353 1835 354
rect 112 325 114 353
rect 144 343 146 353
rect 264 343 266 353
rect 400 343 402 353
rect 536 343 538 353
rect 672 343 674 353
rect 792 343 794 353
rect 912 343 914 353
rect 1024 343 1026 353
rect 1128 343 1130 353
rect 1232 343 1234 353
rect 1336 343 1338 353
rect 1440 343 1442 353
rect 142 342 148 343
rect 142 338 143 342
rect 147 338 148 342
rect 142 337 148 338
rect 262 342 268 343
rect 262 338 263 342
rect 267 338 268 342
rect 262 337 268 338
rect 398 342 404 343
rect 398 338 399 342
rect 403 338 404 342
rect 398 337 404 338
rect 534 342 540 343
rect 534 338 535 342
rect 539 338 540 342
rect 534 337 540 338
rect 670 342 676 343
rect 670 338 671 342
rect 675 338 676 342
rect 670 337 676 338
rect 790 342 796 343
rect 790 338 791 342
rect 795 338 796 342
rect 790 337 796 338
rect 910 342 916 343
rect 910 338 911 342
rect 915 338 916 342
rect 910 337 916 338
rect 1022 342 1028 343
rect 1022 338 1023 342
rect 1027 338 1028 342
rect 1022 337 1028 338
rect 1126 342 1132 343
rect 1126 338 1127 342
rect 1131 338 1132 342
rect 1126 337 1132 338
rect 1230 342 1236 343
rect 1230 338 1231 342
rect 1235 338 1236 342
rect 1230 337 1236 338
rect 1334 342 1340 343
rect 1334 338 1335 342
rect 1339 338 1340 342
rect 1334 337 1340 338
rect 1438 342 1444 343
rect 1438 338 1439 342
rect 1443 338 1444 342
rect 1438 337 1444 338
rect 1832 325 1834 353
rect 1872 347 1874 379
rect 1982 366 1988 367
rect 1982 362 1983 366
rect 1987 362 1988 366
rect 1982 361 1988 362
rect 2070 366 2076 367
rect 2070 362 2071 366
rect 2075 362 2076 366
rect 2070 361 2076 362
rect 2166 366 2172 367
rect 2166 362 2167 366
rect 2171 362 2172 366
rect 2166 361 2172 362
rect 2262 366 2268 367
rect 2262 362 2263 366
rect 2267 362 2268 366
rect 2262 361 2268 362
rect 2366 366 2372 367
rect 2366 362 2367 366
rect 2371 362 2372 366
rect 2366 361 2372 362
rect 2478 366 2484 367
rect 2478 362 2479 366
rect 2483 362 2484 366
rect 2478 361 2484 362
rect 2614 366 2620 367
rect 2614 362 2615 366
rect 2619 362 2620 366
rect 2614 361 2620 362
rect 2766 366 2772 367
rect 2766 362 2767 366
rect 2771 362 2772 366
rect 2766 361 2772 362
rect 2934 366 2940 367
rect 2934 362 2935 366
rect 2939 362 2940 366
rect 2934 361 2940 362
rect 3118 366 3124 367
rect 3118 362 3119 366
rect 3123 362 3124 366
rect 3118 361 3124 362
rect 3310 366 3316 367
rect 3310 362 3311 366
rect 3315 362 3316 366
rect 3310 361 3316 362
rect 3502 366 3508 367
rect 3502 362 3503 366
rect 3507 362 3508 366
rect 3502 361 3508 362
rect 1984 347 1986 361
rect 2072 347 2074 361
rect 2168 347 2170 361
rect 2264 347 2266 361
rect 2368 347 2370 361
rect 2480 347 2482 361
rect 2616 347 2618 361
rect 2768 347 2770 361
rect 2936 347 2938 361
rect 3120 347 3122 361
rect 3312 347 3314 361
rect 3504 347 3506 361
rect 3592 347 3594 379
rect 1871 346 1875 347
rect 1871 341 1875 342
rect 1983 346 1987 347
rect 1983 341 1987 342
rect 2071 346 2075 347
rect 2071 341 2075 342
rect 2167 346 2171 347
rect 2167 341 2171 342
rect 2215 346 2219 347
rect 2215 341 2219 342
rect 2263 346 2267 347
rect 2263 341 2267 342
rect 2295 346 2299 347
rect 2295 341 2299 342
rect 2367 346 2371 347
rect 2367 341 2371 342
rect 2383 346 2387 347
rect 2383 341 2387 342
rect 2479 346 2483 347
rect 2479 341 2483 342
rect 2591 346 2595 347
rect 2591 341 2595 342
rect 2615 346 2619 347
rect 2615 341 2619 342
rect 2719 346 2723 347
rect 2719 341 2723 342
rect 2767 346 2771 347
rect 2767 341 2771 342
rect 2847 346 2851 347
rect 2847 341 2851 342
rect 2935 346 2939 347
rect 2935 341 2939 342
rect 2983 346 2987 347
rect 2983 341 2987 342
rect 3119 346 3123 347
rect 3119 341 3123 342
rect 3255 346 3259 347
rect 3255 341 3259 342
rect 3311 346 3315 347
rect 3311 341 3315 342
rect 3391 346 3395 347
rect 3391 341 3395 342
rect 3503 346 3507 347
rect 3503 341 3507 342
rect 3511 346 3515 347
rect 3511 341 3515 342
rect 3591 346 3595 347
rect 3591 341 3595 342
rect 110 324 116 325
rect 110 320 111 324
rect 115 320 116 324
rect 110 319 116 320
rect 1830 324 1836 325
rect 1830 320 1831 324
rect 1835 320 1836 324
rect 1830 319 1836 320
rect 1872 313 1874 341
rect 2216 331 2218 341
rect 2296 331 2298 341
rect 2384 331 2386 341
rect 2480 331 2482 341
rect 2592 331 2594 341
rect 2720 331 2722 341
rect 2848 331 2850 341
rect 2984 331 2986 341
rect 3120 331 3122 341
rect 3256 331 3258 341
rect 3392 331 3394 341
rect 3512 331 3514 341
rect 2214 330 2220 331
rect 2214 326 2215 330
rect 2219 326 2220 330
rect 2214 325 2220 326
rect 2294 330 2300 331
rect 2294 326 2295 330
rect 2299 326 2300 330
rect 2294 325 2300 326
rect 2382 330 2388 331
rect 2382 326 2383 330
rect 2387 326 2388 330
rect 2382 325 2388 326
rect 2478 330 2484 331
rect 2478 326 2479 330
rect 2483 326 2484 330
rect 2478 325 2484 326
rect 2590 330 2596 331
rect 2590 326 2591 330
rect 2595 326 2596 330
rect 2590 325 2596 326
rect 2718 330 2724 331
rect 2718 326 2719 330
rect 2723 326 2724 330
rect 2718 325 2724 326
rect 2846 330 2852 331
rect 2846 326 2847 330
rect 2851 326 2852 330
rect 2846 325 2852 326
rect 2982 330 2988 331
rect 2982 326 2983 330
rect 2987 326 2988 330
rect 2982 325 2988 326
rect 3118 330 3124 331
rect 3118 326 3119 330
rect 3123 326 3124 330
rect 3118 325 3124 326
rect 3254 330 3260 331
rect 3254 326 3255 330
rect 3259 326 3260 330
rect 3254 325 3260 326
rect 3390 330 3396 331
rect 3390 326 3391 330
rect 3395 326 3396 330
rect 3390 325 3396 326
rect 3510 330 3516 331
rect 3510 326 3511 330
rect 3515 326 3516 330
rect 3510 325 3516 326
rect 3592 313 3594 341
rect 1870 312 1876 313
rect 1870 308 1871 312
rect 1875 308 1876 312
rect 110 307 116 308
rect 110 303 111 307
rect 115 303 116 307
rect 1830 307 1836 308
rect 1870 307 1876 308
rect 3590 312 3596 313
rect 3590 308 3591 312
rect 3595 308 3596 312
rect 3590 307 3596 308
rect 110 302 116 303
rect 134 304 140 305
rect 112 275 114 302
rect 134 300 135 304
rect 139 300 140 304
rect 134 299 140 300
rect 254 304 260 305
rect 254 300 255 304
rect 259 300 260 304
rect 254 299 260 300
rect 390 304 396 305
rect 390 300 391 304
rect 395 300 396 304
rect 390 299 396 300
rect 526 304 532 305
rect 526 300 527 304
rect 531 300 532 304
rect 526 299 532 300
rect 662 304 668 305
rect 662 300 663 304
rect 667 300 668 304
rect 662 299 668 300
rect 782 304 788 305
rect 782 300 783 304
rect 787 300 788 304
rect 782 299 788 300
rect 902 304 908 305
rect 902 300 903 304
rect 907 300 908 304
rect 902 299 908 300
rect 1014 304 1020 305
rect 1014 300 1015 304
rect 1019 300 1020 304
rect 1014 299 1020 300
rect 1118 304 1124 305
rect 1118 300 1119 304
rect 1123 300 1124 304
rect 1118 299 1124 300
rect 1222 304 1228 305
rect 1222 300 1223 304
rect 1227 300 1228 304
rect 1222 299 1228 300
rect 1326 304 1332 305
rect 1326 300 1327 304
rect 1331 300 1332 304
rect 1326 299 1332 300
rect 1430 304 1436 305
rect 1430 300 1431 304
rect 1435 300 1436 304
rect 1830 303 1831 307
rect 1835 303 1836 307
rect 1830 302 1836 303
rect 1430 299 1436 300
rect 136 275 138 299
rect 256 275 258 299
rect 392 275 394 299
rect 528 275 530 299
rect 664 275 666 299
rect 784 275 786 299
rect 904 275 906 299
rect 1016 275 1018 299
rect 1120 275 1122 299
rect 1224 275 1226 299
rect 1328 275 1330 299
rect 1432 275 1434 299
rect 1832 275 1834 302
rect 1870 295 1876 296
rect 1870 291 1871 295
rect 1875 291 1876 295
rect 3590 295 3596 296
rect 1870 290 1876 291
rect 2206 292 2212 293
rect 111 274 115 275
rect 111 269 115 270
rect 135 274 139 275
rect 135 269 139 270
rect 247 274 251 275
rect 247 269 251 270
rect 255 274 259 275
rect 255 269 259 270
rect 391 274 395 275
rect 391 269 395 270
rect 527 274 531 275
rect 527 269 531 270
rect 543 274 547 275
rect 543 269 547 270
rect 663 274 667 275
rect 663 269 667 270
rect 695 274 699 275
rect 695 269 699 270
rect 783 274 787 275
rect 783 269 787 270
rect 847 274 851 275
rect 847 269 851 270
rect 903 274 907 275
rect 903 269 907 270
rect 991 274 995 275
rect 991 269 995 270
rect 1015 274 1019 275
rect 1015 269 1019 270
rect 1119 274 1123 275
rect 1119 269 1123 270
rect 1223 274 1227 275
rect 1223 269 1227 270
rect 1239 274 1243 275
rect 1239 269 1243 270
rect 1327 274 1331 275
rect 1327 269 1331 270
rect 1359 274 1363 275
rect 1359 269 1363 270
rect 1431 274 1435 275
rect 1431 269 1435 270
rect 1479 274 1483 275
rect 1479 269 1483 270
rect 1599 274 1603 275
rect 1599 269 1603 270
rect 1831 274 1835 275
rect 1831 269 1835 270
rect 112 250 114 269
rect 136 253 138 269
rect 248 253 250 269
rect 392 253 394 269
rect 544 253 546 269
rect 696 253 698 269
rect 848 253 850 269
rect 992 253 994 269
rect 1120 253 1122 269
rect 1240 253 1242 269
rect 1360 253 1362 269
rect 1480 253 1482 269
rect 1600 253 1602 269
rect 134 252 140 253
rect 110 249 116 250
rect 110 245 111 249
rect 115 245 116 249
rect 134 248 135 252
rect 139 248 140 252
rect 134 247 140 248
rect 246 252 252 253
rect 246 248 247 252
rect 251 248 252 252
rect 246 247 252 248
rect 390 252 396 253
rect 390 248 391 252
rect 395 248 396 252
rect 390 247 396 248
rect 542 252 548 253
rect 542 248 543 252
rect 547 248 548 252
rect 542 247 548 248
rect 694 252 700 253
rect 694 248 695 252
rect 699 248 700 252
rect 694 247 700 248
rect 846 252 852 253
rect 846 248 847 252
rect 851 248 852 252
rect 846 247 852 248
rect 990 252 996 253
rect 990 248 991 252
rect 995 248 996 252
rect 990 247 996 248
rect 1118 252 1124 253
rect 1118 248 1119 252
rect 1123 248 1124 252
rect 1118 247 1124 248
rect 1238 252 1244 253
rect 1238 248 1239 252
rect 1243 248 1244 252
rect 1238 247 1244 248
rect 1358 252 1364 253
rect 1358 248 1359 252
rect 1363 248 1364 252
rect 1358 247 1364 248
rect 1478 252 1484 253
rect 1478 248 1479 252
rect 1483 248 1484 252
rect 1478 247 1484 248
rect 1598 252 1604 253
rect 1598 248 1599 252
rect 1603 248 1604 252
rect 1832 250 1834 269
rect 1872 267 1874 290
rect 2206 288 2207 292
rect 2211 288 2212 292
rect 2206 287 2212 288
rect 2286 292 2292 293
rect 2286 288 2287 292
rect 2291 288 2292 292
rect 2286 287 2292 288
rect 2374 292 2380 293
rect 2374 288 2375 292
rect 2379 288 2380 292
rect 2374 287 2380 288
rect 2470 292 2476 293
rect 2470 288 2471 292
rect 2475 288 2476 292
rect 2470 287 2476 288
rect 2582 292 2588 293
rect 2582 288 2583 292
rect 2587 288 2588 292
rect 2582 287 2588 288
rect 2710 292 2716 293
rect 2710 288 2711 292
rect 2715 288 2716 292
rect 2710 287 2716 288
rect 2838 292 2844 293
rect 2838 288 2839 292
rect 2843 288 2844 292
rect 2838 287 2844 288
rect 2974 292 2980 293
rect 2974 288 2975 292
rect 2979 288 2980 292
rect 2974 287 2980 288
rect 3110 292 3116 293
rect 3110 288 3111 292
rect 3115 288 3116 292
rect 3110 287 3116 288
rect 3246 292 3252 293
rect 3246 288 3247 292
rect 3251 288 3252 292
rect 3246 287 3252 288
rect 3382 292 3388 293
rect 3382 288 3383 292
rect 3387 288 3388 292
rect 3382 287 3388 288
rect 3502 292 3508 293
rect 3502 288 3503 292
rect 3507 288 3508 292
rect 3590 291 3591 295
rect 3595 291 3596 295
rect 3590 290 3596 291
rect 3502 287 3508 288
rect 2208 267 2210 287
rect 2288 267 2290 287
rect 2376 267 2378 287
rect 2472 267 2474 287
rect 2584 267 2586 287
rect 2712 267 2714 287
rect 2840 267 2842 287
rect 2976 267 2978 287
rect 3112 267 3114 287
rect 3248 267 3250 287
rect 3384 267 3386 287
rect 3504 267 3506 287
rect 3592 267 3594 290
rect 1871 266 1875 267
rect 1871 261 1875 262
rect 1991 266 1995 267
rect 1991 261 1995 262
rect 2119 266 2123 267
rect 2119 261 2123 262
rect 2207 266 2211 267
rect 2207 261 2211 262
rect 2255 266 2259 267
rect 2255 261 2259 262
rect 2287 266 2291 267
rect 2287 261 2291 262
rect 2375 266 2379 267
rect 2375 261 2379 262
rect 2391 266 2395 267
rect 2391 261 2395 262
rect 2471 266 2475 267
rect 2471 261 2475 262
rect 2535 266 2539 267
rect 2535 261 2539 262
rect 2583 266 2587 267
rect 2583 261 2587 262
rect 2679 266 2683 267
rect 2679 261 2683 262
rect 2711 266 2715 267
rect 2711 261 2715 262
rect 2815 266 2819 267
rect 2815 261 2819 262
rect 2839 266 2843 267
rect 2839 261 2843 262
rect 2951 266 2955 267
rect 2951 261 2955 262
rect 2975 266 2979 267
rect 2975 261 2979 262
rect 3095 266 3099 267
rect 3095 261 3099 262
rect 3111 266 3115 267
rect 3111 261 3115 262
rect 3239 266 3243 267
rect 3239 261 3243 262
rect 3247 266 3251 267
rect 3247 261 3251 262
rect 3383 266 3387 267
rect 3383 261 3387 262
rect 3503 266 3507 267
rect 3503 261 3507 262
rect 3591 266 3595 267
rect 3591 261 3595 262
rect 1598 247 1604 248
rect 1830 249 1836 250
rect 110 244 116 245
rect 1830 245 1831 249
rect 1835 245 1836 249
rect 1830 244 1836 245
rect 1872 242 1874 261
rect 1992 245 1994 261
rect 2120 245 2122 261
rect 2256 245 2258 261
rect 2392 245 2394 261
rect 2536 245 2538 261
rect 2680 245 2682 261
rect 2816 245 2818 261
rect 2952 245 2954 261
rect 3096 245 3098 261
rect 3240 245 3242 261
rect 3384 245 3386 261
rect 3504 245 3506 261
rect 1990 244 1996 245
rect 1870 241 1876 242
rect 1870 237 1871 241
rect 1875 237 1876 241
rect 1990 240 1991 244
rect 1995 240 1996 244
rect 1990 239 1996 240
rect 2118 244 2124 245
rect 2118 240 2119 244
rect 2123 240 2124 244
rect 2118 239 2124 240
rect 2254 244 2260 245
rect 2254 240 2255 244
rect 2259 240 2260 244
rect 2254 239 2260 240
rect 2390 244 2396 245
rect 2390 240 2391 244
rect 2395 240 2396 244
rect 2390 239 2396 240
rect 2534 244 2540 245
rect 2534 240 2535 244
rect 2539 240 2540 244
rect 2534 239 2540 240
rect 2678 244 2684 245
rect 2678 240 2679 244
rect 2683 240 2684 244
rect 2678 239 2684 240
rect 2814 244 2820 245
rect 2814 240 2815 244
rect 2819 240 2820 244
rect 2814 239 2820 240
rect 2950 244 2956 245
rect 2950 240 2951 244
rect 2955 240 2956 244
rect 2950 239 2956 240
rect 3094 244 3100 245
rect 3094 240 3095 244
rect 3099 240 3100 244
rect 3094 239 3100 240
rect 3238 244 3244 245
rect 3238 240 3239 244
rect 3243 240 3244 244
rect 3238 239 3244 240
rect 3382 244 3388 245
rect 3382 240 3383 244
rect 3387 240 3388 244
rect 3382 239 3388 240
rect 3502 244 3508 245
rect 3502 240 3503 244
rect 3507 240 3508 244
rect 3592 242 3594 261
rect 3502 239 3508 240
rect 3590 241 3596 242
rect 1870 236 1876 237
rect 3590 237 3591 241
rect 3595 237 3596 241
rect 3590 236 3596 237
rect 110 232 116 233
rect 110 228 111 232
rect 115 228 116 232
rect 110 227 116 228
rect 1830 232 1836 233
rect 1830 228 1831 232
rect 1835 228 1836 232
rect 1830 227 1836 228
rect 112 163 114 227
rect 142 214 148 215
rect 142 210 143 214
rect 147 210 148 214
rect 142 209 148 210
rect 254 214 260 215
rect 254 210 255 214
rect 259 210 260 214
rect 254 209 260 210
rect 398 214 404 215
rect 398 210 399 214
rect 403 210 404 214
rect 398 209 404 210
rect 550 214 556 215
rect 550 210 551 214
rect 555 210 556 214
rect 550 209 556 210
rect 702 214 708 215
rect 702 210 703 214
rect 707 210 708 214
rect 702 209 708 210
rect 854 214 860 215
rect 854 210 855 214
rect 859 210 860 214
rect 854 209 860 210
rect 998 214 1004 215
rect 998 210 999 214
rect 1003 210 1004 214
rect 998 209 1004 210
rect 1126 214 1132 215
rect 1126 210 1127 214
rect 1131 210 1132 214
rect 1126 209 1132 210
rect 1246 214 1252 215
rect 1246 210 1247 214
rect 1251 210 1252 214
rect 1246 209 1252 210
rect 1366 214 1372 215
rect 1366 210 1367 214
rect 1371 210 1372 214
rect 1366 209 1372 210
rect 1486 214 1492 215
rect 1486 210 1487 214
rect 1491 210 1492 214
rect 1486 209 1492 210
rect 1606 214 1612 215
rect 1606 210 1607 214
rect 1611 210 1612 214
rect 1606 209 1612 210
rect 144 163 146 209
rect 256 163 258 209
rect 400 163 402 209
rect 552 163 554 209
rect 704 163 706 209
rect 856 163 858 209
rect 1000 163 1002 209
rect 1128 163 1130 209
rect 1248 163 1250 209
rect 1368 163 1370 209
rect 1488 163 1490 209
rect 1608 163 1610 209
rect 1832 163 1834 227
rect 1870 224 1876 225
rect 1870 220 1871 224
rect 1875 220 1876 224
rect 1870 219 1876 220
rect 3590 224 3596 225
rect 3590 220 3591 224
rect 3595 220 3596 224
rect 3590 219 3596 220
rect 1872 179 1874 219
rect 1998 206 2004 207
rect 1998 202 1999 206
rect 2003 202 2004 206
rect 1998 201 2004 202
rect 2126 206 2132 207
rect 2126 202 2127 206
rect 2131 202 2132 206
rect 2126 201 2132 202
rect 2262 206 2268 207
rect 2262 202 2263 206
rect 2267 202 2268 206
rect 2262 201 2268 202
rect 2398 206 2404 207
rect 2398 202 2399 206
rect 2403 202 2404 206
rect 2398 201 2404 202
rect 2542 206 2548 207
rect 2542 202 2543 206
rect 2547 202 2548 206
rect 2542 201 2548 202
rect 2686 206 2692 207
rect 2686 202 2687 206
rect 2691 202 2692 206
rect 2686 201 2692 202
rect 2822 206 2828 207
rect 2822 202 2823 206
rect 2827 202 2828 206
rect 2822 201 2828 202
rect 2958 206 2964 207
rect 2958 202 2959 206
rect 2963 202 2964 206
rect 2958 201 2964 202
rect 3102 206 3108 207
rect 3102 202 3103 206
rect 3107 202 3108 206
rect 3102 201 3108 202
rect 3246 206 3252 207
rect 3246 202 3247 206
rect 3251 202 3252 206
rect 3246 201 3252 202
rect 3390 206 3396 207
rect 3390 202 3391 206
rect 3395 202 3396 206
rect 3390 201 3396 202
rect 3510 206 3516 207
rect 3510 202 3511 206
rect 3515 202 3516 206
rect 3510 201 3516 202
rect 2000 179 2002 201
rect 2128 179 2130 201
rect 2264 179 2266 201
rect 2400 179 2402 201
rect 2544 179 2546 201
rect 2688 179 2690 201
rect 2824 179 2826 201
rect 2960 179 2962 201
rect 3104 179 3106 201
rect 3248 179 3250 201
rect 3392 179 3394 201
rect 3512 179 3514 201
rect 3592 179 3594 219
rect 1871 178 1875 179
rect 1871 173 1875 174
rect 1903 178 1907 179
rect 1903 173 1907 174
rect 1983 178 1987 179
rect 1983 173 1987 174
rect 1999 178 2003 179
rect 1999 173 2003 174
rect 2087 178 2091 179
rect 2087 173 2091 174
rect 2127 178 2131 179
rect 2127 173 2131 174
rect 2215 178 2219 179
rect 2215 173 2219 174
rect 2263 178 2267 179
rect 2263 173 2267 174
rect 2351 178 2355 179
rect 2351 173 2355 174
rect 2399 178 2403 179
rect 2399 173 2403 174
rect 2487 178 2491 179
rect 2487 173 2491 174
rect 2543 178 2547 179
rect 2543 173 2547 174
rect 2623 178 2627 179
rect 2623 173 2627 174
rect 2687 178 2691 179
rect 2687 173 2691 174
rect 2743 178 2747 179
rect 2743 173 2747 174
rect 2823 178 2827 179
rect 2823 173 2827 174
rect 2855 178 2859 179
rect 2855 173 2859 174
rect 2959 178 2963 179
rect 2959 173 2963 174
rect 3063 178 3067 179
rect 3063 173 3067 174
rect 3103 178 3107 179
rect 3103 173 3107 174
rect 3159 178 3163 179
rect 3159 173 3163 174
rect 3247 178 3251 179
rect 3247 173 3251 174
rect 3343 178 3347 179
rect 3343 173 3347 174
rect 3391 178 3395 179
rect 3391 173 3395 174
rect 3431 178 3435 179
rect 3431 173 3435 174
rect 3511 178 3515 179
rect 3511 173 3515 174
rect 3591 178 3595 179
rect 3591 173 3595 174
rect 111 162 115 163
rect 111 157 115 158
rect 143 162 147 163
rect 143 157 147 158
rect 223 162 227 163
rect 223 157 227 158
rect 255 162 259 163
rect 255 157 259 158
rect 303 162 307 163
rect 303 157 307 158
rect 383 162 387 163
rect 383 157 387 158
rect 399 162 403 163
rect 399 157 403 158
rect 463 162 467 163
rect 463 157 467 158
rect 543 162 547 163
rect 543 157 547 158
rect 551 162 555 163
rect 551 157 555 158
rect 623 162 627 163
rect 623 157 627 158
rect 703 162 707 163
rect 703 157 707 158
rect 783 162 787 163
rect 783 157 787 158
rect 855 162 859 163
rect 855 157 859 158
rect 863 162 867 163
rect 863 157 867 158
rect 943 162 947 163
rect 943 157 947 158
rect 999 162 1003 163
rect 999 157 1003 158
rect 1023 162 1027 163
rect 1023 157 1027 158
rect 1103 162 1107 163
rect 1103 157 1107 158
rect 1127 162 1131 163
rect 1127 157 1131 158
rect 1183 162 1187 163
rect 1183 157 1187 158
rect 1247 162 1251 163
rect 1247 157 1251 158
rect 1263 162 1267 163
rect 1263 157 1267 158
rect 1343 162 1347 163
rect 1343 157 1347 158
rect 1367 162 1371 163
rect 1367 157 1371 158
rect 1423 162 1427 163
rect 1423 157 1427 158
rect 1487 162 1491 163
rect 1487 157 1491 158
rect 1511 162 1515 163
rect 1511 157 1515 158
rect 1591 162 1595 163
rect 1591 157 1595 158
rect 1607 162 1611 163
rect 1607 157 1611 158
rect 1671 162 1675 163
rect 1671 157 1675 158
rect 1751 162 1755 163
rect 1751 157 1755 158
rect 1831 162 1835 163
rect 1831 157 1835 158
rect 112 129 114 157
rect 144 147 146 157
rect 224 147 226 157
rect 304 147 306 157
rect 384 147 386 157
rect 464 147 466 157
rect 544 147 546 157
rect 624 147 626 157
rect 704 147 706 157
rect 784 147 786 157
rect 864 147 866 157
rect 944 147 946 157
rect 1024 147 1026 157
rect 1104 147 1106 157
rect 1184 147 1186 157
rect 1264 147 1266 157
rect 1344 147 1346 157
rect 1424 147 1426 157
rect 1512 147 1514 157
rect 1592 147 1594 157
rect 1672 147 1674 157
rect 1752 147 1754 157
rect 142 146 148 147
rect 142 142 143 146
rect 147 142 148 146
rect 142 141 148 142
rect 222 146 228 147
rect 222 142 223 146
rect 227 142 228 146
rect 222 141 228 142
rect 302 146 308 147
rect 302 142 303 146
rect 307 142 308 146
rect 302 141 308 142
rect 382 146 388 147
rect 382 142 383 146
rect 387 142 388 146
rect 382 141 388 142
rect 462 146 468 147
rect 462 142 463 146
rect 467 142 468 146
rect 462 141 468 142
rect 542 146 548 147
rect 542 142 543 146
rect 547 142 548 146
rect 542 141 548 142
rect 622 146 628 147
rect 622 142 623 146
rect 627 142 628 146
rect 622 141 628 142
rect 702 146 708 147
rect 702 142 703 146
rect 707 142 708 146
rect 702 141 708 142
rect 782 146 788 147
rect 782 142 783 146
rect 787 142 788 146
rect 782 141 788 142
rect 862 146 868 147
rect 862 142 863 146
rect 867 142 868 146
rect 862 141 868 142
rect 942 146 948 147
rect 942 142 943 146
rect 947 142 948 146
rect 942 141 948 142
rect 1022 146 1028 147
rect 1022 142 1023 146
rect 1027 142 1028 146
rect 1022 141 1028 142
rect 1102 146 1108 147
rect 1102 142 1103 146
rect 1107 142 1108 146
rect 1102 141 1108 142
rect 1182 146 1188 147
rect 1182 142 1183 146
rect 1187 142 1188 146
rect 1182 141 1188 142
rect 1262 146 1268 147
rect 1262 142 1263 146
rect 1267 142 1268 146
rect 1262 141 1268 142
rect 1342 146 1348 147
rect 1342 142 1343 146
rect 1347 142 1348 146
rect 1342 141 1348 142
rect 1422 146 1428 147
rect 1422 142 1423 146
rect 1427 142 1428 146
rect 1422 141 1428 142
rect 1510 146 1516 147
rect 1510 142 1511 146
rect 1515 142 1516 146
rect 1510 141 1516 142
rect 1590 146 1596 147
rect 1590 142 1591 146
rect 1595 142 1596 146
rect 1590 141 1596 142
rect 1670 146 1676 147
rect 1670 142 1671 146
rect 1675 142 1676 146
rect 1670 141 1676 142
rect 1750 146 1756 147
rect 1750 142 1751 146
rect 1755 142 1756 146
rect 1750 141 1756 142
rect 1832 129 1834 157
rect 1872 145 1874 173
rect 1904 163 1906 173
rect 1984 163 1986 173
rect 2088 163 2090 173
rect 2216 163 2218 173
rect 2352 163 2354 173
rect 2488 163 2490 173
rect 2624 163 2626 173
rect 2744 163 2746 173
rect 2856 163 2858 173
rect 2960 163 2962 173
rect 3064 163 3066 173
rect 3160 163 3162 173
rect 3248 163 3250 173
rect 3344 163 3346 173
rect 3432 163 3434 173
rect 3512 163 3514 173
rect 1902 162 1908 163
rect 1902 158 1903 162
rect 1907 158 1908 162
rect 1902 157 1908 158
rect 1982 162 1988 163
rect 1982 158 1983 162
rect 1987 158 1988 162
rect 1982 157 1988 158
rect 2086 162 2092 163
rect 2086 158 2087 162
rect 2091 158 2092 162
rect 2086 157 2092 158
rect 2214 162 2220 163
rect 2214 158 2215 162
rect 2219 158 2220 162
rect 2214 157 2220 158
rect 2350 162 2356 163
rect 2350 158 2351 162
rect 2355 158 2356 162
rect 2350 157 2356 158
rect 2486 162 2492 163
rect 2486 158 2487 162
rect 2491 158 2492 162
rect 2486 157 2492 158
rect 2622 162 2628 163
rect 2622 158 2623 162
rect 2627 158 2628 162
rect 2622 157 2628 158
rect 2742 162 2748 163
rect 2742 158 2743 162
rect 2747 158 2748 162
rect 2742 157 2748 158
rect 2854 162 2860 163
rect 2854 158 2855 162
rect 2859 158 2860 162
rect 2854 157 2860 158
rect 2958 162 2964 163
rect 2958 158 2959 162
rect 2963 158 2964 162
rect 2958 157 2964 158
rect 3062 162 3068 163
rect 3062 158 3063 162
rect 3067 158 3068 162
rect 3062 157 3068 158
rect 3158 162 3164 163
rect 3158 158 3159 162
rect 3163 158 3164 162
rect 3158 157 3164 158
rect 3246 162 3252 163
rect 3246 158 3247 162
rect 3251 158 3252 162
rect 3246 157 3252 158
rect 3342 162 3348 163
rect 3342 158 3343 162
rect 3347 158 3348 162
rect 3342 157 3348 158
rect 3430 162 3436 163
rect 3430 158 3431 162
rect 3435 158 3436 162
rect 3430 157 3436 158
rect 3510 162 3516 163
rect 3510 158 3511 162
rect 3515 158 3516 162
rect 3510 157 3516 158
rect 3592 145 3594 173
rect 1870 144 1876 145
rect 1870 140 1871 144
rect 1875 140 1876 144
rect 1870 139 1876 140
rect 3590 144 3596 145
rect 3590 140 3591 144
rect 3595 140 3596 144
rect 3590 139 3596 140
rect 110 128 116 129
rect 110 124 111 128
rect 115 124 116 128
rect 110 123 116 124
rect 1830 128 1836 129
rect 1830 124 1831 128
rect 1835 124 1836 128
rect 1830 123 1836 124
rect 1870 127 1876 128
rect 1870 123 1871 127
rect 1875 123 1876 127
rect 3590 127 3596 128
rect 1870 122 1876 123
rect 1894 124 1900 125
rect 110 111 116 112
rect 110 107 111 111
rect 115 107 116 111
rect 1830 111 1836 112
rect 110 106 116 107
rect 134 108 140 109
rect 112 87 114 106
rect 134 104 135 108
rect 139 104 140 108
rect 134 103 140 104
rect 214 108 220 109
rect 214 104 215 108
rect 219 104 220 108
rect 214 103 220 104
rect 294 108 300 109
rect 294 104 295 108
rect 299 104 300 108
rect 294 103 300 104
rect 374 108 380 109
rect 374 104 375 108
rect 379 104 380 108
rect 374 103 380 104
rect 454 108 460 109
rect 454 104 455 108
rect 459 104 460 108
rect 454 103 460 104
rect 534 108 540 109
rect 534 104 535 108
rect 539 104 540 108
rect 534 103 540 104
rect 614 108 620 109
rect 614 104 615 108
rect 619 104 620 108
rect 614 103 620 104
rect 694 108 700 109
rect 694 104 695 108
rect 699 104 700 108
rect 694 103 700 104
rect 774 108 780 109
rect 774 104 775 108
rect 779 104 780 108
rect 774 103 780 104
rect 854 108 860 109
rect 854 104 855 108
rect 859 104 860 108
rect 854 103 860 104
rect 934 108 940 109
rect 934 104 935 108
rect 939 104 940 108
rect 934 103 940 104
rect 1014 108 1020 109
rect 1014 104 1015 108
rect 1019 104 1020 108
rect 1014 103 1020 104
rect 1094 108 1100 109
rect 1094 104 1095 108
rect 1099 104 1100 108
rect 1094 103 1100 104
rect 1174 108 1180 109
rect 1174 104 1175 108
rect 1179 104 1180 108
rect 1174 103 1180 104
rect 1254 108 1260 109
rect 1254 104 1255 108
rect 1259 104 1260 108
rect 1254 103 1260 104
rect 1334 108 1340 109
rect 1334 104 1335 108
rect 1339 104 1340 108
rect 1334 103 1340 104
rect 1414 108 1420 109
rect 1414 104 1415 108
rect 1419 104 1420 108
rect 1414 103 1420 104
rect 1502 108 1508 109
rect 1502 104 1503 108
rect 1507 104 1508 108
rect 1502 103 1508 104
rect 1582 108 1588 109
rect 1582 104 1583 108
rect 1587 104 1588 108
rect 1582 103 1588 104
rect 1662 108 1668 109
rect 1662 104 1663 108
rect 1667 104 1668 108
rect 1662 103 1668 104
rect 1742 108 1748 109
rect 1742 104 1743 108
rect 1747 104 1748 108
rect 1830 107 1831 111
rect 1835 107 1836 111
rect 1830 106 1836 107
rect 1742 103 1748 104
rect 136 87 138 103
rect 216 87 218 103
rect 296 87 298 103
rect 376 87 378 103
rect 456 87 458 103
rect 536 87 538 103
rect 616 87 618 103
rect 696 87 698 103
rect 776 87 778 103
rect 856 87 858 103
rect 936 87 938 103
rect 1016 87 1018 103
rect 1096 87 1098 103
rect 1176 87 1178 103
rect 1256 87 1258 103
rect 1336 87 1338 103
rect 1416 87 1418 103
rect 1504 87 1506 103
rect 1584 87 1586 103
rect 1664 87 1666 103
rect 1744 87 1746 103
rect 1832 87 1834 106
rect 1872 103 1874 122
rect 1894 120 1895 124
rect 1899 120 1900 124
rect 1894 119 1900 120
rect 1974 124 1980 125
rect 1974 120 1975 124
rect 1979 120 1980 124
rect 1974 119 1980 120
rect 2078 124 2084 125
rect 2078 120 2079 124
rect 2083 120 2084 124
rect 2078 119 2084 120
rect 2206 124 2212 125
rect 2206 120 2207 124
rect 2211 120 2212 124
rect 2206 119 2212 120
rect 2342 124 2348 125
rect 2342 120 2343 124
rect 2347 120 2348 124
rect 2342 119 2348 120
rect 2478 124 2484 125
rect 2478 120 2479 124
rect 2483 120 2484 124
rect 2478 119 2484 120
rect 2614 124 2620 125
rect 2614 120 2615 124
rect 2619 120 2620 124
rect 2614 119 2620 120
rect 2734 124 2740 125
rect 2734 120 2735 124
rect 2739 120 2740 124
rect 2734 119 2740 120
rect 2846 124 2852 125
rect 2846 120 2847 124
rect 2851 120 2852 124
rect 2846 119 2852 120
rect 2950 124 2956 125
rect 2950 120 2951 124
rect 2955 120 2956 124
rect 2950 119 2956 120
rect 3054 124 3060 125
rect 3054 120 3055 124
rect 3059 120 3060 124
rect 3054 119 3060 120
rect 3150 124 3156 125
rect 3150 120 3151 124
rect 3155 120 3156 124
rect 3150 119 3156 120
rect 3238 124 3244 125
rect 3238 120 3239 124
rect 3243 120 3244 124
rect 3238 119 3244 120
rect 3334 124 3340 125
rect 3334 120 3335 124
rect 3339 120 3340 124
rect 3334 119 3340 120
rect 3422 124 3428 125
rect 3422 120 3423 124
rect 3427 120 3428 124
rect 3422 119 3428 120
rect 3502 124 3508 125
rect 3502 120 3503 124
rect 3507 120 3508 124
rect 3590 123 3591 127
rect 3595 123 3596 127
rect 3590 122 3596 123
rect 3502 119 3508 120
rect 1896 103 1898 119
rect 1976 103 1978 119
rect 2080 103 2082 119
rect 2208 103 2210 119
rect 2344 103 2346 119
rect 2480 103 2482 119
rect 2616 103 2618 119
rect 2736 103 2738 119
rect 2848 103 2850 119
rect 2952 103 2954 119
rect 3056 103 3058 119
rect 3152 103 3154 119
rect 3240 103 3242 119
rect 3336 103 3338 119
rect 3424 103 3426 119
rect 3504 103 3506 119
rect 3592 103 3594 122
rect 1871 102 1875 103
rect 1871 97 1875 98
rect 1895 102 1899 103
rect 1895 97 1899 98
rect 1975 102 1979 103
rect 1975 97 1979 98
rect 2079 102 2083 103
rect 2079 97 2083 98
rect 2207 102 2211 103
rect 2207 97 2211 98
rect 2343 102 2347 103
rect 2343 97 2347 98
rect 2479 102 2483 103
rect 2479 97 2483 98
rect 2615 102 2619 103
rect 2615 97 2619 98
rect 2735 102 2739 103
rect 2735 97 2739 98
rect 2847 102 2851 103
rect 2847 97 2851 98
rect 2951 102 2955 103
rect 2951 97 2955 98
rect 3055 102 3059 103
rect 3055 97 3059 98
rect 3151 102 3155 103
rect 3151 97 3155 98
rect 3239 102 3243 103
rect 3239 97 3243 98
rect 3335 102 3339 103
rect 3335 97 3339 98
rect 3423 102 3427 103
rect 3423 97 3427 98
rect 3503 102 3507 103
rect 3503 97 3507 98
rect 3591 102 3595 103
rect 3591 97 3595 98
rect 111 86 115 87
rect 111 81 115 82
rect 135 86 139 87
rect 135 81 139 82
rect 215 86 219 87
rect 215 81 219 82
rect 295 86 299 87
rect 295 81 299 82
rect 375 86 379 87
rect 375 81 379 82
rect 455 86 459 87
rect 455 81 459 82
rect 535 86 539 87
rect 535 81 539 82
rect 615 86 619 87
rect 615 81 619 82
rect 695 86 699 87
rect 695 81 699 82
rect 775 86 779 87
rect 775 81 779 82
rect 855 86 859 87
rect 855 81 859 82
rect 935 86 939 87
rect 935 81 939 82
rect 1015 86 1019 87
rect 1015 81 1019 82
rect 1095 86 1099 87
rect 1095 81 1099 82
rect 1175 86 1179 87
rect 1175 81 1179 82
rect 1255 86 1259 87
rect 1255 81 1259 82
rect 1335 86 1339 87
rect 1335 81 1339 82
rect 1415 86 1419 87
rect 1415 81 1419 82
rect 1503 86 1507 87
rect 1503 81 1507 82
rect 1583 86 1587 87
rect 1583 81 1587 82
rect 1663 86 1667 87
rect 1663 81 1667 82
rect 1743 86 1747 87
rect 1743 81 1747 82
rect 1831 86 1835 87
rect 1831 81 1835 82
<< m4c >>
rect 111 3666 115 3670
rect 135 3666 139 3670
rect 215 3666 219 3670
rect 295 3666 299 3670
rect 1831 3666 1835 3670
rect 1871 3598 1875 3602
rect 2063 3598 2067 3602
rect 2151 3598 2155 3602
rect 2255 3598 2259 3602
rect 2367 3598 2371 3602
rect 2479 3598 2483 3602
rect 2591 3598 2595 3602
rect 2703 3598 2707 3602
rect 2815 3598 2819 3602
rect 2919 3598 2923 3602
rect 3015 3598 3019 3602
rect 3111 3598 3115 3602
rect 3207 3598 3211 3602
rect 3303 3598 3307 3602
rect 3399 3598 3403 3602
rect 3591 3598 3595 3602
rect 111 3590 115 3594
rect 143 3590 147 3594
rect 223 3590 227 3594
rect 303 3590 307 3594
rect 343 3590 347 3594
rect 471 3590 475 3594
rect 607 3590 611 3594
rect 743 3590 747 3594
rect 879 3590 883 3594
rect 999 3590 1003 3594
rect 1111 3590 1115 3594
rect 1223 3590 1227 3594
rect 1327 3590 1331 3594
rect 1423 3590 1427 3594
rect 1527 3590 1531 3594
rect 1631 3590 1635 3594
rect 1831 3590 1835 3594
rect 1871 3522 1875 3526
rect 2055 3522 2059 3526
rect 2087 3522 2091 3526
rect 2143 3522 2147 3526
rect 2167 3522 2171 3526
rect 2247 3522 2251 3526
rect 2263 3522 2267 3526
rect 2359 3522 2363 3526
rect 2367 3522 2371 3526
rect 2471 3522 2475 3526
rect 2487 3522 2491 3526
rect 2583 3522 2587 3526
rect 2615 3522 2619 3526
rect 2695 3522 2699 3526
rect 2743 3522 2747 3526
rect 2807 3522 2811 3526
rect 2871 3522 2875 3526
rect 2911 3522 2915 3526
rect 2991 3522 2995 3526
rect 3007 3522 3011 3526
rect 3103 3522 3107 3526
rect 3119 3522 3123 3526
rect 3199 3522 3203 3526
rect 3247 3522 3251 3526
rect 3295 3522 3299 3526
rect 3375 3522 3379 3526
rect 3391 3522 3395 3526
rect 3591 3522 3595 3526
rect 111 3514 115 3518
rect 135 3514 139 3518
rect 191 3514 195 3518
rect 215 3514 219 3518
rect 327 3514 331 3518
rect 335 3514 339 3518
rect 463 3514 467 3518
rect 471 3514 475 3518
rect 599 3514 603 3518
rect 623 3514 627 3518
rect 735 3514 739 3518
rect 775 3514 779 3518
rect 871 3514 875 3518
rect 919 3514 923 3518
rect 991 3514 995 3518
rect 1055 3514 1059 3518
rect 1103 3514 1107 3518
rect 1183 3514 1187 3518
rect 1215 3514 1219 3518
rect 1311 3514 1315 3518
rect 1319 3514 1323 3518
rect 1415 3514 1419 3518
rect 1439 3514 1443 3518
rect 1519 3514 1523 3518
rect 1567 3514 1571 3518
rect 1623 3514 1627 3518
rect 1831 3514 1835 3518
rect 111 3438 115 3442
rect 151 3438 155 3442
rect 199 3438 203 3442
rect 295 3438 299 3442
rect 335 3438 339 3442
rect 455 3438 459 3442
rect 479 3438 483 3442
rect 623 3438 627 3442
rect 631 3438 635 3442
rect 783 3438 787 3442
rect 791 3438 795 3442
rect 927 3438 931 3442
rect 959 3438 963 3442
rect 1063 3438 1067 3442
rect 1119 3438 1123 3442
rect 1191 3438 1195 3442
rect 1271 3438 1275 3442
rect 1319 3438 1323 3442
rect 1415 3438 1419 3442
rect 1447 3438 1451 3442
rect 1559 3438 1563 3442
rect 1575 3438 1579 3442
rect 1711 3438 1715 3442
rect 1831 3438 1835 3442
rect 1871 3438 1875 3442
rect 2095 3438 2099 3442
rect 2111 3438 2115 3442
rect 2175 3438 2179 3442
rect 2199 3438 2203 3442
rect 2271 3438 2275 3442
rect 2303 3438 2307 3442
rect 2375 3438 2379 3442
rect 2415 3438 2419 3442
rect 2495 3438 2499 3442
rect 2543 3438 2547 3442
rect 2623 3438 2627 3442
rect 2679 3438 2683 3442
rect 2751 3438 2755 3442
rect 2815 3438 2819 3442
rect 2879 3438 2883 3442
rect 2959 3438 2963 3442
rect 2999 3438 3003 3442
rect 3111 3438 3115 3442
rect 3127 3438 3131 3442
rect 3255 3438 3259 3442
rect 3263 3438 3267 3442
rect 3383 3438 3387 3442
rect 3423 3438 3427 3442
rect 3591 3438 3595 3442
rect 111 3362 115 3366
rect 143 3362 147 3366
rect 207 3362 211 3366
rect 287 3362 291 3366
rect 335 3362 339 3366
rect 447 3362 451 3366
rect 471 3362 475 3366
rect 615 3362 619 3366
rect 623 3362 627 3366
rect 783 3362 787 3366
rect 943 3362 947 3366
rect 951 3362 955 3366
rect 1103 3362 1107 3366
rect 1111 3362 1115 3366
rect 1263 3362 1267 3366
rect 1407 3362 1411 3366
rect 1423 3362 1427 3366
rect 1551 3362 1555 3366
rect 1583 3362 1587 3366
rect 1703 3362 1707 3366
rect 1743 3362 1747 3366
rect 1831 3362 1835 3366
rect 1871 3358 1875 3362
rect 2103 3358 2107 3362
rect 2127 3358 2131 3362
rect 2191 3358 2195 3362
rect 2223 3358 2227 3362
rect 2295 3358 2299 3362
rect 2335 3358 2339 3362
rect 2407 3358 2411 3362
rect 2455 3358 2459 3362
rect 2535 3358 2539 3362
rect 2583 3358 2587 3362
rect 2671 3358 2675 3362
rect 2719 3358 2723 3362
rect 2807 3358 2811 3362
rect 2863 3358 2867 3362
rect 2951 3358 2955 3362
rect 3007 3358 3011 3362
rect 3103 3358 3107 3362
rect 3159 3358 3163 3362
rect 3255 3358 3259 3362
rect 3311 3358 3315 3362
rect 3415 3358 3419 3362
rect 3471 3358 3475 3362
rect 3591 3358 3595 3362
rect 111 3282 115 3286
rect 215 3282 219 3286
rect 343 3282 347 3286
rect 351 3282 355 3286
rect 455 3282 459 3286
rect 479 3282 483 3286
rect 575 3282 579 3286
rect 631 3282 635 3286
rect 703 3282 707 3286
rect 791 3282 795 3286
rect 839 3282 843 3286
rect 951 3282 955 3286
rect 983 3282 987 3286
rect 1111 3282 1115 3286
rect 1119 3282 1123 3286
rect 1255 3282 1259 3286
rect 1271 3282 1275 3286
rect 1383 3282 1387 3286
rect 1431 3282 1435 3286
rect 1511 3282 1515 3286
rect 1591 3282 1595 3286
rect 1639 3282 1643 3286
rect 1751 3282 1755 3286
rect 1831 3282 1835 3286
rect 1871 3270 1875 3274
rect 2135 3270 2139 3274
rect 2231 3270 2235 3274
rect 2279 3270 2283 3274
rect 2343 3270 2347 3274
rect 2415 3270 2419 3274
rect 2463 3270 2467 3274
rect 2551 3270 2555 3274
rect 2591 3270 2595 3274
rect 2687 3270 2691 3274
rect 2727 3270 2731 3274
rect 2823 3270 2827 3274
rect 2871 3270 2875 3274
rect 2959 3270 2963 3274
rect 3015 3270 3019 3274
rect 3095 3270 3099 3274
rect 3167 3270 3171 3274
rect 3231 3270 3235 3274
rect 3319 3270 3323 3274
rect 3375 3270 3379 3274
rect 3479 3270 3483 3274
rect 3511 3270 3515 3274
rect 3591 3270 3595 3274
rect 111 3206 115 3210
rect 343 3206 347 3210
rect 447 3206 451 3210
rect 487 3206 491 3210
rect 567 3206 571 3210
rect 575 3206 579 3210
rect 663 3206 667 3210
rect 695 3206 699 3210
rect 767 3206 771 3210
rect 831 3206 835 3210
rect 887 3206 891 3210
rect 975 3206 979 3210
rect 1023 3206 1027 3210
rect 1111 3206 1115 3210
rect 1191 3206 1195 3210
rect 1247 3206 1251 3210
rect 1375 3206 1379 3210
rect 1503 3206 1507 3210
rect 1567 3206 1571 3210
rect 1631 3206 1635 3210
rect 1743 3206 1747 3210
rect 1831 3206 1835 3210
rect 1871 3190 1875 3194
rect 1895 3190 1899 3194
rect 1991 3190 1995 3194
rect 2119 3190 2123 3194
rect 2127 3190 2131 3194
rect 2247 3190 2251 3194
rect 2271 3190 2275 3194
rect 2383 3190 2387 3194
rect 2407 3190 2411 3194
rect 2511 3190 2515 3194
rect 2543 3190 2547 3194
rect 2639 3190 2643 3194
rect 2679 3190 2683 3194
rect 2767 3190 2771 3194
rect 2815 3190 2819 3194
rect 2895 3190 2899 3194
rect 2951 3190 2955 3194
rect 3031 3190 3035 3194
rect 3087 3190 3091 3194
rect 3175 3190 3179 3194
rect 3223 3190 3227 3194
rect 3327 3190 3331 3194
rect 3367 3190 3371 3194
rect 3487 3190 3491 3194
rect 3503 3190 3507 3194
rect 3591 3190 3595 3194
rect 111 3126 115 3130
rect 495 3126 499 3130
rect 583 3126 587 3130
rect 591 3126 595 3130
rect 671 3126 675 3130
rect 759 3126 763 3130
rect 775 3126 779 3130
rect 847 3126 851 3130
rect 895 3126 899 3130
rect 935 3126 939 3130
rect 1023 3126 1027 3130
rect 1031 3126 1035 3130
rect 1111 3126 1115 3130
rect 1199 3126 1203 3130
rect 1287 3126 1291 3130
rect 1375 3126 1379 3130
rect 1383 3126 1387 3130
rect 1575 3126 1579 3130
rect 1751 3126 1755 3130
rect 1831 3126 1835 3130
rect 1871 3098 1875 3102
rect 1903 3098 1907 3102
rect 1999 3098 2003 3102
rect 2015 3098 2019 3102
rect 2127 3098 2131 3102
rect 2191 3098 2195 3102
rect 2255 3098 2259 3102
rect 2391 3098 2395 3102
rect 2407 3098 2411 3102
rect 2519 3098 2523 3102
rect 2647 3098 2651 3102
rect 2655 3098 2659 3102
rect 2775 3098 2779 3102
rect 2903 3098 2907 3102
rect 2935 3098 2939 3102
rect 3039 3098 3043 3102
rect 3183 3098 3187 3102
rect 3231 3098 3235 3102
rect 3335 3098 3339 3102
rect 3495 3098 3499 3102
rect 3511 3098 3515 3102
rect 3591 3098 3595 3102
rect 111 3046 115 3050
rect 543 3046 547 3050
rect 583 3046 587 3050
rect 623 3046 627 3050
rect 663 3046 667 3050
rect 711 3046 715 3050
rect 751 3046 755 3050
rect 807 3046 811 3050
rect 839 3046 843 3050
rect 903 3046 907 3050
rect 927 3046 931 3050
rect 999 3046 1003 3050
rect 1015 3046 1019 3050
rect 1087 3046 1091 3050
rect 1103 3046 1107 3050
rect 1183 3046 1187 3050
rect 1191 3046 1195 3050
rect 1279 3046 1283 3050
rect 1367 3046 1371 3050
rect 1375 3046 1379 3050
rect 1471 3046 1475 3050
rect 1831 3046 1835 3050
rect 1871 3014 1875 3018
rect 1895 3014 1899 3018
rect 2007 3014 2011 3018
rect 2047 3014 2051 3018
rect 2183 3014 2187 3018
rect 2223 3014 2227 3018
rect 2391 3014 2395 3018
rect 2399 3014 2403 3018
rect 2543 3014 2547 3018
rect 2647 3014 2651 3018
rect 2687 3014 2691 3018
rect 2815 3014 2819 3018
rect 2927 3014 2931 3018
rect 3039 3014 3043 3018
rect 3143 3014 3147 3018
rect 3223 3014 3227 3018
rect 3239 3014 3243 3018
rect 3335 3014 3339 3018
rect 3423 3014 3427 3018
rect 3503 3014 3507 3018
rect 3591 3014 3595 3018
rect 111 2970 115 2974
rect 471 2970 475 2974
rect 551 2970 555 2974
rect 575 2970 579 2974
rect 631 2970 635 2974
rect 687 2970 691 2974
rect 719 2970 723 2974
rect 807 2970 811 2974
rect 815 2970 819 2974
rect 911 2970 915 2974
rect 943 2970 947 2974
rect 1007 2970 1011 2974
rect 1087 2970 1091 2974
rect 1095 2970 1099 2974
rect 1191 2970 1195 2974
rect 1247 2970 1251 2974
rect 1287 2970 1291 2974
rect 1383 2970 1387 2974
rect 1415 2970 1419 2974
rect 1479 2970 1483 2974
rect 1591 2970 1595 2974
rect 1751 2970 1755 2974
rect 1831 2970 1835 2974
rect 1871 2938 1875 2942
rect 1903 2938 1907 2942
rect 2055 2938 2059 2942
rect 2087 2938 2091 2942
rect 2231 2938 2235 2942
rect 2295 2938 2299 2942
rect 2399 2938 2403 2942
rect 2487 2938 2491 2942
rect 2551 2938 2555 2942
rect 2671 2938 2675 2942
rect 2695 2938 2699 2942
rect 2823 2938 2827 2942
rect 2839 2938 2843 2942
rect 2935 2938 2939 2942
rect 2999 2938 3003 2942
rect 3047 2938 3051 2942
rect 3151 2938 3155 2942
rect 3247 2938 3251 2942
rect 3303 2938 3307 2942
rect 3343 2938 3347 2942
rect 3431 2938 3435 2942
rect 3455 2938 3459 2942
rect 3511 2938 3515 2942
rect 3591 2938 3595 2942
rect 111 2894 115 2898
rect 311 2894 315 2898
rect 431 2894 435 2898
rect 463 2894 467 2898
rect 551 2894 555 2898
rect 567 2894 571 2898
rect 679 2894 683 2898
rect 799 2894 803 2898
rect 815 2894 819 2898
rect 935 2894 939 2898
rect 951 2894 955 2898
rect 1079 2894 1083 2898
rect 1087 2894 1091 2898
rect 1223 2894 1227 2898
rect 1239 2894 1243 2898
rect 1359 2894 1363 2898
rect 1407 2894 1411 2898
rect 1495 2894 1499 2898
rect 1583 2894 1587 2898
rect 1631 2894 1635 2898
rect 1743 2894 1747 2898
rect 1831 2894 1835 2898
rect 1871 2854 1875 2858
rect 1895 2854 1899 2858
rect 2079 2854 2083 2858
rect 2135 2854 2139 2858
rect 2263 2854 2267 2858
rect 2287 2854 2291 2858
rect 2391 2854 2395 2858
rect 2479 2854 2483 2858
rect 2519 2854 2523 2858
rect 2647 2854 2651 2858
rect 2663 2854 2667 2858
rect 2767 2854 2771 2858
rect 2831 2854 2835 2858
rect 2887 2854 2891 2858
rect 2991 2854 2995 2858
rect 3007 2854 3011 2858
rect 3135 2854 3139 2858
rect 3143 2854 3147 2858
rect 3295 2854 3299 2858
rect 3447 2854 3451 2858
rect 3591 2854 3595 2858
rect 111 2818 115 2822
rect 167 2818 171 2822
rect 303 2818 307 2822
rect 319 2818 323 2822
rect 439 2818 443 2822
rect 447 2818 451 2822
rect 559 2818 563 2822
rect 607 2818 611 2822
rect 687 2818 691 2822
rect 783 2818 787 2822
rect 823 2818 827 2822
rect 959 2818 963 2822
rect 1095 2818 1099 2822
rect 1143 2818 1147 2822
rect 1231 2818 1235 2822
rect 1335 2818 1339 2822
rect 1367 2818 1371 2822
rect 1503 2818 1507 2822
rect 1535 2818 1539 2822
rect 1639 2818 1643 2822
rect 1735 2818 1739 2822
rect 1751 2818 1755 2822
rect 1831 2818 1835 2822
rect 1871 2770 1875 2774
rect 2143 2770 2147 2774
rect 2231 2770 2235 2774
rect 2271 2770 2275 2774
rect 2311 2770 2315 2774
rect 2391 2770 2395 2774
rect 2399 2770 2403 2774
rect 2471 2770 2475 2774
rect 2527 2770 2531 2774
rect 2551 2770 2555 2774
rect 2639 2770 2643 2774
rect 2655 2770 2659 2774
rect 2727 2770 2731 2774
rect 2775 2770 2779 2774
rect 2815 2770 2819 2774
rect 2895 2770 2899 2774
rect 2903 2770 2907 2774
rect 2991 2770 2995 2774
rect 3015 2770 3019 2774
rect 3143 2770 3147 2774
rect 3591 2770 3595 2774
rect 111 2738 115 2742
rect 135 2738 139 2742
rect 159 2738 163 2742
rect 247 2738 251 2742
rect 295 2738 299 2742
rect 391 2738 395 2742
rect 439 2738 443 2742
rect 551 2738 555 2742
rect 599 2738 603 2742
rect 711 2738 715 2742
rect 775 2738 779 2742
rect 879 2738 883 2742
rect 951 2738 955 2742
rect 1039 2738 1043 2742
rect 1135 2738 1139 2742
rect 1199 2738 1203 2742
rect 1327 2738 1331 2742
rect 1359 2738 1363 2742
rect 1519 2738 1523 2742
rect 1527 2738 1531 2742
rect 1687 2738 1691 2742
rect 1727 2738 1731 2742
rect 1831 2738 1835 2742
rect 1871 2694 1875 2698
rect 2223 2694 2227 2698
rect 2239 2694 2243 2698
rect 2303 2694 2307 2698
rect 2319 2694 2323 2698
rect 2383 2694 2387 2698
rect 2399 2694 2403 2698
rect 2463 2694 2467 2698
rect 2479 2694 2483 2698
rect 2543 2694 2547 2698
rect 2559 2694 2563 2698
rect 2631 2694 2635 2698
rect 2639 2694 2643 2698
rect 2719 2694 2723 2698
rect 2799 2694 2803 2698
rect 2807 2694 2811 2698
rect 2879 2694 2883 2698
rect 2895 2694 2899 2698
rect 2959 2694 2963 2698
rect 2983 2694 2987 2698
rect 3591 2694 3595 2698
rect 111 2662 115 2666
rect 143 2662 147 2666
rect 255 2662 259 2666
rect 399 2662 403 2666
rect 551 2662 555 2666
rect 559 2662 563 2666
rect 711 2662 715 2666
rect 719 2662 723 2666
rect 879 2662 883 2666
rect 887 2662 891 2666
rect 1047 2662 1051 2666
rect 1207 2662 1211 2666
rect 1215 2662 1219 2666
rect 1367 2662 1371 2666
rect 1391 2662 1395 2666
rect 1527 2662 1531 2666
rect 1567 2662 1571 2666
rect 1695 2662 1699 2666
rect 1831 2662 1835 2666
rect 1871 2610 1875 2614
rect 2191 2610 2195 2614
rect 2247 2610 2251 2614
rect 2271 2610 2275 2614
rect 2327 2610 2331 2614
rect 2351 2610 2355 2614
rect 2407 2610 2411 2614
rect 2431 2610 2435 2614
rect 2487 2610 2491 2614
rect 2511 2610 2515 2614
rect 2567 2610 2571 2614
rect 2591 2610 2595 2614
rect 2647 2610 2651 2614
rect 2671 2610 2675 2614
rect 2727 2610 2731 2614
rect 2751 2610 2755 2614
rect 2807 2610 2811 2614
rect 2831 2610 2835 2614
rect 2887 2610 2891 2614
rect 2911 2610 2915 2614
rect 2967 2610 2971 2614
rect 2991 2610 2995 2614
rect 3591 2610 3595 2614
rect 111 2582 115 2586
rect 135 2582 139 2586
rect 159 2582 163 2586
rect 247 2582 251 2586
rect 279 2582 283 2586
rect 391 2582 395 2586
rect 415 2582 419 2586
rect 543 2582 547 2586
rect 559 2582 563 2586
rect 703 2582 707 2586
rect 847 2582 851 2586
rect 871 2582 875 2586
rect 983 2582 987 2586
rect 1039 2582 1043 2586
rect 1119 2582 1123 2586
rect 1207 2582 1211 2586
rect 1255 2582 1259 2586
rect 1383 2582 1387 2586
rect 1391 2582 1395 2586
rect 1527 2582 1531 2586
rect 1559 2582 1563 2586
rect 1831 2582 1835 2586
rect 1871 2526 1875 2530
rect 2119 2526 2123 2530
rect 2183 2526 2187 2530
rect 2207 2526 2211 2530
rect 2263 2526 2267 2530
rect 2303 2526 2307 2530
rect 2343 2526 2347 2530
rect 2399 2526 2403 2530
rect 2423 2526 2427 2530
rect 2495 2526 2499 2530
rect 2503 2526 2507 2530
rect 2583 2526 2587 2530
rect 2591 2526 2595 2530
rect 2663 2526 2667 2530
rect 2687 2526 2691 2530
rect 2743 2526 2747 2530
rect 2783 2526 2787 2530
rect 2823 2526 2827 2530
rect 2879 2526 2883 2530
rect 2903 2526 2907 2530
rect 2975 2526 2979 2530
rect 2983 2526 2987 2530
rect 3079 2526 3083 2530
rect 3591 2526 3595 2530
rect 111 2502 115 2506
rect 167 2502 171 2506
rect 287 2502 291 2506
rect 335 2502 339 2506
rect 415 2502 419 2506
rect 423 2502 427 2506
rect 503 2502 507 2506
rect 567 2502 571 2506
rect 599 2502 603 2506
rect 703 2502 707 2506
rect 711 2502 715 2506
rect 815 2502 819 2506
rect 855 2502 859 2506
rect 935 2502 939 2506
rect 991 2502 995 2506
rect 1063 2502 1067 2506
rect 1127 2502 1131 2506
rect 1191 2502 1195 2506
rect 1263 2502 1267 2506
rect 1327 2502 1331 2506
rect 1399 2502 1403 2506
rect 1471 2502 1475 2506
rect 1535 2502 1539 2506
rect 1831 2502 1835 2506
rect 1871 2446 1875 2450
rect 1903 2446 1907 2450
rect 1991 2446 1995 2450
rect 2111 2446 2115 2450
rect 2127 2446 2131 2450
rect 2215 2446 2219 2450
rect 2247 2446 2251 2450
rect 2311 2446 2315 2450
rect 2391 2446 2395 2450
rect 2407 2446 2411 2450
rect 2503 2446 2507 2450
rect 2535 2446 2539 2450
rect 2599 2446 2603 2450
rect 2671 2446 2675 2450
rect 2695 2446 2699 2450
rect 2791 2446 2795 2450
rect 2807 2446 2811 2450
rect 2887 2446 2891 2450
rect 2943 2446 2947 2450
rect 2983 2446 2987 2450
rect 3079 2446 3083 2450
rect 3087 2446 3091 2450
rect 3215 2446 3219 2450
rect 3591 2446 3595 2450
rect 111 2418 115 2422
rect 327 2418 331 2422
rect 383 2418 387 2422
rect 407 2418 411 2422
rect 463 2418 467 2422
rect 495 2418 499 2422
rect 543 2418 547 2422
rect 591 2418 595 2422
rect 623 2418 627 2422
rect 695 2418 699 2422
rect 703 2418 707 2422
rect 783 2418 787 2422
rect 807 2418 811 2422
rect 863 2418 867 2422
rect 927 2418 931 2422
rect 943 2418 947 2422
rect 1023 2418 1027 2422
rect 1055 2418 1059 2422
rect 1103 2418 1107 2422
rect 1183 2418 1187 2422
rect 1263 2418 1267 2422
rect 1319 2418 1323 2422
rect 1351 2418 1355 2422
rect 1439 2418 1443 2422
rect 1463 2418 1467 2422
rect 1527 2418 1531 2422
rect 1831 2418 1835 2422
rect 1871 2362 1875 2366
rect 1895 2362 1899 2366
rect 1983 2362 1987 2366
rect 2015 2362 2019 2366
rect 2103 2362 2107 2366
rect 2175 2362 2179 2366
rect 2239 2362 2243 2366
rect 2343 2362 2347 2366
rect 2383 2362 2387 2366
rect 2511 2362 2515 2366
rect 2527 2362 2531 2366
rect 2663 2362 2667 2366
rect 2671 2362 2675 2366
rect 2799 2362 2803 2366
rect 2823 2362 2827 2366
rect 2935 2362 2939 2366
rect 2959 2362 2963 2366
rect 3071 2362 3075 2366
rect 3079 2362 3083 2366
rect 3191 2362 3195 2366
rect 3207 2362 3211 2366
rect 3303 2362 3307 2366
rect 3415 2362 3419 2366
rect 3503 2362 3507 2366
rect 3591 2362 3595 2366
rect 111 2342 115 2346
rect 391 2342 395 2346
rect 471 2342 475 2346
rect 551 2342 555 2346
rect 631 2342 635 2346
rect 711 2342 715 2346
rect 791 2342 795 2346
rect 871 2342 875 2346
rect 951 2342 955 2346
rect 1031 2342 1035 2346
rect 1111 2342 1115 2346
rect 1191 2342 1195 2346
rect 1271 2342 1275 2346
rect 1359 2342 1363 2346
rect 1407 2342 1411 2346
rect 1447 2342 1451 2346
rect 1487 2342 1491 2346
rect 1535 2342 1539 2346
rect 1567 2342 1571 2346
rect 1647 2342 1651 2346
rect 1831 2342 1835 2346
rect 1871 2286 1875 2290
rect 1903 2286 1907 2290
rect 2023 2286 2027 2290
rect 2031 2286 2035 2290
rect 2183 2286 2187 2290
rect 2351 2286 2355 2290
rect 2367 2286 2371 2290
rect 2519 2286 2523 2290
rect 2575 2286 2579 2290
rect 2679 2286 2683 2290
rect 2791 2286 2795 2290
rect 2831 2286 2835 2290
rect 2967 2286 2971 2290
rect 3023 2286 3027 2290
rect 3087 2286 3091 2290
rect 3199 2286 3203 2290
rect 3255 2286 3259 2290
rect 3311 2286 3315 2290
rect 3423 2286 3427 2290
rect 3495 2286 3499 2290
rect 3511 2286 3515 2290
rect 3591 2286 3595 2290
rect 111 2258 115 2262
rect 135 2258 139 2262
rect 215 2258 219 2262
rect 295 2258 299 2262
rect 383 2258 387 2262
rect 519 2258 523 2262
rect 671 2258 675 2262
rect 831 2258 835 2262
rect 999 2258 1003 2262
rect 1159 2258 1163 2262
rect 1311 2258 1315 2262
rect 1399 2258 1403 2262
rect 1455 2258 1459 2262
rect 1479 2258 1483 2262
rect 1559 2258 1563 2262
rect 1607 2258 1611 2262
rect 1639 2258 1643 2262
rect 1743 2258 1747 2262
rect 1831 2258 1835 2262
rect 1871 2190 1875 2194
rect 1895 2190 1899 2194
rect 2023 2190 2027 2194
rect 2175 2190 2179 2194
rect 2199 2190 2203 2194
rect 2295 2190 2299 2194
rect 2359 2190 2363 2194
rect 2399 2190 2403 2194
rect 2519 2190 2523 2194
rect 2567 2190 2571 2194
rect 2639 2190 2643 2194
rect 2759 2190 2763 2194
rect 2783 2190 2787 2194
rect 2879 2190 2883 2194
rect 2991 2190 2995 2194
rect 3015 2190 3019 2194
rect 3095 2190 3099 2194
rect 3199 2190 3203 2194
rect 3247 2190 3251 2194
rect 3303 2190 3307 2194
rect 3407 2190 3411 2194
rect 3487 2190 3491 2194
rect 3503 2190 3507 2194
rect 3591 2190 3595 2194
rect 111 2178 115 2182
rect 143 2178 147 2182
rect 191 2178 195 2182
rect 223 2178 227 2182
rect 303 2178 307 2182
rect 311 2178 315 2182
rect 391 2178 395 2182
rect 463 2178 467 2182
rect 527 2178 531 2182
rect 639 2178 643 2182
rect 679 2178 683 2182
rect 823 2178 827 2182
rect 839 2178 843 2182
rect 1007 2178 1011 2182
rect 1015 2178 1019 2182
rect 1167 2178 1171 2182
rect 1199 2178 1203 2182
rect 1319 2178 1323 2182
rect 1391 2178 1395 2182
rect 1463 2178 1467 2182
rect 1583 2178 1587 2182
rect 1615 2178 1619 2182
rect 1751 2178 1755 2182
rect 1831 2178 1835 2182
rect 111 2098 115 2102
rect 183 2098 187 2102
rect 215 2098 219 2102
rect 303 2098 307 2102
rect 359 2098 363 2102
rect 455 2098 459 2102
rect 519 2098 523 2102
rect 631 2098 635 2102
rect 703 2098 707 2102
rect 815 2098 819 2102
rect 895 2098 899 2102
rect 1007 2098 1011 2102
rect 1103 2098 1107 2102
rect 1191 2098 1195 2102
rect 1311 2098 1315 2102
rect 1383 2098 1387 2102
rect 1527 2098 1531 2102
rect 1575 2098 1579 2102
rect 1743 2098 1747 2102
rect 1831 2098 1835 2102
rect 1871 2102 1875 2106
rect 2175 2102 2179 2106
rect 2207 2102 2211 2106
rect 2271 2102 2275 2106
rect 2303 2102 2307 2106
rect 2375 2102 2379 2106
rect 2407 2102 2411 2106
rect 2487 2102 2491 2106
rect 2527 2102 2531 2106
rect 2607 2102 2611 2106
rect 2647 2102 2651 2106
rect 2727 2102 2731 2106
rect 2767 2102 2771 2106
rect 2847 2102 2851 2106
rect 2887 2102 2891 2106
rect 2967 2102 2971 2106
rect 2999 2102 3003 2106
rect 3079 2102 3083 2106
rect 3103 2102 3107 2106
rect 3191 2102 3195 2106
rect 3207 2102 3211 2106
rect 3303 2102 3307 2106
rect 3311 2102 3315 2106
rect 3415 2102 3419 2106
rect 3511 2102 3515 2106
rect 3591 2102 3595 2106
rect 111 2022 115 2026
rect 143 2022 147 2026
rect 223 2022 227 2026
rect 263 2022 267 2026
rect 367 2022 371 2026
rect 383 2022 387 2026
rect 495 2022 499 2026
rect 527 2022 531 2026
rect 607 2022 611 2026
rect 711 2022 715 2026
rect 719 2022 723 2026
rect 823 2022 827 2026
rect 903 2022 907 2026
rect 927 2022 931 2026
rect 1023 2022 1027 2026
rect 1111 2022 1115 2026
rect 1207 2022 1211 2026
rect 1295 2022 1299 2026
rect 1319 2022 1323 2026
rect 1391 2022 1395 2026
rect 1487 2022 1491 2026
rect 1535 2022 1539 2026
rect 1583 2022 1587 2026
rect 1671 2022 1675 2026
rect 1751 2022 1755 2026
rect 1831 2022 1835 2026
rect 1871 2022 1875 2026
rect 2071 2022 2075 2026
rect 2167 2022 2171 2026
rect 2207 2022 2211 2026
rect 2263 2022 2267 2026
rect 2359 2022 2363 2026
rect 2367 2022 2371 2026
rect 2479 2022 2483 2026
rect 2519 2022 2523 2026
rect 2599 2022 2603 2026
rect 2679 2022 2683 2026
rect 2719 2022 2723 2026
rect 2839 2022 2843 2026
rect 2847 2022 2851 2026
rect 2959 2022 2963 2026
rect 3015 2022 3019 2026
rect 3071 2022 3075 2026
rect 3183 2022 3187 2026
rect 3295 2022 3299 2026
rect 3351 2022 3355 2026
rect 3407 2022 3411 2026
rect 3503 2022 3507 2026
rect 3591 2022 3595 2026
rect 1871 1946 1875 1950
rect 1903 1946 1907 1950
rect 2007 1946 2011 1950
rect 2079 1946 2083 1950
rect 2135 1946 2139 1950
rect 2215 1946 2219 1950
rect 2255 1946 2259 1950
rect 2367 1946 2371 1950
rect 2375 1946 2379 1950
rect 2487 1946 2491 1950
rect 2527 1946 2531 1950
rect 2599 1946 2603 1950
rect 2687 1946 2691 1950
rect 2719 1946 2723 1950
rect 2839 1946 2843 1950
rect 2855 1946 2859 1950
rect 3023 1946 3027 1950
rect 3191 1946 3195 1950
rect 3359 1946 3363 1950
rect 3511 1946 3515 1950
rect 3591 1946 3595 1950
rect 111 1938 115 1942
rect 135 1938 139 1942
rect 167 1938 171 1942
rect 255 1938 259 1942
rect 327 1938 331 1942
rect 375 1938 379 1942
rect 487 1938 491 1942
rect 599 1938 603 1942
rect 647 1938 651 1942
rect 711 1938 715 1942
rect 799 1938 803 1942
rect 815 1938 819 1942
rect 919 1938 923 1942
rect 943 1938 947 1942
rect 1015 1938 1019 1942
rect 1079 1938 1083 1942
rect 1103 1938 1107 1942
rect 1199 1938 1203 1942
rect 1215 1938 1219 1942
rect 1287 1938 1291 1942
rect 1351 1938 1355 1942
rect 1383 1938 1387 1942
rect 1479 1938 1483 1942
rect 1487 1938 1491 1942
rect 1575 1938 1579 1942
rect 1623 1938 1627 1942
rect 1663 1938 1667 1942
rect 1743 1938 1747 1942
rect 1831 1938 1835 1942
rect 1871 1870 1875 1874
rect 1895 1870 1899 1874
rect 1991 1870 1995 1874
rect 1999 1870 2003 1874
rect 2119 1870 2123 1874
rect 2127 1870 2131 1874
rect 2247 1870 2251 1874
rect 2367 1870 2371 1874
rect 2383 1870 2387 1874
rect 2479 1870 2483 1874
rect 2519 1870 2523 1874
rect 2591 1870 2595 1874
rect 2655 1870 2659 1874
rect 2711 1870 2715 1874
rect 2807 1870 2811 1874
rect 2831 1870 2835 1874
rect 2975 1870 2979 1874
rect 3151 1870 3155 1874
rect 3335 1870 3339 1874
rect 3503 1870 3507 1874
rect 3591 1870 3595 1874
rect 111 1862 115 1866
rect 159 1862 163 1866
rect 175 1862 179 1866
rect 303 1862 307 1866
rect 335 1862 339 1866
rect 447 1862 451 1866
rect 495 1862 499 1866
rect 599 1862 603 1866
rect 655 1862 659 1866
rect 751 1862 755 1866
rect 807 1862 811 1866
rect 903 1862 907 1866
rect 951 1862 955 1866
rect 1055 1862 1059 1866
rect 1087 1862 1091 1866
rect 1207 1862 1211 1866
rect 1223 1862 1227 1866
rect 1351 1862 1355 1866
rect 1359 1862 1363 1866
rect 1487 1862 1491 1866
rect 1495 1862 1499 1866
rect 1631 1862 1635 1866
rect 1751 1862 1755 1866
rect 1831 1862 1835 1866
rect 111 1782 115 1786
rect 151 1782 155 1786
rect 247 1782 251 1786
rect 295 1782 299 1786
rect 423 1782 427 1786
rect 439 1782 443 1786
rect 591 1782 595 1786
rect 743 1782 747 1786
rect 751 1782 755 1786
rect 895 1782 899 1786
rect 1023 1782 1027 1786
rect 1047 1782 1051 1786
rect 1143 1782 1147 1786
rect 1199 1782 1203 1786
rect 1263 1782 1267 1786
rect 1343 1782 1347 1786
rect 1391 1782 1395 1786
rect 1479 1782 1483 1786
rect 1623 1782 1627 1786
rect 1743 1782 1747 1786
rect 1831 1782 1835 1786
rect 1871 1782 1875 1786
rect 1903 1782 1907 1786
rect 1999 1782 2003 1786
rect 2031 1782 2035 1786
rect 2127 1782 2131 1786
rect 2191 1782 2195 1786
rect 2255 1782 2259 1786
rect 2359 1782 2363 1786
rect 2391 1782 2395 1786
rect 2527 1782 2531 1786
rect 2663 1782 2667 1786
rect 2687 1782 2691 1786
rect 2815 1782 2819 1786
rect 2839 1782 2843 1786
rect 2983 1782 2987 1786
rect 3119 1782 3123 1786
rect 3159 1782 3163 1786
rect 3255 1782 3259 1786
rect 3343 1782 3347 1786
rect 3391 1782 3395 1786
rect 3511 1782 3515 1786
rect 3591 1782 3595 1786
rect 111 1702 115 1706
rect 191 1702 195 1706
rect 255 1702 259 1706
rect 311 1702 315 1706
rect 431 1702 435 1706
rect 447 1702 451 1706
rect 591 1702 595 1706
rect 599 1702 603 1706
rect 743 1702 747 1706
rect 759 1702 763 1706
rect 895 1702 899 1706
rect 903 1702 907 1706
rect 1031 1702 1035 1706
rect 1039 1702 1043 1706
rect 1151 1702 1155 1706
rect 1183 1702 1187 1706
rect 1271 1702 1275 1706
rect 1319 1702 1323 1706
rect 1399 1702 1403 1706
rect 1447 1702 1451 1706
rect 1575 1702 1579 1706
rect 1711 1702 1715 1706
rect 1831 1702 1835 1706
rect 1871 1702 1875 1706
rect 1895 1702 1899 1706
rect 1991 1702 1995 1706
rect 2023 1702 2027 1706
rect 2135 1702 2139 1706
rect 2183 1702 2187 1706
rect 2295 1702 2299 1706
rect 2351 1702 2355 1706
rect 2471 1702 2475 1706
rect 2519 1702 2523 1706
rect 2647 1702 2651 1706
rect 2679 1702 2683 1706
rect 2815 1702 2819 1706
rect 2831 1702 2835 1706
rect 2967 1702 2971 1706
rect 2975 1702 2979 1706
rect 3111 1702 3115 1706
rect 3247 1702 3251 1706
rect 3383 1702 3387 1706
rect 3503 1702 3507 1706
rect 3591 1702 3595 1706
rect 111 1618 115 1622
rect 167 1618 171 1622
rect 183 1618 187 1622
rect 303 1618 307 1622
rect 351 1618 355 1622
rect 439 1618 443 1622
rect 543 1618 547 1622
rect 583 1618 587 1622
rect 727 1618 731 1622
rect 735 1618 739 1622
rect 887 1618 891 1622
rect 903 1618 907 1622
rect 1031 1618 1035 1622
rect 1071 1618 1075 1622
rect 1175 1618 1179 1622
rect 1223 1618 1227 1622
rect 1311 1618 1315 1622
rect 1359 1618 1363 1622
rect 1439 1618 1443 1622
rect 1495 1618 1499 1622
rect 1567 1618 1571 1622
rect 1623 1618 1627 1622
rect 1703 1618 1707 1622
rect 1743 1618 1747 1622
rect 1831 1618 1835 1622
rect 1871 1622 1875 1626
rect 1903 1622 1907 1626
rect 1975 1622 1979 1626
rect 1999 1622 2003 1626
rect 2095 1622 2099 1626
rect 2143 1622 2147 1626
rect 2231 1622 2235 1626
rect 2303 1622 2307 1626
rect 2367 1622 2371 1626
rect 2479 1622 2483 1626
rect 2503 1622 2507 1626
rect 2639 1622 2643 1626
rect 2655 1622 2659 1626
rect 2775 1622 2779 1626
rect 2823 1622 2827 1626
rect 2911 1622 2915 1626
rect 2975 1622 2979 1626
rect 3055 1622 3059 1626
rect 3119 1622 3123 1626
rect 3207 1622 3211 1626
rect 3255 1622 3259 1626
rect 3367 1622 3371 1626
rect 3391 1622 3395 1626
rect 3511 1622 3515 1626
rect 3591 1622 3595 1626
rect 111 1538 115 1542
rect 143 1538 147 1542
rect 175 1538 179 1542
rect 247 1538 251 1542
rect 359 1538 363 1542
rect 383 1538 387 1542
rect 527 1538 531 1542
rect 551 1538 555 1542
rect 671 1538 675 1542
rect 735 1538 739 1542
rect 815 1538 819 1542
rect 911 1538 915 1542
rect 951 1538 955 1542
rect 1079 1538 1083 1542
rect 1207 1538 1211 1542
rect 1231 1538 1235 1542
rect 1335 1538 1339 1542
rect 1367 1538 1371 1542
rect 1471 1538 1475 1542
rect 1503 1538 1507 1542
rect 1631 1538 1635 1542
rect 1751 1538 1755 1542
rect 1831 1538 1835 1542
rect 1871 1542 1875 1546
rect 1967 1542 1971 1546
rect 2087 1542 2091 1546
rect 2167 1542 2171 1546
rect 2223 1542 2227 1546
rect 2255 1542 2259 1546
rect 2343 1542 2347 1546
rect 2359 1542 2363 1546
rect 2439 1542 2443 1546
rect 2495 1542 2499 1546
rect 2535 1542 2539 1546
rect 2631 1542 2635 1546
rect 2647 1542 2651 1546
rect 2767 1542 2771 1546
rect 2783 1542 2787 1546
rect 2903 1542 2907 1546
rect 2943 1542 2947 1546
rect 3047 1542 3051 1546
rect 3119 1542 3123 1546
rect 3199 1542 3203 1546
rect 3303 1542 3307 1546
rect 3359 1542 3363 1546
rect 3495 1542 3499 1546
rect 3503 1542 3507 1546
rect 3591 1542 3595 1546
rect 111 1458 115 1462
rect 135 1458 139 1462
rect 231 1458 235 1462
rect 239 1458 243 1462
rect 359 1458 363 1462
rect 375 1458 379 1462
rect 479 1458 483 1462
rect 519 1458 523 1462
rect 599 1458 603 1462
rect 663 1458 667 1462
rect 719 1458 723 1462
rect 807 1458 811 1462
rect 831 1458 835 1462
rect 935 1458 939 1462
rect 943 1458 947 1462
rect 1039 1458 1043 1462
rect 1071 1458 1075 1462
rect 1143 1458 1147 1462
rect 1199 1458 1203 1462
rect 1255 1458 1259 1462
rect 1327 1458 1331 1462
rect 1463 1458 1467 1462
rect 1831 1458 1835 1462
rect 1871 1462 1875 1466
rect 2095 1462 2099 1466
rect 2175 1462 2179 1466
rect 2263 1462 2267 1466
rect 2343 1462 2347 1466
rect 2351 1462 2355 1466
rect 2423 1462 2427 1466
rect 2447 1462 2451 1466
rect 2503 1462 2507 1466
rect 2543 1462 2547 1466
rect 2607 1462 2611 1466
rect 2655 1462 2659 1466
rect 2735 1462 2739 1466
rect 2791 1462 2795 1466
rect 2895 1462 2899 1466
rect 2951 1462 2955 1466
rect 3079 1462 3083 1466
rect 3127 1462 3131 1466
rect 3279 1462 3283 1466
rect 3311 1462 3315 1466
rect 3479 1462 3483 1466
rect 3503 1462 3507 1466
rect 3591 1462 3595 1466
rect 1871 1386 1875 1390
rect 2255 1386 2259 1390
rect 2263 1386 2267 1390
rect 2335 1386 2339 1390
rect 2343 1386 2347 1390
rect 2415 1386 2419 1390
rect 2423 1386 2427 1390
rect 2495 1386 2499 1390
rect 2503 1386 2507 1390
rect 2591 1386 2595 1390
rect 2599 1386 2603 1390
rect 2695 1386 2699 1390
rect 2727 1386 2731 1390
rect 2807 1386 2811 1390
rect 2887 1386 2891 1390
rect 2919 1386 2923 1390
rect 3039 1386 3043 1390
rect 3071 1386 3075 1390
rect 3159 1386 3163 1390
rect 3271 1386 3275 1390
rect 3279 1386 3283 1390
rect 3399 1386 3403 1390
rect 3471 1386 3475 1390
rect 3503 1386 3507 1390
rect 3591 1386 3595 1390
rect 111 1366 115 1370
rect 143 1366 147 1370
rect 239 1366 243 1370
rect 287 1366 291 1370
rect 367 1366 371 1370
rect 431 1366 435 1370
rect 487 1366 491 1370
rect 583 1366 587 1370
rect 607 1366 611 1370
rect 727 1366 731 1370
rect 735 1366 739 1370
rect 839 1366 843 1370
rect 879 1366 883 1370
rect 943 1366 947 1370
rect 1023 1366 1027 1370
rect 1047 1366 1051 1370
rect 1151 1366 1155 1370
rect 1167 1366 1171 1370
rect 1263 1366 1267 1370
rect 1319 1366 1323 1370
rect 1471 1366 1475 1370
rect 1623 1366 1627 1370
rect 1831 1366 1835 1370
rect 1871 1298 1875 1302
rect 2215 1298 2219 1302
rect 2271 1298 2275 1302
rect 2295 1298 2299 1302
rect 2351 1298 2355 1302
rect 2375 1298 2379 1302
rect 2431 1298 2435 1302
rect 2455 1298 2459 1302
rect 2511 1298 2515 1302
rect 2551 1298 2555 1302
rect 2599 1298 2603 1302
rect 2663 1298 2667 1302
rect 2703 1298 2707 1302
rect 2791 1298 2795 1302
rect 2815 1298 2819 1302
rect 2927 1298 2931 1302
rect 3047 1298 3051 1302
rect 3071 1298 3075 1302
rect 3167 1298 3171 1302
rect 3215 1298 3219 1302
rect 3287 1298 3291 1302
rect 3367 1298 3371 1302
rect 3407 1298 3411 1302
rect 3511 1298 3515 1302
rect 3591 1298 3595 1302
rect 111 1286 115 1290
rect 135 1286 139 1290
rect 263 1286 267 1290
rect 279 1286 283 1290
rect 423 1286 427 1290
rect 575 1286 579 1290
rect 591 1286 595 1290
rect 727 1286 731 1290
rect 759 1286 763 1290
rect 871 1286 875 1290
rect 927 1286 931 1290
rect 1015 1286 1019 1290
rect 1079 1286 1083 1290
rect 1159 1286 1163 1290
rect 1223 1286 1227 1290
rect 1311 1286 1315 1290
rect 1351 1286 1355 1290
rect 1463 1286 1467 1290
rect 1479 1286 1483 1290
rect 1607 1286 1611 1290
rect 1615 1286 1619 1290
rect 1735 1286 1739 1290
rect 1831 1286 1835 1290
rect 1871 1218 1875 1222
rect 2111 1218 2115 1222
rect 2207 1218 2211 1222
rect 2287 1218 2291 1222
rect 2303 1218 2307 1222
rect 2367 1218 2371 1222
rect 2407 1218 2411 1222
rect 2447 1218 2451 1222
rect 2527 1218 2531 1222
rect 2543 1218 2547 1222
rect 2647 1218 2651 1222
rect 2655 1218 2659 1222
rect 2775 1218 2779 1222
rect 2783 1218 2787 1222
rect 2911 1218 2915 1222
rect 2919 1218 2923 1222
rect 3055 1218 3059 1222
rect 3063 1218 3067 1222
rect 3199 1218 3203 1222
rect 3207 1218 3211 1222
rect 3343 1218 3347 1222
rect 3359 1218 3363 1222
rect 3495 1218 3499 1222
rect 3503 1218 3507 1222
rect 3591 1218 3595 1222
rect 111 1202 115 1206
rect 143 1202 147 1206
rect 271 1202 275 1206
rect 311 1202 315 1206
rect 431 1202 435 1206
rect 487 1202 491 1206
rect 599 1202 603 1206
rect 671 1202 675 1206
rect 767 1202 771 1206
rect 847 1202 851 1206
rect 935 1202 939 1206
rect 1007 1202 1011 1206
rect 1087 1202 1091 1206
rect 1159 1202 1163 1206
rect 1231 1202 1235 1206
rect 1295 1202 1299 1206
rect 1359 1202 1363 1206
rect 1415 1202 1419 1206
rect 1487 1202 1491 1206
rect 1535 1202 1539 1206
rect 1615 1202 1619 1206
rect 1655 1202 1659 1206
rect 1743 1202 1747 1206
rect 1751 1202 1755 1206
rect 1831 1202 1835 1206
rect 1871 1134 1875 1138
rect 1903 1134 1907 1138
rect 2119 1134 2123 1138
rect 2127 1134 2131 1138
rect 2215 1134 2219 1138
rect 2311 1134 2315 1138
rect 2359 1134 2363 1138
rect 2415 1134 2419 1138
rect 2535 1134 2539 1138
rect 2575 1134 2579 1138
rect 2655 1134 2659 1138
rect 2775 1134 2779 1138
rect 2783 1134 2787 1138
rect 2919 1134 2923 1138
rect 2967 1134 2971 1138
rect 3063 1134 3067 1138
rect 3159 1134 3163 1138
rect 3207 1134 3211 1138
rect 3343 1134 3347 1138
rect 3351 1134 3355 1138
rect 3503 1134 3507 1138
rect 3511 1134 3515 1138
rect 3591 1134 3595 1138
rect 111 1126 115 1130
rect 135 1126 139 1130
rect 247 1126 251 1130
rect 303 1126 307 1130
rect 383 1126 387 1130
rect 479 1126 483 1130
rect 519 1126 523 1130
rect 647 1126 651 1130
rect 663 1126 667 1130
rect 775 1126 779 1130
rect 839 1126 843 1130
rect 895 1126 899 1130
rect 999 1126 1003 1130
rect 1015 1126 1019 1130
rect 1135 1126 1139 1130
rect 1151 1126 1155 1130
rect 1255 1126 1259 1130
rect 1287 1126 1291 1130
rect 1375 1126 1379 1130
rect 1407 1126 1411 1130
rect 1503 1126 1507 1130
rect 1527 1126 1531 1130
rect 1631 1126 1635 1130
rect 1647 1126 1651 1130
rect 1743 1126 1747 1130
rect 1831 1126 1835 1130
rect 1871 1058 1875 1062
rect 1895 1058 1899 1062
rect 2015 1058 2019 1062
rect 2119 1058 2123 1062
rect 2167 1058 2171 1062
rect 2327 1058 2331 1062
rect 2351 1058 2355 1062
rect 2487 1058 2491 1062
rect 2567 1058 2571 1062
rect 2639 1058 2643 1062
rect 2767 1058 2771 1062
rect 2791 1058 2795 1062
rect 2935 1058 2939 1062
rect 2959 1058 2963 1062
rect 3079 1058 3083 1062
rect 3151 1058 3155 1062
rect 3223 1058 3227 1062
rect 3335 1058 3339 1062
rect 3375 1058 3379 1062
rect 3503 1058 3507 1062
rect 3591 1058 3595 1062
rect 111 1038 115 1042
rect 143 1038 147 1042
rect 239 1038 243 1042
rect 255 1038 259 1042
rect 359 1038 363 1042
rect 391 1038 395 1042
rect 471 1038 475 1042
rect 527 1038 531 1042
rect 575 1038 579 1042
rect 655 1038 659 1042
rect 671 1038 675 1042
rect 767 1038 771 1042
rect 783 1038 787 1042
rect 855 1038 859 1042
rect 903 1038 907 1042
rect 943 1038 947 1042
rect 1023 1038 1027 1042
rect 1031 1038 1035 1042
rect 1127 1038 1131 1042
rect 1143 1038 1147 1042
rect 1223 1038 1227 1042
rect 1263 1038 1267 1042
rect 1383 1038 1387 1042
rect 1511 1038 1515 1042
rect 1639 1038 1643 1042
rect 1751 1038 1755 1042
rect 1831 1038 1835 1042
rect 1871 978 1875 982
rect 1903 978 1907 982
rect 1983 978 1987 982
rect 2023 978 2027 982
rect 2079 978 2083 982
rect 2175 978 2179 982
rect 2199 978 2203 982
rect 2335 978 2339 982
rect 2479 978 2483 982
rect 2495 978 2499 982
rect 2631 978 2635 982
rect 2647 978 2651 982
rect 2791 978 2795 982
rect 2799 978 2803 982
rect 2943 978 2947 982
rect 2967 978 2971 982
rect 3087 978 3091 982
rect 3151 978 3155 982
rect 3231 978 3235 982
rect 3343 978 3347 982
rect 3383 978 3387 982
rect 3511 978 3515 982
rect 3591 978 3595 982
rect 111 950 115 954
rect 135 950 139 954
rect 231 950 235 954
rect 263 950 267 954
rect 351 950 355 954
rect 415 950 419 954
rect 463 950 467 954
rect 559 950 563 954
rect 567 950 571 954
rect 663 950 667 954
rect 703 950 707 954
rect 759 950 763 954
rect 839 950 843 954
rect 847 950 851 954
rect 935 950 939 954
rect 975 950 979 954
rect 1023 950 1027 954
rect 1103 950 1107 954
rect 1119 950 1123 954
rect 1215 950 1219 954
rect 1223 950 1227 954
rect 1335 950 1339 954
rect 1439 950 1443 954
rect 1543 950 1547 954
rect 1655 950 1659 954
rect 1743 950 1747 954
rect 1831 950 1835 954
rect 1871 890 1875 894
rect 1895 890 1899 894
rect 1919 890 1923 894
rect 1975 890 1979 894
rect 2071 890 2075 894
rect 2095 890 2099 894
rect 2191 890 2195 894
rect 2271 890 2275 894
rect 2327 890 2331 894
rect 2455 890 2459 894
rect 2471 890 2475 894
rect 2623 890 2627 894
rect 2655 890 2659 894
rect 2783 890 2787 894
rect 2863 890 2867 894
rect 2959 890 2963 894
rect 3079 890 3083 894
rect 3143 890 3147 894
rect 3303 890 3307 894
rect 3335 890 3339 894
rect 3503 890 3507 894
rect 3591 890 3595 894
rect 111 870 115 874
rect 143 870 147 874
rect 247 870 251 874
rect 271 870 275 874
rect 383 870 387 874
rect 423 870 427 874
rect 519 870 523 874
rect 567 870 571 874
rect 663 870 667 874
rect 711 870 715 874
rect 815 870 819 874
rect 847 870 851 874
rect 959 870 963 874
rect 983 870 987 874
rect 1103 870 1107 874
rect 1111 870 1115 874
rect 1231 870 1235 874
rect 1247 870 1251 874
rect 1343 870 1347 874
rect 1383 870 1387 874
rect 1447 870 1451 874
rect 1511 870 1515 874
rect 1551 870 1555 874
rect 1639 870 1643 874
rect 1663 870 1667 874
rect 1751 870 1755 874
rect 1831 870 1835 874
rect 1871 814 1875 818
rect 1903 814 1907 818
rect 1927 814 1931 818
rect 2015 814 2019 818
rect 2103 814 2107 818
rect 2167 814 2171 818
rect 2279 814 2283 818
rect 2327 814 2331 818
rect 2463 814 2467 818
rect 2487 814 2491 818
rect 2647 814 2651 818
rect 2663 814 2667 818
rect 2807 814 2811 818
rect 2871 814 2875 818
rect 2959 814 2963 818
rect 3087 814 3091 818
rect 3103 814 3107 818
rect 3247 814 3251 818
rect 3311 814 3315 818
rect 3391 814 3395 818
rect 3511 814 3515 818
rect 3591 814 3595 818
rect 111 782 115 786
rect 135 782 139 786
rect 215 782 219 786
rect 239 782 243 786
rect 303 782 307 786
rect 375 782 379 786
rect 415 782 419 786
rect 511 782 515 786
rect 543 782 547 786
rect 655 782 659 786
rect 687 782 691 786
rect 807 782 811 786
rect 839 782 843 786
rect 951 782 955 786
rect 991 782 995 786
rect 1095 782 1099 786
rect 1143 782 1147 786
rect 1239 782 1243 786
rect 1295 782 1299 786
rect 1375 782 1379 786
rect 1447 782 1451 786
rect 1503 782 1507 786
rect 1607 782 1611 786
rect 1631 782 1635 786
rect 1743 782 1747 786
rect 1831 782 1835 786
rect 1871 738 1875 742
rect 1895 738 1899 742
rect 1967 738 1971 742
rect 2007 738 2011 742
rect 2063 738 2067 742
rect 2159 738 2163 742
rect 2175 738 2179 742
rect 2303 738 2307 742
rect 2319 738 2323 742
rect 2447 738 2451 742
rect 2479 738 2483 742
rect 2599 738 2603 742
rect 2639 738 2643 742
rect 2751 738 2755 742
rect 2799 738 2803 742
rect 2903 738 2907 742
rect 2951 738 2955 742
rect 3055 738 3059 742
rect 3095 738 3099 742
rect 3207 738 3211 742
rect 3239 738 3243 742
rect 3359 738 3363 742
rect 3383 738 3387 742
rect 3503 738 3507 742
rect 3591 738 3595 742
rect 111 698 115 702
rect 143 698 147 702
rect 223 698 227 702
rect 231 698 235 702
rect 311 698 315 702
rect 319 698 323 702
rect 423 698 427 702
rect 543 698 547 702
rect 551 698 555 702
rect 679 698 683 702
rect 695 698 699 702
rect 815 698 819 702
rect 847 698 851 702
rect 951 698 955 702
rect 999 698 1003 702
rect 1087 698 1091 702
rect 1151 698 1155 702
rect 1215 698 1219 702
rect 1303 698 1307 702
rect 1335 698 1339 702
rect 1455 698 1459 702
rect 1583 698 1587 702
rect 1615 698 1619 702
rect 1831 698 1835 702
rect 1871 662 1875 666
rect 1975 662 1979 666
rect 2071 662 2075 666
rect 2175 662 2179 666
rect 2183 662 2187 666
rect 2271 662 2275 666
rect 2311 662 2315 666
rect 2375 662 2379 666
rect 2455 662 2459 666
rect 2487 662 2491 666
rect 2607 662 2611 666
rect 2735 662 2739 666
rect 2759 662 2763 666
rect 2863 662 2867 666
rect 2911 662 2915 666
rect 2991 662 2995 666
rect 3063 662 3067 666
rect 3119 662 3123 666
rect 3215 662 3219 666
rect 3247 662 3251 666
rect 3367 662 3371 666
rect 3375 662 3379 666
rect 3511 662 3515 666
rect 3591 662 3595 666
rect 111 614 115 618
rect 223 614 227 618
rect 311 614 315 618
rect 415 614 419 618
rect 447 614 451 618
rect 527 614 531 618
rect 535 614 539 618
rect 607 614 611 618
rect 671 614 675 618
rect 687 614 691 618
rect 775 614 779 618
rect 807 614 811 618
rect 871 614 875 618
rect 943 614 947 618
rect 959 614 963 618
rect 1047 614 1051 618
rect 1079 614 1083 618
rect 1143 614 1147 618
rect 1207 614 1211 618
rect 1239 614 1243 618
rect 1327 614 1331 618
rect 1335 614 1339 618
rect 1431 614 1435 618
rect 1447 614 1451 618
rect 1575 614 1579 618
rect 1831 614 1835 618
rect 1871 586 1875 590
rect 2167 586 2171 590
rect 2263 586 2267 590
rect 2343 586 2347 590
rect 2367 586 2371 590
rect 2423 586 2427 590
rect 2479 586 2483 590
rect 2503 586 2507 590
rect 2591 586 2595 590
rect 2599 586 2603 590
rect 2695 586 2699 590
rect 2727 586 2731 590
rect 2815 586 2819 590
rect 2855 586 2859 590
rect 2959 586 2963 590
rect 2983 586 2987 590
rect 3111 586 3115 590
rect 3239 586 3243 590
rect 3279 586 3283 590
rect 3367 586 3371 590
rect 3447 586 3451 590
rect 3503 586 3507 590
rect 3591 586 3595 590
rect 111 526 115 530
rect 335 526 339 530
rect 423 526 427 530
rect 455 526 459 530
rect 511 526 515 530
rect 535 526 539 530
rect 591 526 595 530
rect 615 526 619 530
rect 671 526 675 530
rect 695 526 699 530
rect 751 526 755 530
rect 783 526 787 530
rect 839 526 843 530
rect 879 526 883 530
rect 927 526 931 530
rect 967 526 971 530
rect 1015 526 1019 530
rect 1055 526 1059 530
rect 1103 526 1107 530
rect 1151 526 1155 530
rect 1191 526 1195 530
rect 1247 526 1251 530
rect 1279 526 1283 530
rect 1343 526 1347 530
rect 1439 526 1443 530
rect 1831 526 1835 530
rect 1871 502 1875 506
rect 2191 502 2195 506
rect 2271 502 2275 506
rect 2287 502 2291 506
rect 2351 502 2355 506
rect 2383 502 2387 506
rect 2431 502 2435 506
rect 2487 502 2491 506
rect 2511 502 2515 506
rect 2583 502 2587 506
rect 2599 502 2603 506
rect 2687 502 2691 506
rect 2703 502 2707 506
rect 2791 502 2795 506
rect 2823 502 2827 506
rect 2911 502 2915 506
rect 2967 502 2971 506
rect 3039 502 3043 506
rect 3119 502 3123 506
rect 3175 502 3179 506
rect 3287 502 3291 506
rect 3319 502 3323 506
rect 3455 502 3459 506
rect 3471 502 3475 506
rect 3591 502 3595 506
rect 111 442 115 446
rect 223 442 227 446
rect 327 442 331 446
rect 335 442 339 446
rect 415 442 419 446
rect 447 442 451 446
rect 503 442 507 446
rect 559 442 563 446
rect 583 442 587 446
rect 663 442 667 446
rect 743 442 747 446
rect 759 442 763 446
rect 831 442 835 446
rect 847 442 851 446
rect 919 442 923 446
rect 935 442 939 446
rect 1007 442 1011 446
rect 1023 442 1027 446
rect 1095 442 1099 446
rect 1111 442 1115 446
rect 1183 442 1187 446
rect 1199 442 1203 446
rect 1271 442 1275 446
rect 1295 442 1299 446
rect 1831 442 1835 446
rect 1871 422 1875 426
rect 1975 422 1979 426
rect 2063 422 2067 426
rect 2159 422 2163 426
rect 2183 422 2187 426
rect 2255 422 2259 426
rect 2279 422 2283 426
rect 2359 422 2363 426
rect 2375 422 2379 426
rect 2471 422 2475 426
rect 2479 422 2483 426
rect 2575 422 2579 426
rect 2607 422 2611 426
rect 2679 422 2683 426
rect 2759 422 2763 426
rect 2783 422 2787 426
rect 2903 422 2907 426
rect 2927 422 2931 426
rect 3031 422 3035 426
rect 3111 422 3115 426
rect 3167 422 3171 426
rect 3303 422 3307 426
rect 3311 422 3315 426
rect 3463 422 3467 426
rect 3495 422 3499 426
rect 3591 422 3595 426
rect 111 354 115 358
rect 143 354 147 358
rect 231 354 235 358
rect 263 354 267 358
rect 343 354 347 358
rect 399 354 403 358
rect 455 354 459 358
rect 535 354 539 358
rect 567 354 571 358
rect 671 354 675 358
rect 767 354 771 358
rect 791 354 795 358
rect 855 354 859 358
rect 911 354 915 358
rect 943 354 947 358
rect 1023 354 1027 358
rect 1031 354 1035 358
rect 1119 354 1123 358
rect 1127 354 1131 358
rect 1207 354 1211 358
rect 1231 354 1235 358
rect 1303 354 1307 358
rect 1335 354 1339 358
rect 1439 354 1443 358
rect 1831 354 1835 358
rect 1871 342 1875 346
rect 1983 342 1987 346
rect 2071 342 2075 346
rect 2167 342 2171 346
rect 2215 342 2219 346
rect 2263 342 2267 346
rect 2295 342 2299 346
rect 2367 342 2371 346
rect 2383 342 2387 346
rect 2479 342 2483 346
rect 2591 342 2595 346
rect 2615 342 2619 346
rect 2719 342 2723 346
rect 2767 342 2771 346
rect 2847 342 2851 346
rect 2935 342 2939 346
rect 2983 342 2987 346
rect 3119 342 3123 346
rect 3255 342 3259 346
rect 3311 342 3315 346
rect 3391 342 3395 346
rect 3503 342 3507 346
rect 3511 342 3515 346
rect 3591 342 3595 346
rect 111 270 115 274
rect 135 270 139 274
rect 247 270 251 274
rect 255 270 259 274
rect 391 270 395 274
rect 527 270 531 274
rect 543 270 547 274
rect 663 270 667 274
rect 695 270 699 274
rect 783 270 787 274
rect 847 270 851 274
rect 903 270 907 274
rect 991 270 995 274
rect 1015 270 1019 274
rect 1119 270 1123 274
rect 1223 270 1227 274
rect 1239 270 1243 274
rect 1327 270 1331 274
rect 1359 270 1363 274
rect 1431 270 1435 274
rect 1479 270 1483 274
rect 1599 270 1603 274
rect 1831 270 1835 274
rect 1871 262 1875 266
rect 1991 262 1995 266
rect 2119 262 2123 266
rect 2207 262 2211 266
rect 2255 262 2259 266
rect 2287 262 2291 266
rect 2375 262 2379 266
rect 2391 262 2395 266
rect 2471 262 2475 266
rect 2535 262 2539 266
rect 2583 262 2587 266
rect 2679 262 2683 266
rect 2711 262 2715 266
rect 2815 262 2819 266
rect 2839 262 2843 266
rect 2951 262 2955 266
rect 2975 262 2979 266
rect 3095 262 3099 266
rect 3111 262 3115 266
rect 3239 262 3243 266
rect 3247 262 3251 266
rect 3383 262 3387 266
rect 3503 262 3507 266
rect 3591 262 3595 266
rect 1871 174 1875 178
rect 1903 174 1907 178
rect 1983 174 1987 178
rect 1999 174 2003 178
rect 2087 174 2091 178
rect 2127 174 2131 178
rect 2215 174 2219 178
rect 2263 174 2267 178
rect 2351 174 2355 178
rect 2399 174 2403 178
rect 2487 174 2491 178
rect 2543 174 2547 178
rect 2623 174 2627 178
rect 2687 174 2691 178
rect 2743 174 2747 178
rect 2823 174 2827 178
rect 2855 174 2859 178
rect 2959 174 2963 178
rect 3063 174 3067 178
rect 3103 174 3107 178
rect 3159 174 3163 178
rect 3247 174 3251 178
rect 3343 174 3347 178
rect 3391 174 3395 178
rect 3431 174 3435 178
rect 3511 174 3515 178
rect 3591 174 3595 178
rect 111 158 115 162
rect 143 158 147 162
rect 223 158 227 162
rect 255 158 259 162
rect 303 158 307 162
rect 383 158 387 162
rect 399 158 403 162
rect 463 158 467 162
rect 543 158 547 162
rect 551 158 555 162
rect 623 158 627 162
rect 703 158 707 162
rect 783 158 787 162
rect 855 158 859 162
rect 863 158 867 162
rect 943 158 947 162
rect 999 158 1003 162
rect 1023 158 1027 162
rect 1103 158 1107 162
rect 1127 158 1131 162
rect 1183 158 1187 162
rect 1247 158 1251 162
rect 1263 158 1267 162
rect 1343 158 1347 162
rect 1367 158 1371 162
rect 1423 158 1427 162
rect 1487 158 1491 162
rect 1511 158 1515 162
rect 1591 158 1595 162
rect 1607 158 1611 162
rect 1671 158 1675 162
rect 1751 158 1755 162
rect 1831 158 1835 162
rect 1871 98 1875 102
rect 1895 98 1899 102
rect 1975 98 1979 102
rect 2079 98 2083 102
rect 2207 98 2211 102
rect 2343 98 2347 102
rect 2479 98 2483 102
rect 2615 98 2619 102
rect 2735 98 2739 102
rect 2847 98 2851 102
rect 2951 98 2955 102
rect 3055 98 3059 102
rect 3151 98 3155 102
rect 3239 98 3243 102
rect 3335 98 3339 102
rect 3423 98 3427 102
rect 3503 98 3507 102
rect 3591 98 3595 102
rect 111 82 115 86
rect 135 82 139 86
rect 215 82 219 86
rect 295 82 299 86
rect 375 82 379 86
rect 455 82 459 86
rect 535 82 539 86
rect 615 82 619 86
rect 695 82 699 86
rect 775 82 779 86
rect 855 82 859 86
rect 935 82 939 86
rect 1015 82 1019 86
rect 1095 82 1099 86
rect 1175 82 1179 86
rect 1255 82 1259 86
rect 1335 82 1339 86
rect 1415 82 1419 86
rect 1503 82 1507 86
rect 1583 82 1587 86
rect 1663 82 1667 86
rect 1743 82 1747 86
rect 1831 82 1835 86
<< m4 >>
rect 84 3665 85 3671
rect 91 3670 1843 3671
rect 91 3666 111 3670
rect 115 3666 135 3670
rect 139 3666 215 3670
rect 219 3666 295 3670
rect 299 3666 1831 3670
rect 1835 3666 1843 3670
rect 91 3665 1843 3666
rect 1849 3665 1850 3671
rect 1854 3597 1855 3603
rect 1861 3602 3631 3603
rect 1861 3598 1871 3602
rect 1875 3598 2063 3602
rect 2067 3598 2151 3602
rect 2155 3598 2255 3602
rect 2259 3598 2367 3602
rect 2371 3598 2479 3602
rect 2483 3598 2591 3602
rect 2595 3598 2703 3602
rect 2707 3598 2815 3602
rect 2819 3598 2919 3602
rect 2923 3598 3015 3602
rect 3019 3598 3111 3602
rect 3115 3598 3207 3602
rect 3211 3598 3303 3602
rect 3307 3598 3399 3602
rect 3403 3598 3591 3602
rect 3595 3598 3631 3602
rect 1861 3597 3631 3598
rect 3637 3597 3638 3603
rect 1854 3595 1862 3597
rect 96 3589 97 3595
rect 103 3594 1855 3595
rect 103 3590 111 3594
rect 115 3590 143 3594
rect 147 3590 223 3594
rect 227 3590 303 3594
rect 307 3590 343 3594
rect 347 3590 471 3594
rect 475 3590 607 3594
rect 611 3590 743 3594
rect 747 3590 879 3594
rect 883 3590 999 3594
rect 1003 3590 1111 3594
rect 1115 3590 1223 3594
rect 1227 3590 1327 3594
rect 1331 3590 1423 3594
rect 1427 3590 1527 3594
rect 1531 3590 1631 3594
rect 1635 3590 1831 3594
rect 1835 3590 1855 3594
rect 103 3589 1855 3590
rect 1861 3589 1862 3595
rect 1842 3521 1843 3527
rect 1849 3526 3619 3527
rect 1849 3522 1871 3526
rect 1875 3522 2055 3526
rect 2059 3522 2087 3526
rect 2091 3522 2143 3526
rect 2147 3522 2167 3526
rect 2171 3522 2247 3526
rect 2251 3522 2263 3526
rect 2267 3522 2359 3526
rect 2363 3522 2367 3526
rect 2371 3522 2471 3526
rect 2475 3522 2487 3526
rect 2491 3522 2583 3526
rect 2587 3522 2615 3526
rect 2619 3522 2695 3526
rect 2699 3522 2743 3526
rect 2747 3522 2807 3526
rect 2811 3522 2871 3526
rect 2875 3522 2911 3526
rect 2915 3522 2991 3526
rect 2995 3522 3007 3526
rect 3011 3522 3103 3526
rect 3107 3522 3119 3526
rect 3123 3522 3199 3526
rect 3203 3522 3247 3526
rect 3251 3522 3295 3526
rect 3299 3522 3375 3526
rect 3379 3522 3391 3526
rect 3395 3522 3591 3526
rect 3595 3522 3619 3526
rect 1849 3521 3619 3522
rect 3625 3521 3626 3527
rect 1842 3519 1850 3521
rect 84 3513 85 3519
rect 91 3518 1843 3519
rect 91 3514 111 3518
rect 115 3514 135 3518
rect 139 3514 191 3518
rect 195 3514 215 3518
rect 219 3514 327 3518
rect 331 3514 335 3518
rect 339 3514 463 3518
rect 467 3514 471 3518
rect 475 3514 599 3518
rect 603 3514 623 3518
rect 627 3514 735 3518
rect 739 3514 775 3518
rect 779 3514 871 3518
rect 875 3514 919 3518
rect 923 3514 991 3518
rect 995 3514 1055 3518
rect 1059 3514 1103 3518
rect 1107 3514 1183 3518
rect 1187 3514 1215 3518
rect 1219 3514 1311 3518
rect 1315 3514 1319 3518
rect 1323 3514 1415 3518
rect 1419 3514 1439 3518
rect 1443 3514 1519 3518
rect 1523 3514 1567 3518
rect 1571 3514 1623 3518
rect 1627 3514 1831 3518
rect 1835 3514 1843 3518
rect 91 3513 1843 3514
rect 1849 3513 1850 3519
rect 96 3437 97 3443
rect 103 3442 1855 3443
rect 103 3438 111 3442
rect 115 3438 151 3442
rect 155 3438 199 3442
rect 203 3438 295 3442
rect 299 3438 335 3442
rect 339 3438 455 3442
rect 459 3438 479 3442
rect 483 3438 623 3442
rect 627 3438 631 3442
rect 635 3438 783 3442
rect 787 3438 791 3442
rect 795 3438 927 3442
rect 931 3438 959 3442
rect 963 3438 1063 3442
rect 1067 3438 1119 3442
rect 1123 3438 1191 3442
rect 1195 3438 1271 3442
rect 1275 3438 1319 3442
rect 1323 3438 1415 3442
rect 1419 3438 1447 3442
rect 1451 3438 1559 3442
rect 1563 3438 1575 3442
rect 1579 3438 1711 3442
rect 1715 3438 1831 3442
rect 1835 3438 1855 3442
rect 103 3437 1855 3438
rect 1861 3442 3638 3443
rect 1861 3438 1871 3442
rect 1875 3438 2095 3442
rect 2099 3438 2111 3442
rect 2115 3438 2175 3442
rect 2179 3438 2199 3442
rect 2203 3438 2271 3442
rect 2275 3438 2303 3442
rect 2307 3438 2375 3442
rect 2379 3438 2415 3442
rect 2419 3438 2495 3442
rect 2499 3438 2543 3442
rect 2547 3438 2623 3442
rect 2627 3438 2679 3442
rect 2683 3438 2751 3442
rect 2755 3438 2815 3442
rect 2819 3438 2879 3442
rect 2883 3438 2959 3442
rect 2963 3438 2999 3442
rect 3003 3438 3111 3442
rect 3115 3438 3127 3442
rect 3131 3438 3255 3442
rect 3259 3438 3263 3442
rect 3267 3438 3383 3442
rect 3387 3438 3423 3442
rect 3427 3438 3591 3442
rect 3595 3438 3638 3442
rect 1861 3437 3638 3438
rect 84 3361 85 3367
rect 91 3366 1843 3367
rect 91 3362 111 3366
rect 115 3362 143 3366
rect 147 3362 207 3366
rect 211 3362 287 3366
rect 291 3362 335 3366
rect 339 3362 447 3366
rect 451 3362 471 3366
rect 475 3362 615 3366
rect 619 3362 623 3366
rect 627 3362 783 3366
rect 787 3362 943 3366
rect 947 3362 951 3366
rect 955 3362 1103 3366
rect 1107 3362 1111 3366
rect 1115 3362 1263 3366
rect 1267 3362 1407 3366
rect 1411 3362 1423 3366
rect 1427 3362 1551 3366
rect 1555 3362 1583 3366
rect 1587 3362 1703 3366
rect 1707 3362 1743 3366
rect 1747 3362 1831 3366
rect 1835 3362 1843 3366
rect 91 3361 1843 3362
rect 1849 3363 1850 3367
rect 1849 3362 3626 3363
rect 1849 3361 1871 3362
rect 1842 3358 1871 3361
rect 1875 3358 2103 3362
rect 2107 3358 2127 3362
rect 2131 3358 2191 3362
rect 2195 3358 2223 3362
rect 2227 3358 2295 3362
rect 2299 3358 2335 3362
rect 2339 3358 2407 3362
rect 2411 3358 2455 3362
rect 2459 3358 2535 3362
rect 2539 3358 2583 3362
rect 2587 3358 2671 3362
rect 2675 3358 2719 3362
rect 2723 3358 2807 3362
rect 2811 3358 2863 3362
rect 2867 3358 2951 3362
rect 2955 3358 3007 3362
rect 3011 3358 3103 3362
rect 3107 3358 3159 3362
rect 3163 3358 3255 3362
rect 3259 3358 3311 3362
rect 3315 3358 3415 3362
rect 3419 3358 3471 3362
rect 3475 3358 3591 3362
rect 3595 3358 3626 3362
rect 1842 3357 3626 3358
rect 96 3281 97 3287
rect 103 3286 1855 3287
rect 103 3282 111 3286
rect 115 3282 215 3286
rect 219 3282 343 3286
rect 347 3282 351 3286
rect 355 3282 455 3286
rect 459 3282 479 3286
rect 483 3282 575 3286
rect 579 3282 631 3286
rect 635 3282 703 3286
rect 707 3282 791 3286
rect 795 3282 839 3286
rect 843 3282 951 3286
rect 955 3282 983 3286
rect 987 3282 1111 3286
rect 1115 3282 1119 3286
rect 1123 3282 1255 3286
rect 1259 3282 1271 3286
rect 1275 3282 1383 3286
rect 1387 3282 1431 3286
rect 1435 3282 1511 3286
rect 1515 3282 1591 3286
rect 1595 3282 1639 3286
rect 1643 3282 1751 3286
rect 1755 3282 1831 3286
rect 1835 3282 1855 3286
rect 103 3281 1855 3282
rect 1861 3281 1862 3287
rect 1854 3269 1855 3275
rect 1861 3274 3631 3275
rect 1861 3270 1871 3274
rect 1875 3270 2135 3274
rect 2139 3270 2231 3274
rect 2235 3270 2279 3274
rect 2283 3270 2343 3274
rect 2347 3270 2415 3274
rect 2419 3270 2463 3274
rect 2467 3270 2551 3274
rect 2555 3270 2591 3274
rect 2595 3270 2687 3274
rect 2691 3270 2727 3274
rect 2731 3270 2823 3274
rect 2827 3270 2871 3274
rect 2875 3270 2959 3274
rect 2963 3270 3015 3274
rect 3019 3270 3095 3274
rect 3099 3270 3167 3274
rect 3171 3270 3231 3274
rect 3235 3270 3319 3274
rect 3323 3270 3375 3274
rect 3379 3270 3479 3274
rect 3483 3270 3511 3274
rect 3515 3270 3591 3274
rect 3595 3270 3631 3274
rect 1861 3269 3631 3270
rect 3637 3269 3638 3275
rect 84 3205 85 3211
rect 91 3210 1843 3211
rect 91 3206 111 3210
rect 115 3206 343 3210
rect 347 3206 447 3210
rect 451 3206 487 3210
rect 491 3206 567 3210
rect 571 3206 575 3210
rect 579 3206 663 3210
rect 667 3206 695 3210
rect 699 3206 767 3210
rect 771 3206 831 3210
rect 835 3206 887 3210
rect 891 3206 975 3210
rect 979 3206 1023 3210
rect 1027 3206 1111 3210
rect 1115 3206 1191 3210
rect 1195 3206 1247 3210
rect 1251 3206 1375 3210
rect 1379 3206 1503 3210
rect 1507 3206 1567 3210
rect 1571 3206 1631 3210
rect 1635 3206 1743 3210
rect 1747 3206 1831 3210
rect 1835 3206 1843 3210
rect 91 3205 1843 3206
rect 1849 3205 1850 3211
rect 1842 3189 1843 3195
rect 1849 3194 3619 3195
rect 1849 3190 1871 3194
rect 1875 3190 1895 3194
rect 1899 3190 1991 3194
rect 1995 3190 2119 3194
rect 2123 3190 2127 3194
rect 2131 3190 2247 3194
rect 2251 3190 2271 3194
rect 2275 3190 2383 3194
rect 2387 3190 2407 3194
rect 2411 3190 2511 3194
rect 2515 3190 2543 3194
rect 2547 3190 2639 3194
rect 2643 3190 2679 3194
rect 2683 3190 2767 3194
rect 2771 3190 2815 3194
rect 2819 3190 2895 3194
rect 2899 3190 2951 3194
rect 2955 3190 3031 3194
rect 3035 3190 3087 3194
rect 3091 3190 3175 3194
rect 3179 3190 3223 3194
rect 3227 3190 3327 3194
rect 3331 3190 3367 3194
rect 3371 3190 3487 3194
rect 3491 3190 3503 3194
rect 3507 3190 3591 3194
rect 3595 3190 3619 3194
rect 1849 3189 3619 3190
rect 3625 3189 3626 3195
rect 96 3125 97 3131
rect 103 3130 1855 3131
rect 103 3126 111 3130
rect 115 3126 495 3130
rect 499 3126 583 3130
rect 587 3126 591 3130
rect 595 3126 671 3130
rect 675 3126 759 3130
rect 763 3126 775 3130
rect 779 3126 847 3130
rect 851 3126 895 3130
rect 899 3126 935 3130
rect 939 3126 1023 3130
rect 1027 3126 1031 3130
rect 1035 3126 1111 3130
rect 1115 3126 1199 3130
rect 1203 3126 1287 3130
rect 1291 3126 1375 3130
rect 1379 3126 1383 3130
rect 1387 3126 1575 3130
rect 1579 3126 1751 3130
rect 1755 3126 1831 3130
rect 1835 3126 1855 3130
rect 103 3125 1855 3126
rect 1861 3125 1862 3131
rect 1854 3097 1855 3103
rect 1861 3102 3631 3103
rect 1861 3098 1871 3102
rect 1875 3098 1903 3102
rect 1907 3098 1999 3102
rect 2003 3098 2015 3102
rect 2019 3098 2127 3102
rect 2131 3098 2191 3102
rect 2195 3098 2255 3102
rect 2259 3098 2391 3102
rect 2395 3098 2407 3102
rect 2411 3098 2519 3102
rect 2523 3098 2647 3102
rect 2651 3098 2655 3102
rect 2659 3098 2775 3102
rect 2779 3098 2903 3102
rect 2907 3098 2935 3102
rect 2939 3098 3039 3102
rect 3043 3098 3183 3102
rect 3187 3098 3231 3102
rect 3235 3098 3335 3102
rect 3339 3098 3495 3102
rect 3499 3098 3511 3102
rect 3515 3098 3591 3102
rect 3595 3098 3631 3102
rect 1861 3097 3631 3098
rect 3637 3097 3638 3103
rect 84 3045 85 3051
rect 91 3050 1843 3051
rect 91 3046 111 3050
rect 115 3046 543 3050
rect 547 3046 583 3050
rect 587 3046 623 3050
rect 627 3046 663 3050
rect 667 3046 711 3050
rect 715 3046 751 3050
rect 755 3046 807 3050
rect 811 3046 839 3050
rect 843 3046 903 3050
rect 907 3046 927 3050
rect 931 3046 999 3050
rect 1003 3046 1015 3050
rect 1019 3046 1087 3050
rect 1091 3046 1103 3050
rect 1107 3046 1183 3050
rect 1187 3046 1191 3050
rect 1195 3046 1279 3050
rect 1283 3046 1367 3050
rect 1371 3046 1375 3050
rect 1379 3046 1471 3050
rect 1475 3046 1831 3050
rect 1835 3046 1843 3050
rect 91 3045 1843 3046
rect 1849 3045 1850 3051
rect 1842 3013 1843 3019
rect 1849 3018 3619 3019
rect 1849 3014 1871 3018
rect 1875 3014 1895 3018
rect 1899 3014 2007 3018
rect 2011 3014 2047 3018
rect 2051 3014 2183 3018
rect 2187 3014 2223 3018
rect 2227 3014 2391 3018
rect 2395 3014 2399 3018
rect 2403 3014 2543 3018
rect 2547 3014 2647 3018
rect 2651 3014 2687 3018
rect 2691 3014 2815 3018
rect 2819 3014 2927 3018
rect 2931 3014 3039 3018
rect 3043 3014 3143 3018
rect 3147 3014 3223 3018
rect 3227 3014 3239 3018
rect 3243 3014 3335 3018
rect 3339 3014 3423 3018
rect 3427 3014 3503 3018
rect 3507 3014 3591 3018
rect 3595 3014 3619 3018
rect 1849 3013 3619 3014
rect 3625 3013 3626 3019
rect 96 2969 97 2975
rect 103 2974 1855 2975
rect 103 2970 111 2974
rect 115 2970 471 2974
rect 475 2970 551 2974
rect 555 2970 575 2974
rect 579 2970 631 2974
rect 635 2970 687 2974
rect 691 2970 719 2974
rect 723 2970 807 2974
rect 811 2970 815 2974
rect 819 2970 911 2974
rect 915 2970 943 2974
rect 947 2970 1007 2974
rect 1011 2970 1087 2974
rect 1091 2970 1095 2974
rect 1099 2970 1191 2974
rect 1195 2970 1247 2974
rect 1251 2970 1287 2974
rect 1291 2970 1383 2974
rect 1387 2970 1415 2974
rect 1419 2970 1479 2974
rect 1483 2970 1591 2974
rect 1595 2970 1751 2974
rect 1755 2970 1831 2974
rect 1835 2970 1855 2974
rect 103 2969 1855 2970
rect 1861 2969 1862 2975
rect 1854 2937 1855 2943
rect 1861 2942 3631 2943
rect 1861 2938 1871 2942
rect 1875 2938 1903 2942
rect 1907 2938 2055 2942
rect 2059 2938 2087 2942
rect 2091 2938 2231 2942
rect 2235 2938 2295 2942
rect 2299 2938 2399 2942
rect 2403 2938 2487 2942
rect 2491 2938 2551 2942
rect 2555 2938 2671 2942
rect 2675 2938 2695 2942
rect 2699 2938 2823 2942
rect 2827 2938 2839 2942
rect 2843 2938 2935 2942
rect 2939 2938 2999 2942
rect 3003 2938 3047 2942
rect 3051 2938 3151 2942
rect 3155 2938 3247 2942
rect 3251 2938 3303 2942
rect 3307 2938 3343 2942
rect 3347 2938 3431 2942
rect 3435 2938 3455 2942
rect 3459 2938 3511 2942
rect 3515 2938 3591 2942
rect 3595 2938 3631 2942
rect 1861 2937 3631 2938
rect 3637 2937 3638 2943
rect 84 2893 85 2899
rect 91 2898 1843 2899
rect 91 2894 111 2898
rect 115 2894 311 2898
rect 315 2894 431 2898
rect 435 2894 463 2898
rect 467 2894 551 2898
rect 555 2894 567 2898
rect 571 2894 679 2898
rect 683 2894 799 2898
rect 803 2894 815 2898
rect 819 2894 935 2898
rect 939 2894 951 2898
rect 955 2894 1079 2898
rect 1083 2894 1087 2898
rect 1091 2894 1223 2898
rect 1227 2894 1239 2898
rect 1243 2894 1359 2898
rect 1363 2894 1407 2898
rect 1411 2894 1495 2898
rect 1499 2894 1583 2898
rect 1587 2894 1631 2898
rect 1635 2894 1743 2898
rect 1747 2894 1831 2898
rect 1835 2894 1843 2898
rect 91 2893 1843 2894
rect 1849 2893 1850 2899
rect 1842 2853 1843 2859
rect 1849 2858 3619 2859
rect 1849 2854 1871 2858
rect 1875 2854 1895 2858
rect 1899 2854 2079 2858
rect 2083 2854 2135 2858
rect 2139 2854 2263 2858
rect 2267 2854 2287 2858
rect 2291 2854 2391 2858
rect 2395 2854 2479 2858
rect 2483 2854 2519 2858
rect 2523 2854 2647 2858
rect 2651 2854 2663 2858
rect 2667 2854 2767 2858
rect 2771 2854 2831 2858
rect 2835 2854 2887 2858
rect 2891 2854 2991 2858
rect 2995 2854 3007 2858
rect 3011 2854 3135 2858
rect 3139 2854 3143 2858
rect 3147 2854 3295 2858
rect 3299 2854 3447 2858
rect 3451 2854 3591 2858
rect 3595 2854 3619 2858
rect 1849 2853 3619 2854
rect 3625 2853 3626 2859
rect 96 2817 97 2823
rect 103 2822 1855 2823
rect 103 2818 111 2822
rect 115 2818 167 2822
rect 171 2818 303 2822
rect 307 2818 319 2822
rect 323 2818 439 2822
rect 443 2818 447 2822
rect 451 2818 559 2822
rect 563 2818 607 2822
rect 611 2818 687 2822
rect 691 2818 783 2822
rect 787 2818 823 2822
rect 827 2818 959 2822
rect 963 2818 1095 2822
rect 1099 2818 1143 2822
rect 1147 2818 1231 2822
rect 1235 2818 1335 2822
rect 1339 2818 1367 2822
rect 1371 2818 1503 2822
rect 1507 2818 1535 2822
rect 1539 2818 1639 2822
rect 1643 2818 1735 2822
rect 1739 2818 1751 2822
rect 1755 2818 1831 2822
rect 1835 2818 1855 2822
rect 103 2817 1855 2818
rect 1861 2817 1862 2823
rect 1854 2769 1855 2775
rect 1861 2774 3631 2775
rect 1861 2770 1871 2774
rect 1875 2770 2143 2774
rect 2147 2770 2231 2774
rect 2235 2770 2271 2774
rect 2275 2770 2311 2774
rect 2315 2770 2391 2774
rect 2395 2770 2399 2774
rect 2403 2770 2471 2774
rect 2475 2770 2527 2774
rect 2531 2770 2551 2774
rect 2555 2770 2639 2774
rect 2643 2770 2655 2774
rect 2659 2770 2727 2774
rect 2731 2770 2775 2774
rect 2779 2770 2815 2774
rect 2819 2770 2895 2774
rect 2899 2770 2903 2774
rect 2907 2770 2991 2774
rect 2995 2770 3015 2774
rect 3019 2770 3143 2774
rect 3147 2770 3591 2774
rect 3595 2770 3631 2774
rect 1861 2769 3631 2770
rect 3637 2769 3638 2775
rect 84 2737 85 2743
rect 91 2742 1843 2743
rect 91 2738 111 2742
rect 115 2738 135 2742
rect 139 2738 159 2742
rect 163 2738 247 2742
rect 251 2738 295 2742
rect 299 2738 391 2742
rect 395 2738 439 2742
rect 443 2738 551 2742
rect 555 2738 599 2742
rect 603 2738 711 2742
rect 715 2738 775 2742
rect 779 2738 879 2742
rect 883 2738 951 2742
rect 955 2738 1039 2742
rect 1043 2738 1135 2742
rect 1139 2738 1199 2742
rect 1203 2738 1327 2742
rect 1331 2738 1359 2742
rect 1363 2738 1519 2742
rect 1523 2738 1527 2742
rect 1531 2738 1687 2742
rect 1691 2738 1727 2742
rect 1731 2738 1831 2742
rect 1835 2738 1843 2742
rect 91 2737 1843 2738
rect 1849 2737 1850 2743
rect 1842 2693 1843 2699
rect 1849 2698 3619 2699
rect 1849 2694 1871 2698
rect 1875 2694 2223 2698
rect 2227 2694 2239 2698
rect 2243 2694 2303 2698
rect 2307 2694 2319 2698
rect 2323 2694 2383 2698
rect 2387 2694 2399 2698
rect 2403 2694 2463 2698
rect 2467 2694 2479 2698
rect 2483 2694 2543 2698
rect 2547 2694 2559 2698
rect 2563 2694 2631 2698
rect 2635 2694 2639 2698
rect 2643 2694 2719 2698
rect 2723 2694 2799 2698
rect 2803 2694 2807 2698
rect 2811 2694 2879 2698
rect 2883 2694 2895 2698
rect 2899 2694 2959 2698
rect 2963 2694 2983 2698
rect 2987 2694 3591 2698
rect 3595 2694 3619 2698
rect 1849 2693 3619 2694
rect 3625 2693 3626 2699
rect 96 2661 97 2667
rect 103 2666 1855 2667
rect 103 2662 111 2666
rect 115 2662 143 2666
rect 147 2662 255 2666
rect 259 2662 399 2666
rect 403 2662 551 2666
rect 555 2662 559 2666
rect 563 2662 711 2666
rect 715 2662 719 2666
rect 723 2662 879 2666
rect 883 2662 887 2666
rect 891 2662 1047 2666
rect 1051 2662 1207 2666
rect 1211 2662 1215 2666
rect 1219 2662 1367 2666
rect 1371 2662 1391 2666
rect 1395 2662 1527 2666
rect 1531 2662 1567 2666
rect 1571 2662 1695 2666
rect 1699 2662 1831 2666
rect 1835 2662 1855 2666
rect 103 2661 1855 2662
rect 1861 2661 1862 2667
rect 1854 2609 1855 2615
rect 1861 2614 3631 2615
rect 1861 2610 1871 2614
rect 1875 2610 2191 2614
rect 2195 2610 2247 2614
rect 2251 2610 2271 2614
rect 2275 2610 2327 2614
rect 2331 2610 2351 2614
rect 2355 2610 2407 2614
rect 2411 2610 2431 2614
rect 2435 2610 2487 2614
rect 2491 2610 2511 2614
rect 2515 2610 2567 2614
rect 2571 2610 2591 2614
rect 2595 2610 2647 2614
rect 2651 2610 2671 2614
rect 2675 2610 2727 2614
rect 2731 2610 2751 2614
rect 2755 2610 2807 2614
rect 2811 2610 2831 2614
rect 2835 2610 2887 2614
rect 2891 2610 2911 2614
rect 2915 2610 2967 2614
rect 2971 2610 2991 2614
rect 2995 2610 3591 2614
rect 3595 2610 3631 2614
rect 1861 2609 3631 2610
rect 3637 2609 3638 2615
rect 84 2581 85 2587
rect 91 2586 1843 2587
rect 91 2582 111 2586
rect 115 2582 135 2586
rect 139 2582 159 2586
rect 163 2582 247 2586
rect 251 2582 279 2586
rect 283 2582 391 2586
rect 395 2582 415 2586
rect 419 2582 543 2586
rect 547 2582 559 2586
rect 563 2582 703 2586
rect 707 2582 847 2586
rect 851 2582 871 2586
rect 875 2582 983 2586
rect 987 2582 1039 2586
rect 1043 2582 1119 2586
rect 1123 2582 1207 2586
rect 1211 2582 1255 2586
rect 1259 2582 1383 2586
rect 1387 2582 1391 2586
rect 1395 2582 1527 2586
rect 1531 2582 1559 2586
rect 1563 2582 1831 2586
rect 1835 2582 1843 2586
rect 91 2581 1843 2582
rect 1849 2581 1850 2587
rect 1842 2525 1843 2531
rect 1849 2530 3619 2531
rect 1849 2526 1871 2530
rect 1875 2526 2119 2530
rect 2123 2526 2183 2530
rect 2187 2526 2207 2530
rect 2211 2526 2263 2530
rect 2267 2526 2303 2530
rect 2307 2526 2343 2530
rect 2347 2526 2399 2530
rect 2403 2526 2423 2530
rect 2427 2526 2495 2530
rect 2499 2526 2503 2530
rect 2507 2526 2583 2530
rect 2587 2526 2591 2530
rect 2595 2526 2663 2530
rect 2667 2526 2687 2530
rect 2691 2526 2743 2530
rect 2747 2526 2783 2530
rect 2787 2526 2823 2530
rect 2827 2526 2879 2530
rect 2883 2526 2903 2530
rect 2907 2526 2975 2530
rect 2979 2526 2983 2530
rect 2987 2526 3079 2530
rect 3083 2526 3591 2530
rect 3595 2526 3619 2530
rect 1849 2525 3619 2526
rect 3625 2525 3626 2531
rect 96 2501 97 2507
rect 103 2506 1855 2507
rect 103 2502 111 2506
rect 115 2502 167 2506
rect 171 2502 287 2506
rect 291 2502 335 2506
rect 339 2502 415 2506
rect 419 2502 423 2506
rect 427 2502 503 2506
rect 507 2502 567 2506
rect 571 2502 599 2506
rect 603 2502 703 2506
rect 707 2502 711 2506
rect 715 2502 815 2506
rect 819 2502 855 2506
rect 859 2502 935 2506
rect 939 2502 991 2506
rect 995 2502 1063 2506
rect 1067 2502 1127 2506
rect 1131 2502 1191 2506
rect 1195 2502 1263 2506
rect 1267 2502 1327 2506
rect 1331 2502 1399 2506
rect 1403 2502 1471 2506
rect 1475 2502 1535 2506
rect 1539 2502 1831 2506
rect 1835 2502 1855 2506
rect 103 2501 1855 2502
rect 1861 2501 1862 2507
rect 1854 2445 1855 2451
rect 1861 2450 3631 2451
rect 1861 2446 1871 2450
rect 1875 2446 1903 2450
rect 1907 2446 1991 2450
rect 1995 2446 2111 2450
rect 2115 2446 2127 2450
rect 2131 2446 2215 2450
rect 2219 2446 2247 2450
rect 2251 2446 2311 2450
rect 2315 2446 2391 2450
rect 2395 2446 2407 2450
rect 2411 2446 2503 2450
rect 2507 2446 2535 2450
rect 2539 2446 2599 2450
rect 2603 2446 2671 2450
rect 2675 2446 2695 2450
rect 2699 2446 2791 2450
rect 2795 2446 2807 2450
rect 2811 2446 2887 2450
rect 2891 2446 2943 2450
rect 2947 2446 2983 2450
rect 2987 2446 3079 2450
rect 3083 2446 3087 2450
rect 3091 2446 3215 2450
rect 3219 2446 3591 2450
rect 3595 2446 3631 2450
rect 1861 2445 3631 2446
rect 3637 2445 3638 2451
rect 84 2417 85 2423
rect 91 2422 1843 2423
rect 91 2418 111 2422
rect 115 2418 327 2422
rect 331 2418 383 2422
rect 387 2418 407 2422
rect 411 2418 463 2422
rect 467 2418 495 2422
rect 499 2418 543 2422
rect 547 2418 591 2422
rect 595 2418 623 2422
rect 627 2418 695 2422
rect 699 2418 703 2422
rect 707 2418 783 2422
rect 787 2418 807 2422
rect 811 2418 863 2422
rect 867 2418 927 2422
rect 931 2418 943 2422
rect 947 2418 1023 2422
rect 1027 2418 1055 2422
rect 1059 2418 1103 2422
rect 1107 2418 1183 2422
rect 1187 2418 1263 2422
rect 1267 2418 1319 2422
rect 1323 2418 1351 2422
rect 1355 2418 1439 2422
rect 1443 2418 1463 2422
rect 1467 2418 1527 2422
rect 1531 2418 1831 2422
rect 1835 2418 1843 2422
rect 91 2417 1843 2418
rect 1849 2417 1850 2423
rect 1842 2361 1843 2367
rect 1849 2366 3619 2367
rect 1849 2362 1871 2366
rect 1875 2362 1895 2366
rect 1899 2362 1983 2366
rect 1987 2362 2015 2366
rect 2019 2362 2103 2366
rect 2107 2362 2175 2366
rect 2179 2362 2239 2366
rect 2243 2362 2343 2366
rect 2347 2362 2383 2366
rect 2387 2362 2511 2366
rect 2515 2362 2527 2366
rect 2531 2362 2663 2366
rect 2667 2362 2671 2366
rect 2675 2362 2799 2366
rect 2803 2362 2823 2366
rect 2827 2362 2935 2366
rect 2939 2362 2959 2366
rect 2963 2362 3071 2366
rect 3075 2362 3079 2366
rect 3083 2362 3191 2366
rect 3195 2362 3207 2366
rect 3211 2362 3303 2366
rect 3307 2362 3415 2366
rect 3419 2362 3503 2366
rect 3507 2362 3591 2366
rect 3595 2362 3619 2366
rect 1849 2361 3619 2362
rect 3625 2361 3626 2367
rect 96 2341 97 2347
rect 103 2346 1855 2347
rect 103 2342 111 2346
rect 115 2342 391 2346
rect 395 2342 471 2346
rect 475 2342 551 2346
rect 555 2342 631 2346
rect 635 2342 711 2346
rect 715 2342 791 2346
rect 795 2342 871 2346
rect 875 2342 951 2346
rect 955 2342 1031 2346
rect 1035 2342 1111 2346
rect 1115 2342 1191 2346
rect 1195 2342 1271 2346
rect 1275 2342 1359 2346
rect 1363 2342 1407 2346
rect 1411 2342 1447 2346
rect 1451 2342 1487 2346
rect 1491 2342 1535 2346
rect 1539 2342 1567 2346
rect 1571 2342 1647 2346
rect 1651 2342 1831 2346
rect 1835 2342 1855 2346
rect 103 2341 1855 2342
rect 1861 2341 1862 2347
rect 1854 2285 1855 2291
rect 1861 2290 3631 2291
rect 1861 2286 1871 2290
rect 1875 2286 1903 2290
rect 1907 2286 2023 2290
rect 2027 2286 2031 2290
rect 2035 2286 2183 2290
rect 2187 2286 2351 2290
rect 2355 2286 2367 2290
rect 2371 2286 2519 2290
rect 2523 2286 2575 2290
rect 2579 2286 2679 2290
rect 2683 2286 2791 2290
rect 2795 2286 2831 2290
rect 2835 2286 2967 2290
rect 2971 2286 3023 2290
rect 3027 2286 3087 2290
rect 3091 2286 3199 2290
rect 3203 2286 3255 2290
rect 3259 2286 3311 2290
rect 3315 2286 3423 2290
rect 3427 2286 3495 2290
rect 3499 2286 3511 2290
rect 3515 2286 3591 2290
rect 3595 2286 3631 2290
rect 1861 2285 3631 2286
rect 3637 2285 3638 2291
rect 84 2257 85 2263
rect 91 2262 1843 2263
rect 91 2258 111 2262
rect 115 2258 135 2262
rect 139 2258 215 2262
rect 219 2258 295 2262
rect 299 2258 383 2262
rect 387 2258 519 2262
rect 523 2258 671 2262
rect 675 2258 831 2262
rect 835 2258 999 2262
rect 1003 2258 1159 2262
rect 1163 2258 1311 2262
rect 1315 2258 1399 2262
rect 1403 2258 1455 2262
rect 1459 2258 1479 2262
rect 1483 2258 1559 2262
rect 1563 2258 1607 2262
rect 1611 2258 1639 2262
rect 1643 2258 1743 2262
rect 1747 2258 1831 2262
rect 1835 2258 1843 2262
rect 91 2257 1843 2258
rect 1849 2257 1850 2263
rect 1842 2189 1843 2195
rect 1849 2194 3619 2195
rect 1849 2190 1871 2194
rect 1875 2190 1895 2194
rect 1899 2190 2023 2194
rect 2027 2190 2175 2194
rect 2179 2190 2199 2194
rect 2203 2190 2295 2194
rect 2299 2190 2359 2194
rect 2363 2190 2399 2194
rect 2403 2190 2519 2194
rect 2523 2190 2567 2194
rect 2571 2190 2639 2194
rect 2643 2190 2759 2194
rect 2763 2190 2783 2194
rect 2787 2190 2879 2194
rect 2883 2190 2991 2194
rect 2995 2190 3015 2194
rect 3019 2190 3095 2194
rect 3099 2190 3199 2194
rect 3203 2190 3247 2194
rect 3251 2190 3303 2194
rect 3307 2190 3407 2194
rect 3411 2190 3487 2194
rect 3491 2190 3503 2194
rect 3507 2190 3591 2194
rect 3595 2190 3619 2194
rect 1849 2189 3619 2190
rect 3625 2189 3626 2195
rect 96 2177 97 2183
rect 103 2182 1855 2183
rect 103 2178 111 2182
rect 115 2178 143 2182
rect 147 2178 191 2182
rect 195 2178 223 2182
rect 227 2178 303 2182
rect 307 2178 311 2182
rect 315 2178 391 2182
rect 395 2178 463 2182
rect 467 2178 527 2182
rect 531 2178 639 2182
rect 643 2178 679 2182
rect 683 2178 823 2182
rect 827 2178 839 2182
rect 843 2178 1007 2182
rect 1011 2178 1015 2182
rect 1019 2178 1167 2182
rect 1171 2178 1199 2182
rect 1203 2178 1319 2182
rect 1323 2178 1391 2182
rect 1395 2178 1463 2182
rect 1467 2178 1583 2182
rect 1587 2178 1615 2182
rect 1619 2178 1751 2182
rect 1755 2178 1831 2182
rect 1835 2178 1855 2182
rect 103 2177 1855 2178
rect 1861 2177 1862 2183
rect 84 2097 85 2103
rect 91 2102 1843 2103
rect 91 2098 111 2102
rect 115 2098 183 2102
rect 187 2098 215 2102
rect 219 2098 303 2102
rect 307 2098 359 2102
rect 363 2098 455 2102
rect 459 2098 519 2102
rect 523 2098 631 2102
rect 635 2098 703 2102
rect 707 2098 815 2102
rect 819 2098 895 2102
rect 899 2098 1007 2102
rect 1011 2098 1103 2102
rect 1107 2098 1191 2102
rect 1195 2098 1311 2102
rect 1315 2098 1383 2102
rect 1387 2098 1527 2102
rect 1531 2098 1575 2102
rect 1579 2098 1743 2102
rect 1747 2098 1831 2102
rect 1835 2098 1843 2102
rect 91 2097 1843 2098
rect 1849 2097 1850 2103
rect 1854 2101 1855 2107
rect 1861 2106 3631 2107
rect 1861 2102 1871 2106
rect 1875 2102 2175 2106
rect 2179 2102 2207 2106
rect 2211 2102 2271 2106
rect 2275 2102 2303 2106
rect 2307 2102 2375 2106
rect 2379 2102 2407 2106
rect 2411 2102 2487 2106
rect 2491 2102 2527 2106
rect 2531 2102 2607 2106
rect 2611 2102 2647 2106
rect 2651 2102 2727 2106
rect 2731 2102 2767 2106
rect 2771 2102 2847 2106
rect 2851 2102 2887 2106
rect 2891 2102 2967 2106
rect 2971 2102 2999 2106
rect 3003 2102 3079 2106
rect 3083 2102 3103 2106
rect 3107 2102 3191 2106
rect 3195 2102 3207 2106
rect 3211 2102 3303 2106
rect 3307 2102 3311 2106
rect 3315 2102 3415 2106
rect 3419 2102 3511 2106
rect 3515 2102 3591 2106
rect 3595 2102 3631 2106
rect 1861 2101 3631 2102
rect 3637 2101 3638 2107
rect 1842 2031 1843 2037
rect 1849 2031 1874 2037
rect 1868 2027 1874 2031
rect 96 2021 97 2027
rect 103 2026 1855 2027
rect 103 2022 111 2026
rect 115 2022 143 2026
rect 147 2022 223 2026
rect 227 2022 263 2026
rect 267 2022 367 2026
rect 371 2022 383 2026
rect 387 2022 495 2026
rect 499 2022 527 2026
rect 531 2022 607 2026
rect 611 2022 711 2026
rect 715 2022 719 2026
rect 723 2022 823 2026
rect 827 2022 903 2026
rect 907 2022 927 2026
rect 931 2022 1023 2026
rect 1027 2022 1111 2026
rect 1115 2022 1207 2026
rect 1211 2022 1295 2026
rect 1299 2022 1319 2026
rect 1323 2022 1391 2026
rect 1395 2022 1487 2026
rect 1491 2022 1535 2026
rect 1539 2022 1583 2026
rect 1587 2022 1671 2026
rect 1675 2022 1751 2026
rect 1755 2022 1831 2026
rect 1835 2022 1855 2026
rect 103 2021 1855 2022
rect 1861 2021 1862 2027
rect 1868 2026 3619 2027
rect 1868 2022 1871 2026
rect 1875 2022 2071 2026
rect 2075 2022 2167 2026
rect 2171 2022 2207 2026
rect 2211 2022 2263 2026
rect 2267 2022 2359 2026
rect 2363 2022 2367 2026
rect 2371 2022 2479 2026
rect 2483 2022 2519 2026
rect 2523 2022 2599 2026
rect 2603 2022 2679 2026
rect 2683 2022 2719 2026
rect 2723 2022 2839 2026
rect 2843 2022 2847 2026
rect 2851 2022 2959 2026
rect 2963 2022 3015 2026
rect 3019 2022 3071 2026
rect 3075 2022 3183 2026
rect 3187 2022 3295 2026
rect 3299 2022 3351 2026
rect 3355 2022 3407 2026
rect 3411 2022 3503 2026
rect 3507 2022 3591 2026
rect 3595 2022 3619 2026
rect 1868 2021 3619 2022
rect 3625 2021 3626 2027
rect 1854 1945 1855 1951
rect 1861 1950 3631 1951
rect 1861 1946 1871 1950
rect 1875 1946 1903 1950
rect 1907 1946 2007 1950
rect 2011 1946 2079 1950
rect 2083 1946 2135 1950
rect 2139 1946 2215 1950
rect 2219 1946 2255 1950
rect 2259 1946 2367 1950
rect 2371 1946 2375 1950
rect 2379 1946 2487 1950
rect 2491 1946 2527 1950
rect 2531 1946 2599 1950
rect 2603 1946 2687 1950
rect 2691 1946 2719 1950
rect 2723 1946 2839 1950
rect 2843 1946 2855 1950
rect 2859 1946 3023 1950
rect 3027 1946 3191 1950
rect 3195 1946 3359 1950
rect 3363 1946 3511 1950
rect 3515 1946 3591 1950
rect 3595 1946 3631 1950
rect 1861 1945 3631 1946
rect 3637 1945 3638 1951
rect 84 1937 85 1943
rect 91 1942 1843 1943
rect 91 1938 111 1942
rect 115 1938 135 1942
rect 139 1938 167 1942
rect 171 1938 255 1942
rect 259 1938 327 1942
rect 331 1938 375 1942
rect 379 1938 487 1942
rect 491 1938 599 1942
rect 603 1938 647 1942
rect 651 1938 711 1942
rect 715 1938 799 1942
rect 803 1938 815 1942
rect 819 1938 919 1942
rect 923 1938 943 1942
rect 947 1938 1015 1942
rect 1019 1938 1079 1942
rect 1083 1938 1103 1942
rect 1107 1938 1199 1942
rect 1203 1938 1215 1942
rect 1219 1938 1287 1942
rect 1291 1938 1351 1942
rect 1355 1938 1383 1942
rect 1387 1938 1479 1942
rect 1483 1938 1487 1942
rect 1491 1938 1575 1942
rect 1579 1938 1623 1942
rect 1627 1938 1663 1942
rect 1667 1938 1743 1942
rect 1747 1938 1831 1942
rect 1835 1938 1843 1942
rect 91 1937 1843 1938
rect 1849 1937 1850 1943
rect 1842 1871 1843 1877
rect 1849 1875 1874 1877
rect 1849 1874 3619 1875
rect 1849 1871 1871 1874
rect 1868 1870 1871 1871
rect 1875 1870 1895 1874
rect 1899 1870 1991 1874
rect 1995 1870 1999 1874
rect 2003 1870 2119 1874
rect 2123 1870 2127 1874
rect 2131 1870 2247 1874
rect 2251 1870 2367 1874
rect 2371 1870 2383 1874
rect 2387 1870 2479 1874
rect 2483 1870 2519 1874
rect 2523 1870 2591 1874
rect 2595 1870 2655 1874
rect 2659 1870 2711 1874
rect 2715 1870 2807 1874
rect 2811 1870 2831 1874
rect 2835 1870 2975 1874
rect 2979 1870 3151 1874
rect 3155 1870 3335 1874
rect 3339 1870 3503 1874
rect 3507 1870 3591 1874
rect 3595 1870 3619 1874
rect 1868 1869 3619 1870
rect 3625 1869 3626 1875
rect 96 1861 97 1867
rect 103 1866 1855 1867
rect 103 1862 111 1866
rect 115 1862 159 1866
rect 163 1862 175 1866
rect 179 1862 303 1866
rect 307 1862 335 1866
rect 339 1862 447 1866
rect 451 1862 495 1866
rect 499 1862 599 1866
rect 603 1862 655 1866
rect 659 1862 751 1866
rect 755 1862 807 1866
rect 811 1862 903 1866
rect 907 1862 951 1866
rect 955 1862 1055 1866
rect 1059 1862 1087 1866
rect 1091 1862 1207 1866
rect 1211 1862 1223 1866
rect 1227 1862 1351 1866
rect 1355 1862 1359 1866
rect 1363 1862 1487 1866
rect 1491 1862 1495 1866
rect 1499 1862 1631 1866
rect 1635 1862 1751 1866
rect 1755 1862 1831 1866
rect 1835 1862 1855 1866
rect 103 1861 1855 1862
rect 1861 1861 1862 1867
rect 84 1781 85 1787
rect 91 1786 1843 1787
rect 91 1782 111 1786
rect 115 1782 151 1786
rect 155 1782 247 1786
rect 251 1782 295 1786
rect 299 1782 423 1786
rect 427 1782 439 1786
rect 443 1782 591 1786
rect 595 1782 743 1786
rect 747 1782 751 1786
rect 755 1782 895 1786
rect 899 1782 1023 1786
rect 1027 1782 1047 1786
rect 1051 1782 1143 1786
rect 1147 1782 1199 1786
rect 1203 1782 1263 1786
rect 1267 1782 1343 1786
rect 1347 1782 1391 1786
rect 1395 1782 1479 1786
rect 1483 1782 1623 1786
rect 1627 1782 1743 1786
rect 1747 1782 1831 1786
rect 1835 1782 1843 1786
rect 91 1781 1843 1782
rect 1849 1781 1850 1787
rect 1854 1781 1855 1787
rect 1861 1786 3631 1787
rect 1861 1782 1871 1786
rect 1875 1782 1903 1786
rect 1907 1782 1999 1786
rect 2003 1782 2031 1786
rect 2035 1782 2127 1786
rect 2131 1782 2191 1786
rect 2195 1782 2255 1786
rect 2259 1782 2359 1786
rect 2363 1782 2391 1786
rect 2395 1782 2527 1786
rect 2531 1782 2663 1786
rect 2667 1782 2687 1786
rect 2691 1782 2815 1786
rect 2819 1782 2839 1786
rect 2843 1782 2983 1786
rect 2987 1782 3119 1786
rect 3123 1782 3159 1786
rect 3163 1782 3255 1786
rect 3259 1782 3343 1786
rect 3347 1782 3391 1786
rect 3395 1782 3511 1786
rect 3515 1782 3591 1786
rect 3595 1782 3631 1786
rect 1861 1781 3631 1782
rect 3637 1781 3638 1787
rect 1842 1711 1843 1717
rect 1849 1711 1874 1717
rect 1868 1707 1874 1711
rect 96 1701 97 1707
rect 103 1706 1855 1707
rect 103 1702 111 1706
rect 115 1702 191 1706
rect 195 1702 255 1706
rect 259 1702 311 1706
rect 315 1702 431 1706
rect 435 1702 447 1706
rect 451 1702 591 1706
rect 595 1702 599 1706
rect 603 1702 743 1706
rect 747 1702 759 1706
rect 763 1702 895 1706
rect 899 1702 903 1706
rect 907 1702 1031 1706
rect 1035 1702 1039 1706
rect 1043 1702 1151 1706
rect 1155 1702 1183 1706
rect 1187 1702 1271 1706
rect 1275 1702 1319 1706
rect 1323 1702 1399 1706
rect 1403 1702 1447 1706
rect 1451 1702 1575 1706
rect 1579 1702 1711 1706
rect 1715 1702 1831 1706
rect 1835 1702 1855 1706
rect 103 1701 1855 1702
rect 1861 1701 1862 1707
rect 1868 1706 3619 1707
rect 1868 1702 1871 1706
rect 1875 1702 1895 1706
rect 1899 1702 1991 1706
rect 1995 1702 2023 1706
rect 2027 1702 2135 1706
rect 2139 1702 2183 1706
rect 2187 1702 2295 1706
rect 2299 1702 2351 1706
rect 2355 1702 2471 1706
rect 2475 1702 2519 1706
rect 2523 1702 2647 1706
rect 2651 1702 2679 1706
rect 2683 1702 2815 1706
rect 2819 1702 2831 1706
rect 2835 1702 2967 1706
rect 2971 1702 2975 1706
rect 2979 1702 3111 1706
rect 3115 1702 3247 1706
rect 3251 1702 3383 1706
rect 3387 1702 3503 1706
rect 3507 1702 3591 1706
rect 3595 1702 3619 1706
rect 1868 1701 3619 1702
rect 3625 1701 3626 1707
rect 84 1617 85 1623
rect 91 1622 1843 1623
rect 91 1618 111 1622
rect 115 1618 167 1622
rect 171 1618 183 1622
rect 187 1618 303 1622
rect 307 1618 351 1622
rect 355 1618 439 1622
rect 443 1618 543 1622
rect 547 1618 583 1622
rect 587 1618 727 1622
rect 731 1618 735 1622
rect 739 1618 887 1622
rect 891 1618 903 1622
rect 907 1618 1031 1622
rect 1035 1618 1071 1622
rect 1075 1618 1175 1622
rect 1179 1618 1223 1622
rect 1227 1618 1311 1622
rect 1315 1618 1359 1622
rect 1363 1618 1439 1622
rect 1443 1618 1495 1622
rect 1499 1618 1567 1622
rect 1571 1618 1623 1622
rect 1627 1618 1703 1622
rect 1707 1618 1743 1622
rect 1747 1618 1831 1622
rect 1835 1618 1843 1622
rect 91 1617 1843 1618
rect 1849 1617 1850 1623
rect 1854 1621 1855 1627
rect 1861 1626 3631 1627
rect 1861 1622 1871 1626
rect 1875 1622 1903 1626
rect 1907 1622 1975 1626
rect 1979 1622 1999 1626
rect 2003 1622 2095 1626
rect 2099 1622 2143 1626
rect 2147 1622 2231 1626
rect 2235 1622 2303 1626
rect 2307 1622 2367 1626
rect 2371 1622 2479 1626
rect 2483 1622 2503 1626
rect 2507 1622 2639 1626
rect 2643 1622 2655 1626
rect 2659 1622 2775 1626
rect 2779 1622 2823 1626
rect 2827 1622 2911 1626
rect 2915 1622 2975 1626
rect 2979 1622 3055 1626
rect 3059 1622 3119 1626
rect 3123 1622 3207 1626
rect 3211 1622 3255 1626
rect 3259 1622 3367 1626
rect 3371 1622 3391 1626
rect 3395 1622 3511 1626
rect 3515 1622 3591 1626
rect 3595 1622 3631 1626
rect 1861 1621 3631 1622
rect 3637 1621 3638 1627
rect 1842 1547 1843 1553
rect 1849 1547 1874 1553
rect 1868 1546 3619 1547
rect 96 1537 97 1543
rect 103 1542 1855 1543
rect 103 1538 111 1542
rect 115 1538 143 1542
rect 147 1538 175 1542
rect 179 1538 247 1542
rect 251 1538 359 1542
rect 363 1538 383 1542
rect 387 1538 527 1542
rect 531 1538 551 1542
rect 555 1538 671 1542
rect 675 1538 735 1542
rect 739 1538 815 1542
rect 819 1538 911 1542
rect 915 1538 951 1542
rect 955 1538 1079 1542
rect 1083 1538 1207 1542
rect 1211 1538 1231 1542
rect 1235 1538 1335 1542
rect 1339 1538 1367 1542
rect 1371 1538 1471 1542
rect 1475 1538 1503 1542
rect 1507 1538 1631 1542
rect 1635 1538 1751 1542
rect 1755 1538 1831 1542
rect 1835 1538 1855 1542
rect 103 1537 1855 1538
rect 1861 1537 1862 1543
rect 1868 1542 1871 1546
rect 1875 1542 1967 1546
rect 1971 1542 2087 1546
rect 2091 1542 2167 1546
rect 2171 1542 2223 1546
rect 2227 1542 2255 1546
rect 2259 1542 2343 1546
rect 2347 1542 2359 1546
rect 2363 1542 2439 1546
rect 2443 1542 2495 1546
rect 2499 1542 2535 1546
rect 2539 1542 2631 1546
rect 2635 1542 2647 1546
rect 2651 1542 2767 1546
rect 2771 1542 2783 1546
rect 2787 1542 2903 1546
rect 2907 1542 2943 1546
rect 2947 1542 3047 1546
rect 3051 1542 3119 1546
rect 3123 1542 3199 1546
rect 3203 1542 3303 1546
rect 3307 1542 3359 1546
rect 3363 1542 3495 1546
rect 3499 1542 3503 1546
rect 3507 1542 3591 1546
rect 3595 1542 3619 1546
rect 1868 1541 3619 1542
rect 3625 1541 3626 1547
rect 84 1457 85 1463
rect 91 1462 1843 1463
rect 91 1458 111 1462
rect 115 1458 135 1462
rect 139 1458 231 1462
rect 235 1458 239 1462
rect 243 1458 359 1462
rect 363 1458 375 1462
rect 379 1458 479 1462
rect 483 1458 519 1462
rect 523 1458 599 1462
rect 603 1458 663 1462
rect 667 1458 719 1462
rect 723 1458 807 1462
rect 811 1458 831 1462
rect 835 1458 935 1462
rect 939 1458 943 1462
rect 947 1458 1039 1462
rect 1043 1458 1071 1462
rect 1075 1458 1143 1462
rect 1147 1458 1199 1462
rect 1203 1458 1255 1462
rect 1259 1458 1327 1462
rect 1331 1458 1463 1462
rect 1467 1458 1831 1462
rect 1835 1458 1843 1462
rect 91 1457 1843 1458
rect 1849 1457 1850 1463
rect 1854 1461 1855 1467
rect 1861 1466 3631 1467
rect 1861 1462 1871 1466
rect 1875 1462 2095 1466
rect 2099 1462 2175 1466
rect 2179 1462 2263 1466
rect 2267 1462 2343 1466
rect 2347 1462 2351 1466
rect 2355 1462 2423 1466
rect 2427 1462 2447 1466
rect 2451 1462 2503 1466
rect 2507 1462 2543 1466
rect 2547 1462 2607 1466
rect 2611 1462 2655 1466
rect 2659 1462 2735 1466
rect 2739 1462 2791 1466
rect 2795 1462 2895 1466
rect 2899 1462 2951 1466
rect 2955 1462 3079 1466
rect 3083 1462 3127 1466
rect 3131 1462 3279 1466
rect 3283 1462 3311 1466
rect 3315 1462 3479 1466
rect 3483 1462 3503 1466
rect 3507 1462 3591 1466
rect 3595 1462 3631 1466
rect 1861 1461 3631 1462
rect 3637 1461 3638 1467
rect 1842 1385 1843 1391
rect 1849 1390 3619 1391
rect 1849 1386 1871 1390
rect 1875 1386 2255 1390
rect 2259 1386 2263 1390
rect 2267 1386 2335 1390
rect 2339 1386 2343 1390
rect 2347 1386 2415 1390
rect 2419 1386 2423 1390
rect 2427 1386 2495 1390
rect 2499 1386 2503 1390
rect 2507 1386 2591 1390
rect 2595 1386 2599 1390
rect 2603 1386 2695 1390
rect 2699 1386 2727 1390
rect 2731 1386 2807 1390
rect 2811 1386 2887 1390
rect 2891 1386 2919 1390
rect 2923 1386 3039 1390
rect 3043 1386 3071 1390
rect 3075 1386 3159 1390
rect 3163 1386 3271 1390
rect 3275 1386 3279 1390
rect 3283 1386 3399 1390
rect 3403 1386 3471 1390
rect 3475 1386 3503 1390
rect 3507 1386 3591 1390
rect 3595 1386 3619 1390
rect 1849 1385 3619 1386
rect 3625 1385 3626 1391
rect 96 1365 97 1371
rect 103 1370 1855 1371
rect 103 1366 111 1370
rect 115 1366 143 1370
rect 147 1366 239 1370
rect 243 1366 287 1370
rect 291 1366 367 1370
rect 371 1366 431 1370
rect 435 1366 487 1370
rect 491 1366 583 1370
rect 587 1366 607 1370
rect 611 1366 727 1370
rect 731 1366 735 1370
rect 739 1366 839 1370
rect 843 1366 879 1370
rect 883 1366 943 1370
rect 947 1366 1023 1370
rect 1027 1366 1047 1370
rect 1051 1366 1151 1370
rect 1155 1366 1167 1370
rect 1171 1366 1263 1370
rect 1267 1366 1319 1370
rect 1323 1366 1471 1370
rect 1475 1366 1623 1370
rect 1627 1366 1831 1370
rect 1835 1366 1855 1370
rect 103 1365 1855 1366
rect 1861 1365 1862 1371
rect 1854 1297 1855 1303
rect 1861 1302 3631 1303
rect 1861 1298 1871 1302
rect 1875 1298 2215 1302
rect 2219 1298 2271 1302
rect 2275 1298 2295 1302
rect 2299 1298 2351 1302
rect 2355 1298 2375 1302
rect 2379 1298 2431 1302
rect 2435 1298 2455 1302
rect 2459 1298 2511 1302
rect 2515 1298 2551 1302
rect 2555 1298 2599 1302
rect 2603 1298 2663 1302
rect 2667 1298 2703 1302
rect 2707 1298 2791 1302
rect 2795 1298 2815 1302
rect 2819 1298 2927 1302
rect 2931 1298 3047 1302
rect 3051 1298 3071 1302
rect 3075 1298 3167 1302
rect 3171 1298 3215 1302
rect 3219 1298 3287 1302
rect 3291 1298 3367 1302
rect 3371 1298 3407 1302
rect 3411 1298 3511 1302
rect 3515 1298 3591 1302
rect 3595 1298 3631 1302
rect 1861 1297 3631 1298
rect 3637 1297 3638 1303
rect 84 1285 85 1291
rect 91 1290 1843 1291
rect 91 1286 111 1290
rect 115 1286 135 1290
rect 139 1286 263 1290
rect 267 1286 279 1290
rect 283 1286 423 1290
rect 427 1286 575 1290
rect 579 1286 591 1290
rect 595 1286 727 1290
rect 731 1286 759 1290
rect 763 1286 871 1290
rect 875 1286 927 1290
rect 931 1286 1015 1290
rect 1019 1286 1079 1290
rect 1083 1286 1159 1290
rect 1163 1286 1223 1290
rect 1227 1286 1311 1290
rect 1315 1286 1351 1290
rect 1355 1286 1463 1290
rect 1467 1286 1479 1290
rect 1483 1286 1607 1290
rect 1611 1286 1615 1290
rect 1619 1286 1735 1290
rect 1739 1286 1831 1290
rect 1835 1286 1843 1290
rect 91 1285 1843 1286
rect 1849 1285 1850 1291
rect 1842 1217 1843 1223
rect 1849 1222 3619 1223
rect 1849 1218 1871 1222
rect 1875 1218 2111 1222
rect 2115 1218 2207 1222
rect 2211 1218 2287 1222
rect 2291 1218 2303 1222
rect 2307 1218 2367 1222
rect 2371 1218 2407 1222
rect 2411 1218 2447 1222
rect 2451 1218 2527 1222
rect 2531 1218 2543 1222
rect 2547 1218 2647 1222
rect 2651 1218 2655 1222
rect 2659 1218 2775 1222
rect 2779 1218 2783 1222
rect 2787 1218 2911 1222
rect 2915 1218 2919 1222
rect 2923 1218 3055 1222
rect 3059 1218 3063 1222
rect 3067 1218 3199 1222
rect 3203 1218 3207 1222
rect 3211 1218 3343 1222
rect 3347 1218 3359 1222
rect 3363 1218 3495 1222
rect 3499 1218 3503 1222
rect 3507 1218 3591 1222
rect 3595 1218 3619 1222
rect 1849 1217 3619 1218
rect 3625 1217 3626 1223
rect 96 1201 97 1207
rect 103 1206 1855 1207
rect 103 1202 111 1206
rect 115 1202 143 1206
rect 147 1202 271 1206
rect 275 1202 311 1206
rect 315 1202 431 1206
rect 435 1202 487 1206
rect 491 1202 599 1206
rect 603 1202 671 1206
rect 675 1202 767 1206
rect 771 1202 847 1206
rect 851 1202 935 1206
rect 939 1202 1007 1206
rect 1011 1202 1087 1206
rect 1091 1202 1159 1206
rect 1163 1202 1231 1206
rect 1235 1202 1295 1206
rect 1299 1202 1359 1206
rect 1363 1202 1415 1206
rect 1419 1202 1487 1206
rect 1491 1202 1535 1206
rect 1539 1202 1615 1206
rect 1619 1202 1655 1206
rect 1659 1202 1743 1206
rect 1747 1202 1751 1206
rect 1755 1202 1831 1206
rect 1835 1202 1855 1206
rect 103 1201 1855 1202
rect 1861 1201 1862 1207
rect 1854 1133 1855 1139
rect 1861 1138 3631 1139
rect 1861 1134 1871 1138
rect 1875 1134 1903 1138
rect 1907 1134 2119 1138
rect 2123 1134 2127 1138
rect 2131 1134 2215 1138
rect 2219 1134 2311 1138
rect 2315 1134 2359 1138
rect 2363 1134 2415 1138
rect 2419 1134 2535 1138
rect 2539 1134 2575 1138
rect 2579 1134 2655 1138
rect 2659 1134 2775 1138
rect 2779 1134 2783 1138
rect 2787 1134 2919 1138
rect 2923 1134 2967 1138
rect 2971 1134 3063 1138
rect 3067 1134 3159 1138
rect 3163 1134 3207 1138
rect 3211 1134 3343 1138
rect 3347 1134 3351 1138
rect 3355 1134 3503 1138
rect 3507 1134 3511 1138
rect 3515 1134 3591 1138
rect 3595 1134 3631 1138
rect 1861 1133 3631 1134
rect 3637 1133 3638 1139
rect 84 1125 85 1131
rect 91 1130 1843 1131
rect 91 1126 111 1130
rect 115 1126 135 1130
rect 139 1126 247 1130
rect 251 1126 303 1130
rect 307 1126 383 1130
rect 387 1126 479 1130
rect 483 1126 519 1130
rect 523 1126 647 1130
rect 651 1126 663 1130
rect 667 1126 775 1130
rect 779 1126 839 1130
rect 843 1126 895 1130
rect 899 1126 999 1130
rect 1003 1126 1015 1130
rect 1019 1126 1135 1130
rect 1139 1126 1151 1130
rect 1155 1126 1255 1130
rect 1259 1126 1287 1130
rect 1291 1126 1375 1130
rect 1379 1126 1407 1130
rect 1411 1126 1503 1130
rect 1507 1126 1527 1130
rect 1531 1126 1631 1130
rect 1635 1126 1647 1130
rect 1651 1126 1743 1130
rect 1747 1126 1831 1130
rect 1835 1126 1843 1130
rect 91 1125 1843 1126
rect 1849 1125 1850 1131
rect 1842 1057 1843 1063
rect 1849 1062 3619 1063
rect 1849 1058 1871 1062
rect 1875 1058 1895 1062
rect 1899 1058 2015 1062
rect 2019 1058 2119 1062
rect 2123 1058 2167 1062
rect 2171 1058 2327 1062
rect 2331 1058 2351 1062
rect 2355 1058 2487 1062
rect 2491 1058 2567 1062
rect 2571 1058 2639 1062
rect 2643 1058 2767 1062
rect 2771 1058 2791 1062
rect 2795 1058 2935 1062
rect 2939 1058 2959 1062
rect 2963 1058 3079 1062
rect 3083 1058 3151 1062
rect 3155 1058 3223 1062
rect 3227 1058 3335 1062
rect 3339 1058 3375 1062
rect 3379 1058 3503 1062
rect 3507 1058 3591 1062
rect 3595 1058 3619 1062
rect 1849 1057 3619 1058
rect 3625 1057 3626 1063
rect 96 1037 97 1043
rect 103 1042 1855 1043
rect 103 1038 111 1042
rect 115 1038 143 1042
rect 147 1038 239 1042
rect 243 1038 255 1042
rect 259 1038 359 1042
rect 363 1038 391 1042
rect 395 1038 471 1042
rect 475 1038 527 1042
rect 531 1038 575 1042
rect 579 1038 655 1042
rect 659 1038 671 1042
rect 675 1038 767 1042
rect 771 1038 783 1042
rect 787 1038 855 1042
rect 859 1038 903 1042
rect 907 1038 943 1042
rect 947 1038 1023 1042
rect 1027 1038 1031 1042
rect 1035 1038 1127 1042
rect 1131 1038 1143 1042
rect 1147 1038 1223 1042
rect 1227 1038 1263 1042
rect 1267 1038 1383 1042
rect 1387 1038 1511 1042
rect 1515 1038 1639 1042
rect 1643 1038 1751 1042
rect 1755 1038 1831 1042
rect 1835 1038 1855 1042
rect 103 1037 1855 1038
rect 1861 1037 1862 1043
rect 1854 977 1855 983
rect 1861 982 3631 983
rect 1861 978 1871 982
rect 1875 978 1903 982
rect 1907 978 1983 982
rect 1987 978 2023 982
rect 2027 978 2079 982
rect 2083 978 2175 982
rect 2179 978 2199 982
rect 2203 978 2335 982
rect 2339 978 2479 982
rect 2483 978 2495 982
rect 2499 978 2631 982
rect 2635 978 2647 982
rect 2651 978 2791 982
rect 2795 978 2799 982
rect 2803 978 2943 982
rect 2947 978 2967 982
rect 2971 978 3087 982
rect 3091 978 3151 982
rect 3155 978 3231 982
rect 3235 978 3343 982
rect 3347 978 3383 982
rect 3387 978 3511 982
rect 3515 978 3591 982
rect 3595 978 3631 982
rect 1861 977 3631 978
rect 3637 977 3638 983
rect 84 949 85 955
rect 91 954 1843 955
rect 91 950 111 954
rect 115 950 135 954
rect 139 950 231 954
rect 235 950 263 954
rect 267 950 351 954
rect 355 950 415 954
rect 419 950 463 954
rect 467 950 559 954
rect 563 950 567 954
rect 571 950 663 954
rect 667 950 703 954
rect 707 950 759 954
rect 763 950 839 954
rect 843 950 847 954
rect 851 950 935 954
rect 939 950 975 954
rect 979 950 1023 954
rect 1027 950 1103 954
rect 1107 950 1119 954
rect 1123 950 1215 954
rect 1219 950 1223 954
rect 1227 950 1335 954
rect 1339 950 1439 954
rect 1443 950 1543 954
rect 1547 950 1655 954
rect 1659 950 1743 954
rect 1747 950 1831 954
rect 1835 950 1843 954
rect 91 949 1843 950
rect 1849 949 1850 955
rect 1842 889 1843 895
rect 1849 894 3619 895
rect 1849 890 1871 894
rect 1875 890 1895 894
rect 1899 890 1919 894
rect 1923 890 1975 894
rect 1979 890 2071 894
rect 2075 890 2095 894
rect 2099 890 2191 894
rect 2195 890 2271 894
rect 2275 890 2327 894
rect 2331 890 2455 894
rect 2459 890 2471 894
rect 2475 890 2623 894
rect 2627 890 2655 894
rect 2659 890 2783 894
rect 2787 890 2863 894
rect 2867 890 2959 894
rect 2963 890 3079 894
rect 3083 890 3143 894
rect 3147 890 3303 894
rect 3307 890 3335 894
rect 3339 890 3503 894
rect 3507 890 3591 894
rect 3595 890 3619 894
rect 1849 889 3619 890
rect 3625 889 3626 895
rect 96 869 97 875
rect 103 874 1855 875
rect 103 870 111 874
rect 115 870 143 874
rect 147 870 247 874
rect 251 870 271 874
rect 275 870 383 874
rect 387 870 423 874
rect 427 870 519 874
rect 523 870 567 874
rect 571 870 663 874
rect 667 870 711 874
rect 715 870 815 874
rect 819 870 847 874
rect 851 870 959 874
rect 963 870 983 874
rect 987 870 1103 874
rect 1107 870 1111 874
rect 1115 870 1231 874
rect 1235 870 1247 874
rect 1251 870 1343 874
rect 1347 870 1383 874
rect 1387 870 1447 874
rect 1451 870 1511 874
rect 1515 870 1551 874
rect 1555 870 1639 874
rect 1643 870 1663 874
rect 1667 870 1751 874
rect 1755 870 1831 874
rect 1835 870 1855 874
rect 103 869 1855 870
rect 1861 869 1862 875
rect 1854 813 1855 819
rect 1861 818 3631 819
rect 1861 814 1871 818
rect 1875 814 1903 818
rect 1907 814 1927 818
rect 1931 814 2015 818
rect 2019 814 2103 818
rect 2107 814 2167 818
rect 2171 814 2279 818
rect 2283 814 2327 818
rect 2331 814 2463 818
rect 2467 814 2487 818
rect 2491 814 2647 818
rect 2651 814 2663 818
rect 2667 814 2807 818
rect 2811 814 2871 818
rect 2875 814 2959 818
rect 2963 814 3087 818
rect 3091 814 3103 818
rect 3107 814 3247 818
rect 3251 814 3311 818
rect 3315 814 3391 818
rect 3395 814 3511 818
rect 3515 814 3591 818
rect 3595 814 3631 818
rect 1861 813 3631 814
rect 3637 813 3638 819
rect 84 781 85 787
rect 91 786 1843 787
rect 91 782 111 786
rect 115 782 135 786
rect 139 782 215 786
rect 219 782 239 786
rect 243 782 303 786
rect 307 782 375 786
rect 379 782 415 786
rect 419 782 511 786
rect 515 782 543 786
rect 547 782 655 786
rect 659 782 687 786
rect 691 782 807 786
rect 811 782 839 786
rect 843 782 951 786
rect 955 782 991 786
rect 995 782 1095 786
rect 1099 782 1143 786
rect 1147 782 1239 786
rect 1243 782 1295 786
rect 1299 782 1375 786
rect 1379 782 1447 786
rect 1451 782 1503 786
rect 1507 782 1607 786
rect 1611 782 1631 786
rect 1635 782 1743 786
rect 1747 782 1831 786
rect 1835 782 1843 786
rect 91 781 1843 782
rect 1849 781 1850 787
rect 1842 737 1843 743
rect 1849 742 3619 743
rect 1849 738 1871 742
rect 1875 738 1895 742
rect 1899 738 1967 742
rect 1971 738 2007 742
rect 2011 738 2063 742
rect 2067 738 2159 742
rect 2163 738 2175 742
rect 2179 738 2303 742
rect 2307 738 2319 742
rect 2323 738 2447 742
rect 2451 738 2479 742
rect 2483 738 2599 742
rect 2603 738 2639 742
rect 2643 738 2751 742
rect 2755 738 2799 742
rect 2803 738 2903 742
rect 2907 738 2951 742
rect 2955 738 3055 742
rect 3059 738 3095 742
rect 3099 738 3207 742
rect 3211 738 3239 742
rect 3243 738 3359 742
rect 3363 738 3383 742
rect 3387 738 3503 742
rect 3507 738 3591 742
rect 3595 738 3619 742
rect 1849 737 3619 738
rect 3625 737 3626 743
rect 96 697 97 703
rect 103 702 1855 703
rect 103 698 111 702
rect 115 698 143 702
rect 147 698 223 702
rect 227 698 231 702
rect 235 698 311 702
rect 315 698 319 702
rect 323 698 423 702
rect 427 698 543 702
rect 547 698 551 702
rect 555 698 679 702
rect 683 698 695 702
rect 699 698 815 702
rect 819 698 847 702
rect 851 698 951 702
rect 955 698 999 702
rect 1003 698 1087 702
rect 1091 698 1151 702
rect 1155 698 1215 702
rect 1219 698 1303 702
rect 1307 698 1335 702
rect 1339 698 1455 702
rect 1459 698 1583 702
rect 1587 698 1615 702
rect 1619 698 1831 702
rect 1835 698 1855 702
rect 103 697 1855 698
rect 1861 697 1862 703
rect 1854 661 1855 667
rect 1861 666 3631 667
rect 1861 662 1871 666
rect 1875 662 1975 666
rect 1979 662 2071 666
rect 2075 662 2175 666
rect 2179 662 2183 666
rect 2187 662 2271 666
rect 2275 662 2311 666
rect 2315 662 2375 666
rect 2379 662 2455 666
rect 2459 662 2487 666
rect 2491 662 2607 666
rect 2611 662 2735 666
rect 2739 662 2759 666
rect 2763 662 2863 666
rect 2867 662 2911 666
rect 2915 662 2991 666
rect 2995 662 3063 666
rect 3067 662 3119 666
rect 3123 662 3215 666
rect 3219 662 3247 666
rect 3251 662 3367 666
rect 3371 662 3375 666
rect 3379 662 3511 666
rect 3515 662 3591 666
rect 3595 662 3631 666
rect 1861 661 3631 662
rect 3637 661 3638 667
rect 84 613 85 619
rect 91 618 1843 619
rect 91 614 111 618
rect 115 614 223 618
rect 227 614 311 618
rect 315 614 415 618
rect 419 614 447 618
rect 451 614 527 618
rect 531 614 535 618
rect 539 614 607 618
rect 611 614 671 618
rect 675 614 687 618
rect 691 614 775 618
rect 779 614 807 618
rect 811 614 871 618
rect 875 614 943 618
rect 947 614 959 618
rect 963 614 1047 618
rect 1051 614 1079 618
rect 1083 614 1143 618
rect 1147 614 1207 618
rect 1211 614 1239 618
rect 1243 614 1327 618
rect 1331 614 1335 618
rect 1339 614 1431 618
rect 1435 614 1447 618
rect 1451 614 1575 618
rect 1579 614 1831 618
rect 1835 614 1843 618
rect 91 613 1843 614
rect 1849 613 1850 619
rect 1842 585 1843 591
rect 1849 590 3619 591
rect 1849 586 1871 590
rect 1875 586 2167 590
rect 2171 586 2263 590
rect 2267 586 2343 590
rect 2347 586 2367 590
rect 2371 586 2423 590
rect 2427 586 2479 590
rect 2483 586 2503 590
rect 2507 586 2591 590
rect 2595 586 2599 590
rect 2603 586 2695 590
rect 2699 586 2727 590
rect 2731 586 2815 590
rect 2819 586 2855 590
rect 2859 586 2959 590
rect 2963 586 2983 590
rect 2987 586 3111 590
rect 3115 586 3239 590
rect 3243 586 3279 590
rect 3283 586 3367 590
rect 3371 586 3447 590
rect 3451 586 3503 590
rect 3507 586 3591 590
rect 3595 586 3619 590
rect 1849 585 3619 586
rect 3625 585 3626 591
rect 96 525 97 531
rect 103 530 1855 531
rect 103 526 111 530
rect 115 526 335 530
rect 339 526 423 530
rect 427 526 455 530
rect 459 526 511 530
rect 515 526 535 530
rect 539 526 591 530
rect 595 526 615 530
rect 619 526 671 530
rect 675 526 695 530
rect 699 526 751 530
rect 755 526 783 530
rect 787 526 839 530
rect 843 526 879 530
rect 883 526 927 530
rect 931 526 967 530
rect 971 526 1015 530
rect 1019 526 1055 530
rect 1059 526 1103 530
rect 1107 526 1151 530
rect 1155 526 1191 530
rect 1195 526 1247 530
rect 1251 526 1279 530
rect 1283 526 1343 530
rect 1347 526 1439 530
rect 1443 526 1831 530
rect 1835 526 1855 530
rect 103 525 1855 526
rect 1861 525 1862 531
rect 1854 501 1855 507
rect 1861 506 3631 507
rect 1861 502 1871 506
rect 1875 502 2191 506
rect 2195 502 2271 506
rect 2275 502 2287 506
rect 2291 502 2351 506
rect 2355 502 2383 506
rect 2387 502 2431 506
rect 2435 502 2487 506
rect 2491 502 2511 506
rect 2515 502 2583 506
rect 2587 502 2599 506
rect 2603 502 2687 506
rect 2691 502 2703 506
rect 2707 502 2791 506
rect 2795 502 2823 506
rect 2827 502 2911 506
rect 2915 502 2967 506
rect 2971 502 3039 506
rect 3043 502 3119 506
rect 3123 502 3175 506
rect 3179 502 3287 506
rect 3291 502 3319 506
rect 3323 502 3455 506
rect 3459 502 3471 506
rect 3475 502 3591 506
rect 3595 502 3631 506
rect 1861 501 3631 502
rect 3637 501 3638 507
rect 84 441 85 447
rect 91 446 1843 447
rect 91 442 111 446
rect 115 442 223 446
rect 227 442 327 446
rect 331 442 335 446
rect 339 442 415 446
rect 419 442 447 446
rect 451 442 503 446
rect 507 442 559 446
rect 563 442 583 446
rect 587 442 663 446
rect 667 442 743 446
rect 747 442 759 446
rect 763 442 831 446
rect 835 442 847 446
rect 851 442 919 446
rect 923 442 935 446
rect 939 442 1007 446
rect 1011 442 1023 446
rect 1027 442 1095 446
rect 1099 442 1111 446
rect 1115 442 1183 446
rect 1187 442 1199 446
rect 1203 442 1271 446
rect 1275 442 1295 446
rect 1299 442 1831 446
rect 1835 442 1843 446
rect 91 441 1843 442
rect 1849 441 1850 447
rect 1842 421 1843 427
rect 1849 426 3619 427
rect 1849 422 1871 426
rect 1875 422 1975 426
rect 1979 422 2063 426
rect 2067 422 2159 426
rect 2163 422 2183 426
rect 2187 422 2255 426
rect 2259 422 2279 426
rect 2283 422 2359 426
rect 2363 422 2375 426
rect 2379 422 2471 426
rect 2475 422 2479 426
rect 2483 422 2575 426
rect 2579 422 2607 426
rect 2611 422 2679 426
rect 2683 422 2759 426
rect 2763 422 2783 426
rect 2787 422 2903 426
rect 2907 422 2927 426
rect 2931 422 3031 426
rect 3035 422 3111 426
rect 3115 422 3167 426
rect 3171 422 3303 426
rect 3307 422 3311 426
rect 3315 422 3463 426
rect 3467 422 3495 426
rect 3499 422 3591 426
rect 3595 422 3619 426
rect 1849 421 3619 422
rect 3625 421 3626 427
rect 96 353 97 359
rect 103 358 1855 359
rect 103 354 111 358
rect 115 354 143 358
rect 147 354 231 358
rect 235 354 263 358
rect 267 354 343 358
rect 347 354 399 358
rect 403 354 455 358
rect 459 354 535 358
rect 539 354 567 358
rect 571 354 671 358
rect 675 354 767 358
rect 771 354 791 358
rect 795 354 855 358
rect 859 354 911 358
rect 915 354 943 358
rect 947 354 1023 358
rect 1027 354 1031 358
rect 1035 354 1119 358
rect 1123 354 1127 358
rect 1131 354 1207 358
rect 1211 354 1231 358
rect 1235 354 1303 358
rect 1307 354 1335 358
rect 1339 354 1439 358
rect 1443 354 1831 358
rect 1835 354 1855 358
rect 103 353 1855 354
rect 1861 353 1862 359
rect 1854 341 1855 347
rect 1861 346 3631 347
rect 1861 342 1871 346
rect 1875 342 1983 346
rect 1987 342 2071 346
rect 2075 342 2167 346
rect 2171 342 2215 346
rect 2219 342 2263 346
rect 2267 342 2295 346
rect 2299 342 2367 346
rect 2371 342 2383 346
rect 2387 342 2479 346
rect 2483 342 2591 346
rect 2595 342 2615 346
rect 2619 342 2719 346
rect 2723 342 2767 346
rect 2771 342 2847 346
rect 2851 342 2935 346
rect 2939 342 2983 346
rect 2987 342 3119 346
rect 3123 342 3255 346
rect 3259 342 3311 346
rect 3315 342 3391 346
rect 3395 342 3503 346
rect 3507 342 3511 346
rect 3515 342 3591 346
rect 3595 342 3631 346
rect 1861 341 3631 342
rect 3637 341 3638 347
rect 84 269 85 275
rect 91 274 1843 275
rect 91 270 111 274
rect 115 270 135 274
rect 139 270 247 274
rect 251 270 255 274
rect 259 270 391 274
rect 395 270 527 274
rect 531 270 543 274
rect 547 270 663 274
rect 667 270 695 274
rect 699 270 783 274
rect 787 270 847 274
rect 851 270 903 274
rect 907 270 991 274
rect 995 270 1015 274
rect 1019 270 1119 274
rect 1123 270 1223 274
rect 1227 270 1239 274
rect 1243 270 1327 274
rect 1331 270 1359 274
rect 1363 270 1431 274
rect 1435 270 1479 274
rect 1483 270 1599 274
rect 1603 270 1831 274
rect 1835 270 1843 274
rect 91 269 1843 270
rect 1849 269 1850 275
rect 1842 267 1850 269
rect 1842 261 1843 267
rect 1849 266 3619 267
rect 1849 262 1871 266
rect 1875 262 1991 266
rect 1995 262 2119 266
rect 2123 262 2207 266
rect 2211 262 2255 266
rect 2259 262 2287 266
rect 2291 262 2375 266
rect 2379 262 2391 266
rect 2395 262 2471 266
rect 2475 262 2535 266
rect 2539 262 2583 266
rect 2587 262 2679 266
rect 2683 262 2711 266
rect 2715 262 2815 266
rect 2819 262 2839 266
rect 2843 262 2951 266
rect 2955 262 2975 266
rect 2979 262 3095 266
rect 3099 262 3111 266
rect 3115 262 3239 266
rect 3243 262 3247 266
rect 3251 262 3383 266
rect 3387 262 3503 266
rect 3507 262 3591 266
rect 3595 262 3619 266
rect 1849 261 3619 262
rect 3625 261 3626 267
rect 1854 173 1855 179
rect 1861 178 3631 179
rect 1861 174 1871 178
rect 1875 174 1903 178
rect 1907 174 1983 178
rect 1987 174 1999 178
rect 2003 174 2087 178
rect 2091 174 2127 178
rect 2131 174 2215 178
rect 2219 174 2263 178
rect 2267 174 2351 178
rect 2355 174 2399 178
rect 2403 174 2487 178
rect 2491 174 2543 178
rect 2547 174 2623 178
rect 2627 174 2687 178
rect 2691 174 2743 178
rect 2747 174 2823 178
rect 2827 174 2855 178
rect 2859 174 2959 178
rect 2963 174 3063 178
rect 3067 174 3103 178
rect 3107 174 3159 178
rect 3163 174 3247 178
rect 3251 174 3343 178
rect 3347 174 3391 178
rect 3395 174 3431 178
rect 3435 174 3511 178
rect 3515 174 3591 178
rect 3595 174 3631 178
rect 1861 173 3631 174
rect 3637 173 3638 179
rect 96 157 97 163
rect 103 162 1855 163
rect 103 158 111 162
rect 115 158 143 162
rect 147 158 223 162
rect 227 158 255 162
rect 259 158 303 162
rect 307 158 383 162
rect 387 158 399 162
rect 403 158 463 162
rect 467 158 543 162
rect 547 158 551 162
rect 555 158 623 162
rect 627 158 703 162
rect 707 158 783 162
rect 787 158 855 162
rect 859 158 863 162
rect 867 158 943 162
rect 947 158 999 162
rect 1003 158 1023 162
rect 1027 158 1103 162
rect 1107 158 1127 162
rect 1131 158 1183 162
rect 1187 158 1247 162
rect 1251 158 1263 162
rect 1267 158 1343 162
rect 1347 158 1367 162
rect 1371 158 1423 162
rect 1427 158 1487 162
rect 1491 158 1511 162
rect 1515 158 1591 162
rect 1595 158 1607 162
rect 1611 158 1671 162
rect 1675 158 1751 162
rect 1755 158 1831 162
rect 1835 158 1855 162
rect 103 157 1855 158
rect 1861 157 1862 163
rect 1842 97 1843 103
rect 1849 102 3619 103
rect 1849 98 1871 102
rect 1875 98 1895 102
rect 1899 98 1975 102
rect 1979 98 2079 102
rect 2083 98 2207 102
rect 2211 98 2343 102
rect 2347 98 2479 102
rect 2483 98 2615 102
rect 2619 98 2735 102
rect 2739 98 2847 102
rect 2851 98 2951 102
rect 2955 98 3055 102
rect 3059 98 3151 102
rect 3155 98 3239 102
rect 3243 98 3335 102
rect 3339 98 3423 102
rect 3427 98 3503 102
rect 3507 98 3591 102
rect 3595 98 3619 102
rect 1849 97 3619 98
rect 3625 97 3626 103
rect 84 81 85 87
rect 91 86 1843 87
rect 91 82 111 86
rect 115 82 135 86
rect 139 82 215 86
rect 219 82 295 86
rect 299 82 375 86
rect 379 82 455 86
rect 459 82 535 86
rect 539 82 615 86
rect 619 82 695 86
rect 699 82 775 86
rect 779 82 855 86
rect 859 82 935 86
rect 939 82 1015 86
rect 1019 82 1095 86
rect 1099 82 1175 86
rect 1179 82 1255 86
rect 1259 82 1335 86
rect 1339 82 1415 86
rect 1419 82 1503 86
rect 1507 82 1583 86
rect 1587 82 1663 86
rect 1667 82 1743 86
rect 1747 82 1831 86
rect 1835 82 1843 86
rect 91 81 1843 82
rect 1849 81 1850 87
<< m5c >>
rect 85 3665 91 3671
rect 1843 3665 1849 3671
rect 1855 3597 1861 3603
rect 3631 3597 3637 3603
rect 97 3589 103 3595
rect 1855 3589 1861 3595
rect 1843 3521 1849 3527
rect 3619 3521 3625 3527
rect 85 3513 91 3519
rect 1843 3513 1849 3519
rect 97 3437 103 3443
rect 1855 3437 1861 3443
rect 85 3361 91 3367
rect 1843 3361 1849 3367
rect 97 3281 103 3287
rect 1855 3281 1861 3287
rect 1855 3269 1861 3275
rect 3631 3269 3637 3275
rect 85 3205 91 3211
rect 1843 3205 1849 3211
rect 1843 3189 1849 3195
rect 3619 3189 3625 3195
rect 97 3125 103 3131
rect 1855 3125 1861 3131
rect 1855 3097 1861 3103
rect 3631 3097 3637 3103
rect 85 3045 91 3051
rect 1843 3045 1849 3051
rect 1843 3013 1849 3019
rect 3619 3013 3625 3019
rect 97 2969 103 2975
rect 1855 2969 1861 2975
rect 1855 2937 1861 2943
rect 3631 2937 3637 2943
rect 85 2893 91 2899
rect 1843 2893 1849 2899
rect 1843 2853 1849 2859
rect 3619 2853 3625 2859
rect 97 2817 103 2823
rect 1855 2817 1861 2823
rect 1855 2769 1861 2775
rect 3631 2769 3637 2775
rect 85 2737 91 2743
rect 1843 2737 1849 2743
rect 1843 2693 1849 2699
rect 3619 2693 3625 2699
rect 97 2661 103 2667
rect 1855 2661 1861 2667
rect 1855 2609 1861 2615
rect 3631 2609 3637 2615
rect 85 2581 91 2587
rect 1843 2581 1849 2587
rect 1843 2525 1849 2531
rect 3619 2525 3625 2531
rect 97 2501 103 2507
rect 1855 2501 1861 2507
rect 1855 2445 1861 2451
rect 3631 2445 3637 2451
rect 85 2417 91 2423
rect 1843 2417 1849 2423
rect 1843 2361 1849 2367
rect 3619 2361 3625 2367
rect 97 2341 103 2347
rect 1855 2341 1861 2347
rect 1855 2285 1861 2291
rect 3631 2285 3637 2291
rect 85 2257 91 2263
rect 1843 2257 1849 2263
rect 1843 2189 1849 2195
rect 3619 2189 3625 2195
rect 97 2177 103 2183
rect 1855 2177 1861 2183
rect 85 2097 91 2103
rect 1843 2097 1849 2103
rect 1855 2101 1861 2107
rect 3631 2101 3637 2107
rect 1843 2031 1849 2037
rect 97 2021 103 2027
rect 1855 2021 1861 2027
rect 3619 2021 3625 2027
rect 1855 1945 1861 1951
rect 3631 1945 3637 1951
rect 85 1937 91 1943
rect 1843 1937 1849 1943
rect 1843 1871 1849 1877
rect 3619 1869 3625 1875
rect 97 1861 103 1867
rect 1855 1861 1861 1867
rect 85 1781 91 1787
rect 1843 1781 1849 1787
rect 1855 1781 1861 1787
rect 3631 1781 3637 1787
rect 1843 1711 1849 1717
rect 97 1701 103 1707
rect 1855 1701 1861 1707
rect 3619 1701 3625 1707
rect 85 1617 91 1623
rect 1843 1617 1849 1623
rect 1855 1621 1861 1627
rect 3631 1621 3637 1627
rect 1843 1547 1849 1553
rect 97 1537 103 1543
rect 1855 1537 1861 1543
rect 3619 1541 3625 1547
rect 85 1457 91 1463
rect 1843 1457 1849 1463
rect 1855 1461 1861 1467
rect 3631 1461 3637 1467
rect 1843 1385 1849 1391
rect 3619 1385 3625 1391
rect 97 1365 103 1371
rect 1855 1365 1861 1371
rect 1855 1297 1861 1303
rect 3631 1297 3637 1303
rect 85 1285 91 1291
rect 1843 1285 1849 1291
rect 1843 1217 1849 1223
rect 3619 1217 3625 1223
rect 97 1201 103 1207
rect 1855 1201 1861 1207
rect 1855 1133 1861 1139
rect 3631 1133 3637 1139
rect 85 1125 91 1131
rect 1843 1125 1849 1131
rect 1843 1057 1849 1063
rect 3619 1057 3625 1063
rect 97 1037 103 1043
rect 1855 1037 1861 1043
rect 1855 977 1861 983
rect 3631 977 3637 983
rect 85 949 91 955
rect 1843 949 1849 955
rect 1843 889 1849 895
rect 3619 889 3625 895
rect 97 869 103 875
rect 1855 869 1861 875
rect 1855 813 1861 819
rect 3631 813 3637 819
rect 85 781 91 787
rect 1843 781 1849 787
rect 1843 737 1849 743
rect 3619 737 3625 743
rect 97 697 103 703
rect 1855 697 1861 703
rect 1855 661 1861 667
rect 3631 661 3637 667
rect 85 613 91 619
rect 1843 613 1849 619
rect 1843 585 1849 591
rect 3619 585 3625 591
rect 97 525 103 531
rect 1855 525 1861 531
rect 1855 501 1861 507
rect 3631 501 3637 507
rect 85 441 91 447
rect 1843 441 1849 447
rect 1843 421 1849 427
rect 3619 421 3625 427
rect 97 353 103 359
rect 1855 353 1861 359
rect 1855 341 1861 347
rect 3631 341 3637 347
rect 85 269 91 275
rect 1843 269 1849 275
rect 1843 261 1849 267
rect 3619 261 3625 267
rect 1855 173 1861 179
rect 3631 173 3637 179
rect 97 157 103 163
rect 1855 157 1861 163
rect 1843 97 1849 103
rect 3619 97 3625 103
rect 85 81 91 87
rect 1843 81 1849 87
<< m5 >>
rect 84 3671 92 3672
rect 84 3665 85 3671
rect 91 3665 92 3671
rect 84 3519 92 3665
rect 84 3513 85 3519
rect 91 3513 92 3519
rect 84 3367 92 3513
rect 84 3361 85 3367
rect 91 3361 92 3367
rect 84 3211 92 3361
rect 84 3205 85 3211
rect 91 3205 92 3211
rect 84 3051 92 3205
rect 84 3045 85 3051
rect 91 3045 92 3051
rect 84 2899 92 3045
rect 84 2893 85 2899
rect 91 2893 92 2899
rect 84 2743 92 2893
rect 84 2737 85 2743
rect 91 2737 92 2743
rect 84 2587 92 2737
rect 84 2581 85 2587
rect 91 2581 92 2587
rect 84 2423 92 2581
rect 84 2417 85 2423
rect 91 2417 92 2423
rect 84 2263 92 2417
rect 84 2257 85 2263
rect 91 2257 92 2263
rect 84 2103 92 2257
rect 84 2097 85 2103
rect 91 2097 92 2103
rect 84 1943 92 2097
rect 84 1937 85 1943
rect 91 1937 92 1943
rect 84 1787 92 1937
rect 84 1781 85 1787
rect 91 1781 92 1787
rect 84 1623 92 1781
rect 84 1617 85 1623
rect 91 1617 92 1623
rect 84 1463 92 1617
rect 84 1457 85 1463
rect 91 1457 92 1463
rect 84 1291 92 1457
rect 84 1285 85 1291
rect 91 1285 92 1291
rect 84 1131 92 1285
rect 84 1125 85 1131
rect 91 1125 92 1131
rect 84 955 92 1125
rect 84 949 85 955
rect 91 949 92 955
rect 84 787 92 949
rect 84 781 85 787
rect 91 781 92 787
rect 84 619 92 781
rect 84 613 85 619
rect 91 613 92 619
rect 84 447 92 613
rect 84 441 85 447
rect 91 441 92 447
rect 84 275 92 441
rect 84 269 85 275
rect 91 269 92 275
rect 84 87 92 269
rect 84 81 85 87
rect 91 81 92 87
rect 84 72 92 81
rect 96 3595 104 3672
rect 96 3589 97 3595
rect 103 3589 104 3595
rect 96 3443 104 3589
rect 96 3437 97 3443
rect 103 3437 104 3443
rect 96 3287 104 3437
rect 96 3281 97 3287
rect 103 3281 104 3287
rect 96 3131 104 3281
rect 96 3125 97 3131
rect 103 3125 104 3131
rect 96 2975 104 3125
rect 96 2969 97 2975
rect 103 2969 104 2975
rect 96 2823 104 2969
rect 96 2817 97 2823
rect 103 2817 104 2823
rect 96 2667 104 2817
rect 96 2661 97 2667
rect 103 2661 104 2667
rect 96 2507 104 2661
rect 96 2501 97 2507
rect 103 2501 104 2507
rect 96 2347 104 2501
rect 96 2341 97 2347
rect 103 2341 104 2347
rect 96 2183 104 2341
rect 96 2177 97 2183
rect 103 2177 104 2183
rect 96 2027 104 2177
rect 96 2021 97 2027
rect 103 2021 104 2027
rect 96 1867 104 2021
rect 96 1861 97 1867
rect 103 1861 104 1867
rect 96 1707 104 1861
rect 96 1701 97 1707
rect 103 1701 104 1707
rect 96 1543 104 1701
rect 96 1537 97 1543
rect 103 1537 104 1543
rect 96 1371 104 1537
rect 96 1365 97 1371
rect 103 1365 104 1371
rect 96 1207 104 1365
rect 96 1201 97 1207
rect 103 1201 104 1207
rect 96 1043 104 1201
rect 96 1037 97 1043
rect 103 1037 104 1043
rect 96 875 104 1037
rect 96 869 97 875
rect 103 869 104 875
rect 96 703 104 869
rect 96 697 97 703
rect 103 697 104 703
rect 96 531 104 697
rect 96 525 97 531
rect 103 525 104 531
rect 96 359 104 525
rect 96 353 97 359
rect 103 353 104 359
rect 96 163 104 353
rect 96 157 97 163
rect 103 157 104 163
rect 96 72 104 157
rect 1842 3671 1850 3672
rect 1842 3665 1843 3671
rect 1849 3665 1850 3671
rect 1842 3527 1850 3665
rect 1842 3521 1843 3527
rect 1849 3521 1850 3527
rect 1842 3519 1850 3521
rect 1842 3513 1843 3519
rect 1849 3513 1850 3519
rect 1842 3367 1850 3513
rect 1842 3361 1843 3367
rect 1849 3361 1850 3367
rect 1842 3211 1850 3361
rect 1842 3205 1843 3211
rect 1849 3205 1850 3211
rect 1842 3195 1850 3205
rect 1842 3189 1843 3195
rect 1849 3189 1850 3195
rect 1842 3051 1850 3189
rect 1842 3045 1843 3051
rect 1849 3045 1850 3051
rect 1842 3019 1850 3045
rect 1842 3013 1843 3019
rect 1849 3013 1850 3019
rect 1842 2899 1850 3013
rect 1842 2893 1843 2899
rect 1849 2893 1850 2899
rect 1842 2859 1850 2893
rect 1842 2853 1843 2859
rect 1849 2853 1850 2859
rect 1842 2743 1850 2853
rect 1842 2737 1843 2743
rect 1849 2737 1850 2743
rect 1842 2699 1850 2737
rect 1842 2693 1843 2699
rect 1849 2693 1850 2699
rect 1842 2587 1850 2693
rect 1842 2581 1843 2587
rect 1849 2581 1850 2587
rect 1842 2531 1850 2581
rect 1842 2525 1843 2531
rect 1849 2525 1850 2531
rect 1842 2423 1850 2525
rect 1842 2417 1843 2423
rect 1849 2417 1850 2423
rect 1842 2367 1850 2417
rect 1842 2361 1843 2367
rect 1849 2361 1850 2367
rect 1842 2263 1850 2361
rect 1842 2257 1843 2263
rect 1849 2257 1850 2263
rect 1842 2195 1850 2257
rect 1842 2189 1843 2195
rect 1849 2189 1850 2195
rect 1842 2103 1850 2189
rect 1842 2097 1843 2103
rect 1849 2097 1850 2103
rect 1842 2037 1850 2097
rect 1842 2031 1843 2037
rect 1849 2031 1850 2037
rect 1842 1943 1850 2031
rect 1842 1937 1843 1943
rect 1849 1937 1850 1943
rect 1842 1877 1850 1937
rect 1842 1871 1843 1877
rect 1849 1871 1850 1877
rect 1842 1787 1850 1871
rect 1842 1781 1843 1787
rect 1849 1781 1850 1787
rect 1842 1717 1850 1781
rect 1842 1711 1843 1717
rect 1849 1711 1850 1717
rect 1842 1623 1850 1711
rect 1842 1617 1843 1623
rect 1849 1617 1850 1623
rect 1842 1553 1850 1617
rect 1842 1547 1843 1553
rect 1849 1547 1850 1553
rect 1842 1463 1850 1547
rect 1842 1457 1843 1463
rect 1849 1457 1850 1463
rect 1842 1391 1850 1457
rect 1842 1385 1843 1391
rect 1849 1385 1850 1391
rect 1842 1291 1850 1385
rect 1842 1285 1843 1291
rect 1849 1285 1850 1291
rect 1842 1223 1850 1285
rect 1842 1217 1843 1223
rect 1849 1217 1850 1223
rect 1842 1131 1850 1217
rect 1842 1125 1843 1131
rect 1849 1125 1850 1131
rect 1842 1063 1850 1125
rect 1842 1057 1843 1063
rect 1849 1057 1850 1063
rect 1842 955 1850 1057
rect 1842 949 1843 955
rect 1849 949 1850 955
rect 1842 895 1850 949
rect 1842 889 1843 895
rect 1849 889 1850 895
rect 1842 787 1850 889
rect 1842 781 1843 787
rect 1849 781 1850 787
rect 1842 743 1850 781
rect 1842 737 1843 743
rect 1849 737 1850 743
rect 1842 619 1850 737
rect 1842 613 1843 619
rect 1849 613 1850 619
rect 1842 591 1850 613
rect 1842 585 1843 591
rect 1849 585 1850 591
rect 1842 447 1850 585
rect 1842 441 1843 447
rect 1849 441 1850 447
rect 1842 427 1850 441
rect 1842 421 1843 427
rect 1849 421 1850 427
rect 1842 275 1850 421
rect 1842 269 1843 275
rect 1849 269 1850 275
rect 1842 267 1850 269
rect 1842 261 1843 267
rect 1849 261 1850 267
rect 1842 103 1850 261
rect 1842 97 1843 103
rect 1849 97 1850 103
rect 1842 87 1850 97
rect 1842 81 1843 87
rect 1849 81 1850 87
rect 1842 72 1850 81
rect 1854 3603 1862 3672
rect 1854 3597 1855 3603
rect 1861 3597 1862 3603
rect 1854 3595 1862 3597
rect 1854 3589 1855 3595
rect 1861 3589 1862 3595
rect 1854 3443 1862 3589
rect 1854 3437 1855 3443
rect 1861 3437 1862 3443
rect 1854 3287 1862 3437
rect 1854 3281 1855 3287
rect 1861 3281 1862 3287
rect 1854 3275 1862 3281
rect 1854 3269 1855 3275
rect 1861 3269 1862 3275
rect 1854 3131 1862 3269
rect 1854 3125 1855 3131
rect 1861 3125 1862 3131
rect 1854 3103 1862 3125
rect 1854 3097 1855 3103
rect 1861 3097 1862 3103
rect 1854 2975 1862 3097
rect 1854 2969 1855 2975
rect 1861 2969 1862 2975
rect 1854 2943 1862 2969
rect 1854 2937 1855 2943
rect 1861 2937 1862 2943
rect 1854 2823 1862 2937
rect 1854 2817 1855 2823
rect 1861 2817 1862 2823
rect 1854 2775 1862 2817
rect 1854 2769 1855 2775
rect 1861 2769 1862 2775
rect 1854 2667 1862 2769
rect 1854 2661 1855 2667
rect 1861 2661 1862 2667
rect 1854 2615 1862 2661
rect 1854 2609 1855 2615
rect 1861 2609 1862 2615
rect 1854 2507 1862 2609
rect 1854 2501 1855 2507
rect 1861 2501 1862 2507
rect 1854 2451 1862 2501
rect 1854 2445 1855 2451
rect 1861 2445 1862 2451
rect 1854 2347 1862 2445
rect 1854 2341 1855 2347
rect 1861 2341 1862 2347
rect 1854 2291 1862 2341
rect 1854 2285 1855 2291
rect 1861 2285 1862 2291
rect 1854 2183 1862 2285
rect 1854 2177 1855 2183
rect 1861 2177 1862 2183
rect 1854 2107 1862 2177
rect 1854 2101 1855 2107
rect 1861 2101 1862 2107
rect 1854 2027 1862 2101
rect 1854 2021 1855 2027
rect 1861 2021 1862 2027
rect 1854 1951 1862 2021
rect 1854 1945 1855 1951
rect 1861 1945 1862 1951
rect 1854 1867 1862 1945
rect 1854 1861 1855 1867
rect 1861 1861 1862 1867
rect 1854 1787 1862 1861
rect 1854 1781 1855 1787
rect 1861 1781 1862 1787
rect 1854 1707 1862 1781
rect 1854 1701 1855 1707
rect 1861 1701 1862 1707
rect 1854 1627 1862 1701
rect 1854 1621 1855 1627
rect 1861 1621 1862 1627
rect 1854 1543 1862 1621
rect 1854 1537 1855 1543
rect 1861 1537 1862 1543
rect 1854 1467 1862 1537
rect 1854 1461 1855 1467
rect 1861 1461 1862 1467
rect 1854 1371 1862 1461
rect 1854 1365 1855 1371
rect 1861 1365 1862 1371
rect 1854 1303 1862 1365
rect 1854 1297 1855 1303
rect 1861 1297 1862 1303
rect 1854 1207 1862 1297
rect 1854 1201 1855 1207
rect 1861 1201 1862 1207
rect 1854 1139 1862 1201
rect 1854 1133 1855 1139
rect 1861 1133 1862 1139
rect 1854 1043 1862 1133
rect 1854 1037 1855 1043
rect 1861 1037 1862 1043
rect 1854 983 1862 1037
rect 1854 977 1855 983
rect 1861 977 1862 983
rect 1854 875 1862 977
rect 1854 869 1855 875
rect 1861 869 1862 875
rect 1854 819 1862 869
rect 1854 813 1855 819
rect 1861 813 1862 819
rect 1854 703 1862 813
rect 1854 697 1855 703
rect 1861 697 1862 703
rect 1854 667 1862 697
rect 1854 661 1855 667
rect 1861 661 1862 667
rect 1854 531 1862 661
rect 1854 525 1855 531
rect 1861 525 1862 531
rect 1854 507 1862 525
rect 1854 501 1855 507
rect 1861 501 1862 507
rect 1854 359 1862 501
rect 1854 353 1855 359
rect 1861 353 1862 359
rect 1854 347 1862 353
rect 1854 341 1855 347
rect 1861 341 1862 347
rect 1854 179 1862 341
rect 1854 173 1855 179
rect 1861 173 1862 179
rect 1854 163 1862 173
rect 1854 157 1855 163
rect 1861 157 1862 163
rect 1854 72 1862 157
rect 3618 3527 3626 3672
rect 3618 3521 3619 3527
rect 3625 3521 3626 3527
rect 3618 3195 3626 3521
rect 3618 3189 3619 3195
rect 3625 3189 3626 3195
rect 3618 3019 3626 3189
rect 3618 3013 3619 3019
rect 3625 3013 3626 3019
rect 3618 2859 3626 3013
rect 3618 2853 3619 2859
rect 3625 2853 3626 2859
rect 3618 2699 3626 2853
rect 3618 2693 3619 2699
rect 3625 2693 3626 2699
rect 3618 2531 3626 2693
rect 3618 2525 3619 2531
rect 3625 2525 3626 2531
rect 3618 2367 3626 2525
rect 3618 2361 3619 2367
rect 3625 2361 3626 2367
rect 3618 2195 3626 2361
rect 3618 2189 3619 2195
rect 3625 2189 3626 2195
rect 3618 2027 3626 2189
rect 3618 2021 3619 2027
rect 3625 2021 3626 2027
rect 3618 1875 3626 2021
rect 3618 1869 3619 1875
rect 3625 1869 3626 1875
rect 3618 1707 3626 1869
rect 3618 1701 3619 1707
rect 3625 1701 3626 1707
rect 3618 1547 3626 1701
rect 3618 1541 3619 1547
rect 3625 1541 3626 1547
rect 3618 1391 3626 1541
rect 3618 1385 3619 1391
rect 3625 1385 3626 1391
rect 3618 1223 3626 1385
rect 3618 1217 3619 1223
rect 3625 1217 3626 1223
rect 3618 1063 3626 1217
rect 3618 1057 3619 1063
rect 3625 1057 3626 1063
rect 3618 895 3626 1057
rect 3618 889 3619 895
rect 3625 889 3626 895
rect 3618 743 3626 889
rect 3618 737 3619 743
rect 3625 737 3626 743
rect 3618 591 3626 737
rect 3618 585 3619 591
rect 3625 585 3626 591
rect 3618 427 3626 585
rect 3618 421 3619 427
rect 3625 421 3626 427
rect 3618 267 3626 421
rect 3618 261 3619 267
rect 3625 261 3626 267
rect 3618 103 3626 261
rect 3618 97 3619 103
rect 3625 97 3626 103
rect 3618 72 3626 97
rect 3630 3603 3638 3672
rect 3630 3597 3631 3603
rect 3637 3597 3638 3603
rect 3630 3275 3638 3597
rect 3630 3269 3631 3275
rect 3637 3269 3638 3275
rect 3630 3103 3638 3269
rect 3630 3097 3631 3103
rect 3637 3097 3638 3103
rect 3630 2943 3638 3097
rect 3630 2937 3631 2943
rect 3637 2937 3638 2943
rect 3630 2775 3638 2937
rect 3630 2769 3631 2775
rect 3637 2769 3638 2775
rect 3630 2615 3638 2769
rect 3630 2609 3631 2615
rect 3637 2609 3638 2615
rect 3630 2451 3638 2609
rect 3630 2445 3631 2451
rect 3637 2445 3638 2451
rect 3630 2291 3638 2445
rect 3630 2285 3631 2291
rect 3637 2285 3638 2291
rect 3630 2107 3638 2285
rect 3630 2101 3631 2107
rect 3637 2101 3638 2107
rect 3630 1951 3638 2101
rect 3630 1945 3631 1951
rect 3637 1945 3638 1951
rect 3630 1787 3638 1945
rect 3630 1781 3631 1787
rect 3637 1781 3638 1787
rect 3630 1627 3638 1781
rect 3630 1621 3631 1627
rect 3637 1621 3638 1627
rect 3630 1467 3638 1621
rect 3630 1461 3631 1467
rect 3637 1461 3638 1467
rect 3630 1303 3638 1461
rect 3630 1297 3631 1303
rect 3637 1297 3638 1303
rect 3630 1139 3638 1297
rect 3630 1133 3631 1139
rect 3637 1133 3638 1139
rect 3630 983 3638 1133
rect 3630 977 3631 983
rect 3637 977 3638 983
rect 3630 819 3638 977
rect 3630 813 3631 819
rect 3637 813 3638 819
rect 3630 667 3638 813
rect 3630 661 3631 667
rect 3637 661 3638 667
rect 3630 507 3638 661
rect 3630 501 3631 507
rect 3637 501 3638 507
rect 3630 347 3638 501
rect 3630 341 3631 347
rect 3637 341 3638 347
rect 3630 179 3638 341
rect 3630 173 3631 179
rect 3637 173 3638 179
rect 3630 72 3638 173
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__173
timestamp 1731220558
transform 1 0 3584 0 1 3544
box 7 3 12 24
use welltap_svt  __well_tap__172
timestamp 1731220558
transform 1 0 1864 0 1 3544
box 7 3 12 24
use welltap_svt  __well_tap__171
timestamp 1731220558
transform 1 0 3584 0 -1 3504
box 7 3 12 24
use welltap_svt  __well_tap__170
timestamp 1731220558
transform 1 0 1864 0 -1 3504
box 7 3 12 24
use welltap_svt  __well_tap__169
timestamp 1731220558
transform 1 0 3584 0 1 3384
box 7 3 12 24
use welltap_svt  __well_tap__168
timestamp 1731220558
transform 1 0 1864 0 1 3384
box 7 3 12 24
use welltap_svt  __well_tap__167
timestamp 1731220558
transform 1 0 3584 0 -1 3340
box 7 3 12 24
use welltap_svt  __well_tap__166
timestamp 1731220558
transform 1 0 1864 0 -1 3340
box 7 3 12 24
use welltap_svt  __well_tap__165
timestamp 1731220558
transform 1 0 3584 0 1 3216
box 7 3 12 24
use welltap_svt  __well_tap__164
timestamp 1731220558
transform 1 0 1864 0 1 3216
box 7 3 12 24
use welltap_svt  __well_tap__163
timestamp 1731220558
transform 1 0 3584 0 -1 3172
box 7 3 12 24
use welltap_svt  __well_tap__162
timestamp 1731220558
transform 1 0 1864 0 -1 3172
box 7 3 12 24
use welltap_svt  __well_tap__161
timestamp 1731220558
transform 1 0 3584 0 1 3044
box 7 3 12 24
use welltap_svt  __well_tap__160
timestamp 1731220558
transform 1 0 1864 0 1 3044
box 7 3 12 24
use welltap_svt  __well_tap__159
timestamp 1731220558
transform 1 0 3584 0 -1 2996
box 7 3 12 24
use welltap_svt  __well_tap__158
timestamp 1731220558
transform 1 0 1864 0 -1 2996
box 7 3 12 24
use welltap_svt  __well_tap__157
timestamp 1731220558
transform 1 0 3584 0 1 2884
box 7 3 12 24
use welltap_svt  __well_tap__156
timestamp 1731220558
transform 1 0 1864 0 1 2884
box 7 3 12 24
use welltap_svt  __well_tap__155
timestamp 1731220558
transform 1 0 3584 0 -1 2836
box 7 3 12 24
use welltap_svt  __well_tap__154
timestamp 1731220558
transform 1 0 1864 0 -1 2836
box 7 3 12 24
use welltap_svt  __well_tap__153
timestamp 1731220558
transform 1 0 3584 0 1 2716
box 7 3 12 24
use welltap_svt  __well_tap__152
timestamp 1731220558
transform 1 0 1864 0 1 2716
box 7 3 12 24
use welltap_svt  __well_tap__151
timestamp 1731220558
transform 1 0 3584 0 -1 2676
box 7 3 12 24
use welltap_svt  __well_tap__150
timestamp 1731220558
transform 1 0 1864 0 -1 2676
box 7 3 12 24
use welltap_svt  __well_tap__149
timestamp 1731220558
transform 1 0 3584 0 1 2556
box 7 3 12 24
use welltap_svt  __well_tap__148
timestamp 1731220558
transform 1 0 1864 0 1 2556
box 7 3 12 24
use welltap_svt  __well_tap__147
timestamp 1731220558
transform 1 0 3584 0 -1 2508
box 7 3 12 24
use welltap_svt  __well_tap__146
timestamp 1731220558
transform 1 0 1864 0 -1 2508
box 7 3 12 24
use welltap_svt  __well_tap__145
timestamp 1731220558
transform 1 0 3584 0 1 2392
box 7 3 12 24
use welltap_svt  __well_tap__144
timestamp 1731220558
transform 1 0 1864 0 1 2392
box 7 3 12 24
use welltap_svt  __well_tap__143
timestamp 1731220558
transform 1 0 3584 0 -1 2344
box 7 3 12 24
use welltap_svt  __well_tap__142
timestamp 1731220558
transform 1 0 1864 0 -1 2344
box 7 3 12 24
use welltap_svt  __well_tap__141
timestamp 1731220558
transform 1 0 3584 0 1 2232
box 7 3 12 24
use welltap_svt  __well_tap__140
timestamp 1731220558
transform 1 0 1864 0 1 2232
box 7 3 12 24
use welltap_svt  __well_tap__139
timestamp 1731220558
transform 1 0 3584 0 -1 2172
box 7 3 12 24
use welltap_svt  __well_tap__138
timestamp 1731220558
transform 1 0 1864 0 -1 2172
box 7 3 12 24
use welltap_svt  __well_tap__137
timestamp 1731220558
transform 1 0 3584 0 1 2048
box 7 3 12 24
use welltap_svt  __well_tap__136
timestamp 1731220558
transform 1 0 1864 0 1 2048
box 7 3 12 24
use welltap_svt  __well_tap__135
timestamp 1731220558
transform 1 0 3584 0 -1 2004
box 7 3 12 24
use welltap_svt  __well_tap__134
timestamp 1731220558
transform 1 0 1864 0 -1 2004
box 7 3 12 24
use welltap_svt  __well_tap__133
timestamp 1731220558
transform 1 0 3584 0 1 1892
box 7 3 12 24
use welltap_svt  __well_tap__132
timestamp 1731220558
transform 1 0 1864 0 1 1892
box 7 3 12 24
use welltap_svt  __well_tap__131
timestamp 1731220558
transform 1 0 3584 0 -1 1852
box 7 3 12 24
use welltap_svt  __well_tap__130
timestamp 1731220558
transform 1 0 1864 0 -1 1852
box 7 3 12 24
use welltap_svt  __well_tap__129
timestamp 1731220558
transform 1 0 3584 0 1 1728
box 7 3 12 24
use welltap_svt  __well_tap__128
timestamp 1731220558
transform 1 0 1864 0 1 1728
box 7 3 12 24
use welltap_svt  __well_tap__127
timestamp 1731220558
transform 1 0 3584 0 -1 1684
box 7 3 12 24
use welltap_svt  __well_tap__126
timestamp 1731220558
transform 1 0 1864 0 -1 1684
box 7 3 12 24
use welltap_svt  __well_tap__125
timestamp 1731220558
transform 1 0 3584 0 1 1568
box 7 3 12 24
use welltap_svt  __well_tap__124
timestamp 1731220558
transform 1 0 1864 0 1 1568
box 7 3 12 24
use welltap_svt  __well_tap__123
timestamp 1731220558
transform 1 0 3584 0 -1 1524
box 7 3 12 24
use welltap_svt  __well_tap__122
timestamp 1731220558
transform 1 0 1864 0 -1 1524
box 7 3 12 24
use welltap_svt  __well_tap__121
timestamp 1731220558
transform 1 0 3584 0 1 1408
box 7 3 12 24
use welltap_svt  __well_tap__120
timestamp 1731220558
transform 1 0 1864 0 1 1408
box 7 3 12 24
use welltap_svt  __well_tap__119
timestamp 1731220558
transform 1 0 3584 0 -1 1368
box 7 3 12 24
use welltap_svt  __well_tap__118
timestamp 1731220558
transform 1 0 1864 0 -1 1368
box 7 3 12 24
use welltap_svt  __well_tap__117
timestamp 1731220558
transform 1 0 3584 0 1 1244
box 7 3 12 24
use welltap_svt  __well_tap__116
timestamp 1731220558
transform 1 0 1864 0 1 1244
box 7 3 12 24
use welltap_svt  __well_tap__115
timestamp 1731220558
transform 1 0 3584 0 -1 1200
box 7 3 12 24
use welltap_svt  __well_tap__114
timestamp 1731220558
transform 1 0 1864 0 -1 1200
box 7 3 12 24
use welltap_svt  __well_tap__113
timestamp 1731220558
transform 1 0 3584 0 1 1080
box 7 3 12 24
use welltap_svt  __well_tap__112
timestamp 1731220558
transform 1 0 1864 0 1 1080
box 7 3 12 24
use welltap_svt  __well_tap__111
timestamp 1731220558
transform 1 0 3584 0 -1 1040
box 7 3 12 24
use welltap_svt  __well_tap__110
timestamp 1731220558
transform 1 0 1864 0 -1 1040
box 7 3 12 24
use welltap_svt  __well_tap__109
timestamp 1731220558
transform 1 0 3584 0 1 924
box 7 3 12 24
use welltap_svt  __well_tap__108
timestamp 1731220558
transform 1 0 1864 0 1 924
box 7 3 12 24
use welltap_svt  __well_tap__107
timestamp 1731220558
transform 1 0 3584 0 -1 872
box 7 3 12 24
use welltap_svt  __well_tap__106
timestamp 1731220558
transform 1 0 1864 0 -1 872
box 7 3 12 24
use welltap_svt  __well_tap__105
timestamp 1731220558
transform 1 0 3584 0 1 760
box 7 3 12 24
use welltap_svt  __well_tap__104
timestamp 1731220558
transform 1 0 1864 0 1 760
box 7 3 12 24
use welltap_svt  __well_tap__103
timestamp 1731220558
transform 1 0 3584 0 -1 720
box 7 3 12 24
use welltap_svt  __well_tap__102
timestamp 1731220558
transform 1 0 1864 0 -1 720
box 7 3 12 24
use welltap_svt  __well_tap__101
timestamp 1731220558
transform 1 0 3584 0 1 608
box 7 3 12 24
use welltap_svt  __well_tap__100
timestamp 1731220558
transform 1 0 1864 0 1 608
box 7 3 12 24
use welltap_svt  __well_tap__99
timestamp 1731220558
transform 1 0 3584 0 -1 568
box 7 3 12 24
use welltap_svt  __well_tap__98
timestamp 1731220558
transform 1 0 1864 0 -1 568
box 7 3 12 24
use welltap_svt  __well_tap__97
timestamp 1731220558
transform 1 0 3584 0 1 448
box 7 3 12 24
use welltap_svt  __well_tap__96
timestamp 1731220558
transform 1 0 1864 0 1 448
box 7 3 12 24
use welltap_svt  __well_tap__95
timestamp 1731220558
transform 1 0 3584 0 -1 404
box 7 3 12 24
use welltap_svt  __well_tap__94
timestamp 1731220558
transform 1 0 1864 0 -1 404
box 7 3 12 24
use welltap_svt  __well_tap__93
timestamp 1731220558
transform 1 0 3584 0 1 288
box 7 3 12 24
use welltap_svt  __well_tap__92
timestamp 1731220558
transform 1 0 1864 0 1 288
box 7 3 12 24
use welltap_svt  __well_tap__91
timestamp 1731220558
transform 1 0 3584 0 -1 244
box 7 3 12 24
use welltap_svt  __well_tap__90
timestamp 1731220558
transform 1 0 1864 0 -1 244
box 7 3 12 24
use welltap_svt  __well_tap__89
timestamp 1731220558
transform 1 0 3584 0 1 120
box 7 3 12 24
use welltap_svt  __well_tap__88
timestamp 1731220558
transform 1 0 1864 0 1 120
box 7 3 12 24
use welltap_svt  __well_tap__87
timestamp 1731220558
transform 1 0 1824 0 -1 3648
box 7 3 12 24
use welltap_svt  __well_tap__86
timestamp 1731220558
transform 1 0 104 0 -1 3648
box 7 3 12 24
use welltap_svt  __well_tap__85
timestamp 1731220558
transform 1 0 1824 0 1 3536
box 7 3 12 24
use welltap_svt  __well_tap__84
timestamp 1731220558
transform 1 0 104 0 1 3536
box 7 3 12 24
use welltap_svt  __well_tap__83
timestamp 1731220558
transform 1 0 1824 0 -1 3496
box 7 3 12 24
use welltap_svt  __well_tap__82
timestamp 1731220558
transform 1 0 104 0 -1 3496
box 7 3 12 24
use welltap_svt  __well_tap__81
timestamp 1731220558
transform 1 0 1824 0 1 3384
box 7 3 12 24
use welltap_svt  __well_tap__80
timestamp 1731220558
transform 1 0 104 0 1 3384
box 7 3 12 24
use welltap_svt  __well_tap__79
timestamp 1731220558
transform 1 0 1824 0 -1 3344
box 7 3 12 24
use welltap_svt  __well_tap__78
timestamp 1731220558
transform 1 0 104 0 -1 3344
box 7 3 12 24
use welltap_svt  __well_tap__77
timestamp 1731220558
transform 1 0 1824 0 1 3228
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220558
transform 1 0 104 0 1 3228
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220558
transform 1 0 1824 0 -1 3188
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220558
transform 1 0 104 0 -1 3188
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220558
transform 1 0 1824 0 1 3072
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220558
transform 1 0 104 0 1 3072
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220558
transform 1 0 1824 0 -1 3028
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220558
transform 1 0 104 0 -1 3028
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220558
transform 1 0 1824 0 1 2916
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220558
transform 1 0 104 0 1 2916
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220558
transform 1 0 1824 0 -1 2876
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220558
transform 1 0 104 0 -1 2876
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220558
transform 1 0 1824 0 1 2764
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220558
transform 1 0 104 0 1 2764
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220558
transform 1 0 1824 0 -1 2720
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220558
transform 1 0 104 0 -1 2720
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220558
transform 1 0 1824 0 1 2608
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220558
transform 1 0 104 0 1 2608
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220558
transform 1 0 1824 0 -1 2564
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220558
transform 1 0 104 0 -1 2564
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220558
transform 1 0 1824 0 1 2448
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220558
transform 1 0 104 0 1 2448
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220558
transform 1 0 1824 0 -1 2400
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220558
transform 1 0 104 0 -1 2400
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220558
transform 1 0 1824 0 1 2288
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220558
transform 1 0 104 0 1 2288
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220558
transform 1 0 1824 0 -1 2240
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220558
transform 1 0 104 0 -1 2240
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220558
transform 1 0 1824 0 1 2124
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220558
transform 1 0 104 0 1 2124
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220558
transform 1 0 1824 0 -1 2080
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220558
transform 1 0 104 0 -1 2080
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220558
transform 1 0 1824 0 1 1968
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220558
transform 1 0 104 0 1 1968
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220558
transform 1 0 1824 0 -1 1920
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220558
transform 1 0 104 0 -1 1920
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220558
transform 1 0 1824 0 1 1808
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220558
transform 1 0 104 0 1 1808
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220558
transform 1 0 1824 0 -1 1764
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220558
transform 1 0 104 0 -1 1764
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220558
transform 1 0 1824 0 1 1648
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220558
transform 1 0 104 0 1 1648
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220558
transform 1 0 1824 0 -1 1600
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220558
transform 1 0 104 0 -1 1600
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220558
transform 1 0 1824 0 1 1484
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220558
transform 1 0 104 0 1 1484
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220558
transform 1 0 1824 0 -1 1440
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220558
transform 1 0 104 0 -1 1440
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220558
transform 1 0 1824 0 1 1312
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220558
transform 1 0 104 0 1 1312
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220558
transform 1 0 1824 0 -1 1268
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220558
transform 1 0 104 0 -1 1268
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220558
transform 1 0 1824 0 1 1148
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220558
transform 1 0 104 0 1 1148
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220558
transform 1 0 1824 0 -1 1108
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220558
transform 1 0 104 0 -1 1108
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220558
transform 1 0 1824 0 1 984
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220558
transform 1 0 104 0 1 984
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220558
transform 1 0 1824 0 -1 932
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220558
transform 1 0 104 0 -1 932
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220558
transform 1 0 1824 0 1 816
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220558
transform 1 0 104 0 1 816
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220558
transform 1 0 1824 0 -1 764
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220558
transform 1 0 104 0 -1 764
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220558
transform 1 0 1824 0 1 644
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220558
transform 1 0 104 0 1 644
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220558
transform 1 0 1824 0 -1 596
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220558
transform 1 0 104 0 -1 596
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220558
transform 1 0 1824 0 1 472
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220558
transform 1 0 104 0 1 472
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220558
transform 1 0 1824 0 -1 424
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220558
transform 1 0 104 0 -1 424
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220558
transform 1 0 1824 0 1 300
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220558
transform 1 0 104 0 1 300
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220558
transform 1 0 1824 0 -1 252
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220558
transform 1 0 104 0 -1 252
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220558
transform 1 0 1824 0 1 104
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220558
transform 1 0 104 0 1 104
box 7 3 12 24
use _0_0std_0_0cells_0_0LATCHINV  tst_5999_6
timestamp 1731220558
transform 1 0 3416 0 1 100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5998_6
timestamp 1731220558
transform 1 0 3496 0 1 100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5997_6
timestamp 1731220558
transform 1 0 3496 0 -1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5996_6
timestamp 1731220558
transform 1 0 3496 0 1 268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5995_6
timestamp 1731220558
transform 1 0 3488 0 -1 424
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5994_6
timestamp 1731220558
transform 1 0 3456 0 1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5993_6
timestamp 1731220558
transform 1 0 3296 0 -1 424
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5992_6
timestamp 1731220558
transform 1 0 3376 0 1 268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5991_6
timestamp 1731220558
transform 1 0 3240 0 1 268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5990_6
timestamp 1731220558
transform 1 0 3104 0 1 268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5989_6
timestamp 1731220558
transform 1 0 3088 0 -1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5988_6
timestamp 1731220558
transform 1 0 3232 0 -1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5987_6
timestamp 1731220558
transform 1 0 3376 0 -1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5986_6
timestamp 1731220558
transform 1 0 3328 0 1 100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5985_6
timestamp 1731220558
transform 1 0 3232 0 1 100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5984_6
timestamp 1731220558
transform 1 0 3144 0 1 100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5983_6
timestamp 1731220558
transform 1 0 3048 0 1 100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5982_6
timestamp 1731220558
transform 1 0 2944 0 1 100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5981_6
timestamp 1731220558
transform 1 0 2840 0 1 100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5980_6
timestamp 1731220558
transform 1 0 2728 0 1 100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5979_6
timestamp 1731220558
transform 1 0 2608 0 1 100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5978_6
timestamp 1731220558
transform 1 0 2672 0 -1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5977_6
timestamp 1731220558
transform 1 0 2808 0 -1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5976_6
timestamp 1731220558
transform 1 0 2944 0 -1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5975_6
timestamp 1731220558
transform 1 0 2832 0 1 268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5974_6
timestamp 1731220558
transform 1 0 2968 0 1 268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5973_6
timestamp 1731220558
transform 1 0 3104 0 -1 424
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5972_6
timestamp 1731220558
transform 1 0 2920 0 -1 424
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5971_6
timestamp 1731220558
transform 1 0 2752 0 -1 424
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5970_6
timestamp 1731220558
transform 1 0 2600 0 -1 424
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5969_6
timestamp 1731220558
transform 1 0 2464 0 -1 424
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5968_6
timestamp 1731220558
transform 1 0 2568 0 1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5967_6
timestamp 1731220558
transform 1 0 2672 0 1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5966_6
timestamp 1731220558
transform 1 0 2952 0 -1 588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5965_6
timestamp 1731220558
transform 1 0 2808 0 -1 588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5964_6
timestamp 1731220558
transform 1 0 2720 0 1 588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5963_6
timestamp 1731220558
transform 1 0 2896 0 -1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5962_6
timestamp 1731220558
transform 1 0 2792 0 1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5961_6
timestamp 1731220558
transform 1 0 3072 0 -1 892
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5960_6
timestamp 1731220558
transform 1 0 3296 0 -1 892
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5959_6
timestamp 1731220558
transform 1 0 3136 0 1 904
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5958_6
timestamp 1731220558
transform 1 0 3328 0 1 904
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5957_6
timestamp 1731220558
transform 1 0 3368 0 -1 1060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5956_6
timestamp 1731220558
transform 1 0 3216 0 -1 1060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5955_6
timestamp 1731220558
transform 1 0 3144 0 1 1060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5954_6
timestamp 1731220558
transform 1 0 3328 0 1 1060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5953_6
timestamp 1731220558
transform 1 0 3192 0 -1 1220
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5952_6
timestamp 1731220558
transform 1 0 3336 0 -1 1220
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5951_6
timestamp 1731220558
transform 1 0 3352 0 1 1224
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5950_6
timestamp 1731220558
transform 1 0 3200 0 1 1224
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5949_6
timestamp 1731220558
transform 1 0 3152 0 -1 1388
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5948_6
timestamp 1731220558
transform 1 0 3272 0 -1 1388
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5947_6
timestamp 1731220558
transform 1 0 3392 0 -1 1388
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5946_6
timestamp 1731220558
transform 1 0 3464 0 1 1388
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5945_6
timestamp 1731220558
transform 1 0 3488 0 -1 1544
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5944_6
timestamp 1731220558
transform 1 0 3496 0 -1 1704
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5943_6
timestamp 1731220558
transform 1 0 3496 0 1 1708
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5942_6
timestamp 1731220558
transform 1 0 3496 0 -1 1872
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5941_6
timestamp 1731220558
transform 1 0 3496 0 1 1548
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5940_6
timestamp 1731220558
transform 1 0 3496 0 -1 1388
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5939_6
timestamp 1731220558
transform 1 0 3496 0 1 1224
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5938_6
timestamp 1731220558
transform 1 0 3488 0 -1 1220
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5937_6
timestamp 1731220558
transform 1 0 3496 0 1 1060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5936_6
timestamp 1731220558
transform 1 0 3496 0 -1 1060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5935_6
timestamp 1731220558
transform 1 0 3496 0 1 904
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5934_6
timestamp 1731220558
transform 1 0 3496 0 -1 892
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5933_6
timestamp 1731220558
transform 1 0 3496 0 1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5932_6
timestamp 1731220558
transform 1 0 3496 0 -1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5931_6
timestamp 1731220558
transform 1 0 3496 0 1 588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5930_6
timestamp 1731220558
transform 1 0 3440 0 -1 588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5929_6
timestamp 1731220558
transform 1 0 3360 0 1 588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5928_6
timestamp 1731220558
transform 1 0 3232 0 1 588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5927_6
timestamp 1731220558
transform 1 0 3200 0 -1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5926_6
timestamp 1731220558
transform 1 0 3352 0 -1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5925_6
timestamp 1731220558
transform 1 0 3376 0 1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5924_6
timestamp 1731220558
transform 1 0 3232 0 1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5923_6
timestamp 1731220558
transform 1 0 3088 0 1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5922_6
timestamp 1731220558
transform 1 0 2944 0 1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5921_6
timestamp 1731220558
transform 1 0 3048 0 -1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5920_6
timestamp 1731220558
transform 1 0 3104 0 1 588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5919_6
timestamp 1731220558
transform 1 0 3272 0 -1 588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5918_6
timestamp 1731220558
transform 1 0 3304 0 1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5917_6
timestamp 1731220558
transform 1 0 3160 0 1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5916_6
timestamp 1731220558
transform 1 0 3024 0 1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5915_6
timestamp 1731220558
transform 1 0 2896 0 1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5914_6
timestamp 1731220558
transform 1 0 2776 0 1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5913_6
timestamp 1731220558
transform 1 0 3104 0 -1 588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5912_6
timestamp 1731220558
transform 1 0 2976 0 1 588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5911_6
timestamp 1731220558
transform 1 0 2848 0 1 588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5910_6
timestamp 1731220558
transform 1 0 2744 0 -1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5909_6
timestamp 1731220558
transform 1 0 2632 0 1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5908_6
timestamp 1731220558
transform 1 0 2448 0 -1 892
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5907_6
timestamp 1731220558
transform 1 0 2648 0 -1 892
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5906_6
timestamp 1731220558
transform 1 0 2856 0 -1 892
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5905_6
timestamp 1731220558
transform 1 0 2952 0 1 904
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5904_6
timestamp 1731220558
transform 1 0 2776 0 1 904
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5903_6
timestamp 1731220558
transform 1 0 2616 0 1 904
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5902_6
timestamp 1731220558
transform 1 0 2632 0 -1 1060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5901_6
timestamp 1731220558
transform 1 0 2784 0 -1 1060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5900_6
timestamp 1731220558
transform 1 0 2928 0 -1 1060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5899_6
timestamp 1731220558
transform 1 0 3072 0 -1 1060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5898_6
timestamp 1731220558
transform 1 0 2952 0 1 1060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5897_6
timestamp 1731220558
transform 1 0 2760 0 1 1060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5896_6
timestamp 1731220558
transform 1 0 2560 0 1 1060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5895_6
timestamp 1731220558
transform 1 0 3048 0 -1 1220
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5894_6
timestamp 1731220558
transform 1 0 2904 0 -1 1220
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5893_6
timestamp 1731220558
transform 1 0 2768 0 -1 1220
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5892_6
timestamp 1731220558
transform 1 0 2640 0 -1 1220
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5891_6
timestamp 1731220558
transform 1 0 2776 0 1 1224
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5890_6
timestamp 1731220558
transform 1 0 2912 0 1 1224
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5889_6
timestamp 1731220558
transform 1 0 3056 0 1 1224
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5888_6
timestamp 1731220558
transform 1 0 3032 0 -1 1388
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5887_6
timestamp 1731220558
transform 1 0 2912 0 -1 1388
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5886_6
timestamp 1731220558
transform 1 0 2496 0 -1 1388
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5885_6
timestamp 1731220558
transform 1 0 2336 0 -1 1388
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5884_6
timestamp 1731220558
transform 1 0 2256 0 -1 1388
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5883_6
timestamp 1731220558
transform 1 0 2800 0 -1 1388
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5882_6
timestamp 1731220558
transform 1 0 2688 0 -1 1388
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5881_6
timestamp 1731220558
transform 1 0 2584 0 -1 1388
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5880_6
timestamp 1731220558
transform 1 0 2592 0 1 1388
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5879_6
timestamp 1731220558
transform 1 0 2720 0 1 1388
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5878_6
timestamp 1731220558
transform 1 0 3264 0 1 1388
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5877_6
timestamp 1731220558
transform 1 0 3064 0 1 1388
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5876_6
timestamp 1731220558
transform 1 0 2880 0 1 1388
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5875_6
timestamp 1731220558
transform 1 0 2776 0 -1 1544
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5874_6
timestamp 1731220558
transform 1 0 2640 0 -1 1544
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5873_6
timestamp 1731220558
transform 1 0 3296 0 -1 1544
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5872_6
timestamp 1731220558
transform 1 0 3112 0 -1 1544
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5871_6
timestamp 1731220558
transform 1 0 2936 0 -1 1544
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5870_6
timestamp 1731220558
transform 1 0 2896 0 1 1548
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5869_6
timestamp 1731220558
transform 1 0 2760 0 1 1548
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5868_6
timestamp 1731220558
transform 1 0 2624 0 1 1548
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5867_6
timestamp 1731220558
transform 1 0 3040 0 1 1548
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5866_6
timestamp 1731220558
transform 1 0 3352 0 1 1548
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5865_6
timestamp 1731220558
transform 1 0 3192 0 1 1548
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5864_6
timestamp 1731220558
transform 1 0 3104 0 -1 1704
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5863_6
timestamp 1731220558
transform 1 0 2960 0 -1 1704
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5862_6
timestamp 1731220558
transform 1 0 2808 0 -1 1704
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5861_6
timestamp 1731220558
transform 1 0 3240 0 -1 1704
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5860_6
timestamp 1731220558
transform 1 0 3376 0 -1 1704
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5859_6
timestamp 1731220558
transform 1 0 3376 0 1 1708
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5858_6
timestamp 1731220558
transform 1 0 3240 0 1 1708
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5857_6
timestamp 1731220558
transform 1 0 3104 0 1 1708
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5856_6
timestamp 1731220558
transform 1 0 2968 0 1 1708
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5855_6
timestamp 1731220558
transform 1 0 2824 0 1 1708
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5854_6
timestamp 1731220558
transform 1 0 2672 0 1 1708
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5853_6
timestamp 1731220558
transform 1 0 3328 0 -1 1872
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5852_6
timestamp 1731220558
transform 1 0 3144 0 -1 1872
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5851_6
timestamp 1731220558
transform 1 0 2968 0 -1 1872
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5850_6
timestamp 1731220558
transform 1 0 2800 0 -1 1872
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5849_6
timestamp 1731220558
transform 1 0 2648 0 -1 1872
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5848_6
timestamp 1731220558
transform 1 0 2512 0 -1 1872
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5847_6
timestamp 1731220558
transform 1 0 2824 0 1 1872
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5846_6
timestamp 1731220558
transform 1 0 2704 0 1 1872
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5845_6
timestamp 1731220558
transform 1 0 2584 0 1 1872
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5844_6
timestamp 1731220558
transform 1 0 2472 0 1 1872
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5843_6
timestamp 1731220558
transform 1 0 2360 0 1 1872
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5842_6
timestamp 1731220558
transform 1 0 2672 0 -1 2024
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5841_6
timestamp 1731220558
transform 1 0 2840 0 -1 2024
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5840_6
timestamp 1731220558
transform 1 0 3008 0 -1 2024
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5839_6
timestamp 1731220558
transform 1 0 3064 0 1 2028
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5838_6
timestamp 1731220558
transform 1 0 2952 0 1 2028
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5837_6
timestamp 1731220558
transform 1 0 2832 0 1 2028
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5836_6
timestamp 1731220558
transform 1 0 2872 0 -1 2192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5835_6
timestamp 1731220558
transform 1 0 2984 0 -1 2192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5834_6
timestamp 1731220558
transform 1 0 3088 0 -1 2192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5833_6
timestamp 1731220558
transform 1 0 3192 0 -1 2192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5832_6
timestamp 1731220558
transform 1 0 3296 0 -1 2192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5831_6
timestamp 1731220558
transform 1 0 3288 0 1 2028
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5830_6
timestamp 1731220558
transform 1 0 3176 0 1 2028
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5829_6
timestamp 1731220558
transform 1 0 3400 0 1 2028
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5828_6
timestamp 1731220558
transform 1 0 3344 0 -1 2024
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5827_6
timestamp 1731220558
transform 1 0 3176 0 -1 2024
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5826_6
timestamp 1731220558
transform 1 0 3496 0 -1 2024
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5825_6
timestamp 1731220558
transform 1 0 3496 0 1 2028
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5824_6
timestamp 1731220558
transform 1 0 3496 0 -1 2192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5823_6
timestamp 1731220558
transform 1 0 3400 0 -1 2192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5822_6
timestamp 1731220558
transform 1 0 3240 0 1 2212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5821_6
timestamp 1731220558
transform 1 0 3008 0 1 2212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5820_6
timestamp 1731220558
transform 1 0 3480 0 1 2212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5819_6
timestamp 1731220558
transform 1 0 3496 0 -1 2364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5818_6
timestamp 1731220558
transform 1 0 3408 0 -1 2364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5817_6
timestamp 1731220558
transform 1 0 3296 0 -1 2364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5816_6
timestamp 1731220558
transform 1 0 3184 0 -1 2364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5815_6
timestamp 1731220558
transform 1 0 3072 0 -1 2364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5814_6
timestamp 1731220558
transform 1 0 2952 0 -1 2364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5813_6
timestamp 1731220558
transform 1 0 2816 0 -1 2364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5812_6
timestamp 1731220558
transform 1 0 2664 0 -1 2364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5811_6
timestamp 1731220558
transform 1 0 3200 0 1 2372
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5810_6
timestamp 1731220558
transform 1 0 3064 0 1 2372
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5809_6
timestamp 1731220558
transform 1 0 2928 0 1 2372
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5808_6
timestamp 1731220558
transform 1 0 2792 0 1 2372
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5807_6
timestamp 1731220558
transform 1 0 2656 0 1 2372
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5806_6
timestamp 1731220558
transform 1 0 3072 0 -1 2528
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5805_6
timestamp 1731220558
transform 1 0 2968 0 -1 2528
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5804_6
timestamp 1731220558
transform 1 0 2872 0 -1 2528
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5803_6
timestamp 1731220558
transform 1 0 2776 0 -1 2528
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5802_6
timestamp 1731220558
transform 1 0 2680 0 -1 2528
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5801_6
timestamp 1731220558
transform 1 0 2584 0 -1 2528
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5800_6
timestamp 1731220558
transform 1 0 2976 0 1 2536
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5799_6
timestamp 1731220558
transform 1 0 2896 0 1 2536
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5798_6
timestamp 1731220558
transform 1 0 2816 0 1 2536
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5797_6
timestamp 1731220558
transform 1 0 2736 0 1 2536
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5796_6
timestamp 1731220558
transform 1 0 2656 0 1 2536
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5795_6
timestamp 1731220558
transform 1 0 2632 0 -1 2696
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5794_6
timestamp 1731220558
transform 1 0 2712 0 -1 2696
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5793_6
timestamp 1731220558
transform 1 0 2952 0 -1 2696
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5792_6
timestamp 1731220558
transform 1 0 2872 0 -1 2696
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5791_6
timestamp 1731220558
transform 1 0 2792 0 -1 2696
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5790_6
timestamp 1731220558
transform 1 0 2712 0 1 2696
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5789_6
timestamp 1731220558
transform 1 0 2624 0 1 2696
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5788_6
timestamp 1731220558
transform 1 0 2976 0 1 2696
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5787_6
timestamp 1731220558
transform 1 0 2888 0 1 2696
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5786_6
timestamp 1731220558
transform 1 0 2800 0 1 2696
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5785_6
timestamp 1731220558
transform 1 0 2760 0 -1 2856
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5784_6
timestamp 1731220558
transform 1 0 2640 0 -1 2856
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5783_6
timestamp 1731220558
transform 1 0 3128 0 -1 2856
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5782_6
timestamp 1731220558
transform 1 0 3000 0 -1 2856
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5781_6
timestamp 1731220558
transform 1 0 2880 0 -1 2856
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5780_6
timestamp 1731220558
transform 1 0 2824 0 1 2864
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5779_6
timestamp 1731220558
transform 1 0 2656 0 1 2864
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5778_6
timestamp 1731220558
transform 1 0 3288 0 1 2864
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5777_6
timestamp 1731220558
transform 1 0 3136 0 1 2864
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5776_6
timestamp 1731220558
transform 1 0 2984 0 1 2864
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5775_6
timestamp 1731220558
transform 1 0 2808 0 -1 3016
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5774_6
timestamp 1731220558
transform 1 0 2680 0 -1 3016
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5773_6
timestamp 1731220558
transform 1 0 2536 0 -1 3016
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5772_6
timestamp 1731220558
transform 1 0 2920 0 -1 3016
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5771_6
timestamp 1731220558
transform 1 0 3032 0 -1 3016
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5770_6
timestamp 1731220558
transform 1 0 3136 0 -1 3016
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5769_6
timestamp 1731220558
transform 1 0 3232 0 -1 3016
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5768_6
timestamp 1731220558
transform 1 0 3440 0 1 2864
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5767_6
timestamp 1731220558
transform 1 0 3416 0 -1 3016
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5766_6
timestamp 1731220558
transform 1 0 3328 0 -1 3016
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5765_6
timestamp 1731220558
transform 1 0 3496 0 -1 3016
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5764_6
timestamp 1731220558
transform 1 0 3496 0 1 3024
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5763_6
timestamp 1731220558
transform 1 0 3216 0 1 3024
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5762_6
timestamp 1731220558
transform 1 0 3480 0 -1 3192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5761_6
timestamp 1731220558
transform 1 0 3360 0 1 3196
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5760_6
timestamp 1731220558
transform 1 0 3496 0 1 3196
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5759_6
timestamp 1731220558
transform 1 0 3464 0 -1 3360
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5758_6
timestamp 1731220558
transform 1 0 3304 0 -1 3360
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5757_6
timestamp 1731220558
transform 1 0 3248 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5756_6
timestamp 1731220558
transform 1 0 3408 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5755_6
timestamp 1731220558
transform 1 0 3368 0 -1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5754_6
timestamp 1731220558
transform 1 0 3240 0 -1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5753_6
timestamp 1731220558
transform 1 0 3112 0 -1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5752_6
timestamp 1731220558
transform 1 0 3384 0 1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5751_6
timestamp 1731220558
transform 1 0 3288 0 1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5750_6
timestamp 1731220558
transform 1 0 3192 0 1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5749_6
timestamp 1731220558
transform 1 0 3096 0 1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5748_6
timestamp 1731220558
transform 1 0 3000 0 1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5747_6
timestamp 1731220558
transform 1 0 2904 0 1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5746_6
timestamp 1731220558
transform 1 0 2800 0 1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5745_6
timestamp 1731220558
transform 1 0 2688 0 1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5744_6
timestamp 1731220558
transform 1 0 2864 0 -1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5743_6
timestamp 1731220558
transform 1 0 2984 0 -1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5742_6
timestamp 1731220558
transform 1 0 2944 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5741_6
timestamp 1731220558
transform 1 0 3096 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5740_6
timestamp 1731220558
transform 1 0 3152 0 -1 3360
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5739_6
timestamp 1731220558
transform 1 0 3000 0 -1 3360
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5738_6
timestamp 1731220558
transform 1 0 2944 0 1 3196
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5737_6
timestamp 1731220558
transform 1 0 3080 0 1 3196
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5736_6
timestamp 1731220558
transform 1 0 3216 0 1 3196
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5735_6
timestamp 1731220558
transform 1 0 3320 0 -1 3192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5734_6
timestamp 1731220558
transform 1 0 3168 0 -1 3192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5733_6
timestamp 1731220558
transform 1 0 3024 0 -1 3192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5732_6
timestamp 1731220558
transform 1 0 2888 0 -1 3192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5731_6
timestamp 1731220558
transform 1 0 2760 0 -1 3192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5730_6
timestamp 1731220558
transform 1 0 2632 0 -1 3192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5729_6
timestamp 1731220558
transform 1 0 2504 0 -1 3192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5728_6
timestamp 1731220558
transform 1 0 2536 0 1 3196
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5727_6
timestamp 1731220558
transform 1 0 2672 0 1 3196
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5726_6
timestamp 1731220558
transform 1 0 2808 0 1 3196
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5725_6
timestamp 1731220558
transform 1 0 2856 0 -1 3360
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5724_6
timestamp 1731220558
transform 1 0 2712 0 -1 3360
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5723_6
timestamp 1731220558
transform 1 0 2576 0 -1 3360
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5722_6
timestamp 1731220558
transform 1 0 2528 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5721_6
timestamp 1731220558
transform 1 0 2664 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5720_6
timestamp 1731220558
transform 1 0 2800 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5719_6
timestamp 1731220558
transform 1 0 2736 0 -1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5718_6
timestamp 1731220558
transform 1 0 2608 0 -1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5717_6
timestamp 1731220558
transform 1 0 2480 0 -1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5716_6
timestamp 1731220558
transform 1 0 2360 0 -1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5715_6
timestamp 1731220558
transform 1 0 2576 0 1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5714_6
timestamp 1731220558
transform 1 0 2464 0 1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5713_6
timestamp 1731220558
transform 1 0 2352 0 1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5712_6
timestamp 1731220558
transform 1 0 2240 0 1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5711_6
timestamp 1731220558
transform 1 0 2136 0 1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5710_6
timestamp 1731220558
transform 1 0 2048 0 1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5709_6
timestamp 1731220558
transform 1 0 2080 0 -1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5708_6
timestamp 1731220558
transform 1 0 2160 0 -1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5707_6
timestamp 1731220558
transform 1 0 2256 0 -1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5706_6
timestamp 1731220558
transform 1 0 2184 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5705_6
timestamp 1731220558
transform 1 0 2096 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5704_6
timestamp 1731220558
transform 1 0 2288 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5703_6
timestamp 1731220558
transform 1 0 2400 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5702_6
timestamp 1731220558
transform 1 0 2448 0 -1 3360
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5701_6
timestamp 1731220558
transform 1 0 2328 0 -1 3360
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5700_6
timestamp 1731220558
transform 1 0 2216 0 -1 3360
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5699_6
timestamp 1731220558
transform 1 0 2120 0 -1 3360
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5698_6
timestamp 1731220558
transform 1 0 2120 0 1 3196
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5697_6
timestamp 1731220558
transform 1 0 2400 0 1 3196
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5696_6
timestamp 1731220558
transform 1 0 2264 0 1 3196
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5695_6
timestamp 1731220558
transform 1 0 2240 0 -1 3192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5694_6
timestamp 1731220558
transform 1 0 2376 0 -1 3192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5693_6
timestamp 1731220558
transform 1 0 2920 0 1 3024
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5692_6
timestamp 1731220558
transform 1 0 2640 0 1 3024
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5691_6
timestamp 1731220558
transform 1 0 2392 0 1 3024
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5690_6
timestamp 1731220558
transform 1 0 2216 0 -1 3016
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5689_6
timestamp 1731220558
transform 1 0 2384 0 -1 3016
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5688_6
timestamp 1731220558
transform 1 0 2472 0 1 2864
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5687_6
timestamp 1731220558
transform 1 0 2280 0 1 2864
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5686_6
timestamp 1731220558
transform 1 0 2072 0 1 2864
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5685_6
timestamp 1731220558
transform 1 0 2128 0 -1 2856
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5684_6
timestamp 1731220558
transform 1 0 2256 0 -1 2856
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5683_6
timestamp 1731220558
transform 1 0 2384 0 -1 2856
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5682_6
timestamp 1731220558
transform 1 0 2512 0 -1 2856
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5681_6
timestamp 1731220558
transform 1 0 2536 0 1 2696
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5680_6
timestamp 1731220558
transform 1 0 2456 0 1 2696
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5679_6
timestamp 1731220558
transform 1 0 2376 0 1 2696
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5678_6
timestamp 1731220558
transform 1 0 2296 0 1 2696
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5677_6
timestamp 1731220558
transform 1 0 2216 0 1 2696
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5676_6
timestamp 1731220558
transform 1 0 2232 0 -1 2696
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5675_6
timestamp 1731220558
transform 1 0 2312 0 -1 2696
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5674_6
timestamp 1731220558
transform 1 0 2392 0 -1 2696
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5673_6
timestamp 1731220558
transform 1 0 2472 0 -1 2696
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5672_6
timestamp 1731220558
transform 1 0 2552 0 -1 2696
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5671_6
timestamp 1731220558
transform 1 0 2576 0 1 2536
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5670_6
timestamp 1731220558
transform 1 0 2496 0 1 2536
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5669_6
timestamp 1731220558
transform 1 0 2416 0 1 2536
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5668_6
timestamp 1731220558
transform 1 0 2336 0 1 2536
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5667_6
timestamp 1731220558
transform 1 0 2256 0 1 2536
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5666_6
timestamp 1731220558
transform 1 0 2176 0 1 2536
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5665_6
timestamp 1731220558
transform 1 0 2488 0 -1 2528
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5664_6
timestamp 1731220558
transform 1 0 2392 0 -1 2528
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5663_6
timestamp 1731220558
transform 1 0 2296 0 -1 2528
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5662_6
timestamp 1731220558
transform 1 0 2200 0 -1 2528
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5661_6
timestamp 1731220558
transform 1 0 2112 0 -1 2528
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5660_6
timestamp 1731220558
transform 1 0 2520 0 1 2372
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5659_6
timestamp 1731220558
transform 1 0 2376 0 1 2372
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5658_6
timestamp 1731220558
transform 1 0 2232 0 1 2372
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5657_6
timestamp 1731220558
transform 1 0 2096 0 1 2372
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5656_6
timestamp 1731220558
transform 1 0 1976 0 1 2372
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5655_6
timestamp 1731220558
transform 1 0 1888 0 1 2372
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5654_6
timestamp 1731220558
transform 1 0 2504 0 -1 2364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5653_6
timestamp 1731220558
transform 1 0 2336 0 -1 2364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5652_6
timestamp 1731220558
transform 1 0 2168 0 -1 2364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5651_6
timestamp 1731220558
transform 1 0 2008 0 -1 2364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5650_6
timestamp 1731220558
transform 1 0 1888 0 -1 2364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5649_6
timestamp 1731220558
transform 1 0 1888 0 1 2212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5648_6
timestamp 1731220558
transform 1 0 2016 0 1 2212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5647_6
timestamp 1731220558
transform 1 0 2168 0 1 2212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5646_6
timestamp 1731220558
transform 1 0 2352 0 1 2212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5645_6
timestamp 1731220558
transform 1 0 2776 0 1 2212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5644_6
timestamp 1731220558
transform 1 0 2560 0 1 2212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5643_6
timestamp 1731220558
transform 1 0 2392 0 -1 2192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5642_6
timestamp 1731220558
transform 1 0 2288 0 -1 2192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5641_6
timestamp 1731220558
transform 1 0 2192 0 -1 2192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5640_6
timestamp 1731220558
transform 1 0 2512 0 -1 2192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5639_6
timestamp 1731220558
transform 1 0 2632 0 -1 2192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5638_6
timestamp 1731220558
transform 1 0 2752 0 -1 2192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5637_6
timestamp 1731220558
transform 1 0 2712 0 1 2028
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5636_6
timestamp 1731220558
transform 1 0 2592 0 1 2028
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5635_6
timestamp 1731220558
transform 1 0 2472 0 1 2028
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5634_6
timestamp 1731220558
transform 1 0 2360 0 1 2028
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5633_6
timestamp 1731220558
transform 1 0 2256 0 1 2028
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5632_6
timestamp 1731220558
transform 1 0 2160 0 1 2028
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5631_6
timestamp 1731220558
transform 1 0 2512 0 -1 2024
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5630_6
timestamp 1731220558
transform 1 0 2352 0 -1 2024
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5629_6
timestamp 1731220558
transform 1 0 2200 0 -1 2024
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5628_6
timestamp 1731220558
transform 1 0 2064 0 -1 2024
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5627_6
timestamp 1731220558
transform 1 0 1992 0 1 1872
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5626_6
timestamp 1731220558
transform 1 0 2120 0 1 1872
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5625_6
timestamp 1731220558
transform 1 0 2240 0 1 1872
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5624_6
timestamp 1731220558
transform 1 0 2376 0 -1 1872
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5623_6
timestamp 1731220558
transform 1 0 2240 0 -1 1872
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5622_6
timestamp 1731220558
transform 1 0 2112 0 -1 1872
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5621_6
timestamp 1731220558
transform 1 0 1736 0 1 1788
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5620_6
timestamp 1731220558
transform 1 0 1616 0 1 1788
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5619_6
timestamp 1731220558
transform 1 0 1472 0 1 1788
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5618_6
timestamp 1731220558
transform 1 0 1336 0 1 1788
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5617_6
timestamp 1731220558
transform 1 0 1616 0 -1 1940
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5616_6
timestamp 1731220558
transform 1 0 1480 0 -1 1940
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5615_6
timestamp 1731220558
transform 1 0 1344 0 -1 1940
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5614_6
timestamp 1731220558
transform 1 0 1208 0 -1 1940
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5613_6
timestamp 1731220558
transform 1 0 1472 0 1 1948
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5612_6
timestamp 1731220558
transform 1 0 1376 0 1 1948
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5611_6
timestamp 1731220558
transform 1 0 1280 0 1 1948
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5610_6
timestamp 1731220558
transform 1 0 1192 0 1 1948
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5609_6
timestamp 1731220558
transform 1 0 1096 0 1 1948
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5608_6
timestamp 1731220558
transform 1 0 1304 0 -1 2100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5607_6
timestamp 1731220558
transform 1 0 1096 0 -1 2100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5606_6
timestamp 1731220558
transform 1 0 1008 0 1 1948
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5605_6
timestamp 1731220558
transform 1 0 912 0 1 1948
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5604_6
timestamp 1731220558
transform 1 0 808 0 1 1948
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5603_6
timestamp 1731220558
transform 1 0 936 0 -1 1940
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5602_6
timestamp 1731220558
transform 1 0 1072 0 -1 1940
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5601_6
timestamp 1731220558
transform 1 0 1040 0 1 1788
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5600_6
timestamp 1731220558
transform 1 0 1192 0 1 1788
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5599_6
timestamp 1731220558
transform 1 0 1136 0 -1 1784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5598_6
timestamp 1731220558
transform 1 0 1016 0 -1 1784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5597_6
timestamp 1731220558
transform 1 0 888 0 -1 1784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5596_6
timestamp 1731220558
transform 1 0 1384 0 -1 1784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5595_6
timestamp 1731220558
transform 1 0 1256 0 -1 1784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5594_6
timestamp 1731220558
transform 1 0 1168 0 1 1628
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5593_6
timestamp 1731220558
transform 1 0 1304 0 1 1628
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5592_6
timestamp 1731220558
transform 1 0 1432 0 1 1628
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5591_6
timestamp 1731220558
transform 1 0 1560 0 1 1628
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5590_6
timestamp 1731220558
transform 1 0 1696 0 1 1628
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5589_6
timestamp 1731220558
transform 1 0 1736 0 -1 1620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5588_6
timestamp 1731220558
transform 1 0 1616 0 -1 1620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5587_6
timestamp 1731220558
transform 1 0 1488 0 -1 1620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5586_6
timestamp 1731220558
transform 1 0 1352 0 -1 1620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5585_6
timestamp 1731220558
transform 1 0 1216 0 -1 1620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5584_6
timestamp 1731220558
transform 1 0 1064 0 -1 1620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5583_6
timestamp 1731220558
transform 1 0 1456 0 1 1464
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5582_6
timestamp 1731220558
transform 1 0 1320 0 1 1464
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5581_6
timestamp 1731220558
transform 1 0 1192 0 1 1464
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5580_6
timestamp 1731220558
transform 1 0 1064 0 1 1464
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5579_6
timestamp 1731220558
transform 1 0 936 0 1 1464
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5578_6
timestamp 1731220558
transform 1 0 1248 0 -1 1460
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5577_6
timestamp 1731220558
transform 1 0 1136 0 -1 1460
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5576_6
timestamp 1731220558
transform 1 0 1032 0 -1 1460
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5575_6
timestamp 1731220558
transform 1 0 928 0 -1 1460
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5574_6
timestamp 1731220558
transform 1 0 824 0 -1 1460
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5573_6
timestamp 1731220558
transform 1 0 712 0 -1 1460
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5572_6
timestamp 1731220558
transform 1 0 1152 0 1 1292
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5571_6
timestamp 1731220558
transform 1 0 1008 0 1 1292
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5570_6
timestamp 1731220558
transform 1 0 864 0 1 1292
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5569_6
timestamp 1731220558
transform 1 0 720 0 1 1292
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5568_6
timestamp 1731220558
transform 1 0 568 0 1 1292
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5567_6
timestamp 1731220558
transform 1 0 752 0 -1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5566_6
timestamp 1731220558
transform 1 0 920 0 -1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5565_6
timestamp 1731220558
transform 1 0 832 0 1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5564_6
timestamp 1731220558
transform 1 0 768 0 -1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5563_6
timestamp 1731220558
transform 1 0 640 0 -1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5562_6
timestamp 1731220558
transform 1 0 560 0 1 964
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5561_6
timestamp 1731220558
transform 1 0 456 0 1 964
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5560_6
timestamp 1731220558
transform 1 0 656 0 1 964
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5559_6
timestamp 1731220558
transform 1 0 696 0 -1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5558_6
timestamp 1731220558
transform 1 0 832 0 -1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5557_6
timestamp 1731220558
transform 1 0 800 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5556_6
timestamp 1731220558
transform 1 0 648 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5555_6
timestamp 1731220558
transform 1 0 552 0 -1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5554_6
timestamp 1731220558
transform 1 0 408 0 -1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5553_6
timestamp 1731220558
transform 1 0 256 0 -1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5552_6
timestamp 1731220558
transform 1 0 224 0 1 964
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5551_6
timestamp 1731220558
transform 1 0 344 0 1 964
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5550_6
timestamp 1731220558
transform 1 0 512 0 -1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5549_6
timestamp 1731220558
transform 1 0 376 0 -1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5548_6
timestamp 1731220558
transform 1 0 240 0 -1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5547_6
timestamp 1731220558
transform 1 0 296 0 1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5546_6
timestamp 1731220558
transform 1 0 656 0 1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5545_6
timestamp 1731220558
transform 1 0 472 0 1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5544_6
timestamp 1731220558
transform 1 0 584 0 -1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5543_6
timestamp 1731220558
transform 1 0 416 0 -1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5542_6
timestamp 1731220558
transform 1 0 416 0 1 1292
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5541_6
timestamp 1731220558
transform 1 0 272 0 1 1292
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5540_6
timestamp 1731220558
transform 1 0 352 0 -1 1460
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5539_6
timestamp 1731220558
transform 1 0 472 0 -1 1460
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5538_6
timestamp 1731220558
transform 1 0 592 0 -1 1460
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5537_6
timestamp 1731220558
transform 1 0 800 0 1 1464
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5536_6
timestamp 1731220558
transform 1 0 656 0 1 1464
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5535_6
timestamp 1731220558
transform 1 0 512 0 1 1464
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5534_6
timestamp 1731220558
transform 1 0 368 0 1 1464
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5533_6
timestamp 1731220558
transform 1 0 536 0 -1 1620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5532_6
timestamp 1731220558
transform 1 0 720 0 -1 1620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5531_6
timestamp 1731220558
transform 1 0 896 0 -1 1620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5530_6
timestamp 1731220558
transform 1 0 1024 0 1 1628
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5529_6
timestamp 1731220558
transform 1 0 880 0 1 1628
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5528_6
timestamp 1731220558
transform 1 0 728 0 1 1628
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5527_6
timestamp 1731220558
transform 1 0 576 0 1 1628
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5526_6
timestamp 1731220558
transform 1 0 584 0 -1 1784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5525_6
timestamp 1731220558
transform 1 0 744 0 -1 1784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5524_6
timestamp 1731220558
transform 1 0 888 0 1 1788
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5523_6
timestamp 1731220558
transform 1 0 736 0 1 1788
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5522_6
timestamp 1731220558
transform 1 0 584 0 1 1788
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5521_6
timestamp 1731220558
transform 1 0 480 0 -1 1940
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5520_6
timestamp 1731220558
transform 1 0 640 0 -1 1940
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5519_6
timestamp 1731220558
transform 1 0 792 0 -1 1940
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5518_6
timestamp 1731220558
transform 1 0 704 0 1 1948
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5517_6
timestamp 1731220558
transform 1 0 592 0 1 1948
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5516_6
timestamp 1731220558
transform 1 0 480 0 1 1948
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5515_6
timestamp 1731220558
transform 1 0 512 0 -1 2100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5514_6
timestamp 1731220558
transform 1 0 696 0 -1 2100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5513_6
timestamp 1731220558
transform 1 0 888 0 -1 2100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5512_6
timestamp 1731220558
transform 1 0 808 0 1 2104
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5511_6
timestamp 1731220558
transform 1 0 624 0 1 2104
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5510_6
timestamp 1731220558
transform 1 0 1000 0 1 2104
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5509_6
timestamp 1731220558
transform 1 0 992 0 -1 2260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5508_6
timestamp 1731220558
transform 1 0 824 0 -1 2260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5507_6
timestamp 1731220558
transform 1 0 664 0 -1 2260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5506_6
timestamp 1731220558
transform 1 0 512 0 -1 2260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5505_6
timestamp 1731220558
transform 1 0 376 0 -1 2260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5504_6
timestamp 1731220558
transform 1 0 288 0 -1 2260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5503_6
timestamp 1731220558
transform 1 0 208 0 -1 2260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5502_6
timestamp 1731220558
transform 1 0 128 0 -1 2260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5501_6
timestamp 1731220558
transform 1 0 176 0 1 2104
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5500_6
timestamp 1731220558
transform 1 0 448 0 1 2104
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5499_6
timestamp 1731220558
transform 1 0 296 0 1 2104
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5498_6
timestamp 1731220558
transform 1 0 208 0 -1 2100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5497_6
timestamp 1731220558
transform 1 0 352 0 -1 2100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5496_6
timestamp 1731220558
transform 1 0 368 0 1 1948
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5495_6
timestamp 1731220558
transform 1 0 248 0 1 1948
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5494_6
timestamp 1731220558
transform 1 0 128 0 1 1948
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5493_6
timestamp 1731220558
transform 1 0 160 0 -1 1940
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5492_6
timestamp 1731220558
transform 1 0 320 0 -1 1940
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5491_6
timestamp 1731220558
transform 1 0 288 0 1 1788
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5490_6
timestamp 1731220558
transform 1 0 144 0 1 1788
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5489_6
timestamp 1731220558
transform 1 0 432 0 1 1788
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5488_6
timestamp 1731220558
transform 1 0 416 0 -1 1784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5487_6
timestamp 1731220558
transform 1 0 240 0 -1 1784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5486_6
timestamp 1731220558
transform 1 0 432 0 1 1628
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5485_6
timestamp 1731220558
transform 1 0 296 0 1 1628
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5484_6
timestamp 1731220558
transform 1 0 176 0 1 1628
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5483_6
timestamp 1731220558
transform 1 0 160 0 -1 1620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5482_6
timestamp 1731220558
transform 1 0 344 0 -1 1620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5481_6
timestamp 1731220558
transform 1 0 232 0 1 1464
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5480_6
timestamp 1731220558
transform 1 0 128 0 1 1464
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5479_6
timestamp 1731220558
transform 1 0 128 0 -1 1460
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5478_6
timestamp 1731220558
transform 1 0 224 0 -1 1460
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5477_6
timestamp 1731220558
transform 1 0 128 0 1 1292
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5476_6
timestamp 1731220558
transform 1 0 128 0 -1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5475_6
timestamp 1731220558
transform 1 0 256 0 -1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5474_6
timestamp 1731220558
transform 1 0 128 0 1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5473_6
timestamp 1731220558
transform 1 0 128 0 -1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5472_6
timestamp 1731220558
transform 1 0 128 0 1 964
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5471_6
timestamp 1731220558
transform 1 0 128 0 -1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5470_6
timestamp 1731220558
transform 1 0 128 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5469_6
timestamp 1731220558
transform 1 0 232 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5468_6
timestamp 1731220558
transform 1 0 504 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5467_6
timestamp 1731220558
transform 1 0 368 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5466_6
timestamp 1731220558
transform 1 0 296 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5465_6
timestamp 1731220558
transform 1 0 208 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5464_6
timestamp 1731220558
transform 1 0 128 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5463_6
timestamp 1731220558
transform 1 0 680 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5462_6
timestamp 1731220558
transform 1 0 536 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5461_6
timestamp 1731220558
transform 1 0 408 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5460_6
timestamp 1731220558
transform 1 0 408 0 1 624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5459_6
timestamp 1731220558
transform 1 0 304 0 1 624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5458_6
timestamp 1731220558
transform 1 0 216 0 1 624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5457_6
timestamp 1731220558
transform 1 0 528 0 1 624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5456_6
timestamp 1731220558
transform 1 0 664 0 1 624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5455_6
timestamp 1731220558
transform 1 0 800 0 1 624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5454_6
timestamp 1731220558
transform 1 0 768 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5453_6
timestamp 1731220558
transform 1 0 680 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5452_6
timestamp 1731220558
transform 1 0 600 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5451_6
timestamp 1731220558
transform 1 0 520 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5450_6
timestamp 1731220558
transform 1 0 440 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5449_6
timestamp 1731220558
transform 1 0 576 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5448_6
timestamp 1731220558
transform 1 0 496 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5447_6
timestamp 1731220558
transform 1 0 408 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5446_6
timestamp 1731220558
transform 1 0 320 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5445_6
timestamp 1731220558
transform 1 0 216 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5444_6
timestamp 1731220558
transform 1 0 328 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5443_6
timestamp 1731220558
transform 1 0 440 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5442_6
timestamp 1731220558
transform 1 0 384 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5441_6
timestamp 1731220558
transform 1 0 248 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5440_6
timestamp 1731220558
transform 1 0 128 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5439_6
timestamp 1731220558
transform 1 0 128 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5438_6
timestamp 1731220558
transform 1 0 240 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5437_6
timestamp 1731220558
transform 1 0 384 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5436_6
timestamp 1731220558
transform 1 0 288 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5435_6
timestamp 1731220558
transform 1 0 208 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5434_6
timestamp 1731220558
transform 1 0 128 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5433_6
timestamp 1731220558
transform 1 0 368 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5432_6
timestamp 1731220558
transform 1 0 448 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5431_6
timestamp 1731220558
transform 1 0 528 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5430_6
timestamp 1731220558
transform 1 0 768 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5429_6
timestamp 1731220558
transform 1 0 688 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5428_6
timestamp 1731220558
transform 1 0 608 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5427_6
timestamp 1731220558
transform 1 0 536 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5426_6
timestamp 1731220558
transform 1 0 688 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5425_6
timestamp 1731220558
transform 1 0 840 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5424_6
timestamp 1731220558
transform 1 0 776 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5423_6
timestamp 1731220558
transform 1 0 656 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5422_6
timestamp 1731220558
transform 1 0 520 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5421_6
timestamp 1731220558
transform 1 0 552 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5420_6
timestamp 1731220558
transform 1 0 656 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5419_6
timestamp 1731220558
transform 1 0 752 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5418_6
timestamp 1731220558
transform 1 0 736 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5417_6
timestamp 1731220558
transform 1 0 656 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5416_6
timestamp 1731220558
transform 1 0 864 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5415_6
timestamp 1731220558
transform 1 0 952 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5414_6
timestamp 1731220558
transform 1 0 936 0 1 624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5413_6
timestamp 1731220558
transform 1 0 832 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5412_6
timestamp 1731220558
transform 1 0 984 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5411_6
timestamp 1731220558
transform 1 0 1136 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5410_6
timestamp 1731220558
transform 1 0 1232 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5409_6
timestamp 1731220558
transform 1 0 1088 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5408_6
timestamp 1731220558
transform 1 0 944 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5407_6
timestamp 1731220558
transform 1 0 968 0 -1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5406_6
timestamp 1731220558
transform 1 0 1096 0 -1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5405_6
timestamp 1731220558
transform 1 0 1216 0 -1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5404_6
timestamp 1731220558
transform 1 0 1208 0 1 964
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5403_6
timestamp 1731220558
transform 1 0 1112 0 1 964
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5402_6
timestamp 1731220558
transform 1 0 1016 0 1 964
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5401_6
timestamp 1731220558
transform 1 0 928 0 1 964
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5400_6
timestamp 1731220558
transform 1 0 840 0 1 964
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5399_6
timestamp 1731220558
transform 1 0 752 0 1 964
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5398_6
timestamp 1731220558
transform 1 0 888 0 -1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5397_6
timestamp 1731220558
transform 1 0 1008 0 -1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5396_6
timestamp 1731220558
transform 1 0 1128 0 -1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5395_6
timestamp 1731220558
transform 1 0 1496 0 -1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5394_6
timestamp 1731220558
transform 1 0 1368 0 -1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5393_6
timestamp 1731220558
transform 1 0 1248 0 -1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5392_6
timestamp 1731220558
transform 1 0 1144 0 1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5391_6
timestamp 1731220558
transform 1 0 992 0 1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5390_6
timestamp 1731220558
transform 1 0 1280 0 1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5389_6
timestamp 1731220558
transform 1 0 1216 0 -1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5388_6
timestamp 1731220558
transform 1 0 1072 0 -1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5387_6
timestamp 1731220558
transform 1 0 1344 0 -1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5386_6
timestamp 1731220558
transform 1 0 1304 0 1 1292
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5385_6
timestamp 1731220558
transform 1 0 1456 0 1 1292
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5384_6
timestamp 1731220558
transform 1 0 1608 0 1 1292
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5383_6
timestamp 1731220558
transform 1 0 1600 0 -1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5382_6
timestamp 1731220558
transform 1 0 1472 0 -1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5381_6
timestamp 1731220558
transform 1 0 1728 0 -1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5380_6
timestamp 1731220558
transform 1 0 1736 0 1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5379_6
timestamp 1731220558
transform 1 0 1640 0 1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5378_6
timestamp 1731220558
transform 1 0 1520 0 1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5377_6
timestamp 1731220558
transform 1 0 1400 0 1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5376_6
timestamp 1731220558
transform 1 0 1624 0 -1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5375_6
timestamp 1731220558
transform 1 0 1736 0 -1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5374_6
timestamp 1731220558
transform 1 0 1888 0 1 1060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5373_6
timestamp 1731220558
transform 1 0 1888 0 -1 1060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5372_6
timestamp 1731220558
transform 1 0 2008 0 -1 1060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5371_6
timestamp 1731220558
transform 1 0 2160 0 -1 1060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5370_6
timestamp 1731220558
transform 1 0 2184 0 1 904
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5369_6
timestamp 1731220558
transform 1 0 2064 0 1 904
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5368_6
timestamp 1731220558
transform 1 0 1968 0 1 904
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5367_6
timestamp 1731220558
transform 1 0 1888 0 1 904
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5366_6
timestamp 1731220558
transform 1 0 1736 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5365_6
timestamp 1731220558
transform 1 0 1736 0 -1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5364_6
timestamp 1731220558
transform 1 0 1648 0 -1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5363_6
timestamp 1731220558
transform 1 0 1536 0 -1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5362_6
timestamp 1731220558
transform 1 0 1432 0 -1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5361_6
timestamp 1731220558
transform 1 0 1328 0 -1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5360_6
timestamp 1731220558
transform 1 0 1368 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5359_6
timestamp 1731220558
transform 1 0 1624 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5358_6
timestamp 1731220558
transform 1 0 1496 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5357_6
timestamp 1731220558
transform 1 0 1440 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5356_6
timestamp 1731220558
transform 1 0 1288 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5355_6
timestamp 1731220558
transform 1 0 1600 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5354_6
timestamp 1731220558
transform 1 0 1568 0 1 624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5353_6
timestamp 1731220558
transform 1 0 1440 0 1 624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5352_6
timestamp 1731220558
transform 1 0 1320 0 1 624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5351_6
timestamp 1731220558
transform 1 0 1200 0 1 624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5350_6
timestamp 1731220558
transform 1 0 1072 0 1 624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5349_6
timestamp 1731220558
transform 1 0 1424 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5348_6
timestamp 1731220558
transform 1 0 1328 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5347_6
timestamp 1731220558
transform 1 0 1232 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5346_6
timestamp 1731220558
transform 1 0 1136 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5345_6
timestamp 1731220558
transform 1 0 1040 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5344_6
timestamp 1731220558
transform 1 0 1264 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5343_6
timestamp 1731220558
transform 1 0 1176 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5342_6
timestamp 1731220558
transform 1 0 1088 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5341_6
timestamp 1731220558
transform 1 0 1000 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5340_6
timestamp 1731220558
transform 1 0 912 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5339_6
timestamp 1731220558
transform 1 0 824 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5338_6
timestamp 1731220558
transform 1 0 840 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5337_6
timestamp 1731220558
transform 1 0 928 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5336_6
timestamp 1731220558
transform 1 0 1016 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5335_6
timestamp 1731220558
transform 1 0 1104 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5334_6
timestamp 1731220558
transform 1 0 1288 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5333_6
timestamp 1731220558
transform 1 0 1192 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5332_6
timestamp 1731220558
transform 1 0 1112 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5331_6
timestamp 1731220558
transform 1 0 1008 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5330_6
timestamp 1731220558
transform 1 0 896 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5329_6
timestamp 1731220558
transform 1 0 1216 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5328_6
timestamp 1731220558
transform 1 0 1424 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5327_6
timestamp 1731220558
transform 1 0 1320 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5326_6
timestamp 1731220558
transform 1 0 1232 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5325_6
timestamp 1731220558
transform 1 0 1112 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5324_6
timestamp 1731220558
transform 1 0 984 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5323_6
timestamp 1731220558
transform 1 0 1592 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5322_6
timestamp 1731220558
transform 1 0 1472 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5321_6
timestamp 1731220558
transform 1 0 1352 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5320_6
timestamp 1731220558
transform 1 0 1008 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5319_6
timestamp 1731220558
transform 1 0 928 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5318_6
timestamp 1731220558
transform 1 0 848 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5317_6
timestamp 1731220558
transform 1 0 1088 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5316_6
timestamp 1731220558
transform 1 0 1168 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5315_6
timestamp 1731220558
transform 1 0 1248 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5314_6
timestamp 1731220558
transform 1 0 1328 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5313_6
timestamp 1731220558
transform 1 0 1408 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5312_6
timestamp 1731220558
transform 1 0 1496 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5311_6
timestamp 1731220558
transform 1 0 1576 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5310_6
timestamp 1731220558
transform 1 0 1656 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5309_6
timestamp 1731220558
transform 1 0 1736 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5308_6
timestamp 1731220558
transform 1 0 1888 0 1 100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5307_6
timestamp 1731220558
transform 1 0 1968 0 1 100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5306_6
timestamp 1731220558
transform 1 0 2072 0 1 100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5305_6
timestamp 1731220558
transform 1 0 2472 0 1 100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5304_6
timestamp 1731220558
transform 1 0 2336 0 1 100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5303_6
timestamp 1731220558
transform 1 0 2200 0 1 100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5302_6
timestamp 1731220558
transform 1 0 2112 0 -1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5301_6
timestamp 1731220558
transform 1 0 1984 0 -1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5300_6
timestamp 1731220558
transform 1 0 2248 0 -1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5299_6
timestamp 1731220558
transform 1 0 2384 0 -1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5298_6
timestamp 1731220558
transform 1 0 2528 0 -1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5297_6
timestamp 1731220558
transform 1 0 2704 0 1 268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5296_6
timestamp 1731220558
transform 1 0 2576 0 1 268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5295_6
timestamp 1731220558
transform 1 0 2464 0 1 268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5294_6
timestamp 1731220558
transform 1 0 2368 0 1 268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5293_6
timestamp 1731220558
transform 1 0 2280 0 1 268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5292_6
timestamp 1731220558
transform 1 0 2200 0 1 268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5291_6
timestamp 1731220558
transform 1 0 2352 0 -1 424
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5290_6
timestamp 1731220558
transform 1 0 2248 0 -1 424
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5289_6
timestamp 1731220558
transform 1 0 2152 0 -1 424
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5288_6
timestamp 1731220558
transform 1 0 2056 0 -1 424
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5287_6
timestamp 1731220558
transform 1 0 1968 0 -1 424
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5286_6
timestamp 1731220558
transform 1 0 2176 0 1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5285_6
timestamp 1731220558
transform 1 0 2272 0 1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5284_6
timestamp 1731220558
transform 1 0 2368 0 1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5283_6
timestamp 1731220558
transform 1 0 2472 0 1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5282_6
timestamp 1731220558
transform 1 0 2688 0 -1 588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5281_6
timestamp 1731220558
transform 1 0 2584 0 -1 588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5280_6
timestamp 1731220558
transform 1 0 2496 0 -1 588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5279_6
timestamp 1731220558
transform 1 0 2416 0 -1 588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5278_6
timestamp 1731220558
transform 1 0 2336 0 -1 588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5277_6
timestamp 1731220558
transform 1 0 2256 0 -1 588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5276_6
timestamp 1731220558
transform 1 0 2592 0 1 588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5275_6
timestamp 1731220558
transform 1 0 2472 0 1 588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5274_6
timestamp 1731220558
transform 1 0 2360 0 1 588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5273_6
timestamp 1731220558
transform 1 0 2256 0 1 588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5272_6
timestamp 1731220558
transform 1 0 2160 0 1 588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5271_6
timestamp 1731220558
transform 1 0 2592 0 -1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5270_6
timestamp 1731220558
transform 1 0 2440 0 -1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5269_6
timestamp 1731220558
transform 1 0 2296 0 -1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5268_6
timestamp 1731220558
transform 1 0 2168 0 -1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5267_6
timestamp 1731220558
transform 1 0 2056 0 -1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5266_6
timestamp 1731220558
transform 1 0 1960 0 -1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5265_6
timestamp 1731220558
transform 1 0 2472 0 1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5264_6
timestamp 1731220558
transform 1 0 2312 0 1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5263_6
timestamp 1731220558
transform 1 0 2152 0 1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5262_6
timestamp 1731220558
transform 1 0 2000 0 1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5261_6
timestamp 1731220558
transform 1 0 1888 0 1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5260_6
timestamp 1731220558
transform 1 0 1912 0 -1 892
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5259_6
timestamp 1731220558
transform 1 0 2088 0 -1 892
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5258_6
timestamp 1731220558
transform 1 0 2264 0 -1 892
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5257_6
timestamp 1731220558
transform 1 0 2320 0 1 904
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5256_6
timestamp 1731220558
transform 1 0 2464 0 1 904
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5255_6
timestamp 1731220558
transform 1 0 2480 0 -1 1060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5254_6
timestamp 1731220558
transform 1 0 2320 0 -1 1060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5253_6
timestamp 1731220558
transform 1 0 2112 0 1 1060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5252_6
timestamp 1731220558
transform 1 0 2344 0 1 1060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5251_6
timestamp 1731220558
transform 1 0 2520 0 -1 1220
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5250_6
timestamp 1731220558
transform 1 0 2400 0 -1 1220
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5249_6
timestamp 1731220558
transform 1 0 2296 0 -1 1220
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5248_6
timestamp 1731220558
transform 1 0 2200 0 -1 1220
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5247_6
timestamp 1731220558
transform 1 0 2104 0 -1 1220
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5246_6
timestamp 1731220558
transform 1 0 2200 0 1 1224
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5245_6
timestamp 1731220558
transform 1 0 2280 0 1 1224
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5244_6
timestamp 1731220558
transform 1 0 2360 0 1 1224
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5243_6
timestamp 1731220558
transform 1 0 2648 0 1 1224
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5242_6
timestamp 1731220558
transform 1 0 2536 0 1 1224
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5241_6
timestamp 1731220558
transform 1 0 2440 0 1 1224
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5240_6
timestamp 1731220558
transform 1 0 2416 0 -1 1388
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5239_6
timestamp 1731220558
transform 1 0 2488 0 1 1388
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5238_6
timestamp 1731220558
transform 1 0 2408 0 1 1388
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5237_6
timestamp 1731220558
transform 1 0 2328 0 1 1388
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5236_6
timestamp 1731220558
transform 1 0 2248 0 1 1388
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5235_6
timestamp 1731220558
transform 1 0 2528 0 -1 1544
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5234_6
timestamp 1731220558
transform 1 0 2432 0 -1 1544
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5233_6
timestamp 1731220558
transform 1 0 2336 0 -1 1544
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5232_6
timestamp 1731220558
transform 1 0 2248 0 -1 1544
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5231_6
timestamp 1731220558
transform 1 0 2160 0 -1 1544
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5230_6
timestamp 1731220558
transform 1 0 2080 0 -1 1544
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5229_6
timestamp 1731220558
transform 1 0 2488 0 1 1548
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5228_6
timestamp 1731220558
transform 1 0 2352 0 1 1548
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5227_6
timestamp 1731220558
transform 1 0 2216 0 1 1548
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5226_6
timestamp 1731220558
transform 1 0 2080 0 1 1548
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5225_6
timestamp 1731220558
transform 1 0 1960 0 1 1548
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5224_6
timestamp 1731220558
transform 1 0 2640 0 -1 1704
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5223_6
timestamp 1731220558
transform 1 0 2464 0 -1 1704
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5222_6
timestamp 1731220558
transform 1 0 2288 0 -1 1704
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5221_6
timestamp 1731220558
transform 1 0 2128 0 -1 1704
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5220_6
timestamp 1731220558
transform 1 0 1984 0 -1 1704
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5219_6
timestamp 1731220558
transform 1 0 1888 0 -1 1704
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5218_6
timestamp 1731220558
transform 1 0 2512 0 1 1708
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5217_6
timestamp 1731220558
transform 1 0 2344 0 1 1708
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5216_6
timestamp 1731220558
transform 1 0 2176 0 1 1708
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5215_6
timestamp 1731220558
transform 1 0 2016 0 1 1708
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5214_6
timestamp 1731220558
transform 1 0 1888 0 1 1708
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5213_6
timestamp 1731220558
transform 1 0 1984 0 -1 1872
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5212_6
timestamp 1731220558
transform 1 0 1888 0 -1 1872
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5211_6
timestamp 1731220558
transform 1 0 1888 0 1 1872
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5210_6
timestamp 1731220558
transform 1 0 1736 0 -1 1940
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5209_6
timestamp 1731220558
transform 1 0 1736 0 1 1948
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5208_6
timestamp 1731220558
transform 1 0 1656 0 1 1948
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5207_6
timestamp 1731220558
transform 1 0 1568 0 1 1948
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5206_6
timestamp 1731220558
transform 1 0 1520 0 -1 2100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5205_6
timestamp 1731220558
transform 1 0 1736 0 -1 2100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5204_6
timestamp 1731220558
transform 1 0 1736 0 1 2104
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5203_6
timestamp 1731220558
transform 1 0 1568 0 1 2104
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5202_6
timestamp 1731220558
transform 1 0 1376 0 1 2104
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5201_6
timestamp 1731220558
transform 1 0 1184 0 1 2104
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5200_6
timestamp 1731220558
transform 1 0 1736 0 -1 2260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5199_6
timestamp 1731220558
transform 1 0 1600 0 -1 2260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5198_6
timestamp 1731220558
transform 1 0 1448 0 -1 2260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5197_6
timestamp 1731220558
transform 1 0 1304 0 -1 2260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5196_6
timestamp 1731220558
transform 1 0 1152 0 -1 2260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5195_6
timestamp 1731220558
transform 1 0 1632 0 1 2268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5194_6
timestamp 1731220558
transform 1 0 1552 0 1 2268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5193_6
timestamp 1731220558
transform 1 0 1472 0 1 2268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5192_6
timestamp 1731220558
transform 1 0 1392 0 1 2268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5191_6
timestamp 1731220558
transform 1 0 1344 0 -1 2420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5190_6
timestamp 1731220558
transform 1 0 1432 0 -1 2420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5189_6
timestamp 1731220558
transform 1 0 1520 0 -1 2420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5188_6
timestamp 1731220558
transform 1 0 1456 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5187_6
timestamp 1731220558
transform 1 0 1312 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5186_6
timestamp 1731220558
transform 1 0 1248 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5185_6
timestamp 1731220558
transform 1 0 1384 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5184_6
timestamp 1731220558
transform 1 0 1520 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5183_6
timestamp 1731220558
transform 1 0 1552 0 1 2588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5182_6
timestamp 1731220558
transform 1 0 1376 0 1 2588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5181_6
timestamp 1731220558
transform 1 0 1352 0 -1 2740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5180_6
timestamp 1731220558
transform 1 0 1512 0 -1 2740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5179_6
timestamp 1731220558
transform 1 0 1680 0 -1 2740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5178_6
timestamp 1731220558
transform 1 0 1720 0 1 2744
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5177_6
timestamp 1731220558
transform 1 0 1520 0 1 2744
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5176_6
timestamp 1731220558
transform 1 0 1488 0 -1 2896
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5175_6
timestamp 1731220558
transform 1 0 1624 0 -1 2896
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5174_6
timestamp 1731220558
transform 1 0 1736 0 -1 2896
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5173_6
timestamp 1731220558
transform 1 0 1736 0 1 2896
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5172_6
timestamp 1731220558
transform 1 0 1888 0 1 2864
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5171_6
timestamp 1731220558
transform 1 0 1888 0 -1 3016
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5170_6
timestamp 1731220558
transform 1 0 2040 0 -1 3016
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5169_6
timestamp 1731220558
transform 1 0 2000 0 1 3024
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5168_6
timestamp 1731220558
transform 1 0 1888 0 1 3024
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5167_6
timestamp 1731220558
transform 1 0 2176 0 1 3024
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5166_6
timestamp 1731220558
transform 1 0 2112 0 -1 3192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5165_6
timestamp 1731220558
transform 1 0 1984 0 -1 3192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5164_6
timestamp 1731220558
transform 1 0 1888 0 -1 3192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5163_6
timestamp 1731220558
transform 1 0 1736 0 -1 3208
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5162_6
timestamp 1731220558
transform 1 0 1736 0 1 3208
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5161_6
timestamp 1731220558
transform 1 0 1624 0 1 3208
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5160_6
timestamp 1731220558
transform 1 0 1496 0 1 3208
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5159_6
timestamp 1731220558
transform 1 0 1368 0 1 3208
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5158_6
timestamp 1731220558
transform 1 0 1416 0 -1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5157_6
timestamp 1731220558
transform 1 0 1576 0 -1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5156_6
timestamp 1731220558
transform 1 0 1736 0 -1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5155_6
timestamp 1731220558
transform 1 0 1696 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5154_6
timestamp 1731220558
transform 1 0 1544 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5153_6
timestamp 1731220558
transform 1 0 1400 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5152_6
timestamp 1731220558
transform 1 0 1256 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5151_6
timestamp 1731220558
transform 1 0 1304 0 -1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5150_6
timestamp 1731220558
transform 1 0 1432 0 -1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5149_6
timestamp 1731220558
transform 1 0 1560 0 -1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5148_6
timestamp 1731220558
transform 1 0 1616 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5147_6
timestamp 1731220558
transform 1 0 1512 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5146_6
timestamp 1731220558
transform 1 0 1408 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5145_6
timestamp 1731220558
transform 1 0 1312 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5144_6
timestamp 1731220558
transform 1 0 1208 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5143_6
timestamp 1731220558
transform 1 0 1096 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5142_6
timestamp 1731220558
transform 1 0 984 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5141_6
timestamp 1731220558
transform 1 0 864 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5140_6
timestamp 1731220558
transform 1 0 912 0 -1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5139_6
timestamp 1731220558
transform 1 0 1048 0 -1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5138_6
timestamp 1731220558
transform 1 0 1176 0 -1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5137_6
timestamp 1731220558
transform 1 0 1104 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5136_6
timestamp 1731220558
transform 1 0 944 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5135_6
timestamp 1731220558
transform 1 0 936 0 -1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5134_6
timestamp 1731220558
transform 1 0 1096 0 -1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5133_6
timestamp 1731220558
transform 1 0 1256 0 -1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5132_6
timestamp 1731220558
transform 1 0 1240 0 1 3208
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5131_6
timestamp 1731220558
transform 1 0 1104 0 1 3208
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5130_6
timestamp 1731220558
transform 1 0 968 0 1 3208
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5129_6
timestamp 1731220558
transform 1 0 1016 0 -1 3208
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5128_6
timestamp 1731220558
transform 1 0 1184 0 -1 3208
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5127_6
timestamp 1731220558
transform 1 0 1560 0 -1 3208
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5126_6
timestamp 1731220558
transform 1 0 1368 0 -1 3208
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5125_6
timestamp 1731220558
transform 1 0 1360 0 1 3052
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5124_6
timestamp 1731220558
transform 1 0 1272 0 1 3052
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5123_6
timestamp 1731220558
transform 1 0 1184 0 1 3052
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5122_6
timestamp 1731220558
transform 1 0 1096 0 1 3052
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5121_6
timestamp 1731220558
transform 1 0 1008 0 1 3052
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5120_6
timestamp 1731220558
transform 1 0 1080 0 -1 3048
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5119_6
timestamp 1731220558
transform 1 0 1176 0 -1 3048
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5118_6
timestamp 1731220558
transform 1 0 1272 0 -1 3048
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5117_6
timestamp 1731220558
transform 1 0 1368 0 -1 3048
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5116_6
timestamp 1731220558
transform 1 0 1464 0 -1 3048
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5115_6
timestamp 1731220558
transform 1 0 1576 0 1 2896
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5114_6
timestamp 1731220558
transform 1 0 1400 0 1 2896
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5113_6
timestamp 1731220558
transform 1 0 1232 0 1 2896
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5112_6
timestamp 1731220558
transform 1 0 1072 0 1 2896
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5111_6
timestamp 1731220558
transform 1 0 1352 0 -1 2896
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5110_6
timestamp 1731220558
transform 1 0 1216 0 -1 2896
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5109_6
timestamp 1731220558
transform 1 0 1080 0 -1 2896
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5108_6
timestamp 1731220558
transform 1 0 944 0 -1 2896
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5107_6
timestamp 1731220558
transform 1 0 944 0 1 2744
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5106_6
timestamp 1731220558
transform 1 0 1128 0 1 2744
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5105_6
timestamp 1731220558
transform 1 0 1320 0 1 2744
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5104_6
timestamp 1731220558
transform 1 0 1192 0 -1 2740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5103_6
timestamp 1731220558
transform 1 0 1032 0 -1 2740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5102_6
timestamp 1731220558
transform 1 0 872 0 -1 2740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5101_6
timestamp 1731220558
transform 1 0 864 0 1 2588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5100_6
timestamp 1731220558
transform 1 0 1032 0 1 2588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_599_6
timestamp 1731220558
transform 1 0 1200 0 1 2588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_598_6
timestamp 1731220558
transform 1 0 1112 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_597_6
timestamp 1731220558
transform 1 0 976 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_596_6
timestamp 1731220558
transform 1 0 840 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_595_6
timestamp 1731220558
transform 1 0 920 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_594_6
timestamp 1731220558
transform 1 0 1048 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_593_6
timestamp 1731220558
transform 1 0 1176 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_592_6
timestamp 1731220558
transform 1 0 1256 0 -1 2420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_591_6
timestamp 1731220558
transform 1 0 1176 0 -1 2420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_590_6
timestamp 1731220558
transform 1 0 1096 0 -1 2420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_589_6
timestamp 1731220558
transform 1 0 1016 0 -1 2420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_588_6
timestamp 1731220558
transform 1 0 936 0 -1 2420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_587_6
timestamp 1731220558
transform 1 0 856 0 -1 2420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_586_6
timestamp 1731220558
transform 1 0 776 0 -1 2420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_585_6
timestamp 1731220558
transform 1 0 696 0 -1 2420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_584_6
timestamp 1731220558
transform 1 0 616 0 -1 2420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_583_6
timestamp 1731220558
transform 1 0 536 0 -1 2420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_582_6
timestamp 1731220558
transform 1 0 456 0 -1 2420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_581_6
timestamp 1731220558
transform 1 0 376 0 -1 2420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_580_6
timestamp 1731220558
transform 1 0 800 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_579_6
timestamp 1731220558
transform 1 0 688 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_578_6
timestamp 1731220558
transform 1 0 584 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_577_6
timestamp 1731220558
transform 1 0 488 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_576_6
timestamp 1731220558
transform 1 0 400 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_575_6
timestamp 1731220558
transform 1 0 320 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_574_6
timestamp 1731220558
transform 1 0 696 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_573_6
timestamp 1731220558
transform 1 0 552 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_572_6
timestamp 1731220558
transform 1 0 408 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_571_6
timestamp 1731220558
transform 1 0 272 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_570_6
timestamp 1731220558
transform 1 0 152 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_569_6
timestamp 1731220558
transform 1 0 696 0 1 2588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_568_6
timestamp 1731220558
transform 1 0 536 0 1 2588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_567_6
timestamp 1731220558
transform 1 0 384 0 1 2588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_566_6
timestamp 1731220558
transform 1 0 240 0 1 2588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_565_6
timestamp 1731220558
transform 1 0 128 0 1 2588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_564_6
timestamp 1731220558
transform 1 0 128 0 -1 2740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_563_6
timestamp 1731220558
transform 1 0 240 0 -1 2740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_562_6
timestamp 1731220558
transform 1 0 704 0 -1 2740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_561_6
timestamp 1731220558
transform 1 0 544 0 -1 2740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_560_6
timestamp 1731220558
transform 1 0 384 0 -1 2740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_559_6
timestamp 1731220558
transform 1 0 288 0 1 2744
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_558_6
timestamp 1731220558
transform 1 0 152 0 1 2744
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_557_6
timestamp 1731220558
transform 1 0 768 0 1 2744
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_556_6
timestamp 1731220558
transform 1 0 592 0 1 2744
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_555_6
timestamp 1731220558
transform 1 0 432 0 1 2744
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_554_6
timestamp 1731220558
transform 1 0 424 0 -1 2896
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_553_6
timestamp 1731220558
transform 1 0 304 0 -1 2896
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_552_6
timestamp 1731220558
transform 1 0 808 0 -1 2896
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_551_6
timestamp 1731220558
transform 1 0 672 0 -1 2896
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_550_6
timestamp 1731220558
transform 1 0 544 0 -1 2896
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_549_6
timestamp 1731220558
transform 1 0 456 0 1 2896
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_548_6
timestamp 1731220558
transform 1 0 560 0 1 2896
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_547_6
timestamp 1731220558
transform 1 0 928 0 1 2896
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_546_6
timestamp 1731220558
transform 1 0 792 0 1 2896
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_545_6
timestamp 1731220558
transform 1 0 672 0 1 2896
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_544_6
timestamp 1731220558
transform 1 0 616 0 -1 3048
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_543_6
timestamp 1731220558
transform 1 0 536 0 -1 3048
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_542_6
timestamp 1731220558
transform 1 0 704 0 -1 3048
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_541_6
timestamp 1731220558
transform 1 0 800 0 -1 3048
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_540_6
timestamp 1731220558
transform 1 0 896 0 -1 3048
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_539_6
timestamp 1731220558
transform 1 0 992 0 -1 3048
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_538_6
timestamp 1731220558
transform 1 0 920 0 1 3052
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_537_6
timestamp 1731220558
transform 1 0 832 0 1 3052
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_536_6
timestamp 1731220558
transform 1 0 744 0 1 3052
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_535_6
timestamp 1731220558
transform 1 0 656 0 1 3052
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_534_6
timestamp 1731220558
transform 1 0 576 0 1 3052
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_533_6
timestamp 1731220558
transform 1 0 880 0 -1 3208
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_532_6
timestamp 1731220558
transform 1 0 760 0 -1 3208
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_531_6
timestamp 1731220558
transform 1 0 656 0 -1 3208
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_530_6
timestamp 1731220558
transform 1 0 568 0 -1 3208
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_529_6
timestamp 1731220558
transform 1 0 480 0 -1 3208
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_528_6
timestamp 1731220558
transform 1 0 824 0 1 3208
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_527_6
timestamp 1731220558
transform 1 0 688 0 1 3208
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_526_6
timestamp 1731220558
transform 1 0 560 0 1 3208
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_525_6
timestamp 1731220558
transform 1 0 440 0 1 3208
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_524_6
timestamp 1731220558
transform 1 0 336 0 1 3208
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_523_6
timestamp 1731220558
transform 1 0 776 0 -1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_522_6
timestamp 1731220558
transform 1 0 616 0 -1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_521_6
timestamp 1731220558
transform 1 0 464 0 -1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_520_6
timestamp 1731220558
transform 1 0 328 0 -1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_519_6
timestamp 1731220558
transform 1 0 200 0 -1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_518_6
timestamp 1731220558
transform 1 0 776 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_517_6
timestamp 1731220558
transform 1 0 608 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_516_6
timestamp 1731220558
transform 1 0 440 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_515_6
timestamp 1731220558
transform 1 0 280 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_514_6
timestamp 1731220558
transform 1 0 136 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_513_6
timestamp 1731220558
transform 1 0 184 0 -1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_512_6
timestamp 1731220558
transform 1 0 320 0 -1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_511_6
timestamp 1731220558
transform 1 0 464 0 -1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_510_6
timestamp 1731220558
transform 1 0 616 0 -1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_59_6
timestamp 1731220558
transform 1 0 768 0 -1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_58_6
timestamp 1731220558
transform 1 0 728 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_57_6
timestamp 1731220558
transform 1 0 592 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_56_6
timestamp 1731220558
transform 1 0 456 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_55_6
timestamp 1731220558
transform 1 0 328 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_54_6
timestamp 1731220558
transform 1 0 208 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_53_6
timestamp 1731220558
transform 1 0 128 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_52_6
timestamp 1731220558
transform 1 0 128 0 -1 3668
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_51_6
timestamp 1731220558
transform 1 0 208 0 -1 3668
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_50_6
timestamp 1731220558
transform 1 0 288 0 -1 3668
box 8 4 70 72
<< end >>
