magic
tech sky130l
timestamp 1731220559
<< m2 >>
rect 2150 3648 2156 3649
rect 1870 3645 1876 3646
rect 1870 3641 1871 3645
rect 1875 3641 1876 3645
rect 2150 3644 2151 3648
rect 2155 3644 2156 3648
rect 2150 3643 2156 3644
rect 2438 3648 2444 3649
rect 2438 3644 2439 3648
rect 2443 3644 2444 3648
rect 2438 3643 2444 3644
rect 2726 3648 2732 3649
rect 2726 3644 2727 3648
rect 2731 3644 2732 3648
rect 2726 3643 2732 3644
rect 3014 3648 3020 3649
rect 3014 3644 3015 3648
rect 3019 3644 3020 3648
rect 3014 3643 3020 3644
rect 3590 3645 3596 3646
rect 1870 3640 1876 3641
rect 3590 3641 3591 3645
rect 3595 3641 3596 3645
rect 3590 3640 3596 3641
rect 1870 3628 1876 3629
rect 142 3626 148 3627
rect 142 3622 143 3626
rect 147 3622 148 3626
rect 142 3621 148 3622
rect 238 3626 244 3627
rect 238 3622 239 3626
rect 243 3622 244 3626
rect 238 3621 244 3622
rect 366 3626 372 3627
rect 366 3622 367 3626
rect 371 3622 372 3626
rect 366 3621 372 3622
rect 502 3626 508 3627
rect 502 3622 503 3626
rect 507 3622 508 3626
rect 502 3621 508 3622
rect 638 3626 644 3627
rect 638 3622 639 3626
rect 643 3622 644 3626
rect 638 3621 644 3622
rect 774 3626 780 3627
rect 774 3622 775 3626
rect 779 3622 780 3626
rect 774 3621 780 3622
rect 910 3626 916 3627
rect 910 3622 911 3626
rect 915 3622 916 3626
rect 910 3621 916 3622
rect 1054 3626 1060 3627
rect 1054 3622 1055 3626
rect 1059 3622 1060 3626
rect 1054 3621 1060 3622
rect 1198 3626 1204 3627
rect 1198 3622 1199 3626
rect 1203 3622 1204 3626
rect 1870 3624 1871 3628
rect 1875 3624 1876 3628
rect 1870 3623 1876 3624
rect 3590 3628 3596 3629
rect 3590 3624 3591 3628
rect 3595 3624 3596 3628
rect 3590 3623 3596 3624
rect 1198 3621 1204 3622
rect 2158 3610 2164 3611
rect 110 3608 116 3609
rect 110 3604 111 3608
rect 115 3604 116 3608
rect 110 3603 116 3604
rect 1830 3608 1836 3609
rect 1830 3604 1831 3608
rect 1835 3604 1836 3608
rect 2158 3606 2159 3610
rect 2163 3606 2164 3610
rect 2158 3605 2164 3606
rect 2446 3610 2452 3611
rect 2446 3606 2447 3610
rect 2451 3606 2452 3610
rect 2446 3605 2452 3606
rect 2734 3610 2740 3611
rect 2734 3606 2735 3610
rect 2739 3606 2740 3610
rect 2734 3605 2740 3606
rect 3022 3610 3028 3611
rect 3022 3606 3023 3610
rect 3027 3606 3028 3610
rect 3022 3605 3028 3606
rect 1830 3603 1836 3604
rect 110 3591 116 3592
rect 110 3587 111 3591
rect 115 3587 116 3591
rect 1830 3591 1836 3592
rect 110 3586 116 3587
rect 134 3588 140 3589
rect 134 3584 135 3588
rect 139 3584 140 3588
rect 134 3583 140 3584
rect 230 3588 236 3589
rect 230 3584 231 3588
rect 235 3584 236 3588
rect 230 3583 236 3584
rect 358 3588 364 3589
rect 358 3584 359 3588
rect 363 3584 364 3588
rect 358 3583 364 3584
rect 494 3588 500 3589
rect 494 3584 495 3588
rect 499 3584 500 3588
rect 494 3583 500 3584
rect 630 3588 636 3589
rect 630 3584 631 3588
rect 635 3584 636 3588
rect 630 3583 636 3584
rect 766 3588 772 3589
rect 766 3584 767 3588
rect 771 3584 772 3588
rect 766 3583 772 3584
rect 902 3588 908 3589
rect 902 3584 903 3588
rect 907 3584 908 3588
rect 902 3583 908 3584
rect 1046 3588 1052 3589
rect 1046 3584 1047 3588
rect 1051 3584 1052 3588
rect 1046 3583 1052 3584
rect 1190 3588 1196 3589
rect 1190 3584 1191 3588
rect 1195 3584 1196 3588
rect 1830 3587 1831 3591
rect 1835 3587 1836 3591
rect 1830 3586 1836 3587
rect 1190 3583 1196 3584
rect 1902 3578 1908 3579
rect 1902 3574 1903 3578
rect 1907 3574 1908 3578
rect 1902 3573 1908 3574
rect 1982 3578 1988 3579
rect 1982 3574 1983 3578
rect 1987 3574 1988 3578
rect 1982 3573 1988 3574
rect 2070 3578 2076 3579
rect 2070 3574 2071 3578
rect 2075 3574 2076 3578
rect 2070 3573 2076 3574
rect 2174 3578 2180 3579
rect 2174 3574 2175 3578
rect 2179 3574 2180 3578
rect 2174 3573 2180 3574
rect 2294 3578 2300 3579
rect 2294 3574 2295 3578
rect 2299 3574 2300 3578
rect 2294 3573 2300 3574
rect 2422 3578 2428 3579
rect 2422 3574 2423 3578
rect 2427 3574 2428 3578
rect 2422 3573 2428 3574
rect 2558 3578 2564 3579
rect 2558 3574 2559 3578
rect 2563 3574 2564 3578
rect 2558 3573 2564 3574
rect 2694 3578 2700 3579
rect 2694 3574 2695 3578
rect 2699 3574 2700 3578
rect 2694 3573 2700 3574
rect 2830 3578 2836 3579
rect 2830 3574 2831 3578
rect 2835 3574 2836 3578
rect 2830 3573 2836 3574
rect 2974 3578 2980 3579
rect 2974 3574 2975 3578
rect 2979 3574 2980 3578
rect 2974 3573 2980 3574
rect 3118 3578 3124 3579
rect 3118 3574 3119 3578
rect 3123 3574 3124 3578
rect 3118 3573 3124 3574
rect 3262 3578 3268 3579
rect 3262 3574 3263 3578
rect 3267 3574 3268 3578
rect 3262 3573 3268 3574
rect 1870 3560 1876 3561
rect 1870 3556 1871 3560
rect 1875 3556 1876 3560
rect 1870 3555 1876 3556
rect 3590 3560 3596 3561
rect 3590 3556 3591 3560
rect 3595 3556 3596 3560
rect 3590 3555 3596 3556
rect 182 3544 188 3545
rect 110 3541 116 3542
rect 110 3537 111 3541
rect 115 3537 116 3541
rect 182 3540 183 3544
rect 187 3540 188 3544
rect 182 3539 188 3540
rect 302 3544 308 3545
rect 302 3540 303 3544
rect 307 3540 308 3544
rect 302 3539 308 3540
rect 414 3544 420 3545
rect 414 3540 415 3544
rect 419 3540 420 3544
rect 414 3539 420 3540
rect 526 3544 532 3545
rect 526 3540 527 3544
rect 531 3540 532 3544
rect 526 3539 532 3540
rect 630 3544 636 3545
rect 630 3540 631 3544
rect 635 3540 636 3544
rect 630 3539 636 3540
rect 734 3544 740 3545
rect 734 3540 735 3544
rect 739 3540 740 3544
rect 734 3539 740 3540
rect 830 3544 836 3545
rect 830 3540 831 3544
rect 835 3540 836 3544
rect 830 3539 836 3540
rect 918 3544 924 3545
rect 918 3540 919 3544
rect 923 3540 924 3544
rect 918 3539 924 3540
rect 1006 3544 1012 3545
rect 1006 3540 1007 3544
rect 1011 3540 1012 3544
rect 1006 3539 1012 3540
rect 1094 3544 1100 3545
rect 1094 3540 1095 3544
rect 1099 3540 1100 3544
rect 1094 3539 1100 3540
rect 1182 3544 1188 3545
rect 1182 3540 1183 3544
rect 1187 3540 1188 3544
rect 1182 3539 1188 3540
rect 1270 3544 1276 3545
rect 1270 3540 1271 3544
rect 1275 3540 1276 3544
rect 1270 3539 1276 3540
rect 1358 3544 1364 3545
rect 1358 3540 1359 3544
rect 1363 3540 1364 3544
rect 1358 3539 1364 3540
rect 1446 3544 1452 3545
rect 1446 3540 1447 3544
rect 1451 3540 1452 3544
rect 1870 3543 1876 3544
rect 1446 3539 1452 3540
rect 1830 3541 1836 3542
rect 110 3536 116 3537
rect 1830 3537 1831 3541
rect 1835 3537 1836 3541
rect 1870 3539 1871 3543
rect 1875 3539 1876 3543
rect 3590 3543 3596 3544
rect 1870 3538 1876 3539
rect 1894 3540 1900 3541
rect 1830 3536 1836 3537
rect 1894 3536 1895 3540
rect 1899 3536 1900 3540
rect 1894 3535 1900 3536
rect 1974 3540 1980 3541
rect 1974 3536 1975 3540
rect 1979 3536 1980 3540
rect 1974 3535 1980 3536
rect 2062 3540 2068 3541
rect 2062 3536 2063 3540
rect 2067 3536 2068 3540
rect 2062 3535 2068 3536
rect 2166 3540 2172 3541
rect 2166 3536 2167 3540
rect 2171 3536 2172 3540
rect 2166 3535 2172 3536
rect 2286 3540 2292 3541
rect 2286 3536 2287 3540
rect 2291 3536 2292 3540
rect 2286 3535 2292 3536
rect 2414 3540 2420 3541
rect 2414 3536 2415 3540
rect 2419 3536 2420 3540
rect 2414 3535 2420 3536
rect 2550 3540 2556 3541
rect 2550 3536 2551 3540
rect 2555 3536 2556 3540
rect 2550 3535 2556 3536
rect 2686 3540 2692 3541
rect 2686 3536 2687 3540
rect 2691 3536 2692 3540
rect 2686 3535 2692 3536
rect 2822 3540 2828 3541
rect 2822 3536 2823 3540
rect 2827 3536 2828 3540
rect 2822 3535 2828 3536
rect 2966 3540 2972 3541
rect 2966 3536 2967 3540
rect 2971 3536 2972 3540
rect 2966 3535 2972 3536
rect 3110 3540 3116 3541
rect 3110 3536 3111 3540
rect 3115 3536 3116 3540
rect 3110 3535 3116 3536
rect 3254 3540 3260 3541
rect 3254 3536 3255 3540
rect 3259 3536 3260 3540
rect 3590 3539 3591 3543
rect 3595 3539 3596 3543
rect 3590 3538 3596 3539
rect 3254 3535 3260 3536
rect 110 3524 116 3525
rect 110 3520 111 3524
rect 115 3520 116 3524
rect 110 3519 116 3520
rect 1830 3524 1836 3525
rect 1830 3520 1831 3524
rect 1835 3520 1836 3524
rect 1830 3519 1836 3520
rect 190 3506 196 3507
rect 190 3502 191 3506
rect 195 3502 196 3506
rect 190 3501 196 3502
rect 310 3506 316 3507
rect 310 3502 311 3506
rect 315 3502 316 3506
rect 310 3501 316 3502
rect 422 3506 428 3507
rect 422 3502 423 3506
rect 427 3502 428 3506
rect 422 3501 428 3502
rect 534 3506 540 3507
rect 534 3502 535 3506
rect 539 3502 540 3506
rect 534 3501 540 3502
rect 638 3506 644 3507
rect 638 3502 639 3506
rect 643 3502 644 3506
rect 638 3501 644 3502
rect 742 3506 748 3507
rect 742 3502 743 3506
rect 747 3502 748 3506
rect 742 3501 748 3502
rect 838 3506 844 3507
rect 838 3502 839 3506
rect 843 3502 844 3506
rect 838 3501 844 3502
rect 926 3506 932 3507
rect 926 3502 927 3506
rect 931 3502 932 3506
rect 926 3501 932 3502
rect 1014 3506 1020 3507
rect 1014 3502 1015 3506
rect 1019 3502 1020 3506
rect 1014 3501 1020 3502
rect 1102 3506 1108 3507
rect 1102 3502 1103 3506
rect 1107 3502 1108 3506
rect 1102 3501 1108 3502
rect 1190 3506 1196 3507
rect 1190 3502 1191 3506
rect 1195 3502 1196 3506
rect 1190 3501 1196 3502
rect 1278 3506 1284 3507
rect 1278 3502 1279 3506
rect 1283 3502 1284 3506
rect 1278 3501 1284 3502
rect 1366 3506 1372 3507
rect 1366 3502 1367 3506
rect 1371 3502 1372 3506
rect 1366 3501 1372 3502
rect 1454 3506 1460 3507
rect 1454 3502 1455 3506
rect 1459 3502 1460 3506
rect 1454 3501 1460 3502
rect 1966 3496 1972 3497
rect 1870 3493 1876 3494
rect 1870 3489 1871 3493
rect 1875 3489 1876 3493
rect 1966 3492 1967 3496
rect 1971 3492 1972 3496
rect 1966 3491 1972 3492
rect 2150 3496 2156 3497
rect 2150 3492 2151 3496
rect 2155 3492 2156 3496
rect 2150 3491 2156 3492
rect 2334 3496 2340 3497
rect 2334 3492 2335 3496
rect 2339 3492 2340 3496
rect 2334 3491 2340 3492
rect 2510 3496 2516 3497
rect 2510 3492 2511 3496
rect 2515 3492 2516 3496
rect 2510 3491 2516 3492
rect 2670 3496 2676 3497
rect 2670 3492 2671 3496
rect 2675 3492 2676 3496
rect 2670 3491 2676 3492
rect 2822 3496 2828 3497
rect 2822 3492 2823 3496
rect 2827 3492 2828 3496
rect 2822 3491 2828 3492
rect 2958 3496 2964 3497
rect 2958 3492 2959 3496
rect 2963 3492 2964 3496
rect 2958 3491 2964 3492
rect 3078 3496 3084 3497
rect 3078 3492 3079 3496
rect 3083 3492 3084 3496
rect 3078 3491 3084 3492
rect 3190 3496 3196 3497
rect 3190 3492 3191 3496
rect 3195 3492 3196 3496
rect 3190 3491 3196 3492
rect 3302 3496 3308 3497
rect 3302 3492 3303 3496
rect 3307 3492 3308 3496
rect 3302 3491 3308 3492
rect 3414 3496 3420 3497
rect 3414 3492 3415 3496
rect 3419 3492 3420 3496
rect 3414 3491 3420 3492
rect 3502 3496 3508 3497
rect 3502 3492 3503 3496
rect 3507 3492 3508 3496
rect 3502 3491 3508 3492
rect 3590 3493 3596 3494
rect 1870 3488 1876 3489
rect 3590 3489 3591 3493
rect 3595 3489 3596 3493
rect 3590 3488 3596 3489
rect 1870 3476 1876 3477
rect 1870 3472 1871 3476
rect 1875 3472 1876 3476
rect 1870 3471 1876 3472
rect 3590 3476 3596 3477
rect 3590 3472 3591 3476
rect 3595 3472 3596 3476
rect 3590 3471 3596 3472
rect 230 3466 236 3467
rect 230 3462 231 3466
rect 235 3462 236 3466
rect 230 3461 236 3462
rect 366 3466 372 3467
rect 366 3462 367 3466
rect 371 3462 372 3466
rect 366 3461 372 3462
rect 502 3466 508 3467
rect 502 3462 503 3466
rect 507 3462 508 3466
rect 502 3461 508 3462
rect 622 3466 628 3467
rect 622 3462 623 3466
rect 627 3462 628 3466
rect 622 3461 628 3462
rect 734 3466 740 3467
rect 734 3462 735 3466
rect 739 3462 740 3466
rect 734 3461 740 3462
rect 838 3466 844 3467
rect 838 3462 839 3466
rect 843 3462 844 3466
rect 838 3461 844 3462
rect 942 3466 948 3467
rect 942 3462 943 3466
rect 947 3462 948 3466
rect 942 3461 948 3462
rect 1038 3466 1044 3467
rect 1038 3462 1039 3466
rect 1043 3462 1044 3466
rect 1038 3461 1044 3462
rect 1134 3466 1140 3467
rect 1134 3462 1135 3466
rect 1139 3462 1140 3466
rect 1134 3461 1140 3462
rect 1230 3466 1236 3467
rect 1230 3462 1231 3466
rect 1235 3462 1236 3466
rect 1230 3461 1236 3462
rect 1326 3466 1332 3467
rect 1326 3462 1327 3466
rect 1331 3462 1332 3466
rect 1326 3461 1332 3462
rect 1974 3458 1980 3459
rect 1974 3454 1975 3458
rect 1979 3454 1980 3458
rect 1974 3453 1980 3454
rect 2158 3458 2164 3459
rect 2158 3454 2159 3458
rect 2163 3454 2164 3458
rect 2158 3453 2164 3454
rect 2342 3458 2348 3459
rect 2342 3454 2343 3458
rect 2347 3454 2348 3458
rect 2342 3453 2348 3454
rect 2518 3458 2524 3459
rect 2518 3454 2519 3458
rect 2523 3454 2524 3458
rect 2518 3453 2524 3454
rect 2678 3458 2684 3459
rect 2678 3454 2679 3458
rect 2683 3454 2684 3458
rect 2678 3453 2684 3454
rect 2830 3458 2836 3459
rect 2830 3454 2831 3458
rect 2835 3454 2836 3458
rect 2830 3453 2836 3454
rect 2966 3458 2972 3459
rect 2966 3454 2967 3458
rect 2971 3454 2972 3458
rect 2966 3453 2972 3454
rect 3086 3458 3092 3459
rect 3086 3454 3087 3458
rect 3091 3454 3092 3458
rect 3086 3453 3092 3454
rect 3198 3458 3204 3459
rect 3198 3454 3199 3458
rect 3203 3454 3204 3458
rect 3198 3453 3204 3454
rect 3310 3458 3316 3459
rect 3310 3454 3311 3458
rect 3315 3454 3316 3458
rect 3310 3453 3316 3454
rect 3422 3458 3428 3459
rect 3422 3454 3423 3458
rect 3427 3454 3428 3458
rect 3422 3453 3428 3454
rect 3510 3458 3516 3459
rect 3510 3454 3511 3458
rect 3515 3454 3516 3458
rect 3510 3453 3516 3454
rect 110 3448 116 3449
rect 110 3444 111 3448
rect 115 3444 116 3448
rect 110 3443 116 3444
rect 1830 3448 1836 3449
rect 1830 3444 1831 3448
rect 1835 3444 1836 3448
rect 1830 3443 1836 3444
rect 110 3431 116 3432
rect 110 3427 111 3431
rect 115 3427 116 3431
rect 1830 3431 1836 3432
rect 110 3426 116 3427
rect 222 3428 228 3429
rect 222 3424 223 3428
rect 227 3424 228 3428
rect 222 3423 228 3424
rect 358 3428 364 3429
rect 358 3424 359 3428
rect 363 3424 364 3428
rect 358 3423 364 3424
rect 494 3428 500 3429
rect 494 3424 495 3428
rect 499 3424 500 3428
rect 494 3423 500 3424
rect 614 3428 620 3429
rect 614 3424 615 3428
rect 619 3424 620 3428
rect 614 3423 620 3424
rect 726 3428 732 3429
rect 726 3424 727 3428
rect 731 3424 732 3428
rect 726 3423 732 3424
rect 830 3428 836 3429
rect 830 3424 831 3428
rect 835 3424 836 3428
rect 830 3423 836 3424
rect 934 3428 940 3429
rect 934 3424 935 3428
rect 939 3424 940 3428
rect 934 3423 940 3424
rect 1030 3428 1036 3429
rect 1030 3424 1031 3428
rect 1035 3424 1036 3428
rect 1030 3423 1036 3424
rect 1126 3428 1132 3429
rect 1126 3424 1127 3428
rect 1131 3424 1132 3428
rect 1126 3423 1132 3424
rect 1222 3428 1228 3429
rect 1222 3424 1223 3428
rect 1227 3424 1228 3428
rect 1222 3423 1228 3424
rect 1318 3428 1324 3429
rect 1318 3424 1319 3428
rect 1323 3424 1324 3428
rect 1830 3427 1831 3431
rect 1835 3427 1836 3431
rect 1830 3426 1836 3427
rect 2006 3426 2012 3427
rect 1318 3423 1324 3424
rect 2006 3422 2007 3426
rect 2011 3422 2012 3426
rect 2006 3421 2012 3422
rect 2126 3426 2132 3427
rect 2126 3422 2127 3426
rect 2131 3422 2132 3426
rect 2126 3421 2132 3422
rect 2254 3426 2260 3427
rect 2254 3422 2255 3426
rect 2259 3422 2260 3426
rect 2254 3421 2260 3422
rect 2390 3426 2396 3427
rect 2390 3422 2391 3426
rect 2395 3422 2396 3426
rect 2390 3421 2396 3422
rect 2534 3426 2540 3427
rect 2534 3422 2535 3426
rect 2539 3422 2540 3426
rect 2534 3421 2540 3422
rect 2678 3426 2684 3427
rect 2678 3422 2679 3426
rect 2683 3422 2684 3426
rect 2678 3421 2684 3422
rect 2830 3426 2836 3427
rect 2830 3422 2831 3426
rect 2835 3422 2836 3426
rect 2830 3421 2836 3422
rect 2998 3426 3004 3427
rect 2998 3422 2999 3426
rect 3003 3422 3004 3426
rect 2998 3421 3004 3422
rect 3166 3426 3172 3427
rect 3166 3422 3167 3426
rect 3171 3422 3172 3426
rect 3166 3421 3172 3422
rect 3342 3426 3348 3427
rect 3342 3422 3343 3426
rect 3347 3422 3348 3426
rect 3342 3421 3348 3422
rect 3510 3426 3516 3427
rect 3510 3422 3511 3426
rect 3515 3422 3516 3426
rect 3510 3421 3516 3422
rect 1870 3408 1876 3409
rect 1870 3404 1871 3408
rect 1875 3404 1876 3408
rect 1870 3403 1876 3404
rect 3590 3408 3596 3409
rect 3590 3404 3591 3408
rect 3595 3404 3596 3408
rect 3590 3403 3596 3404
rect 1870 3391 1876 3392
rect 1870 3387 1871 3391
rect 1875 3387 1876 3391
rect 3590 3391 3596 3392
rect 1870 3386 1876 3387
rect 1998 3388 2004 3389
rect 1998 3384 1999 3388
rect 2003 3384 2004 3388
rect 1998 3383 2004 3384
rect 2118 3388 2124 3389
rect 2118 3384 2119 3388
rect 2123 3384 2124 3388
rect 2118 3383 2124 3384
rect 2246 3388 2252 3389
rect 2246 3384 2247 3388
rect 2251 3384 2252 3388
rect 2246 3383 2252 3384
rect 2382 3388 2388 3389
rect 2382 3384 2383 3388
rect 2387 3384 2388 3388
rect 2382 3383 2388 3384
rect 2526 3388 2532 3389
rect 2526 3384 2527 3388
rect 2531 3384 2532 3388
rect 2526 3383 2532 3384
rect 2670 3388 2676 3389
rect 2670 3384 2671 3388
rect 2675 3384 2676 3388
rect 2670 3383 2676 3384
rect 2822 3388 2828 3389
rect 2822 3384 2823 3388
rect 2827 3384 2828 3388
rect 2822 3383 2828 3384
rect 2990 3388 2996 3389
rect 2990 3384 2991 3388
rect 2995 3384 2996 3388
rect 2990 3383 2996 3384
rect 3158 3388 3164 3389
rect 3158 3384 3159 3388
rect 3163 3384 3164 3388
rect 3158 3383 3164 3384
rect 3334 3388 3340 3389
rect 3334 3384 3335 3388
rect 3339 3384 3340 3388
rect 3334 3383 3340 3384
rect 3502 3388 3508 3389
rect 3502 3384 3503 3388
rect 3507 3384 3508 3388
rect 3590 3387 3591 3391
rect 3595 3387 3596 3391
rect 3590 3386 3596 3387
rect 3502 3383 3508 3384
rect 214 3380 220 3381
rect 110 3377 116 3378
rect 110 3373 111 3377
rect 115 3373 116 3377
rect 214 3376 215 3380
rect 219 3376 220 3380
rect 214 3375 220 3376
rect 366 3380 372 3381
rect 366 3376 367 3380
rect 371 3376 372 3380
rect 366 3375 372 3376
rect 510 3380 516 3381
rect 510 3376 511 3380
rect 515 3376 516 3380
rect 510 3375 516 3376
rect 646 3380 652 3381
rect 646 3376 647 3380
rect 651 3376 652 3380
rect 646 3375 652 3376
rect 774 3380 780 3381
rect 774 3376 775 3380
rect 779 3376 780 3380
rect 774 3375 780 3376
rect 894 3380 900 3381
rect 894 3376 895 3380
rect 899 3376 900 3380
rect 894 3375 900 3376
rect 1014 3380 1020 3381
rect 1014 3376 1015 3380
rect 1019 3376 1020 3380
rect 1014 3375 1020 3376
rect 1126 3380 1132 3381
rect 1126 3376 1127 3380
rect 1131 3376 1132 3380
rect 1126 3375 1132 3376
rect 1238 3380 1244 3381
rect 1238 3376 1239 3380
rect 1243 3376 1244 3380
rect 1238 3375 1244 3376
rect 1350 3380 1356 3381
rect 1350 3376 1351 3380
rect 1355 3376 1356 3380
rect 1350 3375 1356 3376
rect 1830 3377 1836 3378
rect 110 3372 116 3373
rect 1830 3373 1831 3377
rect 1835 3373 1836 3377
rect 1830 3372 1836 3373
rect 110 3360 116 3361
rect 110 3356 111 3360
rect 115 3356 116 3360
rect 110 3355 116 3356
rect 1830 3360 1836 3361
rect 1830 3356 1831 3360
rect 1835 3356 1836 3360
rect 1830 3355 1836 3356
rect 2014 3344 2020 3345
rect 222 3342 228 3343
rect 222 3338 223 3342
rect 227 3338 228 3342
rect 222 3337 228 3338
rect 374 3342 380 3343
rect 374 3338 375 3342
rect 379 3338 380 3342
rect 374 3337 380 3338
rect 518 3342 524 3343
rect 518 3338 519 3342
rect 523 3338 524 3342
rect 518 3337 524 3338
rect 654 3342 660 3343
rect 654 3338 655 3342
rect 659 3338 660 3342
rect 654 3337 660 3338
rect 782 3342 788 3343
rect 782 3338 783 3342
rect 787 3338 788 3342
rect 782 3337 788 3338
rect 902 3342 908 3343
rect 902 3338 903 3342
rect 907 3338 908 3342
rect 902 3337 908 3338
rect 1022 3342 1028 3343
rect 1022 3338 1023 3342
rect 1027 3338 1028 3342
rect 1022 3337 1028 3338
rect 1134 3342 1140 3343
rect 1134 3338 1135 3342
rect 1139 3338 1140 3342
rect 1134 3337 1140 3338
rect 1246 3342 1252 3343
rect 1246 3338 1247 3342
rect 1251 3338 1252 3342
rect 1246 3337 1252 3338
rect 1358 3342 1364 3343
rect 1358 3338 1359 3342
rect 1363 3338 1364 3342
rect 1358 3337 1364 3338
rect 1870 3341 1876 3342
rect 1870 3337 1871 3341
rect 1875 3337 1876 3341
rect 2014 3340 2015 3344
rect 2019 3340 2020 3344
rect 2014 3339 2020 3340
rect 2150 3344 2156 3345
rect 2150 3340 2151 3344
rect 2155 3340 2156 3344
rect 2150 3339 2156 3340
rect 2294 3344 2300 3345
rect 2294 3340 2295 3344
rect 2299 3340 2300 3344
rect 2294 3339 2300 3340
rect 2438 3344 2444 3345
rect 2438 3340 2439 3344
rect 2443 3340 2444 3344
rect 2438 3339 2444 3340
rect 2582 3344 2588 3345
rect 2582 3340 2583 3344
rect 2587 3340 2588 3344
rect 2582 3339 2588 3340
rect 2726 3344 2732 3345
rect 2726 3340 2727 3344
rect 2731 3340 2732 3344
rect 2726 3339 2732 3340
rect 2870 3344 2876 3345
rect 2870 3340 2871 3344
rect 2875 3340 2876 3344
rect 2870 3339 2876 3340
rect 3022 3344 3028 3345
rect 3022 3340 3023 3344
rect 3027 3340 3028 3344
rect 3022 3339 3028 3340
rect 3182 3344 3188 3345
rect 3182 3340 3183 3344
rect 3187 3340 3188 3344
rect 3182 3339 3188 3340
rect 3350 3344 3356 3345
rect 3350 3340 3351 3344
rect 3355 3340 3356 3344
rect 3350 3339 3356 3340
rect 3502 3344 3508 3345
rect 3502 3340 3503 3344
rect 3507 3340 3508 3344
rect 3502 3339 3508 3340
rect 3590 3341 3596 3342
rect 1870 3336 1876 3337
rect 3590 3337 3591 3341
rect 3595 3337 3596 3341
rect 3590 3336 3596 3337
rect 1870 3324 1876 3325
rect 1870 3320 1871 3324
rect 1875 3320 1876 3324
rect 1870 3319 1876 3320
rect 3590 3324 3596 3325
rect 3590 3320 3591 3324
rect 3595 3320 3596 3324
rect 3590 3319 3596 3320
rect 206 3306 212 3307
rect 206 3302 207 3306
rect 211 3302 212 3306
rect 206 3301 212 3302
rect 366 3306 372 3307
rect 366 3302 367 3306
rect 371 3302 372 3306
rect 366 3301 372 3302
rect 518 3306 524 3307
rect 518 3302 519 3306
rect 523 3302 524 3306
rect 518 3301 524 3302
rect 670 3306 676 3307
rect 670 3302 671 3306
rect 675 3302 676 3306
rect 670 3301 676 3302
rect 814 3306 820 3307
rect 814 3302 815 3306
rect 819 3302 820 3306
rect 814 3301 820 3302
rect 950 3306 956 3307
rect 950 3302 951 3306
rect 955 3302 956 3306
rect 950 3301 956 3302
rect 1086 3306 1092 3307
rect 1086 3302 1087 3306
rect 1091 3302 1092 3306
rect 1086 3301 1092 3302
rect 1214 3306 1220 3307
rect 1214 3302 1215 3306
rect 1219 3302 1220 3306
rect 1214 3301 1220 3302
rect 1342 3306 1348 3307
rect 1342 3302 1343 3306
rect 1347 3302 1348 3306
rect 1342 3301 1348 3302
rect 1470 3306 1476 3307
rect 1470 3302 1471 3306
rect 1475 3302 1476 3306
rect 1470 3301 1476 3302
rect 2022 3306 2028 3307
rect 2022 3302 2023 3306
rect 2027 3302 2028 3306
rect 2022 3301 2028 3302
rect 2158 3306 2164 3307
rect 2158 3302 2159 3306
rect 2163 3302 2164 3306
rect 2158 3301 2164 3302
rect 2302 3306 2308 3307
rect 2302 3302 2303 3306
rect 2307 3302 2308 3306
rect 2302 3301 2308 3302
rect 2446 3306 2452 3307
rect 2446 3302 2447 3306
rect 2451 3302 2452 3306
rect 2446 3301 2452 3302
rect 2590 3306 2596 3307
rect 2590 3302 2591 3306
rect 2595 3302 2596 3306
rect 2590 3301 2596 3302
rect 2734 3306 2740 3307
rect 2734 3302 2735 3306
rect 2739 3302 2740 3306
rect 2734 3301 2740 3302
rect 2878 3306 2884 3307
rect 2878 3302 2879 3306
rect 2883 3302 2884 3306
rect 2878 3301 2884 3302
rect 3030 3306 3036 3307
rect 3030 3302 3031 3306
rect 3035 3302 3036 3306
rect 3030 3301 3036 3302
rect 3190 3306 3196 3307
rect 3190 3302 3191 3306
rect 3195 3302 3196 3306
rect 3190 3301 3196 3302
rect 3358 3306 3364 3307
rect 3358 3302 3359 3306
rect 3363 3302 3364 3306
rect 3358 3301 3364 3302
rect 3510 3306 3516 3307
rect 3510 3302 3511 3306
rect 3515 3302 3516 3306
rect 3510 3301 3516 3302
rect 110 3288 116 3289
rect 110 3284 111 3288
rect 115 3284 116 3288
rect 110 3283 116 3284
rect 1830 3288 1836 3289
rect 1830 3284 1831 3288
rect 1835 3284 1836 3288
rect 1830 3283 1836 3284
rect 1926 3274 1932 3275
rect 110 3271 116 3272
rect 110 3267 111 3271
rect 115 3267 116 3271
rect 1830 3271 1836 3272
rect 110 3266 116 3267
rect 198 3268 204 3269
rect 198 3264 199 3268
rect 203 3264 204 3268
rect 198 3263 204 3264
rect 358 3268 364 3269
rect 358 3264 359 3268
rect 363 3264 364 3268
rect 358 3263 364 3264
rect 510 3268 516 3269
rect 510 3264 511 3268
rect 515 3264 516 3268
rect 510 3263 516 3264
rect 662 3268 668 3269
rect 662 3264 663 3268
rect 667 3264 668 3268
rect 662 3263 668 3264
rect 806 3268 812 3269
rect 806 3264 807 3268
rect 811 3264 812 3268
rect 806 3263 812 3264
rect 942 3268 948 3269
rect 942 3264 943 3268
rect 947 3264 948 3268
rect 942 3263 948 3264
rect 1078 3268 1084 3269
rect 1078 3264 1079 3268
rect 1083 3264 1084 3268
rect 1078 3263 1084 3264
rect 1206 3268 1212 3269
rect 1206 3264 1207 3268
rect 1211 3264 1212 3268
rect 1206 3263 1212 3264
rect 1334 3268 1340 3269
rect 1334 3264 1335 3268
rect 1339 3264 1340 3268
rect 1334 3263 1340 3264
rect 1462 3268 1468 3269
rect 1462 3264 1463 3268
rect 1467 3264 1468 3268
rect 1830 3267 1831 3271
rect 1835 3267 1836 3271
rect 1926 3270 1927 3274
rect 1931 3270 1932 3274
rect 1926 3269 1932 3270
rect 2062 3274 2068 3275
rect 2062 3270 2063 3274
rect 2067 3270 2068 3274
rect 2062 3269 2068 3270
rect 2190 3274 2196 3275
rect 2190 3270 2191 3274
rect 2195 3270 2196 3274
rect 2190 3269 2196 3270
rect 2318 3274 2324 3275
rect 2318 3270 2319 3274
rect 2323 3270 2324 3274
rect 2318 3269 2324 3270
rect 2446 3274 2452 3275
rect 2446 3270 2447 3274
rect 2451 3270 2452 3274
rect 2446 3269 2452 3270
rect 2590 3274 2596 3275
rect 2590 3270 2591 3274
rect 2595 3270 2596 3274
rect 2590 3269 2596 3270
rect 2742 3274 2748 3275
rect 2742 3270 2743 3274
rect 2747 3270 2748 3274
rect 2742 3269 2748 3270
rect 2918 3274 2924 3275
rect 2918 3270 2919 3274
rect 2923 3270 2924 3274
rect 2918 3269 2924 3270
rect 3110 3274 3116 3275
rect 3110 3270 3111 3274
rect 3115 3270 3116 3274
rect 3110 3269 3116 3270
rect 3310 3274 3316 3275
rect 3310 3270 3311 3274
rect 3315 3270 3316 3274
rect 3310 3269 3316 3270
rect 3510 3274 3516 3275
rect 3510 3270 3511 3274
rect 3515 3270 3516 3274
rect 3510 3269 3516 3270
rect 1830 3266 1836 3267
rect 1462 3263 1468 3264
rect 1870 3256 1876 3257
rect 1870 3252 1871 3256
rect 1875 3252 1876 3256
rect 1870 3251 1876 3252
rect 3590 3256 3596 3257
rect 3590 3252 3591 3256
rect 3595 3252 3596 3256
rect 3590 3251 3596 3252
rect 1870 3239 1876 3240
rect 1870 3235 1871 3239
rect 1875 3235 1876 3239
rect 3590 3239 3596 3240
rect 1870 3234 1876 3235
rect 1918 3236 1924 3237
rect 1918 3232 1919 3236
rect 1923 3232 1924 3236
rect 1918 3231 1924 3232
rect 2054 3236 2060 3237
rect 2054 3232 2055 3236
rect 2059 3232 2060 3236
rect 2054 3231 2060 3232
rect 2182 3236 2188 3237
rect 2182 3232 2183 3236
rect 2187 3232 2188 3236
rect 2182 3231 2188 3232
rect 2310 3236 2316 3237
rect 2310 3232 2311 3236
rect 2315 3232 2316 3236
rect 2310 3231 2316 3232
rect 2438 3236 2444 3237
rect 2438 3232 2439 3236
rect 2443 3232 2444 3236
rect 2438 3231 2444 3232
rect 2582 3236 2588 3237
rect 2582 3232 2583 3236
rect 2587 3232 2588 3236
rect 2582 3231 2588 3232
rect 2734 3236 2740 3237
rect 2734 3232 2735 3236
rect 2739 3232 2740 3236
rect 2734 3231 2740 3232
rect 2910 3236 2916 3237
rect 2910 3232 2911 3236
rect 2915 3232 2916 3236
rect 2910 3231 2916 3232
rect 3102 3236 3108 3237
rect 3102 3232 3103 3236
rect 3107 3232 3108 3236
rect 3102 3231 3108 3232
rect 3302 3236 3308 3237
rect 3302 3232 3303 3236
rect 3307 3232 3308 3236
rect 3302 3231 3308 3232
rect 3502 3236 3508 3237
rect 3502 3232 3503 3236
rect 3507 3232 3508 3236
rect 3590 3235 3591 3239
rect 3595 3235 3596 3239
rect 3590 3234 3596 3235
rect 3502 3231 3508 3232
rect 134 3224 140 3225
rect 110 3221 116 3222
rect 110 3217 111 3221
rect 115 3217 116 3221
rect 134 3220 135 3224
rect 139 3220 140 3224
rect 134 3219 140 3220
rect 270 3224 276 3225
rect 270 3220 271 3224
rect 275 3220 276 3224
rect 270 3219 276 3220
rect 414 3224 420 3225
rect 414 3220 415 3224
rect 419 3220 420 3224
rect 414 3219 420 3220
rect 574 3224 580 3225
rect 574 3220 575 3224
rect 579 3220 580 3224
rect 574 3219 580 3220
rect 734 3224 740 3225
rect 734 3220 735 3224
rect 739 3220 740 3224
rect 734 3219 740 3220
rect 894 3224 900 3225
rect 894 3220 895 3224
rect 899 3220 900 3224
rect 894 3219 900 3220
rect 1046 3224 1052 3225
rect 1046 3220 1047 3224
rect 1051 3220 1052 3224
rect 1046 3219 1052 3220
rect 1190 3224 1196 3225
rect 1190 3220 1191 3224
rect 1195 3220 1196 3224
rect 1190 3219 1196 3220
rect 1326 3224 1332 3225
rect 1326 3220 1327 3224
rect 1331 3220 1332 3224
rect 1326 3219 1332 3220
rect 1462 3224 1468 3225
rect 1462 3220 1463 3224
rect 1467 3220 1468 3224
rect 1462 3219 1468 3220
rect 1606 3224 1612 3225
rect 1606 3220 1607 3224
rect 1611 3220 1612 3224
rect 1606 3219 1612 3220
rect 1830 3221 1836 3222
rect 110 3216 116 3217
rect 1830 3217 1831 3221
rect 1835 3217 1836 3221
rect 1830 3216 1836 3217
rect 110 3204 116 3205
rect 110 3200 111 3204
rect 115 3200 116 3204
rect 110 3199 116 3200
rect 1830 3204 1836 3205
rect 1830 3200 1831 3204
rect 1835 3200 1836 3204
rect 1830 3199 1836 3200
rect 1894 3192 1900 3193
rect 1870 3189 1876 3190
rect 142 3186 148 3187
rect 142 3182 143 3186
rect 147 3182 148 3186
rect 142 3181 148 3182
rect 278 3186 284 3187
rect 278 3182 279 3186
rect 283 3182 284 3186
rect 278 3181 284 3182
rect 422 3186 428 3187
rect 422 3182 423 3186
rect 427 3182 428 3186
rect 422 3181 428 3182
rect 582 3186 588 3187
rect 582 3182 583 3186
rect 587 3182 588 3186
rect 582 3181 588 3182
rect 742 3186 748 3187
rect 742 3182 743 3186
rect 747 3182 748 3186
rect 742 3181 748 3182
rect 902 3186 908 3187
rect 902 3182 903 3186
rect 907 3182 908 3186
rect 902 3181 908 3182
rect 1054 3186 1060 3187
rect 1054 3182 1055 3186
rect 1059 3182 1060 3186
rect 1054 3181 1060 3182
rect 1198 3186 1204 3187
rect 1198 3182 1199 3186
rect 1203 3182 1204 3186
rect 1198 3181 1204 3182
rect 1334 3186 1340 3187
rect 1334 3182 1335 3186
rect 1339 3182 1340 3186
rect 1334 3181 1340 3182
rect 1470 3186 1476 3187
rect 1470 3182 1471 3186
rect 1475 3182 1476 3186
rect 1470 3181 1476 3182
rect 1614 3186 1620 3187
rect 1614 3182 1615 3186
rect 1619 3182 1620 3186
rect 1870 3185 1871 3189
rect 1875 3185 1876 3189
rect 1894 3188 1895 3192
rect 1899 3188 1900 3192
rect 1894 3187 1900 3188
rect 2006 3192 2012 3193
rect 2006 3188 2007 3192
rect 2011 3188 2012 3192
rect 2006 3187 2012 3188
rect 2142 3192 2148 3193
rect 2142 3188 2143 3192
rect 2147 3188 2148 3192
rect 2142 3187 2148 3188
rect 2294 3192 2300 3193
rect 2294 3188 2295 3192
rect 2299 3188 2300 3192
rect 2294 3187 2300 3188
rect 2454 3192 2460 3193
rect 2454 3188 2455 3192
rect 2459 3188 2460 3192
rect 2454 3187 2460 3188
rect 2622 3192 2628 3193
rect 2622 3188 2623 3192
rect 2627 3188 2628 3192
rect 2622 3187 2628 3188
rect 2798 3192 2804 3193
rect 2798 3188 2799 3192
rect 2803 3188 2804 3192
rect 2798 3187 2804 3188
rect 2974 3192 2980 3193
rect 2974 3188 2975 3192
rect 2979 3188 2980 3192
rect 2974 3187 2980 3188
rect 3150 3192 3156 3193
rect 3150 3188 3151 3192
rect 3155 3188 3156 3192
rect 3150 3187 3156 3188
rect 3326 3192 3332 3193
rect 3326 3188 3327 3192
rect 3331 3188 3332 3192
rect 3326 3187 3332 3188
rect 3502 3192 3508 3193
rect 3502 3188 3503 3192
rect 3507 3188 3508 3192
rect 3502 3187 3508 3188
rect 3590 3189 3596 3190
rect 1870 3184 1876 3185
rect 3590 3185 3591 3189
rect 3595 3185 3596 3189
rect 3590 3184 3596 3185
rect 1614 3181 1620 3182
rect 1870 3172 1876 3173
rect 1870 3168 1871 3172
rect 1875 3168 1876 3172
rect 1870 3167 1876 3168
rect 3590 3172 3596 3173
rect 3590 3168 3591 3172
rect 3595 3168 3596 3172
rect 3590 3167 3596 3168
rect 1902 3154 1908 3155
rect 1902 3150 1903 3154
rect 1907 3150 1908 3154
rect 1902 3149 1908 3150
rect 2014 3154 2020 3155
rect 2014 3150 2015 3154
rect 2019 3150 2020 3154
rect 2014 3149 2020 3150
rect 2150 3154 2156 3155
rect 2150 3150 2151 3154
rect 2155 3150 2156 3154
rect 2150 3149 2156 3150
rect 2302 3154 2308 3155
rect 2302 3150 2303 3154
rect 2307 3150 2308 3154
rect 2302 3149 2308 3150
rect 2462 3154 2468 3155
rect 2462 3150 2463 3154
rect 2467 3150 2468 3154
rect 2462 3149 2468 3150
rect 2630 3154 2636 3155
rect 2630 3150 2631 3154
rect 2635 3150 2636 3154
rect 2630 3149 2636 3150
rect 2806 3154 2812 3155
rect 2806 3150 2807 3154
rect 2811 3150 2812 3154
rect 2806 3149 2812 3150
rect 2982 3154 2988 3155
rect 2982 3150 2983 3154
rect 2987 3150 2988 3154
rect 2982 3149 2988 3150
rect 3158 3154 3164 3155
rect 3158 3150 3159 3154
rect 3163 3150 3164 3154
rect 3158 3149 3164 3150
rect 3334 3154 3340 3155
rect 3334 3150 3335 3154
rect 3339 3150 3340 3154
rect 3334 3149 3340 3150
rect 3510 3154 3516 3155
rect 3510 3150 3511 3154
rect 3515 3150 3516 3154
rect 3510 3149 3516 3150
rect 174 3146 180 3147
rect 174 3142 175 3146
rect 179 3142 180 3146
rect 174 3141 180 3142
rect 318 3146 324 3147
rect 318 3142 319 3146
rect 323 3142 324 3146
rect 318 3141 324 3142
rect 462 3146 468 3147
rect 462 3142 463 3146
rect 467 3142 468 3146
rect 462 3141 468 3142
rect 606 3146 612 3147
rect 606 3142 607 3146
rect 611 3142 612 3146
rect 606 3141 612 3142
rect 742 3146 748 3147
rect 742 3142 743 3146
rect 747 3142 748 3146
rect 742 3141 748 3142
rect 870 3146 876 3147
rect 870 3142 871 3146
rect 875 3142 876 3146
rect 870 3141 876 3142
rect 990 3146 996 3147
rect 990 3142 991 3146
rect 995 3142 996 3146
rect 990 3141 996 3142
rect 1102 3146 1108 3147
rect 1102 3142 1103 3146
rect 1107 3142 1108 3146
rect 1102 3141 1108 3142
rect 1206 3146 1212 3147
rect 1206 3142 1207 3146
rect 1211 3142 1212 3146
rect 1206 3141 1212 3142
rect 1310 3146 1316 3147
rect 1310 3142 1311 3146
rect 1315 3142 1316 3146
rect 1310 3141 1316 3142
rect 1406 3146 1412 3147
rect 1406 3142 1407 3146
rect 1411 3142 1412 3146
rect 1406 3141 1412 3142
rect 1494 3146 1500 3147
rect 1494 3142 1495 3146
rect 1499 3142 1500 3146
rect 1494 3141 1500 3142
rect 1582 3146 1588 3147
rect 1582 3142 1583 3146
rect 1587 3142 1588 3146
rect 1582 3141 1588 3142
rect 1670 3146 1676 3147
rect 1670 3142 1671 3146
rect 1675 3142 1676 3146
rect 1670 3141 1676 3142
rect 1750 3146 1756 3147
rect 1750 3142 1751 3146
rect 1755 3142 1756 3146
rect 1750 3141 1756 3142
rect 110 3128 116 3129
rect 110 3124 111 3128
rect 115 3124 116 3128
rect 110 3123 116 3124
rect 1830 3128 1836 3129
rect 1830 3124 1831 3128
rect 1835 3124 1836 3128
rect 1830 3123 1836 3124
rect 1902 3122 1908 3123
rect 1902 3118 1903 3122
rect 1907 3118 1908 3122
rect 1902 3117 1908 3118
rect 2070 3122 2076 3123
rect 2070 3118 2071 3122
rect 2075 3118 2076 3122
rect 2070 3117 2076 3118
rect 2262 3122 2268 3123
rect 2262 3118 2263 3122
rect 2267 3118 2268 3122
rect 2262 3117 2268 3118
rect 2454 3122 2460 3123
rect 2454 3118 2455 3122
rect 2459 3118 2460 3122
rect 2454 3117 2460 3118
rect 2646 3122 2652 3123
rect 2646 3118 2647 3122
rect 2651 3118 2652 3122
rect 2646 3117 2652 3118
rect 2830 3122 2836 3123
rect 2830 3118 2831 3122
rect 2835 3118 2836 3122
rect 2830 3117 2836 3118
rect 3014 3122 3020 3123
rect 3014 3118 3015 3122
rect 3019 3118 3020 3122
rect 3014 3117 3020 3118
rect 3198 3122 3204 3123
rect 3198 3118 3199 3122
rect 3203 3118 3204 3122
rect 3198 3117 3204 3118
rect 3390 3122 3396 3123
rect 3390 3118 3391 3122
rect 3395 3118 3396 3122
rect 3390 3117 3396 3118
rect 110 3111 116 3112
rect 110 3107 111 3111
rect 115 3107 116 3111
rect 1830 3111 1836 3112
rect 110 3106 116 3107
rect 166 3108 172 3109
rect 166 3104 167 3108
rect 171 3104 172 3108
rect 166 3103 172 3104
rect 310 3108 316 3109
rect 310 3104 311 3108
rect 315 3104 316 3108
rect 310 3103 316 3104
rect 454 3108 460 3109
rect 454 3104 455 3108
rect 459 3104 460 3108
rect 454 3103 460 3104
rect 598 3108 604 3109
rect 598 3104 599 3108
rect 603 3104 604 3108
rect 598 3103 604 3104
rect 734 3108 740 3109
rect 734 3104 735 3108
rect 739 3104 740 3108
rect 734 3103 740 3104
rect 862 3108 868 3109
rect 862 3104 863 3108
rect 867 3104 868 3108
rect 862 3103 868 3104
rect 982 3108 988 3109
rect 982 3104 983 3108
rect 987 3104 988 3108
rect 982 3103 988 3104
rect 1094 3108 1100 3109
rect 1094 3104 1095 3108
rect 1099 3104 1100 3108
rect 1094 3103 1100 3104
rect 1198 3108 1204 3109
rect 1198 3104 1199 3108
rect 1203 3104 1204 3108
rect 1198 3103 1204 3104
rect 1302 3108 1308 3109
rect 1302 3104 1303 3108
rect 1307 3104 1308 3108
rect 1302 3103 1308 3104
rect 1398 3108 1404 3109
rect 1398 3104 1399 3108
rect 1403 3104 1404 3108
rect 1398 3103 1404 3104
rect 1486 3108 1492 3109
rect 1486 3104 1487 3108
rect 1491 3104 1492 3108
rect 1486 3103 1492 3104
rect 1574 3108 1580 3109
rect 1574 3104 1575 3108
rect 1579 3104 1580 3108
rect 1574 3103 1580 3104
rect 1662 3108 1668 3109
rect 1662 3104 1663 3108
rect 1667 3104 1668 3108
rect 1662 3103 1668 3104
rect 1742 3108 1748 3109
rect 1742 3104 1743 3108
rect 1747 3104 1748 3108
rect 1830 3107 1831 3111
rect 1835 3107 1836 3111
rect 1830 3106 1836 3107
rect 1742 3103 1748 3104
rect 1870 3104 1876 3105
rect 1870 3100 1871 3104
rect 1875 3100 1876 3104
rect 1870 3099 1876 3100
rect 3590 3104 3596 3105
rect 3590 3100 3591 3104
rect 3595 3100 3596 3104
rect 3590 3099 3596 3100
rect 1870 3087 1876 3088
rect 1870 3083 1871 3087
rect 1875 3083 1876 3087
rect 3590 3087 3596 3088
rect 1870 3082 1876 3083
rect 1894 3084 1900 3085
rect 1894 3080 1895 3084
rect 1899 3080 1900 3084
rect 1894 3079 1900 3080
rect 2062 3084 2068 3085
rect 2062 3080 2063 3084
rect 2067 3080 2068 3084
rect 2062 3079 2068 3080
rect 2254 3084 2260 3085
rect 2254 3080 2255 3084
rect 2259 3080 2260 3084
rect 2254 3079 2260 3080
rect 2446 3084 2452 3085
rect 2446 3080 2447 3084
rect 2451 3080 2452 3084
rect 2446 3079 2452 3080
rect 2638 3084 2644 3085
rect 2638 3080 2639 3084
rect 2643 3080 2644 3084
rect 2638 3079 2644 3080
rect 2822 3084 2828 3085
rect 2822 3080 2823 3084
rect 2827 3080 2828 3084
rect 2822 3079 2828 3080
rect 3006 3084 3012 3085
rect 3006 3080 3007 3084
rect 3011 3080 3012 3084
rect 3006 3079 3012 3080
rect 3190 3084 3196 3085
rect 3190 3080 3191 3084
rect 3195 3080 3196 3084
rect 3190 3079 3196 3080
rect 3382 3084 3388 3085
rect 3382 3080 3383 3084
rect 3387 3080 3388 3084
rect 3590 3083 3591 3087
rect 3595 3083 3596 3087
rect 3590 3082 3596 3083
rect 3382 3079 3388 3080
rect 134 3052 140 3053
rect 110 3049 116 3050
rect 110 3045 111 3049
rect 115 3045 116 3049
rect 134 3048 135 3052
rect 139 3048 140 3052
rect 134 3047 140 3048
rect 222 3052 228 3053
rect 222 3048 223 3052
rect 227 3048 228 3052
rect 222 3047 228 3048
rect 326 3052 332 3053
rect 326 3048 327 3052
rect 331 3048 332 3052
rect 326 3047 332 3048
rect 438 3052 444 3053
rect 438 3048 439 3052
rect 443 3048 444 3052
rect 438 3047 444 3048
rect 550 3052 556 3053
rect 550 3048 551 3052
rect 555 3048 556 3052
rect 550 3047 556 3048
rect 662 3052 668 3053
rect 662 3048 663 3052
rect 667 3048 668 3052
rect 662 3047 668 3048
rect 1830 3049 1836 3050
rect 110 3044 116 3045
rect 1830 3045 1831 3049
rect 1835 3045 1836 3049
rect 1830 3044 1836 3045
rect 110 3032 116 3033
rect 110 3028 111 3032
rect 115 3028 116 3032
rect 110 3027 116 3028
rect 1830 3032 1836 3033
rect 1830 3028 1831 3032
rect 1835 3028 1836 3032
rect 1830 3027 1836 3028
rect 2198 3028 2204 3029
rect 1870 3025 1876 3026
rect 1870 3021 1871 3025
rect 1875 3021 1876 3025
rect 2198 3024 2199 3028
rect 2203 3024 2204 3028
rect 2198 3023 2204 3024
rect 2334 3028 2340 3029
rect 2334 3024 2335 3028
rect 2339 3024 2340 3028
rect 2334 3023 2340 3024
rect 2478 3028 2484 3029
rect 2478 3024 2479 3028
rect 2483 3024 2484 3028
rect 2478 3023 2484 3024
rect 2622 3028 2628 3029
rect 2622 3024 2623 3028
rect 2627 3024 2628 3028
rect 2622 3023 2628 3024
rect 2766 3028 2772 3029
rect 2766 3024 2767 3028
rect 2771 3024 2772 3028
rect 2766 3023 2772 3024
rect 2902 3028 2908 3029
rect 2902 3024 2903 3028
rect 2907 3024 2908 3028
rect 2902 3023 2908 3024
rect 3038 3028 3044 3029
rect 3038 3024 3039 3028
rect 3043 3024 3044 3028
rect 3038 3023 3044 3024
rect 3182 3028 3188 3029
rect 3182 3024 3183 3028
rect 3187 3024 3188 3028
rect 3182 3023 3188 3024
rect 3326 3028 3332 3029
rect 3326 3024 3327 3028
rect 3331 3024 3332 3028
rect 3326 3023 3332 3024
rect 3590 3025 3596 3026
rect 1870 3020 1876 3021
rect 3590 3021 3591 3025
rect 3595 3021 3596 3025
rect 3590 3020 3596 3021
rect 142 3014 148 3015
rect 142 3010 143 3014
rect 147 3010 148 3014
rect 142 3009 148 3010
rect 230 3014 236 3015
rect 230 3010 231 3014
rect 235 3010 236 3014
rect 230 3009 236 3010
rect 334 3014 340 3015
rect 334 3010 335 3014
rect 339 3010 340 3014
rect 334 3009 340 3010
rect 446 3014 452 3015
rect 446 3010 447 3014
rect 451 3010 452 3014
rect 446 3009 452 3010
rect 558 3014 564 3015
rect 558 3010 559 3014
rect 563 3010 564 3014
rect 558 3009 564 3010
rect 670 3014 676 3015
rect 670 3010 671 3014
rect 675 3010 676 3014
rect 670 3009 676 3010
rect 1870 3008 1876 3009
rect 1870 3004 1871 3008
rect 1875 3004 1876 3008
rect 1870 3003 1876 3004
rect 3590 3008 3596 3009
rect 3590 3004 3591 3008
rect 3595 3004 3596 3008
rect 3590 3003 3596 3004
rect 2206 2990 2212 2991
rect 2206 2986 2207 2990
rect 2211 2986 2212 2990
rect 2206 2985 2212 2986
rect 2342 2990 2348 2991
rect 2342 2986 2343 2990
rect 2347 2986 2348 2990
rect 2342 2985 2348 2986
rect 2486 2990 2492 2991
rect 2486 2986 2487 2990
rect 2491 2986 2492 2990
rect 2486 2985 2492 2986
rect 2630 2990 2636 2991
rect 2630 2986 2631 2990
rect 2635 2986 2636 2990
rect 2630 2985 2636 2986
rect 2774 2990 2780 2991
rect 2774 2986 2775 2990
rect 2779 2986 2780 2990
rect 2774 2985 2780 2986
rect 2910 2990 2916 2991
rect 2910 2986 2911 2990
rect 2915 2986 2916 2990
rect 2910 2985 2916 2986
rect 3046 2990 3052 2991
rect 3046 2986 3047 2990
rect 3051 2986 3052 2990
rect 3046 2985 3052 2986
rect 3190 2990 3196 2991
rect 3190 2986 3191 2990
rect 3195 2986 3196 2990
rect 3190 2985 3196 2986
rect 3334 2990 3340 2991
rect 3334 2986 3335 2990
rect 3339 2986 3340 2990
rect 3334 2985 3340 2986
rect 158 2970 164 2971
rect 158 2966 159 2970
rect 163 2966 164 2970
rect 158 2965 164 2966
rect 318 2970 324 2971
rect 318 2966 319 2970
rect 323 2966 324 2970
rect 318 2965 324 2966
rect 486 2970 492 2971
rect 486 2966 487 2970
rect 491 2966 492 2970
rect 486 2965 492 2966
rect 646 2970 652 2971
rect 646 2966 647 2970
rect 651 2966 652 2970
rect 646 2965 652 2966
rect 798 2970 804 2971
rect 798 2966 799 2970
rect 803 2966 804 2970
rect 798 2965 804 2966
rect 942 2970 948 2971
rect 942 2966 943 2970
rect 947 2966 948 2970
rect 942 2965 948 2966
rect 1078 2970 1084 2971
rect 1078 2966 1079 2970
rect 1083 2966 1084 2970
rect 1078 2965 1084 2966
rect 1198 2970 1204 2971
rect 1198 2966 1199 2970
rect 1203 2966 1204 2970
rect 1198 2965 1204 2966
rect 1310 2970 1316 2971
rect 1310 2966 1311 2970
rect 1315 2966 1316 2970
rect 1310 2965 1316 2966
rect 1422 2970 1428 2971
rect 1422 2966 1423 2970
rect 1427 2966 1428 2970
rect 1422 2965 1428 2966
rect 1534 2970 1540 2971
rect 1534 2966 1535 2970
rect 1539 2966 1540 2970
rect 1534 2965 1540 2966
rect 1646 2970 1652 2971
rect 1646 2966 1647 2970
rect 1651 2966 1652 2970
rect 1646 2965 1652 2966
rect 110 2952 116 2953
rect 110 2948 111 2952
rect 115 2948 116 2952
rect 110 2947 116 2948
rect 1830 2952 1836 2953
rect 1830 2948 1831 2952
rect 1835 2948 1836 2952
rect 1830 2947 1836 2948
rect 2126 2946 2132 2947
rect 2126 2942 2127 2946
rect 2131 2942 2132 2946
rect 2126 2941 2132 2942
rect 2206 2946 2212 2947
rect 2206 2942 2207 2946
rect 2211 2942 2212 2946
rect 2206 2941 2212 2942
rect 2286 2946 2292 2947
rect 2286 2942 2287 2946
rect 2291 2942 2292 2946
rect 2286 2941 2292 2942
rect 2366 2946 2372 2947
rect 2366 2942 2367 2946
rect 2371 2942 2372 2946
rect 2366 2941 2372 2942
rect 2446 2946 2452 2947
rect 2446 2942 2447 2946
rect 2451 2942 2452 2946
rect 2446 2941 2452 2942
rect 2526 2946 2532 2947
rect 2526 2942 2527 2946
rect 2531 2942 2532 2946
rect 2526 2941 2532 2942
rect 2606 2946 2612 2947
rect 2606 2942 2607 2946
rect 2611 2942 2612 2946
rect 2606 2941 2612 2942
rect 2694 2946 2700 2947
rect 2694 2942 2695 2946
rect 2699 2942 2700 2946
rect 2694 2941 2700 2942
rect 2790 2946 2796 2947
rect 2790 2942 2791 2946
rect 2795 2942 2796 2946
rect 2790 2941 2796 2942
rect 2910 2946 2916 2947
rect 2910 2942 2911 2946
rect 2915 2942 2916 2946
rect 2910 2941 2916 2942
rect 3038 2946 3044 2947
rect 3038 2942 3039 2946
rect 3043 2942 3044 2946
rect 3038 2941 3044 2942
rect 3182 2946 3188 2947
rect 3182 2942 3183 2946
rect 3187 2942 3188 2946
rect 3182 2941 3188 2942
rect 3334 2946 3340 2947
rect 3334 2942 3335 2946
rect 3339 2942 3340 2946
rect 3334 2941 3340 2942
rect 3494 2946 3500 2947
rect 3494 2942 3495 2946
rect 3499 2942 3500 2946
rect 3494 2941 3500 2942
rect 110 2935 116 2936
rect 110 2931 111 2935
rect 115 2931 116 2935
rect 1830 2935 1836 2936
rect 110 2930 116 2931
rect 150 2932 156 2933
rect 150 2928 151 2932
rect 155 2928 156 2932
rect 150 2927 156 2928
rect 310 2932 316 2933
rect 310 2928 311 2932
rect 315 2928 316 2932
rect 310 2927 316 2928
rect 478 2932 484 2933
rect 478 2928 479 2932
rect 483 2928 484 2932
rect 478 2927 484 2928
rect 638 2932 644 2933
rect 638 2928 639 2932
rect 643 2928 644 2932
rect 638 2927 644 2928
rect 790 2932 796 2933
rect 790 2928 791 2932
rect 795 2928 796 2932
rect 790 2927 796 2928
rect 934 2932 940 2933
rect 934 2928 935 2932
rect 939 2928 940 2932
rect 934 2927 940 2928
rect 1070 2932 1076 2933
rect 1070 2928 1071 2932
rect 1075 2928 1076 2932
rect 1070 2927 1076 2928
rect 1190 2932 1196 2933
rect 1190 2928 1191 2932
rect 1195 2928 1196 2932
rect 1190 2927 1196 2928
rect 1302 2932 1308 2933
rect 1302 2928 1303 2932
rect 1307 2928 1308 2932
rect 1302 2927 1308 2928
rect 1414 2932 1420 2933
rect 1414 2928 1415 2932
rect 1419 2928 1420 2932
rect 1414 2927 1420 2928
rect 1526 2932 1532 2933
rect 1526 2928 1527 2932
rect 1531 2928 1532 2932
rect 1526 2927 1532 2928
rect 1638 2932 1644 2933
rect 1638 2928 1639 2932
rect 1643 2928 1644 2932
rect 1830 2931 1831 2935
rect 1835 2931 1836 2935
rect 1830 2930 1836 2931
rect 1638 2927 1644 2928
rect 1870 2928 1876 2929
rect 1870 2924 1871 2928
rect 1875 2924 1876 2928
rect 1870 2923 1876 2924
rect 3590 2928 3596 2929
rect 3590 2924 3591 2928
rect 3595 2924 3596 2928
rect 3590 2923 3596 2924
rect 1870 2911 1876 2912
rect 1870 2907 1871 2911
rect 1875 2907 1876 2911
rect 3590 2911 3596 2912
rect 1870 2906 1876 2907
rect 2118 2908 2124 2909
rect 2118 2904 2119 2908
rect 2123 2904 2124 2908
rect 2118 2903 2124 2904
rect 2198 2908 2204 2909
rect 2198 2904 2199 2908
rect 2203 2904 2204 2908
rect 2198 2903 2204 2904
rect 2278 2908 2284 2909
rect 2278 2904 2279 2908
rect 2283 2904 2284 2908
rect 2278 2903 2284 2904
rect 2358 2908 2364 2909
rect 2358 2904 2359 2908
rect 2363 2904 2364 2908
rect 2358 2903 2364 2904
rect 2438 2908 2444 2909
rect 2438 2904 2439 2908
rect 2443 2904 2444 2908
rect 2438 2903 2444 2904
rect 2518 2908 2524 2909
rect 2518 2904 2519 2908
rect 2523 2904 2524 2908
rect 2518 2903 2524 2904
rect 2598 2908 2604 2909
rect 2598 2904 2599 2908
rect 2603 2904 2604 2908
rect 2598 2903 2604 2904
rect 2686 2908 2692 2909
rect 2686 2904 2687 2908
rect 2691 2904 2692 2908
rect 2686 2903 2692 2904
rect 2782 2908 2788 2909
rect 2782 2904 2783 2908
rect 2787 2904 2788 2908
rect 2782 2903 2788 2904
rect 2902 2908 2908 2909
rect 2902 2904 2903 2908
rect 2907 2904 2908 2908
rect 2902 2903 2908 2904
rect 3030 2908 3036 2909
rect 3030 2904 3031 2908
rect 3035 2904 3036 2908
rect 3030 2903 3036 2904
rect 3174 2908 3180 2909
rect 3174 2904 3175 2908
rect 3179 2904 3180 2908
rect 3174 2903 3180 2904
rect 3326 2908 3332 2909
rect 3326 2904 3327 2908
rect 3331 2904 3332 2908
rect 3326 2903 3332 2904
rect 3486 2908 3492 2909
rect 3486 2904 3487 2908
rect 3491 2904 3492 2908
rect 3590 2907 3591 2911
rect 3595 2907 3596 2911
rect 3590 2906 3596 2907
rect 3486 2903 3492 2904
rect 150 2888 156 2889
rect 110 2885 116 2886
rect 110 2881 111 2885
rect 115 2881 116 2885
rect 150 2884 151 2888
rect 155 2884 156 2888
rect 150 2883 156 2884
rect 310 2888 316 2889
rect 310 2884 311 2888
rect 315 2884 316 2888
rect 310 2883 316 2884
rect 470 2888 476 2889
rect 470 2884 471 2888
rect 475 2884 476 2888
rect 470 2883 476 2884
rect 630 2888 636 2889
rect 630 2884 631 2888
rect 635 2884 636 2888
rect 630 2883 636 2884
rect 782 2888 788 2889
rect 782 2884 783 2888
rect 787 2884 788 2888
rect 782 2883 788 2884
rect 926 2888 932 2889
rect 926 2884 927 2888
rect 931 2884 932 2888
rect 926 2883 932 2884
rect 1054 2888 1060 2889
rect 1054 2884 1055 2888
rect 1059 2884 1060 2888
rect 1054 2883 1060 2884
rect 1174 2888 1180 2889
rect 1174 2884 1175 2888
rect 1179 2884 1180 2888
rect 1174 2883 1180 2884
rect 1286 2888 1292 2889
rect 1286 2884 1287 2888
rect 1291 2884 1292 2888
rect 1286 2883 1292 2884
rect 1390 2888 1396 2889
rect 1390 2884 1391 2888
rect 1395 2884 1396 2888
rect 1390 2883 1396 2884
rect 1486 2888 1492 2889
rect 1486 2884 1487 2888
rect 1491 2884 1492 2888
rect 1486 2883 1492 2884
rect 1590 2888 1596 2889
rect 1590 2884 1591 2888
rect 1595 2884 1596 2888
rect 1590 2883 1596 2884
rect 1694 2888 1700 2889
rect 1694 2884 1695 2888
rect 1699 2884 1700 2888
rect 1694 2883 1700 2884
rect 1830 2885 1836 2886
rect 110 2880 116 2881
rect 1830 2881 1831 2885
rect 1835 2881 1836 2885
rect 1830 2880 1836 2881
rect 110 2868 116 2869
rect 110 2864 111 2868
rect 115 2864 116 2868
rect 110 2863 116 2864
rect 1830 2868 1836 2869
rect 1830 2864 1831 2868
rect 1835 2864 1836 2868
rect 1830 2863 1836 2864
rect 2046 2864 2052 2865
rect 1870 2861 1876 2862
rect 1870 2857 1871 2861
rect 1875 2857 1876 2861
rect 2046 2860 2047 2864
rect 2051 2860 2052 2864
rect 2046 2859 2052 2860
rect 2134 2864 2140 2865
rect 2134 2860 2135 2864
rect 2139 2860 2140 2864
rect 2134 2859 2140 2860
rect 2238 2864 2244 2865
rect 2238 2860 2239 2864
rect 2243 2860 2244 2864
rect 2238 2859 2244 2860
rect 2342 2864 2348 2865
rect 2342 2860 2343 2864
rect 2347 2860 2348 2864
rect 2342 2859 2348 2860
rect 2462 2864 2468 2865
rect 2462 2860 2463 2864
rect 2467 2860 2468 2864
rect 2462 2859 2468 2860
rect 2590 2864 2596 2865
rect 2590 2860 2591 2864
rect 2595 2860 2596 2864
rect 2590 2859 2596 2860
rect 2726 2864 2732 2865
rect 2726 2860 2727 2864
rect 2731 2860 2732 2864
rect 2726 2859 2732 2860
rect 2878 2864 2884 2865
rect 2878 2860 2879 2864
rect 2883 2860 2884 2864
rect 2878 2859 2884 2860
rect 3030 2864 3036 2865
rect 3030 2860 3031 2864
rect 3035 2860 3036 2864
rect 3030 2859 3036 2860
rect 3190 2864 3196 2865
rect 3190 2860 3191 2864
rect 3195 2860 3196 2864
rect 3190 2859 3196 2860
rect 3358 2864 3364 2865
rect 3358 2860 3359 2864
rect 3363 2860 3364 2864
rect 3358 2859 3364 2860
rect 3502 2864 3508 2865
rect 3502 2860 3503 2864
rect 3507 2860 3508 2864
rect 3502 2859 3508 2860
rect 3590 2861 3596 2862
rect 1870 2856 1876 2857
rect 3590 2857 3591 2861
rect 3595 2857 3596 2861
rect 3590 2856 3596 2857
rect 158 2850 164 2851
rect 158 2846 159 2850
rect 163 2846 164 2850
rect 158 2845 164 2846
rect 318 2850 324 2851
rect 318 2846 319 2850
rect 323 2846 324 2850
rect 318 2845 324 2846
rect 478 2850 484 2851
rect 478 2846 479 2850
rect 483 2846 484 2850
rect 478 2845 484 2846
rect 638 2850 644 2851
rect 638 2846 639 2850
rect 643 2846 644 2850
rect 638 2845 644 2846
rect 790 2850 796 2851
rect 790 2846 791 2850
rect 795 2846 796 2850
rect 790 2845 796 2846
rect 934 2850 940 2851
rect 934 2846 935 2850
rect 939 2846 940 2850
rect 934 2845 940 2846
rect 1062 2850 1068 2851
rect 1062 2846 1063 2850
rect 1067 2846 1068 2850
rect 1062 2845 1068 2846
rect 1182 2850 1188 2851
rect 1182 2846 1183 2850
rect 1187 2846 1188 2850
rect 1182 2845 1188 2846
rect 1294 2850 1300 2851
rect 1294 2846 1295 2850
rect 1299 2846 1300 2850
rect 1294 2845 1300 2846
rect 1398 2850 1404 2851
rect 1398 2846 1399 2850
rect 1403 2846 1404 2850
rect 1398 2845 1404 2846
rect 1494 2850 1500 2851
rect 1494 2846 1495 2850
rect 1499 2846 1500 2850
rect 1494 2845 1500 2846
rect 1598 2850 1604 2851
rect 1598 2846 1599 2850
rect 1603 2846 1604 2850
rect 1598 2845 1604 2846
rect 1702 2850 1708 2851
rect 1702 2846 1703 2850
rect 1707 2846 1708 2850
rect 1702 2845 1708 2846
rect 1870 2844 1876 2845
rect 1870 2840 1871 2844
rect 1875 2840 1876 2844
rect 1870 2839 1876 2840
rect 3590 2844 3596 2845
rect 3590 2840 3591 2844
rect 3595 2840 3596 2844
rect 3590 2839 3596 2840
rect 2054 2826 2060 2827
rect 2054 2822 2055 2826
rect 2059 2822 2060 2826
rect 2054 2821 2060 2822
rect 2142 2826 2148 2827
rect 2142 2822 2143 2826
rect 2147 2822 2148 2826
rect 2142 2821 2148 2822
rect 2246 2826 2252 2827
rect 2246 2822 2247 2826
rect 2251 2822 2252 2826
rect 2246 2821 2252 2822
rect 2350 2826 2356 2827
rect 2350 2822 2351 2826
rect 2355 2822 2356 2826
rect 2350 2821 2356 2822
rect 2470 2826 2476 2827
rect 2470 2822 2471 2826
rect 2475 2822 2476 2826
rect 2470 2821 2476 2822
rect 2598 2826 2604 2827
rect 2598 2822 2599 2826
rect 2603 2822 2604 2826
rect 2598 2821 2604 2822
rect 2734 2826 2740 2827
rect 2734 2822 2735 2826
rect 2739 2822 2740 2826
rect 2734 2821 2740 2822
rect 2886 2826 2892 2827
rect 2886 2822 2887 2826
rect 2891 2822 2892 2826
rect 2886 2821 2892 2822
rect 3038 2826 3044 2827
rect 3038 2822 3039 2826
rect 3043 2822 3044 2826
rect 3038 2821 3044 2822
rect 3198 2826 3204 2827
rect 3198 2822 3199 2826
rect 3203 2822 3204 2826
rect 3198 2821 3204 2822
rect 3366 2826 3372 2827
rect 3366 2822 3367 2826
rect 3371 2822 3372 2826
rect 3366 2821 3372 2822
rect 3510 2826 3516 2827
rect 3510 2822 3511 2826
rect 3515 2822 3516 2826
rect 3510 2821 3516 2822
rect 142 2814 148 2815
rect 142 2810 143 2814
rect 147 2810 148 2814
rect 142 2809 148 2810
rect 246 2814 252 2815
rect 246 2810 247 2814
rect 251 2810 252 2814
rect 246 2809 252 2810
rect 382 2814 388 2815
rect 382 2810 383 2814
rect 387 2810 388 2814
rect 382 2809 388 2810
rect 534 2814 540 2815
rect 534 2810 535 2814
rect 539 2810 540 2814
rect 534 2809 540 2810
rect 686 2814 692 2815
rect 686 2810 687 2814
rect 691 2810 692 2814
rect 686 2809 692 2810
rect 846 2814 852 2815
rect 846 2810 847 2814
rect 851 2810 852 2814
rect 846 2809 852 2810
rect 998 2814 1004 2815
rect 998 2810 999 2814
rect 1003 2810 1004 2814
rect 998 2809 1004 2810
rect 1142 2814 1148 2815
rect 1142 2810 1143 2814
rect 1147 2810 1148 2814
rect 1142 2809 1148 2810
rect 1278 2814 1284 2815
rect 1278 2810 1279 2814
rect 1283 2810 1284 2814
rect 1278 2809 1284 2810
rect 1406 2814 1412 2815
rect 1406 2810 1407 2814
rect 1411 2810 1412 2814
rect 1406 2809 1412 2810
rect 1526 2814 1532 2815
rect 1526 2810 1527 2814
rect 1531 2810 1532 2814
rect 1526 2809 1532 2810
rect 1646 2814 1652 2815
rect 1646 2810 1647 2814
rect 1651 2810 1652 2814
rect 1646 2809 1652 2810
rect 1750 2814 1756 2815
rect 1750 2810 1751 2814
rect 1755 2810 1756 2814
rect 1750 2809 1756 2810
rect 110 2796 116 2797
rect 110 2792 111 2796
rect 115 2792 116 2796
rect 110 2791 116 2792
rect 1830 2796 1836 2797
rect 1830 2792 1831 2796
rect 1835 2792 1836 2796
rect 1830 2791 1836 2792
rect 1902 2782 1908 2783
rect 110 2779 116 2780
rect 110 2775 111 2779
rect 115 2775 116 2779
rect 1830 2779 1836 2780
rect 110 2774 116 2775
rect 134 2776 140 2777
rect 134 2772 135 2776
rect 139 2772 140 2776
rect 134 2771 140 2772
rect 238 2776 244 2777
rect 238 2772 239 2776
rect 243 2772 244 2776
rect 238 2771 244 2772
rect 374 2776 380 2777
rect 374 2772 375 2776
rect 379 2772 380 2776
rect 374 2771 380 2772
rect 526 2776 532 2777
rect 526 2772 527 2776
rect 531 2772 532 2776
rect 526 2771 532 2772
rect 678 2776 684 2777
rect 678 2772 679 2776
rect 683 2772 684 2776
rect 678 2771 684 2772
rect 838 2776 844 2777
rect 838 2772 839 2776
rect 843 2772 844 2776
rect 838 2771 844 2772
rect 990 2776 996 2777
rect 990 2772 991 2776
rect 995 2772 996 2776
rect 990 2771 996 2772
rect 1134 2776 1140 2777
rect 1134 2772 1135 2776
rect 1139 2772 1140 2776
rect 1134 2771 1140 2772
rect 1270 2776 1276 2777
rect 1270 2772 1271 2776
rect 1275 2772 1276 2776
rect 1270 2771 1276 2772
rect 1398 2776 1404 2777
rect 1398 2772 1399 2776
rect 1403 2772 1404 2776
rect 1398 2771 1404 2772
rect 1518 2776 1524 2777
rect 1518 2772 1519 2776
rect 1523 2772 1524 2776
rect 1518 2771 1524 2772
rect 1638 2776 1644 2777
rect 1638 2772 1639 2776
rect 1643 2772 1644 2776
rect 1638 2771 1644 2772
rect 1742 2776 1748 2777
rect 1742 2772 1743 2776
rect 1747 2772 1748 2776
rect 1830 2775 1831 2779
rect 1835 2775 1836 2779
rect 1902 2778 1903 2782
rect 1907 2778 1908 2782
rect 1902 2777 1908 2778
rect 2014 2782 2020 2783
rect 2014 2778 2015 2782
rect 2019 2778 2020 2782
rect 2014 2777 2020 2778
rect 2166 2782 2172 2783
rect 2166 2778 2167 2782
rect 2171 2778 2172 2782
rect 2166 2777 2172 2778
rect 2326 2782 2332 2783
rect 2326 2778 2327 2782
rect 2331 2778 2332 2782
rect 2326 2777 2332 2778
rect 2486 2782 2492 2783
rect 2486 2778 2487 2782
rect 2491 2778 2492 2782
rect 2486 2777 2492 2778
rect 2638 2782 2644 2783
rect 2638 2778 2639 2782
rect 2643 2778 2644 2782
rect 2638 2777 2644 2778
rect 2790 2782 2796 2783
rect 2790 2778 2791 2782
rect 2795 2778 2796 2782
rect 2790 2777 2796 2778
rect 2942 2782 2948 2783
rect 2942 2778 2943 2782
rect 2947 2778 2948 2782
rect 2942 2777 2948 2778
rect 3086 2782 3092 2783
rect 3086 2778 3087 2782
rect 3091 2778 3092 2782
rect 3086 2777 3092 2778
rect 3230 2782 3236 2783
rect 3230 2778 3231 2782
rect 3235 2778 3236 2782
rect 3230 2777 3236 2778
rect 3382 2782 3388 2783
rect 3382 2778 3383 2782
rect 3387 2778 3388 2782
rect 3382 2777 3388 2778
rect 3510 2782 3516 2783
rect 3510 2778 3511 2782
rect 3515 2778 3516 2782
rect 3510 2777 3516 2778
rect 1830 2774 1836 2775
rect 1742 2771 1748 2772
rect 1870 2764 1876 2765
rect 1870 2760 1871 2764
rect 1875 2760 1876 2764
rect 1870 2759 1876 2760
rect 3590 2764 3596 2765
rect 3590 2760 3591 2764
rect 3595 2760 3596 2764
rect 3590 2759 3596 2760
rect 1870 2747 1876 2748
rect 1870 2743 1871 2747
rect 1875 2743 1876 2747
rect 3590 2747 3596 2748
rect 1870 2742 1876 2743
rect 1894 2744 1900 2745
rect 1894 2740 1895 2744
rect 1899 2740 1900 2744
rect 1894 2739 1900 2740
rect 2006 2744 2012 2745
rect 2006 2740 2007 2744
rect 2011 2740 2012 2744
rect 2006 2739 2012 2740
rect 2158 2744 2164 2745
rect 2158 2740 2159 2744
rect 2163 2740 2164 2744
rect 2158 2739 2164 2740
rect 2318 2744 2324 2745
rect 2318 2740 2319 2744
rect 2323 2740 2324 2744
rect 2318 2739 2324 2740
rect 2478 2744 2484 2745
rect 2478 2740 2479 2744
rect 2483 2740 2484 2744
rect 2478 2739 2484 2740
rect 2630 2744 2636 2745
rect 2630 2740 2631 2744
rect 2635 2740 2636 2744
rect 2630 2739 2636 2740
rect 2782 2744 2788 2745
rect 2782 2740 2783 2744
rect 2787 2740 2788 2744
rect 2782 2739 2788 2740
rect 2934 2744 2940 2745
rect 2934 2740 2935 2744
rect 2939 2740 2940 2744
rect 2934 2739 2940 2740
rect 3078 2744 3084 2745
rect 3078 2740 3079 2744
rect 3083 2740 3084 2744
rect 3078 2739 3084 2740
rect 3222 2744 3228 2745
rect 3222 2740 3223 2744
rect 3227 2740 3228 2744
rect 3222 2739 3228 2740
rect 3374 2744 3380 2745
rect 3374 2740 3375 2744
rect 3379 2740 3380 2744
rect 3374 2739 3380 2740
rect 3502 2744 3508 2745
rect 3502 2740 3503 2744
rect 3507 2740 3508 2744
rect 3590 2743 3591 2747
rect 3595 2743 3596 2747
rect 3590 2742 3596 2743
rect 3502 2739 3508 2740
rect 134 2728 140 2729
rect 110 2725 116 2726
rect 110 2721 111 2725
rect 115 2721 116 2725
rect 134 2724 135 2728
rect 139 2724 140 2728
rect 134 2723 140 2724
rect 230 2728 236 2729
rect 230 2724 231 2728
rect 235 2724 236 2728
rect 230 2723 236 2724
rect 366 2728 372 2729
rect 366 2724 367 2728
rect 371 2724 372 2728
rect 366 2723 372 2724
rect 510 2728 516 2729
rect 510 2724 511 2728
rect 515 2724 516 2728
rect 510 2723 516 2724
rect 662 2728 668 2729
rect 662 2724 663 2728
rect 667 2724 668 2728
rect 662 2723 668 2724
rect 814 2728 820 2729
rect 814 2724 815 2728
rect 819 2724 820 2728
rect 814 2723 820 2724
rect 974 2728 980 2729
rect 974 2724 975 2728
rect 979 2724 980 2728
rect 974 2723 980 2724
rect 1134 2728 1140 2729
rect 1134 2724 1135 2728
rect 1139 2724 1140 2728
rect 1134 2723 1140 2724
rect 1286 2728 1292 2729
rect 1286 2724 1287 2728
rect 1291 2724 1292 2728
rect 1286 2723 1292 2724
rect 1446 2728 1452 2729
rect 1446 2724 1447 2728
rect 1451 2724 1452 2728
rect 1446 2723 1452 2724
rect 1606 2728 1612 2729
rect 1606 2724 1607 2728
rect 1611 2724 1612 2728
rect 1606 2723 1612 2724
rect 1742 2728 1748 2729
rect 1742 2724 1743 2728
rect 1747 2724 1748 2728
rect 1742 2723 1748 2724
rect 1830 2725 1836 2726
rect 110 2720 116 2721
rect 1830 2721 1831 2725
rect 1835 2721 1836 2725
rect 1830 2720 1836 2721
rect 110 2708 116 2709
rect 110 2704 111 2708
rect 115 2704 116 2708
rect 110 2703 116 2704
rect 1830 2708 1836 2709
rect 1830 2704 1831 2708
rect 1835 2704 1836 2708
rect 1830 2703 1836 2704
rect 1894 2700 1900 2701
rect 1870 2697 1876 2698
rect 1870 2693 1871 2697
rect 1875 2693 1876 2697
rect 1894 2696 1895 2700
rect 1899 2696 1900 2700
rect 1894 2695 1900 2696
rect 2102 2700 2108 2701
rect 2102 2696 2103 2700
rect 2107 2696 2108 2700
rect 2102 2695 2108 2696
rect 2326 2700 2332 2701
rect 2326 2696 2327 2700
rect 2331 2696 2332 2700
rect 2326 2695 2332 2696
rect 2534 2700 2540 2701
rect 2534 2696 2535 2700
rect 2539 2696 2540 2700
rect 2534 2695 2540 2696
rect 2734 2700 2740 2701
rect 2734 2696 2735 2700
rect 2739 2696 2740 2700
rect 2734 2695 2740 2696
rect 2910 2700 2916 2701
rect 2910 2696 2911 2700
rect 2915 2696 2916 2700
rect 2910 2695 2916 2696
rect 3070 2700 3076 2701
rect 3070 2696 3071 2700
rect 3075 2696 3076 2700
rect 3070 2695 3076 2696
rect 3222 2700 3228 2701
rect 3222 2696 3223 2700
rect 3227 2696 3228 2700
rect 3222 2695 3228 2696
rect 3374 2700 3380 2701
rect 3374 2696 3375 2700
rect 3379 2696 3380 2700
rect 3374 2695 3380 2696
rect 3502 2700 3508 2701
rect 3502 2696 3503 2700
rect 3507 2696 3508 2700
rect 3502 2695 3508 2696
rect 3590 2697 3596 2698
rect 1870 2692 1876 2693
rect 3590 2693 3591 2697
rect 3595 2693 3596 2697
rect 3590 2692 3596 2693
rect 142 2690 148 2691
rect 142 2686 143 2690
rect 147 2686 148 2690
rect 142 2685 148 2686
rect 238 2690 244 2691
rect 238 2686 239 2690
rect 243 2686 244 2690
rect 238 2685 244 2686
rect 374 2690 380 2691
rect 374 2686 375 2690
rect 379 2686 380 2690
rect 374 2685 380 2686
rect 518 2690 524 2691
rect 518 2686 519 2690
rect 523 2686 524 2690
rect 518 2685 524 2686
rect 670 2690 676 2691
rect 670 2686 671 2690
rect 675 2686 676 2690
rect 670 2685 676 2686
rect 822 2690 828 2691
rect 822 2686 823 2690
rect 827 2686 828 2690
rect 822 2685 828 2686
rect 982 2690 988 2691
rect 982 2686 983 2690
rect 987 2686 988 2690
rect 982 2685 988 2686
rect 1142 2690 1148 2691
rect 1142 2686 1143 2690
rect 1147 2686 1148 2690
rect 1142 2685 1148 2686
rect 1294 2690 1300 2691
rect 1294 2686 1295 2690
rect 1299 2686 1300 2690
rect 1294 2685 1300 2686
rect 1454 2690 1460 2691
rect 1454 2686 1455 2690
rect 1459 2686 1460 2690
rect 1454 2685 1460 2686
rect 1614 2690 1620 2691
rect 1614 2686 1615 2690
rect 1619 2686 1620 2690
rect 1614 2685 1620 2686
rect 1750 2690 1756 2691
rect 1750 2686 1751 2690
rect 1755 2686 1756 2690
rect 1750 2685 1756 2686
rect 1870 2680 1876 2681
rect 1870 2676 1871 2680
rect 1875 2676 1876 2680
rect 1870 2675 1876 2676
rect 3590 2680 3596 2681
rect 3590 2676 3591 2680
rect 3595 2676 3596 2680
rect 3590 2675 3596 2676
rect 1902 2662 1908 2663
rect 1902 2658 1903 2662
rect 1907 2658 1908 2662
rect 1902 2657 1908 2658
rect 2110 2662 2116 2663
rect 2110 2658 2111 2662
rect 2115 2658 2116 2662
rect 2110 2657 2116 2658
rect 2334 2662 2340 2663
rect 2334 2658 2335 2662
rect 2339 2658 2340 2662
rect 2334 2657 2340 2658
rect 2542 2662 2548 2663
rect 2542 2658 2543 2662
rect 2547 2658 2548 2662
rect 2542 2657 2548 2658
rect 2742 2662 2748 2663
rect 2742 2658 2743 2662
rect 2747 2658 2748 2662
rect 2742 2657 2748 2658
rect 2918 2662 2924 2663
rect 2918 2658 2919 2662
rect 2923 2658 2924 2662
rect 2918 2657 2924 2658
rect 3078 2662 3084 2663
rect 3078 2658 3079 2662
rect 3083 2658 3084 2662
rect 3078 2657 3084 2658
rect 3230 2662 3236 2663
rect 3230 2658 3231 2662
rect 3235 2658 3236 2662
rect 3230 2657 3236 2658
rect 3382 2662 3388 2663
rect 3382 2658 3383 2662
rect 3387 2658 3388 2662
rect 3382 2657 3388 2658
rect 3510 2662 3516 2663
rect 3510 2658 3511 2662
rect 3515 2658 3516 2662
rect 3510 2657 3516 2658
rect 142 2650 148 2651
rect 142 2646 143 2650
rect 147 2646 148 2650
rect 142 2645 148 2646
rect 278 2650 284 2651
rect 278 2646 279 2650
rect 283 2646 284 2650
rect 278 2645 284 2646
rect 446 2650 452 2651
rect 446 2646 447 2650
rect 451 2646 452 2650
rect 446 2645 452 2646
rect 622 2650 628 2651
rect 622 2646 623 2650
rect 627 2646 628 2650
rect 622 2645 628 2646
rect 790 2650 796 2651
rect 790 2646 791 2650
rect 795 2646 796 2650
rect 790 2645 796 2646
rect 950 2650 956 2651
rect 950 2646 951 2650
rect 955 2646 956 2650
rect 950 2645 956 2646
rect 1102 2650 1108 2651
rect 1102 2646 1103 2650
rect 1107 2646 1108 2650
rect 1102 2645 1108 2646
rect 1246 2650 1252 2651
rect 1246 2646 1247 2650
rect 1251 2646 1252 2650
rect 1246 2645 1252 2646
rect 1398 2650 1404 2651
rect 1398 2646 1399 2650
rect 1403 2646 1404 2650
rect 1398 2645 1404 2646
rect 1550 2650 1556 2651
rect 1550 2646 1551 2650
rect 1555 2646 1556 2650
rect 1550 2645 1556 2646
rect 110 2632 116 2633
rect 110 2628 111 2632
rect 115 2628 116 2632
rect 110 2627 116 2628
rect 1830 2632 1836 2633
rect 1830 2628 1831 2632
rect 1835 2628 1836 2632
rect 1830 2627 1836 2628
rect 1902 2622 1908 2623
rect 1902 2618 1903 2622
rect 1907 2618 1908 2622
rect 1902 2617 1908 2618
rect 2054 2622 2060 2623
rect 2054 2618 2055 2622
rect 2059 2618 2060 2622
rect 2054 2617 2060 2618
rect 2262 2622 2268 2623
rect 2262 2618 2263 2622
rect 2267 2618 2268 2622
rect 2262 2617 2268 2618
rect 2494 2622 2500 2623
rect 2494 2618 2495 2622
rect 2499 2618 2500 2622
rect 2494 2617 2500 2618
rect 2750 2622 2756 2623
rect 2750 2618 2751 2622
rect 2755 2618 2756 2622
rect 2750 2617 2756 2618
rect 3014 2622 3020 2623
rect 3014 2618 3015 2622
rect 3019 2618 3020 2622
rect 3014 2617 3020 2618
rect 3286 2622 3292 2623
rect 3286 2618 3287 2622
rect 3291 2618 3292 2622
rect 3286 2617 3292 2618
rect 110 2615 116 2616
rect 110 2611 111 2615
rect 115 2611 116 2615
rect 1830 2615 1836 2616
rect 110 2610 116 2611
rect 134 2612 140 2613
rect 134 2608 135 2612
rect 139 2608 140 2612
rect 134 2607 140 2608
rect 270 2612 276 2613
rect 270 2608 271 2612
rect 275 2608 276 2612
rect 270 2607 276 2608
rect 438 2612 444 2613
rect 438 2608 439 2612
rect 443 2608 444 2612
rect 438 2607 444 2608
rect 614 2612 620 2613
rect 614 2608 615 2612
rect 619 2608 620 2612
rect 614 2607 620 2608
rect 782 2612 788 2613
rect 782 2608 783 2612
rect 787 2608 788 2612
rect 782 2607 788 2608
rect 942 2612 948 2613
rect 942 2608 943 2612
rect 947 2608 948 2612
rect 942 2607 948 2608
rect 1094 2612 1100 2613
rect 1094 2608 1095 2612
rect 1099 2608 1100 2612
rect 1094 2607 1100 2608
rect 1238 2612 1244 2613
rect 1238 2608 1239 2612
rect 1243 2608 1244 2612
rect 1238 2607 1244 2608
rect 1390 2612 1396 2613
rect 1390 2608 1391 2612
rect 1395 2608 1396 2612
rect 1390 2607 1396 2608
rect 1542 2612 1548 2613
rect 1542 2608 1543 2612
rect 1547 2608 1548 2612
rect 1830 2611 1831 2615
rect 1835 2611 1836 2615
rect 1830 2610 1836 2611
rect 1542 2607 1548 2608
rect 1870 2604 1876 2605
rect 1870 2600 1871 2604
rect 1875 2600 1876 2604
rect 1870 2599 1876 2600
rect 3590 2604 3596 2605
rect 3590 2600 3591 2604
rect 3595 2600 3596 2604
rect 3590 2599 3596 2600
rect 1870 2587 1876 2588
rect 1870 2583 1871 2587
rect 1875 2583 1876 2587
rect 3590 2587 3596 2588
rect 1870 2582 1876 2583
rect 1894 2584 1900 2585
rect 1894 2580 1895 2584
rect 1899 2580 1900 2584
rect 1894 2579 1900 2580
rect 2046 2584 2052 2585
rect 2046 2580 2047 2584
rect 2051 2580 2052 2584
rect 2046 2579 2052 2580
rect 2254 2584 2260 2585
rect 2254 2580 2255 2584
rect 2259 2580 2260 2584
rect 2254 2579 2260 2580
rect 2486 2584 2492 2585
rect 2486 2580 2487 2584
rect 2491 2580 2492 2584
rect 2486 2579 2492 2580
rect 2742 2584 2748 2585
rect 2742 2580 2743 2584
rect 2747 2580 2748 2584
rect 2742 2579 2748 2580
rect 3006 2584 3012 2585
rect 3006 2580 3007 2584
rect 3011 2580 3012 2584
rect 3006 2579 3012 2580
rect 3278 2584 3284 2585
rect 3278 2580 3279 2584
rect 3283 2580 3284 2584
rect 3590 2583 3591 2587
rect 3595 2583 3596 2587
rect 3590 2582 3596 2583
rect 3278 2579 3284 2580
rect 134 2564 140 2565
rect 110 2561 116 2562
rect 110 2557 111 2561
rect 115 2557 116 2561
rect 134 2560 135 2564
rect 139 2560 140 2564
rect 134 2559 140 2560
rect 222 2564 228 2565
rect 222 2560 223 2564
rect 227 2560 228 2564
rect 222 2559 228 2560
rect 366 2564 372 2565
rect 366 2560 367 2564
rect 371 2560 372 2564
rect 366 2559 372 2560
rect 526 2564 532 2565
rect 526 2560 527 2564
rect 531 2560 532 2564
rect 526 2559 532 2560
rect 702 2564 708 2565
rect 702 2560 703 2564
rect 707 2560 708 2564
rect 702 2559 708 2560
rect 878 2564 884 2565
rect 878 2560 879 2564
rect 883 2560 884 2564
rect 878 2559 884 2560
rect 1046 2564 1052 2565
rect 1046 2560 1047 2564
rect 1051 2560 1052 2564
rect 1046 2559 1052 2560
rect 1206 2564 1212 2565
rect 1206 2560 1207 2564
rect 1211 2560 1212 2564
rect 1206 2559 1212 2560
rect 1358 2564 1364 2565
rect 1358 2560 1359 2564
rect 1363 2560 1364 2564
rect 1358 2559 1364 2560
rect 1510 2564 1516 2565
rect 1510 2560 1511 2564
rect 1515 2560 1516 2564
rect 1510 2559 1516 2560
rect 1670 2564 1676 2565
rect 1670 2560 1671 2564
rect 1675 2560 1676 2564
rect 1670 2559 1676 2560
rect 1830 2561 1836 2562
rect 110 2556 116 2557
rect 1830 2557 1831 2561
rect 1835 2557 1836 2561
rect 1830 2556 1836 2557
rect 110 2544 116 2545
rect 110 2540 111 2544
rect 115 2540 116 2544
rect 110 2539 116 2540
rect 1830 2544 1836 2545
rect 1830 2540 1831 2544
rect 1835 2540 1836 2544
rect 1830 2539 1836 2540
rect 1894 2540 1900 2541
rect 1870 2537 1876 2538
rect 1870 2533 1871 2537
rect 1875 2533 1876 2537
rect 1894 2536 1895 2540
rect 1899 2536 1900 2540
rect 1894 2535 1900 2536
rect 2006 2540 2012 2541
rect 2006 2536 2007 2540
rect 2011 2536 2012 2540
rect 2006 2535 2012 2536
rect 2158 2540 2164 2541
rect 2158 2536 2159 2540
rect 2163 2536 2164 2540
rect 2158 2535 2164 2536
rect 2318 2540 2324 2541
rect 2318 2536 2319 2540
rect 2323 2536 2324 2540
rect 2318 2535 2324 2536
rect 2470 2540 2476 2541
rect 2470 2536 2471 2540
rect 2475 2536 2476 2540
rect 2470 2535 2476 2536
rect 2622 2540 2628 2541
rect 2622 2536 2623 2540
rect 2627 2536 2628 2540
rect 2622 2535 2628 2536
rect 2758 2540 2764 2541
rect 2758 2536 2759 2540
rect 2763 2536 2764 2540
rect 2758 2535 2764 2536
rect 2886 2540 2892 2541
rect 2886 2536 2887 2540
rect 2891 2536 2892 2540
rect 2886 2535 2892 2536
rect 3006 2540 3012 2541
rect 3006 2536 3007 2540
rect 3011 2536 3012 2540
rect 3006 2535 3012 2536
rect 3118 2540 3124 2541
rect 3118 2536 3119 2540
rect 3123 2536 3124 2540
rect 3118 2535 3124 2536
rect 3222 2540 3228 2541
rect 3222 2536 3223 2540
rect 3227 2536 3228 2540
rect 3222 2535 3228 2536
rect 3318 2540 3324 2541
rect 3318 2536 3319 2540
rect 3323 2536 3324 2540
rect 3318 2535 3324 2536
rect 3422 2540 3428 2541
rect 3422 2536 3423 2540
rect 3427 2536 3428 2540
rect 3422 2535 3428 2536
rect 3502 2540 3508 2541
rect 3502 2536 3503 2540
rect 3507 2536 3508 2540
rect 3502 2535 3508 2536
rect 3590 2537 3596 2538
rect 1870 2532 1876 2533
rect 3590 2533 3591 2537
rect 3595 2533 3596 2537
rect 3590 2532 3596 2533
rect 142 2526 148 2527
rect 142 2522 143 2526
rect 147 2522 148 2526
rect 142 2521 148 2522
rect 230 2526 236 2527
rect 230 2522 231 2526
rect 235 2522 236 2526
rect 230 2521 236 2522
rect 374 2526 380 2527
rect 374 2522 375 2526
rect 379 2522 380 2526
rect 374 2521 380 2522
rect 534 2526 540 2527
rect 534 2522 535 2526
rect 539 2522 540 2526
rect 534 2521 540 2522
rect 710 2526 716 2527
rect 710 2522 711 2526
rect 715 2522 716 2526
rect 710 2521 716 2522
rect 886 2526 892 2527
rect 886 2522 887 2526
rect 891 2522 892 2526
rect 886 2521 892 2522
rect 1054 2526 1060 2527
rect 1054 2522 1055 2526
rect 1059 2522 1060 2526
rect 1054 2521 1060 2522
rect 1214 2526 1220 2527
rect 1214 2522 1215 2526
rect 1219 2522 1220 2526
rect 1214 2521 1220 2522
rect 1366 2526 1372 2527
rect 1366 2522 1367 2526
rect 1371 2522 1372 2526
rect 1366 2521 1372 2522
rect 1518 2526 1524 2527
rect 1518 2522 1519 2526
rect 1523 2522 1524 2526
rect 1518 2521 1524 2522
rect 1678 2526 1684 2527
rect 1678 2522 1679 2526
rect 1683 2522 1684 2526
rect 1678 2521 1684 2522
rect 1870 2520 1876 2521
rect 1870 2516 1871 2520
rect 1875 2516 1876 2520
rect 1870 2515 1876 2516
rect 3590 2520 3596 2521
rect 3590 2516 3591 2520
rect 3595 2516 3596 2520
rect 3590 2515 3596 2516
rect 1902 2502 1908 2503
rect 1902 2498 1903 2502
rect 1907 2498 1908 2502
rect 1902 2497 1908 2498
rect 2014 2502 2020 2503
rect 2014 2498 2015 2502
rect 2019 2498 2020 2502
rect 2014 2497 2020 2498
rect 2166 2502 2172 2503
rect 2166 2498 2167 2502
rect 2171 2498 2172 2502
rect 2166 2497 2172 2498
rect 2326 2502 2332 2503
rect 2326 2498 2327 2502
rect 2331 2498 2332 2502
rect 2326 2497 2332 2498
rect 2478 2502 2484 2503
rect 2478 2498 2479 2502
rect 2483 2498 2484 2502
rect 2478 2497 2484 2498
rect 2630 2502 2636 2503
rect 2630 2498 2631 2502
rect 2635 2498 2636 2502
rect 2630 2497 2636 2498
rect 2766 2502 2772 2503
rect 2766 2498 2767 2502
rect 2771 2498 2772 2502
rect 2766 2497 2772 2498
rect 2894 2502 2900 2503
rect 2894 2498 2895 2502
rect 2899 2498 2900 2502
rect 2894 2497 2900 2498
rect 3014 2502 3020 2503
rect 3014 2498 3015 2502
rect 3019 2498 3020 2502
rect 3014 2497 3020 2498
rect 3126 2502 3132 2503
rect 3126 2498 3127 2502
rect 3131 2498 3132 2502
rect 3126 2497 3132 2498
rect 3230 2502 3236 2503
rect 3230 2498 3231 2502
rect 3235 2498 3236 2502
rect 3230 2497 3236 2498
rect 3326 2502 3332 2503
rect 3326 2498 3327 2502
rect 3331 2498 3332 2502
rect 3326 2497 3332 2498
rect 3430 2502 3436 2503
rect 3430 2498 3431 2502
rect 3435 2498 3436 2502
rect 3430 2497 3436 2498
rect 3510 2502 3516 2503
rect 3510 2498 3511 2502
rect 3515 2498 3516 2502
rect 3510 2497 3516 2498
rect 142 2490 148 2491
rect 142 2486 143 2490
rect 147 2486 148 2490
rect 142 2485 148 2486
rect 222 2490 228 2491
rect 222 2486 223 2490
rect 227 2486 228 2490
rect 222 2485 228 2486
rect 302 2490 308 2491
rect 302 2486 303 2490
rect 307 2486 308 2490
rect 302 2485 308 2486
rect 390 2490 396 2491
rect 390 2486 391 2490
rect 395 2486 396 2490
rect 390 2485 396 2486
rect 510 2490 516 2491
rect 510 2486 511 2490
rect 515 2486 516 2490
rect 510 2485 516 2486
rect 646 2490 652 2491
rect 646 2486 647 2490
rect 651 2486 652 2490
rect 646 2485 652 2486
rect 782 2490 788 2491
rect 782 2486 783 2490
rect 787 2486 788 2490
rect 782 2485 788 2486
rect 926 2490 932 2491
rect 926 2486 927 2490
rect 931 2486 932 2490
rect 926 2485 932 2486
rect 1062 2490 1068 2491
rect 1062 2486 1063 2490
rect 1067 2486 1068 2490
rect 1062 2485 1068 2486
rect 1190 2490 1196 2491
rect 1190 2486 1191 2490
rect 1195 2486 1196 2490
rect 1190 2485 1196 2486
rect 1310 2490 1316 2491
rect 1310 2486 1311 2490
rect 1315 2486 1316 2490
rect 1310 2485 1316 2486
rect 1430 2490 1436 2491
rect 1430 2486 1431 2490
rect 1435 2486 1436 2490
rect 1430 2485 1436 2486
rect 1550 2490 1556 2491
rect 1550 2486 1551 2490
rect 1555 2486 1556 2490
rect 1550 2485 1556 2486
rect 1670 2490 1676 2491
rect 1670 2486 1671 2490
rect 1675 2486 1676 2490
rect 1670 2485 1676 2486
rect 110 2472 116 2473
rect 110 2468 111 2472
rect 115 2468 116 2472
rect 110 2467 116 2468
rect 1830 2472 1836 2473
rect 1830 2468 1831 2472
rect 1835 2468 1836 2472
rect 1830 2467 1836 2468
rect 1998 2462 2004 2463
rect 1998 2458 1999 2462
rect 2003 2458 2004 2462
rect 1998 2457 2004 2458
rect 2126 2462 2132 2463
rect 2126 2458 2127 2462
rect 2131 2458 2132 2462
rect 2126 2457 2132 2458
rect 2262 2462 2268 2463
rect 2262 2458 2263 2462
rect 2267 2458 2268 2462
rect 2262 2457 2268 2458
rect 2406 2462 2412 2463
rect 2406 2458 2407 2462
rect 2411 2458 2412 2462
rect 2406 2457 2412 2458
rect 2550 2462 2556 2463
rect 2550 2458 2551 2462
rect 2555 2458 2556 2462
rect 2550 2457 2556 2458
rect 2702 2462 2708 2463
rect 2702 2458 2703 2462
rect 2707 2458 2708 2462
rect 2702 2457 2708 2458
rect 2862 2462 2868 2463
rect 2862 2458 2863 2462
rect 2867 2458 2868 2462
rect 2862 2457 2868 2458
rect 3022 2462 3028 2463
rect 3022 2458 3023 2462
rect 3027 2458 3028 2462
rect 3022 2457 3028 2458
rect 3190 2462 3196 2463
rect 3190 2458 3191 2462
rect 3195 2458 3196 2462
rect 3190 2457 3196 2458
rect 3358 2462 3364 2463
rect 3358 2458 3359 2462
rect 3363 2458 3364 2462
rect 3358 2457 3364 2458
rect 3510 2462 3516 2463
rect 3510 2458 3511 2462
rect 3515 2458 3516 2462
rect 3510 2457 3516 2458
rect 110 2455 116 2456
rect 110 2451 111 2455
rect 115 2451 116 2455
rect 1830 2455 1836 2456
rect 110 2450 116 2451
rect 134 2452 140 2453
rect 134 2448 135 2452
rect 139 2448 140 2452
rect 134 2447 140 2448
rect 214 2452 220 2453
rect 214 2448 215 2452
rect 219 2448 220 2452
rect 214 2447 220 2448
rect 294 2452 300 2453
rect 294 2448 295 2452
rect 299 2448 300 2452
rect 294 2447 300 2448
rect 382 2452 388 2453
rect 382 2448 383 2452
rect 387 2448 388 2452
rect 382 2447 388 2448
rect 502 2452 508 2453
rect 502 2448 503 2452
rect 507 2448 508 2452
rect 502 2447 508 2448
rect 638 2452 644 2453
rect 638 2448 639 2452
rect 643 2448 644 2452
rect 638 2447 644 2448
rect 774 2452 780 2453
rect 774 2448 775 2452
rect 779 2448 780 2452
rect 774 2447 780 2448
rect 918 2452 924 2453
rect 918 2448 919 2452
rect 923 2448 924 2452
rect 918 2447 924 2448
rect 1054 2452 1060 2453
rect 1054 2448 1055 2452
rect 1059 2448 1060 2452
rect 1054 2447 1060 2448
rect 1182 2452 1188 2453
rect 1182 2448 1183 2452
rect 1187 2448 1188 2452
rect 1182 2447 1188 2448
rect 1302 2452 1308 2453
rect 1302 2448 1303 2452
rect 1307 2448 1308 2452
rect 1302 2447 1308 2448
rect 1422 2452 1428 2453
rect 1422 2448 1423 2452
rect 1427 2448 1428 2452
rect 1422 2447 1428 2448
rect 1542 2452 1548 2453
rect 1542 2448 1543 2452
rect 1547 2448 1548 2452
rect 1542 2447 1548 2448
rect 1662 2452 1668 2453
rect 1662 2448 1663 2452
rect 1667 2448 1668 2452
rect 1830 2451 1831 2455
rect 1835 2451 1836 2455
rect 1830 2450 1836 2451
rect 1662 2447 1668 2448
rect 1870 2444 1876 2445
rect 1870 2440 1871 2444
rect 1875 2440 1876 2444
rect 1870 2439 1876 2440
rect 3590 2444 3596 2445
rect 3590 2440 3591 2444
rect 3595 2440 3596 2444
rect 3590 2439 3596 2440
rect 1870 2427 1876 2428
rect 1870 2423 1871 2427
rect 1875 2423 1876 2427
rect 3590 2427 3596 2428
rect 1870 2422 1876 2423
rect 1990 2424 1996 2425
rect 1990 2420 1991 2424
rect 1995 2420 1996 2424
rect 1990 2419 1996 2420
rect 2118 2424 2124 2425
rect 2118 2420 2119 2424
rect 2123 2420 2124 2424
rect 2118 2419 2124 2420
rect 2254 2424 2260 2425
rect 2254 2420 2255 2424
rect 2259 2420 2260 2424
rect 2254 2419 2260 2420
rect 2398 2424 2404 2425
rect 2398 2420 2399 2424
rect 2403 2420 2404 2424
rect 2398 2419 2404 2420
rect 2542 2424 2548 2425
rect 2542 2420 2543 2424
rect 2547 2420 2548 2424
rect 2542 2419 2548 2420
rect 2694 2424 2700 2425
rect 2694 2420 2695 2424
rect 2699 2420 2700 2424
rect 2694 2419 2700 2420
rect 2854 2424 2860 2425
rect 2854 2420 2855 2424
rect 2859 2420 2860 2424
rect 2854 2419 2860 2420
rect 3014 2424 3020 2425
rect 3014 2420 3015 2424
rect 3019 2420 3020 2424
rect 3014 2419 3020 2420
rect 3182 2424 3188 2425
rect 3182 2420 3183 2424
rect 3187 2420 3188 2424
rect 3182 2419 3188 2420
rect 3350 2424 3356 2425
rect 3350 2420 3351 2424
rect 3355 2420 3356 2424
rect 3350 2419 3356 2420
rect 3502 2424 3508 2425
rect 3502 2420 3503 2424
rect 3507 2420 3508 2424
rect 3590 2423 3591 2427
rect 3595 2423 3596 2427
rect 3590 2422 3596 2423
rect 3502 2419 3508 2420
rect 1062 2396 1068 2397
rect 110 2393 116 2394
rect 110 2389 111 2393
rect 115 2389 116 2393
rect 1062 2392 1063 2396
rect 1067 2392 1068 2396
rect 1062 2391 1068 2392
rect 1142 2396 1148 2397
rect 1142 2392 1143 2396
rect 1147 2392 1148 2396
rect 1142 2391 1148 2392
rect 1222 2396 1228 2397
rect 1222 2392 1223 2396
rect 1227 2392 1228 2396
rect 1222 2391 1228 2392
rect 1302 2396 1308 2397
rect 1302 2392 1303 2396
rect 1307 2392 1308 2396
rect 1302 2391 1308 2392
rect 1382 2396 1388 2397
rect 1382 2392 1383 2396
rect 1387 2392 1388 2396
rect 1382 2391 1388 2392
rect 1462 2396 1468 2397
rect 1462 2392 1463 2396
rect 1467 2392 1468 2396
rect 1462 2391 1468 2392
rect 1830 2393 1836 2394
rect 110 2388 116 2389
rect 1830 2389 1831 2393
rect 1835 2389 1836 2393
rect 1830 2388 1836 2389
rect 110 2376 116 2377
rect 110 2372 111 2376
rect 115 2372 116 2376
rect 110 2371 116 2372
rect 1830 2376 1836 2377
rect 1830 2372 1831 2376
rect 1835 2372 1836 2376
rect 2142 2376 2148 2377
rect 1830 2371 1836 2372
rect 1870 2373 1876 2374
rect 1870 2369 1871 2373
rect 1875 2369 1876 2373
rect 2142 2372 2143 2376
rect 2147 2372 2148 2376
rect 2142 2371 2148 2372
rect 2238 2376 2244 2377
rect 2238 2372 2239 2376
rect 2243 2372 2244 2376
rect 2238 2371 2244 2372
rect 2342 2376 2348 2377
rect 2342 2372 2343 2376
rect 2347 2372 2348 2376
rect 2342 2371 2348 2372
rect 2454 2376 2460 2377
rect 2454 2372 2455 2376
rect 2459 2372 2460 2376
rect 2454 2371 2460 2372
rect 2574 2376 2580 2377
rect 2574 2372 2575 2376
rect 2579 2372 2580 2376
rect 2574 2371 2580 2372
rect 2702 2376 2708 2377
rect 2702 2372 2703 2376
rect 2707 2372 2708 2376
rect 2702 2371 2708 2372
rect 2846 2376 2852 2377
rect 2846 2372 2847 2376
rect 2851 2372 2852 2376
rect 2846 2371 2852 2372
rect 3006 2376 3012 2377
rect 3006 2372 3007 2376
rect 3011 2372 3012 2376
rect 3006 2371 3012 2372
rect 3174 2376 3180 2377
rect 3174 2372 3175 2376
rect 3179 2372 3180 2376
rect 3174 2371 3180 2372
rect 3350 2376 3356 2377
rect 3350 2372 3351 2376
rect 3355 2372 3356 2376
rect 3350 2371 3356 2372
rect 3502 2376 3508 2377
rect 3502 2372 3503 2376
rect 3507 2372 3508 2376
rect 3502 2371 3508 2372
rect 3590 2373 3596 2374
rect 1870 2368 1876 2369
rect 3590 2369 3591 2373
rect 3595 2369 3596 2373
rect 3590 2368 3596 2369
rect 1070 2358 1076 2359
rect 1070 2354 1071 2358
rect 1075 2354 1076 2358
rect 1070 2353 1076 2354
rect 1150 2358 1156 2359
rect 1150 2354 1151 2358
rect 1155 2354 1156 2358
rect 1150 2353 1156 2354
rect 1230 2358 1236 2359
rect 1230 2354 1231 2358
rect 1235 2354 1236 2358
rect 1230 2353 1236 2354
rect 1310 2358 1316 2359
rect 1310 2354 1311 2358
rect 1315 2354 1316 2358
rect 1310 2353 1316 2354
rect 1390 2358 1396 2359
rect 1390 2354 1391 2358
rect 1395 2354 1396 2358
rect 1390 2353 1396 2354
rect 1470 2358 1476 2359
rect 1470 2354 1471 2358
rect 1475 2354 1476 2358
rect 1470 2353 1476 2354
rect 1870 2356 1876 2357
rect 1870 2352 1871 2356
rect 1875 2352 1876 2356
rect 1870 2351 1876 2352
rect 3590 2356 3596 2357
rect 3590 2352 3591 2356
rect 3595 2352 3596 2356
rect 3590 2351 3596 2352
rect 2150 2338 2156 2339
rect 2150 2334 2151 2338
rect 2155 2334 2156 2338
rect 2150 2333 2156 2334
rect 2246 2338 2252 2339
rect 2246 2334 2247 2338
rect 2251 2334 2252 2338
rect 2246 2333 2252 2334
rect 2350 2338 2356 2339
rect 2350 2334 2351 2338
rect 2355 2334 2356 2338
rect 2350 2333 2356 2334
rect 2462 2338 2468 2339
rect 2462 2334 2463 2338
rect 2467 2334 2468 2338
rect 2462 2333 2468 2334
rect 2582 2338 2588 2339
rect 2582 2334 2583 2338
rect 2587 2334 2588 2338
rect 2582 2333 2588 2334
rect 2710 2338 2716 2339
rect 2710 2334 2711 2338
rect 2715 2334 2716 2338
rect 2710 2333 2716 2334
rect 2854 2338 2860 2339
rect 2854 2334 2855 2338
rect 2859 2334 2860 2338
rect 2854 2333 2860 2334
rect 3014 2338 3020 2339
rect 3014 2334 3015 2338
rect 3019 2334 3020 2338
rect 3014 2333 3020 2334
rect 3182 2338 3188 2339
rect 3182 2334 3183 2338
rect 3187 2334 3188 2338
rect 3182 2333 3188 2334
rect 3358 2338 3364 2339
rect 3358 2334 3359 2338
rect 3363 2334 3364 2338
rect 3358 2333 3364 2334
rect 3510 2338 3516 2339
rect 3510 2334 3511 2338
rect 3515 2334 3516 2338
rect 3510 2333 3516 2334
rect 358 2318 364 2319
rect 358 2314 359 2318
rect 363 2314 364 2318
rect 358 2313 364 2314
rect 438 2318 444 2319
rect 438 2314 439 2318
rect 443 2314 444 2318
rect 438 2313 444 2314
rect 518 2318 524 2319
rect 518 2314 519 2318
rect 523 2314 524 2318
rect 518 2313 524 2314
rect 598 2318 604 2319
rect 598 2314 599 2318
rect 603 2314 604 2318
rect 598 2313 604 2314
rect 678 2318 684 2319
rect 678 2314 679 2318
rect 683 2314 684 2318
rect 678 2313 684 2314
rect 758 2318 764 2319
rect 758 2314 759 2318
rect 763 2314 764 2318
rect 758 2313 764 2314
rect 838 2318 844 2319
rect 838 2314 839 2318
rect 843 2314 844 2318
rect 838 2313 844 2314
rect 918 2318 924 2319
rect 918 2314 919 2318
rect 923 2314 924 2318
rect 918 2313 924 2314
rect 998 2318 1004 2319
rect 998 2314 999 2318
rect 1003 2314 1004 2318
rect 998 2313 1004 2314
rect 1078 2318 1084 2319
rect 1078 2314 1079 2318
rect 1083 2314 1084 2318
rect 1078 2313 1084 2314
rect 1158 2318 1164 2319
rect 1158 2314 1159 2318
rect 1163 2314 1164 2318
rect 1158 2313 1164 2314
rect 1238 2318 1244 2319
rect 1238 2314 1239 2318
rect 1243 2314 1244 2318
rect 1238 2313 1244 2314
rect 1318 2318 1324 2319
rect 1318 2314 1319 2318
rect 1323 2314 1324 2318
rect 1318 2313 1324 2314
rect 2278 2302 2284 2303
rect 110 2300 116 2301
rect 110 2296 111 2300
rect 115 2296 116 2300
rect 110 2295 116 2296
rect 1830 2300 1836 2301
rect 1830 2296 1831 2300
rect 1835 2296 1836 2300
rect 2278 2298 2279 2302
rect 2283 2298 2284 2302
rect 2278 2297 2284 2298
rect 2358 2302 2364 2303
rect 2358 2298 2359 2302
rect 2363 2298 2364 2302
rect 2358 2297 2364 2298
rect 2438 2302 2444 2303
rect 2438 2298 2439 2302
rect 2443 2298 2444 2302
rect 2438 2297 2444 2298
rect 2518 2302 2524 2303
rect 2518 2298 2519 2302
rect 2523 2298 2524 2302
rect 2518 2297 2524 2298
rect 2598 2302 2604 2303
rect 2598 2298 2599 2302
rect 2603 2298 2604 2302
rect 2598 2297 2604 2298
rect 2678 2302 2684 2303
rect 2678 2298 2679 2302
rect 2683 2298 2684 2302
rect 2678 2297 2684 2298
rect 2758 2302 2764 2303
rect 2758 2298 2759 2302
rect 2763 2298 2764 2302
rect 2758 2297 2764 2298
rect 2846 2302 2852 2303
rect 2846 2298 2847 2302
rect 2851 2298 2852 2302
rect 2846 2297 2852 2298
rect 2934 2302 2940 2303
rect 2934 2298 2935 2302
rect 2939 2298 2940 2302
rect 2934 2297 2940 2298
rect 1830 2295 1836 2296
rect 1870 2284 1876 2285
rect 110 2283 116 2284
rect 110 2279 111 2283
rect 115 2279 116 2283
rect 1830 2283 1836 2284
rect 110 2278 116 2279
rect 350 2280 356 2281
rect 350 2276 351 2280
rect 355 2276 356 2280
rect 350 2275 356 2276
rect 430 2280 436 2281
rect 430 2276 431 2280
rect 435 2276 436 2280
rect 430 2275 436 2276
rect 510 2280 516 2281
rect 510 2276 511 2280
rect 515 2276 516 2280
rect 510 2275 516 2276
rect 590 2280 596 2281
rect 590 2276 591 2280
rect 595 2276 596 2280
rect 590 2275 596 2276
rect 670 2280 676 2281
rect 670 2276 671 2280
rect 675 2276 676 2280
rect 670 2275 676 2276
rect 750 2280 756 2281
rect 750 2276 751 2280
rect 755 2276 756 2280
rect 750 2275 756 2276
rect 830 2280 836 2281
rect 830 2276 831 2280
rect 835 2276 836 2280
rect 830 2275 836 2276
rect 910 2280 916 2281
rect 910 2276 911 2280
rect 915 2276 916 2280
rect 910 2275 916 2276
rect 990 2280 996 2281
rect 990 2276 991 2280
rect 995 2276 996 2280
rect 990 2275 996 2276
rect 1070 2280 1076 2281
rect 1070 2276 1071 2280
rect 1075 2276 1076 2280
rect 1070 2275 1076 2276
rect 1150 2280 1156 2281
rect 1150 2276 1151 2280
rect 1155 2276 1156 2280
rect 1150 2275 1156 2276
rect 1230 2280 1236 2281
rect 1230 2276 1231 2280
rect 1235 2276 1236 2280
rect 1230 2275 1236 2276
rect 1310 2280 1316 2281
rect 1310 2276 1311 2280
rect 1315 2276 1316 2280
rect 1830 2279 1831 2283
rect 1835 2279 1836 2283
rect 1870 2280 1871 2284
rect 1875 2280 1876 2284
rect 1870 2279 1876 2280
rect 3590 2284 3596 2285
rect 3590 2280 3591 2284
rect 3595 2280 3596 2284
rect 3590 2279 3596 2280
rect 1830 2278 1836 2279
rect 1310 2275 1316 2276
rect 1870 2267 1876 2268
rect 1870 2263 1871 2267
rect 1875 2263 1876 2267
rect 3590 2267 3596 2268
rect 1870 2262 1876 2263
rect 2270 2264 2276 2265
rect 2270 2260 2271 2264
rect 2275 2260 2276 2264
rect 2270 2259 2276 2260
rect 2350 2264 2356 2265
rect 2350 2260 2351 2264
rect 2355 2260 2356 2264
rect 2350 2259 2356 2260
rect 2430 2264 2436 2265
rect 2430 2260 2431 2264
rect 2435 2260 2436 2264
rect 2430 2259 2436 2260
rect 2510 2264 2516 2265
rect 2510 2260 2511 2264
rect 2515 2260 2516 2264
rect 2510 2259 2516 2260
rect 2590 2264 2596 2265
rect 2590 2260 2591 2264
rect 2595 2260 2596 2264
rect 2590 2259 2596 2260
rect 2670 2264 2676 2265
rect 2670 2260 2671 2264
rect 2675 2260 2676 2264
rect 2670 2259 2676 2260
rect 2750 2264 2756 2265
rect 2750 2260 2751 2264
rect 2755 2260 2756 2264
rect 2750 2259 2756 2260
rect 2838 2264 2844 2265
rect 2838 2260 2839 2264
rect 2843 2260 2844 2264
rect 2838 2259 2844 2260
rect 2926 2264 2932 2265
rect 2926 2260 2927 2264
rect 2931 2260 2932 2264
rect 3590 2263 3591 2267
rect 3595 2263 3596 2267
rect 3590 2262 3596 2263
rect 2926 2259 2932 2260
rect 374 2236 380 2237
rect 110 2233 116 2234
rect 110 2229 111 2233
rect 115 2229 116 2233
rect 374 2232 375 2236
rect 379 2232 380 2236
rect 374 2231 380 2232
rect 454 2236 460 2237
rect 454 2232 455 2236
rect 459 2232 460 2236
rect 454 2231 460 2232
rect 534 2236 540 2237
rect 534 2232 535 2236
rect 539 2232 540 2236
rect 534 2231 540 2232
rect 614 2236 620 2237
rect 614 2232 615 2236
rect 619 2232 620 2236
rect 614 2231 620 2232
rect 694 2236 700 2237
rect 694 2232 695 2236
rect 699 2232 700 2236
rect 694 2231 700 2232
rect 774 2236 780 2237
rect 774 2232 775 2236
rect 779 2232 780 2236
rect 774 2231 780 2232
rect 854 2236 860 2237
rect 854 2232 855 2236
rect 859 2232 860 2236
rect 854 2231 860 2232
rect 934 2236 940 2237
rect 934 2232 935 2236
rect 939 2232 940 2236
rect 934 2231 940 2232
rect 1014 2236 1020 2237
rect 1014 2232 1015 2236
rect 1019 2232 1020 2236
rect 1014 2231 1020 2232
rect 1094 2236 1100 2237
rect 1094 2232 1095 2236
rect 1099 2232 1100 2236
rect 1094 2231 1100 2232
rect 1174 2236 1180 2237
rect 1174 2232 1175 2236
rect 1179 2232 1180 2236
rect 1174 2231 1180 2232
rect 1254 2236 1260 2237
rect 1254 2232 1255 2236
rect 1259 2232 1260 2236
rect 1254 2231 1260 2232
rect 1830 2233 1836 2234
rect 110 2228 116 2229
rect 1830 2229 1831 2233
rect 1835 2229 1836 2233
rect 1830 2228 1836 2229
rect 2310 2220 2316 2221
rect 1870 2217 1876 2218
rect 110 2216 116 2217
rect 110 2212 111 2216
rect 115 2212 116 2216
rect 110 2211 116 2212
rect 1830 2216 1836 2217
rect 1830 2212 1831 2216
rect 1835 2212 1836 2216
rect 1870 2213 1871 2217
rect 1875 2213 1876 2217
rect 2310 2216 2311 2220
rect 2315 2216 2316 2220
rect 2310 2215 2316 2216
rect 2398 2220 2404 2221
rect 2398 2216 2399 2220
rect 2403 2216 2404 2220
rect 2398 2215 2404 2216
rect 2494 2220 2500 2221
rect 2494 2216 2495 2220
rect 2499 2216 2500 2220
rect 2494 2215 2500 2216
rect 2598 2220 2604 2221
rect 2598 2216 2599 2220
rect 2603 2216 2604 2220
rect 2598 2215 2604 2216
rect 2718 2220 2724 2221
rect 2718 2216 2719 2220
rect 2723 2216 2724 2220
rect 2718 2215 2724 2216
rect 2854 2220 2860 2221
rect 2854 2216 2855 2220
rect 2859 2216 2860 2220
rect 2854 2215 2860 2216
rect 3006 2220 3012 2221
rect 3006 2216 3007 2220
rect 3011 2216 3012 2220
rect 3006 2215 3012 2216
rect 3174 2220 3180 2221
rect 3174 2216 3175 2220
rect 3179 2216 3180 2220
rect 3174 2215 3180 2216
rect 3350 2220 3356 2221
rect 3350 2216 3351 2220
rect 3355 2216 3356 2220
rect 3350 2215 3356 2216
rect 3502 2220 3508 2221
rect 3502 2216 3503 2220
rect 3507 2216 3508 2220
rect 3502 2215 3508 2216
rect 3590 2217 3596 2218
rect 1870 2212 1876 2213
rect 3590 2213 3591 2217
rect 3595 2213 3596 2217
rect 3590 2212 3596 2213
rect 1830 2211 1836 2212
rect 1870 2200 1876 2201
rect 382 2198 388 2199
rect 382 2194 383 2198
rect 387 2194 388 2198
rect 382 2193 388 2194
rect 462 2198 468 2199
rect 462 2194 463 2198
rect 467 2194 468 2198
rect 462 2193 468 2194
rect 542 2198 548 2199
rect 542 2194 543 2198
rect 547 2194 548 2198
rect 542 2193 548 2194
rect 622 2198 628 2199
rect 622 2194 623 2198
rect 627 2194 628 2198
rect 622 2193 628 2194
rect 702 2198 708 2199
rect 702 2194 703 2198
rect 707 2194 708 2198
rect 702 2193 708 2194
rect 782 2198 788 2199
rect 782 2194 783 2198
rect 787 2194 788 2198
rect 782 2193 788 2194
rect 862 2198 868 2199
rect 862 2194 863 2198
rect 867 2194 868 2198
rect 862 2193 868 2194
rect 942 2198 948 2199
rect 942 2194 943 2198
rect 947 2194 948 2198
rect 942 2193 948 2194
rect 1022 2198 1028 2199
rect 1022 2194 1023 2198
rect 1027 2194 1028 2198
rect 1022 2193 1028 2194
rect 1102 2198 1108 2199
rect 1102 2194 1103 2198
rect 1107 2194 1108 2198
rect 1102 2193 1108 2194
rect 1182 2198 1188 2199
rect 1182 2194 1183 2198
rect 1187 2194 1188 2198
rect 1182 2193 1188 2194
rect 1262 2198 1268 2199
rect 1262 2194 1263 2198
rect 1267 2194 1268 2198
rect 1870 2196 1871 2200
rect 1875 2196 1876 2200
rect 1870 2195 1876 2196
rect 3590 2200 3596 2201
rect 3590 2196 3591 2200
rect 3595 2196 3596 2200
rect 3590 2195 3596 2196
rect 1262 2193 1268 2194
rect 2318 2182 2324 2183
rect 2318 2178 2319 2182
rect 2323 2178 2324 2182
rect 2318 2177 2324 2178
rect 2406 2182 2412 2183
rect 2406 2178 2407 2182
rect 2411 2178 2412 2182
rect 2406 2177 2412 2178
rect 2502 2182 2508 2183
rect 2502 2178 2503 2182
rect 2507 2178 2508 2182
rect 2502 2177 2508 2178
rect 2606 2182 2612 2183
rect 2606 2178 2607 2182
rect 2611 2178 2612 2182
rect 2606 2177 2612 2178
rect 2726 2182 2732 2183
rect 2726 2178 2727 2182
rect 2731 2178 2732 2182
rect 2726 2177 2732 2178
rect 2862 2182 2868 2183
rect 2862 2178 2863 2182
rect 2867 2178 2868 2182
rect 2862 2177 2868 2178
rect 3014 2182 3020 2183
rect 3014 2178 3015 2182
rect 3019 2178 3020 2182
rect 3014 2177 3020 2178
rect 3182 2182 3188 2183
rect 3182 2178 3183 2182
rect 3187 2178 3188 2182
rect 3182 2177 3188 2178
rect 3358 2182 3364 2183
rect 3358 2178 3359 2182
rect 3363 2178 3364 2182
rect 3358 2177 3364 2178
rect 3510 2182 3516 2183
rect 3510 2178 3511 2182
rect 3515 2178 3516 2182
rect 3510 2177 3516 2178
rect 310 2154 316 2155
rect 310 2150 311 2154
rect 315 2150 316 2154
rect 310 2149 316 2150
rect 406 2154 412 2155
rect 406 2150 407 2154
rect 411 2150 412 2154
rect 406 2149 412 2150
rect 502 2154 508 2155
rect 502 2150 503 2154
rect 507 2150 508 2154
rect 502 2149 508 2150
rect 598 2154 604 2155
rect 598 2150 599 2154
rect 603 2150 604 2154
rect 598 2149 604 2150
rect 686 2154 692 2155
rect 686 2150 687 2154
rect 691 2150 692 2154
rect 686 2149 692 2150
rect 774 2154 780 2155
rect 774 2150 775 2154
rect 779 2150 780 2154
rect 774 2149 780 2150
rect 862 2154 868 2155
rect 862 2150 863 2154
rect 867 2150 868 2154
rect 862 2149 868 2150
rect 950 2154 956 2155
rect 950 2150 951 2154
rect 955 2150 956 2154
rect 950 2149 956 2150
rect 1038 2154 1044 2155
rect 1038 2150 1039 2154
rect 1043 2150 1044 2154
rect 1038 2149 1044 2150
rect 1126 2154 1132 2155
rect 1126 2150 1127 2154
rect 1131 2150 1132 2154
rect 1126 2149 1132 2150
rect 1222 2154 1228 2155
rect 1222 2150 1223 2154
rect 1227 2150 1228 2154
rect 1222 2149 1228 2150
rect 1902 2146 1908 2147
rect 1902 2142 1903 2146
rect 1907 2142 1908 2146
rect 1902 2141 1908 2142
rect 1982 2146 1988 2147
rect 1982 2142 1983 2146
rect 1987 2142 1988 2146
rect 1982 2141 1988 2142
rect 2110 2146 2116 2147
rect 2110 2142 2111 2146
rect 2115 2142 2116 2146
rect 2110 2141 2116 2142
rect 2246 2146 2252 2147
rect 2246 2142 2247 2146
rect 2251 2142 2252 2146
rect 2246 2141 2252 2142
rect 2390 2146 2396 2147
rect 2390 2142 2391 2146
rect 2395 2142 2396 2146
rect 2390 2141 2396 2142
rect 2542 2146 2548 2147
rect 2542 2142 2543 2146
rect 2547 2142 2548 2146
rect 2542 2141 2548 2142
rect 2694 2146 2700 2147
rect 2694 2142 2695 2146
rect 2699 2142 2700 2146
rect 2694 2141 2700 2142
rect 2846 2146 2852 2147
rect 2846 2142 2847 2146
rect 2851 2142 2852 2146
rect 2846 2141 2852 2142
rect 3006 2146 3012 2147
rect 3006 2142 3007 2146
rect 3011 2142 3012 2146
rect 3006 2141 3012 2142
rect 3174 2146 3180 2147
rect 3174 2142 3175 2146
rect 3179 2142 3180 2146
rect 3174 2141 3180 2142
rect 3350 2146 3356 2147
rect 3350 2142 3351 2146
rect 3355 2142 3356 2146
rect 3350 2141 3356 2142
rect 3510 2146 3516 2147
rect 3510 2142 3511 2146
rect 3515 2142 3516 2146
rect 3510 2141 3516 2142
rect 110 2136 116 2137
rect 110 2132 111 2136
rect 115 2132 116 2136
rect 110 2131 116 2132
rect 1830 2136 1836 2137
rect 1830 2132 1831 2136
rect 1835 2132 1836 2136
rect 1830 2131 1836 2132
rect 1870 2128 1876 2129
rect 1870 2124 1871 2128
rect 1875 2124 1876 2128
rect 1870 2123 1876 2124
rect 3590 2128 3596 2129
rect 3590 2124 3591 2128
rect 3595 2124 3596 2128
rect 3590 2123 3596 2124
rect 110 2119 116 2120
rect 110 2115 111 2119
rect 115 2115 116 2119
rect 1830 2119 1836 2120
rect 110 2114 116 2115
rect 302 2116 308 2117
rect 302 2112 303 2116
rect 307 2112 308 2116
rect 302 2111 308 2112
rect 398 2116 404 2117
rect 398 2112 399 2116
rect 403 2112 404 2116
rect 398 2111 404 2112
rect 494 2116 500 2117
rect 494 2112 495 2116
rect 499 2112 500 2116
rect 494 2111 500 2112
rect 590 2116 596 2117
rect 590 2112 591 2116
rect 595 2112 596 2116
rect 590 2111 596 2112
rect 678 2116 684 2117
rect 678 2112 679 2116
rect 683 2112 684 2116
rect 678 2111 684 2112
rect 766 2116 772 2117
rect 766 2112 767 2116
rect 771 2112 772 2116
rect 766 2111 772 2112
rect 854 2116 860 2117
rect 854 2112 855 2116
rect 859 2112 860 2116
rect 854 2111 860 2112
rect 942 2116 948 2117
rect 942 2112 943 2116
rect 947 2112 948 2116
rect 942 2111 948 2112
rect 1030 2116 1036 2117
rect 1030 2112 1031 2116
rect 1035 2112 1036 2116
rect 1030 2111 1036 2112
rect 1118 2116 1124 2117
rect 1118 2112 1119 2116
rect 1123 2112 1124 2116
rect 1118 2111 1124 2112
rect 1214 2116 1220 2117
rect 1214 2112 1215 2116
rect 1219 2112 1220 2116
rect 1830 2115 1831 2119
rect 1835 2115 1836 2119
rect 1830 2114 1836 2115
rect 1214 2111 1220 2112
rect 1870 2111 1876 2112
rect 1870 2107 1871 2111
rect 1875 2107 1876 2111
rect 3590 2111 3596 2112
rect 1870 2106 1876 2107
rect 1894 2108 1900 2109
rect 1894 2104 1895 2108
rect 1899 2104 1900 2108
rect 1894 2103 1900 2104
rect 1974 2108 1980 2109
rect 1974 2104 1975 2108
rect 1979 2104 1980 2108
rect 1974 2103 1980 2104
rect 2102 2108 2108 2109
rect 2102 2104 2103 2108
rect 2107 2104 2108 2108
rect 2102 2103 2108 2104
rect 2238 2108 2244 2109
rect 2238 2104 2239 2108
rect 2243 2104 2244 2108
rect 2238 2103 2244 2104
rect 2382 2108 2388 2109
rect 2382 2104 2383 2108
rect 2387 2104 2388 2108
rect 2382 2103 2388 2104
rect 2534 2108 2540 2109
rect 2534 2104 2535 2108
rect 2539 2104 2540 2108
rect 2534 2103 2540 2104
rect 2686 2108 2692 2109
rect 2686 2104 2687 2108
rect 2691 2104 2692 2108
rect 2686 2103 2692 2104
rect 2838 2108 2844 2109
rect 2838 2104 2839 2108
rect 2843 2104 2844 2108
rect 2838 2103 2844 2104
rect 2998 2108 3004 2109
rect 2998 2104 2999 2108
rect 3003 2104 3004 2108
rect 2998 2103 3004 2104
rect 3166 2108 3172 2109
rect 3166 2104 3167 2108
rect 3171 2104 3172 2108
rect 3166 2103 3172 2104
rect 3342 2108 3348 2109
rect 3342 2104 3343 2108
rect 3347 2104 3348 2108
rect 3342 2103 3348 2104
rect 3502 2108 3508 2109
rect 3502 2104 3503 2108
rect 3507 2104 3508 2108
rect 3590 2107 3591 2111
rect 3595 2107 3596 2111
rect 3590 2106 3596 2107
rect 3502 2103 3508 2104
rect 206 2060 212 2061
rect 110 2057 116 2058
rect 110 2053 111 2057
rect 115 2053 116 2057
rect 206 2056 207 2060
rect 211 2056 212 2060
rect 206 2055 212 2056
rect 326 2060 332 2061
rect 326 2056 327 2060
rect 331 2056 332 2060
rect 326 2055 332 2056
rect 446 2060 452 2061
rect 446 2056 447 2060
rect 451 2056 452 2060
rect 446 2055 452 2056
rect 574 2060 580 2061
rect 574 2056 575 2060
rect 579 2056 580 2060
rect 574 2055 580 2056
rect 702 2060 708 2061
rect 702 2056 703 2060
rect 707 2056 708 2060
rect 702 2055 708 2056
rect 822 2060 828 2061
rect 822 2056 823 2060
rect 827 2056 828 2060
rect 822 2055 828 2056
rect 942 2060 948 2061
rect 942 2056 943 2060
rect 947 2056 948 2060
rect 942 2055 948 2056
rect 1062 2060 1068 2061
rect 1062 2056 1063 2060
rect 1067 2056 1068 2060
rect 1062 2055 1068 2056
rect 1174 2060 1180 2061
rect 1174 2056 1175 2060
rect 1179 2056 1180 2060
rect 1174 2055 1180 2056
rect 1278 2060 1284 2061
rect 1278 2056 1279 2060
rect 1283 2056 1284 2060
rect 1278 2055 1284 2056
rect 1374 2060 1380 2061
rect 1374 2056 1375 2060
rect 1379 2056 1380 2060
rect 1374 2055 1380 2056
rect 1470 2060 1476 2061
rect 1470 2056 1471 2060
rect 1475 2056 1476 2060
rect 1470 2055 1476 2056
rect 1566 2060 1572 2061
rect 1566 2056 1567 2060
rect 1571 2056 1572 2060
rect 1566 2055 1572 2056
rect 1662 2060 1668 2061
rect 1662 2056 1663 2060
rect 1667 2056 1668 2060
rect 1662 2055 1668 2056
rect 1742 2060 1748 2061
rect 1742 2056 1743 2060
rect 1747 2056 1748 2060
rect 1742 2055 1748 2056
rect 1830 2057 1836 2058
rect 110 2052 116 2053
rect 1830 2053 1831 2057
rect 1835 2053 1836 2057
rect 1966 2056 1972 2057
rect 1830 2052 1836 2053
rect 1870 2053 1876 2054
rect 1870 2049 1871 2053
rect 1875 2049 1876 2053
rect 1966 2052 1967 2056
rect 1971 2052 1972 2056
rect 1966 2051 1972 2052
rect 2214 2056 2220 2057
rect 2214 2052 2215 2056
rect 2219 2052 2220 2056
rect 2214 2051 2220 2052
rect 2446 2056 2452 2057
rect 2446 2052 2447 2056
rect 2451 2052 2452 2056
rect 2446 2051 2452 2052
rect 2654 2056 2660 2057
rect 2654 2052 2655 2056
rect 2659 2052 2660 2056
rect 2654 2051 2660 2052
rect 2838 2056 2844 2057
rect 2838 2052 2839 2056
rect 2843 2052 2844 2056
rect 2838 2051 2844 2052
rect 2998 2056 3004 2057
rect 2998 2052 2999 2056
rect 3003 2052 3004 2056
rect 2998 2051 3004 2052
rect 3142 2056 3148 2057
rect 3142 2052 3143 2056
rect 3147 2052 3148 2056
rect 3142 2051 3148 2052
rect 3270 2056 3276 2057
rect 3270 2052 3271 2056
rect 3275 2052 3276 2056
rect 3270 2051 3276 2052
rect 3398 2056 3404 2057
rect 3398 2052 3399 2056
rect 3403 2052 3404 2056
rect 3398 2051 3404 2052
rect 3502 2056 3508 2057
rect 3502 2052 3503 2056
rect 3507 2052 3508 2056
rect 3502 2051 3508 2052
rect 3590 2053 3596 2054
rect 1870 2048 1876 2049
rect 3590 2049 3591 2053
rect 3595 2049 3596 2053
rect 3590 2048 3596 2049
rect 110 2040 116 2041
rect 110 2036 111 2040
rect 115 2036 116 2040
rect 110 2035 116 2036
rect 1830 2040 1836 2041
rect 1830 2036 1831 2040
rect 1835 2036 1836 2040
rect 1830 2035 1836 2036
rect 1870 2036 1876 2037
rect 1870 2032 1871 2036
rect 1875 2032 1876 2036
rect 1870 2031 1876 2032
rect 3590 2036 3596 2037
rect 3590 2032 3591 2036
rect 3595 2032 3596 2036
rect 3590 2031 3596 2032
rect 214 2022 220 2023
rect 214 2018 215 2022
rect 219 2018 220 2022
rect 214 2017 220 2018
rect 334 2022 340 2023
rect 334 2018 335 2022
rect 339 2018 340 2022
rect 334 2017 340 2018
rect 454 2022 460 2023
rect 454 2018 455 2022
rect 459 2018 460 2022
rect 454 2017 460 2018
rect 582 2022 588 2023
rect 582 2018 583 2022
rect 587 2018 588 2022
rect 582 2017 588 2018
rect 710 2022 716 2023
rect 710 2018 711 2022
rect 715 2018 716 2022
rect 710 2017 716 2018
rect 830 2022 836 2023
rect 830 2018 831 2022
rect 835 2018 836 2022
rect 830 2017 836 2018
rect 950 2022 956 2023
rect 950 2018 951 2022
rect 955 2018 956 2022
rect 950 2017 956 2018
rect 1070 2022 1076 2023
rect 1070 2018 1071 2022
rect 1075 2018 1076 2022
rect 1070 2017 1076 2018
rect 1182 2022 1188 2023
rect 1182 2018 1183 2022
rect 1187 2018 1188 2022
rect 1182 2017 1188 2018
rect 1286 2022 1292 2023
rect 1286 2018 1287 2022
rect 1291 2018 1292 2022
rect 1286 2017 1292 2018
rect 1382 2022 1388 2023
rect 1382 2018 1383 2022
rect 1387 2018 1388 2022
rect 1382 2017 1388 2018
rect 1478 2022 1484 2023
rect 1478 2018 1479 2022
rect 1483 2018 1484 2022
rect 1478 2017 1484 2018
rect 1574 2022 1580 2023
rect 1574 2018 1575 2022
rect 1579 2018 1580 2022
rect 1574 2017 1580 2018
rect 1670 2022 1676 2023
rect 1670 2018 1671 2022
rect 1675 2018 1676 2022
rect 1670 2017 1676 2018
rect 1750 2022 1756 2023
rect 1750 2018 1751 2022
rect 1755 2018 1756 2022
rect 1750 2017 1756 2018
rect 1974 2018 1980 2019
rect 1974 2014 1975 2018
rect 1979 2014 1980 2018
rect 1974 2013 1980 2014
rect 2222 2018 2228 2019
rect 2222 2014 2223 2018
rect 2227 2014 2228 2018
rect 2222 2013 2228 2014
rect 2454 2018 2460 2019
rect 2454 2014 2455 2018
rect 2459 2014 2460 2018
rect 2454 2013 2460 2014
rect 2662 2018 2668 2019
rect 2662 2014 2663 2018
rect 2667 2014 2668 2018
rect 2662 2013 2668 2014
rect 2846 2018 2852 2019
rect 2846 2014 2847 2018
rect 2851 2014 2852 2018
rect 2846 2013 2852 2014
rect 3006 2018 3012 2019
rect 3006 2014 3007 2018
rect 3011 2014 3012 2018
rect 3006 2013 3012 2014
rect 3150 2018 3156 2019
rect 3150 2014 3151 2018
rect 3155 2014 3156 2018
rect 3150 2013 3156 2014
rect 3278 2018 3284 2019
rect 3278 2014 3279 2018
rect 3283 2014 3284 2018
rect 3278 2013 3284 2014
rect 3406 2018 3412 2019
rect 3406 2014 3407 2018
rect 3411 2014 3412 2018
rect 3406 2013 3412 2014
rect 3510 2018 3516 2019
rect 3510 2014 3511 2018
rect 3515 2014 3516 2018
rect 3510 2013 3516 2014
rect 190 1986 196 1987
rect 190 1982 191 1986
rect 195 1982 196 1986
rect 190 1981 196 1982
rect 350 1986 356 1987
rect 350 1982 351 1986
rect 355 1982 356 1986
rect 350 1981 356 1982
rect 518 1986 524 1987
rect 518 1982 519 1986
rect 523 1982 524 1986
rect 518 1981 524 1982
rect 686 1986 692 1987
rect 686 1982 687 1986
rect 691 1982 692 1986
rect 686 1981 692 1982
rect 854 1986 860 1987
rect 854 1982 855 1986
rect 859 1982 860 1986
rect 854 1981 860 1982
rect 1014 1986 1020 1987
rect 1014 1982 1015 1986
rect 1019 1982 1020 1986
rect 1014 1981 1020 1982
rect 1166 1986 1172 1987
rect 1166 1982 1167 1986
rect 1171 1982 1172 1986
rect 1166 1981 1172 1982
rect 1310 1986 1316 1987
rect 1310 1982 1311 1986
rect 1315 1982 1316 1986
rect 1310 1981 1316 1982
rect 1446 1986 1452 1987
rect 1446 1982 1447 1986
rect 1451 1982 1452 1986
rect 1446 1981 1452 1982
rect 1582 1986 1588 1987
rect 1582 1982 1583 1986
rect 1587 1982 1588 1986
rect 1582 1981 1588 1982
rect 1718 1986 1724 1987
rect 1718 1982 1719 1986
rect 1723 1982 1724 1986
rect 1718 1981 1724 1982
rect 1958 1986 1964 1987
rect 1958 1982 1959 1986
rect 1963 1982 1964 1986
rect 1958 1981 1964 1982
rect 2078 1986 2084 1987
rect 2078 1982 2079 1986
rect 2083 1982 2084 1986
rect 2078 1981 2084 1982
rect 2198 1986 2204 1987
rect 2198 1982 2199 1986
rect 2203 1982 2204 1986
rect 2198 1981 2204 1982
rect 2318 1986 2324 1987
rect 2318 1982 2319 1986
rect 2323 1982 2324 1986
rect 2318 1981 2324 1982
rect 2446 1986 2452 1987
rect 2446 1982 2447 1986
rect 2451 1982 2452 1986
rect 2446 1981 2452 1982
rect 2582 1986 2588 1987
rect 2582 1982 2583 1986
rect 2587 1982 2588 1986
rect 2582 1981 2588 1982
rect 2742 1986 2748 1987
rect 2742 1982 2743 1986
rect 2747 1982 2748 1986
rect 2742 1981 2748 1982
rect 2918 1986 2924 1987
rect 2918 1982 2919 1986
rect 2923 1982 2924 1986
rect 2918 1981 2924 1982
rect 3118 1986 3124 1987
rect 3118 1982 3119 1986
rect 3123 1982 3124 1986
rect 3118 1981 3124 1982
rect 3326 1986 3332 1987
rect 3326 1982 3327 1986
rect 3331 1982 3332 1986
rect 3326 1981 3332 1982
rect 3510 1986 3516 1987
rect 3510 1982 3511 1986
rect 3515 1982 3516 1986
rect 3510 1981 3516 1982
rect 110 1968 116 1969
rect 110 1964 111 1968
rect 115 1964 116 1968
rect 110 1963 116 1964
rect 1830 1968 1836 1969
rect 1830 1964 1831 1968
rect 1835 1964 1836 1968
rect 1830 1963 1836 1964
rect 1870 1968 1876 1969
rect 1870 1964 1871 1968
rect 1875 1964 1876 1968
rect 1870 1963 1876 1964
rect 3590 1968 3596 1969
rect 3590 1964 3591 1968
rect 3595 1964 3596 1968
rect 3590 1963 3596 1964
rect 110 1951 116 1952
rect 110 1947 111 1951
rect 115 1947 116 1951
rect 1830 1951 1836 1952
rect 110 1946 116 1947
rect 182 1948 188 1949
rect 182 1944 183 1948
rect 187 1944 188 1948
rect 182 1943 188 1944
rect 342 1948 348 1949
rect 342 1944 343 1948
rect 347 1944 348 1948
rect 342 1943 348 1944
rect 510 1948 516 1949
rect 510 1944 511 1948
rect 515 1944 516 1948
rect 510 1943 516 1944
rect 678 1948 684 1949
rect 678 1944 679 1948
rect 683 1944 684 1948
rect 678 1943 684 1944
rect 846 1948 852 1949
rect 846 1944 847 1948
rect 851 1944 852 1948
rect 846 1943 852 1944
rect 1006 1948 1012 1949
rect 1006 1944 1007 1948
rect 1011 1944 1012 1948
rect 1006 1943 1012 1944
rect 1158 1948 1164 1949
rect 1158 1944 1159 1948
rect 1163 1944 1164 1948
rect 1158 1943 1164 1944
rect 1302 1948 1308 1949
rect 1302 1944 1303 1948
rect 1307 1944 1308 1948
rect 1302 1943 1308 1944
rect 1438 1948 1444 1949
rect 1438 1944 1439 1948
rect 1443 1944 1444 1948
rect 1438 1943 1444 1944
rect 1574 1948 1580 1949
rect 1574 1944 1575 1948
rect 1579 1944 1580 1948
rect 1574 1943 1580 1944
rect 1710 1948 1716 1949
rect 1710 1944 1711 1948
rect 1715 1944 1716 1948
rect 1830 1947 1831 1951
rect 1835 1947 1836 1951
rect 1830 1946 1836 1947
rect 1870 1951 1876 1952
rect 1870 1947 1871 1951
rect 1875 1947 1876 1951
rect 3590 1951 3596 1952
rect 1870 1946 1876 1947
rect 1950 1948 1956 1949
rect 1710 1943 1716 1944
rect 1950 1944 1951 1948
rect 1955 1944 1956 1948
rect 1950 1943 1956 1944
rect 2070 1948 2076 1949
rect 2070 1944 2071 1948
rect 2075 1944 2076 1948
rect 2070 1943 2076 1944
rect 2190 1948 2196 1949
rect 2190 1944 2191 1948
rect 2195 1944 2196 1948
rect 2190 1943 2196 1944
rect 2310 1948 2316 1949
rect 2310 1944 2311 1948
rect 2315 1944 2316 1948
rect 2310 1943 2316 1944
rect 2438 1948 2444 1949
rect 2438 1944 2439 1948
rect 2443 1944 2444 1948
rect 2438 1943 2444 1944
rect 2574 1948 2580 1949
rect 2574 1944 2575 1948
rect 2579 1944 2580 1948
rect 2574 1943 2580 1944
rect 2734 1948 2740 1949
rect 2734 1944 2735 1948
rect 2739 1944 2740 1948
rect 2734 1943 2740 1944
rect 2910 1948 2916 1949
rect 2910 1944 2911 1948
rect 2915 1944 2916 1948
rect 2910 1943 2916 1944
rect 3110 1948 3116 1949
rect 3110 1944 3111 1948
rect 3115 1944 3116 1948
rect 3110 1943 3116 1944
rect 3318 1948 3324 1949
rect 3318 1944 3319 1948
rect 3323 1944 3324 1948
rect 3318 1943 3324 1944
rect 3502 1948 3508 1949
rect 3502 1944 3503 1948
rect 3507 1944 3508 1948
rect 3590 1947 3591 1951
rect 3595 1947 3596 1951
rect 3590 1946 3596 1947
rect 3502 1943 3508 1944
rect 134 1900 140 1901
rect 110 1897 116 1898
rect 110 1893 111 1897
rect 115 1893 116 1897
rect 134 1896 135 1900
rect 139 1896 140 1900
rect 134 1895 140 1896
rect 238 1900 244 1901
rect 238 1896 239 1900
rect 243 1896 244 1900
rect 238 1895 244 1896
rect 374 1900 380 1901
rect 374 1896 375 1900
rect 379 1896 380 1900
rect 374 1895 380 1896
rect 526 1900 532 1901
rect 526 1896 527 1900
rect 531 1896 532 1900
rect 526 1895 532 1896
rect 686 1900 692 1901
rect 686 1896 687 1900
rect 691 1896 692 1900
rect 686 1895 692 1896
rect 846 1900 852 1901
rect 846 1896 847 1900
rect 851 1896 852 1900
rect 846 1895 852 1896
rect 1006 1900 1012 1901
rect 1006 1896 1007 1900
rect 1011 1896 1012 1900
rect 1006 1895 1012 1896
rect 1158 1900 1164 1901
rect 1158 1896 1159 1900
rect 1163 1896 1164 1900
rect 1158 1895 1164 1896
rect 1302 1900 1308 1901
rect 1302 1896 1303 1900
rect 1307 1896 1308 1900
rect 1302 1895 1308 1896
rect 1454 1900 1460 1901
rect 1454 1896 1455 1900
rect 1459 1896 1460 1900
rect 1454 1895 1460 1896
rect 1606 1900 1612 1901
rect 1606 1896 1607 1900
rect 1611 1896 1612 1900
rect 1606 1895 1612 1896
rect 1830 1897 1836 1898
rect 110 1892 116 1893
rect 1830 1893 1831 1897
rect 1835 1893 1836 1897
rect 2062 1896 2068 1897
rect 1830 1892 1836 1893
rect 1870 1893 1876 1894
rect 1870 1889 1871 1893
rect 1875 1889 1876 1893
rect 2062 1892 2063 1896
rect 2067 1892 2068 1896
rect 2062 1891 2068 1892
rect 2150 1896 2156 1897
rect 2150 1892 2151 1896
rect 2155 1892 2156 1896
rect 2150 1891 2156 1892
rect 2238 1896 2244 1897
rect 2238 1892 2239 1896
rect 2243 1892 2244 1896
rect 2238 1891 2244 1892
rect 2318 1896 2324 1897
rect 2318 1892 2319 1896
rect 2323 1892 2324 1896
rect 2318 1891 2324 1892
rect 2398 1896 2404 1897
rect 2398 1892 2399 1896
rect 2403 1892 2404 1896
rect 2398 1891 2404 1892
rect 2486 1896 2492 1897
rect 2486 1892 2487 1896
rect 2491 1892 2492 1896
rect 2486 1891 2492 1892
rect 2574 1896 2580 1897
rect 2574 1892 2575 1896
rect 2579 1892 2580 1896
rect 2574 1891 2580 1892
rect 2662 1896 2668 1897
rect 2662 1892 2663 1896
rect 2667 1892 2668 1896
rect 2662 1891 2668 1892
rect 2758 1896 2764 1897
rect 2758 1892 2759 1896
rect 2763 1892 2764 1896
rect 2758 1891 2764 1892
rect 2870 1896 2876 1897
rect 2870 1892 2871 1896
rect 2875 1892 2876 1896
rect 2870 1891 2876 1892
rect 2990 1896 2996 1897
rect 2990 1892 2991 1896
rect 2995 1892 2996 1896
rect 2990 1891 2996 1892
rect 3118 1896 3124 1897
rect 3118 1892 3119 1896
rect 3123 1892 3124 1896
rect 3118 1891 3124 1892
rect 3246 1896 3252 1897
rect 3246 1892 3247 1896
rect 3251 1892 3252 1896
rect 3246 1891 3252 1892
rect 3382 1896 3388 1897
rect 3382 1892 3383 1896
rect 3387 1892 3388 1896
rect 3382 1891 3388 1892
rect 3502 1896 3508 1897
rect 3502 1892 3503 1896
rect 3507 1892 3508 1896
rect 3502 1891 3508 1892
rect 3590 1893 3596 1894
rect 1870 1888 1876 1889
rect 3590 1889 3591 1893
rect 3595 1889 3596 1893
rect 3590 1888 3596 1889
rect 110 1880 116 1881
rect 110 1876 111 1880
rect 115 1876 116 1880
rect 110 1875 116 1876
rect 1830 1880 1836 1881
rect 1830 1876 1831 1880
rect 1835 1876 1836 1880
rect 1830 1875 1836 1876
rect 1870 1876 1876 1877
rect 1870 1872 1871 1876
rect 1875 1872 1876 1876
rect 1870 1871 1876 1872
rect 3590 1876 3596 1877
rect 3590 1872 3591 1876
rect 3595 1872 3596 1876
rect 3590 1871 3596 1872
rect 142 1862 148 1863
rect 142 1858 143 1862
rect 147 1858 148 1862
rect 142 1857 148 1858
rect 246 1862 252 1863
rect 246 1858 247 1862
rect 251 1858 252 1862
rect 246 1857 252 1858
rect 382 1862 388 1863
rect 382 1858 383 1862
rect 387 1858 388 1862
rect 382 1857 388 1858
rect 534 1862 540 1863
rect 534 1858 535 1862
rect 539 1858 540 1862
rect 534 1857 540 1858
rect 694 1862 700 1863
rect 694 1858 695 1862
rect 699 1858 700 1862
rect 694 1857 700 1858
rect 854 1862 860 1863
rect 854 1858 855 1862
rect 859 1858 860 1862
rect 854 1857 860 1858
rect 1014 1862 1020 1863
rect 1014 1858 1015 1862
rect 1019 1858 1020 1862
rect 1014 1857 1020 1858
rect 1166 1862 1172 1863
rect 1166 1858 1167 1862
rect 1171 1858 1172 1862
rect 1166 1857 1172 1858
rect 1310 1862 1316 1863
rect 1310 1858 1311 1862
rect 1315 1858 1316 1862
rect 1310 1857 1316 1858
rect 1462 1862 1468 1863
rect 1462 1858 1463 1862
rect 1467 1858 1468 1862
rect 1462 1857 1468 1858
rect 1614 1862 1620 1863
rect 1614 1858 1615 1862
rect 1619 1858 1620 1862
rect 1614 1857 1620 1858
rect 2070 1858 2076 1859
rect 2070 1854 2071 1858
rect 2075 1854 2076 1858
rect 2070 1853 2076 1854
rect 2158 1858 2164 1859
rect 2158 1854 2159 1858
rect 2163 1854 2164 1858
rect 2158 1853 2164 1854
rect 2246 1858 2252 1859
rect 2246 1854 2247 1858
rect 2251 1854 2252 1858
rect 2246 1853 2252 1854
rect 2326 1858 2332 1859
rect 2326 1854 2327 1858
rect 2331 1854 2332 1858
rect 2326 1853 2332 1854
rect 2406 1858 2412 1859
rect 2406 1854 2407 1858
rect 2411 1854 2412 1858
rect 2406 1853 2412 1854
rect 2494 1858 2500 1859
rect 2494 1854 2495 1858
rect 2499 1854 2500 1858
rect 2494 1853 2500 1854
rect 2582 1858 2588 1859
rect 2582 1854 2583 1858
rect 2587 1854 2588 1858
rect 2582 1853 2588 1854
rect 2670 1858 2676 1859
rect 2670 1854 2671 1858
rect 2675 1854 2676 1858
rect 2670 1853 2676 1854
rect 2766 1858 2772 1859
rect 2766 1854 2767 1858
rect 2771 1854 2772 1858
rect 2766 1853 2772 1854
rect 2878 1858 2884 1859
rect 2878 1854 2879 1858
rect 2883 1854 2884 1858
rect 2878 1853 2884 1854
rect 2998 1858 3004 1859
rect 2998 1854 2999 1858
rect 3003 1854 3004 1858
rect 2998 1853 3004 1854
rect 3126 1858 3132 1859
rect 3126 1854 3127 1858
rect 3131 1854 3132 1858
rect 3126 1853 3132 1854
rect 3254 1858 3260 1859
rect 3254 1854 3255 1858
rect 3259 1854 3260 1858
rect 3254 1853 3260 1854
rect 3390 1858 3396 1859
rect 3390 1854 3391 1858
rect 3395 1854 3396 1858
rect 3390 1853 3396 1854
rect 3510 1858 3516 1859
rect 3510 1854 3511 1858
rect 3515 1854 3516 1858
rect 3510 1853 3516 1854
rect 142 1826 148 1827
rect 142 1822 143 1826
rect 147 1822 148 1826
rect 142 1821 148 1822
rect 286 1826 292 1827
rect 286 1822 287 1826
rect 291 1822 292 1826
rect 286 1821 292 1822
rect 470 1826 476 1827
rect 470 1822 471 1826
rect 475 1822 476 1826
rect 470 1821 476 1822
rect 662 1826 668 1827
rect 662 1822 663 1826
rect 667 1822 668 1826
rect 662 1821 668 1822
rect 846 1826 852 1827
rect 846 1822 847 1826
rect 851 1822 852 1826
rect 846 1821 852 1822
rect 1022 1826 1028 1827
rect 1022 1822 1023 1826
rect 1027 1822 1028 1826
rect 1022 1821 1028 1822
rect 1190 1826 1196 1827
rect 1190 1822 1191 1826
rect 1195 1822 1196 1826
rect 1190 1821 1196 1822
rect 1350 1826 1356 1827
rect 1350 1822 1351 1826
rect 1355 1822 1356 1826
rect 1350 1821 1356 1822
rect 1510 1826 1516 1827
rect 1510 1822 1511 1826
rect 1515 1822 1516 1826
rect 1510 1821 1516 1822
rect 1678 1826 1684 1827
rect 1678 1822 1679 1826
rect 1683 1822 1684 1826
rect 1678 1821 1684 1822
rect 2094 1810 2100 1811
rect 110 1808 116 1809
rect 110 1804 111 1808
rect 115 1804 116 1808
rect 110 1803 116 1804
rect 1830 1808 1836 1809
rect 1830 1804 1831 1808
rect 1835 1804 1836 1808
rect 2094 1806 2095 1810
rect 2099 1806 2100 1810
rect 2094 1805 2100 1806
rect 2238 1810 2244 1811
rect 2238 1806 2239 1810
rect 2243 1806 2244 1810
rect 2238 1805 2244 1806
rect 2398 1810 2404 1811
rect 2398 1806 2399 1810
rect 2403 1806 2404 1810
rect 2398 1805 2404 1806
rect 2558 1810 2564 1811
rect 2558 1806 2559 1810
rect 2563 1806 2564 1810
rect 2558 1805 2564 1806
rect 2718 1810 2724 1811
rect 2718 1806 2719 1810
rect 2723 1806 2724 1810
rect 2718 1805 2724 1806
rect 2878 1810 2884 1811
rect 2878 1806 2879 1810
rect 2883 1806 2884 1810
rect 2878 1805 2884 1806
rect 3030 1810 3036 1811
rect 3030 1806 3031 1810
rect 3035 1806 3036 1810
rect 3030 1805 3036 1806
rect 3174 1810 3180 1811
rect 3174 1806 3175 1810
rect 3179 1806 3180 1810
rect 3174 1805 3180 1806
rect 3318 1810 3324 1811
rect 3318 1806 3319 1810
rect 3323 1806 3324 1810
rect 3318 1805 3324 1806
rect 3470 1810 3476 1811
rect 3470 1806 3471 1810
rect 3475 1806 3476 1810
rect 3470 1805 3476 1806
rect 1830 1803 1836 1804
rect 1870 1792 1876 1793
rect 110 1791 116 1792
rect 110 1787 111 1791
rect 115 1787 116 1791
rect 1830 1791 1836 1792
rect 110 1786 116 1787
rect 134 1788 140 1789
rect 134 1784 135 1788
rect 139 1784 140 1788
rect 134 1783 140 1784
rect 278 1788 284 1789
rect 278 1784 279 1788
rect 283 1784 284 1788
rect 278 1783 284 1784
rect 462 1788 468 1789
rect 462 1784 463 1788
rect 467 1784 468 1788
rect 462 1783 468 1784
rect 654 1788 660 1789
rect 654 1784 655 1788
rect 659 1784 660 1788
rect 654 1783 660 1784
rect 838 1788 844 1789
rect 838 1784 839 1788
rect 843 1784 844 1788
rect 838 1783 844 1784
rect 1014 1788 1020 1789
rect 1014 1784 1015 1788
rect 1019 1784 1020 1788
rect 1014 1783 1020 1784
rect 1182 1788 1188 1789
rect 1182 1784 1183 1788
rect 1187 1784 1188 1788
rect 1182 1783 1188 1784
rect 1342 1788 1348 1789
rect 1342 1784 1343 1788
rect 1347 1784 1348 1788
rect 1342 1783 1348 1784
rect 1502 1788 1508 1789
rect 1502 1784 1503 1788
rect 1507 1784 1508 1788
rect 1502 1783 1508 1784
rect 1670 1788 1676 1789
rect 1670 1784 1671 1788
rect 1675 1784 1676 1788
rect 1830 1787 1831 1791
rect 1835 1787 1836 1791
rect 1870 1788 1871 1792
rect 1875 1788 1876 1792
rect 1870 1787 1876 1788
rect 3590 1792 3596 1793
rect 3590 1788 3591 1792
rect 3595 1788 3596 1792
rect 3590 1787 3596 1788
rect 1830 1786 1836 1787
rect 1670 1783 1676 1784
rect 1870 1775 1876 1776
rect 1870 1771 1871 1775
rect 1875 1771 1876 1775
rect 3590 1775 3596 1776
rect 1870 1770 1876 1771
rect 2086 1772 2092 1773
rect 2086 1768 2087 1772
rect 2091 1768 2092 1772
rect 2086 1767 2092 1768
rect 2230 1772 2236 1773
rect 2230 1768 2231 1772
rect 2235 1768 2236 1772
rect 2230 1767 2236 1768
rect 2390 1772 2396 1773
rect 2390 1768 2391 1772
rect 2395 1768 2396 1772
rect 2390 1767 2396 1768
rect 2550 1772 2556 1773
rect 2550 1768 2551 1772
rect 2555 1768 2556 1772
rect 2550 1767 2556 1768
rect 2710 1772 2716 1773
rect 2710 1768 2711 1772
rect 2715 1768 2716 1772
rect 2710 1767 2716 1768
rect 2870 1772 2876 1773
rect 2870 1768 2871 1772
rect 2875 1768 2876 1772
rect 2870 1767 2876 1768
rect 3022 1772 3028 1773
rect 3022 1768 3023 1772
rect 3027 1768 3028 1772
rect 3022 1767 3028 1768
rect 3166 1772 3172 1773
rect 3166 1768 3167 1772
rect 3171 1768 3172 1772
rect 3166 1767 3172 1768
rect 3310 1772 3316 1773
rect 3310 1768 3311 1772
rect 3315 1768 3316 1772
rect 3310 1767 3316 1768
rect 3462 1772 3468 1773
rect 3462 1768 3463 1772
rect 3467 1768 3468 1772
rect 3590 1771 3591 1775
rect 3595 1771 3596 1775
rect 3590 1770 3596 1771
rect 3462 1767 3468 1768
rect 134 1736 140 1737
rect 110 1733 116 1734
rect 110 1729 111 1733
rect 115 1729 116 1733
rect 134 1732 135 1736
rect 139 1732 140 1736
rect 134 1731 140 1732
rect 214 1736 220 1737
rect 214 1732 215 1736
rect 219 1732 220 1736
rect 214 1731 220 1732
rect 342 1736 348 1737
rect 342 1732 343 1736
rect 347 1732 348 1736
rect 342 1731 348 1732
rect 494 1736 500 1737
rect 494 1732 495 1736
rect 499 1732 500 1736
rect 494 1731 500 1732
rect 662 1736 668 1737
rect 662 1732 663 1736
rect 667 1732 668 1736
rect 662 1731 668 1732
rect 838 1736 844 1737
rect 838 1732 839 1736
rect 843 1732 844 1736
rect 838 1731 844 1732
rect 1006 1736 1012 1737
rect 1006 1732 1007 1736
rect 1011 1732 1012 1736
rect 1006 1731 1012 1732
rect 1166 1736 1172 1737
rect 1166 1732 1167 1736
rect 1171 1732 1172 1736
rect 1166 1731 1172 1732
rect 1318 1736 1324 1737
rect 1318 1732 1319 1736
rect 1323 1732 1324 1736
rect 1318 1731 1324 1732
rect 1462 1736 1468 1737
rect 1462 1732 1463 1736
rect 1467 1732 1468 1736
rect 1462 1731 1468 1732
rect 1606 1736 1612 1737
rect 1606 1732 1607 1736
rect 1611 1732 1612 1736
rect 1606 1731 1612 1732
rect 1742 1736 1748 1737
rect 1742 1732 1743 1736
rect 1747 1732 1748 1736
rect 1742 1731 1748 1732
rect 1830 1733 1836 1734
rect 110 1728 116 1729
rect 1830 1729 1831 1733
rect 1835 1729 1836 1733
rect 1830 1728 1836 1729
rect 2102 1724 2108 1725
rect 1870 1721 1876 1722
rect 1870 1717 1871 1721
rect 1875 1717 1876 1721
rect 2102 1720 2103 1724
rect 2107 1720 2108 1724
rect 2102 1719 2108 1720
rect 2238 1724 2244 1725
rect 2238 1720 2239 1724
rect 2243 1720 2244 1724
rect 2238 1719 2244 1720
rect 2382 1724 2388 1725
rect 2382 1720 2383 1724
rect 2387 1720 2388 1724
rect 2382 1719 2388 1720
rect 2526 1724 2532 1725
rect 2526 1720 2527 1724
rect 2531 1720 2532 1724
rect 2526 1719 2532 1720
rect 2662 1724 2668 1725
rect 2662 1720 2663 1724
rect 2667 1720 2668 1724
rect 2662 1719 2668 1720
rect 2798 1724 2804 1725
rect 2798 1720 2799 1724
rect 2803 1720 2804 1724
rect 2798 1719 2804 1720
rect 2926 1724 2932 1725
rect 2926 1720 2927 1724
rect 2931 1720 2932 1724
rect 2926 1719 2932 1720
rect 3046 1724 3052 1725
rect 3046 1720 3047 1724
rect 3051 1720 3052 1724
rect 3046 1719 3052 1720
rect 3158 1724 3164 1725
rect 3158 1720 3159 1724
rect 3163 1720 3164 1724
rect 3158 1719 3164 1720
rect 3270 1724 3276 1725
rect 3270 1720 3271 1724
rect 3275 1720 3276 1724
rect 3270 1719 3276 1720
rect 3390 1724 3396 1725
rect 3390 1720 3391 1724
rect 3395 1720 3396 1724
rect 3390 1719 3396 1720
rect 3502 1724 3508 1725
rect 3502 1720 3503 1724
rect 3507 1720 3508 1724
rect 3502 1719 3508 1720
rect 3590 1721 3596 1722
rect 110 1716 116 1717
rect 110 1712 111 1716
rect 115 1712 116 1716
rect 110 1711 116 1712
rect 1830 1716 1836 1717
rect 1870 1716 1876 1717
rect 3590 1717 3591 1721
rect 3595 1717 3596 1721
rect 3590 1716 3596 1717
rect 1830 1712 1831 1716
rect 1835 1712 1836 1716
rect 1830 1711 1836 1712
rect 1870 1704 1876 1705
rect 1870 1700 1871 1704
rect 1875 1700 1876 1704
rect 1870 1699 1876 1700
rect 3590 1704 3596 1705
rect 3590 1700 3591 1704
rect 3595 1700 3596 1704
rect 3590 1699 3596 1700
rect 142 1698 148 1699
rect 142 1694 143 1698
rect 147 1694 148 1698
rect 142 1693 148 1694
rect 222 1698 228 1699
rect 222 1694 223 1698
rect 227 1694 228 1698
rect 222 1693 228 1694
rect 350 1698 356 1699
rect 350 1694 351 1698
rect 355 1694 356 1698
rect 350 1693 356 1694
rect 502 1698 508 1699
rect 502 1694 503 1698
rect 507 1694 508 1698
rect 502 1693 508 1694
rect 670 1698 676 1699
rect 670 1694 671 1698
rect 675 1694 676 1698
rect 670 1693 676 1694
rect 846 1698 852 1699
rect 846 1694 847 1698
rect 851 1694 852 1698
rect 846 1693 852 1694
rect 1014 1698 1020 1699
rect 1014 1694 1015 1698
rect 1019 1694 1020 1698
rect 1014 1693 1020 1694
rect 1174 1698 1180 1699
rect 1174 1694 1175 1698
rect 1179 1694 1180 1698
rect 1174 1693 1180 1694
rect 1326 1698 1332 1699
rect 1326 1694 1327 1698
rect 1331 1694 1332 1698
rect 1326 1693 1332 1694
rect 1470 1698 1476 1699
rect 1470 1694 1471 1698
rect 1475 1694 1476 1698
rect 1470 1693 1476 1694
rect 1614 1698 1620 1699
rect 1614 1694 1615 1698
rect 1619 1694 1620 1698
rect 1614 1693 1620 1694
rect 1750 1698 1756 1699
rect 1750 1694 1751 1698
rect 1755 1694 1756 1698
rect 1750 1693 1756 1694
rect 2110 1686 2116 1687
rect 2110 1682 2111 1686
rect 2115 1682 2116 1686
rect 2110 1681 2116 1682
rect 2246 1686 2252 1687
rect 2246 1682 2247 1686
rect 2251 1682 2252 1686
rect 2246 1681 2252 1682
rect 2390 1686 2396 1687
rect 2390 1682 2391 1686
rect 2395 1682 2396 1686
rect 2390 1681 2396 1682
rect 2534 1686 2540 1687
rect 2534 1682 2535 1686
rect 2539 1682 2540 1686
rect 2534 1681 2540 1682
rect 2670 1686 2676 1687
rect 2670 1682 2671 1686
rect 2675 1682 2676 1686
rect 2670 1681 2676 1682
rect 2806 1686 2812 1687
rect 2806 1682 2807 1686
rect 2811 1682 2812 1686
rect 2806 1681 2812 1682
rect 2934 1686 2940 1687
rect 2934 1682 2935 1686
rect 2939 1682 2940 1686
rect 2934 1681 2940 1682
rect 3054 1686 3060 1687
rect 3054 1682 3055 1686
rect 3059 1682 3060 1686
rect 3054 1681 3060 1682
rect 3166 1686 3172 1687
rect 3166 1682 3167 1686
rect 3171 1682 3172 1686
rect 3166 1681 3172 1682
rect 3278 1686 3284 1687
rect 3278 1682 3279 1686
rect 3283 1682 3284 1686
rect 3278 1681 3284 1682
rect 3398 1686 3404 1687
rect 3398 1682 3399 1686
rect 3403 1682 3404 1686
rect 3398 1681 3404 1682
rect 3510 1686 3516 1687
rect 3510 1682 3511 1686
rect 3515 1682 3516 1686
rect 3510 1681 3516 1682
rect 142 1662 148 1663
rect 142 1658 143 1662
rect 147 1658 148 1662
rect 142 1657 148 1658
rect 294 1662 300 1663
rect 294 1658 295 1662
rect 299 1658 300 1662
rect 294 1657 300 1658
rect 478 1662 484 1663
rect 478 1658 479 1662
rect 483 1658 484 1662
rect 478 1657 484 1658
rect 670 1662 676 1663
rect 670 1658 671 1662
rect 675 1658 676 1662
rect 670 1657 676 1658
rect 854 1662 860 1663
rect 854 1658 855 1662
rect 859 1658 860 1662
rect 854 1657 860 1658
rect 1030 1662 1036 1663
rect 1030 1658 1031 1662
rect 1035 1658 1036 1662
rect 1030 1657 1036 1658
rect 1198 1662 1204 1663
rect 1198 1658 1199 1662
rect 1203 1658 1204 1662
rect 1198 1657 1204 1658
rect 1358 1662 1364 1663
rect 1358 1658 1359 1662
rect 1363 1658 1364 1662
rect 1358 1657 1364 1658
rect 1518 1662 1524 1663
rect 1518 1658 1519 1662
rect 1523 1658 1524 1662
rect 1518 1657 1524 1658
rect 1678 1662 1684 1663
rect 1678 1658 1679 1662
rect 1683 1658 1684 1662
rect 1678 1657 1684 1658
rect 1966 1650 1972 1651
rect 1966 1646 1967 1650
rect 1971 1646 1972 1650
rect 1966 1645 1972 1646
rect 2086 1650 2092 1651
rect 2086 1646 2087 1650
rect 2091 1646 2092 1650
rect 2086 1645 2092 1646
rect 2214 1650 2220 1651
rect 2214 1646 2215 1650
rect 2219 1646 2220 1650
rect 2214 1645 2220 1646
rect 2350 1650 2356 1651
rect 2350 1646 2351 1650
rect 2355 1646 2356 1650
rect 2350 1645 2356 1646
rect 2494 1650 2500 1651
rect 2494 1646 2495 1650
rect 2499 1646 2500 1650
rect 2494 1645 2500 1646
rect 2638 1650 2644 1651
rect 2638 1646 2639 1650
rect 2643 1646 2644 1650
rect 2638 1645 2644 1646
rect 2782 1650 2788 1651
rect 2782 1646 2783 1650
rect 2787 1646 2788 1650
rect 2782 1645 2788 1646
rect 2926 1650 2932 1651
rect 2926 1646 2927 1650
rect 2931 1646 2932 1650
rect 2926 1645 2932 1646
rect 3070 1650 3076 1651
rect 3070 1646 3071 1650
rect 3075 1646 3076 1650
rect 3070 1645 3076 1646
rect 3222 1650 3228 1651
rect 3222 1646 3223 1650
rect 3227 1646 3228 1650
rect 3222 1645 3228 1646
rect 3374 1650 3380 1651
rect 3374 1646 3375 1650
rect 3379 1646 3380 1650
rect 3374 1645 3380 1646
rect 3510 1650 3516 1651
rect 3510 1646 3511 1650
rect 3515 1646 3516 1650
rect 3510 1645 3516 1646
rect 110 1644 116 1645
rect 110 1640 111 1644
rect 115 1640 116 1644
rect 110 1639 116 1640
rect 1830 1644 1836 1645
rect 1830 1640 1831 1644
rect 1835 1640 1836 1644
rect 1830 1639 1836 1640
rect 1870 1632 1876 1633
rect 1870 1628 1871 1632
rect 1875 1628 1876 1632
rect 110 1627 116 1628
rect 110 1623 111 1627
rect 115 1623 116 1627
rect 1830 1627 1836 1628
rect 1870 1627 1876 1628
rect 3590 1632 3596 1633
rect 3590 1628 3591 1632
rect 3595 1628 3596 1632
rect 3590 1627 3596 1628
rect 110 1622 116 1623
rect 134 1624 140 1625
rect 134 1620 135 1624
rect 139 1620 140 1624
rect 134 1619 140 1620
rect 286 1624 292 1625
rect 286 1620 287 1624
rect 291 1620 292 1624
rect 286 1619 292 1620
rect 470 1624 476 1625
rect 470 1620 471 1624
rect 475 1620 476 1624
rect 470 1619 476 1620
rect 662 1624 668 1625
rect 662 1620 663 1624
rect 667 1620 668 1624
rect 662 1619 668 1620
rect 846 1624 852 1625
rect 846 1620 847 1624
rect 851 1620 852 1624
rect 846 1619 852 1620
rect 1022 1624 1028 1625
rect 1022 1620 1023 1624
rect 1027 1620 1028 1624
rect 1022 1619 1028 1620
rect 1190 1624 1196 1625
rect 1190 1620 1191 1624
rect 1195 1620 1196 1624
rect 1190 1619 1196 1620
rect 1350 1624 1356 1625
rect 1350 1620 1351 1624
rect 1355 1620 1356 1624
rect 1350 1619 1356 1620
rect 1510 1624 1516 1625
rect 1510 1620 1511 1624
rect 1515 1620 1516 1624
rect 1510 1619 1516 1620
rect 1670 1624 1676 1625
rect 1670 1620 1671 1624
rect 1675 1620 1676 1624
rect 1830 1623 1831 1627
rect 1835 1623 1836 1627
rect 1830 1622 1836 1623
rect 1670 1619 1676 1620
rect 1870 1615 1876 1616
rect 1870 1611 1871 1615
rect 1875 1611 1876 1615
rect 3590 1615 3596 1616
rect 1870 1610 1876 1611
rect 1958 1612 1964 1613
rect 1958 1608 1959 1612
rect 1963 1608 1964 1612
rect 1958 1607 1964 1608
rect 2078 1612 2084 1613
rect 2078 1608 2079 1612
rect 2083 1608 2084 1612
rect 2078 1607 2084 1608
rect 2206 1612 2212 1613
rect 2206 1608 2207 1612
rect 2211 1608 2212 1612
rect 2206 1607 2212 1608
rect 2342 1612 2348 1613
rect 2342 1608 2343 1612
rect 2347 1608 2348 1612
rect 2342 1607 2348 1608
rect 2486 1612 2492 1613
rect 2486 1608 2487 1612
rect 2491 1608 2492 1612
rect 2486 1607 2492 1608
rect 2630 1612 2636 1613
rect 2630 1608 2631 1612
rect 2635 1608 2636 1612
rect 2630 1607 2636 1608
rect 2774 1612 2780 1613
rect 2774 1608 2775 1612
rect 2779 1608 2780 1612
rect 2774 1607 2780 1608
rect 2918 1612 2924 1613
rect 2918 1608 2919 1612
rect 2923 1608 2924 1612
rect 2918 1607 2924 1608
rect 3062 1612 3068 1613
rect 3062 1608 3063 1612
rect 3067 1608 3068 1612
rect 3062 1607 3068 1608
rect 3214 1612 3220 1613
rect 3214 1608 3215 1612
rect 3219 1608 3220 1612
rect 3214 1607 3220 1608
rect 3366 1612 3372 1613
rect 3366 1608 3367 1612
rect 3371 1608 3372 1612
rect 3366 1607 3372 1608
rect 3502 1612 3508 1613
rect 3502 1608 3503 1612
rect 3507 1608 3508 1612
rect 3590 1611 3591 1615
rect 3595 1611 3596 1615
rect 3590 1610 3596 1611
rect 3502 1607 3508 1608
rect 158 1580 164 1581
rect 110 1577 116 1578
rect 110 1573 111 1577
rect 115 1573 116 1577
rect 158 1576 159 1580
rect 163 1576 164 1580
rect 158 1575 164 1576
rect 286 1580 292 1581
rect 286 1576 287 1580
rect 291 1576 292 1580
rect 286 1575 292 1576
rect 422 1580 428 1581
rect 422 1576 423 1580
rect 427 1576 428 1580
rect 422 1575 428 1576
rect 566 1580 572 1581
rect 566 1576 567 1580
rect 571 1576 572 1580
rect 566 1575 572 1576
rect 710 1580 716 1581
rect 710 1576 711 1580
rect 715 1576 716 1580
rect 710 1575 716 1576
rect 846 1580 852 1581
rect 846 1576 847 1580
rect 851 1576 852 1580
rect 846 1575 852 1576
rect 982 1580 988 1581
rect 982 1576 983 1580
rect 987 1576 988 1580
rect 982 1575 988 1576
rect 1118 1580 1124 1581
rect 1118 1576 1119 1580
rect 1123 1576 1124 1580
rect 1118 1575 1124 1576
rect 1246 1580 1252 1581
rect 1246 1576 1247 1580
rect 1251 1576 1252 1580
rect 1246 1575 1252 1576
rect 1374 1580 1380 1581
rect 1374 1576 1375 1580
rect 1379 1576 1380 1580
rect 1374 1575 1380 1576
rect 1510 1580 1516 1581
rect 1510 1576 1511 1580
rect 1515 1576 1516 1580
rect 1510 1575 1516 1576
rect 1830 1577 1836 1578
rect 110 1572 116 1573
rect 1830 1573 1831 1577
rect 1835 1573 1836 1577
rect 1830 1572 1836 1573
rect 110 1560 116 1561
rect 110 1556 111 1560
rect 115 1556 116 1560
rect 110 1555 116 1556
rect 1830 1560 1836 1561
rect 1830 1556 1831 1560
rect 1835 1556 1836 1560
rect 1894 1560 1900 1561
rect 1830 1555 1836 1556
rect 1870 1557 1876 1558
rect 1870 1553 1871 1557
rect 1875 1553 1876 1557
rect 1894 1556 1895 1560
rect 1899 1556 1900 1560
rect 1894 1555 1900 1556
rect 2046 1560 2052 1561
rect 2046 1556 2047 1560
rect 2051 1556 2052 1560
rect 2046 1555 2052 1556
rect 2206 1560 2212 1561
rect 2206 1556 2207 1560
rect 2211 1556 2212 1560
rect 2206 1555 2212 1556
rect 2366 1560 2372 1561
rect 2366 1556 2367 1560
rect 2371 1556 2372 1560
rect 2366 1555 2372 1556
rect 2526 1560 2532 1561
rect 2526 1556 2527 1560
rect 2531 1556 2532 1560
rect 2526 1555 2532 1556
rect 2686 1560 2692 1561
rect 2686 1556 2687 1560
rect 2691 1556 2692 1560
rect 2686 1555 2692 1556
rect 2838 1560 2844 1561
rect 2838 1556 2839 1560
rect 2843 1556 2844 1560
rect 2838 1555 2844 1556
rect 2982 1560 2988 1561
rect 2982 1556 2983 1560
rect 2987 1556 2988 1560
rect 2982 1555 2988 1556
rect 3118 1560 3124 1561
rect 3118 1556 3119 1560
rect 3123 1556 3124 1560
rect 3118 1555 3124 1556
rect 3254 1560 3260 1561
rect 3254 1556 3255 1560
rect 3259 1556 3260 1560
rect 3254 1555 3260 1556
rect 3390 1560 3396 1561
rect 3390 1556 3391 1560
rect 3395 1556 3396 1560
rect 3390 1555 3396 1556
rect 3502 1560 3508 1561
rect 3502 1556 3503 1560
rect 3507 1556 3508 1560
rect 3502 1555 3508 1556
rect 3590 1557 3596 1558
rect 1870 1552 1876 1553
rect 3590 1553 3591 1557
rect 3595 1553 3596 1557
rect 3590 1552 3596 1553
rect 166 1542 172 1543
rect 166 1538 167 1542
rect 171 1538 172 1542
rect 166 1537 172 1538
rect 294 1542 300 1543
rect 294 1538 295 1542
rect 299 1538 300 1542
rect 294 1537 300 1538
rect 430 1542 436 1543
rect 430 1538 431 1542
rect 435 1538 436 1542
rect 430 1537 436 1538
rect 574 1542 580 1543
rect 574 1538 575 1542
rect 579 1538 580 1542
rect 574 1537 580 1538
rect 718 1542 724 1543
rect 718 1538 719 1542
rect 723 1538 724 1542
rect 718 1537 724 1538
rect 854 1542 860 1543
rect 854 1538 855 1542
rect 859 1538 860 1542
rect 854 1537 860 1538
rect 990 1542 996 1543
rect 990 1538 991 1542
rect 995 1538 996 1542
rect 990 1537 996 1538
rect 1126 1542 1132 1543
rect 1126 1538 1127 1542
rect 1131 1538 1132 1542
rect 1126 1537 1132 1538
rect 1254 1542 1260 1543
rect 1254 1538 1255 1542
rect 1259 1538 1260 1542
rect 1254 1537 1260 1538
rect 1382 1542 1388 1543
rect 1382 1538 1383 1542
rect 1387 1538 1388 1542
rect 1382 1537 1388 1538
rect 1518 1542 1524 1543
rect 1518 1538 1519 1542
rect 1523 1538 1524 1542
rect 1518 1537 1524 1538
rect 1870 1540 1876 1541
rect 1870 1536 1871 1540
rect 1875 1536 1876 1540
rect 1870 1535 1876 1536
rect 3590 1540 3596 1541
rect 3590 1536 3591 1540
rect 3595 1536 3596 1540
rect 3590 1535 3596 1536
rect 1902 1522 1908 1523
rect 1902 1518 1903 1522
rect 1907 1518 1908 1522
rect 1902 1517 1908 1518
rect 2054 1522 2060 1523
rect 2054 1518 2055 1522
rect 2059 1518 2060 1522
rect 2054 1517 2060 1518
rect 2214 1522 2220 1523
rect 2214 1518 2215 1522
rect 2219 1518 2220 1522
rect 2214 1517 2220 1518
rect 2374 1522 2380 1523
rect 2374 1518 2375 1522
rect 2379 1518 2380 1522
rect 2374 1517 2380 1518
rect 2534 1522 2540 1523
rect 2534 1518 2535 1522
rect 2539 1518 2540 1522
rect 2534 1517 2540 1518
rect 2694 1522 2700 1523
rect 2694 1518 2695 1522
rect 2699 1518 2700 1522
rect 2694 1517 2700 1518
rect 2846 1522 2852 1523
rect 2846 1518 2847 1522
rect 2851 1518 2852 1522
rect 2846 1517 2852 1518
rect 2990 1522 2996 1523
rect 2990 1518 2991 1522
rect 2995 1518 2996 1522
rect 2990 1517 2996 1518
rect 3126 1522 3132 1523
rect 3126 1518 3127 1522
rect 3131 1518 3132 1522
rect 3126 1517 3132 1518
rect 3262 1522 3268 1523
rect 3262 1518 3263 1522
rect 3267 1518 3268 1522
rect 3262 1517 3268 1518
rect 3398 1522 3404 1523
rect 3398 1518 3399 1522
rect 3403 1518 3404 1522
rect 3398 1517 3404 1518
rect 3510 1522 3516 1523
rect 3510 1518 3511 1522
rect 3515 1518 3516 1522
rect 3510 1517 3516 1518
rect 230 1506 236 1507
rect 230 1502 231 1506
rect 235 1502 236 1506
rect 230 1501 236 1502
rect 374 1506 380 1507
rect 374 1502 375 1506
rect 379 1502 380 1506
rect 374 1501 380 1502
rect 518 1506 524 1507
rect 518 1502 519 1506
rect 523 1502 524 1506
rect 518 1501 524 1502
rect 654 1506 660 1507
rect 654 1502 655 1506
rect 659 1502 660 1506
rect 654 1501 660 1502
rect 782 1506 788 1507
rect 782 1502 783 1506
rect 787 1502 788 1506
rect 782 1501 788 1502
rect 902 1506 908 1507
rect 902 1502 903 1506
rect 907 1502 908 1506
rect 902 1501 908 1502
rect 1014 1506 1020 1507
rect 1014 1502 1015 1506
rect 1019 1502 1020 1506
rect 1014 1501 1020 1502
rect 1118 1506 1124 1507
rect 1118 1502 1119 1506
rect 1123 1502 1124 1506
rect 1118 1501 1124 1502
rect 1214 1506 1220 1507
rect 1214 1502 1215 1506
rect 1219 1502 1220 1506
rect 1214 1501 1220 1502
rect 1318 1506 1324 1507
rect 1318 1502 1319 1506
rect 1323 1502 1324 1506
rect 1318 1501 1324 1502
rect 1422 1506 1428 1507
rect 1422 1502 1423 1506
rect 1427 1502 1428 1506
rect 1422 1501 1428 1502
rect 110 1488 116 1489
rect 110 1484 111 1488
rect 115 1484 116 1488
rect 110 1483 116 1484
rect 1830 1488 1836 1489
rect 1830 1484 1831 1488
rect 1835 1484 1836 1488
rect 1830 1483 1836 1484
rect 1902 1482 1908 1483
rect 1902 1478 1903 1482
rect 1907 1478 1908 1482
rect 1902 1477 1908 1478
rect 2006 1482 2012 1483
rect 2006 1478 2007 1482
rect 2011 1478 2012 1482
rect 2006 1477 2012 1478
rect 2134 1482 2140 1483
rect 2134 1478 2135 1482
rect 2139 1478 2140 1482
rect 2134 1477 2140 1478
rect 2270 1482 2276 1483
rect 2270 1478 2271 1482
rect 2275 1478 2276 1482
rect 2270 1477 2276 1478
rect 2414 1482 2420 1483
rect 2414 1478 2415 1482
rect 2419 1478 2420 1482
rect 2414 1477 2420 1478
rect 2566 1482 2572 1483
rect 2566 1478 2567 1482
rect 2571 1478 2572 1482
rect 2566 1477 2572 1478
rect 2718 1482 2724 1483
rect 2718 1478 2719 1482
rect 2723 1478 2724 1482
rect 2718 1477 2724 1478
rect 2878 1482 2884 1483
rect 2878 1478 2879 1482
rect 2883 1478 2884 1482
rect 2878 1477 2884 1478
rect 3038 1482 3044 1483
rect 3038 1478 3039 1482
rect 3043 1478 3044 1482
rect 3038 1477 3044 1478
rect 3198 1482 3204 1483
rect 3198 1478 3199 1482
rect 3203 1478 3204 1482
rect 3198 1477 3204 1478
rect 3366 1482 3372 1483
rect 3366 1478 3367 1482
rect 3371 1478 3372 1482
rect 3366 1477 3372 1478
rect 3510 1482 3516 1483
rect 3510 1478 3511 1482
rect 3515 1478 3516 1482
rect 3510 1477 3516 1478
rect 110 1471 116 1472
rect 110 1467 111 1471
rect 115 1467 116 1471
rect 1830 1471 1836 1472
rect 110 1466 116 1467
rect 222 1468 228 1469
rect 222 1464 223 1468
rect 227 1464 228 1468
rect 222 1463 228 1464
rect 366 1468 372 1469
rect 366 1464 367 1468
rect 371 1464 372 1468
rect 366 1463 372 1464
rect 510 1468 516 1469
rect 510 1464 511 1468
rect 515 1464 516 1468
rect 510 1463 516 1464
rect 646 1468 652 1469
rect 646 1464 647 1468
rect 651 1464 652 1468
rect 646 1463 652 1464
rect 774 1468 780 1469
rect 774 1464 775 1468
rect 779 1464 780 1468
rect 774 1463 780 1464
rect 894 1468 900 1469
rect 894 1464 895 1468
rect 899 1464 900 1468
rect 894 1463 900 1464
rect 1006 1468 1012 1469
rect 1006 1464 1007 1468
rect 1011 1464 1012 1468
rect 1006 1463 1012 1464
rect 1110 1468 1116 1469
rect 1110 1464 1111 1468
rect 1115 1464 1116 1468
rect 1110 1463 1116 1464
rect 1206 1468 1212 1469
rect 1206 1464 1207 1468
rect 1211 1464 1212 1468
rect 1206 1463 1212 1464
rect 1310 1468 1316 1469
rect 1310 1464 1311 1468
rect 1315 1464 1316 1468
rect 1310 1463 1316 1464
rect 1414 1468 1420 1469
rect 1414 1464 1415 1468
rect 1419 1464 1420 1468
rect 1830 1467 1831 1471
rect 1835 1467 1836 1471
rect 1830 1466 1836 1467
rect 1414 1463 1420 1464
rect 1870 1464 1876 1465
rect 1870 1460 1871 1464
rect 1875 1460 1876 1464
rect 1870 1459 1876 1460
rect 3590 1464 3596 1465
rect 3590 1460 3591 1464
rect 3595 1460 3596 1464
rect 3590 1459 3596 1460
rect 1870 1447 1876 1448
rect 1870 1443 1871 1447
rect 1875 1443 1876 1447
rect 3590 1447 3596 1448
rect 1870 1442 1876 1443
rect 1894 1444 1900 1445
rect 1894 1440 1895 1444
rect 1899 1440 1900 1444
rect 1894 1439 1900 1440
rect 1998 1444 2004 1445
rect 1998 1440 1999 1444
rect 2003 1440 2004 1444
rect 1998 1439 2004 1440
rect 2126 1444 2132 1445
rect 2126 1440 2127 1444
rect 2131 1440 2132 1444
rect 2126 1439 2132 1440
rect 2262 1444 2268 1445
rect 2262 1440 2263 1444
rect 2267 1440 2268 1444
rect 2262 1439 2268 1440
rect 2406 1444 2412 1445
rect 2406 1440 2407 1444
rect 2411 1440 2412 1444
rect 2406 1439 2412 1440
rect 2558 1444 2564 1445
rect 2558 1440 2559 1444
rect 2563 1440 2564 1444
rect 2558 1439 2564 1440
rect 2710 1444 2716 1445
rect 2710 1440 2711 1444
rect 2715 1440 2716 1444
rect 2710 1439 2716 1440
rect 2870 1444 2876 1445
rect 2870 1440 2871 1444
rect 2875 1440 2876 1444
rect 2870 1439 2876 1440
rect 3030 1444 3036 1445
rect 3030 1440 3031 1444
rect 3035 1440 3036 1444
rect 3030 1439 3036 1440
rect 3190 1444 3196 1445
rect 3190 1440 3191 1444
rect 3195 1440 3196 1444
rect 3190 1439 3196 1440
rect 3358 1444 3364 1445
rect 3358 1440 3359 1444
rect 3363 1440 3364 1444
rect 3358 1439 3364 1440
rect 3502 1444 3508 1445
rect 3502 1440 3503 1444
rect 3507 1440 3508 1444
rect 3590 1443 3591 1447
rect 3595 1443 3596 1447
rect 3590 1442 3596 1443
rect 3502 1439 3508 1440
rect 254 1416 260 1417
rect 110 1413 116 1414
rect 110 1409 111 1413
rect 115 1409 116 1413
rect 254 1412 255 1416
rect 259 1412 260 1416
rect 254 1411 260 1412
rect 350 1416 356 1417
rect 350 1412 351 1416
rect 355 1412 356 1416
rect 350 1411 356 1412
rect 446 1416 452 1417
rect 446 1412 447 1416
rect 451 1412 452 1416
rect 446 1411 452 1412
rect 542 1416 548 1417
rect 542 1412 543 1416
rect 547 1412 548 1416
rect 542 1411 548 1412
rect 630 1416 636 1417
rect 630 1412 631 1416
rect 635 1412 636 1416
rect 630 1411 636 1412
rect 718 1416 724 1417
rect 718 1412 719 1416
rect 723 1412 724 1416
rect 718 1411 724 1412
rect 806 1416 812 1417
rect 806 1412 807 1416
rect 811 1412 812 1416
rect 806 1411 812 1412
rect 918 1416 924 1417
rect 918 1412 919 1416
rect 923 1412 924 1416
rect 918 1411 924 1412
rect 1046 1416 1052 1417
rect 1046 1412 1047 1416
rect 1051 1412 1052 1416
rect 1046 1411 1052 1412
rect 1206 1416 1212 1417
rect 1206 1412 1207 1416
rect 1211 1412 1212 1416
rect 1206 1411 1212 1412
rect 1382 1416 1388 1417
rect 1382 1412 1383 1416
rect 1387 1412 1388 1416
rect 1382 1411 1388 1412
rect 1574 1416 1580 1417
rect 1574 1412 1575 1416
rect 1579 1412 1580 1416
rect 1574 1411 1580 1412
rect 1742 1416 1748 1417
rect 1742 1412 1743 1416
rect 1747 1412 1748 1416
rect 1742 1411 1748 1412
rect 1830 1413 1836 1414
rect 110 1408 116 1409
rect 1830 1409 1831 1413
rect 1835 1409 1836 1413
rect 1830 1408 1836 1409
rect 1894 1400 1900 1401
rect 1870 1397 1876 1398
rect 110 1396 116 1397
rect 110 1392 111 1396
rect 115 1392 116 1396
rect 110 1391 116 1392
rect 1830 1396 1836 1397
rect 1830 1392 1831 1396
rect 1835 1392 1836 1396
rect 1870 1393 1871 1397
rect 1875 1393 1876 1397
rect 1894 1396 1895 1400
rect 1899 1396 1900 1400
rect 1894 1395 1900 1396
rect 2022 1400 2028 1401
rect 2022 1396 2023 1400
rect 2027 1396 2028 1400
rect 2022 1395 2028 1396
rect 2166 1400 2172 1401
rect 2166 1396 2167 1400
rect 2171 1396 2172 1400
rect 2166 1395 2172 1396
rect 2302 1400 2308 1401
rect 2302 1396 2303 1400
rect 2307 1396 2308 1400
rect 2302 1395 2308 1396
rect 2430 1400 2436 1401
rect 2430 1396 2431 1400
rect 2435 1396 2436 1400
rect 2430 1395 2436 1396
rect 2550 1400 2556 1401
rect 2550 1396 2551 1400
rect 2555 1396 2556 1400
rect 2550 1395 2556 1396
rect 2670 1400 2676 1401
rect 2670 1396 2671 1400
rect 2675 1396 2676 1400
rect 2670 1395 2676 1396
rect 2790 1400 2796 1401
rect 2790 1396 2791 1400
rect 2795 1396 2796 1400
rect 2790 1395 2796 1396
rect 2910 1400 2916 1401
rect 2910 1396 2911 1400
rect 2915 1396 2916 1400
rect 2910 1395 2916 1396
rect 3590 1397 3596 1398
rect 1870 1392 1876 1393
rect 3590 1393 3591 1397
rect 3595 1393 3596 1397
rect 3590 1392 3596 1393
rect 1830 1391 1836 1392
rect 1870 1380 1876 1381
rect 262 1378 268 1379
rect 262 1374 263 1378
rect 267 1374 268 1378
rect 262 1373 268 1374
rect 358 1378 364 1379
rect 358 1374 359 1378
rect 363 1374 364 1378
rect 358 1373 364 1374
rect 454 1378 460 1379
rect 454 1374 455 1378
rect 459 1374 460 1378
rect 454 1373 460 1374
rect 550 1378 556 1379
rect 550 1374 551 1378
rect 555 1374 556 1378
rect 550 1373 556 1374
rect 638 1378 644 1379
rect 638 1374 639 1378
rect 643 1374 644 1378
rect 638 1373 644 1374
rect 726 1378 732 1379
rect 726 1374 727 1378
rect 731 1374 732 1378
rect 726 1373 732 1374
rect 814 1378 820 1379
rect 814 1374 815 1378
rect 819 1374 820 1378
rect 814 1373 820 1374
rect 926 1378 932 1379
rect 926 1374 927 1378
rect 931 1374 932 1378
rect 926 1373 932 1374
rect 1054 1378 1060 1379
rect 1054 1374 1055 1378
rect 1059 1374 1060 1378
rect 1054 1373 1060 1374
rect 1214 1378 1220 1379
rect 1214 1374 1215 1378
rect 1219 1374 1220 1378
rect 1214 1373 1220 1374
rect 1390 1378 1396 1379
rect 1390 1374 1391 1378
rect 1395 1374 1396 1378
rect 1390 1373 1396 1374
rect 1582 1378 1588 1379
rect 1582 1374 1583 1378
rect 1587 1374 1588 1378
rect 1582 1373 1588 1374
rect 1750 1378 1756 1379
rect 1750 1374 1751 1378
rect 1755 1374 1756 1378
rect 1870 1376 1871 1380
rect 1875 1376 1876 1380
rect 1870 1375 1876 1376
rect 3590 1380 3596 1381
rect 3590 1376 3591 1380
rect 3595 1376 3596 1380
rect 3590 1375 3596 1376
rect 1750 1373 1756 1374
rect 1902 1362 1908 1363
rect 1902 1358 1903 1362
rect 1907 1358 1908 1362
rect 1902 1357 1908 1358
rect 2030 1362 2036 1363
rect 2030 1358 2031 1362
rect 2035 1358 2036 1362
rect 2030 1357 2036 1358
rect 2174 1362 2180 1363
rect 2174 1358 2175 1362
rect 2179 1358 2180 1362
rect 2174 1357 2180 1358
rect 2310 1362 2316 1363
rect 2310 1358 2311 1362
rect 2315 1358 2316 1362
rect 2310 1357 2316 1358
rect 2438 1362 2444 1363
rect 2438 1358 2439 1362
rect 2443 1358 2444 1362
rect 2438 1357 2444 1358
rect 2558 1362 2564 1363
rect 2558 1358 2559 1362
rect 2563 1358 2564 1362
rect 2558 1357 2564 1358
rect 2678 1362 2684 1363
rect 2678 1358 2679 1362
rect 2683 1358 2684 1362
rect 2678 1357 2684 1358
rect 2798 1362 2804 1363
rect 2798 1358 2799 1362
rect 2803 1358 2804 1362
rect 2798 1357 2804 1358
rect 2918 1362 2924 1363
rect 2918 1358 2919 1362
rect 2923 1358 2924 1362
rect 2918 1357 2924 1358
rect 358 1346 364 1347
rect 358 1342 359 1346
rect 363 1342 364 1346
rect 358 1341 364 1342
rect 470 1346 476 1347
rect 470 1342 471 1346
rect 475 1342 476 1346
rect 470 1341 476 1342
rect 590 1346 596 1347
rect 590 1342 591 1346
rect 595 1342 596 1346
rect 590 1341 596 1342
rect 726 1346 732 1347
rect 726 1342 727 1346
rect 731 1342 732 1346
rect 726 1341 732 1342
rect 862 1346 868 1347
rect 862 1342 863 1346
rect 867 1342 868 1346
rect 862 1341 868 1342
rect 1006 1346 1012 1347
rect 1006 1342 1007 1346
rect 1011 1342 1012 1346
rect 1006 1341 1012 1342
rect 1142 1346 1148 1347
rect 1142 1342 1143 1346
rect 1147 1342 1148 1346
rect 1142 1341 1148 1342
rect 1278 1346 1284 1347
rect 1278 1342 1279 1346
rect 1283 1342 1284 1346
rect 1278 1341 1284 1342
rect 1406 1346 1412 1347
rect 1406 1342 1407 1346
rect 1411 1342 1412 1346
rect 1406 1341 1412 1342
rect 1526 1346 1532 1347
rect 1526 1342 1527 1346
rect 1531 1342 1532 1346
rect 1526 1341 1532 1342
rect 1646 1346 1652 1347
rect 1646 1342 1647 1346
rect 1651 1342 1652 1346
rect 1646 1341 1652 1342
rect 1750 1346 1756 1347
rect 1750 1342 1751 1346
rect 1755 1342 1756 1346
rect 1750 1341 1756 1342
rect 110 1328 116 1329
rect 110 1324 111 1328
rect 115 1324 116 1328
rect 110 1323 116 1324
rect 1830 1328 1836 1329
rect 1830 1324 1831 1328
rect 1835 1324 1836 1328
rect 1830 1323 1836 1324
rect 1926 1322 1932 1323
rect 1926 1318 1927 1322
rect 1931 1318 1932 1322
rect 1926 1317 1932 1318
rect 2046 1322 2052 1323
rect 2046 1318 2047 1322
rect 2051 1318 2052 1322
rect 2046 1317 2052 1318
rect 2182 1322 2188 1323
rect 2182 1318 2183 1322
rect 2187 1318 2188 1322
rect 2182 1317 2188 1318
rect 2318 1322 2324 1323
rect 2318 1318 2319 1322
rect 2323 1318 2324 1322
rect 2318 1317 2324 1318
rect 2454 1322 2460 1323
rect 2454 1318 2455 1322
rect 2459 1318 2460 1322
rect 2454 1317 2460 1318
rect 2590 1322 2596 1323
rect 2590 1318 2591 1322
rect 2595 1318 2596 1322
rect 2590 1317 2596 1318
rect 2718 1322 2724 1323
rect 2718 1318 2719 1322
rect 2723 1318 2724 1322
rect 2718 1317 2724 1318
rect 2838 1322 2844 1323
rect 2838 1318 2839 1322
rect 2843 1318 2844 1322
rect 2838 1317 2844 1318
rect 2950 1322 2956 1323
rect 2950 1318 2951 1322
rect 2955 1318 2956 1322
rect 2950 1317 2956 1318
rect 3062 1322 3068 1323
rect 3062 1318 3063 1322
rect 3067 1318 3068 1322
rect 3062 1317 3068 1318
rect 3182 1322 3188 1323
rect 3182 1318 3183 1322
rect 3187 1318 3188 1322
rect 3182 1317 3188 1318
rect 110 1311 116 1312
rect 110 1307 111 1311
rect 115 1307 116 1311
rect 1830 1311 1836 1312
rect 110 1306 116 1307
rect 350 1308 356 1309
rect 350 1304 351 1308
rect 355 1304 356 1308
rect 350 1303 356 1304
rect 462 1308 468 1309
rect 462 1304 463 1308
rect 467 1304 468 1308
rect 462 1303 468 1304
rect 582 1308 588 1309
rect 582 1304 583 1308
rect 587 1304 588 1308
rect 582 1303 588 1304
rect 718 1308 724 1309
rect 718 1304 719 1308
rect 723 1304 724 1308
rect 718 1303 724 1304
rect 854 1308 860 1309
rect 854 1304 855 1308
rect 859 1304 860 1308
rect 854 1303 860 1304
rect 998 1308 1004 1309
rect 998 1304 999 1308
rect 1003 1304 1004 1308
rect 998 1303 1004 1304
rect 1134 1308 1140 1309
rect 1134 1304 1135 1308
rect 1139 1304 1140 1308
rect 1134 1303 1140 1304
rect 1270 1308 1276 1309
rect 1270 1304 1271 1308
rect 1275 1304 1276 1308
rect 1270 1303 1276 1304
rect 1398 1308 1404 1309
rect 1398 1304 1399 1308
rect 1403 1304 1404 1308
rect 1398 1303 1404 1304
rect 1518 1308 1524 1309
rect 1518 1304 1519 1308
rect 1523 1304 1524 1308
rect 1518 1303 1524 1304
rect 1638 1308 1644 1309
rect 1638 1304 1639 1308
rect 1643 1304 1644 1308
rect 1638 1303 1644 1304
rect 1742 1308 1748 1309
rect 1742 1304 1743 1308
rect 1747 1304 1748 1308
rect 1830 1307 1831 1311
rect 1835 1307 1836 1311
rect 1830 1306 1836 1307
rect 1742 1303 1748 1304
rect 1870 1304 1876 1305
rect 1870 1300 1871 1304
rect 1875 1300 1876 1304
rect 1870 1299 1876 1300
rect 3590 1304 3596 1305
rect 3590 1300 3591 1304
rect 3595 1300 3596 1304
rect 3590 1299 3596 1300
rect 1870 1287 1876 1288
rect 1870 1283 1871 1287
rect 1875 1283 1876 1287
rect 3590 1287 3596 1288
rect 1870 1282 1876 1283
rect 1918 1284 1924 1285
rect 1918 1280 1919 1284
rect 1923 1280 1924 1284
rect 1918 1279 1924 1280
rect 2038 1284 2044 1285
rect 2038 1280 2039 1284
rect 2043 1280 2044 1284
rect 2038 1279 2044 1280
rect 2174 1284 2180 1285
rect 2174 1280 2175 1284
rect 2179 1280 2180 1284
rect 2174 1279 2180 1280
rect 2310 1284 2316 1285
rect 2310 1280 2311 1284
rect 2315 1280 2316 1284
rect 2310 1279 2316 1280
rect 2446 1284 2452 1285
rect 2446 1280 2447 1284
rect 2451 1280 2452 1284
rect 2446 1279 2452 1280
rect 2582 1284 2588 1285
rect 2582 1280 2583 1284
rect 2587 1280 2588 1284
rect 2582 1279 2588 1280
rect 2710 1284 2716 1285
rect 2710 1280 2711 1284
rect 2715 1280 2716 1284
rect 2710 1279 2716 1280
rect 2830 1284 2836 1285
rect 2830 1280 2831 1284
rect 2835 1280 2836 1284
rect 2830 1279 2836 1280
rect 2942 1284 2948 1285
rect 2942 1280 2943 1284
rect 2947 1280 2948 1284
rect 2942 1279 2948 1280
rect 3054 1284 3060 1285
rect 3054 1280 3055 1284
rect 3059 1280 3060 1284
rect 3054 1279 3060 1280
rect 3174 1284 3180 1285
rect 3174 1280 3175 1284
rect 3179 1280 3180 1284
rect 3590 1283 3591 1287
rect 3595 1283 3596 1287
rect 3590 1282 3596 1283
rect 3174 1279 3180 1280
rect 310 1260 316 1261
rect 110 1257 116 1258
rect 110 1253 111 1257
rect 115 1253 116 1257
rect 310 1256 311 1260
rect 315 1256 316 1260
rect 310 1255 316 1256
rect 414 1260 420 1261
rect 414 1256 415 1260
rect 419 1256 420 1260
rect 414 1255 420 1256
rect 534 1260 540 1261
rect 534 1256 535 1260
rect 539 1256 540 1260
rect 534 1255 540 1256
rect 670 1260 676 1261
rect 670 1256 671 1260
rect 675 1256 676 1260
rect 670 1255 676 1256
rect 814 1260 820 1261
rect 814 1256 815 1260
rect 819 1256 820 1260
rect 814 1255 820 1256
rect 958 1260 964 1261
rect 958 1256 959 1260
rect 963 1256 964 1260
rect 958 1255 964 1256
rect 1102 1260 1108 1261
rect 1102 1256 1103 1260
rect 1107 1256 1108 1260
rect 1102 1255 1108 1256
rect 1238 1260 1244 1261
rect 1238 1256 1239 1260
rect 1243 1256 1244 1260
rect 1238 1255 1244 1256
rect 1374 1260 1380 1261
rect 1374 1256 1375 1260
rect 1379 1256 1380 1260
rect 1374 1255 1380 1256
rect 1502 1260 1508 1261
rect 1502 1256 1503 1260
rect 1507 1256 1508 1260
rect 1502 1255 1508 1256
rect 1630 1260 1636 1261
rect 1630 1256 1631 1260
rect 1635 1256 1636 1260
rect 1630 1255 1636 1256
rect 1742 1260 1748 1261
rect 1742 1256 1743 1260
rect 1747 1256 1748 1260
rect 1742 1255 1748 1256
rect 1830 1257 1836 1258
rect 110 1252 116 1253
rect 1830 1253 1831 1257
rect 1835 1253 1836 1257
rect 1830 1252 1836 1253
rect 110 1240 116 1241
rect 110 1236 111 1240
rect 115 1236 116 1240
rect 110 1235 116 1236
rect 1830 1240 1836 1241
rect 1830 1236 1831 1240
rect 1835 1236 1836 1240
rect 1830 1235 1836 1236
rect 1894 1232 1900 1233
rect 1870 1229 1876 1230
rect 1870 1225 1871 1229
rect 1875 1225 1876 1229
rect 1894 1228 1895 1232
rect 1899 1228 1900 1232
rect 1894 1227 1900 1228
rect 2070 1232 2076 1233
rect 2070 1228 2071 1232
rect 2075 1228 2076 1232
rect 2070 1227 2076 1228
rect 2270 1232 2276 1233
rect 2270 1228 2271 1232
rect 2275 1228 2276 1232
rect 2270 1227 2276 1228
rect 2470 1232 2476 1233
rect 2470 1228 2471 1232
rect 2475 1228 2476 1232
rect 2470 1227 2476 1228
rect 2662 1232 2668 1233
rect 2662 1228 2663 1232
rect 2667 1228 2668 1232
rect 2662 1227 2668 1228
rect 2846 1232 2852 1233
rect 2846 1228 2847 1232
rect 2851 1228 2852 1232
rect 2846 1227 2852 1228
rect 3022 1232 3028 1233
rect 3022 1228 3023 1232
rect 3027 1228 3028 1232
rect 3022 1227 3028 1228
rect 3190 1232 3196 1233
rect 3190 1228 3191 1232
rect 3195 1228 3196 1232
rect 3190 1227 3196 1228
rect 3358 1232 3364 1233
rect 3358 1228 3359 1232
rect 3363 1228 3364 1232
rect 3358 1227 3364 1228
rect 3502 1232 3508 1233
rect 3502 1228 3503 1232
rect 3507 1228 3508 1232
rect 3502 1227 3508 1228
rect 3590 1229 3596 1230
rect 1870 1224 1876 1225
rect 3590 1225 3591 1229
rect 3595 1225 3596 1229
rect 3590 1224 3596 1225
rect 318 1222 324 1223
rect 318 1218 319 1222
rect 323 1218 324 1222
rect 318 1217 324 1218
rect 422 1222 428 1223
rect 422 1218 423 1222
rect 427 1218 428 1222
rect 422 1217 428 1218
rect 542 1222 548 1223
rect 542 1218 543 1222
rect 547 1218 548 1222
rect 542 1217 548 1218
rect 678 1222 684 1223
rect 678 1218 679 1222
rect 683 1218 684 1222
rect 678 1217 684 1218
rect 822 1222 828 1223
rect 822 1218 823 1222
rect 827 1218 828 1222
rect 822 1217 828 1218
rect 966 1222 972 1223
rect 966 1218 967 1222
rect 971 1218 972 1222
rect 966 1217 972 1218
rect 1110 1222 1116 1223
rect 1110 1218 1111 1222
rect 1115 1218 1116 1222
rect 1110 1217 1116 1218
rect 1246 1222 1252 1223
rect 1246 1218 1247 1222
rect 1251 1218 1252 1222
rect 1246 1217 1252 1218
rect 1382 1222 1388 1223
rect 1382 1218 1383 1222
rect 1387 1218 1388 1222
rect 1382 1217 1388 1218
rect 1510 1222 1516 1223
rect 1510 1218 1511 1222
rect 1515 1218 1516 1222
rect 1510 1217 1516 1218
rect 1638 1222 1644 1223
rect 1638 1218 1639 1222
rect 1643 1218 1644 1222
rect 1638 1217 1644 1218
rect 1750 1222 1756 1223
rect 1750 1218 1751 1222
rect 1755 1218 1756 1222
rect 1750 1217 1756 1218
rect 1870 1212 1876 1213
rect 1870 1208 1871 1212
rect 1875 1208 1876 1212
rect 1870 1207 1876 1208
rect 3590 1212 3596 1213
rect 3590 1208 3591 1212
rect 3595 1208 3596 1212
rect 3590 1207 3596 1208
rect 1902 1194 1908 1195
rect 238 1190 244 1191
rect 238 1186 239 1190
rect 243 1186 244 1190
rect 238 1185 244 1186
rect 414 1190 420 1191
rect 414 1186 415 1190
rect 419 1186 420 1190
rect 414 1185 420 1186
rect 590 1190 596 1191
rect 590 1186 591 1190
rect 595 1186 596 1190
rect 590 1185 596 1186
rect 758 1190 764 1191
rect 758 1186 759 1190
rect 763 1186 764 1190
rect 758 1185 764 1186
rect 926 1190 932 1191
rect 926 1186 927 1190
rect 931 1186 932 1190
rect 926 1185 932 1186
rect 1078 1190 1084 1191
rect 1078 1186 1079 1190
rect 1083 1186 1084 1190
rect 1078 1185 1084 1186
rect 1222 1190 1228 1191
rect 1222 1186 1223 1190
rect 1227 1186 1228 1190
rect 1222 1185 1228 1186
rect 1366 1190 1372 1191
rect 1366 1186 1367 1190
rect 1371 1186 1372 1190
rect 1366 1185 1372 1186
rect 1502 1190 1508 1191
rect 1502 1186 1503 1190
rect 1507 1186 1508 1190
rect 1502 1185 1508 1186
rect 1638 1190 1644 1191
rect 1638 1186 1639 1190
rect 1643 1186 1644 1190
rect 1638 1185 1644 1186
rect 1750 1190 1756 1191
rect 1750 1186 1751 1190
rect 1755 1186 1756 1190
rect 1902 1190 1903 1194
rect 1907 1190 1908 1194
rect 1902 1189 1908 1190
rect 2078 1194 2084 1195
rect 2078 1190 2079 1194
rect 2083 1190 2084 1194
rect 2078 1189 2084 1190
rect 2278 1194 2284 1195
rect 2278 1190 2279 1194
rect 2283 1190 2284 1194
rect 2278 1189 2284 1190
rect 2478 1194 2484 1195
rect 2478 1190 2479 1194
rect 2483 1190 2484 1194
rect 2478 1189 2484 1190
rect 2670 1194 2676 1195
rect 2670 1190 2671 1194
rect 2675 1190 2676 1194
rect 2670 1189 2676 1190
rect 2854 1194 2860 1195
rect 2854 1190 2855 1194
rect 2859 1190 2860 1194
rect 2854 1189 2860 1190
rect 3030 1194 3036 1195
rect 3030 1190 3031 1194
rect 3035 1190 3036 1194
rect 3030 1189 3036 1190
rect 3198 1194 3204 1195
rect 3198 1190 3199 1194
rect 3203 1190 3204 1194
rect 3198 1189 3204 1190
rect 3366 1194 3372 1195
rect 3366 1190 3367 1194
rect 3371 1190 3372 1194
rect 3366 1189 3372 1190
rect 3510 1194 3516 1195
rect 3510 1190 3511 1194
rect 3515 1190 3516 1194
rect 3510 1189 3516 1190
rect 1750 1185 1756 1186
rect 110 1172 116 1173
rect 110 1168 111 1172
rect 115 1168 116 1172
rect 110 1167 116 1168
rect 1830 1172 1836 1173
rect 1830 1168 1831 1172
rect 1835 1168 1836 1172
rect 1830 1167 1836 1168
rect 1902 1158 1908 1159
rect 110 1155 116 1156
rect 110 1151 111 1155
rect 115 1151 116 1155
rect 1830 1155 1836 1156
rect 110 1150 116 1151
rect 230 1152 236 1153
rect 230 1148 231 1152
rect 235 1148 236 1152
rect 230 1147 236 1148
rect 406 1152 412 1153
rect 406 1148 407 1152
rect 411 1148 412 1152
rect 406 1147 412 1148
rect 582 1152 588 1153
rect 582 1148 583 1152
rect 587 1148 588 1152
rect 582 1147 588 1148
rect 750 1152 756 1153
rect 750 1148 751 1152
rect 755 1148 756 1152
rect 750 1147 756 1148
rect 918 1152 924 1153
rect 918 1148 919 1152
rect 923 1148 924 1152
rect 918 1147 924 1148
rect 1070 1152 1076 1153
rect 1070 1148 1071 1152
rect 1075 1148 1076 1152
rect 1070 1147 1076 1148
rect 1214 1152 1220 1153
rect 1214 1148 1215 1152
rect 1219 1148 1220 1152
rect 1214 1147 1220 1148
rect 1358 1152 1364 1153
rect 1358 1148 1359 1152
rect 1363 1148 1364 1152
rect 1358 1147 1364 1148
rect 1494 1152 1500 1153
rect 1494 1148 1495 1152
rect 1499 1148 1500 1152
rect 1494 1147 1500 1148
rect 1630 1152 1636 1153
rect 1630 1148 1631 1152
rect 1635 1148 1636 1152
rect 1630 1147 1636 1148
rect 1742 1152 1748 1153
rect 1742 1148 1743 1152
rect 1747 1148 1748 1152
rect 1830 1151 1831 1155
rect 1835 1151 1836 1155
rect 1902 1154 1903 1158
rect 1907 1154 1908 1158
rect 1902 1153 1908 1154
rect 1982 1158 1988 1159
rect 1982 1154 1983 1158
rect 1987 1154 1988 1158
rect 1982 1153 1988 1154
rect 2086 1158 2092 1159
rect 2086 1154 2087 1158
rect 2091 1154 2092 1158
rect 2086 1153 2092 1154
rect 2214 1158 2220 1159
rect 2214 1154 2215 1158
rect 2219 1154 2220 1158
rect 2214 1153 2220 1154
rect 2366 1158 2372 1159
rect 2366 1154 2367 1158
rect 2371 1154 2372 1158
rect 2366 1153 2372 1154
rect 2526 1158 2532 1159
rect 2526 1154 2527 1158
rect 2531 1154 2532 1158
rect 2526 1153 2532 1154
rect 2686 1158 2692 1159
rect 2686 1154 2687 1158
rect 2691 1154 2692 1158
rect 2686 1153 2692 1154
rect 2838 1158 2844 1159
rect 2838 1154 2839 1158
rect 2843 1154 2844 1158
rect 2838 1153 2844 1154
rect 2982 1158 2988 1159
rect 2982 1154 2983 1158
rect 2987 1154 2988 1158
rect 2982 1153 2988 1154
rect 3126 1158 3132 1159
rect 3126 1154 3127 1158
rect 3131 1154 3132 1158
rect 3126 1153 3132 1154
rect 3262 1158 3268 1159
rect 3262 1154 3263 1158
rect 3267 1154 3268 1158
rect 3262 1153 3268 1154
rect 3398 1158 3404 1159
rect 3398 1154 3399 1158
rect 3403 1154 3404 1158
rect 3398 1153 3404 1154
rect 3510 1158 3516 1159
rect 3510 1154 3511 1158
rect 3515 1154 3516 1158
rect 3510 1153 3516 1154
rect 1830 1150 1836 1151
rect 1742 1147 1748 1148
rect 1870 1140 1876 1141
rect 1870 1136 1871 1140
rect 1875 1136 1876 1140
rect 1870 1135 1876 1136
rect 3590 1140 3596 1141
rect 3590 1136 3591 1140
rect 3595 1136 3596 1140
rect 3590 1135 3596 1136
rect 1870 1123 1876 1124
rect 1870 1119 1871 1123
rect 1875 1119 1876 1123
rect 3590 1123 3596 1124
rect 1870 1118 1876 1119
rect 1894 1120 1900 1121
rect 1894 1116 1895 1120
rect 1899 1116 1900 1120
rect 1894 1115 1900 1116
rect 1974 1120 1980 1121
rect 1974 1116 1975 1120
rect 1979 1116 1980 1120
rect 1974 1115 1980 1116
rect 2078 1120 2084 1121
rect 2078 1116 2079 1120
rect 2083 1116 2084 1120
rect 2078 1115 2084 1116
rect 2206 1120 2212 1121
rect 2206 1116 2207 1120
rect 2211 1116 2212 1120
rect 2206 1115 2212 1116
rect 2358 1120 2364 1121
rect 2358 1116 2359 1120
rect 2363 1116 2364 1120
rect 2358 1115 2364 1116
rect 2518 1120 2524 1121
rect 2518 1116 2519 1120
rect 2523 1116 2524 1120
rect 2518 1115 2524 1116
rect 2678 1120 2684 1121
rect 2678 1116 2679 1120
rect 2683 1116 2684 1120
rect 2678 1115 2684 1116
rect 2830 1120 2836 1121
rect 2830 1116 2831 1120
rect 2835 1116 2836 1120
rect 2830 1115 2836 1116
rect 2974 1120 2980 1121
rect 2974 1116 2975 1120
rect 2979 1116 2980 1120
rect 2974 1115 2980 1116
rect 3118 1120 3124 1121
rect 3118 1116 3119 1120
rect 3123 1116 3124 1120
rect 3118 1115 3124 1116
rect 3254 1120 3260 1121
rect 3254 1116 3255 1120
rect 3259 1116 3260 1120
rect 3254 1115 3260 1116
rect 3390 1120 3396 1121
rect 3390 1116 3391 1120
rect 3395 1116 3396 1120
rect 3390 1115 3396 1116
rect 3502 1120 3508 1121
rect 3502 1116 3503 1120
rect 3507 1116 3508 1120
rect 3590 1119 3591 1123
rect 3595 1119 3596 1123
rect 3590 1118 3596 1119
rect 3502 1115 3508 1116
rect 142 1104 148 1105
rect 110 1101 116 1102
rect 110 1097 111 1101
rect 115 1097 116 1101
rect 142 1100 143 1104
rect 147 1100 148 1104
rect 142 1099 148 1100
rect 278 1104 284 1105
rect 278 1100 279 1104
rect 283 1100 284 1104
rect 278 1099 284 1100
rect 422 1104 428 1105
rect 422 1100 423 1104
rect 427 1100 428 1104
rect 422 1099 428 1100
rect 566 1104 572 1105
rect 566 1100 567 1104
rect 571 1100 572 1104
rect 566 1099 572 1100
rect 710 1104 716 1105
rect 710 1100 711 1104
rect 715 1100 716 1104
rect 710 1099 716 1100
rect 846 1104 852 1105
rect 846 1100 847 1104
rect 851 1100 852 1104
rect 846 1099 852 1100
rect 974 1104 980 1105
rect 974 1100 975 1104
rect 979 1100 980 1104
rect 974 1099 980 1100
rect 1102 1104 1108 1105
rect 1102 1100 1103 1104
rect 1107 1100 1108 1104
rect 1102 1099 1108 1100
rect 1222 1104 1228 1105
rect 1222 1100 1223 1104
rect 1227 1100 1228 1104
rect 1222 1099 1228 1100
rect 1342 1104 1348 1105
rect 1342 1100 1343 1104
rect 1347 1100 1348 1104
rect 1342 1099 1348 1100
rect 1470 1104 1476 1105
rect 1470 1100 1471 1104
rect 1475 1100 1476 1104
rect 1470 1099 1476 1100
rect 1830 1101 1836 1102
rect 110 1096 116 1097
rect 1830 1097 1831 1101
rect 1835 1097 1836 1101
rect 1830 1096 1836 1097
rect 110 1084 116 1085
rect 110 1080 111 1084
rect 115 1080 116 1084
rect 110 1079 116 1080
rect 1830 1084 1836 1085
rect 1830 1080 1831 1084
rect 1835 1080 1836 1084
rect 1830 1079 1836 1080
rect 2166 1068 2172 1069
rect 150 1066 156 1067
rect 150 1062 151 1066
rect 155 1062 156 1066
rect 150 1061 156 1062
rect 286 1066 292 1067
rect 286 1062 287 1066
rect 291 1062 292 1066
rect 286 1061 292 1062
rect 430 1066 436 1067
rect 430 1062 431 1066
rect 435 1062 436 1066
rect 430 1061 436 1062
rect 574 1066 580 1067
rect 574 1062 575 1066
rect 579 1062 580 1066
rect 574 1061 580 1062
rect 718 1066 724 1067
rect 718 1062 719 1066
rect 723 1062 724 1066
rect 718 1061 724 1062
rect 854 1066 860 1067
rect 854 1062 855 1066
rect 859 1062 860 1066
rect 854 1061 860 1062
rect 982 1066 988 1067
rect 982 1062 983 1066
rect 987 1062 988 1066
rect 982 1061 988 1062
rect 1110 1066 1116 1067
rect 1110 1062 1111 1066
rect 1115 1062 1116 1066
rect 1110 1061 1116 1062
rect 1230 1066 1236 1067
rect 1230 1062 1231 1066
rect 1235 1062 1236 1066
rect 1230 1061 1236 1062
rect 1350 1066 1356 1067
rect 1350 1062 1351 1066
rect 1355 1062 1356 1066
rect 1350 1061 1356 1062
rect 1478 1066 1484 1067
rect 1478 1062 1479 1066
rect 1483 1062 1484 1066
rect 1478 1061 1484 1062
rect 1870 1065 1876 1066
rect 1870 1061 1871 1065
rect 1875 1061 1876 1065
rect 2166 1064 2167 1068
rect 2171 1064 2172 1068
rect 2166 1063 2172 1064
rect 2254 1068 2260 1069
rect 2254 1064 2255 1068
rect 2259 1064 2260 1068
rect 2254 1063 2260 1064
rect 2358 1068 2364 1069
rect 2358 1064 2359 1068
rect 2363 1064 2364 1068
rect 2358 1063 2364 1064
rect 2478 1068 2484 1069
rect 2478 1064 2479 1068
rect 2483 1064 2484 1068
rect 2478 1063 2484 1064
rect 2606 1068 2612 1069
rect 2606 1064 2607 1068
rect 2611 1064 2612 1068
rect 2606 1063 2612 1064
rect 2750 1068 2756 1069
rect 2750 1064 2751 1068
rect 2755 1064 2756 1068
rect 2750 1063 2756 1064
rect 2894 1068 2900 1069
rect 2894 1064 2895 1068
rect 2899 1064 2900 1068
rect 2894 1063 2900 1064
rect 3046 1068 3052 1069
rect 3046 1064 3047 1068
rect 3051 1064 3052 1068
rect 3046 1063 3052 1064
rect 3206 1068 3212 1069
rect 3206 1064 3207 1068
rect 3211 1064 3212 1068
rect 3206 1063 3212 1064
rect 3366 1068 3372 1069
rect 3366 1064 3367 1068
rect 3371 1064 3372 1068
rect 3366 1063 3372 1064
rect 3502 1068 3508 1069
rect 3502 1064 3503 1068
rect 3507 1064 3508 1068
rect 3502 1063 3508 1064
rect 3590 1065 3596 1066
rect 1870 1060 1876 1061
rect 3590 1061 3591 1065
rect 3595 1061 3596 1065
rect 3590 1060 3596 1061
rect 1870 1048 1876 1049
rect 1870 1044 1871 1048
rect 1875 1044 1876 1048
rect 1870 1043 1876 1044
rect 3590 1048 3596 1049
rect 3590 1044 3591 1048
rect 3595 1044 3596 1048
rect 3590 1043 3596 1044
rect 2174 1030 2180 1031
rect 142 1026 148 1027
rect 142 1022 143 1026
rect 147 1022 148 1026
rect 142 1021 148 1022
rect 262 1026 268 1027
rect 262 1022 263 1026
rect 267 1022 268 1026
rect 262 1021 268 1022
rect 406 1026 412 1027
rect 406 1022 407 1026
rect 411 1022 412 1026
rect 406 1021 412 1022
rect 550 1026 556 1027
rect 550 1022 551 1026
rect 555 1022 556 1026
rect 550 1021 556 1022
rect 686 1026 692 1027
rect 686 1022 687 1026
rect 691 1022 692 1026
rect 686 1021 692 1022
rect 806 1026 812 1027
rect 806 1022 807 1026
rect 811 1022 812 1026
rect 806 1021 812 1022
rect 926 1026 932 1027
rect 926 1022 927 1026
rect 931 1022 932 1026
rect 926 1021 932 1022
rect 1038 1026 1044 1027
rect 1038 1022 1039 1026
rect 1043 1022 1044 1026
rect 1038 1021 1044 1022
rect 1142 1026 1148 1027
rect 1142 1022 1143 1026
rect 1147 1022 1148 1026
rect 1142 1021 1148 1022
rect 1246 1026 1252 1027
rect 1246 1022 1247 1026
rect 1251 1022 1252 1026
rect 1246 1021 1252 1022
rect 1358 1026 1364 1027
rect 1358 1022 1359 1026
rect 1363 1022 1364 1026
rect 2174 1026 2175 1030
rect 2179 1026 2180 1030
rect 2174 1025 2180 1026
rect 2262 1030 2268 1031
rect 2262 1026 2263 1030
rect 2267 1026 2268 1030
rect 2262 1025 2268 1026
rect 2366 1030 2372 1031
rect 2366 1026 2367 1030
rect 2371 1026 2372 1030
rect 2366 1025 2372 1026
rect 2486 1030 2492 1031
rect 2486 1026 2487 1030
rect 2491 1026 2492 1030
rect 2486 1025 2492 1026
rect 2614 1030 2620 1031
rect 2614 1026 2615 1030
rect 2619 1026 2620 1030
rect 2614 1025 2620 1026
rect 2758 1030 2764 1031
rect 2758 1026 2759 1030
rect 2763 1026 2764 1030
rect 2758 1025 2764 1026
rect 2902 1030 2908 1031
rect 2902 1026 2903 1030
rect 2907 1026 2908 1030
rect 2902 1025 2908 1026
rect 3054 1030 3060 1031
rect 3054 1026 3055 1030
rect 3059 1026 3060 1030
rect 3054 1025 3060 1026
rect 3214 1030 3220 1031
rect 3214 1026 3215 1030
rect 3219 1026 3220 1030
rect 3214 1025 3220 1026
rect 3374 1030 3380 1031
rect 3374 1026 3375 1030
rect 3379 1026 3380 1030
rect 3374 1025 3380 1026
rect 3510 1030 3516 1031
rect 3510 1026 3511 1030
rect 3515 1026 3516 1030
rect 3510 1025 3516 1026
rect 1358 1021 1364 1022
rect 110 1008 116 1009
rect 110 1004 111 1008
rect 115 1004 116 1008
rect 110 1003 116 1004
rect 1830 1008 1836 1009
rect 1830 1004 1831 1008
rect 1835 1004 1836 1008
rect 1830 1003 1836 1004
rect 2302 998 2308 999
rect 2302 994 2303 998
rect 2307 994 2308 998
rect 2302 993 2308 994
rect 2382 998 2388 999
rect 2382 994 2383 998
rect 2387 994 2388 998
rect 2382 993 2388 994
rect 2470 998 2476 999
rect 2470 994 2471 998
rect 2475 994 2476 998
rect 2470 993 2476 994
rect 2566 998 2572 999
rect 2566 994 2567 998
rect 2571 994 2572 998
rect 2566 993 2572 994
rect 2670 998 2676 999
rect 2670 994 2671 998
rect 2675 994 2676 998
rect 2670 993 2676 994
rect 2782 998 2788 999
rect 2782 994 2783 998
rect 2787 994 2788 998
rect 2782 993 2788 994
rect 2910 998 2916 999
rect 2910 994 2911 998
rect 2915 994 2916 998
rect 2910 993 2916 994
rect 3054 998 3060 999
rect 3054 994 3055 998
rect 3059 994 3060 998
rect 3054 993 3060 994
rect 3206 998 3212 999
rect 3206 994 3207 998
rect 3211 994 3212 998
rect 3206 993 3212 994
rect 3366 998 3372 999
rect 3366 994 3367 998
rect 3371 994 3372 998
rect 3366 993 3372 994
rect 3510 998 3516 999
rect 3510 994 3511 998
rect 3515 994 3516 998
rect 3510 993 3516 994
rect 110 991 116 992
rect 110 987 111 991
rect 115 987 116 991
rect 1830 991 1836 992
rect 110 986 116 987
rect 134 988 140 989
rect 134 984 135 988
rect 139 984 140 988
rect 134 983 140 984
rect 254 988 260 989
rect 254 984 255 988
rect 259 984 260 988
rect 254 983 260 984
rect 398 988 404 989
rect 398 984 399 988
rect 403 984 404 988
rect 398 983 404 984
rect 542 988 548 989
rect 542 984 543 988
rect 547 984 548 988
rect 542 983 548 984
rect 678 988 684 989
rect 678 984 679 988
rect 683 984 684 988
rect 678 983 684 984
rect 798 988 804 989
rect 798 984 799 988
rect 803 984 804 988
rect 798 983 804 984
rect 918 988 924 989
rect 918 984 919 988
rect 923 984 924 988
rect 918 983 924 984
rect 1030 988 1036 989
rect 1030 984 1031 988
rect 1035 984 1036 988
rect 1030 983 1036 984
rect 1134 988 1140 989
rect 1134 984 1135 988
rect 1139 984 1140 988
rect 1134 983 1140 984
rect 1238 988 1244 989
rect 1238 984 1239 988
rect 1243 984 1244 988
rect 1238 983 1244 984
rect 1350 988 1356 989
rect 1350 984 1351 988
rect 1355 984 1356 988
rect 1830 987 1831 991
rect 1835 987 1836 991
rect 1830 986 1836 987
rect 1350 983 1356 984
rect 1870 980 1876 981
rect 1870 976 1871 980
rect 1875 976 1876 980
rect 1870 975 1876 976
rect 3590 980 3596 981
rect 3590 976 3591 980
rect 3595 976 3596 980
rect 3590 975 3596 976
rect 1870 963 1876 964
rect 1870 959 1871 963
rect 1875 959 1876 963
rect 3590 963 3596 964
rect 1870 958 1876 959
rect 2294 960 2300 961
rect 2294 956 2295 960
rect 2299 956 2300 960
rect 2294 955 2300 956
rect 2374 960 2380 961
rect 2374 956 2375 960
rect 2379 956 2380 960
rect 2374 955 2380 956
rect 2462 960 2468 961
rect 2462 956 2463 960
rect 2467 956 2468 960
rect 2462 955 2468 956
rect 2558 960 2564 961
rect 2558 956 2559 960
rect 2563 956 2564 960
rect 2558 955 2564 956
rect 2662 960 2668 961
rect 2662 956 2663 960
rect 2667 956 2668 960
rect 2662 955 2668 956
rect 2774 960 2780 961
rect 2774 956 2775 960
rect 2779 956 2780 960
rect 2774 955 2780 956
rect 2902 960 2908 961
rect 2902 956 2903 960
rect 2907 956 2908 960
rect 2902 955 2908 956
rect 3046 960 3052 961
rect 3046 956 3047 960
rect 3051 956 3052 960
rect 3046 955 3052 956
rect 3198 960 3204 961
rect 3198 956 3199 960
rect 3203 956 3204 960
rect 3198 955 3204 956
rect 3358 960 3364 961
rect 3358 956 3359 960
rect 3363 956 3364 960
rect 3358 955 3364 956
rect 3502 960 3508 961
rect 3502 956 3503 960
rect 3507 956 3508 960
rect 3590 959 3591 963
rect 3595 959 3596 963
rect 3590 958 3596 959
rect 3502 955 3508 956
rect 134 936 140 937
rect 110 933 116 934
rect 110 929 111 933
rect 115 929 116 933
rect 134 932 135 936
rect 139 932 140 936
rect 134 931 140 932
rect 214 936 220 937
rect 214 932 215 936
rect 219 932 220 936
rect 214 931 220 932
rect 326 936 332 937
rect 326 932 327 936
rect 331 932 332 936
rect 326 931 332 932
rect 446 936 452 937
rect 446 932 447 936
rect 451 932 452 936
rect 446 931 452 932
rect 566 936 572 937
rect 566 932 567 936
rect 571 932 572 936
rect 566 931 572 932
rect 686 936 692 937
rect 686 932 687 936
rect 691 932 692 936
rect 686 931 692 932
rect 798 936 804 937
rect 798 932 799 936
rect 803 932 804 936
rect 798 931 804 932
rect 910 936 916 937
rect 910 932 911 936
rect 915 932 916 936
rect 910 931 916 932
rect 1014 936 1020 937
rect 1014 932 1015 936
rect 1019 932 1020 936
rect 1014 931 1020 932
rect 1118 936 1124 937
rect 1118 932 1119 936
rect 1123 932 1124 936
rect 1118 931 1124 932
rect 1222 936 1228 937
rect 1222 932 1223 936
rect 1227 932 1228 936
rect 1222 931 1228 932
rect 1326 936 1332 937
rect 1326 932 1327 936
rect 1331 932 1332 936
rect 1326 931 1332 932
rect 1830 933 1836 934
rect 110 928 116 929
rect 1830 929 1831 933
rect 1835 929 1836 933
rect 1830 928 1836 929
rect 110 916 116 917
rect 110 912 111 916
rect 115 912 116 916
rect 110 911 116 912
rect 1830 916 1836 917
rect 1830 912 1831 916
rect 1835 912 1836 916
rect 1830 911 1836 912
rect 2278 908 2284 909
rect 1870 905 1876 906
rect 1870 901 1871 905
rect 1875 901 1876 905
rect 2278 904 2279 908
rect 2283 904 2284 908
rect 2278 903 2284 904
rect 2358 908 2364 909
rect 2358 904 2359 908
rect 2363 904 2364 908
rect 2358 903 2364 904
rect 2438 908 2444 909
rect 2438 904 2439 908
rect 2443 904 2444 908
rect 2438 903 2444 904
rect 2518 908 2524 909
rect 2518 904 2519 908
rect 2523 904 2524 908
rect 2518 903 2524 904
rect 2606 908 2612 909
rect 2606 904 2607 908
rect 2611 904 2612 908
rect 2606 903 2612 904
rect 2702 908 2708 909
rect 2702 904 2703 908
rect 2707 904 2708 908
rect 2702 903 2708 904
rect 2806 908 2812 909
rect 2806 904 2807 908
rect 2811 904 2812 908
rect 2806 903 2812 904
rect 2910 908 2916 909
rect 2910 904 2911 908
rect 2915 904 2916 908
rect 2910 903 2916 904
rect 3014 908 3020 909
rect 3014 904 3015 908
rect 3019 904 3020 908
rect 3014 903 3020 904
rect 3110 908 3116 909
rect 3110 904 3111 908
rect 3115 904 3116 908
rect 3110 903 3116 904
rect 3214 908 3220 909
rect 3214 904 3215 908
rect 3219 904 3220 908
rect 3214 903 3220 904
rect 3318 908 3324 909
rect 3318 904 3319 908
rect 3323 904 3324 908
rect 3318 903 3324 904
rect 3422 908 3428 909
rect 3422 904 3423 908
rect 3427 904 3428 908
rect 3422 903 3428 904
rect 3502 908 3508 909
rect 3502 904 3503 908
rect 3507 904 3508 908
rect 3502 903 3508 904
rect 3590 905 3596 906
rect 1870 900 1876 901
rect 3590 901 3591 905
rect 3595 901 3596 905
rect 3590 900 3596 901
rect 142 898 148 899
rect 142 894 143 898
rect 147 894 148 898
rect 142 893 148 894
rect 222 898 228 899
rect 222 894 223 898
rect 227 894 228 898
rect 222 893 228 894
rect 334 898 340 899
rect 334 894 335 898
rect 339 894 340 898
rect 334 893 340 894
rect 454 898 460 899
rect 454 894 455 898
rect 459 894 460 898
rect 454 893 460 894
rect 574 898 580 899
rect 574 894 575 898
rect 579 894 580 898
rect 574 893 580 894
rect 694 898 700 899
rect 694 894 695 898
rect 699 894 700 898
rect 694 893 700 894
rect 806 898 812 899
rect 806 894 807 898
rect 811 894 812 898
rect 806 893 812 894
rect 918 898 924 899
rect 918 894 919 898
rect 923 894 924 898
rect 918 893 924 894
rect 1022 898 1028 899
rect 1022 894 1023 898
rect 1027 894 1028 898
rect 1022 893 1028 894
rect 1126 898 1132 899
rect 1126 894 1127 898
rect 1131 894 1132 898
rect 1126 893 1132 894
rect 1230 898 1236 899
rect 1230 894 1231 898
rect 1235 894 1236 898
rect 1230 893 1236 894
rect 1334 898 1340 899
rect 1334 894 1335 898
rect 1339 894 1340 898
rect 1334 893 1340 894
rect 1870 888 1876 889
rect 1870 884 1871 888
rect 1875 884 1876 888
rect 1870 883 1876 884
rect 3590 888 3596 889
rect 3590 884 3591 888
rect 3595 884 3596 888
rect 3590 883 3596 884
rect 2286 870 2292 871
rect 2286 866 2287 870
rect 2291 866 2292 870
rect 2286 865 2292 866
rect 2366 870 2372 871
rect 2366 866 2367 870
rect 2371 866 2372 870
rect 2366 865 2372 866
rect 2446 870 2452 871
rect 2446 866 2447 870
rect 2451 866 2452 870
rect 2446 865 2452 866
rect 2526 870 2532 871
rect 2526 866 2527 870
rect 2531 866 2532 870
rect 2526 865 2532 866
rect 2614 870 2620 871
rect 2614 866 2615 870
rect 2619 866 2620 870
rect 2614 865 2620 866
rect 2710 870 2716 871
rect 2710 866 2711 870
rect 2715 866 2716 870
rect 2710 865 2716 866
rect 2814 870 2820 871
rect 2814 866 2815 870
rect 2819 866 2820 870
rect 2814 865 2820 866
rect 2918 870 2924 871
rect 2918 866 2919 870
rect 2923 866 2924 870
rect 2918 865 2924 866
rect 3022 870 3028 871
rect 3022 866 3023 870
rect 3027 866 3028 870
rect 3022 865 3028 866
rect 3118 870 3124 871
rect 3118 866 3119 870
rect 3123 866 3124 870
rect 3118 865 3124 866
rect 3222 870 3228 871
rect 3222 866 3223 870
rect 3227 866 3228 870
rect 3222 865 3228 866
rect 3326 870 3332 871
rect 3326 866 3327 870
rect 3331 866 3332 870
rect 3326 865 3332 866
rect 3430 870 3436 871
rect 3430 866 3431 870
rect 3435 866 3436 870
rect 3430 865 3436 866
rect 3510 870 3516 871
rect 3510 866 3511 870
rect 3515 866 3516 870
rect 3510 865 3516 866
rect 142 858 148 859
rect 142 854 143 858
rect 147 854 148 858
rect 142 853 148 854
rect 254 858 260 859
rect 254 854 255 858
rect 259 854 260 858
rect 254 853 260 854
rect 398 858 404 859
rect 398 854 399 858
rect 403 854 404 858
rect 398 853 404 854
rect 558 858 564 859
rect 558 854 559 858
rect 563 854 564 858
rect 558 853 564 854
rect 718 858 724 859
rect 718 854 719 858
rect 723 854 724 858
rect 718 853 724 854
rect 870 858 876 859
rect 870 854 871 858
rect 875 854 876 858
rect 870 853 876 854
rect 1014 858 1020 859
rect 1014 854 1015 858
rect 1019 854 1020 858
rect 1014 853 1020 854
rect 1150 858 1156 859
rect 1150 854 1151 858
rect 1155 854 1156 858
rect 1150 853 1156 854
rect 1278 858 1284 859
rect 1278 854 1279 858
rect 1283 854 1284 858
rect 1278 853 1284 854
rect 1398 858 1404 859
rect 1398 854 1399 858
rect 1403 854 1404 858
rect 1398 853 1404 854
rect 1518 858 1524 859
rect 1518 854 1519 858
rect 1523 854 1524 858
rect 1518 853 1524 854
rect 1646 858 1652 859
rect 1646 854 1647 858
rect 1651 854 1652 858
rect 1646 853 1652 854
rect 110 840 116 841
rect 110 836 111 840
rect 115 836 116 840
rect 110 835 116 836
rect 1830 840 1836 841
rect 1830 836 1831 840
rect 1835 836 1836 840
rect 1830 835 1836 836
rect 2166 826 2172 827
rect 110 823 116 824
rect 110 819 111 823
rect 115 819 116 823
rect 1830 823 1836 824
rect 110 818 116 819
rect 134 820 140 821
rect 134 816 135 820
rect 139 816 140 820
rect 134 815 140 816
rect 246 820 252 821
rect 246 816 247 820
rect 251 816 252 820
rect 246 815 252 816
rect 390 820 396 821
rect 390 816 391 820
rect 395 816 396 820
rect 390 815 396 816
rect 550 820 556 821
rect 550 816 551 820
rect 555 816 556 820
rect 550 815 556 816
rect 710 820 716 821
rect 710 816 711 820
rect 715 816 716 820
rect 710 815 716 816
rect 862 820 868 821
rect 862 816 863 820
rect 867 816 868 820
rect 862 815 868 816
rect 1006 820 1012 821
rect 1006 816 1007 820
rect 1011 816 1012 820
rect 1006 815 1012 816
rect 1142 820 1148 821
rect 1142 816 1143 820
rect 1147 816 1148 820
rect 1142 815 1148 816
rect 1270 820 1276 821
rect 1270 816 1271 820
rect 1275 816 1276 820
rect 1270 815 1276 816
rect 1390 820 1396 821
rect 1390 816 1391 820
rect 1395 816 1396 820
rect 1390 815 1396 816
rect 1510 820 1516 821
rect 1510 816 1511 820
rect 1515 816 1516 820
rect 1510 815 1516 816
rect 1638 820 1644 821
rect 1638 816 1639 820
rect 1643 816 1644 820
rect 1830 819 1831 823
rect 1835 819 1836 823
rect 2166 822 2167 826
rect 2171 822 2172 826
rect 2166 821 2172 822
rect 2246 826 2252 827
rect 2246 822 2247 826
rect 2251 822 2252 826
rect 2246 821 2252 822
rect 2326 826 2332 827
rect 2326 822 2327 826
rect 2331 822 2332 826
rect 2326 821 2332 822
rect 2422 826 2428 827
rect 2422 822 2423 826
rect 2427 822 2428 826
rect 2422 821 2428 822
rect 2534 826 2540 827
rect 2534 822 2535 826
rect 2539 822 2540 826
rect 2534 821 2540 822
rect 2654 826 2660 827
rect 2654 822 2655 826
rect 2659 822 2660 826
rect 2654 821 2660 822
rect 2782 826 2788 827
rect 2782 822 2783 826
rect 2787 822 2788 826
rect 2782 821 2788 822
rect 2910 826 2916 827
rect 2910 822 2911 826
rect 2915 822 2916 826
rect 2910 821 2916 822
rect 3038 826 3044 827
rect 3038 822 3039 826
rect 3043 822 3044 826
rect 3038 821 3044 822
rect 3158 826 3164 827
rect 3158 822 3159 826
rect 3163 822 3164 826
rect 3158 821 3164 822
rect 3278 826 3284 827
rect 3278 822 3279 826
rect 3283 822 3284 826
rect 3278 821 3284 822
rect 3406 826 3412 827
rect 3406 822 3407 826
rect 3411 822 3412 826
rect 3406 821 3412 822
rect 3510 826 3516 827
rect 3510 822 3511 826
rect 3515 822 3516 826
rect 3510 821 3516 822
rect 1830 818 1836 819
rect 1638 815 1644 816
rect 1870 808 1876 809
rect 1870 804 1871 808
rect 1875 804 1876 808
rect 1870 803 1876 804
rect 3590 808 3596 809
rect 3590 804 3591 808
rect 3595 804 3596 808
rect 3590 803 3596 804
rect 1870 791 1876 792
rect 1870 787 1871 791
rect 1875 787 1876 791
rect 3590 791 3596 792
rect 1870 786 1876 787
rect 2158 788 2164 789
rect 2158 784 2159 788
rect 2163 784 2164 788
rect 2158 783 2164 784
rect 2238 788 2244 789
rect 2238 784 2239 788
rect 2243 784 2244 788
rect 2238 783 2244 784
rect 2318 788 2324 789
rect 2318 784 2319 788
rect 2323 784 2324 788
rect 2318 783 2324 784
rect 2414 788 2420 789
rect 2414 784 2415 788
rect 2419 784 2420 788
rect 2414 783 2420 784
rect 2526 788 2532 789
rect 2526 784 2527 788
rect 2531 784 2532 788
rect 2526 783 2532 784
rect 2646 788 2652 789
rect 2646 784 2647 788
rect 2651 784 2652 788
rect 2646 783 2652 784
rect 2774 788 2780 789
rect 2774 784 2775 788
rect 2779 784 2780 788
rect 2774 783 2780 784
rect 2902 788 2908 789
rect 2902 784 2903 788
rect 2907 784 2908 788
rect 2902 783 2908 784
rect 3030 788 3036 789
rect 3030 784 3031 788
rect 3035 784 3036 788
rect 3030 783 3036 784
rect 3150 788 3156 789
rect 3150 784 3151 788
rect 3155 784 3156 788
rect 3150 783 3156 784
rect 3270 788 3276 789
rect 3270 784 3271 788
rect 3275 784 3276 788
rect 3270 783 3276 784
rect 3398 788 3404 789
rect 3398 784 3399 788
rect 3403 784 3404 788
rect 3398 783 3404 784
rect 3502 788 3508 789
rect 3502 784 3503 788
rect 3507 784 3508 788
rect 3590 787 3591 791
rect 3595 787 3596 791
rect 3590 786 3596 787
rect 3502 783 3508 784
rect 134 764 140 765
rect 110 761 116 762
rect 110 757 111 761
rect 115 757 116 761
rect 134 760 135 764
rect 139 760 140 764
rect 134 759 140 760
rect 262 764 268 765
rect 262 760 263 764
rect 267 760 268 764
rect 262 759 268 760
rect 430 764 436 765
rect 430 760 431 764
rect 435 760 436 764
rect 430 759 436 760
rect 606 764 612 765
rect 606 760 607 764
rect 611 760 612 764
rect 606 759 612 760
rect 782 764 788 765
rect 782 760 783 764
rect 787 760 788 764
rect 782 759 788 760
rect 950 764 956 765
rect 950 760 951 764
rect 955 760 956 764
rect 950 759 956 760
rect 1102 764 1108 765
rect 1102 760 1103 764
rect 1107 760 1108 764
rect 1102 759 1108 760
rect 1246 764 1252 765
rect 1246 760 1247 764
rect 1251 760 1252 764
rect 1246 759 1252 760
rect 1382 764 1388 765
rect 1382 760 1383 764
rect 1387 760 1388 764
rect 1382 759 1388 760
rect 1510 764 1516 765
rect 1510 760 1511 764
rect 1515 760 1516 764
rect 1510 759 1516 760
rect 1638 764 1644 765
rect 1638 760 1639 764
rect 1643 760 1644 764
rect 1638 759 1644 760
rect 1742 764 1748 765
rect 1742 760 1743 764
rect 1747 760 1748 764
rect 1742 759 1748 760
rect 1830 761 1836 762
rect 110 756 116 757
rect 1830 757 1831 761
rect 1835 757 1836 761
rect 1830 756 1836 757
rect 110 744 116 745
rect 110 740 111 744
rect 115 740 116 744
rect 110 739 116 740
rect 1830 744 1836 745
rect 1830 740 1831 744
rect 1835 740 1836 744
rect 1830 739 1836 740
rect 1894 736 1900 737
rect 1870 733 1876 734
rect 1870 729 1871 733
rect 1875 729 1876 733
rect 1894 732 1895 736
rect 1899 732 1900 736
rect 1894 731 1900 732
rect 1974 736 1980 737
rect 1974 732 1975 736
rect 1979 732 1980 736
rect 1974 731 1980 732
rect 2070 736 2076 737
rect 2070 732 2071 736
rect 2075 732 2076 736
rect 2070 731 2076 732
rect 2182 736 2188 737
rect 2182 732 2183 736
rect 2187 732 2188 736
rect 2182 731 2188 732
rect 2310 736 2316 737
rect 2310 732 2311 736
rect 2315 732 2316 736
rect 2310 731 2316 732
rect 2446 736 2452 737
rect 2446 732 2447 736
rect 2451 732 2452 736
rect 2446 731 2452 732
rect 2590 736 2596 737
rect 2590 732 2591 736
rect 2595 732 2596 736
rect 2590 731 2596 732
rect 2742 736 2748 737
rect 2742 732 2743 736
rect 2747 732 2748 736
rect 2742 731 2748 732
rect 2894 736 2900 737
rect 2894 732 2895 736
rect 2899 732 2900 736
rect 2894 731 2900 732
rect 3046 736 3052 737
rect 3046 732 3047 736
rect 3051 732 3052 736
rect 3046 731 3052 732
rect 3198 736 3204 737
rect 3198 732 3199 736
rect 3203 732 3204 736
rect 3198 731 3204 732
rect 3358 736 3364 737
rect 3358 732 3359 736
rect 3363 732 3364 736
rect 3358 731 3364 732
rect 3502 736 3508 737
rect 3502 732 3503 736
rect 3507 732 3508 736
rect 3502 731 3508 732
rect 3590 733 3596 734
rect 1870 728 1876 729
rect 3590 729 3591 733
rect 3595 729 3596 733
rect 3590 728 3596 729
rect 142 726 148 727
rect 142 722 143 726
rect 147 722 148 726
rect 142 721 148 722
rect 270 726 276 727
rect 270 722 271 726
rect 275 722 276 726
rect 270 721 276 722
rect 438 726 444 727
rect 438 722 439 726
rect 443 722 444 726
rect 438 721 444 722
rect 614 726 620 727
rect 614 722 615 726
rect 619 722 620 726
rect 614 721 620 722
rect 790 726 796 727
rect 790 722 791 726
rect 795 722 796 726
rect 790 721 796 722
rect 958 726 964 727
rect 958 722 959 726
rect 963 722 964 726
rect 958 721 964 722
rect 1110 726 1116 727
rect 1110 722 1111 726
rect 1115 722 1116 726
rect 1110 721 1116 722
rect 1254 726 1260 727
rect 1254 722 1255 726
rect 1259 722 1260 726
rect 1254 721 1260 722
rect 1390 726 1396 727
rect 1390 722 1391 726
rect 1395 722 1396 726
rect 1390 721 1396 722
rect 1518 726 1524 727
rect 1518 722 1519 726
rect 1523 722 1524 726
rect 1518 721 1524 722
rect 1646 726 1652 727
rect 1646 722 1647 726
rect 1651 722 1652 726
rect 1646 721 1652 722
rect 1750 726 1756 727
rect 1750 722 1751 726
rect 1755 722 1756 726
rect 1750 721 1756 722
rect 1870 716 1876 717
rect 1870 712 1871 716
rect 1875 712 1876 716
rect 1870 711 1876 712
rect 3590 716 3596 717
rect 3590 712 3591 716
rect 3595 712 3596 716
rect 3590 711 3596 712
rect 1902 698 1908 699
rect 1902 694 1903 698
rect 1907 694 1908 698
rect 1902 693 1908 694
rect 1982 698 1988 699
rect 1982 694 1983 698
rect 1987 694 1988 698
rect 1982 693 1988 694
rect 2078 698 2084 699
rect 2078 694 2079 698
rect 2083 694 2084 698
rect 2078 693 2084 694
rect 2190 698 2196 699
rect 2190 694 2191 698
rect 2195 694 2196 698
rect 2190 693 2196 694
rect 2318 698 2324 699
rect 2318 694 2319 698
rect 2323 694 2324 698
rect 2318 693 2324 694
rect 2454 698 2460 699
rect 2454 694 2455 698
rect 2459 694 2460 698
rect 2454 693 2460 694
rect 2598 698 2604 699
rect 2598 694 2599 698
rect 2603 694 2604 698
rect 2598 693 2604 694
rect 2750 698 2756 699
rect 2750 694 2751 698
rect 2755 694 2756 698
rect 2750 693 2756 694
rect 2902 698 2908 699
rect 2902 694 2903 698
rect 2907 694 2908 698
rect 2902 693 2908 694
rect 3054 698 3060 699
rect 3054 694 3055 698
rect 3059 694 3060 698
rect 3054 693 3060 694
rect 3206 698 3212 699
rect 3206 694 3207 698
rect 3211 694 3212 698
rect 3206 693 3212 694
rect 3366 698 3372 699
rect 3366 694 3367 698
rect 3371 694 3372 698
rect 3366 693 3372 694
rect 3510 698 3516 699
rect 3510 694 3511 698
rect 3515 694 3516 698
rect 3510 693 3516 694
rect 294 682 300 683
rect 294 678 295 682
rect 299 678 300 682
rect 294 677 300 678
rect 406 682 412 683
rect 406 678 407 682
rect 411 678 412 682
rect 406 677 412 678
rect 526 682 532 683
rect 526 678 527 682
rect 531 678 532 682
rect 526 677 532 678
rect 654 682 660 683
rect 654 678 655 682
rect 659 678 660 682
rect 654 677 660 678
rect 782 682 788 683
rect 782 678 783 682
rect 787 678 788 682
rect 782 677 788 678
rect 902 682 908 683
rect 902 678 903 682
rect 907 678 908 682
rect 902 677 908 678
rect 1022 682 1028 683
rect 1022 678 1023 682
rect 1027 678 1028 682
rect 1022 677 1028 678
rect 1134 682 1140 683
rect 1134 678 1135 682
rect 1139 678 1140 682
rect 1134 677 1140 678
rect 1246 682 1252 683
rect 1246 678 1247 682
rect 1251 678 1252 682
rect 1246 677 1252 678
rect 1350 682 1356 683
rect 1350 678 1351 682
rect 1355 678 1356 682
rect 1350 677 1356 678
rect 1454 682 1460 683
rect 1454 678 1455 682
rect 1459 678 1460 682
rect 1454 677 1460 678
rect 1558 682 1564 683
rect 1558 678 1559 682
rect 1563 678 1564 682
rect 1558 677 1564 678
rect 1662 682 1668 683
rect 1662 678 1663 682
rect 1667 678 1668 682
rect 1662 677 1668 678
rect 1750 682 1756 683
rect 1750 678 1751 682
rect 1755 678 1756 682
rect 1750 677 1756 678
rect 110 664 116 665
rect 110 660 111 664
rect 115 660 116 664
rect 110 659 116 660
rect 1830 664 1836 665
rect 1830 660 1831 664
rect 1835 660 1836 664
rect 1830 659 1836 660
rect 1902 662 1908 663
rect 1902 658 1903 662
rect 1907 658 1908 662
rect 1902 657 1908 658
rect 2094 662 2100 663
rect 2094 658 2095 662
rect 2099 658 2100 662
rect 2094 657 2100 658
rect 2294 662 2300 663
rect 2294 658 2295 662
rect 2299 658 2300 662
rect 2294 657 2300 658
rect 2478 662 2484 663
rect 2478 658 2479 662
rect 2483 658 2484 662
rect 2478 657 2484 658
rect 2654 662 2660 663
rect 2654 658 2655 662
rect 2659 658 2660 662
rect 2654 657 2660 658
rect 2830 662 2836 663
rect 2830 658 2831 662
rect 2835 658 2836 662
rect 2830 657 2836 658
rect 3006 662 3012 663
rect 3006 658 3007 662
rect 3011 658 3012 662
rect 3006 657 3012 658
rect 3182 662 3188 663
rect 3182 658 3183 662
rect 3187 658 3188 662
rect 3182 657 3188 658
rect 3358 662 3364 663
rect 3358 658 3359 662
rect 3363 658 3364 662
rect 3358 657 3364 658
rect 3510 662 3516 663
rect 3510 658 3511 662
rect 3515 658 3516 662
rect 3510 657 3516 658
rect 110 647 116 648
rect 110 643 111 647
rect 115 643 116 647
rect 1830 647 1836 648
rect 110 642 116 643
rect 286 644 292 645
rect 286 640 287 644
rect 291 640 292 644
rect 286 639 292 640
rect 398 644 404 645
rect 398 640 399 644
rect 403 640 404 644
rect 398 639 404 640
rect 518 644 524 645
rect 518 640 519 644
rect 523 640 524 644
rect 518 639 524 640
rect 646 644 652 645
rect 646 640 647 644
rect 651 640 652 644
rect 646 639 652 640
rect 774 644 780 645
rect 774 640 775 644
rect 779 640 780 644
rect 774 639 780 640
rect 894 644 900 645
rect 894 640 895 644
rect 899 640 900 644
rect 894 639 900 640
rect 1014 644 1020 645
rect 1014 640 1015 644
rect 1019 640 1020 644
rect 1014 639 1020 640
rect 1126 644 1132 645
rect 1126 640 1127 644
rect 1131 640 1132 644
rect 1126 639 1132 640
rect 1238 644 1244 645
rect 1238 640 1239 644
rect 1243 640 1244 644
rect 1238 639 1244 640
rect 1342 644 1348 645
rect 1342 640 1343 644
rect 1347 640 1348 644
rect 1342 639 1348 640
rect 1446 644 1452 645
rect 1446 640 1447 644
rect 1451 640 1452 644
rect 1446 639 1452 640
rect 1550 644 1556 645
rect 1550 640 1551 644
rect 1555 640 1556 644
rect 1550 639 1556 640
rect 1654 644 1660 645
rect 1654 640 1655 644
rect 1659 640 1660 644
rect 1654 639 1660 640
rect 1742 644 1748 645
rect 1742 640 1743 644
rect 1747 640 1748 644
rect 1830 643 1831 647
rect 1835 643 1836 647
rect 1830 642 1836 643
rect 1870 644 1876 645
rect 1742 639 1748 640
rect 1870 640 1871 644
rect 1875 640 1876 644
rect 1870 639 1876 640
rect 3590 644 3596 645
rect 3590 640 3591 644
rect 3595 640 3596 644
rect 3590 639 3596 640
rect 1870 627 1876 628
rect 1870 623 1871 627
rect 1875 623 1876 627
rect 3590 627 3596 628
rect 1870 622 1876 623
rect 1894 624 1900 625
rect 1894 620 1895 624
rect 1899 620 1900 624
rect 1894 619 1900 620
rect 2086 624 2092 625
rect 2086 620 2087 624
rect 2091 620 2092 624
rect 2086 619 2092 620
rect 2286 624 2292 625
rect 2286 620 2287 624
rect 2291 620 2292 624
rect 2286 619 2292 620
rect 2470 624 2476 625
rect 2470 620 2471 624
rect 2475 620 2476 624
rect 2470 619 2476 620
rect 2646 624 2652 625
rect 2646 620 2647 624
rect 2651 620 2652 624
rect 2646 619 2652 620
rect 2822 624 2828 625
rect 2822 620 2823 624
rect 2827 620 2828 624
rect 2822 619 2828 620
rect 2998 624 3004 625
rect 2998 620 2999 624
rect 3003 620 3004 624
rect 2998 619 3004 620
rect 3174 624 3180 625
rect 3174 620 3175 624
rect 3179 620 3180 624
rect 3174 619 3180 620
rect 3350 624 3356 625
rect 3350 620 3351 624
rect 3355 620 3356 624
rect 3350 619 3356 620
rect 3502 624 3508 625
rect 3502 620 3503 624
rect 3507 620 3508 624
rect 3590 623 3591 627
rect 3595 623 3596 627
rect 3590 622 3596 623
rect 3502 619 3508 620
rect 310 596 316 597
rect 110 593 116 594
rect 110 589 111 593
rect 115 589 116 593
rect 310 592 311 596
rect 315 592 316 596
rect 310 591 316 592
rect 390 596 396 597
rect 390 592 391 596
rect 395 592 396 596
rect 390 591 396 592
rect 470 596 476 597
rect 470 592 471 596
rect 475 592 476 596
rect 470 591 476 592
rect 558 596 564 597
rect 558 592 559 596
rect 563 592 564 596
rect 558 591 564 592
rect 646 596 652 597
rect 646 592 647 596
rect 651 592 652 596
rect 646 591 652 592
rect 734 596 740 597
rect 734 592 735 596
rect 739 592 740 596
rect 734 591 740 592
rect 822 596 828 597
rect 822 592 823 596
rect 827 592 828 596
rect 822 591 828 592
rect 910 596 916 597
rect 910 592 911 596
rect 915 592 916 596
rect 910 591 916 592
rect 998 596 1004 597
rect 998 592 999 596
rect 1003 592 1004 596
rect 998 591 1004 592
rect 1086 596 1092 597
rect 1086 592 1087 596
rect 1091 592 1092 596
rect 1086 591 1092 592
rect 1174 596 1180 597
rect 1174 592 1175 596
rect 1179 592 1180 596
rect 1174 591 1180 592
rect 1262 596 1268 597
rect 1262 592 1263 596
rect 1267 592 1268 596
rect 1262 591 1268 592
rect 1830 593 1836 594
rect 110 588 116 589
rect 1830 589 1831 593
rect 1835 589 1836 593
rect 1830 588 1836 589
rect 110 576 116 577
rect 110 572 111 576
rect 115 572 116 576
rect 110 571 116 572
rect 1830 576 1836 577
rect 1830 572 1831 576
rect 1835 572 1836 576
rect 1894 576 1900 577
rect 1830 571 1836 572
rect 1870 573 1876 574
rect 1870 569 1871 573
rect 1875 569 1876 573
rect 1894 572 1895 576
rect 1899 572 1900 576
rect 1894 571 1900 572
rect 1974 576 1980 577
rect 1974 572 1975 576
rect 1979 572 1980 576
rect 1974 571 1980 572
rect 2086 576 2092 577
rect 2086 572 2087 576
rect 2091 572 2092 576
rect 2086 571 2092 572
rect 2214 576 2220 577
rect 2214 572 2215 576
rect 2219 572 2220 576
rect 2214 571 2220 572
rect 2350 576 2356 577
rect 2350 572 2351 576
rect 2355 572 2356 576
rect 2350 571 2356 572
rect 2494 576 2500 577
rect 2494 572 2495 576
rect 2499 572 2500 576
rect 2494 571 2500 572
rect 2646 576 2652 577
rect 2646 572 2647 576
rect 2651 572 2652 576
rect 2646 571 2652 572
rect 2806 576 2812 577
rect 2806 572 2807 576
rect 2811 572 2812 576
rect 2806 571 2812 572
rect 2974 576 2980 577
rect 2974 572 2975 576
rect 2979 572 2980 576
rect 2974 571 2980 572
rect 3150 576 3156 577
rect 3150 572 3151 576
rect 3155 572 3156 576
rect 3150 571 3156 572
rect 3334 576 3340 577
rect 3334 572 3335 576
rect 3339 572 3340 576
rect 3334 571 3340 572
rect 3502 576 3508 577
rect 3502 572 3503 576
rect 3507 572 3508 576
rect 3502 571 3508 572
rect 3590 573 3596 574
rect 1870 568 1876 569
rect 3590 569 3591 573
rect 3595 569 3596 573
rect 3590 568 3596 569
rect 318 558 324 559
rect 318 554 319 558
rect 323 554 324 558
rect 318 553 324 554
rect 398 558 404 559
rect 398 554 399 558
rect 403 554 404 558
rect 398 553 404 554
rect 478 558 484 559
rect 478 554 479 558
rect 483 554 484 558
rect 478 553 484 554
rect 566 558 572 559
rect 566 554 567 558
rect 571 554 572 558
rect 566 553 572 554
rect 654 558 660 559
rect 654 554 655 558
rect 659 554 660 558
rect 654 553 660 554
rect 742 558 748 559
rect 742 554 743 558
rect 747 554 748 558
rect 742 553 748 554
rect 830 558 836 559
rect 830 554 831 558
rect 835 554 836 558
rect 830 553 836 554
rect 918 558 924 559
rect 918 554 919 558
rect 923 554 924 558
rect 918 553 924 554
rect 1006 558 1012 559
rect 1006 554 1007 558
rect 1011 554 1012 558
rect 1006 553 1012 554
rect 1094 558 1100 559
rect 1094 554 1095 558
rect 1099 554 1100 558
rect 1094 553 1100 554
rect 1182 558 1188 559
rect 1182 554 1183 558
rect 1187 554 1188 558
rect 1182 553 1188 554
rect 1270 558 1276 559
rect 1270 554 1271 558
rect 1275 554 1276 558
rect 1270 553 1276 554
rect 1870 556 1876 557
rect 1870 552 1871 556
rect 1875 552 1876 556
rect 1870 551 1876 552
rect 3590 556 3596 557
rect 3590 552 3591 556
rect 3595 552 3596 556
rect 3590 551 3596 552
rect 1902 538 1908 539
rect 1902 534 1903 538
rect 1907 534 1908 538
rect 1902 533 1908 534
rect 1982 538 1988 539
rect 1982 534 1983 538
rect 1987 534 1988 538
rect 1982 533 1988 534
rect 2094 538 2100 539
rect 2094 534 2095 538
rect 2099 534 2100 538
rect 2094 533 2100 534
rect 2222 538 2228 539
rect 2222 534 2223 538
rect 2227 534 2228 538
rect 2222 533 2228 534
rect 2358 538 2364 539
rect 2358 534 2359 538
rect 2363 534 2364 538
rect 2358 533 2364 534
rect 2502 538 2508 539
rect 2502 534 2503 538
rect 2507 534 2508 538
rect 2502 533 2508 534
rect 2654 538 2660 539
rect 2654 534 2655 538
rect 2659 534 2660 538
rect 2654 533 2660 534
rect 2814 538 2820 539
rect 2814 534 2815 538
rect 2819 534 2820 538
rect 2814 533 2820 534
rect 2982 538 2988 539
rect 2982 534 2983 538
rect 2987 534 2988 538
rect 2982 533 2988 534
rect 3158 538 3164 539
rect 3158 534 3159 538
rect 3163 534 3164 538
rect 3158 533 3164 534
rect 3342 538 3348 539
rect 3342 534 3343 538
rect 3347 534 3348 538
rect 3342 533 3348 534
rect 3510 538 3516 539
rect 3510 534 3511 538
rect 3515 534 3516 538
rect 3510 533 3516 534
rect 238 514 244 515
rect 238 510 239 514
rect 243 510 244 514
rect 238 509 244 510
rect 342 514 348 515
rect 342 510 343 514
rect 347 510 348 514
rect 342 509 348 510
rect 438 514 444 515
rect 438 510 439 514
rect 443 510 444 514
rect 438 509 444 510
rect 534 514 540 515
rect 534 510 535 514
rect 539 510 540 514
rect 534 509 540 510
rect 630 514 636 515
rect 630 510 631 514
rect 635 510 636 514
rect 630 509 636 510
rect 718 514 724 515
rect 718 510 719 514
rect 723 510 724 514
rect 718 509 724 510
rect 806 514 812 515
rect 806 510 807 514
rect 811 510 812 514
rect 806 509 812 510
rect 894 514 900 515
rect 894 510 895 514
rect 899 510 900 514
rect 894 509 900 510
rect 982 514 988 515
rect 982 510 983 514
rect 987 510 988 514
rect 982 509 988 510
rect 1070 514 1076 515
rect 1070 510 1071 514
rect 1075 510 1076 514
rect 1070 509 1076 510
rect 1158 514 1164 515
rect 1158 510 1159 514
rect 1163 510 1164 514
rect 1158 509 1164 510
rect 1246 514 1252 515
rect 1246 510 1247 514
rect 1251 510 1252 514
rect 1246 509 1252 510
rect 2150 506 2156 507
rect 2150 502 2151 506
rect 2155 502 2156 506
rect 2150 501 2156 502
rect 2230 506 2236 507
rect 2230 502 2231 506
rect 2235 502 2236 506
rect 2230 501 2236 502
rect 2326 506 2332 507
rect 2326 502 2327 506
rect 2331 502 2332 506
rect 2326 501 2332 502
rect 2430 506 2436 507
rect 2430 502 2431 506
rect 2435 502 2436 506
rect 2430 501 2436 502
rect 2550 506 2556 507
rect 2550 502 2551 506
rect 2555 502 2556 506
rect 2550 501 2556 502
rect 2686 506 2692 507
rect 2686 502 2687 506
rect 2691 502 2692 506
rect 2686 501 2692 502
rect 2838 506 2844 507
rect 2838 502 2839 506
rect 2843 502 2844 506
rect 2838 501 2844 502
rect 2998 506 3004 507
rect 2998 502 2999 506
rect 3003 502 3004 506
rect 2998 501 3004 502
rect 3174 506 3180 507
rect 3174 502 3175 506
rect 3179 502 3180 506
rect 3174 501 3180 502
rect 3350 506 3356 507
rect 3350 502 3351 506
rect 3355 502 3356 506
rect 3350 501 3356 502
rect 3510 506 3516 507
rect 3510 502 3511 506
rect 3515 502 3516 506
rect 3510 501 3516 502
rect 110 496 116 497
rect 110 492 111 496
rect 115 492 116 496
rect 110 491 116 492
rect 1830 496 1836 497
rect 1830 492 1831 496
rect 1835 492 1836 496
rect 1830 491 1836 492
rect 1870 488 1876 489
rect 1870 484 1871 488
rect 1875 484 1876 488
rect 1870 483 1876 484
rect 3590 488 3596 489
rect 3590 484 3591 488
rect 3595 484 3596 488
rect 3590 483 3596 484
rect 110 479 116 480
rect 110 475 111 479
rect 115 475 116 479
rect 1830 479 1836 480
rect 110 474 116 475
rect 230 476 236 477
rect 230 472 231 476
rect 235 472 236 476
rect 230 471 236 472
rect 334 476 340 477
rect 334 472 335 476
rect 339 472 340 476
rect 334 471 340 472
rect 430 476 436 477
rect 430 472 431 476
rect 435 472 436 476
rect 430 471 436 472
rect 526 476 532 477
rect 526 472 527 476
rect 531 472 532 476
rect 526 471 532 472
rect 622 476 628 477
rect 622 472 623 476
rect 627 472 628 476
rect 622 471 628 472
rect 710 476 716 477
rect 710 472 711 476
rect 715 472 716 476
rect 710 471 716 472
rect 798 476 804 477
rect 798 472 799 476
rect 803 472 804 476
rect 798 471 804 472
rect 886 476 892 477
rect 886 472 887 476
rect 891 472 892 476
rect 886 471 892 472
rect 974 476 980 477
rect 974 472 975 476
rect 979 472 980 476
rect 974 471 980 472
rect 1062 476 1068 477
rect 1062 472 1063 476
rect 1067 472 1068 476
rect 1062 471 1068 472
rect 1150 476 1156 477
rect 1150 472 1151 476
rect 1155 472 1156 476
rect 1150 471 1156 472
rect 1238 476 1244 477
rect 1238 472 1239 476
rect 1243 472 1244 476
rect 1830 475 1831 479
rect 1835 475 1836 479
rect 1830 474 1836 475
rect 1238 471 1244 472
rect 1870 471 1876 472
rect 1870 467 1871 471
rect 1875 467 1876 471
rect 3590 471 3596 472
rect 1870 466 1876 467
rect 2142 468 2148 469
rect 2142 464 2143 468
rect 2147 464 2148 468
rect 2142 463 2148 464
rect 2222 468 2228 469
rect 2222 464 2223 468
rect 2227 464 2228 468
rect 2222 463 2228 464
rect 2318 468 2324 469
rect 2318 464 2319 468
rect 2323 464 2324 468
rect 2318 463 2324 464
rect 2422 468 2428 469
rect 2422 464 2423 468
rect 2427 464 2428 468
rect 2422 463 2428 464
rect 2542 468 2548 469
rect 2542 464 2543 468
rect 2547 464 2548 468
rect 2542 463 2548 464
rect 2678 468 2684 469
rect 2678 464 2679 468
rect 2683 464 2684 468
rect 2678 463 2684 464
rect 2830 468 2836 469
rect 2830 464 2831 468
rect 2835 464 2836 468
rect 2830 463 2836 464
rect 2990 468 2996 469
rect 2990 464 2991 468
rect 2995 464 2996 468
rect 2990 463 2996 464
rect 3166 468 3172 469
rect 3166 464 3167 468
rect 3171 464 3172 468
rect 3166 463 3172 464
rect 3342 468 3348 469
rect 3342 464 3343 468
rect 3347 464 3348 468
rect 3342 463 3348 464
rect 3502 468 3508 469
rect 3502 464 3503 468
rect 3507 464 3508 468
rect 3590 467 3591 471
rect 3595 467 3596 471
rect 3590 466 3596 467
rect 3502 463 3508 464
rect 134 424 140 425
rect 110 421 116 422
rect 110 417 111 421
rect 115 417 116 421
rect 134 420 135 424
rect 139 420 140 424
rect 134 419 140 420
rect 246 424 252 425
rect 246 420 247 424
rect 251 420 252 424
rect 246 419 252 420
rect 374 424 380 425
rect 374 420 375 424
rect 379 420 380 424
rect 374 419 380 420
rect 494 424 500 425
rect 494 420 495 424
rect 499 420 500 424
rect 494 419 500 420
rect 606 424 612 425
rect 606 420 607 424
rect 611 420 612 424
rect 606 419 612 420
rect 718 424 724 425
rect 718 420 719 424
rect 723 420 724 424
rect 718 419 724 420
rect 822 424 828 425
rect 822 420 823 424
rect 827 420 828 424
rect 822 419 828 420
rect 918 424 924 425
rect 918 420 919 424
rect 923 420 924 424
rect 918 419 924 420
rect 1006 424 1012 425
rect 1006 420 1007 424
rect 1011 420 1012 424
rect 1006 419 1012 420
rect 1102 424 1108 425
rect 1102 420 1103 424
rect 1107 420 1108 424
rect 1102 419 1108 420
rect 1198 424 1204 425
rect 1198 420 1199 424
rect 1203 420 1204 424
rect 1198 419 1204 420
rect 1294 424 1300 425
rect 1294 420 1295 424
rect 1299 420 1300 424
rect 1294 419 1300 420
rect 1830 421 1836 422
rect 110 416 116 417
rect 1830 417 1831 421
rect 1835 417 1836 421
rect 2334 420 2340 421
rect 1830 416 1836 417
rect 1870 417 1876 418
rect 1870 413 1871 417
rect 1875 413 1876 417
rect 2334 416 2335 420
rect 2339 416 2340 420
rect 2334 415 2340 416
rect 2414 420 2420 421
rect 2414 416 2415 420
rect 2419 416 2420 420
rect 2414 415 2420 416
rect 2494 420 2500 421
rect 2494 416 2495 420
rect 2499 416 2500 420
rect 2494 415 2500 416
rect 2582 420 2588 421
rect 2582 416 2583 420
rect 2587 416 2588 420
rect 2582 415 2588 416
rect 2686 420 2692 421
rect 2686 416 2687 420
rect 2691 416 2692 420
rect 2686 415 2692 416
rect 2798 420 2804 421
rect 2798 416 2799 420
rect 2803 416 2804 420
rect 2798 415 2804 416
rect 2926 420 2932 421
rect 2926 416 2927 420
rect 2931 416 2932 420
rect 2926 415 2932 416
rect 3070 420 3076 421
rect 3070 416 3071 420
rect 3075 416 3076 420
rect 3070 415 3076 416
rect 3214 420 3220 421
rect 3214 416 3215 420
rect 3219 416 3220 420
rect 3214 415 3220 416
rect 3366 420 3372 421
rect 3366 416 3367 420
rect 3371 416 3372 420
rect 3366 415 3372 416
rect 3502 420 3508 421
rect 3502 416 3503 420
rect 3507 416 3508 420
rect 3502 415 3508 416
rect 3590 417 3596 418
rect 1870 412 1876 413
rect 3590 413 3591 417
rect 3595 413 3596 417
rect 3590 412 3596 413
rect 110 404 116 405
rect 110 400 111 404
rect 115 400 116 404
rect 110 399 116 400
rect 1830 404 1836 405
rect 1830 400 1831 404
rect 1835 400 1836 404
rect 1830 399 1836 400
rect 1870 400 1876 401
rect 1870 396 1871 400
rect 1875 396 1876 400
rect 1870 395 1876 396
rect 3590 400 3596 401
rect 3590 396 3591 400
rect 3595 396 3596 400
rect 3590 395 3596 396
rect 142 386 148 387
rect 142 382 143 386
rect 147 382 148 386
rect 142 381 148 382
rect 254 386 260 387
rect 254 382 255 386
rect 259 382 260 386
rect 254 381 260 382
rect 382 386 388 387
rect 382 382 383 386
rect 387 382 388 386
rect 382 381 388 382
rect 502 386 508 387
rect 502 382 503 386
rect 507 382 508 386
rect 502 381 508 382
rect 614 386 620 387
rect 614 382 615 386
rect 619 382 620 386
rect 614 381 620 382
rect 726 386 732 387
rect 726 382 727 386
rect 731 382 732 386
rect 726 381 732 382
rect 830 386 836 387
rect 830 382 831 386
rect 835 382 836 386
rect 830 381 836 382
rect 926 386 932 387
rect 926 382 927 386
rect 931 382 932 386
rect 926 381 932 382
rect 1014 386 1020 387
rect 1014 382 1015 386
rect 1019 382 1020 386
rect 1014 381 1020 382
rect 1110 386 1116 387
rect 1110 382 1111 386
rect 1115 382 1116 386
rect 1110 381 1116 382
rect 1206 386 1212 387
rect 1206 382 1207 386
rect 1211 382 1212 386
rect 1206 381 1212 382
rect 1302 386 1308 387
rect 1302 382 1303 386
rect 1307 382 1308 386
rect 1302 381 1308 382
rect 2342 382 2348 383
rect 2342 378 2343 382
rect 2347 378 2348 382
rect 2342 377 2348 378
rect 2422 382 2428 383
rect 2422 378 2423 382
rect 2427 378 2428 382
rect 2422 377 2428 378
rect 2502 382 2508 383
rect 2502 378 2503 382
rect 2507 378 2508 382
rect 2502 377 2508 378
rect 2590 382 2596 383
rect 2590 378 2591 382
rect 2595 378 2596 382
rect 2590 377 2596 378
rect 2694 382 2700 383
rect 2694 378 2695 382
rect 2699 378 2700 382
rect 2694 377 2700 378
rect 2806 382 2812 383
rect 2806 378 2807 382
rect 2811 378 2812 382
rect 2806 377 2812 378
rect 2934 382 2940 383
rect 2934 378 2935 382
rect 2939 378 2940 382
rect 2934 377 2940 378
rect 3078 382 3084 383
rect 3078 378 3079 382
rect 3083 378 3084 382
rect 3078 377 3084 378
rect 3222 382 3228 383
rect 3222 378 3223 382
rect 3227 378 3228 382
rect 3222 377 3228 378
rect 3374 382 3380 383
rect 3374 378 3375 382
rect 3379 378 3380 382
rect 3374 377 3380 378
rect 3510 382 3516 383
rect 3510 378 3511 382
rect 3515 378 3516 382
rect 3510 377 3516 378
rect 142 342 148 343
rect 142 338 143 342
rect 147 338 148 342
rect 142 337 148 338
rect 246 342 252 343
rect 246 338 247 342
rect 251 338 252 342
rect 246 337 252 338
rect 374 342 380 343
rect 374 338 375 342
rect 379 338 380 342
rect 374 337 380 338
rect 510 342 516 343
rect 510 338 511 342
rect 515 338 516 342
rect 510 337 516 338
rect 646 342 652 343
rect 646 338 647 342
rect 651 338 652 342
rect 646 337 652 338
rect 774 342 780 343
rect 774 338 775 342
rect 779 338 780 342
rect 774 337 780 338
rect 894 342 900 343
rect 894 338 895 342
rect 899 338 900 342
rect 894 337 900 338
rect 1006 342 1012 343
rect 1006 338 1007 342
rect 1011 338 1012 342
rect 1006 337 1012 338
rect 1118 342 1124 343
rect 1118 338 1119 342
rect 1123 338 1124 342
rect 1118 337 1124 338
rect 1222 342 1228 343
rect 1222 338 1223 342
rect 1227 338 1228 342
rect 1222 337 1228 338
rect 1326 342 1332 343
rect 1326 338 1327 342
rect 1331 338 1332 342
rect 1326 337 1332 338
rect 1438 342 1444 343
rect 1438 338 1439 342
rect 1443 338 1444 342
rect 1438 337 1444 338
rect 2078 342 2084 343
rect 2078 338 2079 342
rect 2083 338 2084 342
rect 2078 337 2084 338
rect 2166 342 2172 343
rect 2166 338 2167 342
rect 2171 338 2172 342
rect 2166 337 2172 338
rect 2262 342 2268 343
rect 2262 338 2263 342
rect 2267 338 2268 342
rect 2262 337 2268 338
rect 2374 342 2380 343
rect 2374 338 2375 342
rect 2379 338 2380 342
rect 2374 337 2380 338
rect 2502 342 2508 343
rect 2502 338 2503 342
rect 2507 338 2508 342
rect 2502 337 2508 338
rect 2638 342 2644 343
rect 2638 338 2639 342
rect 2643 338 2644 342
rect 2638 337 2644 338
rect 2774 342 2780 343
rect 2774 338 2775 342
rect 2779 338 2780 342
rect 2774 337 2780 338
rect 2910 342 2916 343
rect 2910 338 2911 342
rect 2915 338 2916 342
rect 2910 337 2916 338
rect 3038 342 3044 343
rect 3038 338 3039 342
rect 3043 338 3044 342
rect 3038 337 3044 338
rect 3166 342 3172 343
rect 3166 338 3167 342
rect 3171 338 3172 342
rect 3166 337 3172 338
rect 3286 342 3292 343
rect 3286 338 3287 342
rect 3291 338 3292 342
rect 3286 337 3292 338
rect 3406 342 3412 343
rect 3406 338 3407 342
rect 3411 338 3412 342
rect 3406 337 3412 338
rect 3510 342 3516 343
rect 3510 338 3511 342
rect 3515 338 3516 342
rect 3510 337 3516 338
rect 110 324 116 325
rect 110 320 111 324
rect 115 320 116 324
rect 110 319 116 320
rect 1830 324 1836 325
rect 1830 320 1831 324
rect 1835 320 1836 324
rect 1830 319 1836 320
rect 1870 324 1876 325
rect 1870 320 1871 324
rect 1875 320 1876 324
rect 1870 319 1876 320
rect 3590 324 3596 325
rect 3590 320 3591 324
rect 3595 320 3596 324
rect 3590 319 3596 320
rect 110 307 116 308
rect 110 303 111 307
rect 115 303 116 307
rect 1830 307 1836 308
rect 110 302 116 303
rect 134 304 140 305
rect 134 300 135 304
rect 139 300 140 304
rect 134 299 140 300
rect 238 304 244 305
rect 238 300 239 304
rect 243 300 244 304
rect 238 299 244 300
rect 366 304 372 305
rect 366 300 367 304
rect 371 300 372 304
rect 366 299 372 300
rect 502 304 508 305
rect 502 300 503 304
rect 507 300 508 304
rect 502 299 508 300
rect 638 304 644 305
rect 638 300 639 304
rect 643 300 644 304
rect 638 299 644 300
rect 766 304 772 305
rect 766 300 767 304
rect 771 300 772 304
rect 766 299 772 300
rect 886 304 892 305
rect 886 300 887 304
rect 891 300 892 304
rect 886 299 892 300
rect 998 304 1004 305
rect 998 300 999 304
rect 1003 300 1004 304
rect 998 299 1004 300
rect 1110 304 1116 305
rect 1110 300 1111 304
rect 1115 300 1116 304
rect 1110 299 1116 300
rect 1214 304 1220 305
rect 1214 300 1215 304
rect 1219 300 1220 304
rect 1214 299 1220 300
rect 1318 304 1324 305
rect 1318 300 1319 304
rect 1323 300 1324 304
rect 1318 299 1324 300
rect 1430 304 1436 305
rect 1430 300 1431 304
rect 1435 300 1436 304
rect 1830 303 1831 307
rect 1835 303 1836 307
rect 1830 302 1836 303
rect 1870 307 1876 308
rect 1870 303 1871 307
rect 1875 303 1876 307
rect 3590 307 3596 308
rect 1870 302 1876 303
rect 2070 304 2076 305
rect 1430 299 1436 300
rect 2070 300 2071 304
rect 2075 300 2076 304
rect 2070 299 2076 300
rect 2158 304 2164 305
rect 2158 300 2159 304
rect 2163 300 2164 304
rect 2158 299 2164 300
rect 2254 304 2260 305
rect 2254 300 2255 304
rect 2259 300 2260 304
rect 2254 299 2260 300
rect 2366 304 2372 305
rect 2366 300 2367 304
rect 2371 300 2372 304
rect 2366 299 2372 300
rect 2494 304 2500 305
rect 2494 300 2495 304
rect 2499 300 2500 304
rect 2494 299 2500 300
rect 2630 304 2636 305
rect 2630 300 2631 304
rect 2635 300 2636 304
rect 2630 299 2636 300
rect 2766 304 2772 305
rect 2766 300 2767 304
rect 2771 300 2772 304
rect 2766 299 2772 300
rect 2902 304 2908 305
rect 2902 300 2903 304
rect 2907 300 2908 304
rect 2902 299 2908 300
rect 3030 304 3036 305
rect 3030 300 3031 304
rect 3035 300 3036 304
rect 3030 299 3036 300
rect 3158 304 3164 305
rect 3158 300 3159 304
rect 3163 300 3164 304
rect 3158 299 3164 300
rect 3278 304 3284 305
rect 3278 300 3279 304
rect 3283 300 3284 304
rect 3278 299 3284 300
rect 3398 304 3404 305
rect 3398 300 3399 304
rect 3403 300 3404 304
rect 3398 299 3404 300
rect 3502 304 3508 305
rect 3502 300 3503 304
rect 3507 300 3508 304
rect 3590 303 3591 307
rect 3595 303 3596 307
rect 3590 302 3596 303
rect 3502 299 3508 300
rect 222 252 228 253
rect 110 249 116 250
rect 110 245 111 249
rect 115 245 116 249
rect 222 248 223 252
rect 227 248 228 252
rect 222 247 228 248
rect 334 252 340 253
rect 334 248 335 252
rect 339 248 340 252
rect 334 247 340 248
rect 462 252 468 253
rect 462 248 463 252
rect 467 248 468 252
rect 462 247 468 248
rect 598 252 604 253
rect 598 248 599 252
rect 603 248 604 252
rect 598 247 604 248
rect 734 252 740 253
rect 734 248 735 252
rect 739 248 740 252
rect 734 247 740 248
rect 870 252 876 253
rect 870 248 871 252
rect 875 248 876 252
rect 870 247 876 248
rect 1006 252 1012 253
rect 1006 248 1007 252
rect 1011 248 1012 252
rect 1006 247 1012 248
rect 1134 252 1140 253
rect 1134 248 1135 252
rect 1139 248 1140 252
rect 1134 247 1140 248
rect 1254 252 1260 253
rect 1254 248 1255 252
rect 1259 248 1260 252
rect 1254 247 1260 248
rect 1366 252 1372 253
rect 1366 248 1367 252
rect 1371 248 1372 252
rect 1366 247 1372 248
rect 1478 252 1484 253
rect 1478 248 1479 252
rect 1483 248 1484 252
rect 1478 247 1484 248
rect 1598 252 1604 253
rect 1598 248 1599 252
rect 1603 248 1604 252
rect 1894 252 1900 253
rect 1598 247 1604 248
rect 1830 249 1836 250
rect 110 244 116 245
rect 1830 245 1831 249
rect 1835 245 1836 249
rect 1830 244 1836 245
rect 1870 249 1876 250
rect 1870 245 1871 249
rect 1875 245 1876 249
rect 1894 248 1895 252
rect 1899 248 1900 252
rect 1894 247 1900 248
rect 1982 252 1988 253
rect 1982 248 1983 252
rect 1987 248 1988 252
rect 1982 247 1988 248
rect 2094 252 2100 253
rect 2094 248 2095 252
rect 2099 248 2100 252
rect 2094 247 2100 248
rect 2222 252 2228 253
rect 2222 248 2223 252
rect 2227 248 2228 252
rect 2222 247 2228 248
rect 2358 252 2364 253
rect 2358 248 2359 252
rect 2363 248 2364 252
rect 2358 247 2364 248
rect 2502 252 2508 253
rect 2502 248 2503 252
rect 2507 248 2508 252
rect 2502 247 2508 248
rect 2646 252 2652 253
rect 2646 248 2647 252
rect 2651 248 2652 252
rect 2646 247 2652 248
rect 2790 252 2796 253
rect 2790 248 2791 252
rect 2795 248 2796 252
rect 2790 247 2796 248
rect 2934 252 2940 253
rect 2934 248 2935 252
rect 2939 248 2940 252
rect 2934 247 2940 248
rect 3078 252 3084 253
rect 3078 248 3079 252
rect 3083 248 3084 252
rect 3078 247 3084 248
rect 3222 252 3228 253
rect 3222 248 3223 252
rect 3227 248 3228 252
rect 3222 247 3228 248
rect 3374 252 3380 253
rect 3374 248 3375 252
rect 3379 248 3380 252
rect 3374 247 3380 248
rect 3502 252 3508 253
rect 3502 248 3503 252
rect 3507 248 3508 252
rect 3502 247 3508 248
rect 3590 249 3596 250
rect 1870 244 1876 245
rect 3590 245 3591 249
rect 3595 245 3596 249
rect 3590 244 3596 245
rect 110 232 116 233
rect 110 228 111 232
rect 115 228 116 232
rect 110 227 116 228
rect 1830 232 1836 233
rect 1830 228 1831 232
rect 1835 228 1836 232
rect 1830 227 1836 228
rect 1870 232 1876 233
rect 1870 228 1871 232
rect 1875 228 1876 232
rect 1870 227 1876 228
rect 3590 232 3596 233
rect 3590 228 3591 232
rect 3595 228 3596 232
rect 3590 227 3596 228
rect 230 214 236 215
rect 230 210 231 214
rect 235 210 236 214
rect 230 209 236 210
rect 342 214 348 215
rect 342 210 343 214
rect 347 210 348 214
rect 342 209 348 210
rect 470 214 476 215
rect 470 210 471 214
rect 475 210 476 214
rect 470 209 476 210
rect 606 214 612 215
rect 606 210 607 214
rect 611 210 612 214
rect 606 209 612 210
rect 742 214 748 215
rect 742 210 743 214
rect 747 210 748 214
rect 742 209 748 210
rect 878 214 884 215
rect 878 210 879 214
rect 883 210 884 214
rect 878 209 884 210
rect 1014 214 1020 215
rect 1014 210 1015 214
rect 1019 210 1020 214
rect 1014 209 1020 210
rect 1142 214 1148 215
rect 1142 210 1143 214
rect 1147 210 1148 214
rect 1142 209 1148 210
rect 1262 214 1268 215
rect 1262 210 1263 214
rect 1267 210 1268 214
rect 1262 209 1268 210
rect 1374 214 1380 215
rect 1374 210 1375 214
rect 1379 210 1380 214
rect 1374 209 1380 210
rect 1486 214 1492 215
rect 1486 210 1487 214
rect 1491 210 1492 214
rect 1486 209 1492 210
rect 1606 214 1612 215
rect 1606 210 1607 214
rect 1611 210 1612 214
rect 1606 209 1612 210
rect 1902 214 1908 215
rect 1902 210 1903 214
rect 1907 210 1908 214
rect 1902 209 1908 210
rect 1990 214 1996 215
rect 1990 210 1991 214
rect 1995 210 1996 214
rect 1990 209 1996 210
rect 2102 214 2108 215
rect 2102 210 2103 214
rect 2107 210 2108 214
rect 2102 209 2108 210
rect 2230 214 2236 215
rect 2230 210 2231 214
rect 2235 210 2236 214
rect 2230 209 2236 210
rect 2366 214 2372 215
rect 2366 210 2367 214
rect 2371 210 2372 214
rect 2366 209 2372 210
rect 2510 214 2516 215
rect 2510 210 2511 214
rect 2515 210 2516 214
rect 2510 209 2516 210
rect 2654 214 2660 215
rect 2654 210 2655 214
rect 2659 210 2660 214
rect 2654 209 2660 210
rect 2798 214 2804 215
rect 2798 210 2799 214
rect 2803 210 2804 214
rect 2798 209 2804 210
rect 2942 214 2948 215
rect 2942 210 2943 214
rect 2947 210 2948 214
rect 2942 209 2948 210
rect 3086 214 3092 215
rect 3086 210 3087 214
rect 3091 210 3092 214
rect 3086 209 3092 210
rect 3230 214 3236 215
rect 3230 210 3231 214
rect 3235 210 3236 214
rect 3230 209 3236 210
rect 3382 214 3388 215
rect 3382 210 3383 214
rect 3387 210 3388 214
rect 3382 209 3388 210
rect 3510 214 3516 215
rect 3510 210 3511 214
rect 3515 210 3516 214
rect 3510 209 3516 210
rect 1902 170 1908 171
rect 1902 166 1903 170
rect 1907 166 1908 170
rect 1902 165 1908 166
rect 1982 170 1988 171
rect 1982 166 1983 170
rect 1987 166 1988 170
rect 1982 165 1988 166
rect 2086 170 2092 171
rect 2086 166 2087 170
rect 2091 166 2092 170
rect 2086 165 2092 166
rect 2206 170 2212 171
rect 2206 166 2207 170
rect 2211 166 2212 170
rect 2206 165 2212 166
rect 2334 170 2340 171
rect 2334 166 2335 170
rect 2339 166 2340 170
rect 2334 165 2340 166
rect 2462 170 2468 171
rect 2462 166 2463 170
rect 2467 166 2468 170
rect 2462 165 2468 166
rect 2582 170 2588 171
rect 2582 166 2583 170
rect 2587 166 2588 170
rect 2582 165 2588 166
rect 2702 170 2708 171
rect 2702 166 2703 170
rect 2707 166 2708 170
rect 2702 165 2708 166
rect 2814 170 2820 171
rect 2814 166 2815 170
rect 2819 166 2820 170
rect 2814 165 2820 166
rect 2918 170 2924 171
rect 2918 166 2919 170
rect 2923 166 2924 170
rect 2918 165 2924 166
rect 3014 170 3020 171
rect 3014 166 3015 170
rect 3019 166 3020 170
rect 3014 165 3020 166
rect 3110 170 3116 171
rect 3110 166 3111 170
rect 3115 166 3116 170
rect 3110 165 3116 166
rect 3206 170 3212 171
rect 3206 166 3207 170
rect 3211 166 3212 170
rect 3206 165 3212 166
rect 3302 170 3308 171
rect 3302 166 3303 170
rect 3307 166 3308 170
rect 3302 165 3308 166
rect 3398 170 3404 171
rect 3398 166 3399 170
rect 3403 166 3404 170
rect 3398 165 3404 166
rect 1870 152 1876 153
rect 158 150 164 151
rect 158 146 159 150
rect 163 146 164 150
rect 158 145 164 146
rect 238 150 244 151
rect 238 146 239 150
rect 243 146 244 150
rect 238 145 244 146
rect 318 150 324 151
rect 318 146 319 150
rect 323 146 324 150
rect 318 145 324 146
rect 398 150 404 151
rect 398 146 399 150
rect 403 146 404 150
rect 398 145 404 146
rect 478 150 484 151
rect 478 146 479 150
rect 483 146 484 150
rect 478 145 484 146
rect 558 150 564 151
rect 558 146 559 150
rect 563 146 564 150
rect 558 145 564 146
rect 646 150 652 151
rect 646 146 647 150
rect 651 146 652 150
rect 646 145 652 146
rect 734 150 740 151
rect 734 146 735 150
rect 739 146 740 150
rect 734 145 740 146
rect 822 150 828 151
rect 822 146 823 150
rect 827 146 828 150
rect 822 145 828 146
rect 910 150 916 151
rect 910 146 911 150
rect 915 146 916 150
rect 910 145 916 146
rect 998 150 1004 151
rect 998 146 999 150
rect 1003 146 1004 150
rect 998 145 1004 146
rect 1086 150 1092 151
rect 1086 146 1087 150
rect 1091 146 1092 150
rect 1086 145 1092 146
rect 1166 150 1172 151
rect 1166 146 1167 150
rect 1171 146 1172 150
rect 1166 145 1172 146
rect 1246 150 1252 151
rect 1246 146 1247 150
rect 1251 146 1252 150
rect 1246 145 1252 146
rect 1334 150 1340 151
rect 1334 146 1335 150
rect 1339 146 1340 150
rect 1334 145 1340 146
rect 1422 150 1428 151
rect 1422 146 1423 150
rect 1427 146 1428 150
rect 1422 145 1428 146
rect 1510 150 1516 151
rect 1510 146 1511 150
rect 1515 146 1516 150
rect 1510 145 1516 146
rect 1590 150 1596 151
rect 1590 146 1591 150
rect 1595 146 1596 150
rect 1590 145 1596 146
rect 1670 150 1676 151
rect 1670 146 1671 150
rect 1675 146 1676 150
rect 1670 145 1676 146
rect 1750 150 1756 151
rect 1750 146 1751 150
rect 1755 146 1756 150
rect 1870 148 1871 152
rect 1875 148 1876 152
rect 1870 147 1876 148
rect 3590 152 3596 153
rect 3590 148 3591 152
rect 3595 148 3596 152
rect 3590 147 3596 148
rect 1750 145 1756 146
rect 1870 135 1876 136
rect 110 132 116 133
rect 110 128 111 132
rect 115 128 116 132
rect 110 127 116 128
rect 1830 132 1836 133
rect 1830 128 1831 132
rect 1835 128 1836 132
rect 1870 131 1871 135
rect 1875 131 1876 135
rect 3590 135 3596 136
rect 1870 130 1876 131
rect 1894 132 1900 133
rect 1830 127 1836 128
rect 1894 128 1895 132
rect 1899 128 1900 132
rect 1894 127 1900 128
rect 1974 132 1980 133
rect 1974 128 1975 132
rect 1979 128 1980 132
rect 1974 127 1980 128
rect 2078 132 2084 133
rect 2078 128 2079 132
rect 2083 128 2084 132
rect 2078 127 2084 128
rect 2198 132 2204 133
rect 2198 128 2199 132
rect 2203 128 2204 132
rect 2198 127 2204 128
rect 2326 132 2332 133
rect 2326 128 2327 132
rect 2331 128 2332 132
rect 2326 127 2332 128
rect 2454 132 2460 133
rect 2454 128 2455 132
rect 2459 128 2460 132
rect 2454 127 2460 128
rect 2574 132 2580 133
rect 2574 128 2575 132
rect 2579 128 2580 132
rect 2574 127 2580 128
rect 2694 132 2700 133
rect 2694 128 2695 132
rect 2699 128 2700 132
rect 2694 127 2700 128
rect 2806 132 2812 133
rect 2806 128 2807 132
rect 2811 128 2812 132
rect 2806 127 2812 128
rect 2910 132 2916 133
rect 2910 128 2911 132
rect 2915 128 2916 132
rect 2910 127 2916 128
rect 3006 132 3012 133
rect 3006 128 3007 132
rect 3011 128 3012 132
rect 3006 127 3012 128
rect 3102 132 3108 133
rect 3102 128 3103 132
rect 3107 128 3108 132
rect 3102 127 3108 128
rect 3198 132 3204 133
rect 3198 128 3199 132
rect 3203 128 3204 132
rect 3198 127 3204 128
rect 3294 132 3300 133
rect 3294 128 3295 132
rect 3299 128 3300 132
rect 3294 127 3300 128
rect 3390 132 3396 133
rect 3390 128 3391 132
rect 3395 128 3396 132
rect 3590 131 3591 135
rect 3595 131 3596 135
rect 3590 130 3596 131
rect 3390 127 3396 128
rect 110 115 116 116
rect 110 111 111 115
rect 115 111 116 115
rect 1830 115 1836 116
rect 110 110 116 111
rect 150 112 156 113
rect 150 108 151 112
rect 155 108 156 112
rect 150 107 156 108
rect 230 112 236 113
rect 230 108 231 112
rect 235 108 236 112
rect 230 107 236 108
rect 310 112 316 113
rect 310 108 311 112
rect 315 108 316 112
rect 310 107 316 108
rect 390 112 396 113
rect 390 108 391 112
rect 395 108 396 112
rect 390 107 396 108
rect 470 112 476 113
rect 470 108 471 112
rect 475 108 476 112
rect 470 107 476 108
rect 550 112 556 113
rect 550 108 551 112
rect 555 108 556 112
rect 550 107 556 108
rect 638 112 644 113
rect 638 108 639 112
rect 643 108 644 112
rect 638 107 644 108
rect 726 112 732 113
rect 726 108 727 112
rect 731 108 732 112
rect 726 107 732 108
rect 814 112 820 113
rect 814 108 815 112
rect 819 108 820 112
rect 814 107 820 108
rect 902 112 908 113
rect 902 108 903 112
rect 907 108 908 112
rect 902 107 908 108
rect 990 112 996 113
rect 990 108 991 112
rect 995 108 996 112
rect 990 107 996 108
rect 1078 112 1084 113
rect 1078 108 1079 112
rect 1083 108 1084 112
rect 1078 107 1084 108
rect 1158 112 1164 113
rect 1158 108 1159 112
rect 1163 108 1164 112
rect 1158 107 1164 108
rect 1238 112 1244 113
rect 1238 108 1239 112
rect 1243 108 1244 112
rect 1238 107 1244 108
rect 1326 112 1332 113
rect 1326 108 1327 112
rect 1331 108 1332 112
rect 1326 107 1332 108
rect 1414 112 1420 113
rect 1414 108 1415 112
rect 1419 108 1420 112
rect 1414 107 1420 108
rect 1502 112 1508 113
rect 1502 108 1503 112
rect 1507 108 1508 112
rect 1502 107 1508 108
rect 1582 112 1588 113
rect 1582 108 1583 112
rect 1587 108 1588 112
rect 1582 107 1588 108
rect 1662 112 1668 113
rect 1662 108 1663 112
rect 1667 108 1668 112
rect 1662 107 1668 108
rect 1742 112 1748 113
rect 1742 108 1743 112
rect 1747 108 1748 112
rect 1830 111 1831 115
rect 1835 111 1836 115
rect 1830 110 1836 111
rect 1742 107 1748 108
<< m3c >>
rect 1871 3641 1875 3645
rect 2151 3644 2155 3648
rect 2439 3644 2443 3648
rect 2727 3644 2731 3648
rect 3015 3644 3019 3648
rect 3591 3641 3595 3645
rect 143 3622 147 3626
rect 239 3622 243 3626
rect 367 3622 371 3626
rect 503 3622 507 3626
rect 639 3622 643 3626
rect 775 3622 779 3626
rect 911 3622 915 3626
rect 1055 3622 1059 3626
rect 1199 3622 1203 3626
rect 1871 3624 1875 3628
rect 3591 3624 3595 3628
rect 111 3604 115 3608
rect 1831 3604 1835 3608
rect 2159 3606 2163 3610
rect 2447 3606 2451 3610
rect 2735 3606 2739 3610
rect 3023 3606 3027 3610
rect 111 3587 115 3591
rect 135 3584 139 3588
rect 231 3584 235 3588
rect 359 3584 363 3588
rect 495 3584 499 3588
rect 631 3584 635 3588
rect 767 3584 771 3588
rect 903 3584 907 3588
rect 1047 3584 1051 3588
rect 1191 3584 1195 3588
rect 1831 3587 1835 3591
rect 1903 3574 1907 3578
rect 1983 3574 1987 3578
rect 2071 3574 2075 3578
rect 2175 3574 2179 3578
rect 2295 3574 2299 3578
rect 2423 3574 2427 3578
rect 2559 3574 2563 3578
rect 2695 3574 2699 3578
rect 2831 3574 2835 3578
rect 2975 3574 2979 3578
rect 3119 3574 3123 3578
rect 3263 3574 3267 3578
rect 1871 3556 1875 3560
rect 3591 3556 3595 3560
rect 111 3537 115 3541
rect 183 3540 187 3544
rect 303 3540 307 3544
rect 415 3540 419 3544
rect 527 3540 531 3544
rect 631 3540 635 3544
rect 735 3540 739 3544
rect 831 3540 835 3544
rect 919 3540 923 3544
rect 1007 3540 1011 3544
rect 1095 3540 1099 3544
rect 1183 3540 1187 3544
rect 1271 3540 1275 3544
rect 1359 3540 1363 3544
rect 1447 3540 1451 3544
rect 1831 3537 1835 3541
rect 1871 3539 1875 3543
rect 1895 3536 1899 3540
rect 1975 3536 1979 3540
rect 2063 3536 2067 3540
rect 2167 3536 2171 3540
rect 2287 3536 2291 3540
rect 2415 3536 2419 3540
rect 2551 3536 2555 3540
rect 2687 3536 2691 3540
rect 2823 3536 2827 3540
rect 2967 3536 2971 3540
rect 3111 3536 3115 3540
rect 3255 3536 3259 3540
rect 3591 3539 3595 3543
rect 111 3520 115 3524
rect 1831 3520 1835 3524
rect 191 3502 195 3506
rect 311 3502 315 3506
rect 423 3502 427 3506
rect 535 3502 539 3506
rect 639 3502 643 3506
rect 743 3502 747 3506
rect 839 3502 843 3506
rect 927 3502 931 3506
rect 1015 3502 1019 3506
rect 1103 3502 1107 3506
rect 1191 3502 1195 3506
rect 1279 3502 1283 3506
rect 1367 3502 1371 3506
rect 1455 3502 1459 3506
rect 1871 3489 1875 3493
rect 1967 3492 1971 3496
rect 2151 3492 2155 3496
rect 2335 3492 2339 3496
rect 2511 3492 2515 3496
rect 2671 3492 2675 3496
rect 2823 3492 2827 3496
rect 2959 3492 2963 3496
rect 3079 3492 3083 3496
rect 3191 3492 3195 3496
rect 3303 3492 3307 3496
rect 3415 3492 3419 3496
rect 3503 3492 3507 3496
rect 3591 3489 3595 3493
rect 1871 3472 1875 3476
rect 3591 3472 3595 3476
rect 231 3462 235 3466
rect 367 3462 371 3466
rect 503 3462 507 3466
rect 623 3462 627 3466
rect 735 3462 739 3466
rect 839 3462 843 3466
rect 943 3462 947 3466
rect 1039 3462 1043 3466
rect 1135 3462 1139 3466
rect 1231 3462 1235 3466
rect 1327 3462 1331 3466
rect 1975 3454 1979 3458
rect 2159 3454 2163 3458
rect 2343 3454 2347 3458
rect 2519 3454 2523 3458
rect 2679 3454 2683 3458
rect 2831 3454 2835 3458
rect 2967 3454 2971 3458
rect 3087 3454 3091 3458
rect 3199 3454 3203 3458
rect 3311 3454 3315 3458
rect 3423 3454 3427 3458
rect 3511 3454 3515 3458
rect 111 3444 115 3448
rect 1831 3444 1835 3448
rect 111 3427 115 3431
rect 223 3424 227 3428
rect 359 3424 363 3428
rect 495 3424 499 3428
rect 615 3424 619 3428
rect 727 3424 731 3428
rect 831 3424 835 3428
rect 935 3424 939 3428
rect 1031 3424 1035 3428
rect 1127 3424 1131 3428
rect 1223 3424 1227 3428
rect 1319 3424 1323 3428
rect 1831 3427 1835 3431
rect 2007 3422 2011 3426
rect 2127 3422 2131 3426
rect 2255 3422 2259 3426
rect 2391 3422 2395 3426
rect 2535 3422 2539 3426
rect 2679 3422 2683 3426
rect 2831 3422 2835 3426
rect 2999 3422 3003 3426
rect 3167 3422 3171 3426
rect 3343 3422 3347 3426
rect 3511 3422 3515 3426
rect 1871 3404 1875 3408
rect 3591 3404 3595 3408
rect 1871 3387 1875 3391
rect 1999 3384 2003 3388
rect 2119 3384 2123 3388
rect 2247 3384 2251 3388
rect 2383 3384 2387 3388
rect 2527 3384 2531 3388
rect 2671 3384 2675 3388
rect 2823 3384 2827 3388
rect 2991 3384 2995 3388
rect 3159 3384 3163 3388
rect 3335 3384 3339 3388
rect 3503 3384 3507 3388
rect 3591 3387 3595 3391
rect 111 3373 115 3377
rect 215 3376 219 3380
rect 367 3376 371 3380
rect 511 3376 515 3380
rect 647 3376 651 3380
rect 775 3376 779 3380
rect 895 3376 899 3380
rect 1015 3376 1019 3380
rect 1127 3376 1131 3380
rect 1239 3376 1243 3380
rect 1351 3376 1355 3380
rect 1831 3373 1835 3377
rect 111 3356 115 3360
rect 1831 3356 1835 3360
rect 223 3338 227 3342
rect 375 3338 379 3342
rect 519 3338 523 3342
rect 655 3338 659 3342
rect 783 3338 787 3342
rect 903 3338 907 3342
rect 1023 3338 1027 3342
rect 1135 3338 1139 3342
rect 1247 3338 1251 3342
rect 1359 3338 1363 3342
rect 1871 3337 1875 3341
rect 2015 3340 2019 3344
rect 2151 3340 2155 3344
rect 2295 3340 2299 3344
rect 2439 3340 2443 3344
rect 2583 3340 2587 3344
rect 2727 3340 2731 3344
rect 2871 3340 2875 3344
rect 3023 3340 3027 3344
rect 3183 3340 3187 3344
rect 3351 3340 3355 3344
rect 3503 3340 3507 3344
rect 3591 3337 3595 3341
rect 1871 3320 1875 3324
rect 3591 3320 3595 3324
rect 207 3302 211 3306
rect 367 3302 371 3306
rect 519 3302 523 3306
rect 671 3302 675 3306
rect 815 3302 819 3306
rect 951 3302 955 3306
rect 1087 3302 1091 3306
rect 1215 3302 1219 3306
rect 1343 3302 1347 3306
rect 1471 3302 1475 3306
rect 2023 3302 2027 3306
rect 2159 3302 2163 3306
rect 2303 3302 2307 3306
rect 2447 3302 2451 3306
rect 2591 3302 2595 3306
rect 2735 3302 2739 3306
rect 2879 3302 2883 3306
rect 3031 3302 3035 3306
rect 3191 3302 3195 3306
rect 3359 3302 3363 3306
rect 3511 3302 3515 3306
rect 111 3284 115 3288
rect 1831 3284 1835 3288
rect 111 3267 115 3271
rect 199 3264 203 3268
rect 359 3264 363 3268
rect 511 3264 515 3268
rect 663 3264 667 3268
rect 807 3264 811 3268
rect 943 3264 947 3268
rect 1079 3264 1083 3268
rect 1207 3264 1211 3268
rect 1335 3264 1339 3268
rect 1463 3264 1467 3268
rect 1831 3267 1835 3271
rect 1927 3270 1931 3274
rect 2063 3270 2067 3274
rect 2191 3270 2195 3274
rect 2319 3270 2323 3274
rect 2447 3270 2451 3274
rect 2591 3270 2595 3274
rect 2743 3270 2747 3274
rect 2919 3270 2923 3274
rect 3111 3270 3115 3274
rect 3311 3270 3315 3274
rect 3511 3270 3515 3274
rect 1871 3252 1875 3256
rect 3591 3252 3595 3256
rect 1871 3235 1875 3239
rect 1919 3232 1923 3236
rect 2055 3232 2059 3236
rect 2183 3232 2187 3236
rect 2311 3232 2315 3236
rect 2439 3232 2443 3236
rect 2583 3232 2587 3236
rect 2735 3232 2739 3236
rect 2911 3232 2915 3236
rect 3103 3232 3107 3236
rect 3303 3232 3307 3236
rect 3503 3232 3507 3236
rect 3591 3235 3595 3239
rect 111 3217 115 3221
rect 135 3220 139 3224
rect 271 3220 275 3224
rect 415 3220 419 3224
rect 575 3220 579 3224
rect 735 3220 739 3224
rect 895 3220 899 3224
rect 1047 3220 1051 3224
rect 1191 3220 1195 3224
rect 1327 3220 1331 3224
rect 1463 3220 1467 3224
rect 1607 3220 1611 3224
rect 1831 3217 1835 3221
rect 111 3200 115 3204
rect 1831 3200 1835 3204
rect 143 3182 147 3186
rect 279 3182 283 3186
rect 423 3182 427 3186
rect 583 3182 587 3186
rect 743 3182 747 3186
rect 903 3182 907 3186
rect 1055 3182 1059 3186
rect 1199 3182 1203 3186
rect 1335 3182 1339 3186
rect 1471 3182 1475 3186
rect 1615 3182 1619 3186
rect 1871 3185 1875 3189
rect 1895 3188 1899 3192
rect 2007 3188 2011 3192
rect 2143 3188 2147 3192
rect 2295 3188 2299 3192
rect 2455 3188 2459 3192
rect 2623 3188 2627 3192
rect 2799 3188 2803 3192
rect 2975 3188 2979 3192
rect 3151 3188 3155 3192
rect 3327 3188 3331 3192
rect 3503 3188 3507 3192
rect 3591 3185 3595 3189
rect 1871 3168 1875 3172
rect 3591 3168 3595 3172
rect 1903 3150 1907 3154
rect 2015 3150 2019 3154
rect 2151 3150 2155 3154
rect 2303 3150 2307 3154
rect 2463 3150 2467 3154
rect 2631 3150 2635 3154
rect 2807 3150 2811 3154
rect 2983 3150 2987 3154
rect 3159 3150 3163 3154
rect 3335 3150 3339 3154
rect 3511 3150 3515 3154
rect 175 3142 179 3146
rect 319 3142 323 3146
rect 463 3142 467 3146
rect 607 3142 611 3146
rect 743 3142 747 3146
rect 871 3142 875 3146
rect 991 3142 995 3146
rect 1103 3142 1107 3146
rect 1207 3142 1211 3146
rect 1311 3142 1315 3146
rect 1407 3142 1411 3146
rect 1495 3142 1499 3146
rect 1583 3142 1587 3146
rect 1671 3142 1675 3146
rect 1751 3142 1755 3146
rect 111 3124 115 3128
rect 1831 3124 1835 3128
rect 1903 3118 1907 3122
rect 2071 3118 2075 3122
rect 2263 3118 2267 3122
rect 2455 3118 2459 3122
rect 2647 3118 2651 3122
rect 2831 3118 2835 3122
rect 3015 3118 3019 3122
rect 3199 3118 3203 3122
rect 3391 3118 3395 3122
rect 111 3107 115 3111
rect 167 3104 171 3108
rect 311 3104 315 3108
rect 455 3104 459 3108
rect 599 3104 603 3108
rect 735 3104 739 3108
rect 863 3104 867 3108
rect 983 3104 987 3108
rect 1095 3104 1099 3108
rect 1199 3104 1203 3108
rect 1303 3104 1307 3108
rect 1399 3104 1403 3108
rect 1487 3104 1491 3108
rect 1575 3104 1579 3108
rect 1663 3104 1667 3108
rect 1743 3104 1747 3108
rect 1831 3107 1835 3111
rect 1871 3100 1875 3104
rect 3591 3100 3595 3104
rect 1871 3083 1875 3087
rect 1895 3080 1899 3084
rect 2063 3080 2067 3084
rect 2255 3080 2259 3084
rect 2447 3080 2451 3084
rect 2639 3080 2643 3084
rect 2823 3080 2827 3084
rect 3007 3080 3011 3084
rect 3191 3080 3195 3084
rect 3383 3080 3387 3084
rect 3591 3083 3595 3087
rect 111 3045 115 3049
rect 135 3048 139 3052
rect 223 3048 227 3052
rect 327 3048 331 3052
rect 439 3048 443 3052
rect 551 3048 555 3052
rect 663 3048 667 3052
rect 1831 3045 1835 3049
rect 111 3028 115 3032
rect 1831 3028 1835 3032
rect 1871 3021 1875 3025
rect 2199 3024 2203 3028
rect 2335 3024 2339 3028
rect 2479 3024 2483 3028
rect 2623 3024 2627 3028
rect 2767 3024 2771 3028
rect 2903 3024 2907 3028
rect 3039 3024 3043 3028
rect 3183 3024 3187 3028
rect 3327 3024 3331 3028
rect 3591 3021 3595 3025
rect 143 3010 147 3014
rect 231 3010 235 3014
rect 335 3010 339 3014
rect 447 3010 451 3014
rect 559 3010 563 3014
rect 671 3010 675 3014
rect 1871 3004 1875 3008
rect 3591 3004 3595 3008
rect 2207 2986 2211 2990
rect 2343 2986 2347 2990
rect 2487 2986 2491 2990
rect 2631 2986 2635 2990
rect 2775 2986 2779 2990
rect 2911 2986 2915 2990
rect 3047 2986 3051 2990
rect 3191 2986 3195 2990
rect 3335 2986 3339 2990
rect 159 2966 163 2970
rect 319 2966 323 2970
rect 487 2966 491 2970
rect 647 2966 651 2970
rect 799 2966 803 2970
rect 943 2966 947 2970
rect 1079 2966 1083 2970
rect 1199 2966 1203 2970
rect 1311 2966 1315 2970
rect 1423 2966 1427 2970
rect 1535 2966 1539 2970
rect 1647 2966 1651 2970
rect 111 2948 115 2952
rect 1831 2948 1835 2952
rect 2127 2942 2131 2946
rect 2207 2942 2211 2946
rect 2287 2942 2291 2946
rect 2367 2942 2371 2946
rect 2447 2942 2451 2946
rect 2527 2942 2531 2946
rect 2607 2942 2611 2946
rect 2695 2942 2699 2946
rect 2791 2942 2795 2946
rect 2911 2942 2915 2946
rect 3039 2942 3043 2946
rect 3183 2942 3187 2946
rect 3335 2942 3339 2946
rect 3495 2942 3499 2946
rect 111 2931 115 2935
rect 151 2928 155 2932
rect 311 2928 315 2932
rect 479 2928 483 2932
rect 639 2928 643 2932
rect 791 2928 795 2932
rect 935 2928 939 2932
rect 1071 2928 1075 2932
rect 1191 2928 1195 2932
rect 1303 2928 1307 2932
rect 1415 2928 1419 2932
rect 1527 2928 1531 2932
rect 1639 2928 1643 2932
rect 1831 2931 1835 2935
rect 1871 2924 1875 2928
rect 3591 2924 3595 2928
rect 1871 2907 1875 2911
rect 2119 2904 2123 2908
rect 2199 2904 2203 2908
rect 2279 2904 2283 2908
rect 2359 2904 2363 2908
rect 2439 2904 2443 2908
rect 2519 2904 2523 2908
rect 2599 2904 2603 2908
rect 2687 2904 2691 2908
rect 2783 2904 2787 2908
rect 2903 2904 2907 2908
rect 3031 2904 3035 2908
rect 3175 2904 3179 2908
rect 3327 2904 3331 2908
rect 3487 2904 3491 2908
rect 3591 2907 3595 2911
rect 111 2881 115 2885
rect 151 2884 155 2888
rect 311 2884 315 2888
rect 471 2884 475 2888
rect 631 2884 635 2888
rect 783 2884 787 2888
rect 927 2884 931 2888
rect 1055 2884 1059 2888
rect 1175 2884 1179 2888
rect 1287 2884 1291 2888
rect 1391 2884 1395 2888
rect 1487 2884 1491 2888
rect 1591 2884 1595 2888
rect 1695 2884 1699 2888
rect 1831 2881 1835 2885
rect 111 2864 115 2868
rect 1831 2864 1835 2868
rect 1871 2857 1875 2861
rect 2047 2860 2051 2864
rect 2135 2860 2139 2864
rect 2239 2860 2243 2864
rect 2343 2860 2347 2864
rect 2463 2860 2467 2864
rect 2591 2860 2595 2864
rect 2727 2860 2731 2864
rect 2879 2860 2883 2864
rect 3031 2860 3035 2864
rect 3191 2860 3195 2864
rect 3359 2860 3363 2864
rect 3503 2860 3507 2864
rect 3591 2857 3595 2861
rect 159 2846 163 2850
rect 319 2846 323 2850
rect 479 2846 483 2850
rect 639 2846 643 2850
rect 791 2846 795 2850
rect 935 2846 939 2850
rect 1063 2846 1067 2850
rect 1183 2846 1187 2850
rect 1295 2846 1299 2850
rect 1399 2846 1403 2850
rect 1495 2846 1499 2850
rect 1599 2846 1603 2850
rect 1703 2846 1707 2850
rect 1871 2840 1875 2844
rect 3591 2840 3595 2844
rect 2055 2822 2059 2826
rect 2143 2822 2147 2826
rect 2247 2822 2251 2826
rect 2351 2822 2355 2826
rect 2471 2822 2475 2826
rect 2599 2822 2603 2826
rect 2735 2822 2739 2826
rect 2887 2822 2891 2826
rect 3039 2822 3043 2826
rect 3199 2822 3203 2826
rect 3367 2822 3371 2826
rect 3511 2822 3515 2826
rect 143 2810 147 2814
rect 247 2810 251 2814
rect 383 2810 387 2814
rect 535 2810 539 2814
rect 687 2810 691 2814
rect 847 2810 851 2814
rect 999 2810 1003 2814
rect 1143 2810 1147 2814
rect 1279 2810 1283 2814
rect 1407 2810 1411 2814
rect 1527 2810 1531 2814
rect 1647 2810 1651 2814
rect 1751 2810 1755 2814
rect 111 2792 115 2796
rect 1831 2792 1835 2796
rect 111 2775 115 2779
rect 135 2772 139 2776
rect 239 2772 243 2776
rect 375 2772 379 2776
rect 527 2772 531 2776
rect 679 2772 683 2776
rect 839 2772 843 2776
rect 991 2772 995 2776
rect 1135 2772 1139 2776
rect 1271 2772 1275 2776
rect 1399 2772 1403 2776
rect 1519 2772 1523 2776
rect 1639 2772 1643 2776
rect 1743 2772 1747 2776
rect 1831 2775 1835 2779
rect 1903 2778 1907 2782
rect 2015 2778 2019 2782
rect 2167 2778 2171 2782
rect 2327 2778 2331 2782
rect 2487 2778 2491 2782
rect 2639 2778 2643 2782
rect 2791 2778 2795 2782
rect 2943 2778 2947 2782
rect 3087 2778 3091 2782
rect 3231 2778 3235 2782
rect 3383 2778 3387 2782
rect 3511 2778 3515 2782
rect 1871 2760 1875 2764
rect 3591 2760 3595 2764
rect 1871 2743 1875 2747
rect 1895 2740 1899 2744
rect 2007 2740 2011 2744
rect 2159 2740 2163 2744
rect 2319 2740 2323 2744
rect 2479 2740 2483 2744
rect 2631 2740 2635 2744
rect 2783 2740 2787 2744
rect 2935 2740 2939 2744
rect 3079 2740 3083 2744
rect 3223 2740 3227 2744
rect 3375 2740 3379 2744
rect 3503 2740 3507 2744
rect 3591 2743 3595 2747
rect 111 2721 115 2725
rect 135 2724 139 2728
rect 231 2724 235 2728
rect 367 2724 371 2728
rect 511 2724 515 2728
rect 663 2724 667 2728
rect 815 2724 819 2728
rect 975 2724 979 2728
rect 1135 2724 1139 2728
rect 1287 2724 1291 2728
rect 1447 2724 1451 2728
rect 1607 2724 1611 2728
rect 1743 2724 1747 2728
rect 1831 2721 1835 2725
rect 111 2704 115 2708
rect 1831 2704 1835 2708
rect 1871 2693 1875 2697
rect 1895 2696 1899 2700
rect 2103 2696 2107 2700
rect 2327 2696 2331 2700
rect 2535 2696 2539 2700
rect 2735 2696 2739 2700
rect 2911 2696 2915 2700
rect 3071 2696 3075 2700
rect 3223 2696 3227 2700
rect 3375 2696 3379 2700
rect 3503 2696 3507 2700
rect 3591 2693 3595 2697
rect 143 2686 147 2690
rect 239 2686 243 2690
rect 375 2686 379 2690
rect 519 2686 523 2690
rect 671 2686 675 2690
rect 823 2686 827 2690
rect 983 2686 987 2690
rect 1143 2686 1147 2690
rect 1295 2686 1299 2690
rect 1455 2686 1459 2690
rect 1615 2686 1619 2690
rect 1751 2686 1755 2690
rect 1871 2676 1875 2680
rect 3591 2676 3595 2680
rect 1903 2658 1907 2662
rect 2111 2658 2115 2662
rect 2335 2658 2339 2662
rect 2543 2658 2547 2662
rect 2743 2658 2747 2662
rect 2919 2658 2923 2662
rect 3079 2658 3083 2662
rect 3231 2658 3235 2662
rect 3383 2658 3387 2662
rect 3511 2658 3515 2662
rect 143 2646 147 2650
rect 279 2646 283 2650
rect 447 2646 451 2650
rect 623 2646 627 2650
rect 791 2646 795 2650
rect 951 2646 955 2650
rect 1103 2646 1107 2650
rect 1247 2646 1251 2650
rect 1399 2646 1403 2650
rect 1551 2646 1555 2650
rect 111 2628 115 2632
rect 1831 2628 1835 2632
rect 1903 2618 1907 2622
rect 2055 2618 2059 2622
rect 2263 2618 2267 2622
rect 2495 2618 2499 2622
rect 2751 2618 2755 2622
rect 3015 2618 3019 2622
rect 3287 2618 3291 2622
rect 111 2611 115 2615
rect 135 2608 139 2612
rect 271 2608 275 2612
rect 439 2608 443 2612
rect 615 2608 619 2612
rect 783 2608 787 2612
rect 943 2608 947 2612
rect 1095 2608 1099 2612
rect 1239 2608 1243 2612
rect 1391 2608 1395 2612
rect 1543 2608 1547 2612
rect 1831 2611 1835 2615
rect 1871 2600 1875 2604
rect 3591 2600 3595 2604
rect 1871 2583 1875 2587
rect 1895 2580 1899 2584
rect 2047 2580 2051 2584
rect 2255 2580 2259 2584
rect 2487 2580 2491 2584
rect 2743 2580 2747 2584
rect 3007 2580 3011 2584
rect 3279 2580 3283 2584
rect 3591 2583 3595 2587
rect 111 2557 115 2561
rect 135 2560 139 2564
rect 223 2560 227 2564
rect 367 2560 371 2564
rect 527 2560 531 2564
rect 703 2560 707 2564
rect 879 2560 883 2564
rect 1047 2560 1051 2564
rect 1207 2560 1211 2564
rect 1359 2560 1363 2564
rect 1511 2560 1515 2564
rect 1671 2560 1675 2564
rect 1831 2557 1835 2561
rect 111 2540 115 2544
rect 1831 2540 1835 2544
rect 1871 2533 1875 2537
rect 1895 2536 1899 2540
rect 2007 2536 2011 2540
rect 2159 2536 2163 2540
rect 2319 2536 2323 2540
rect 2471 2536 2475 2540
rect 2623 2536 2627 2540
rect 2759 2536 2763 2540
rect 2887 2536 2891 2540
rect 3007 2536 3011 2540
rect 3119 2536 3123 2540
rect 3223 2536 3227 2540
rect 3319 2536 3323 2540
rect 3423 2536 3427 2540
rect 3503 2536 3507 2540
rect 3591 2533 3595 2537
rect 143 2522 147 2526
rect 231 2522 235 2526
rect 375 2522 379 2526
rect 535 2522 539 2526
rect 711 2522 715 2526
rect 887 2522 891 2526
rect 1055 2522 1059 2526
rect 1215 2522 1219 2526
rect 1367 2522 1371 2526
rect 1519 2522 1523 2526
rect 1679 2522 1683 2526
rect 1871 2516 1875 2520
rect 3591 2516 3595 2520
rect 1903 2498 1907 2502
rect 2015 2498 2019 2502
rect 2167 2498 2171 2502
rect 2327 2498 2331 2502
rect 2479 2498 2483 2502
rect 2631 2498 2635 2502
rect 2767 2498 2771 2502
rect 2895 2498 2899 2502
rect 3015 2498 3019 2502
rect 3127 2498 3131 2502
rect 3231 2498 3235 2502
rect 3327 2498 3331 2502
rect 3431 2498 3435 2502
rect 3511 2498 3515 2502
rect 143 2486 147 2490
rect 223 2486 227 2490
rect 303 2486 307 2490
rect 391 2486 395 2490
rect 511 2486 515 2490
rect 647 2486 651 2490
rect 783 2486 787 2490
rect 927 2486 931 2490
rect 1063 2486 1067 2490
rect 1191 2486 1195 2490
rect 1311 2486 1315 2490
rect 1431 2486 1435 2490
rect 1551 2486 1555 2490
rect 1671 2486 1675 2490
rect 111 2468 115 2472
rect 1831 2468 1835 2472
rect 1999 2458 2003 2462
rect 2127 2458 2131 2462
rect 2263 2458 2267 2462
rect 2407 2458 2411 2462
rect 2551 2458 2555 2462
rect 2703 2458 2707 2462
rect 2863 2458 2867 2462
rect 3023 2458 3027 2462
rect 3191 2458 3195 2462
rect 3359 2458 3363 2462
rect 3511 2458 3515 2462
rect 111 2451 115 2455
rect 135 2448 139 2452
rect 215 2448 219 2452
rect 295 2448 299 2452
rect 383 2448 387 2452
rect 503 2448 507 2452
rect 639 2448 643 2452
rect 775 2448 779 2452
rect 919 2448 923 2452
rect 1055 2448 1059 2452
rect 1183 2448 1187 2452
rect 1303 2448 1307 2452
rect 1423 2448 1427 2452
rect 1543 2448 1547 2452
rect 1663 2448 1667 2452
rect 1831 2451 1835 2455
rect 1871 2440 1875 2444
rect 3591 2440 3595 2444
rect 1871 2423 1875 2427
rect 1991 2420 1995 2424
rect 2119 2420 2123 2424
rect 2255 2420 2259 2424
rect 2399 2420 2403 2424
rect 2543 2420 2547 2424
rect 2695 2420 2699 2424
rect 2855 2420 2859 2424
rect 3015 2420 3019 2424
rect 3183 2420 3187 2424
rect 3351 2420 3355 2424
rect 3503 2420 3507 2424
rect 3591 2423 3595 2427
rect 111 2389 115 2393
rect 1063 2392 1067 2396
rect 1143 2392 1147 2396
rect 1223 2392 1227 2396
rect 1303 2392 1307 2396
rect 1383 2392 1387 2396
rect 1463 2392 1467 2396
rect 1831 2389 1835 2393
rect 111 2372 115 2376
rect 1831 2372 1835 2376
rect 1871 2369 1875 2373
rect 2143 2372 2147 2376
rect 2239 2372 2243 2376
rect 2343 2372 2347 2376
rect 2455 2372 2459 2376
rect 2575 2372 2579 2376
rect 2703 2372 2707 2376
rect 2847 2372 2851 2376
rect 3007 2372 3011 2376
rect 3175 2372 3179 2376
rect 3351 2372 3355 2376
rect 3503 2372 3507 2376
rect 3591 2369 3595 2373
rect 1071 2354 1075 2358
rect 1151 2354 1155 2358
rect 1231 2354 1235 2358
rect 1311 2354 1315 2358
rect 1391 2354 1395 2358
rect 1471 2354 1475 2358
rect 1871 2352 1875 2356
rect 3591 2352 3595 2356
rect 2151 2334 2155 2338
rect 2247 2334 2251 2338
rect 2351 2334 2355 2338
rect 2463 2334 2467 2338
rect 2583 2334 2587 2338
rect 2711 2334 2715 2338
rect 2855 2334 2859 2338
rect 3015 2334 3019 2338
rect 3183 2334 3187 2338
rect 3359 2334 3363 2338
rect 3511 2334 3515 2338
rect 359 2314 363 2318
rect 439 2314 443 2318
rect 519 2314 523 2318
rect 599 2314 603 2318
rect 679 2314 683 2318
rect 759 2314 763 2318
rect 839 2314 843 2318
rect 919 2314 923 2318
rect 999 2314 1003 2318
rect 1079 2314 1083 2318
rect 1159 2314 1163 2318
rect 1239 2314 1243 2318
rect 1319 2314 1323 2318
rect 111 2296 115 2300
rect 1831 2296 1835 2300
rect 2279 2298 2283 2302
rect 2359 2298 2363 2302
rect 2439 2298 2443 2302
rect 2519 2298 2523 2302
rect 2599 2298 2603 2302
rect 2679 2298 2683 2302
rect 2759 2298 2763 2302
rect 2847 2298 2851 2302
rect 2935 2298 2939 2302
rect 111 2279 115 2283
rect 351 2276 355 2280
rect 431 2276 435 2280
rect 511 2276 515 2280
rect 591 2276 595 2280
rect 671 2276 675 2280
rect 751 2276 755 2280
rect 831 2276 835 2280
rect 911 2276 915 2280
rect 991 2276 995 2280
rect 1071 2276 1075 2280
rect 1151 2276 1155 2280
rect 1231 2276 1235 2280
rect 1311 2276 1315 2280
rect 1831 2279 1835 2283
rect 1871 2280 1875 2284
rect 3591 2280 3595 2284
rect 1871 2263 1875 2267
rect 2271 2260 2275 2264
rect 2351 2260 2355 2264
rect 2431 2260 2435 2264
rect 2511 2260 2515 2264
rect 2591 2260 2595 2264
rect 2671 2260 2675 2264
rect 2751 2260 2755 2264
rect 2839 2260 2843 2264
rect 2927 2260 2931 2264
rect 3591 2263 3595 2267
rect 111 2229 115 2233
rect 375 2232 379 2236
rect 455 2232 459 2236
rect 535 2232 539 2236
rect 615 2232 619 2236
rect 695 2232 699 2236
rect 775 2232 779 2236
rect 855 2232 859 2236
rect 935 2232 939 2236
rect 1015 2232 1019 2236
rect 1095 2232 1099 2236
rect 1175 2232 1179 2236
rect 1255 2232 1259 2236
rect 1831 2229 1835 2233
rect 111 2212 115 2216
rect 1831 2212 1835 2216
rect 1871 2213 1875 2217
rect 2311 2216 2315 2220
rect 2399 2216 2403 2220
rect 2495 2216 2499 2220
rect 2599 2216 2603 2220
rect 2719 2216 2723 2220
rect 2855 2216 2859 2220
rect 3007 2216 3011 2220
rect 3175 2216 3179 2220
rect 3351 2216 3355 2220
rect 3503 2216 3507 2220
rect 3591 2213 3595 2217
rect 383 2194 387 2198
rect 463 2194 467 2198
rect 543 2194 547 2198
rect 623 2194 627 2198
rect 703 2194 707 2198
rect 783 2194 787 2198
rect 863 2194 867 2198
rect 943 2194 947 2198
rect 1023 2194 1027 2198
rect 1103 2194 1107 2198
rect 1183 2194 1187 2198
rect 1263 2194 1267 2198
rect 1871 2196 1875 2200
rect 3591 2196 3595 2200
rect 2319 2178 2323 2182
rect 2407 2178 2411 2182
rect 2503 2178 2507 2182
rect 2607 2178 2611 2182
rect 2727 2178 2731 2182
rect 2863 2178 2867 2182
rect 3015 2178 3019 2182
rect 3183 2178 3187 2182
rect 3359 2178 3363 2182
rect 3511 2178 3515 2182
rect 311 2150 315 2154
rect 407 2150 411 2154
rect 503 2150 507 2154
rect 599 2150 603 2154
rect 687 2150 691 2154
rect 775 2150 779 2154
rect 863 2150 867 2154
rect 951 2150 955 2154
rect 1039 2150 1043 2154
rect 1127 2150 1131 2154
rect 1223 2150 1227 2154
rect 1903 2142 1907 2146
rect 1983 2142 1987 2146
rect 2111 2142 2115 2146
rect 2247 2142 2251 2146
rect 2391 2142 2395 2146
rect 2543 2142 2547 2146
rect 2695 2142 2699 2146
rect 2847 2142 2851 2146
rect 3007 2142 3011 2146
rect 3175 2142 3179 2146
rect 3351 2142 3355 2146
rect 3511 2142 3515 2146
rect 111 2132 115 2136
rect 1831 2132 1835 2136
rect 1871 2124 1875 2128
rect 3591 2124 3595 2128
rect 111 2115 115 2119
rect 303 2112 307 2116
rect 399 2112 403 2116
rect 495 2112 499 2116
rect 591 2112 595 2116
rect 679 2112 683 2116
rect 767 2112 771 2116
rect 855 2112 859 2116
rect 943 2112 947 2116
rect 1031 2112 1035 2116
rect 1119 2112 1123 2116
rect 1215 2112 1219 2116
rect 1831 2115 1835 2119
rect 1871 2107 1875 2111
rect 1895 2104 1899 2108
rect 1975 2104 1979 2108
rect 2103 2104 2107 2108
rect 2239 2104 2243 2108
rect 2383 2104 2387 2108
rect 2535 2104 2539 2108
rect 2687 2104 2691 2108
rect 2839 2104 2843 2108
rect 2999 2104 3003 2108
rect 3167 2104 3171 2108
rect 3343 2104 3347 2108
rect 3503 2104 3507 2108
rect 3591 2107 3595 2111
rect 111 2053 115 2057
rect 207 2056 211 2060
rect 327 2056 331 2060
rect 447 2056 451 2060
rect 575 2056 579 2060
rect 703 2056 707 2060
rect 823 2056 827 2060
rect 943 2056 947 2060
rect 1063 2056 1067 2060
rect 1175 2056 1179 2060
rect 1279 2056 1283 2060
rect 1375 2056 1379 2060
rect 1471 2056 1475 2060
rect 1567 2056 1571 2060
rect 1663 2056 1667 2060
rect 1743 2056 1747 2060
rect 1831 2053 1835 2057
rect 1871 2049 1875 2053
rect 1967 2052 1971 2056
rect 2215 2052 2219 2056
rect 2447 2052 2451 2056
rect 2655 2052 2659 2056
rect 2839 2052 2843 2056
rect 2999 2052 3003 2056
rect 3143 2052 3147 2056
rect 3271 2052 3275 2056
rect 3399 2052 3403 2056
rect 3503 2052 3507 2056
rect 3591 2049 3595 2053
rect 111 2036 115 2040
rect 1831 2036 1835 2040
rect 1871 2032 1875 2036
rect 3591 2032 3595 2036
rect 215 2018 219 2022
rect 335 2018 339 2022
rect 455 2018 459 2022
rect 583 2018 587 2022
rect 711 2018 715 2022
rect 831 2018 835 2022
rect 951 2018 955 2022
rect 1071 2018 1075 2022
rect 1183 2018 1187 2022
rect 1287 2018 1291 2022
rect 1383 2018 1387 2022
rect 1479 2018 1483 2022
rect 1575 2018 1579 2022
rect 1671 2018 1675 2022
rect 1751 2018 1755 2022
rect 1975 2014 1979 2018
rect 2223 2014 2227 2018
rect 2455 2014 2459 2018
rect 2663 2014 2667 2018
rect 2847 2014 2851 2018
rect 3007 2014 3011 2018
rect 3151 2014 3155 2018
rect 3279 2014 3283 2018
rect 3407 2014 3411 2018
rect 3511 2014 3515 2018
rect 191 1982 195 1986
rect 351 1982 355 1986
rect 519 1982 523 1986
rect 687 1982 691 1986
rect 855 1982 859 1986
rect 1015 1982 1019 1986
rect 1167 1982 1171 1986
rect 1311 1982 1315 1986
rect 1447 1982 1451 1986
rect 1583 1982 1587 1986
rect 1719 1982 1723 1986
rect 1959 1982 1963 1986
rect 2079 1982 2083 1986
rect 2199 1982 2203 1986
rect 2319 1982 2323 1986
rect 2447 1982 2451 1986
rect 2583 1982 2587 1986
rect 2743 1982 2747 1986
rect 2919 1982 2923 1986
rect 3119 1982 3123 1986
rect 3327 1982 3331 1986
rect 3511 1982 3515 1986
rect 111 1964 115 1968
rect 1831 1964 1835 1968
rect 1871 1964 1875 1968
rect 3591 1964 3595 1968
rect 111 1947 115 1951
rect 183 1944 187 1948
rect 343 1944 347 1948
rect 511 1944 515 1948
rect 679 1944 683 1948
rect 847 1944 851 1948
rect 1007 1944 1011 1948
rect 1159 1944 1163 1948
rect 1303 1944 1307 1948
rect 1439 1944 1443 1948
rect 1575 1944 1579 1948
rect 1711 1944 1715 1948
rect 1831 1947 1835 1951
rect 1871 1947 1875 1951
rect 1951 1944 1955 1948
rect 2071 1944 2075 1948
rect 2191 1944 2195 1948
rect 2311 1944 2315 1948
rect 2439 1944 2443 1948
rect 2575 1944 2579 1948
rect 2735 1944 2739 1948
rect 2911 1944 2915 1948
rect 3111 1944 3115 1948
rect 3319 1944 3323 1948
rect 3503 1944 3507 1948
rect 3591 1947 3595 1951
rect 111 1893 115 1897
rect 135 1896 139 1900
rect 239 1896 243 1900
rect 375 1896 379 1900
rect 527 1896 531 1900
rect 687 1896 691 1900
rect 847 1896 851 1900
rect 1007 1896 1011 1900
rect 1159 1896 1163 1900
rect 1303 1896 1307 1900
rect 1455 1896 1459 1900
rect 1607 1896 1611 1900
rect 1831 1893 1835 1897
rect 1871 1889 1875 1893
rect 2063 1892 2067 1896
rect 2151 1892 2155 1896
rect 2239 1892 2243 1896
rect 2319 1892 2323 1896
rect 2399 1892 2403 1896
rect 2487 1892 2491 1896
rect 2575 1892 2579 1896
rect 2663 1892 2667 1896
rect 2759 1892 2763 1896
rect 2871 1892 2875 1896
rect 2991 1892 2995 1896
rect 3119 1892 3123 1896
rect 3247 1892 3251 1896
rect 3383 1892 3387 1896
rect 3503 1892 3507 1896
rect 3591 1889 3595 1893
rect 111 1876 115 1880
rect 1831 1876 1835 1880
rect 1871 1872 1875 1876
rect 3591 1872 3595 1876
rect 143 1858 147 1862
rect 247 1858 251 1862
rect 383 1858 387 1862
rect 535 1858 539 1862
rect 695 1858 699 1862
rect 855 1858 859 1862
rect 1015 1858 1019 1862
rect 1167 1858 1171 1862
rect 1311 1858 1315 1862
rect 1463 1858 1467 1862
rect 1615 1858 1619 1862
rect 2071 1854 2075 1858
rect 2159 1854 2163 1858
rect 2247 1854 2251 1858
rect 2327 1854 2331 1858
rect 2407 1854 2411 1858
rect 2495 1854 2499 1858
rect 2583 1854 2587 1858
rect 2671 1854 2675 1858
rect 2767 1854 2771 1858
rect 2879 1854 2883 1858
rect 2999 1854 3003 1858
rect 3127 1854 3131 1858
rect 3255 1854 3259 1858
rect 3391 1854 3395 1858
rect 3511 1854 3515 1858
rect 143 1822 147 1826
rect 287 1822 291 1826
rect 471 1822 475 1826
rect 663 1822 667 1826
rect 847 1822 851 1826
rect 1023 1822 1027 1826
rect 1191 1822 1195 1826
rect 1351 1822 1355 1826
rect 1511 1822 1515 1826
rect 1679 1822 1683 1826
rect 111 1804 115 1808
rect 1831 1804 1835 1808
rect 2095 1806 2099 1810
rect 2239 1806 2243 1810
rect 2399 1806 2403 1810
rect 2559 1806 2563 1810
rect 2719 1806 2723 1810
rect 2879 1806 2883 1810
rect 3031 1806 3035 1810
rect 3175 1806 3179 1810
rect 3319 1806 3323 1810
rect 3471 1806 3475 1810
rect 111 1787 115 1791
rect 135 1784 139 1788
rect 279 1784 283 1788
rect 463 1784 467 1788
rect 655 1784 659 1788
rect 839 1784 843 1788
rect 1015 1784 1019 1788
rect 1183 1784 1187 1788
rect 1343 1784 1347 1788
rect 1503 1784 1507 1788
rect 1671 1784 1675 1788
rect 1831 1787 1835 1791
rect 1871 1788 1875 1792
rect 3591 1788 3595 1792
rect 1871 1771 1875 1775
rect 2087 1768 2091 1772
rect 2231 1768 2235 1772
rect 2391 1768 2395 1772
rect 2551 1768 2555 1772
rect 2711 1768 2715 1772
rect 2871 1768 2875 1772
rect 3023 1768 3027 1772
rect 3167 1768 3171 1772
rect 3311 1768 3315 1772
rect 3463 1768 3467 1772
rect 3591 1771 3595 1775
rect 111 1729 115 1733
rect 135 1732 139 1736
rect 215 1732 219 1736
rect 343 1732 347 1736
rect 495 1732 499 1736
rect 663 1732 667 1736
rect 839 1732 843 1736
rect 1007 1732 1011 1736
rect 1167 1732 1171 1736
rect 1319 1732 1323 1736
rect 1463 1732 1467 1736
rect 1607 1732 1611 1736
rect 1743 1732 1747 1736
rect 1831 1729 1835 1733
rect 1871 1717 1875 1721
rect 2103 1720 2107 1724
rect 2239 1720 2243 1724
rect 2383 1720 2387 1724
rect 2527 1720 2531 1724
rect 2663 1720 2667 1724
rect 2799 1720 2803 1724
rect 2927 1720 2931 1724
rect 3047 1720 3051 1724
rect 3159 1720 3163 1724
rect 3271 1720 3275 1724
rect 3391 1720 3395 1724
rect 3503 1720 3507 1724
rect 111 1712 115 1716
rect 3591 1717 3595 1721
rect 1831 1712 1835 1716
rect 1871 1700 1875 1704
rect 3591 1700 3595 1704
rect 143 1694 147 1698
rect 223 1694 227 1698
rect 351 1694 355 1698
rect 503 1694 507 1698
rect 671 1694 675 1698
rect 847 1694 851 1698
rect 1015 1694 1019 1698
rect 1175 1694 1179 1698
rect 1327 1694 1331 1698
rect 1471 1694 1475 1698
rect 1615 1694 1619 1698
rect 1751 1694 1755 1698
rect 2111 1682 2115 1686
rect 2247 1682 2251 1686
rect 2391 1682 2395 1686
rect 2535 1682 2539 1686
rect 2671 1682 2675 1686
rect 2807 1682 2811 1686
rect 2935 1682 2939 1686
rect 3055 1682 3059 1686
rect 3167 1682 3171 1686
rect 3279 1682 3283 1686
rect 3399 1682 3403 1686
rect 3511 1682 3515 1686
rect 143 1658 147 1662
rect 295 1658 299 1662
rect 479 1658 483 1662
rect 671 1658 675 1662
rect 855 1658 859 1662
rect 1031 1658 1035 1662
rect 1199 1658 1203 1662
rect 1359 1658 1363 1662
rect 1519 1658 1523 1662
rect 1679 1658 1683 1662
rect 1967 1646 1971 1650
rect 2087 1646 2091 1650
rect 2215 1646 2219 1650
rect 2351 1646 2355 1650
rect 2495 1646 2499 1650
rect 2639 1646 2643 1650
rect 2783 1646 2787 1650
rect 2927 1646 2931 1650
rect 3071 1646 3075 1650
rect 3223 1646 3227 1650
rect 3375 1646 3379 1650
rect 3511 1646 3515 1650
rect 111 1640 115 1644
rect 1831 1640 1835 1644
rect 1871 1628 1875 1632
rect 111 1623 115 1627
rect 3591 1628 3595 1632
rect 135 1620 139 1624
rect 287 1620 291 1624
rect 471 1620 475 1624
rect 663 1620 667 1624
rect 847 1620 851 1624
rect 1023 1620 1027 1624
rect 1191 1620 1195 1624
rect 1351 1620 1355 1624
rect 1511 1620 1515 1624
rect 1671 1620 1675 1624
rect 1831 1623 1835 1627
rect 1871 1611 1875 1615
rect 1959 1608 1963 1612
rect 2079 1608 2083 1612
rect 2207 1608 2211 1612
rect 2343 1608 2347 1612
rect 2487 1608 2491 1612
rect 2631 1608 2635 1612
rect 2775 1608 2779 1612
rect 2919 1608 2923 1612
rect 3063 1608 3067 1612
rect 3215 1608 3219 1612
rect 3367 1608 3371 1612
rect 3503 1608 3507 1612
rect 3591 1611 3595 1615
rect 111 1573 115 1577
rect 159 1576 163 1580
rect 287 1576 291 1580
rect 423 1576 427 1580
rect 567 1576 571 1580
rect 711 1576 715 1580
rect 847 1576 851 1580
rect 983 1576 987 1580
rect 1119 1576 1123 1580
rect 1247 1576 1251 1580
rect 1375 1576 1379 1580
rect 1511 1576 1515 1580
rect 1831 1573 1835 1577
rect 111 1556 115 1560
rect 1831 1556 1835 1560
rect 1871 1553 1875 1557
rect 1895 1556 1899 1560
rect 2047 1556 2051 1560
rect 2207 1556 2211 1560
rect 2367 1556 2371 1560
rect 2527 1556 2531 1560
rect 2687 1556 2691 1560
rect 2839 1556 2843 1560
rect 2983 1556 2987 1560
rect 3119 1556 3123 1560
rect 3255 1556 3259 1560
rect 3391 1556 3395 1560
rect 3503 1556 3507 1560
rect 3591 1553 3595 1557
rect 167 1538 171 1542
rect 295 1538 299 1542
rect 431 1538 435 1542
rect 575 1538 579 1542
rect 719 1538 723 1542
rect 855 1538 859 1542
rect 991 1538 995 1542
rect 1127 1538 1131 1542
rect 1255 1538 1259 1542
rect 1383 1538 1387 1542
rect 1519 1538 1523 1542
rect 1871 1536 1875 1540
rect 3591 1536 3595 1540
rect 1903 1518 1907 1522
rect 2055 1518 2059 1522
rect 2215 1518 2219 1522
rect 2375 1518 2379 1522
rect 2535 1518 2539 1522
rect 2695 1518 2699 1522
rect 2847 1518 2851 1522
rect 2991 1518 2995 1522
rect 3127 1518 3131 1522
rect 3263 1518 3267 1522
rect 3399 1518 3403 1522
rect 3511 1518 3515 1522
rect 231 1502 235 1506
rect 375 1502 379 1506
rect 519 1502 523 1506
rect 655 1502 659 1506
rect 783 1502 787 1506
rect 903 1502 907 1506
rect 1015 1502 1019 1506
rect 1119 1502 1123 1506
rect 1215 1502 1219 1506
rect 1319 1502 1323 1506
rect 1423 1502 1427 1506
rect 111 1484 115 1488
rect 1831 1484 1835 1488
rect 1903 1478 1907 1482
rect 2007 1478 2011 1482
rect 2135 1478 2139 1482
rect 2271 1478 2275 1482
rect 2415 1478 2419 1482
rect 2567 1478 2571 1482
rect 2719 1478 2723 1482
rect 2879 1478 2883 1482
rect 3039 1478 3043 1482
rect 3199 1478 3203 1482
rect 3367 1478 3371 1482
rect 3511 1478 3515 1482
rect 111 1467 115 1471
rect 223 1464 227 1468
rect 367 1464 371 1468
rect 511 1464 515 1468
rect 647 1464 651 1468
rect 775 1464 779 1468
rect 895 1464 899 1468
rect 1007 1464 1011 1468
rect 1111 1464 1115 1468
rect 1207 1464 1211 1468
rect 1311 1464 1315 1468
rect 1415 1464 1419 1468
rect 1831 1467 1835 1471
rect 1871 1460 1875 1464
rect 3591 1460 3595 1464
rect 1871 1443 1875 1447
rect 1895 1440 1899 1444
rect 1999 1440 2003 1444
rect 2127 1440 2131 1444
rect 2263 1440 2267 1444
rect 2407 1440 2411 1444
rect 2559 1440 2563 1444
rect 2711 1440 2715 1444
rect 2871 1440 2875 1444
rect 3031 1440 3035 1444
rect 3191 1440 3195 1444
rect 3359 1440 3363 1444
rect 3503 1440 3507 1444
rect 3591 1443 3595 1447
rect 111 1409 115 1413
rect 255 1412 259 1416
rect 351 1412 355 1416
rect 447 1412 451 1416
rect 543 1412 547 1416
rect 631 1412 635 1416
rect 719 1412 723 1416
rect 807 1412 811 1416
rect 919 1412 923 1416
rect 1047 1412 1051 1416
rect 1207 1412 1211 1416
rect 1383 1412 1387 1416
rect 1575 1412 1579 1416
rect 1743 1412 1747 1416
rect 1831 1409 1835 1413
rect 111 1392 115 1396
rect 1831 1392 1835 1396
rect 1871 1393 1875 1397
rect 1895 1396 1899 1400
rect 2023 1396 2027 1400
rect 2167 1396 2171 1400
rect 2303 1396 2307 1400
rect 2431 1396 2435 1400
rect 2551 1396 2555 1400
rect 2671 1396 2675 1400
rect 2791 1396 2795 1400
rect 2911 1396 2915 1400
rect 3591 1393 3595 1397
rect 263 1374 267 1378
rect 359 1374 363 1378
rect 455 1374 459 1378
rect 551 1374 555 1378
rect 639 1374 643 1378
rect 727 1374 731 1378
rect 815 1374 819 1378
rect 927 1374 931 1378
rect 1055 1374 1059 1378
rect 1215 1374 1219 1378
rect 1391 1374 1395 1378
rect 1583 1374 1587 1378
rect 1751 1374 1755 1378
rect 1871 1376 1875 1380
rect 3591 1376 3595 1380
rect 1903 1358 1907 1362
rect 2031 1358 2035 1362
rect 2175 1358 2179 1362
rect 2311 1358 2315 1362
rect 2439 1358 2443 1362
rect 2559 1358 2563 1362
rect 2679 1358 2683 1362
rect 2799 1358 2803 1362
rect 2919 1358 2923 1362
rect 359 1342 363 1346
rect 471 1342 475 1346
rect 591 1342 595 1346
rect 727 1342 731 1346
rect 863 1342 867 1346
rect 1007 1342 1011 1346
rect 1143 1342 1147 1346
rect 1279 1342 1283 1346
rect 1407 1342 1411 1346
rect 1527 1342 1531 1346
rect 1647 1342 1651 1346
rect 1751 1342 1755 1346
rect 111 1324 115 1328
rect 1831 1324 1835 1328
rect 1927 1318 1931 1322
rect 2047 1318 2051 1322
rect 2183 1318 2187 1322
rect 2319 1318 2323 1322
rect 2455 1318 2459 1322
rect 2591 1318 2595 1322
rect 2719 1318 2723 1322
rect 2839 1318 2843 1322
rect 2951 1318 2955 1322
rect 3063 1318 3067 1322
rect 3183 1318 3187 1322
rect 111 1307 115 1311
rect 351 1304 355 1308
rect 463 1304 467 1308
rect 583 1304 587 1308
rect 719 1304 723 1308
rect 855 1304 859 1308
rect 999 1304 1003 1308
rect 1135 1304 1139 1308
rect 1271 1304 1275 1308
rect 1399 1304 1403 1308
rect 1519 1304 1523 1308
rect 1639 1304 1643 1308
rect 1743 1304 1747 1308
rect 1831 1307 1835 1311
rect 1871 1300 1875 1304
rect 3591 1300 3595 1304
rect 1871 1283 1875 1287
rect 1919 1280 1923 1284
rect 2039 1280 2043 1284
rect 2175 1280 2179 1284
rect 2311 1280 2315 1284
rect 2447 1280 2451 1284
rect 2583 1280 2587 1284
rect 2711 1280 2715 1284
rect 2831 1280 2835 1284
rect 2943 1280 2947 1284
rect 3055 1280 3059 1284
rect 3175 1280 3179 1284
rect 3591 1283 3595 1287
rect 111 1253 115 1257
rect 311 1256 315 1260
rect 415 1256 419 1260
rect 535 1256 539 1260
rect 671 1256 675 1260
rect 815 1256 819 1260
rect 959 1256 963 1260
rect 1103 1256 1107 1260
rect 1239 1256 1243 1260
rect 1375 1256 1379 1260
rect 1503 1256 1507 1260
rect 1631 1256 1635 1260
rect 1743 1256 1747 1260
rect 1831 1253 1835 1257
rect 111 1236 115 1240
rect 1831 1236 1835 1240
rect 1871 1225 1875 1229
rect 1895 1228 1899 1232
rect 2071 1228 2075 1232
rect 2271 1228 2275 1232
rect 2471 1228 2475 1232
rect 2663 1228 2667 1232
rect 2847 1228 2851 1232
rect 3023 1228 3027 1232
rect 3191 1228 3195 1232
rect 3359 1228 3363 1232
rect 3503 1228 3507 1232
rect 3591 1225 3595 1229
rect 319 1218 323 1222
rect 423 1218 427 1222
rect 543 1218 547 1222
rect 679 1218 683 1222
rect 823 1218 827 1222
rect 967 1218 971 1222
rect 1111 1218 1115 1222
rect 1247 1218 1251 1222
rect 1383 1218 1387 1222
rect 1511 1218 1515 1222
rect 1639 1218 1643 1222
rect 1751 1218 1755 1222
rect 1871 1208 1875 1212
rect 3591 1208 3595 1212
rect 239 1186 243 1190
rect 415 1186 419 1190
rect 591 1186 595 1190
rect 759 1186 763 1190
rect 927 1186 931 1190
rect 1079 1186 1083 1190
rect 1223 1186 1227 1190
rect 1367 1186 1371 1190
rect 1503 1186 1507 1190
rect 1639 1186 1643 1190
rect 1751 1186 1755 1190
rect 1903 1190 1907 1194
rect 2079 1190 2083 1194
rect 2279 1190 2283 1194
rect 2479 1190 2483 1194
rect 2671 1190 2675 1194
rect 2855 1190 2859 1194
rect 3031 1190 3035 1194
rect 3199 1190 3203 1194
rect 3367 1190 3371 1194
rect 3511 1190 3515 1194
rect 111 1168 115 1172
rect 1831 1168 1835 1172
rect 111 1151 115 1155
rect 231 1148 235 1152
rect 407 1148 411 1152
rect 583 1148 587 1152
rect 751 1148 755 1152
rect 919 1148 923 1152
rect 1071 1148 1075 1152
rect 1215 1148 1219 1152
rect 1359 1148 1363 1152
rect 1495 1148 1499 1152
rect 1631 1148 1635 1152
rect 1743 1148 1747 1152
rect 1831 1151 1835 1155
rect 1903 1154 1907 1158
rect 1983 1154 1987 1158
rect 2087 1154 2091 1158
rect 2215 1154 2219 1158
rect 2367 1154 2371 1158
rect 2527 1154 2531 1158
rect 2687 1154 2691 1158
rect 2839 1154 2843 1158
rect 2983 1154 2987 1158
rect 3127 1154 3131 1158
rect 3263 1154 3267 1158
rect 3399 1154 3403 1158
rect 3511 1154 3515 1158
rect 1871 1136 1875 1140
rect 3591 1136 3595 1140
rect 1871 1119 1875 1123
rect 1895 1116 1899 1120
rect 1975 1116 1979 1120
rect 2079 1116 2083 1120
rect 2207 1116 2211 1120
rect 2359 1116 2363 1120
rect 2519 1116 2523 1120
rect 2679 1116 2683 1120
rect 2831 1116 2835 1120
rect 2975 1116 2979 1120
rect 3119 1116 3123 1120
rect 3255 1116 3259 1120
rect 3391 1116 3395 1120
rect 3503 1116 3507 1120
rect 3591 1119 3595 1123
rect 111 1097 115 1101
rect 143 1100 147 1104
rect 279 1100 283 1104
rect 423 1100 427 1104
rect 567 1100 571 1104
rect 711 1100 715 1104
rect 847 1100 851 1104
rect 975 1100 979 1104
rect 1103 1100 1107 1104
rect 1223 1100 1227 1104
rect 1343 1100 1347 1104
rect 1471 1100 1475 1104
rect 1831 1097 1835 1101
rect 111 1080 115 1084
rect 1831 1080 1835 1084
rect 151 1062 155 1066
rect 287 1062 291 1066
rect 431 1062 435 1066
rect 575 1062 579 1066
rect 719 1062 723 1066
rect 855 1062 859 1066
rect 983 1062 987 1066
rect 1111 1062 1115 1066
rect 1231 1062 1235 1066
rect 1351 1062 1355 1066
rect 1479 1062 1483 1066
rect 1871 1061 1875 1065
rect 2167 1064 2171 1068
rect 2255 1064 2259 1068
rect 2359 1064 2363 1068
rect 2479 1064 2483 1068
rect 2607 1064 2611 1068
rect 2751 1064 2755 1068
rect 2895 1064 2899 1068
rect 3047 1064 3051 1068
rect 3207 1064 3211 1068
rect 3367 1064 3371 1068
rect 3503 1064 3507 1068
rect 3591 1061 3595 1065
rect 1871 1044 1875 1048
rect 3591 1044 3595 1048
rect 143 1022 147 1026
rect 263 1022 267 1026
rect 407 1022 411 1026
rect 551 1022 555 1026
rect 687 1022 691 1026
rect 807 1022 811 1026
rect 927 1022 931 1026
rect 1039 1022 1043 1026
rect 1143 1022 1147 1026
rect 1247 1022 1251 1026
rect 1359 1022 1363 1026
rect 2175 1026 2179 1030
rect 2263 1026 2267 1030
rect 2367 1026 2371 1030
rect 2487 1026 2491 1030
rect 2615 1026 2619 1030
rect 2759 1026 2763 1030
rect 2903 1026 2907 1030
rect 3055 1026 3059 1030
rect 3215 1026 3219 1030
rect 3375 1026 3379 1030
rect 3511 1026 3515 1030
rect 111 1004 115 1008
rect 1831 1004 1835 1008
rect 2303 994 2307 998
rect 2383 994 2387 998
rect 2471 994 2475 998
rect 2567 994 2571 998
rect 2671 994 2675 998
rect 2783 994 2787 998
rect 2911 994 2915 998
rect 3055 994 3059 998
rect 3207 994 3211 998
rect 3367 994 3371 998
rect 3511 994 3515 998
rect 111 987 115 991
rect 135 984 139 988
rect 255 984 259 988
rect 399 984 403 988
rect 543 984 547 988
rect 679 984 683 988
rect 799 984 803 988
rect 919 984 923 988
rect 1031 984 1035 988
rect 1135 984 1139 988
rect 1239 984 1243 988
rect 1351 984 1355 988
rect 1831 987 1835 991
rect 1871 976 1875 980
rect 3591 976 3595 980
rect 1871 959 1875 963
rect 2295 956 2299 960
rect 2375 956 2379 960
rect 2463 956 2467 960
rect 2559 956 2563 960
rect 2663 956 2667 960
rect 2775 956 2779 960
rect 2903 956 2907 960
rect 3047 956 3051 960
rect 3199 956 3203 960
rect 3359 956 3363 960
rect 3503 956 3507 960
rect 3591 959 3595 963
rect 111 929 115 933
rect 135 932 139 936
rect 215 932 219 936
rect 327 932 331 936
rect 447 932 451 936
rect 567 932 571 936
rect 687 932 691 936
rect 799 932 803 936
rect 911 932 915 936
rect 1015 932 1019 936
rect 1119 932 1123 936
rect 1223 932 1227 936
rect 1327 932 1331 936
rect 1831 929 1835 933
rect 111 912 115 916
rect 1831 912 1835 916
rect 1871 901 1875 905
rect 2279 904 2283 908
rect 2359 904 2363 908
rect 2439 904 2443 908
rect 2519 904 2523 908
rect 2607 904 2611 908
rect 2703 904 2707 908
rect 2807 904 2811 908
rect 2911 904 2915 908
rect 3015 904 3019 908
rect 3111 904 3115 908
rect 3215 904 3219 908
rect 3319 904 3323 908
rect 3423 904 3427 908
rect 3503 904 3507 908
rect 3591 901 3595 905
rect 143 894 147 898
rect 223 894 227 898
rect 335 894 339 898
rect 455 894 459 898
rect 575 894 579 898
rect 695 894 699 898
rect 807 894 811 898
rect 919 894 923 898
rect 1023 894 1027 898
rect 1127 894 1131 898
rect 1231 894 1235 898
rect 1335 894 1339 898
rect 1871 884 1875 888
rect 3591 884 3595 888
rect 2287 866 2291 870
rect 2367 866 2371 870
rect 2447 866 2451 870
rect 2527 866 2531 870
rect 2615 866 2619 870
rect 2711 866 2715 870
rect 2815 866 2819 870
rect 2919 866 2923 870
rect 3023 866 3027 870
rect 3119 866 3123 870
rect 3223 866 3227 870
rect 3327 866 3331 870
rect 3431 866 3435 870
rect 3511 866 3515 870
rect 143 854 147 858
rect 255 854 259 858
rect 399 854 403 858
rect 559 854 563 858
rect 719 854 723 858
rect 871 854 875 858
rect 1015 854 1019 858
rect 1151 854 1155 858
rect 1279 854 1283 858
rect 1399 854 1403 858
rect 1519 854 1523 858
rect 1647 854 1651 858
rect 111 836 115 840
rect 1831 836 1835 840
rect 111 819 115 823
rect 135 816 139 820
rect 247 816 251 820
rect 391 816 395 820
rect 551 816 555 820
rect 711 816 715 820
rect 863 816 867 820
rect 1007 816 1011 820
rect 1143 816 1147 820
rect 1271 816 1275 820
rect 1391 816 1395 820
rect 1511 816 1515 820
rect 1639 816 1643 820
rect 1831 819 1835 823
rect 2167 822 2171 826
rect 2247 822 2251 826
rect 2327 822 2331 826
rect 2423 822 2427 826
rect 2535 822 2539 826
rect 2655 822 2659 826
rect 2783 822 2787 826
rect 2911 822 2915 826
rect 3039 822 3043 826
rect 3159 822 3163 826
rect 3279 822 3283 826
rect 3407 822 3411 826
rect 3511 822 3515 826
rect 1871 804 1875 808
rect 3591 804 3595 808
rect 1871 787 1875 791
rect 2159 784 2163 788
rect 2239 784 2243 788
rect 2319 784 2323 788
rect 2415 784 2419 788
rect 2527 784 2531 788
rect 2647 784 2651 788
rect 2775 784 2779 788
rect 2903 784 2907 788
rect 3031 784 3035 788
rect 3151 784 3155 788
rect 3271 784 3275 788
rect 3399 784 3403 788
rect 3503 784 3507 788
rect 3591 787 3595 791
rect 111 757 115 761
rect 135 760 139 764
rect 263 760 267 764
rect 431 760 435 764
rect 607 760 611 764
rect 783 760 787 764
rect 951 760 955 764
rect 1103 760 1107 764
rect 1247 760 1251 764
rect 1383 760 1387 764
rect 1511 760 1515 764
rect 1639 760 1643 764
rect 1743 760 1747 764
rect 1831 757 1835 761
rect 111 740 115 744
rect 1831 740 1835 744
rect 1871 729 1875 733
rect 1895 732 1899 736
rect 1975 732 1979 736
rect 2071 732 2075 736
rect 2183 732 2187 736
rect 2311 732 2315 736
rect 2447 732 2451 736
rect 2591 732 2595 736
rect 2743 732 2747 736
rect 2895 732 2899 736
rect 3047 732 3051 736
rect 3199 732 3203 736
rect 3359 732 3363 736
rect 3503 732 3507 736
rect 3591 729 3595 733
rect 143 722 147 726
rect 271 722 275 726
rect 439 722 443 726
rect 615 722 619 726
rect 791 722 795 726
rect 959 722 963 726
rect 1111 722 1115 726
rect 1255 722 1259 726
rect 1391 722 1395 726
rect 1519 722 1523 726
rect 1647 722 1651 726
rect 1751 722 1755 726
rect 1871 712 1875 716
rect 3591 712 3595 716
rect 1903 694 1907 698
rect 1983 694 1987 698
rect 2079 694 2083 698
rect 2191 694 2195 698
rect 2319 694 2323 698
rect 2455 694 2459 698
rect 2599 694 2603 698
rect 2751 694 2755 698
rect 2903 694 2907 698
rect 3055 694 3059 698
rect 3207 694 3211 698
rect 3367 694 3371 698
rect 3511 694 3515 698
rect 295 678 299 682
rect 407 678 411 682
rect 527 678 531 682
rect 655 678 659 682
rect 783 678 787 682
rect 903 678 907 682
rect 1023 678 1027 682
rect 1135 678 1139 682
rect 1247 678 1251 682
rect 1351 678 1355 682
rect 1455 678 1459 682
rect 1559 678 1563 682
rect 1663 678 1667 682
rect 1751 678 1755 682
rect 111 660 115 664
rect 1831 660 1835 664
rect 1903 658 1907 662
rect 2095 658 2099 662
rect 2295 658 2299 662
rect 2479 658 2483 662
rect 2655 658 2659 662
rect 2831 658 2835 662
rect 3007 658 3011 662
rect 3183 658 3187 662
rect 3359 658 3363 662
rect 3511 658 3515 662
rect 111 643 115 647
rect 287 640 291 644
rect 399 640 403 644
rect 519 640 523 644
rect 647 640 651 644
rect 775 640 779 644
rect 895 640 899 644
rect 1015 640 1019 644
rect 1127 640 1131 644
rect 1239 640 1243 644
rect 1343 640 1347 644
rect 1447 640 1451 644
rect 1551 640 1555 644
rect 1655 640 1659 644
rect 1743 640 1747 644
rect 1831 643 1835 647
rect 1871 640 1875 644
rect 3591 640 3595 644
rect 1871 623 1875 627
rect 1895 620 1899 624
rect 2087 620 2091 624
rect 2287 620 2291 624
rect 2471 620 2475 624
rect 2647 620 2651 624
rect 2823 620 2827 624
rect 2999 620 3003 624
rect 3175 620 3179 624
rect 3351 620 3355 624
rect 3503 620 3507 624
rect 3591 623 3595 627
rect 111 589 115 593
rect 311 592 315 596
rect 391 592 395 596
rect 471 592 475 596
rect 559 592 563 596
rect 647 592 651 596
rect 735 592 739 596
rect 823 592 827 596
rect 911 592 915 596
rect 999 592 1003 596
rect 1087 592 1091 596
rect 1175 592 1179 596
rect 1263 592 1267 596
rect 1831 589 1835 593
rect 111 572 115 576
rect 1831 572 1835 576
rect 1871 569 1875 573
rect 1895 572 1899 576
rect 1975 572 1979 576
rect 2087 572 2091 576
rect 2215 572 2219 576
rect 2351 572 2355 576
rect 2495 572 2499 576
rect 2647 572 2651 576
rect 2807 572 2811 576
rect 2975 572 2979 576
rect 3151 572 3155 576
rect 3335 572 3339 576
rect 3503 572 3507 576
rect 3591 569 3595 573
rect 319 554 323 558
rect 399 554 403 558
rect 479 554 483 558
rect 567 554 571 558
rect 655 554 659 558
rect 743 554 747 558
rect 831 554 835 558
rect 919 554 923 558
rect 1007 554 1011 558
rect 1095 554 1099 558
rect 1183 554 1187 558
rect 1271 554 1275 558
rect 1871 552 1875 556
rect 3591 552 3595 556
rect 1903 534 1907 538
rect 1983 534 1987 538
rect 2095 534 2099 538
rect 2223 534 2227 538
rect 2359 534 2363 538
rect 2503 534 2507 538
rect 2655 534 2659 538
rect 2815 534 2819 538
rect 2983 534 2987 538
rect 3159 534 3163 538
rect 3343 534 3347 538
rect 3511 534 3515 538
rect 239 510 243 514
rect 343 510 347 514
rect 439 510 443 514
rect 535 510 539 514
rect 631 510 635 514
rect 719 510 723 514
rect 807 510 811 514
rect 895 510 899 514
rect 983 510 987 514
rect 1071 510 1075 514
rect 1159 510 1163 514
rect 1247 510 1251 514
rect 2151 502 2155 506
rect 2231 502 2235 506
rect 2327 502 2331 506
rect 2431 502 2435 506
rect 2551 502 2555 506
rect 2687 502 2691 506
rect 2839 502 2843 506
rect 2999 502 3003 506
rect 3175 502 3179 506
rect 3351 502 3355 506
rect 3511 502 3515 506
rect 111 492 115 496
rect 1831 492 1835 496
rect 1871 484 1875 488
rect 3591 484 3595 488
rect 111 475 115 479
rect 231 472 235 476
rect 335 472 339 476
rect 431 472 435 476
rect 527 472 531 476
rect 623 472 627 476
rect 711 472 715 476
rect 799 472 803 476
rect 887 472 891 476
rect 975 472 979 476
rect 1063 472 1067 476
rect 1151 472 1155 476
rect 1239 472 1243 476
rect 1831 475 1835 479
rect 1871 467 1875 471
rect 2143 464 2147 468
rect 2223 464 2227 468
rect 2319 464 2323 468
rect 2423 464 2427 468
rect 2543 464 2547 468
rect 2679 464 2683 468
rect 2831 464 2835 468
rect 2991 464 2995 468
rect 3167 464 3171 468
rect 3343 464 3347 468
rect 3503 464 3507 468
rect 3591 467 3595 471
rect 111 417 115 421
rect 135 420 139 424
rect 247 420 251 424
rect 375 420 379 424
rect 495 420 499 424
rect 607 420 611 424
rect 719 420 723 424
rect 823 420 827 424
rect 919 420 923 424
rect 1007 420 1011 424
rect 1103 420 1107 424
rect 1199 420 1203 424
rect 1295 420 1299 424
rect 1831 417 1835 421
rect 1871 413 1875 417
rect 2335 416 2339 420
rect 2415 416 2419 420
rect 2495 416 2499 420
rect 2583 416 2587 420
rect 2687 416 2691 420
rect 2799 416 2803 420
rect 2927 416 2931 420
rect 3071 416 3075 420
rect 3215 416 3219 420
rect 3367 416 3371 420
rect 3503 416 3507 420
rect 3591 413 3595 417
rect 111 400 115 404
rect 1831 400 1835 404
rect 1871 396 1875 400
rect 3591 396 3595 400
rect 143 382 147 386
rect 255 382 259 386
rect 383 382 387 386
rect 503 382 507 386
rect 615 382 619 386
rect 727 382 731 386
rect 831 382 835 386
rect 927 382 931 386
rect 1015 382 1019 386
rect 1111 382 1115 386
rect 1207 382 1211 386
rect 1303 382 1307 386
rect 2343 378 2347 382
rect 2423 378 2427 382
rect 2503 378 2507 382
rect 2591 378 2595 382
rect 2695 378 2699 382
rect 2807 378 2811 382
rect 2935 378 2939 382
rect 3079 378 3083 382
rect 3223 378 3227 382
rect 3375 378 3379 382
rect 3511 378 3515 382
rect 143 338 147 342
rect 247 338 251 342
rect 375 338 379 342
rect 511 338 515 342
rect 647 338 651 342
rect 775 338 779 342
rect 895 338 899 342
rect 1007 338 1011 342
rect 1119 338 1123 342
rect 1223 338 1227 342
rect 1327 338 1331 342
rect 1439 338 1443 342
rect 2079 338 2083 342
rect 2167 338 2171 342
rect 2263 338 2267 342
rect 2375 338 2379 342
rect 2503 338 2507 342
rect 2639 338 2643 342
rect 2775 338 2779 342
rect 2911 338 2915 342
rect 3039 338 3043 342
rect 3167 338 3171 342
rect 3287 338 3291 342
rect 3407 338 3411 342
rect 3511 338 3515 342
rect 111 320 115 324
rect 1831 320 1835 324
rect 1871 320 1875 324
rect 3591 320 3595 324
rect 111 303 115 307
rect 135 300 139 304
rect 239 300 243 304
rect 367 300 371 304
rect 503 300 507 304
rect 639 300 643 304
rect 767 300 771 304
rect 887 300 891 304
rect 999 300 1003 304
rect 1111 300 1115 304
rect 1215 300 1219 304
rect 1319 300 1323 304
rect 1431 300 1435 304
rect 1831 303 1835 307
rect 1871 303 1875 307
rect 2071 300 2075 304
rect 2159 300 2163 304
rect 2255 300 2259 304
rect 2367 300 2371 304
rect 2495 300 2499 304
rect 2631 300 2635 304
rect 2767 300 2771 304
rect 2903 300 2907 304
rect 3031 300 3035 304
rect 3159 300 3163 304
rect 3279 300 3283 304
rect 3399 300 3403 304
rect 3503 300 3507 304
rect 3591 303 3595 307
rect 111 245 115 249
rect 223 248 227 252
rect 335 248 339 252
rect 463 248 467 252
rect 599 248 603 252
rect 735 248 739 252
rect 871 248 875 252
rect 1007 248 1011 252
rect 1135 248 1139 252
rect 1255 248 1259 252
rect 1367 248 1371 252
rect 1479 248 1483 252
rect 1599 248 1603 252
rect 1831 245 1835 249
rect 1871 245 1875 249
rect 1895 248 1899 252
rect 1983 248 1987 252
rect 2095 248 2099 252
rect 2223 248 2227 252
rect 2359 248 2363 252
rect 2503 248 2507 252
rect 2647 248 2651 252
rect 2791 248 2795 252
rect 2935 248 2939 252
rect 3079 248 3083 252
rect 3223 248 3227 252
rect 3375 248 3379 252
rect 3503 248 3507 252
rect 3591 245 3595 249
rect 111 228 115 232
rect 1831 228 1835 232
rect 1871 228 1875 232
rect 3591 228 3595 232
rect 231 210 235 214
rect 343 210 347 214
rect 471 210 475 214
rect 607 210 611 214
rect 743 210 747 214
rect 879 210 883 214
rect 1015 210 1019 214
rect 1143 210 1147 214
rect 1263 210 1267 214
rect 1375 210 1379 214
rect 1487 210 1491 214
rect 1607 210 1611 214
rect 1903 210 1907 214
rect 1991 210 1995 214
rect 2103 210 2107 214
rect 2231 210 2235 214
rect 2367 210 2371 214
rect 2511 210 2515 214
rect 2655 210 2659 214
rect 2799 210 2803 214
rect 2943 210 2947 214
rect 3087 210 3091 214
rect 3231 210 3235 214
rect 3383 210 3387 214
rect 3511 210 3515 214
rect 1903 166 1907 170
rect 1983 166 1987 170
rect 2087 166 2091 170
rect 2207 166 2211 170
rect 2335 166 2339 170
rect 2463 166 2467 170
rect 2583 166 2587 170
rect 2703 166 2707 170
rect 2815 166 2819 170
rect 2919 166 2923 170
rect 3015 166 3019 170
rect 3111 166 3115 170
rect 3207 166 3211 170
rect 3303 166 3307 170
rect 3399 166 3403 170
rect 159 146 163 150
rect 239 146 243 150
rect 319 146 323 150
rect 399 146 403 150
rect 479 146 483 150
rect 559 146 563 150
rect 647 146 651 150
rect 735 146 739 150
rect 823 146 827 150
rect 911 146 915 150
rect 999 146 1003 150
rect 1087 146 1091 150
rect 1167 146 1171 150
rect 1247 146 1251 150
rect 1335 146 1339 150
rect 1423 146 1427 150
rect 1511 146 1515 150
rect 1591 146 1595 150
rect 1671 146 1675 150
rect 1751 146 1755 150
rect 1871 148 1875 152
rect 3591 148 3595 152
rect 111 128 115 132
rect 1831 128 1835 132
rect 1871 131 1875 135
rect 1895 128 1899 132
rect 1975 128 1979 132
rect 2079 128 2083 132
rect 2199 128 2203 132
rect 2327 128 2331 132
rect 2455 128 2459 132
rect 2575 128 2579 132
rect 2695 128 2699 132
rect 2807 128 2811 132
rect 2911 128 2915 132
rect 3007 128 3011 132
rect 3103 128 3107 132
rect 3199 128 3203 132
rect 3295 128 3299 132
rect 3391 128 3395 132
rect 3591 131 3595 135
rect 111 111 115 115
rect 151 108 155 112
rect 231 108 235 112
rect 311 108 315 112
rect 391 108 395 112
rect 471 108 475 112
rect 551 108 555 112
rect 639 108 643 112
rect 727 108 731 112
rect 815 108 819 112
rect 903 108 907 112
rect 991 108 995 112
rect 1079 108 1083 112
rect 1159 108 1163 112
rect 1239 108 1243 112
rect 1327 108 1331 112
rect 1415 108 1419 112
rect 1503 108 1507 112
rect 1583 108 1587 112
rect 1663 108 1667 112
rect 1743 108 1747 112
rect 1831 111 1835 115
<< m3 >>
rect 1871 3670 1875 3671
rect 1871 3665 1875 3666
rect 2151 3670 2155 3671
rect 2151 3665 2155 3666
rect 2439 3670 2443 3671
rect 2439 3665 2443 3666
rect 2727 3670 2731 3671
rect 2727 3665 2731 3666
rect 3015 3670 3019 3671
rect 3015 3665 3019 3666
rect 3591 3670 3595 3671
rect 3591 3665 3595 3666
rect 1872 3646 1874 3665
rect 2152 3649 2154 3665
rect 2440 3649 2442 3665
rect 2728 3649 2730 3665
rect 3016 3649 3018 3665
rect 2150 3648 2156 3649
rect 1870 3645 1876 3646
rect 111 3642 115 3643
rect 111 3637 115 3638
rect 143 3642 147 3643
rect 143 3637 147 3638
rect 239 3642 243 3643
rect 239 3637 243 3638
rect 367 3642 371 3643
rect 367 3637 371 3638
rect 503 3642 507 3643
rect 503 3637 507 3638
rect 639 3642 643 3643
rect 639 3637 643 3638
rect 775 3642 779 3643
rect 775 3637 779 3638
rect 911 3642 915 3643
rect 911 3637 915 3638
rect 1055 3642 1059 3643
rect 1055 3637 1059 3638
rect 1199 3642 1203 3643
rect 1199 3637 1203 3638
rect 1831 3642 1835 3643
rect 1870 3641 1871 3645
rect 1875 3641 1876 3645
rect 2150 3644 2151 3648
rect 2155 3644 2156 3648
rect 2150 3643 2156 3644
rect 2438 3648 2444 3649
rect 2438 3644 2439 3648
rect 2443 3644 2444 3648
rect 2438 3643 2444 3644
rect 2726 3648 2732 3649
rect 2726 3644 2727 3648
rect 2731 3644 2732 3648
rect 2726 3643 2732 3644
rect 3014 3648 3020 3649
rect 3014 3644 3015 3648
rect 3019 3644 3020 3648
rect 3592 3646 3594 3665
rect 3014 3643 3020 3644
rect 3590 3645 3596 3646
rect 1870 3640 1876 3641
rect 3590 3641 3591 3645
rect 3595 3641 3596 3645
rect 3590 3640 3596 3641
rect 1831 3637 1835 3638
rect 112 3609 114 3637
rect 144 3627 146 3637
rect 240 3627 242 3637
rect 368 3627 370 3637
rect 504 3627 506 3637
rect 640 3627 642 3637
rect 776 3627 778 3637
rect 912 3627 914 3637
rect 1056 3627 1058 3637
rect 1200 3627 1202 3637
rect 142 3626 148 3627
rect 142 3622 143 3626
rect 147 3622 148 3626
rect 142 3621 148 3622
rect 238 3626 244 3627
rect 238 3622 239 3626
rect 243 3622 244 3626
rect 238 3621 244 3622
rect 366 3626 372 3627
rect 366 3622 367 3626
rect 371 3622 372 3626
rect 366 3621 372 3622
rect 502 3626 508 3627
rect 502 3622 503 3626
rect 507 3622 508 3626
rect 502 3621 508 3622
rect 638 3626 644 3627
rect 638 3622 639 3626
rect 643 3622 644 3626
rect 638 3621 644 3622
rect 774 3626 780 3627
rect 774 3622 775 3626
rect 779 3622 780 3626
rect 774 3621 780 3622
rect 910 3626 916 3627
rect 910 3622 911 3626
rect 915 3622 916 3626
rect 910 3621 916 3622
rect 1054 3626 1060 3627
rect 1054 3622 1055 3626
rect 1059 3622 1060 3626
rect 1054 3621 1060 3622
rect 1198 3626 1204 3627
rect 1198 3622 1199 3626
rect 1203 3622 1204 3626
rect 1198 3621 1204 3622
rect 1832 3609 1834 3637
rect 1870 3628 1876 3629
rect 1870 3624 1871 3628
rect 1875 3624 1876 3628
rect 1870 3623 1876 3624
rect 3590 3628 3596 3629
rect 3590 3624 3591 3628
rect 3595 3624 3596 3628
rect 3590 3623 3596 3624
rect 110 3608 116 3609
rect 110 3604 111 3608
rect 115 3604 116 3608
rect 110 3603 116 3604
rect 1830 3608 1836 3609
rect 1830 3604 1831 3608
rect 1835 3604 1836 3608
rect 1830 3603 1836 3604
rect 1872 3595 1874 3623
rect 2158 3610 2164 3611
rect 2158 3606 2159 3610
rect 2163 3606 2164 3610
rect 2158 3605 2164 3606
rect 2446 3610 2452 3611
rect 2446 3606 2447 3610
rect 2451 3606 2452 3610
rect 2446 3605 2452 3606
rect 2734 3610 2740 3611
rect 2734 3606 2735 3610
rect 2739 3606 2740 3610
rect 2734 3605 2740 3606
rect 3022 3610 3028 3611
rect 3022 3606 3023 3610
rect 3027 3606 3028 3610
rect 3022 3605 3028 3606
rect 2160 3595 2162 3605
rect 2448 3595 2450 3605
rect 2736 3595 2738 3605
rect 3024 3595 3026 3605
rect 3592 3595 3594 3623
rect 1871 3594 1875 3595
rect 110 3591 116 3592
rect 110 3587 111 3591
rect 115 3587 116 3591
rect 1830 3591 1836 3592
rect 110 3586 116 3587
rect 134 3588 140 3589
rect 112 3567 114 3586
rect 134 3584 135 3588
rect 139 3584 140 3588
rect 134 3583 140 3584
rect 230 3588 236 3589
rect 230 3584 231 3588
rect 235 3584 236 3588
rect 230 3583 236 3584
rect 358 3588 364 3589
rect 358 3584 359 3588
rect 363 3584 364 3588
rect 358 3583 364 3584
rect 494 3588 500 3589
rect 494 3584 495 3588
rect 499 3584 500 3588
rect 494 3583 500 3584
rect 630 3588 636 3589
rect 630 3584 631 3588
rect 635 3584 636 3588
rect 630 3583 636 3584
rect 766 3588 772 3589
rect 766 3584 767 3588
rect 771 3584 772 3588
rect 766 3583 772 3584
rect 902 3588 908 3589
rect 902 3584 903 3588
rect 907 3584 908 3588
rect 902 3583 908 3584
rect 1046 3588 1052 3589
rect 1046 3584 1047 3588
rect 1051 3584 1052 3588
rect 1046 3583 1052 3584
rect 1190 3588 1196 3589
rect 1190 3584 1191 3588
rect 1195 3584 1196 3588
rect 1830 3587 1831 3591
rect 1835 3587 1836 3591
rect 1871 3589 1875 3590
rect 1903 3594 1907 3595
rect 1903 3589 1907 3590
rect 1983 3594 1987 3595
rect 1983 3589 1987 3590
rect 2071 3594 2075 3595
rect 2071 3589 2075 3590
rect 2159 3594 2163 3595
rect 2159 3589 2163 3590
rect 2175 3594 2179 3595
rect 2175 3589 2179 3590
rect 2295 3594 2299 3595
rect 2295 3589 2299 3590
rect 2423 3594 2427 3595
rect 2423 3589 2427 3590
rect 2447 3594 2451 3595
rect 2447 3589 2451 3590
rect 2559 3594 2563 3595
rect 2559 3589 2563 3590
rect 2695 3594 2699 3595
rect 2695 3589 2699 3590
rect 2735 3594 2739 3595
rect 2735 3589 2739 3590
rect 2831 3594 2835 3595
rect 2831 3589 2835 3590
rect 2975 3594 2979 3595
rect 2975 3589 2979 3590
rect 3023 3594 3027 3595
rect 3023 3589 3027 3590
rect 3119 3594 3123 3595
rect 3119 3589 3123 3590
rect 3263 3594 3267 3595
rect 3263 3589 3267 3590
rect 3591 3594 3595 3595
rect 3591 3589 3595 3590
rect 1830 3586 1836 3587
rect 1190 3583 1196 3584
rect 136 3567 138 3583
rect 232 3567 234 3583
rect 360 3567 362 3583
rect 496 3567 498 3583
rect 632 3567 634 3583
rect 768 3567 770 3583
rect 904 3567 906 3583
rect 1048 3567 1050 3583
rect 1192 3567 1194 3583
rect 1832 3567 1834 3586
rect 111 3566 115 3567
rect 111 3561 115 3562
rect 135 3566 139 3567
rect 135 3561 139 3562
rect 183 3566 187 3567
rect 183 3561 187 3562
rect 231 3566 235 3567
rect 231 3561 235 3562
rect 303 3566 307 3567
rect 303 3561 307 3562
rect 359 3566 363 3567
rect 359 3561 363 3562
rect 415 3566 419 3567
rect 415 3561 419 3562
rect 495 3566 499 3567
rect 495 3561 499 3562
rect 527 3566 531 3567
rect 527 3561 531 3562
rect 631 3566 635 3567
rect 631 3561 635 3562
rect 735 3566 739 3567
rect 735 3561 739 3562
rect 767 3566 771 3567
rect 767 3561 771 3562
rect 831 3566 835 3567
rect 831 3561 835 3562
rect 903 3566 907 3567
rect 903 3561 907 3562
rect 919 3566 923 3567
rect 919 3561 923 3562
rect 1007 3566 1011 3567
rect 1007 3561 1011 3562
rect 1047 3566 1051 3567
rect 1047 3561 1051 3562
rect 1095 3566 1099 3567
rect 1095 3561 1099 3562
rect 1183 3566 1187 3567
rect 1183 3561 1187 3562
rect 1191 3566 1195 3567
rect 1191 3561 1195 3562
rect 1271 3566 1275 3567
rect 1271 3561 1275 3562
rect 1359 3566 1363 3567
rect 1359 3561 1363 3562
rect 1447 3566 1451 3567
rect 1447 3561 1451 3562
rect 1831 3566 1835 3567
rect 1831 3561 1835 3562
rect 1872 3561 1874 3589
rect 1904 3579 1906 3589
rect 1984 3579 1986 3589
rect 2072 3579 2074 3589
rect 2176 3579 2178 3589
rect 2296 3579 2298 3589
rect 2424 3579 2426 3589
rect 2560 3579 2562 3589
rect 2696 3579 2698 3589
rect 2832 3579 2834 3589
rect 2976 3579 2978 3589
rect 3120 3579 3122 3589
rect 3264 3579 3266 3589
rect 1902 3578 1908 3579
rect 1902 3574 1903 3578
rect 1907 3574 1908 3578
rect 1902 3573 1908 3574
rect 1982 3578 1988 3579
rect 1982 3574 1983 3578
rect 1987 3574 1988 3578
rect 1982 3573 1988 3574
rect 2070 3578 2076 3579
rect 2070 3574 2071 3578
rect 2075 3574 2076 3578
rect 2070 3573 2076 3574
rect 2174 3578 2180 3579
rect 2174 3574 2175 3578
rect 2179 3574 2180 3578
rect 2174 3573 2180 3574
rect 2294 3578 2300 3579
rect 2294 3574 2295 3578
rect 2299 3574 2300 3578
rect 2294 3573 2300 3574
rect 2422 3578 2428 3579
rect 2422 3574 2423 3578
rect 2427 3574 2428 3578
rect 2422 3573 2428 3574
rect 2558 3578 2564 3579
rect 2558 3574 2559 3578
rect 2563 3574 2564 3578
rect 2558 3573 2564 3574
rect 2694 3578 2700 3579
rect 2694 3574 2695 3578
rect 2699 3574 2700 3578
rect 2694 3573 2700 3574
rect 2830 3578 2836 3579
rect 2830 3574 2831 3578
rect 2835 3574 2836 3578
rect 2830 3573 2836 3574
rect 2974 3578 2980 3579
rect 2974 3574 2975 3578
rect 2979 3574 2980 3578
rect 2974 3573 2980 3574
rect 3118 3578 3124 3579
rect 3118 3574 3119 3578
rect 3123 3574 3124 3578
rect 3118 3573 3124 3574
rect 3262 3578 3268 3579
rect 3262 3574 3263 3578
rect 3267 3574 3268 3578
rect 3262 3573 3268 3574
rect 3592 3561 3594 3589
rect 112 3542 114 3561
rect 184 3545 186 3561
rect 304 3545 306 3561
rect 416 3545 418 3561
rect 528 3545 530 3561
rect 632 3545 634 3561
rect 736 3545 738 3561
rect 832 3545 834 3561
rect 920 3545 922 3561
rect 1008 3545 1010 3561
rect 1096 3545 1098 3561
rect 1184 3545 1186 3561
rect 1272 3545 1274 3561
rect 1360 3545 1362 3561
rect 1448 3545 1450 3561
rect 182 3544 188 3545
rect 110 3541 116 3542
rect 110 3537 111 3541
rect 115 3537 116 3541
rect 182 3540 183 3544
rect 187 3540 188 3544
rect 182 3539 188 3540
rect 302 3544 308 3545
rect 302 3540 303 3544
rect 307 3540 308 3544
rect 302 3539 308 3540
rect 414 3544 420 3545
rect 414 3540 415 3544
rect 419 3540 420 3544
rect 414 3539 420 3540
rect 526 3544 532 3545
rect 526 3540 527 3544
rect 531 3540 532 3544
rect 526 3539 532 3540
rect 630 3544 636 3545
rect 630 3540 631 3544
rect 635 3540 636 3544
rect 630 3539 636 3540
rect 734 3544 740 3545
rect 734 3540 735 3544
rect 739 3540 740 3544
rect 734 3539 740 3540
rect 830 3544 836 3545
rect 830 3540 831 3544
rect 835 3540 836 3544
rect 830 3539 836 3540
rect 918 3544 924 3545
rect 918 3540 919 3544
rect 923 3540 924 3544
rect 918 3539 924 3540
rect 1006 3544 1012 3545
rect 1006 3540 1007 3544
rect 1011 3540 1012 3544
rect 1006 3539 1012 3540
rect 1094 3544 1100 3545
rect 1094 3540 1095 3544
rect 1099 3540 1100 3544
rect 1094 3539 1100 3540
rect 1182 3544 1188 3545
rect 1182 3540 1183 3544
rect 1187 3540 1188 3544
rect 1182 3539 1188 3540
rect 1270 3544 1276 3545
rect 1270 3540 1271 3544
rect 1275 3540 1276 3544
rect 1270 3539 1276 3540
rect 1358 3544 1364 3545
rect 1358 3540 1359 3544
rect 1363 3540 1364 3544
rect 1358 3539 1364 3540
rect 1446 3544 1452 3545
rect 1446 3540 1447 3544
rect 1451 3540 1452 3544
rect 1832 3542 1834 3561
rect 1870 3560 1876 3561
rect 1870 3556 1871 3560
rect 1875 3556 1876 3560
rect 1870 3555 1876 3556
rect 3590 3560 3596 3561
rect 3590 3556 3591 3560
rect 3595 3556 3596 3560
rect 3590 3555 3596 3556
rect 1870 3543 1876 3544
rect 1446 3539 1452 3540
rect 1830 3541 1836 3542
rect 110 3536 116 3537
rect 1830 3537 1831 3541
rect 1835 3537 1836 3541
rect 1870 3539 1871 3543
rect 1875 3539 1876 3543
rect 3590 3543 3596 3544
rect 1870 3538 1876 3539
rect 1894 3540 1900 3541
rect 1830 3536 1836 3537
rect 110 3524 116 3525
rect 110 3520 111 3524
rect 115 3520 116 3524
rect 110 3519 116 3520
rect 1830 3524 1836 3525
rect 1830 3520 1831 3524
rect 1835 3520 1836 3524
rect 1830 3519 1836 3520
rect 1872 3519 1874 3538
rect 1894 3536 1895 3540
rect 1899 3536 1900 3540
rect 1894 3535 1900 3536
rect 1974 3540 1980 3541
rect 1974 3536 1975 3540
rect 1979 3536 1980 3540
rect 1974 3535 1980 3536
rect 2062 3540 2068 3541
rect 2062 3536 2063 3540
rect 2067 3536 2068 3540
rect 2062 3535 2068 3536
rect 2166 3540 2172 3541
rect 2166 3536 2167 3540
rect 2171 3536 2172 3540
rect 2166 3535 2172 3536
rect 2286 3540 2292 3541
rect 2286 3536 2287 3540
rect 2291 3536 2292 3540
rect 2286 3535 2292 3536
rect 2414 3540 2420 3541
rect 2414 3536 2415 3540
rect 2419 3536 2420 3540
rect 2414 3535 2420 3536
rect 2550 3540 2556 3541
rect 2550 3536 2551 3540
rect 2555 3536 2556 3540
rect 2550 3535 2556 3536
rect 2686 3540 2692 3541
rect 2686 3536 2687 3540
rect 2691 3536 2692 3540
rect 2686 3535 2692 3536
rect 2822 3540 2828 3541
rect 2822 3536 2823 3540
rect 2827 3536 2828 3540
rect 2822 3535 2828 3536
rect 2966 3540 2972 3541
rect 2966 3536 2967 3540
rect 2971 3536 2972 3540
rect 2966 3535 2972 3536
rect 3110 3540 3116 3541
rect 3110 3536 3111 3540
rect 3115 3536 3116 3540
rect 3110 3535 3116 3536
rect 3254 3540 3260 3541
rect 3254 3536 3255 3540
rect 3259 3536 3260 3540
rect 3590 3539 3591 3543
rect 3595 3539 3596 3543
rect 3590 3538 3596 3539
rect 3254 3535 3260 3536
rect 1896 3519 1898 3535
rect 1976 3519 1978 3535
rect 2064 3519 2066 3535
rect 2168 3519 2170 3535
rect 2288 3519 2290 3535
rect 2416 3519 2418 3535
rect 2552 3519 2554 3535
rect 2688 3519 2690 3535
rect 2824 3519 2826 3535
rect 2968 3519 2970 3535
rect 3112 3519 3114 3535
rect 3256 3519 3258 3535
rect 3592 3519 3594 3538
rect 112 3483 114 3519
rect 190 3506 196 3507
rect 190 3502 191 3506
rect 195 3502 196 3506
rect 190 3501 196 3502
rect 310 3506 316 3507
rect 310 3502 311 3506
rect 315 3502 316 3506
rect 310 3501 316 3502
rect 422 3506 428 3507
rect 422 3502 423 3506
rect 427 3502 428 3506
rect 422 3501 428 3502
rect 534 3506 540 3507
rect 534 3502 535 3506
rect 539 3502 540 3506
rect 534 3501 540 3502
rect 638 3506 644 3507
rect 638 3502 639 3506
rect 643 3502 644 3506
rect 638 3501 644 3502
rect 742 3506 748 3507
rect 742 3502 743 3506
rect 747 3502 748 3506
rect 742 3501 748 3502
rect 838 3506 844 3507
rect 838 3502 839 3506
rect 843 3502 844 3506
rect 838 3501 844 3502
rect 926 3506 932 3507
rect 926 3502 927 3506
rect 931 3502 932 3506
rect 926 3501 932 3502
rect 1014 3506 1020 3507
rect 1014 3502 1015 3506
rect 1019 3502 1020 3506
rect 1014 3501 1020 3502
rect 1102 3506 1108 3507
rect 1102 3502 1103 3506
rect 1107 3502 1108 3506
rect 1102 3501 1108 3502
rect 1190 3506 1196 3507
rect 1190 3502 1191 3506
rect 1195 3502 1196 3506
rect 1190 3501 1196 3502
rect 1278 3506 1284 3507
rect 1278 3502 1279 3506
rect 1283 3502 1284 3506
rect 1278 3501 1284 3502
rect 1366 3506 1372 3507
rect 1366 3502 1367 3506
rect 1371 3502 1372 3506
rect 1366 3501 1372 3502
rect 1454 3506 1460 3507
rect 1454 3502 1455 3506
rect 1459 3502 1460 3506
rect 1454 3501 1460 3502
rect 192 3483 194 3501
rect 312 3483 314 3501
rect 424 3483 426 3501
rect 536 3483 538 3501
rect 640 3483 642 3501
rect 744 3483 746 3501
rect 840 3483 842 3501
rect 928 3483 930 3501
rect 1016 3483 1018 3501
rect 1104 3483 1106 3501
rect 1192 3483 1194 3501
rect 1280 3483 1282 3501
rect 1368 3483 1370 3501
rect 1456 3483 1458 3501
rect 1832 3483 1834 3519
rect 1871 3518 1875 3519
rect 1871 3513 1875 3514
rect 1895 3518 1899 3519
rect 1895 3513 1899 3514
rect 1967 3518 1971 3519
rect 1967 3513 1971 3514
rect 1975 3518 1979 3519
rect 1975 3513 1979 3514
rect 2063 3518 2067 3519
rect 2063 3513 2067 3514
rect 2151 3518 2155 3519
rect 2151 3513 2155 3514
rect 2167 3518 2171 3519
rect 2167 3513 2171 3514
rect 2287 3518 2291 3519
rect 2287 3513 2291 3514
rect 2335 3518 2339 3519
rect 2335 3513 2339 3514
rect 2415 3518 2419 3519
rect 2415 3513 2419 3514
rect 2511 3518 2515 3519
rect 2511 3513 2515 3514
rect 2551 3518 2555 3519
rect 2551 3513 2555 3514
rect 2671 3518 2675 3519
rect 2671 3513 2675 3514
rect 2687 3518 2691 3519
rect 2687 3513 2691 3514
rect 2823 3518 2827 3519
rect 2823 3513 2827 3514
rect 2959 3518 2963 3519
rect 2959 3513 2963 3514
rect 2967 3518 2971 3519
rect 2967 3513 2971 3514
rect 3079 3518 3083 3519
rect 3079 3513 3083 3514
rect 3111 3518 3115 3519
rect 3111 3513 3115 3514
rect 3191 3518 3195 3519
rect 3191 3513 3195 3514
rect 3255 3518 3259 3519
rect 3255 3513 3259 3514
rect 3303 3518 3307 3519
rect 3303 3513 3307 3514
rect 3415 3518 3419 3519
rect 3415 3513 3419 3514
rect 3503 3518 3507 3519
rect 3503 3513 3507 3514
rect 3591 3518 3595 3519
rect 3591 3513 3595 3514
rect 1872 3494 1874 3513
rect 1968 3497 1970 3513
rect 2152 3497 2154 3513
rect 2336 3497 2338 3513
rect 2512 3497 2514 3513
rect 2672 3497 2674 3513
rect 2824 3497 2826 3513
rect 2960 3497 2962 3513
rect 3080 3497 3082 3513
rect 3192 3497 3194 3513
rect 3304 3497 3306 3513
rect 3416 3497 3418 3513
rect 3504 3497 3506 3513
rect 1966 3496 1972 3497
rect 1870 3493 1876 3494
rect 1870 3489 1871 3493
rect 1875 3489 1876 3493
rect 1966 3492 1967 3496
rect 1971 3492 1972 3496
rect 1966 3491 1972 3492
rect 2150 3496 2156 3497
rect 2150 3492 2151 3496
rect 2155 3492 2156 3496
rect 2150 3491 2156 3492
rect 2334 3496 2340 3497
rect 2334 3492 2335 3496
rect 2339 3492 2340 3496
rect 2334 3491 2340 3492
rect 2510 3496 2516 3497
rect 2510 3492 2511 3496
rect 2515 3492 2516 3496
rect 2510 3491 2516 3492
rect 2670 3496 2676 3497
rect 2670 3492 2671 3496
rect 2675 3492 2676 3496
rect 2670 3491 2676 3492
rect 2822 3496 2828 3497
rect 2822 3492 2823 3496
rect 2827 3492 2828 3496
rect 2822 3491 2828 3492
rect 2958 3496 2964 3497
rect 2958 3492 2959 3496
rect 2963 3492 2964 3496
rect 2958 3491 2964 3492
rect 3078 3496 3084 3497
rect 3078 3492 3079 3496
rect 3083 3492 3084 3496
rect 3078 3491 3084 3492
rect 3190 3496 3196 3497
rect 3190 3492 3191 3496
rect 3195 3492 3196 3496
rect 3190 3491 3196 3492
rect 3302 3496 3308 3497
rect 3302 3492 3303 3496
rect 3307 3492 3308 3496
rect 3302 3491 3308 3492
rect 3414 3496 3420 3497
rect 3414 3492 3415 3496
rect 3419 3492 3420 3496
rect 3414 3491 3420 3492
rect 3502 3496 3508 3497
rect 3502 3492 3503 3496
rect 3507 3492 3508 3496
rect 3592 3494 3594 3513
rect 3502 3491 3508 3492
rect 3590 3493 3596 3494
rect 1870 3488 1876 3489
rect 3590 3489 3591 3493
rect 3595 3489 3596 3493
rect 3590 3488 3596 3489
rect 111 3482 115 3483
rect 111 3477 115 3478
rect 191 3482 195 3483
rect 191 3477 195 3478
rect 231 3482 235 3483
rect 231 3477 235 3478
rect 311 3482 315 3483
rect 311 3477 315 3478
rect 367 3482 371 3483
rect 367 3477 371 3478
rect 423 3482 427 3483
rect 423 3477 427 3478
rect 503 3482 507 3483
rect 503 3477 507 3478
rect 535 3482 539 3483
rect 535 3477 539 3478
rect 623 3482 627 3483
rect 623 3477 627 3478
rect 639 3482 643 3483
rect 639 3477 643 3478
rect 735 3482 739 3483
rect 735 3477 739 3478
rect 743 3482 747 3483
rect 743 3477 747 3478
rect 839 3482 843 3483
rect 839 3477 843 3478
rect 927 3482 931 3483
rect 927 3477 931 3478
rect 943 3482 947 3483
rect 943 3477 947 3478
rect 1015 3482 1019 3483
rect 1015 3477 1019 3478
rect 1039 3482 1043 3483
rect 1039 3477 1043 3478
rect 1103 3482 1107 3483
rect 1103 3477 1107 3478
rect 1135 3482 1139 3483
rect 1135 3477 1139 3478
rect 1191 3482 1195 3483
rect 1191 3477 1195 3478
rect 1231 3482 1235 3483
rect 1231 3477 1235 3478
rect 1279 3482 1283 3483
rect 1279 3477 1283 3478
rect 1327 3482 1331 3483
rect 1327 3477 1331 3478
rect 1367 3482 1371 3483
rect 1367 3477 1371 3478
rect 1455 3482 1459 3483
rect 1455 3477 1459 3478
rect 1831 3482 1835 3483
rect 1831 3477 1835 3478
rect 112 3449 114 3477
rect 232 3467 234 3477
rect 368 3467 370 3477
rect 504 3467 506 3477
rect 624 3467 626 3477
rect 736 3467 738 3477
rect 840 3467 842 3477
rect 944 3467 946 3477
rect 1040 3467 1042 3477
rect 1136 3467 1138 3477
rect 1232 3467 1234 3477
rect 1328 3467 1330 3477
rect 230 3466 236 3467
rect 230 3462 231 3466
rect 235 3462 236 3466
rect 230 3461 236 3462
rect 366 3466 372 3467
rect 366 3462 367 3466
rect 371 3462 372 3466
rect 366 3461 372 3462
rect 502 3466 508 3467
rect 502 3462 503 3466
rect 507 3462 508 3466
rect 502 3461 508 3462
rect 622 3466 628 3467
rect 622 3462 623 3466
rect 627 3462 628 3466
rect 622 3461 628 3462
rect 734 3466 740 3467
rect 734 3462 735 3466
rect 739 3462 740 3466
rect 734 3461 740 3462
rect 838 3466 844 3467
rect 838 3462 839 3466
rect 843 3462 844 3466
rect 838 3461 844 3462
rect 942 3466 948 3467
rect 942 3462 943 3466
rect 947 3462 948 3466
rect 942 3461 948 3462
rect 1038 3466 1044 3467
rect 1038 3462 1039 3466
rect 1043 3462 1044 3466
rect 1038 3461 1044 3462
rect 1134 3466 1140 3467
rect 1134 3462 1135 3466
rect 1139 3462 1140 3466
rect 1134 3461 1140 3462
rect 1230 3466 1236 3467
rect 1230 3462 1231 3466
rect 1235 3462 1236 3466
rect 1230 3461 1236 3462
rect 1326 3466 1332 3467
rect 1326 3462 1327 3466
rect 1331 3462 1332 3466
rect 1326 3461 1332 3462
rect 1832 3449 1834 3477
rect 1870 3476 1876 3477
rect 1870 3472 1871 3476
rect 1875 3472 1876 3476
rect 1870 3471 1876 3472
rect 3590 3476 3596 3477
rect 3590 3472 3591 3476
rect 3595 3472 3596 3476
rect 3590 3471 3596 3472
rect 110 3448 116 3449
rect 110 3444 111 3448
rect 115 3444 116 3448
rect 110 3443 116 3444
rect 1830 3448 1836 3449
rect 1830 3444 1831 3448
rect 1835 3444 1836 3448
rect 1830 3443 1836 3444
rect 1872 3443 1874 3471
rect 1974 3458 1980 3459
rect 1974 3454 1975 3458
rect 1979 3454 1980 3458
rect 1974 3453 1980 3454
rect 2158 3458 2164 3459
rect 2158 3454 2159 3458
rect 2163 3454 2164 3458
rect 2158 3453 2164 3454
rect 2342 3458 2348 3459
rect 2342 3454 2343 3458
rect 2347 3454 2348 3458
rect 2342 3453 2348 3454
rect 2518 3458 2524 3459
rect 2518 3454 2519 3458
rect 2523 3454 2524 3458
rect 2518 3453 2524 3454
rect 2678 3458 2684 3459
rect 2678 3454 2679 3458
rect 2683 3454 2684 3458
rect 2678 3453 2684 3454
rect 2830 3458 2836 3459
rect 2830 3454 2831 3458
rect 2835 3454 2836 3458
rect 2830 3453 2836 3454
rect 2966 3458 2972 3459
rect 2966 3454 2967 3458
rect 2971 3454 2972 3458
rect 2966 3453 2972 3454
rect 3086 3458 3092 3459
rect 3086 3454 3087 3458
rect 3091 3454 3092 3458
rect 3086 3453 3092 3454
rect 3198 3458 3204 3459
rect 3198 3454 3199 3458
rect 3203 3454 3204 3458
rect 3198 3453 3204 3454
rect 3310 3458 3316 3459
rect 3310 3454 3311 3458
rect 3315 3454 3316 3458
rect 3310 3453 3316 3454
rect 3422 3458 3428 3459
rect 3422 3454 3423 3458
rect 3427 3454 3428 3458
rect 3422 3453 3428 3454
rect 3510 3458 3516 3459
rect 3510 3454 3511 3458
rect 3515 3454 3516 3458
rect 3510 3453 3516 3454
rect 1976 3443 1978 3453
rect 2160 3443 2162 3453
rect 2344 3443 2346 3453
rect 2520 3443 2522 3453
rect 2680 3443 2682 3453
rect 2832 3443 2834 3453
rect 2968 3443 2970 3453
rect 3088 3443 3090 3453
rect 3200 3443 3202 3453
rect 3312 3443 3314 3453
rect 3424 3443 3426 3453
rect 3512 3443 3514 3453
rect 3592 3443 3594 3471
rect 1871 3442 1875 3443
rect 1871 3437 1875 3438
rect 1975 3442 1979 3443
rect 1975 3437 1979 3438
rect 2007 3442 2011 3443
rect 2007 3437 2011 3438
rect 2127 3442 2131 3443
rect 2127 3437 2131 3438
rect 2159 3442 2163 3443
rect 2159 3437 2163 3438
rect 2255 3442 2259 3443
rect 2255 3437 2259 3438
rect 2343 3442 2347 3443
rect 2343 3437 2347 3438
rect 2391 3442 2395 3443
rect 2391 3437 2395 3438
rect 2519 3442 2523 3443
rect 2519 3437 2523 3438
rect 2535 3442 2539 3443
rect 2535 3437 2539 3438
rect 2679 3442 2683 3443
rect 2679 3437 2683 3438
rect 2831 3442 2835 3443
rect 2831 3437 2835 3438
rect 2967 3442 2971 3443
rect 2967 3437 2971 3438
rect 2999 3442 3003 3443
rect 2999 3437 3003 3438
rect 3087 3442 3091 3443
rect 3087 3437 3091 3438
rect 3167 3442 3171 3443
rect 3167 3437 3171 3438
rect 3199 3442 3203 3443
rect 3199 3437 3203 3438
rect 3311 3442 3315 3443
rect 3311 3437 3315 3438
rect 3343 3442 3347 3443
rect 3343 3437 3347 3438
rect 3423 3442 3427 3443
rect 3423 3437 3427 3438
rect 3511 3442 3515 3443
rect 3511 3437 3515 3438
rect 3591 3442 3595 3443
rect 3591 3437 3595 3438
rect 110 3431 116 3432
rect 110 3427 111 3431
rect 115 3427 116 3431
rect 1830 3431 1836 3432
rect 110 3426 116 3427
rect 222 3428 228 3429
rect 112 3403 114 3426
rect 222 3424 223 3428
rect 227 3424 228 3428
rect 222 3423 228 3424
rect 358 3428 364 3429
rect 358 3424 359 3428
rect 363 3424 364 3428
rect 358 3423 364 3424
rect 494 3428 500 3429
rect 494 3424 495 3428
rect 499 3424 500 3428
rect 494 3423 500 3424
rect 614 3428 620 3429
rect 614 3424 615 3428
rect 619 3424 620 3428
rect 614 3423 620 3424
rect 726 3428 732 3429
rect 726 3424 727 3428
rect 731 3424 732 3428
rect 726 3423 732 3424
rect 830 3428 836 3429
rect 830 3424 831 3428
rect 835 3424 836 3428
rect 830 3423 836 3424
rect 934 3428 940 3429
rect 934 3424 935 3428
rect 939 3424 940 3428
rect 934 3423 940 3424
rect 1030 3428 1036 3429
rect 1030 3424 1031 3428
rect 1035 3424 1036 3428
rect 1030 3423 1036 3424
rect 1126 3428 1132 3429
rect 1126 3424 1127 3428
rect 1131 3424 1132 3428
rect 1126 3423 1132 3424
rect 1222 3428 1228 3429
rect 1222 3424 1223 3428
rect 1227 3424 1228 3428
rect 1222 3423 1228 3424
rect 1318 3428 1324 3429
rect 1318 3424 1319 3428
rect 1323 3424 1324 3428
rect 1830 3427 1831 3431
rect 1835 3427 1836 3431
rect 1830 3426 1836 3427
rect 1318 3423 1324 3424
rect 224 3403 226 3423
rect 360 3403 362 3423
rect 496 3403 498 3423
rect 616 3403 618 3423
rect 728 3403 730 3423
rect 832 3403 834 3423
rect 936 3403 938 3423
rect 1032 3403 1034 3423
rect 1128 3403 1130 3423
rect 1224 3403 1226 3423
rect 1320 3403 1322 3423
rect 1832 3403 1834 3426
rect 1872 3409 1874 3437
rect 2008 3427 2010 3437
rect 2128 3427 2130 3437
rect 2256 3427 2258 3437
rect 2392 3427 2394 3437
rect 2536 3427 2538 3437
rect 2680 3427 2682 3437
rect 2832 3427 2834 3437
rect 3000 3427 3002 3437
rect 3168 3427 3170 3437
rect 3344 3427 3346 3437
rect 3512 3427 3514 3437
rect 2006 3426 2012 3427
rect 2006 3422 2007 3426
rect 2011 3422 2012 3426
rect 2006 3421 2012 3422
rect 2126 3426 2132 3427
rect 2126 3422 2127 3426
rect 2131 3422 2132 3426
rect 2126 3421 2132 3422
rect 2254 3426 2260 3427
rect 2254 3422 2255 3426
rect 2259 3422 2260 3426
rect 2254 3421 2260 3422
rect 2390 3426 2396 3427
rect 2390 3422 2391 3426
rect 2395 3422 2396 3426
rect 2390 3421 2396 3422
rect 2534 3426 2540 3427
rect 2534 3422 2535 3426
rect 2539 3422 2540 3426
rect 2534 3421 2540 3422
rect 2678 3426 2684 3427
rect 2678 3422 2679 3426
rect 2683 3422 2684 3426
rect 2678 3421 2684 3422
rect 2830 3426 2836 3427
rect 2830 3422 2831 3426
rect 2835 3422 2836 3426
rect 2830 3421 2836 3422
rect 2998 3426 3004 3427
rect 2998 3422 2999 3426
rect 3003 3422 3004 3426
rect 2998 3421 3004 3422
rect 3166 3426 3172 3427
rect 3166 3422 3167 3426
rect 3171 3422 3172 3426
rect 3166 3421 3172 3422
rect 3342 3426 3348 3427
rect 3342 3422 3343 3426
rect 3347 3422 3348 3426
rect 3342 3421 3348 3422
rect 3510 3426 3516 3427
rect 3510 3422 3511 3426
rect 3515 3422 3516 3426
rect 3510 3421 3516 3422
rect 3592 3409 3594 3437
rect 1870 3408 1876 3409
rect 1870 3404 1871 3408
rect 1875 3404 1876 3408
rect 1870 3403 1876 3404
rect 3590 3408 3596 3409
rect 3590 3404 3591 3408
rect 3595 3404 3596 3408
rect 3590 3403 3596 3404
rect 111 3402 115 3403
rect 111 3397 115 3398
rect 215 3402 219 3403
rect 215 3397 219 3398
rect 223 3402 227 3403
rect 223 3397 227 3398
rect 359 3402 363 3403
rect 359 3397 363 3398
rect 367 3402 371 3403
rect 367 3397 371 3398
rect 495 3402 499 3403
rect 495 3397 499 3398
rect 511 3402 515 3403
rect 511 3397 515 3398
rect 615 3402 619 3403
rect 615 3397 619 3398
rect 647 3402 651 3403
rect 647 3397 651 3398
rect 727 3402 731 3403
rect 727 3397 731 3398
rect 775 3402 779 3403
rect 775 3397 779 3398
rect 831 3402 835 3403
rect 831 3397 835 3398
rect 895 3402 899 3403
rect 895 3397 899 3398
rect 935 3402 939 3403
rect 935 3397 939 3398
rect 1015 3402 1019 3403
rect 1015 3397 1019 3398
rect 1031 3402 1035 3403
rect 1031 3397 1035 3398
rect 1127 3402 1131 3403
rect 1127 3397 1131 3398
rect 1223 3402 1227 3403
rect 1223 3397 1227 3398
rect 1239 3402 1243 3403
rect 1239 3397 1243 3398
rect 1319 3402 1323 3403
rect 1319 3397 1323 3398
rect 1351 3402 1355 3403
rect 1351 3397 1355 3398
rect 1831 3402 1835 3403
rect 1831 3397 1835 3398
rect 112 3378 114 3397
rect 216 3381 218 3397
rect 368 3381 370 3397
rect 512 3381 514 3397
rect 648 3381 650 3397
rect 776 3381 778 3397
rect 896 3381 898 3397
rect 1016 3381 1018 3397
rect 1128 3381 1130 3397
rect 1240 3381 1242 3397
rect 1352 3381 1354 3397
rect 214 3380 220 3381
rect 110 3377 116 3378
rect 110 3373 111 3377
rect 115 3373 116 3377
rect 214 3376 215 3380
rect 219 3376 220 3380
rect 214 3375 220 3376
rect 366 3380 372 3381
rect 366 3376 367 3380
rect 371 3376 372 3380
rect 366 3375 372 3376
rect 510 3380 516 3381
rect 510 3376 511 3380
rect 515 3376 516 3380
rect 510 3375 516 3376
rect 646 3380 652 3381
rect 646 3376 647 3380
rect 651 3376 652 3380
rect 646 3375 652 3376
rect 774 3380 780 3381
rect 774 3376 775 3380
rect 779 3376 780 3380
rect 774 3375 780 3376
rect 894 3380 900 3381
rect 894 3376 895 3380
rect 899 3376 900 3380
rect 894 3375 900 3376
rect 1014 3380 1020 3381
rect 1014 3376 1015 3380
rect 1019 3376 1020 3380
rect 1014 3375 1020 3376
rect 1126 3380 1132 3381
rect 1126 3376 1127 3380
rect 1131 3376 1132 3380
rect 1126 3375 1132 3376
rect 1238 3380 1244 3381
rect 1238 3376 1239 3380
rect 1243 3376 1244 3380
rect 1238 3375 1244 3376
rect 1350 3380 1356 3381
rect 1350 3376 1351 3380
rect 1355 3376 1356 3380
rect 1832 3378 1834 3397
rect 1870 3391 1876 3392
rect 1870 3387 1871 3391
rect 1875 3387 1876 3391
rect 3590 3391 3596 3392
rect 1870 3386 1876 3387
rect 1998 3388 2004 3389
rect 1350 3375 1356 3376
rect 1830 3377 1836 3378
rect 110 3372 116 3373
rect 1830 3373 1831 3377
rect 1835 3373 1836 3377
rect 1830 3372 1836 3373
rect 1872 3367 1874 3386
rect 1998 3384 1999 3388
rect 2003 3384 2004 3388
rect 1998 3383 2004 3384
rect 2118 3388 2124 3389
rect 2118 3384 2119 3388
rect 2123 3384 2124 3388
rect 2118 3383 2124 3384
rect 2246 3388 2252 3389
rect 2246 3384 2247 3388
rect 2251 3384 2252 3388
rect 2246 3383 2252 3384
rect 2382 3388 2388 3389
rect 2382 3384 2383 3388
rect 2387 3384 2388 3388
rect 2382 3383 2388 3384
rect 2526 3388 2532 3389
rect 2526 3384 2527 3388
rect 2531 3384 2532 3388
rect 2526 3383 2532 3384
rect 2670 3388 2676 3389
rect 2670 3384 2671 3388
rect 2675 3384 2676 3388
rect 2670 3383 2676 3384
rect 2822 3388 2828 3389
rect 2822 3384 2823 3388
rect 2827 3384 2828 3388
rect 2822 3383 2828 3384
rect 2990 3388 2996 3389
rect 2990 3384 2991 3388
rect 2995 3384 2996 3388
rect 2990 3383 2996 3384
rect 3158 3388 3164 3389
rect 3158 3384 3159 3388
rect 3163 3384 3164 3388
rect 3158 3383 3164 3384
rect 3334 3388 3340 3389
rect 3334 3384 3335 3388
rect 3339 3384 3340 3388
rect 3334 3383 3340 3384
rect 3502 3388 3508 3389
rect 3502 3384 3503 3388
rect 3507 3384 3508 3388
rect 3590 3387 3591 3391
rect 3595 3387 3596 3391
rect 3590 3386 3596 3387
rect 3502 3383 3508 3384
rect 2000 3367 2002 3383
rect 2120 3367 2122 3383
rect 2248 3367 2250 3383
rect 2384 3367 2386 3383
rect 2528 3367 2530 3383
rect 2672 3367 2674 3383
rect 2824 3367 2826 3383
rect 2992 3367 2994 3383
rect 3160 3367 3162 3383
rect 3336 3367 3338 3383
rect 3504 3367 3506 3383
rect 3592 3367 3594 3386
rect 1871 3366 1875 3367
rect 1871 3361 1875 3362
rect 1999 3366 2003 3367
rect 1999 3361 2003 3362
rect 2015 3366 2019 3367
rect 2015 3361 2019 3362
rect 2119 3366 2123 3367
rect 2119 3361 2123 3362
rect 2151 3366 2155 3367
rect 2151 3361 2155 3362
rect 2247 3366 2251 3367
rect 2247 3361 2251 3362
rect 2295 3366 2299 3367
rect 2295 3361 2299 3362
rect 2383 3366 2387 3367
rect 2383 3361 2387 3362
rect 2439 3366 2443 3367
rect 2439 3361 2443 3362
rect 2527 3366 2531 3367
rect 2527 3361 2531 3362
rect 2583 3366 2587 3367
rect 2583 3361 2587 3362
rect 2671 3366 2675 3367
rect 2671 3361 2675 3362
rect 2727 3366 2731 3367
rect 2727 3361 2731 3362
rect 2823 3366 2827 3367
rect 2823 3361 2827 3362
rect 2871 3366 2875 3367
rect 2871 3361 2875 3362
rect 2991 3366 2995 3367
rect 2991 3361 2995 3362
rect 3023 3366 3027 3367
rect 3023 3361 3027 3362
rect 3159 3366 3163 3367
rect 3159 3361 3163 3362
rect 3183 3366 3187 3367
rect 3183 3361 3187 3362
rect 3335 3366 3339 3367
rect 3335 3361 3339 3362
rect 3351 3366 3355 3367
rect 3351 3361 3355 3362
rect 3503 3366 3507 3367
rect 3503 3361 3507 3362
rect 3591 3366 3595 3367
rect 3591 3361 3595 3362
rect 110 3360 116 3361
rect 110 3356 111 3360
rect 115 3356 116 3360
rect 110 3355 116 3356
rect 1830 3360 1836 3361
rect 1830 3356 1831 3360
rect 1835 3356 1836 3360
rect 1830 3355 1836 3356
rect 112 3323 114 3355
rect 222 3342 228 3343
rect 222 3338 223 3342
rect 227 3338 228 3342
rect 222 3337 228 3338
rect 374 3342 380 3343
rect 374 3338 375 3342
rect 379 3338 380 3342
rect 374 3337 380 3338
rect 518 3342 524 3343
rect 518 3338 519 3342
rect 523 3338 524 3342
rect 518 3337 524 3338
rect 654 3342 660 3343
rect 654 3338 655 3342
rect 659 3338 660 3342
rect 654 3337 660 3338
rect 782 3342 788 3343
rect 782 3338 783 3342
rect 787 3338 788 3342
rect 782 3337 788 3338
rect 902 3342 908 3343
rect 902 3338 903 3342
rect 907 3338 908 3342
rect 902 3337 908 3338
rect 1022 3342 1028 3343
rect 1022 3338 1023 3342
rect 1027 3338 1028 3342
rect 1022 3337 1028 3338
rect 1134 3342 1140 3343
rect 1134 3338 1135 3342
rect 1139 3338 1140 3342
rect 1134 3337 1140 3338
rect 1246 3342 1252 3343
rect 1246 3338 1247 3342
rect 1251 3338 1252 3342
rect 1246 3337 1252 3338
rect 1358 3342 1364 3343
rect 1358 3338 1359 3342
rect 1363 3338 1364 3342
rect 1358 3337 1364 3338
rect 224 3323 226 3337
rect 376 3323 378 3337
rect 520 3323 522 3337
rect 656 3323 658 3337
rect 784 3323 786 3337
rect 904 3323 906 3337
rect 1024 3323 1026 3337
rect 1136 3323 1138 3337
rect 1248 3323 1250 3337
rect 1360 3323 1362 3337
rect 1832 3323 1834 3355
rect 1872 3342 1874 3361
rect 2016 3345 2018 3361
rect 2152 3345 2154 3361
rect 2296 3345 2298 3361
rect 2440 3345 2442 3361
rect 2584 3345 2586 3361
rect 2728 3345 2730 3361
rect 2872 3345 2874 3361
rect 3024 3345 3026 3361
rect 3184 3345 3186 3361
rect 3352 3345 3354 3361
rect 3504 3345 3506 3361
rect 2014 3344 2020 3345
rect 1870 3341 1876 3342
rect 1870 3337 1871 3341
rect 1875 3337 1876 3341
rect 2014 3340 2015 3344
rect 2019 3340 2020 3344
rect 2014 3339 2020 3340
rect 2150 3344 2156 3345
rect 2150 3340 2151 3344
rect 2155 3340 2156 3344
rect 2150 3339 2156 3340
rect 2294 3344 2300 3345
rect 2294 3340 2295 3344
rect 2299 3340 2300 3344
rect 2294 3339 2300 3340
rect 2438 3344 2444 3345
rect 2438 3340 2439 3344
rect 2443 3340 2444 3344
rect 2438 3339 2444 3340
rect 2582 3344 2588 3345
rect 2582 3340 2583 3344
rect 2587 3340 2588 3344
rect 2582 3339 2588 3340
rect 2726 3344 2732 3345
rect 2726 3340 2727 3344
rect 2731 3340 2732 3344
rect 2726 3339 2732 3340
rect 2870 3344 2876 3345
rect 2870 3340 2871 3344
rect 2875 3340 2876 3344
rect 2870 3339 2876 3340
rect 3022 3344 3028 3345
rect 3022 3340 3023 3344
rect 3027 3340 3028 3344
rect 3022 3339 3028 3340
rect 3182 3344 3188 3345
rect 3182 3340 3183 3344
rect 3187 3340 3188 3344
rect 3182 3339 3188 3340
rect 3350 3344 3356 3345
rect 3350 3340 3351 3344
rect 3355 3340 3356 3344
rect 3350 3339 3356 3340
rect 3502 3344 3508 3345
rect 3502 3340 3503 3344
rect 3507 3340 3508 3344
rect 3592 3342 3594 3361
rect 3502 3339 3508 3340
rect 3590 3341 3596 3342
rect 1870 3336 1876 3337
rect 3590 3337 3591 3341
rect 3595 3337 3596 3341
rect 3590 3336 3596 3337
rect 1870 3324 1876 3325
rect 111 3322 115 3323
rect 111 3317 115 3318
rect 207 3322 211 3323
rect 207 3317 211 3318
rect 223 3322 227 3323
rect 223 3317 227 3318
rect 367 3322 371 3323
rect 367 3317 371 3318
rect 375 3322 379 3323
rect 375 3317 379 3318
rect 519 3322 523 3323
rect 519 3317 523 3318
rect 655 3322 659 3323
rect 655 3317 659 3318
rect 671 3322 675 3323
rect 671 3317 675 3318
rect 783 3322 787 3323
rect 783 3317 787 3318
rect 815 3322 819 3323
rect 815 3317 819 3318
rect 903 3322 907 3323
rect 903 3317 907 3318
rect 951 3322 955 3323
rect 951 3317 955 3318
rect 1023 3322 1027 3323
rect 1023 3317 1027 3318
rect 1087 3322 1091 3323
rect 1087 3317 1091 3318
rect 1135 3322 1139 3323
rect 1135 3317 1139 3318
rect 1215 3322 1219 3323
rect 1215 3317 1219 3318
rect 1247 3322 1251 3323
rect 1247 3317 1251 3318
rect 1343 3322 1347 3323
rect 1343 3317 1347 3318
rect 1359 3322 1363 3323
rect 1359 3317 1363 3318
rect 1471 3322 1475 3323
rect 1471 3317 1475 3318
rect 1831 3322 1835 3323
rect 1870 3320 1871 3324
rect 1875 3320 1876 3324
rect 1870 3319 1876 3320
rect 3590 3324 3596 3325
rect 3590 3320 3591 3324
rect 3595 3320 3596 3324
rect 3590 3319 3596 3320
rect 1831 3317 1835 3318
rect 112 3289 114 3317
rect 208 3307 210 3317
rect 368 3307 370 3317
rect 520 3307 522 3317
rect 672 3307 674 3317
rect 816 3307 818 3317
rect 952 3307 954 3317
rect 1088 3307 1090 3317
rect 1216 3307 1218 3317
rect 1344 3307 1346 3317
rect 1472 3307 1474 3317
rect 206 3306 212 3307
rect 206 3302 207 3306
rect 211 3302 212 3306
rect 206 3301 212 3302
rect 366 3306 372 3307
rect 366 3302 367 3306
rect 371 3302 372 3306
rect 366 3301 372 3302
rect 518 3306 524 3307
rect 518 3302 519 3306
rect 523 3302 524 3306
rect 518 3301 524 3302
rect 670 3306 676 3307
rect 670 3302 671 3306
rect 675 3302 676 3306
rect 670 3301 676 3302
rect 814 3306 820 3307
rect 814 3302 815 3306
rect 819 3302 820 3306
rect 814 3301 820 3302
rect 950 3306 956 3307
rect 950 3302 951 3306
rect 955 3302 956 3306
rect 950 3301 956 3302
rect 1086 3306 1092 3307
rect 1086 3302 1087 3306
rect 1091 3302 1092 3306
rect 1086 3301 1092 3302
rect 1214 3306 1220 3307
rect 1214 3302 1215 3306
rect 1219 3302 1220 3306
rect 1214 3301 1220 3302
rect 1342 3306 1348 3307
rect 1342 3302 1343 3306
rect 1347 3302 1348 3306
rect 1342 3301 1348 3302
rect 1470 3306 1476 3307
rect 1470 3302 1471 3306
rect 1475 3302 1476 3306
rect 1470 3301 1476 3302
rect 1832 3289 1834 3317
rect 1872 3291 1874 3319
rect 2022 3306 2028 3307
rect 2022 3302 2023 3306
rect 2027 3302 2028 3306
rect 2022 3301 2028 3302
rect 2158 3306 2164 3307
rect 2158 3302 2159 3306
rect 2163 3302 2164 3306
rect 2158 3301 2164 3302
rect 2302 3306 2308 3307
rect 2302 3302 2303 3306
rect 2307 3302 2308 3306
rect 2302 3301 2308 3302
rect 2446 3306 2452 3307
rect 2446 3302 2447 3306
rect 2451 3302 2452 3306
rect 2446 3301 2452 3302
rect 2590 3306 2596 3307
rect 2590 3302 2591 3306
rect 2595 3302 2596 3306
rect 2590 3301 2596 3302
rect 2734 3306 2740 3307
rect 2734 3302 2735 3306
rect 2739 3302 2740 3306
rect 2734 3301 2740 3302
rect 2878 3306 2884 3307
rect 2878 3302 2879 3306
rect 2883 3302 2884 3306
rect 2878 3301 2884 3302
rect 3030 3306 3036 3307
rect 3030 3302 3031 3306
rect 3035 3302 3036 3306
rect 3030 3301 3036 3302
rect 3190 3306 3196 3307
rect 3190 3302 3191 3306
rect 3195 3302 3196 3306
rect 3190 3301 3196 3302
rect 3358 3306 3364 3307
rect 3358 3302 3359 3306
rect 3363 3302 3364 3306
rect 3358 3301 3364 3302
rect 3510 3306 3516 3307
rect 3510 3302 3511 3306
rect 3515 3302 3516 3306
rect 3510 3301 3516 3302
rect 2024 3291 2026 3301
rect 2160 3291 2162 3301
rect 2304 3291 2306 3301
rect 2448 3291 2450 3301
rect 2592 3291 2594 3301
rect 2736 3291 2738 3301
rect 2880 3291 2882 3301
rect 3032 3291 3034 3301
rect 3192 3291 3194 3301
rect 3360 3291 3362 3301
rect 3512 3291 3514 3301
rect 3592 3291 3594 3319
rect 1871 3290 1875 3291
rect 110 3288 116 3289
rect 110 3284 111 3288
rect 115 3284 116 3288
rect 110 3283 116 3284
rect 1830 3288 1836 3289
rect 1830 3284 1831 3288
rect 1835 3284 1836 3288
rect 1871 3285 1875 3286
rect 1927 3290 1931 3291
rect 1927 3285 1931 3286
rect 2023 3290 2027 3291
rect 2023 3285 2027 3286
rect 2063 3290 2067 3291
rect 2063 3285 2067 3286
rect 2159 3290 2163 3291
rect 2159 3285 2163 3286
rect 2191 3290 2195 3291
rect 2191 3285 2195 3286
rect 2303 3290 2307 3291
rect 2303 3285 2307 3286
rect 2319 3290 2323 3291
rect 2319 3285 2323 3286
rect 2447 3290 2451 3291
rect 2447 3285 2451 3286
rect 2591 3290 2595 3291
rect 2591 3285 2595 3286
rect 2735 3290 2739 3291
rect 2735 3285 2739 3286
rect 2743 3290 2747 3291
rect 2743 3285 2747 3286
rect 2879 3290 2883 3291
rect 2879 3285 2883 3286
rect 2919 3290 2923 3291
rect 2919 3285 2923 3286
rect 3031 3290 3035 3291
rect 3031 3285 3035 3286
rect 3111 3290 3115 3291
rect 3111 3285 3115 3286
rect 3191 3290 3195 3291
rect 3191 3285 3195 3286
rect 3311 3290 3315 3291
rect 3311 3285 3315 3286
rect 3359 3290 3363 3291
rect 3359 3285 3363 3286
rect 3511 3290 3515 3291
rect 3511 3285 3515 3286
rect 3591 3290 3595 3291
rect 3591 3285 3595 3286
rect 1830 3283 1836 3284
rect 110 3271 116 3272
rect 110 3267 111 3271
rect 115 3267 116 3271
rect 1830 3271 1836 3272
rect 110 3266 116 3267
rect 198 3268 204 3269
rect 112 3247 114 3266
rect 198 3264 199 3268
rect 203 3264 204 3268
rect 198 3263 204 3264
rect 358 3268 364 3269
rect 358 3264 359 3268
rect 363 3264 364 3268
rect 358 3263 364 3264
rect 510 3268 516 3269
rect 510 3264 511 3268
rect 515 3264 516 3268
rect 510 3263 516 3264
rect 662 3268 668 3269
rect 662 3264 663 3268
rect 667 3264 668 3268
rect 662 3263 668 3264
rect 806 3268 812 3269
rect 806 3264 807 3268
rect 811 3264 812 3268
rect 806 3263 812 3264
rect 942 3268 948 3269
rect 942 3264 943 3268
rect 947 3264 948 3268
rect 942 3263 948 3264
rect 1078 3268 1084 3269
rect 1078 3264 1079 3268
rect 1083 3264 1084 3268
rect 1078 3263 1084 3264
rect 1206 3268 1212 3269
rect 1206 3264 1207 3268
rect 1211 3264 1212 3268
rect 1206 3263 1212 3264
rect 1334 3268 1340 3269
rect 1334 3264 1335 3268
rect 1339 3264 1340 3268
rect 1334 3263 1340 3264
rect 1462 3268 1468 3269
rect 1462 3264 1463 3268
rect 1467 3264 1468 3268
rect 1830 3267 1831 3271
rect 1835 3267 1836 3271
rect 1830 3266 1836 3267
rect 1462 3263 1468 3264
rect 200 3247 202 3263
rect 360 3247 362 3263
rect 512 3247 514 3263
rect 664 3247 666 3263
rect 808 3247 810 3263
rect 944 3247 946 3263
rect 1080 3247 1082 3263
rect 1208 3247 1210 3263
rect 1336 3247 1338 3263
rect 1464 3247 1466 3263
rect 1832 3247 1834 3266
rect 1872 3257 1874 3285
rect 1928 3275 1930 3285
rect 2064 3275 2066 3285
rect 2192 3275 2194 3285
rect 2320 3275 2322 3285
rect 2448 3275 2450 3285
rect 2592 3275 2594 3285
rect 2744 3275 2746 3285
rect 2920 3275 2922 3285
rect 3112 3275 3114 3285
rect 3312 3275 3314 3285
rect 3512 3275 3514 3285
rect 1926 3274 1932 3275
rect 1926 3270 1927 3274
rect 1931 3270 1932 3274
rect 1926 3269 1932 3270
rect 2062 3274 2068 3275
rect 2062 3270 2063 3274
rect 2067 3270 2068 3274
rect 2062 3269 2068 3270
rect 2190 3274 2196 3275
rect 2190 3270 2191 3274
rect 2195 3270 2196 3274
rect 2190 3269 2196 3270
rect 2318 3274 2324 3275
rect 2318 3270 2319 3274
rect 2323 3270 2324 3274
rect 2318 3269 2324 3270
rect 2446 3274 2452 3275
rect 2446 3270 2447 3274
rect 2451 3270 2452 3274
rect 2446 3269 2452 3270
rect 2590 3274 2596 3275
rect 2590 3270 2591 3274
rect 2595 3270 2596 3274
rect 2590 3269 2596 3270
rect 2742 3274 2748 3275
rect 2742 3270 2743 3274
rect 2747 3270 2748 3274
rect 2742 3269 2748 3270
rect 2918 3274 2924 3275
rect 2918 3270 2919 3274
rect 2923 3270 2924 3274
rect 2918 3269 2924 3270
rect 3110 3274 3116 3275
rect 3110 3270 3111 3274
rect 3115 3270 3116 3274
rect 3110 3269 3116 3270
rect 3310 3274 3316 3275
rect 3310 3270 3311 3274
rect 3315 3270 3316 3274
rect 3310 3269 3316 3270
rect 3510 3274 3516 3275
rect 3510 3270 3511 3274
rect 3515 3270 3516 3274
rect 3510 3269 3516 3270
rect 3592 3257 3594 3285
rect 1870 3256 1876 3257
rect 1870 3252 1871 3256
rect 1875 3252 1876 3256
rect 1870 3251 1876 3252
rect 3590 3256 3596 3257
rect 3590 3252 3591 3256
rect 3595 3252 3596 3256
rect 3590 3251 3596 3252
rect 111 3246 115 3247
rect 111 3241 115 3242
rect 135 3246 139 3247
rect 135 3241 139 3242
rect 199 3246 203 3247
rect 199 3241 203 3242
rect 271 3246 275 3247
rect 271 3241 275 3242
rect 359 3246 363 3247
rect 359 3241 363 3242
rect 415 3246 419 3247
rect 415 3241 419 3242
rect 511 3246 515 3247
rect 511 3241 515 3242
rect 575 3246 579 3247
rect 575 3241 579 3242
rect 663 3246 667 3247
rect 663 3241 667 3242
rect 735 3246 739 3247
rect 735 3241 739 3242
rect 807 3246 811 3247
rect 807 3241 811 3242
rect 895 3246 899 3247
rect 895 3241 899 3242
rect 943 3246 947 3247
rect 943 3241 947 3242
rect 1047 3246 1051 3247
rect 1047 3241 1051 3242
rect 1079 3246 1083 3247
rect 1079 3241 1083 3242
rect 1191 3246 1195 3247
rect 1191 3241 1195 3242
rect 1207 3246 1211 3247
rect 1207 3241 1211 3242
rect 1327 3246 1331 3247
rect 1327 3241 1331 3242
rect 1335 3246 1339 3247
rect 1335 3241 1339 3242
rect 1463 3246 1467 3247
rect 1463 3241 1467 3242
rect 1607 3246 1611 3247
rect 1607 3241 1611 3242
rect 1831 3246 1835 3247
rect 1831 3241 1835 3242
rect 112 3222 114 3241
rect 136 3225 138 3241
rect 272 3225 274 3241
rect 416 3225 418 3241
rect 576 3225 578 3241
rect 736 3225 738 3241
rect 896 3225 898 3241
rect 1048 3225 1050 3241
rect 1192 3225 1194 3241
rect 1328 3225 1330 3241
rect 1464 3225 1466 3241
rect 1608 3225 1610 3241
rect 134 3224 140 3225
rect 110 3221 116 3222
rect 110 3217 111 3221
rect 115 3217 116 3221
rect 134 3220 135 3224
rect 139 3220 140 3224
rect 134 3219 140 3220
rect 270 3224 276 3225
rect 270 3220 271 3224
rect 275 3220 276 3224
rect 270 3219 276 3220
rect 414 3224 420 3225
rect 414 3220 415 3224
rect 419 3220 420 3224
rect 414 3219 420 3220
rect 574 3224 580 3225
rect 574 3220 575 3224
rect 579 3220 580 3224
rect 574 3219 580 3220
rect 734 3224 740 3225
rect 734 3220 735 3224
rect 739 3220 740 3224
rect 734 3219 740 3220
rect 894 3224 900 3225
rect 894 3220 895 3224
rect 899 3220 900 3224
rect 894 3219 900 3220
rect 1046 3224 1052 3225
rect 1046 3220 1047 3224
rect 1051 3220 1052 3224
rect 1046 3219 1052 3220
rect 1190 3224 1196 3225
rect 1190 3220 1191 3224
rect 1195 3220 1196 3224
rect 1190 3219 1196 3220
rect 1326 3224 1332 3225
rect 1326 3220 1327 3224
rect 1331 3220 1332 3224
rect 1326 3219 1332 3220
rect 1462 3224 1468 3225
rect 1462 3220 1463 3224
rect 1467 3220 1468 3224
rect 1462 3219 1468 3220
rect 1606 3224 1612 3225
rect 1606 3220 1607 3224
rect 1611 3220 1612 3224
rect 1832 3222 1834 3241
rect 1870 3239 1876 3240
rect 1870 3235 1871 3239
rect 1875 3235 1876 3239
rect 3590 3239 3596 3240
rect 1870 3234 1876 3235
rect 1918 3236 1924 3237
rect 1606 3219 1612 3220
rect 1830 3221 1836 3222
rect 110 3216 116 3217
rect 1830 3217 1831 3221
rect 1835 3217 1836 3221
rect 1830 3216 1836 3217
rect 1872 3215 1874 3234
rect 1918 3232 1919 3236
rect 1923 3232 1924 3236
rect 1918 3231 1924 3232
rect 2054 3236 2060 3237
rect 2054 3232 2055 3236
rect 2059 3232 2060 3236
rect 2054 3231 2060 3232
rect 2182 3236 2188 3237
rect 2182 3232 2183 3236
rect 2187 3232 2188 3236
rect 2182 3231 2188 3232
rect 2310 3236 2316 3237
rect 2310 3232 2311 3236
rect 2315 3232 2316 3236
rect 2310 3231 2316 3232
rect 2438 3236 2444 3237
rect 2438 3232 2439 3236
rect 2443 3232 2444 3236
rect 2438 3231 2444 3232
rect 2582 3236 2588 3237
rect 2582 3232 2583 3236
rect 2587 3232 2588 3236
rect 2582 3231 2588 3232
rect 2734 3236 2740 3237
rect 2734 3232 2735 3236
rect 2739 3232 2740 3236
rect 2734 3231 2740 3232
rect 2910 3236 2916 3237
rect 2910 3232 2911 3236
rect 2915 3232 2916 3236
rect 2910 3231 2916 3232
rect 3102 3236 3108 3237
rect 3102 3232 3103 3236
rect 3107 3232 3108 3236
rect 3102 3231 3108 3232
rect 3302 3236 3308 3237
rect 3302 3232 3303 3236
rect 3307 3232 3308 3236
rect 3302 3231 3308 3232
rect 3502 3236 3508 3237
rect 3502 3232 3503 3236
rect 3507 3232 3508 3236
rect 3590 3235 3591 3239
rect 3595 3235 3596 3239
rect 3590 3234 3596 3235
rect 3502 3231 3508 3232
rect 1920 3215 1922 3231
rect 2056 3215 2058 3231
rect 2184 3215 2186 3231
rect 2312 3215 2314 3231
rect 2440 3215 2442 3231
rect 2584 3215 2586 3231
rect 2736 3215 2738 3231
rect 2912 3215 2914 3231
rect 3104 3215 3106 3231
rect 3304 3215 3306 3231
rect 3504 3215 3506 3231
rect 3592 3215 3594 3234
rect 1871 3214 1875 3215
rect 1871 3209 1875 3210
rect 1895 3214 1899 3215
rect 1895 3209 1899 3210
rect 1919 3214 1923 3215
rect 1919 3209 1923 3210
rect 2007 3214 2011 3215
rect 2007 3209 2011 3210
rect 2055 3214 2059 3215
rect 2055 3209 2059 3210
rect 2143 3214 2147 3215
rect 2143 3209 2147 3210
rect 2183 3214 2187 3215
rect 2183 3209 2187 3210
rect 2295 3214 2299 3215
rect 2295 3209 2299 3210
rect 2311 3214 2315 3215
rect 2311 3209 2315 3210
rect 2439 3214 2443 3215
rect 2439 3209 2443 3210
rect 2455 3214 2459 3215
rect 2455 3209 2459 3210
rect 2583 3214 2587 3215
rect 2583 3209 2587 3210
rect 2623 3214 2627 3215
rect 2623 3209 2627 3210
rect 2735 3214 2739 3215
rect 2735 3209 2739 3210
rect 2799 3214 2803 3215
rect 2799 3209 2803 3210
rect 2911 3214 2915 3215
rect 2911 3209 2915 3210
rect 2975 3214 2979 3215
rect 2975 3209 2979 3210
rect 3103 3214 3107 3215
rect 3103 3209 3107 3210
rect 3151 3214 3155 3215
rect 3151 3209 3155 3210
rect 3303 3214 3307 3215
rect 3303 3209 3307 3210
rect 3327 3214 3331 3215
rect 3327 3209 3331 3210
rect 3503 3214 3507 3215
rect 3503 3209 3507 3210
rect 3591 3214 3595 3215
rect 3591 3209 3595 3210
rect 110 3204 116 3205
rect 110 3200 111 3204
rect 115 3200 116 3204
rect 110 3199 116 3200
rect 1830 3204 1836 3205
rect 1830 3200 1831 3204
rect 1835 3200 1836 3204
rect 1830 3199 1836 3200
rect 112 3163 114 3199
rect 142 3186 148 3187
rect 142 3182 143 3186
rect 147 3182 148 3186
rect 142 3181 148 3182
rect 278 3186 284 3187
rect 278 3182 279 3186
rect 283 3182 284 3186
rect 278 3181 284 3182
rect 422 3186 428 3187
rect 422 3182 423 3186
rect 427 3182 428 3186
rect 422 3181 428 3182
rect 582 3186 588 3187
rect 582 3182 583 3186
rect 587 3182 588 3186
rect 582 3181 588 3182
rect 742 3186 748 3187
rect 742 3182 743 3186
rect 747 3182 748 3186
rect 742 3181 748 3182
rect 902 3186 908 3187
rect 902 3182 903 3186
rect 907 3182 908 3186
rect 902 3181 908 3182
rect 1054 3186 1060 3187
rect 1054 3182 1055 3186
rect 1059 3182 1060 3186
rect 1054 3181 1060 3182
rect 1198 3186 1204 3187
rect 1198 3182 1199 3186
rect 1203 3182 1204 3186
rect 1198 3181 1204 3182
rect 1334 3186 1340 3187
rect 1334 3182 1335 3186
rect 1339 3182 1340 3186
rect 1334 3181 1340 3182
rect 1470 3186 1476 3187
rect 1470 3182 1471 3186
rect 1475 3182 1476 3186
rect 1470 3181 1476 3182
rect 1614 3186 1620 3187
rect 1614 3182 1615 3186
rect 1619 3182 1620 3186
rect 1614 3181 1620 3182
rect 144 3163 146 3181
rect 280 3163 282 3181
rect 424 3163 426 3181
rect 584 3163 586 3181
rect 744 3163 746 3181
rect 904 3163 906 3181
rect 1056 3163 1058 3181
rect 1200 3163 1202 3181
rect 1336 3163 1338 3181
rect 1472 3163 1474 3181
rect 1616 3163 1618 3181
rect 1832 3163 1834 3199
rect 1872 3190 1874 3209
rect 1896 3193 1898 3209
rect 2008 3193 2010 3209
rect 2144 3193 2146 3209
rect 2296 3193 2298 3209
rect 2456 3193 2458 3209
rect 2624 3193 2626 3209
rect 2800 3193 2802 3209
rect 2976 3193 2978 3209
rect 3152 3193 3154 3209
rect 3328 3193 3330 3209
rect 3504 3193 3506 3209
rect 1894 3192 1900 3193
rect 1870 3189 1876 3190
rect 1870 3185 1871 3189
rect 1875 3185 1876 3189
rect 1894 3188 1895 3192
rect 1899 3188 1900 3192
rect 1894 3187 1900 3188
rect 2006 3192 2012 3193
rect 2006 3188 2007 3192
rect 2011 3188 2012 3192
rect 2006 3187 2012 3188
rect 2142 3192 2148 3193
rect 2142 3188 2143 3192
rect 2147 3188 2148 3192
rect 2142 3187 2148 3188
rect 2294 3192 2300 3193
rect 2294 3188 2295 3192
rect 2299 3188 2300 3192
rect 2294 3187 2300 3188
rect 2454 3192 2460 3193
rect 2454 3188 2455 3192
rect 2459 3188 2460 3192
rect 2454 3187 2460 3188
rect 2622 3192 2628 3193
rect 2622 3188 2623 3192
rect 2627 3188 2628 3192
rect 2622 3187 2628 3188
rect 2798 3192 2804 3193
rect 2798 3188 2799 3192
rect 2803 3188 2804 3192
rect 2798 3187 2804 3188
rect 2974 3192 2980 3193
rect 2974 3188 2975 3192
rect 2979 3188 2980 3192
rect 2974 3187 2980 3188
rect 3150 3192 3156 3193
rect 3150 3188 3151 3192
rect 3155 3188 3156 3192
rect 3150 3187 3156 3188
rect 3326 3192 3332 3193
rect 3326 3188 3327 3192
rect 3331 3188 3332 3192
rect 3326 3187 3332 3188
rect 3502 3192 3508 3193
rect 3502 3188 3503 3192
rect 3507 3188 3508 3192
rect 3592 3190 3594 3209
rect 3502 3187 3508 3188
rect 3590 3189 3596 3190
rect 1870 3184 1876 3185
rect 3590 3185 3591 3189
rect 3595 3185 3596 3189
rect 3590 3184 3596 3185
rect 1870 3172 1876 3173
rect 1870 3168 1871 3172
rect 1875 3168 1876 3172
rect 1870 3167 1876 3168
rect 3590 3172 3596 3173
rect 3590 3168 3591 3172
rect 3595 3168 3596 3172
rect 3590 3167 3596 3168
rect 111 3162 115 3163
rect 111 3157 115 3158
rect 143 3162 147 3163
rect 143 3157 147 3158
rect 175 3162 179 3163
rect 175 3157 179 3158
rect 279 3162 283 3163
rect 279 3157 283 3158
rect 319 3162 323 3163
rect 319 3157 323 3158
rect 423 3162 427 3163
rect 423 3157 427 3158
rect 463 3162 467 3163
rect 463 3157 467 3158
rect 583 3162 587 3163
rect 583 3157 587 3158
rect 607 3162 611 3163
rect 607 3157 611 3158
rect 743 3162 747 3163
rect 743 3157 747 3158
rect 871 3162 875 3163
rect 871 3157 875 3158
rect 903 3162 907 3163
rect 903 3157 907 3158
rect 991 3162 995 3163
rect 991 3157 995 3158
rect 1055 3162 1059 3163
rect 1055 3157 1059 3158
rect 1103 3162 1107 3163
rect 1103 3157 1107 3158
rect 1199 3162 1203 3163
rect 1199 3157 1203 3158
rect 1207 3162 1211 3163
rect 1207 3157 1211 3158
rect 1311 3162 1315 3163
rect 1311 3157 1315 3158
rect 1335 3162 1339 3163
rect 1335 3157 1339 3158
rect 1407 3162 1411 3163
rect 1407 3157 1411 3158
rect 1471 3162 1475 3163
rect 1471 3157 1475 3158
rect 1495 3162 1499 3163
rect 1495 3157 1499 3158
rect 1583 3162 1587 3163
rect 1583 3157 1587 3158
rect 1615 3162 1619 3163
rect 1615 3157 1619 3158
rect 1671 3162 1675 3163
rect 1671 3157 1675 3158
rect 1751 3162 1755 3163
rect 1751 3157 1755 3158
rect 1831 3162 1835 3163
rect 1831 3157 1835 3158
rect 112 3129 114 3157
rect 176 3147 178 3157
rect 320 3147 322 3157
rect 464 3147 466 3157
rect 608 3147 610 3157
rect 744 3147 746 3157
rect 872 3147 874 3157
rect 992 3147 994 3157
rect 1104 3147 1106 3157
rect 1208 3147 1210 3157
rect 1312 3147 1314 3157
rect 1408 3147 1410 3157
rect 1496 3147 1498 3157
rect 1584 3147 1586 3157
rect 1672 3147 1674 3157
rect 1752 3147 1754 3157
rect 174 3146 180 3147
rect 174 3142 175 3146
rect 179 3142 180 3146
rect 174 3141 180 3142
rect 318 3146 324 3147
rect 318 3142 319 3146
rect 323 3142 324 3146
rect 318 3141 324 3142
rect 462 3146 468 3147
rect 462 3142 463 3146
rect 467 3142 468 3146
rect 462 3141 468 3142
rect 606 3146 612 3147
rect 606 3142 607 3146
rect 611 3142 612 3146
rect 606 3141 612 3142
rect 742 3146 748 3147
rect 742 3142 743 3146
rect 747 3142 748 3146
rect 742 3141 748 3142
rect 870 3146 876 3147
rect 870 3142 871 3146
rect 875 3142 876 3146
rect 870 3141 876 3142
rect 990 3146 996 3147
rect 990 3142 991 3146
rect 995 3142 996 3146
rect 990 3141 996 3142
rect 1102 3146 1108 3147
rect 1102 3142 1103 3146
rect 1107 3142 1108 3146
rect 1102 3141 1108 3142
rect 1206 3146 1212 3147
rect 1206 3142 1207 3146
rect 1211 3142 1212 3146
rect 1206 3141 1212 3142
rect 1310 3146 1316 3147
rect 1310 3142 1311 3146
rect 1315 3142 1316 3146
rect 1310 3141 1316 3142
rect 1406 3146 1412 3147
rect 1406 3142 1407 3146
rect 1411 3142 1412 3146
rect 1406 3141 1412 3142
rect 1494 3146 1500 3147
rect 1494 3142 1495 3146
rect 1499 3142 1500 3146
rect 1494 3141 1500 3142
rect 1582 3146 1588 3147
rect 1582 3142 1583 3146
rect 1587 3142 1588 3146
rect 1582 3141 1588 3142
rect 1670 3146 1676 3147
rect 1670 3142 1671 3146
rect 1675 3142 1676 3146
rect 1670 3141 1676 3142
rect 1750 3146 1756 3147
rect 1750 3142 1751 3146
rect 1755 3142 1756 3146
rect 1750 3141 1756 3142
rect 1832 3129 1834 3157
rect 1872 3139 1874 3167
rect 1902 3154 1908 3155
rect 1902 3150 1903 3154
rect 1907 3150 1908 3154
rect 1902 3149 1908 3150
rect 2014 3154 2020 3155
rect 2014 3150 2015 3154
rect 2019 3150 2020 3154
rect 2014 3149 2020 3150
rect 2150 3154 2156 3155
rect 2150 3150 2151 3154
rect 2155 3150 2156 3154
rect 2150 3149 2156 3150
rect 2302 3154 2308 3155
rect 2302 3150 2303 3154
rect 2307 3150 2308 3154
rect 2302 3149 2308 3150
rect 2462 3154 2468 3155
rect 2462 3150 2463 3154
rect 2467 3150 2468 3154
rect 2462 3149 2468 3150
rect 2630 3154 2636 3155
rect 2630 3150 2631 3154
rect 2635 3150 2636 3154
rect 2630 3149 2636 3150
rect 2806 3154 2812 3155
rect 2806 3150 2807 3154
rect 2811 3150 2812 3154
rect 2806 3149 2812 3150
rect 2982 3154 2988 3155
rect 2982 3150 2983 3154
rect 2987 3150 2988 3154
rect 2982 3149 2988 3150
rect 3158 3154 3164 3155
rect 3158 3150 3159 3154
rect 3163 3150 3164 3154
rect 3158 3149 3164 3150
rect 3334 3154 3340 3155
rect 3334 3150 3335 3154
rect 3339 3150 3340 3154
rect 3334 3149 3340 3150
rect 3510 3154 3516 3155
rect 3510 3150 3511 3154
rect 3515 3150 3516 3154
rect 3510 3149 3516 3150
rect 1904 3139 1906 3149
rect 2016 3139 2018 3149
rect 2152 3139 2154 3149
rect 2304 3139 2306 3149
rect 2464 3139 2466 3149
rect 2632 3139 2634 3149
rect 2808 3139 2810 3149
rect 2984 3139 2986 3149
rect 3160 3139 3162 3149
rect 3336 3139 3338 3149
rect 3512 3139 3514 3149
rect 3592 3139 3594 3167
rect 1871 3138 1875 3139
rect 1871 3133 1875 3134
rect 1903 3138 1907 3139
rect 1903 3133 1907 3134
rect 2015 3138 2019 3139
rect 2015 3133 2019 3134
rect 2071 3138 2075 3139
rect 2071 3133 2075 3134
rect 2151 3138 2155 3139
rect 2151 3133 2155 3134
rect 2263 3138 2267 3139
rect 2263 3133 2267 3134
rect 2303 3138 2307 3139
rect 2303 3133 2307 3134
rect 2455 3138 2459 3139
rect 2455 3133 2459 3134
rect 2463 3138 2467 3139
rect 2463 3133 2467 3134
rect 2631 3138 2635 3139
rect 2631 3133 2635 3134
rect 2647 3138 2651 3139
rect 2647 3133 2651 3134
rect 2807 3138 2811 3139
rect 2807 3133 2811 3134
rect 2831 3138 2835 3139
rect 2831 3133 2835 3134
rect 2983 3138 2987 3139
rect 2983 3133 2987 3134
rect 3015 3138 3019 3139
rect 3015 3133 3019 3134
rect 3159 3138 3163 3139
rect 3159 3133 3163 3134
rect 3199 3138 3203 3139
rect 3199 3133 3203 3134
rect 3335 3138 3339 3139
rect 3335 3133 3339 3134
rect 3391 3138 3395 3139
rect 3391 3133 3395 3134
rect 3511 3138 3515 3139
rect 3511 3133 3515 3134
rect 3591 3138 3595 3139
rect 3591 3133 3595 3134
rect 110 3128 116 3129
rect 110 3124 111 3128
rect 115 3124 116 3128
rect 110 3123 116 3124
rect 1830 3128 1836 3129
rect 1830 3124 1831 3128
rect 1835 3124 1836 3128
rect 1830 3123 1836 3124
rect 110 3111 116 3112
rect 110 3107 111 3111
rect 115 3107 116 3111
rect 1830 3111 1836 3112
rect 110 3106 116 3107
rect 166 3108 172 3109
rect 112 3075 114 3106
rect 166 3104 167 3108
rect 171 3104 172 3108
rect 166 3103 172 3104
rect 310 3108 316 3109
rect 310 3104 311 3108
rect 315 3104 316 3108
rect 310 3103 316 3104
rect 454 3108 460 3109
rect 454 3104 455 3108
rect 459 3104 460 3108
rect 454 3103 460 3104
rect 598 3108 604 3109
rect 598 3104 599 3108
rect 603 3104 604 3108
rect 598 3103 604 3104
rect 734 3108 740 3109
rect 734 3104 735 3108
rect 739 3104 740 3108
rect 734 3103 740 3104
rect 862 3108 868 3109
rect 862 3104 863 3108
rect 867 3104 868 3108
rect 862 3103 868 3104
rect 982 3108 988 3109
rect 982 3104 983 3108
rect 987 3104 988 3108
rect 982 3103 988 3104
rect 1094 3108 1100 3109
rect 1094 3104 1095 3108
rect 1099 3104 1100 3108
rect 1094 3103 1100 3104
rect 1198 3108 1204 3109
rect 1198 3104 1199 3108
rect 1203 3104 1204 3108
rect 1198 3103 1204 3104
rect 1302 3108 1308 3109
rect 1302 3104 1303 3108
rect 1307 3104 1308 3108
rect 1302 3103 1308 3104
rect 1398 3108 1404 3109
rect 1398 3104 1399 3108
rect 1403 3104 1404 3108
rect 1398 3103 1404 3104
rect 1486 3108 1492 3109
rect 1486 3104 1487 3108
rect 1491 3104 1492 3108
rect 1486 3103 1492 3104
rect 1574 3108 1580 3109
rect 1574 3104 1575 3108
rect 1579 3104 1580 3108
rect 1574 3103 1580 3104
rect 1662 3108 1668 3109
rect 1662 3104 1663 3108
rect 1667 3104 1668 3108
rect 1662 3103 1668 3104
rect 1742 3108 1748 3109
rect 1742 3104 1743 3108
rect 1747 3104 1748 3108
rect 1830 3107 1831 3111
rect 1835 3107 1836 3111
rect 1830 3106 1836 3107
rect 1742 3103 1748 3104
rect 168 3075 170 3103
rect 312 3075 314 3103
rect 456 3075 458 3103
rect 600 3075 602 3103
rect 736 3075 738 3103
rect 864 3075 866 3103
rect 984 3075 986 3103
rect 1096 3075 1098 3103
rect 1200 3075 1202 3103
rect 1304 3075 1306 3103
rect 1400 3075 1402 3103
rect 1488 3075 1490 3103
rect 1576 3075 1578 3103
rect 1664 3075 1666 3103
rect 1744 3075 1746 3103
rect 1832 3075 1834 3106
rect 1872 3105 1874 3133
rect 1904 3123 1906 3133
rect 2072 3123 2074 3133
rect 2264 3123 2266 3133
rect 2456 3123 2458 3133
rect 2648 3123 2650 3133
rect 2832 3123 2834 3133
rect 3016 3123 3018 3133
rect 3200 3123 3202 3133
rect 3392 3123 3394 3133
rect 1902 3122 1908 3123
rect 1902 3118 1903 3122
rect 1907 3118 1908 3122
rect 1902 3117 1908 3118
rect 2070 3122 2076 3123
rect 2070 3118 2071 3122
rect 2075 3118 2076 3122
rect 2070 3117 2076 3118
rect 2262 3122 2268 3123
rect 2262 3118 2263 3122
rect 2267 3118 2268 3122
rect 2262 3117 2268 3118
rect 2454 3122 2460 3123
rect 2454 3118 2455 3122
rect 2459 3118 2460 3122
rect 2454 3117 2460 3118
rect 2646 3122 2652 3123
rect 2646 3118 2647 3122
rect 2651 3118 2652 3122
rect 2646 3117 2652 3118
rect 2830 3122 2836 3123
rect 2830 3118 2831 3122
rect 2835 3118 2836 3122
rect 2830 3117 2836 3118
rect 3014 3122 3020 3123
rect 3014 3118 3015 3122
rect 3019 3118 3020 3122
rect 3014 3117 3020 3118
rect 3198 3122 3204 3123
rect 3198 3118 3199 3122
rect 3203 3118 3204 3122
rect 3198 3117 3204 3118
rect 3390 3122 3396 3123
rect 3390 3118 3391 3122
rect 3395 3118 3396 3122
rect 3390 3117 3396 3118
rect 3592 3105 3594 3133
rect 1870 3104 1876 3105
rect 1870 3100 1871 3104
rect 1875 3100 1876 3104
rect 1870 3099 1876 3100
rect 3590 3104 3596 3105
rect 3590 3100 3591 3104
rect 3595 3100 3596 3104
rect 3590 3099 3596 3100
rect 1870 3087 1876 3088
rect 1870 3083 1871 3087
rect 1875 3083 1876 3087
rect 3590 3087 3596 3088
rect 1870 3082 1876 3083
rect 1894 3084 1900 3085
rect 111 3074 115 3075
rect 111 3069 115 3070
rect 135 3074 139 3075
rect 135 3069 139 3070
rect 167 3074 171 3075
rect 167 3069 171 3070
rect 223 3074 227 3075
rect 223 3069 227 3070
rect 311 3074 315 3075
rect 311 3069 315 3070
rect 327 3074 331 3075
rect 327 3069 331 3070
rect 439 3074 443 3075
rect 439 3069 443 3070
rect 455 3074 459 3075
rect 455 3069 459 3070
rect 551 3074 555 3075
rect 551 3069 555 3070
rect 599 3074 603 3075
rect 599 3069 603 3070
rect 663 3074 667 3075
rect 663 3069 667 3070
rect 735 3074 739 3075
rect 735 3069 739 3070
rect 863 3074 867 3075
rect 863 3069 867 3070
rect 983 3074 987 3075
rect 983 3069 987 3070
rect 1095 3074 1099 3075
rect 1095 3069 1099 3070
rect 1199 3074 1203 3075
rect 1199 3069 1203 3070
rect 1303 3074 1307 3075
rect 1303 3069 1307 3070
rect 1399 3074 1403 3075
rect 1399 3069 1403 3070
rect 1487 3074 1491 3075
rect 1487 3069 1491 3070
rect 1575 3074 1579 3075
rect 1575 3069 1579 3070
rect 1663 3074 1667 3075
rect 1663 3069 1667 3070
rect 1743 3074 1747 3075
rect 1743 3069 1747 3070
rect 1831 3074 1835 3075
rect 1831 3069 1835 3070
rect 112 3050 114 3069
rect 136 3053 138 3069
rect 224 3053 226 3069
rect 328 3053 330 3069
rect 440 3053 442 3069
rect 552 3053 554 3069
rect 664 3053 666 3069
rect 134 3052 140 3053
rect 110 3049 116 3050
rect 110 3045 111 3049
rect 115 3045 116 3049
rect 134 3048 135 3052
rect 139 3048 140 3052
rect 134 3047 140 3048
rect 222 3052 228 3053
rect 222 3048 223 3052
rect 227 3048 228 3052
rect 222 3047 228 3048
rect 326 3052 332 3053
rect 326 3048 327 3052
rect 331 3048 332 3052
rect 326 3047 332 3048
rect 438 3052 444 3053
rect 438 3048 439 3052
rect 443 3048 444 3052
rect 438 3047 444 3048
rect 550 3052 556 3053
rect 550 3048 551 3052
rect 555 3048 556 3052
rect 550 3047 556 3048
rect 662 3052 668 3053
rect 662 3048 663 3052
rect 667 3048 668 3052
rect 1832 3050 1834 3069
rect 1872 3051 1874 3082
rect 1894 3080 1895 3084
rect 1899 3080 1900 3084
rect 1894 3079 1900 3080
rect 2062 3084 2068 3085
rect 2062 3080 2063 3084
rect 2067 3080 2068 3084
rect 2062 3079 2068 3080
rect 2254 3084 2260 3085
rect 2254 3080 2255 3084
rect 2259 3080 2260 3084
rect 2254 3079 2260 3080
rect 2446 3084 2452 3085
rect 2446 3080 2447 3084
rect 2451 3080 2452 3084
rect 2446 3079 2452 3080
rect 2638 3084 2644 3085
rect 2638 3080 2639 3084
rect 2643 3080 2644 3084
rect 2638 3079 2644 3080
rect 2822 3084 2828 3085
rect 2822 3080 2823 3084
rect 2827 3080 2828 3084
rect 2822 3079 2828 3080
rect 3006 3084 3012 3085
rect 3006 3080 3007 3084
rect 3011 3080 3012 3084
rect 3006 3079 3012 3080
rect 3190 3084 3196 3085
rect 3190 3080 3191 3084
rect 3195 3080 3196 3084
rect 3190 3079 3196 3080
rect 3382 3084 3388 3085
rect 3382 3080 3383 3084
rect 3387 3080 3388 3084
rect 3590 3083 3591 3087
rect 3595 3083 3596 3087
rect 3590 3082 3596 3083
rect 3382 3079 3388 3080
rect 1896 3051 1898 3079
rect 2064 3051 2066 3079
rect 2256 3051 2258 3079
rect 2448 3051 2450 3079
rect 2640 3051 2642 3079
rect 2824 3051 2826 3079
rect 3008 3051 3010 3079
rect 3192 3051 3194 3079
rect 3384 3051 3386 3079
rect 3592 3051 3594 3082
rect 1871 3050 1875 3051
rect 662 3047 668 3048
rect 1830 3049 1836 3050
rect 110 3044 116 3045
rect 1830 3045 1831 3049
rect 1835 3045 1836 3049
rect 1871 3045 1875 3046
rect 1895 3050 1899 3051
rect 1895 3045 1899 3046
rect 2063 3050 2067 3051
rect 2063 3045 2067 3046
rect 2199 3050 2203 3051
rect 2199 3045 2203 3046
rect 2255 3050 2259 3051
rect 2255 3045 2259 3046
rect 2335 3050 2339 3051
rect 2335 3045 2339 3046
rect 2447 3050 2451 3051
rect 2447 3045 2451 3046
rect 2479 3050 2483 3051
rect 2479 3045 2483 3046
rect 2623 3050 2627 3051
rect 2623 3045 2627 3046
rect 2639 3050 2643 3051
rect 2639 3045 2643 3046
rect 2767 3050 2771 3051
rect 2767 3045 2771 3046
rect 2823 3050 2827 3051
rect 2823 3045 2827 3046
rect 2903 3050 2907 3051
rect 2903 3045 2907 3046
rect 3007 3050 3011 3051
rect 3007 3045 3011 3046
rect 3039 3050 3043 3051
rect 3039 3045 3043 3046
rect 3183 3050 3187 3051
rect 3183 3045 3187 3046
rect 3191 3050 3195 3051
rect 3191 3045 3195 3046
rect 3327 3050 3331 3051
rect 3327 3045 3331 3046
rect 3383 3050 3387 3051
rect 3383 3045 3387 3046
rect 3591 3050 3595 3051
rect 3591 3045 3595 3046
rect 1830 3044 1836 3045
rect 110 3032 116 3033
rect 110 3028 111 3032
rect 115 3028 116 3032
rect 110 3027 116 3028
rect 1830 3032 1836 3033
rect 1830 3028 1831 3032
rect 1835 3028 1836 3032
rect 1830 3027 1836 3028
rect 112 2987 114 3027
rect 142 3014 148 3015
rect 142 3010 143 3014
rect 147 3010 148 3014
rect 142 3009 148 3010
rect 230 3014 236 3015
rect 230 3010 231 3014
rect 235 3010 236 3014
rect 230 3009 236 3010
rect 334 3014 340 3015
rect 334 3010 335 3014
rect 339 3010 340 3014
rect 334 3009 340 3010
rect 446 3014 452 3015
rect 446 3010 447 3014
rect 451 3010 452 3014
rect 446 3009 452 3010
rect 558 3014 564 3015
rect 558 3010 559 3014
rect 563 3010 564 3014
rect 558 3009 564 3010
rect 670 3014 676 3015
rect 670 3010 671 3014
rect 675 3010 676 3014
rect 670 3009 676 3010
rect 144 2987 146 3009
rect 232 2987 234 3009
rect 336 2987 338 3009
rect 448 2987 450 3009
rect 560 2987 562 3009
rect 672 2987 674 3009
rect 1832 2987 1834 3027
rect 1872 3026 1874 3045
rect 2200 3029 2202 3045
rect 2336 3029 2338 3045
rect 2480 3029 2482 3045
rect 2624 3029 2626 3045
rect 2768 3029 2770 3045
rect 2904 3029 2906 3045
rect 3040 3029 3042 3045
rect 3184 3029 3186 3045
rect 3328 3029 3330 3045
rect 2198 3028 2204 3029
rect 1870 3025 1876 3026
rect 1870 3021 1871 3025
rect 1875 3021 1876 3025
rect 2198 3024 2199 3028
rect 2203 3024 2204 3028
rect 2198 3023 2204 3024
rect 2334 3028 2340 3029
rect 2334 3024 2335 3028
rect 2339 3024 2340 3028
rect 2334 3023 2340 3024
rect 2478 3028 2484 3029
rect 2478 3024 2479 3028
rect 2483 3024 2484 3028
rect 2478 3023 2484 3024
rect 2622 3028 2628 3029
rect 2622 3024 2623 3028
rect 2627 3024 2628 3028
rect 2622 3023 2628 3024
rect 2766 3028 2772 3029
rect 2766 3024 2767 3028
rect 2771 3024 2772 3028
rect 2766 3023 2772 3024
rect 2902 3028 2908 3029
rect 2902 3024 2903 3028
rect 2907 3024 2908 3028
rect 2902 3023 2908 3024
rect 3038 3028 3044 3029
rect 3038 3024 3039 3028
rect 3043 3024 3044 3028
rect 3038 3023 3044 3024
rect 3182 3028 3188 3029
rect 3182 3024 3183 3028
rect 3187 3024 3188 3028
rect 3182 3023 3188 3024
rect 3326 3028 3332 3029
rect 3326 3024 3327 3028
rect 3331 3024 3332 3028
rect 3592 3026 3594 3045
rect 3326 3023 3332 3024
rect 3590 3025 3596 3026
rect 1870 3020 1876 3021
rect 3590 3021 3591 3025
rect 3595 3021 3596 3025
rect 3590 3020 3596 3021
rect 1870 3008 1876 3009
rect 1870 3004 1871 3008
rect 1875 3004 1876 3008
rect 1870 3003 1876 3004
rect 3590 3008 3596 3009
rect 3590 3004 3591 3008
rect 3595 3004 3596 3008
rect 3590 3003 3596 3004
rect 111 2986 115 2987
rect 111 2981 115 2982
rect 143 2986 147 2987
rect 143 2981 147 2982
rect 159 2986 163 2987
rect 159 2981 163 2982
rect 231 2986 235 2987
rect 231 2981 235 2982
rect 319 2986 323 2987
rect 319 2981 323 2982
rect 335 2986 339 2987
rect 335 2981 339 2982
rect 447 2986 451 2987
rect 447 2981 451 2982
rect 487 2986 491 2987
rect 487 2981 491 2982
rect 559 2986 563 2987
rect 559 2981 563 2982
rect 647 2986 651 2987
rect 647 2981 651 2982
rect 671 2986 675 2987
rect 671 2981 675 2982
rect 799 2986 803 2987
rect 799 2981 803 2982
rect 943 2986 947 2987
rect 943 2981 947 2982
rect 1079 2986 1083 2987
rect 1079 2981 1083 2982
rect 1199 2986 1203 2987
rect 1199 2981 1203 2982
rect 1311 2986 1315 2987
rect 1311 2981 1315 2982
rect 1423 2986 1427 2987
rect 1423 2981 1427 2982
rect 1535 2986 1539 2987
rect 1535 2981 1539 2982
rect 1647 2986 1651 2987
rect 1647 2981 1651 2982
rect 1831 2986 1835 2987
rect 1831 2981 1835 2982
rect 112 2953 114 2981
rect 160 2971 162 2981
rect 320 2971 322 2981
rect 488 2971 490 2981
rect 648 2971 650 2981
rect 800 2971 802 2981
rect 944 2971 946 2981
rect 1080 2971 1082 2981
rect 1200 2971 1202 2981
rect 1312 2971 1314 2981
rect 1424 2971 1426 2981
rect 1536 2971 1538 2981
rect 1648 2971 1650 2981
rect 158 2970 164 2971
rect 158 2966 159 2970
rect 163 2966 164 2970
rect 158 2965 164 2966
rect 318 2970 324 2971
rect 318 2966 319 2970
rect 323 2966 324 2970
rect 318 2965 324 2966
rect 486 2970 492 2971
rect 486 2966 487 2970
rect 491 2966 492 2970
rect 486 2965 492 2966
rect 646 2970 652 2971
rect 646 2966 647 2970
rect 651 2966 652 2970
rect 646 2965 652 2966
rect 798 2970 804 2971
rect 798 2966 799 2970
rect 803 2966 804 2970
rect 798 2965 804 2966
rect 942 2970 948 2971
rect 942 2966 943 2970
rect 947 2966 948 2970
rect 942 2965 948 2966
rect 1078 2970 1084 2971
rect 1078 2966 1079 2970
rect 1083 2966 1084 2970
rect 1078 2965 1084 2966
rect 1198 2970 1204 2971
rect 1198 2966 1199 2970
rect 1203 2966 1204 2970
rect 1198 2965 1204 2966
rect 1310 2970 1316 2971
rect 1310 2966 1311 2970
rect 1315 2966 1316 2970
rect 1310 2965 1316 2966
rect 1422 2970 1428 2971
rect 1422 2966 1423 2970
rect 1427 2966 1428 2970
rect 1422 2965 1428 2966
rect 1534 2970 1540 2971
rect 1534 2966 1535 2970
rect 1539 2966 1540 2970
rect 1534 2965 1540 2966
rect 1646 2970 1652 2971
rect 1646 2966 1647 2970
rect 1651 2966 1652 2970
rect 1646 2965 1652 2966
rect 1832 2953 1834 2981
rect 1872 2963 1874 3003
rect 2206 2990 2212 2991
rect 2206 2986 2207 2990
rect 2211 2986 2212 2990
rect 2206 2985 2212 2986
rect 2342 2990 2348 2991
rect 2342 2986 2343 2990
rect 2347 2986 2348 2990
rect 2342 2985 2348 2986
rect 2486 2990 2492 2991
rect 2486 2986 2487 2990
rect 2491 2986 2492 2990
rect 2486 2985 2492 2986
rect 2630 2990 2636 2991
rect 2630 2986 2631 2990
rect 2635 2986 2636 2990
rect 2630 2985 2636 2986
rect 2774 2990 2780 2991
rect 2774 2986 2775 2990
rect 2779 2986 2780 2990
rect 2774 2985 2780 2986
rect 2910 2990 2916 2991
rect 2910 2986 2911 2990
rect 2915 2986 2916 2990
rect 2910 2985 2916 2986
rect 3046 2990 3052 2991
rect 3046 2986 3047 2990
rect 3051 2986 3052 2990
rect 3046 2985 3052 2986
rect 3190 2990 3196 2991
rect 3190 2986 3191 2990
rect 3195 2986 3196 2990
rect 3190 2985 3196 2986
rect 3334 2990 3340 2991
rect 3334 2986 3335 2990
rect 3339 2986 3340 2990
rect 3334 2985 3340 2986
rect 2208 2963 2210 2985
rect 2344 2963 2346 2985
rect 2488 2963 2490 2985
rect 2632 2963 2634 2985
rect 2776 2963 2778 2985
rect 2912 2963 2914 2985
rect 3048 2963 3050 2985
rect 3192 2963 3194 2985
rect 3336 2963 3338 2985
rect 3592 2963 3594 3003
rect 1871 2962 1875 2963
rect 1871 2957 1875 2958
rect 2127 2962 2131 2963
rect 2127 2957 2131 2958
rect 2207 2962 2211 2963
rect 2207 2957 2211 2958
rect 2287 2962 2291 2963
rect 2287 2957 2291 2958
rect 2343 2962 2347 2963
rect 2343 2957 2347 2958
rect 2367 2962 2371 2963
rect 2367 2957 2371 2958
rect 2447 2962 2451 2963
rect 2447 2957 2451 2958
rect 2487 2962 2491 2963
rect 2487 2957 2491 2958
rect 2527 2962 2531 2963
rect 2527 2957 2531 2958
rect 2607 2962 2611 2963
rect 2607 2957 2611 2958
rect 2631 2962 2635 2963
rect 2631 2957 2635 2958
rect 2695 2962 2699 2963
rect 2695 2957 2699 2958
rect 2775 2962 2779 2963
rect 2775 2957 2779 2958
rect 2791 2962 2795 2963
rect 2791 2957 2795 2958
rect 2911 2962 2915 2963
rect 2911 2957 2915 2958
rect 3039 2962 3043 2963
rect 3039 2957 3043 2958
rect 3047 2962 3051 2963
rect 3047 2957 3051 2958
rect 3183 2962 3187 2963
rect 3183 2957 3187 2958
rect 3191 2962 3195 2963
rect 3191 2957 3195 2958
rect 3335 2962 3339 2963
rect 3335 2957 3339 2958
rect 3495 2962 3499 2963
rect 3495 2957 3499 2958
rect 3591 2962 3595 2963
rect 3591 2957 3595 2958
rect 110 2952 116 2953
rect 110 2948 111 2952
rect 115 2948 116 2952
rect 110 2947 116 2948
rect 1830 2952 1836 2953
rect 1830 2948 1831 2952
rect 1835 2948 1836 2952
rect 1830 2947 1836 2948
rect 110 2935 116 2936
rect 110 2931 111 2935
rect 115 2931 116 2935
rect 1830 2935 1836 2936
rect 110 2930 116 2931
rect 150 2932 156 2933
rect 112 2911 114 2930
rect 150 2928 151 2932
rect 155 2928 156 2932
rect 150 2927 156 2928
rect 310 2932 316 2933
rect 310 2928 311 2932
rect 315 2928 316 2932
rect 310 2927 316 2928
rect 478 2932 484 2933
rect 478 2928 479 2932
rect 483 2928 484 2932
rect 478 2927 484 2928
rect 638 2932 644 2933
rect 638 2928 639 2932
rect 643 2928 644 2932
rect 638 2927 644 2928
rect 790 2932 796 2933
rect 790 2928 791 2932
rect 795 2928 796 2932
rect 790 2927 796 2928
rect 934 2932 940 2933
rect 934 2928 935 2932
rect 939 2928 940 2932
rect 934 2927 940 2928
rect 1070 2932 1076 2933
rect 1070 2928 1071 2932
rect 1075 2928 1076 2932
rect 1070 2927 1076 2928
rect 1190 2932 1196 2933
rect 1190 2928 1191 2932
rect 1195 2928 1196 2932
rect 1190 2927 1196 2928
rect 1302 2932 1308 2933
rect 1302 2928 1303 2932
rect 1307 2928 1308 2932
rect 1302 2927 1308 2928
rect 1414 2932 1420 2933
rect 1414 2928 1415 2932
rect 1419 2928 1420 2932
rect 1414 2927 1420 2928
rect 1526 2932 1532 2933
rect 1526 2928 1527 2932
rect 1531 2928 1532 2932
rect 1526 2927 1532 2928
rect 1638 2932 1644 2933
rect 1638 2928 1639 2932
rect 1643 2928 1644 2932
rect 1830 2931 1831 2935
rect 1835 2931 1836 2935
rect 1830 2930 1836 2931
rect 1638 2927 1644 2928
rect 152 2911 154 2927
rect 312 2911 314 2927
rect 480 2911 482 2927
rect 640 2911 642 2927
rect 792 2911 794 2927
rect 936 2911 938 2927
rect 1072 2911 1074 2927
rect 1192 2911 1194 2927
rect 1304 2911 1306 2927
rect 1416 2911 1418 2927
rect 1528 2911 1530 2927
rect 1640 2911 1642 2927
rect 1832 2911 1834 2930
rect 1872 2929 1874 2957
rect 2128 2947 2130 2957
rect 2208 2947 2210 2957
rect 2288 2947 2290 2957
rect 2368 2947 2370 2957
rect 2448 2947 2450 2957
rect 2528 2947 2530 2957
rect 2608 2947 2610 2957
rect 2696 2947 2698 2957
rect 2792 2947 2794 2957
rect 2912 2947 2914 2957
rect 3040 2947 3042 2957
rect 3184 2947 3186 2957
rect 3336 2947 3338 2957
rect 3496 2947 3498 2957
rect 2126 2946 2132 2947
rect 2126 2942 2127 2946
rect 2131 2942 2132 2946
rect 2126 2941 2132 2942
rect 2206 2946 2212 2947
rect 2206 2942 2207 2946
rect 2211 2942 2212 2946
rect 2206 2941 2212 2942
rect 2286 2946 2292 2947
rect 2286 2942 2287 2946
rect 2291 2942 2292 2946
rect 2286 2941 2292 2942
rect 2366 2946 2372 2947
rect 2366 2942 2367 2946
rect 2371 2942 2372 2946
rect 2366 2941 2372 2942
rect 2446 2946 2452 2947
rect 2446 2942 2447 2946
rect 2451 2942 2452 2946
rect 2446 2941 2452 2942
rect 2526 2946 2532 2947
rect 2526 2942 2527 2946
rect 2531 2942 2532 2946
rect 2526 2941 2532 2942
rect 2606 2946 2612 2947
rect 2606 2942 2607 2946
rect 2611 2942 2612 2946
rect 2606 2941 2612 2942
rect 2694 2946 2700 2947
rect 2694 2942 2695 2946
rect 2699 2942 2700 2946
rect 2694 2941 2700 2942
rect 2790 2946 2796 2947
rect 2790 2942 2791 2946
rect 2795 2942 2796 2946
rect 2790 2941 2796 2942
rect 2910 2946 2916 2947
rect 2910 2942 2911 2946
rect 2915 2942 2916 2946
rect 2910 2941 2916 2942
rect 3038 2946 3044 2947
rect 3038 2942 3039 2946
rect 3043 2942 3044 2946
rect 3038 2941 3044 2942
rect 3182 2946 3188 2947
rect 3182 2942 3183 2946
rect 3187 2942 3188 2946
rect 3182 2941 3188 2942
rect 3334 2946 3340 2947
rect 3334 2942 3335 2946
rect 3339 2942 3340 2946
rect 3334 2941 3340 2942
rect 3494 2946 3500 2947
rect 3494 2942 3495 2946
rect 3499 2942 3500 2946
rect 3494 2941 3500 2942
rect 3592 2929 3594 2957
rect 1870 2928 1876 2929
rect 1870 2924 1871 2928
rect 1875 2924 1876 2928
rect 1870 2923 1876 2924
rect 3590 2928 3596 2929
rect 3590 2924 3591 2928
rect 3595 2924 3596 2928
rect 3590 2923 3596 2924
rect 1870 2911 1876 2912
rect 111 2910 115 2911
rect 111 2905 115 2906
rect 151 2910 155 2911
rect 151 2905 155 2906
rect 311 2910 315 2911
rect 311 2905 315 2906
rect 471 2910 475 2911
rect 471 2905 475 2906
rect 479 2910 483 2911
rect 479 2905 483 2906
rect 631 2910 635 2911
rect 631 2905 635 2906
rect 639 2910 643 2911
rect 639 2905 643 2906
rect 783 2910 787 2911
rect 783 2905 787 2906
rect 791 2910 795 2911
rect 791 2905 795 2906
rect 927 2910 931 2911
rect 927 2905 931 2906
rect 935 2910 939 2911
rect 935 2905 939 2906
rect 1055 2910 1059 2911
rect 1055 2905 1059 2906
rect 1071 2910 1075 2911
rect 1071 2905 1075 2906
rect 1175 2910 1179 2911
rect 1175 2905 1179 2906
rect 1191 2910 1195 2911
rect 1191 2905 1195 2906
rect 1287 2910 1291 2911
rect 1287 2905 1291 2906
rect 1303 2910 1307 2911
rect 1303 2905 1307 2906
rect 1391 2910 1395 2911
rect 1391 2905 1395 2906
rect 1415 2910 1419 2911
rect 1415 2905 1419 2906
rect 1487 2910 1491 2911
rect 1487 2905 1491 2906
rect 1527 2910 1531 2911
rect 1527 2905 1531 2906
rect 1591 2910 1595 2911
rect 1591 2905 1595 2906
rect 1639 2910 1643 2911
rect 1639 2905 1643 2906
rect 1695 2910 1699 2911
rect 1695 2905 1699 2906
rect 1831 2910 1835 2911
rect 1870 2907 1871 2911
rect 1875 2907 1876 2911
rect 3590 2911 3596 2912
rect 1870 2906 1876 2907
rect 2118 2908 2124 2909
rect 1831 2905 1835 2906
rect 112 2886 114 2905
rect 152 2889 154 2905
rect 312 2889 314 2905
rect 472 2889 474 2905
rect 632 2889 634 2905
rect 784 2889 786 2905
rect 928 2889 930 2905
rect 1056 2889 1058 2905
rect 1176 2889 1178 2905
rect 1288 2889 1290 2905
rect 1392 2889 1394 2905
rect 1488 2889 1490 2905
rect 1592 2889 1594 2905
rect 1696 2889 1698 2905
rect 150 2888 156 2889
rect 110 2885 116 2886
rect 110 2881 111 2885
rect 115 2881 116 2885
rect 150 2884 151 2888
rect 155 2884 156 2888
rect 150 2883 156 2884
rect 310 2888 316 2889
rect 310 2884 311 2888
rect 315 2884 316 2888
rect 310 2883 316 2884
rect 470 2888 476 2889
rect 470 2884 471 2888
rect 475 2884 476 2888
rect 470 2883 476 2884
rect 630 2888 636 2889
rect 630 2884 631 2888
rect 635 2884 636 2888
rect 630 2883 636 2884
rect 782 2888 788 2889
rect 782 2884 783 2888
rect 787 2884 788 2888
rect 782 2883 788 2884
rect 926 2888 932 2889
rect 926 2884 927 2888
rect 931 2884 932 2888
rect 926 2883 932 2884
rect 1054 2888 1060 2889
rect 1054 2884 1055 2888
rect 1059 2884 1060 2888
rect 1054 2883 1060 2884
rect 1174 2888 1180 2889
rect 1174 2884 1175 2888
rect 1179 2884 1180 2888
rect 1174 2883 1180 2884
rect 1286 2888 1292 2889
rect 1286 2884 1287 2888
rect 1291 2884 1292 2888
rect 1286 2883 1292 2884
rect 1390 2888 1396 2889
rect 1390 2884 1391 2888
rect 1395 2884 1396 2888
rect 1390 2883 1396 2884
rect 1486 2888 1492 2889
rect 1486 2884 1487 2888
rect 1491 2884 1492 2888
rect 1486 2883 1492 2884
rect 1590 2888 1596 2889
rect 1590 2884 1591 2888
rect 1595 2884 1596 2888
rect 1590 2883 1596 2884
rect 1694 2888 1700 2889
rect 1694 2884 1695 2888
rect 1699 2884 1700 2888
rect 1832 2886 1834 2905
rect 1872 2887 1874 2906
rect 2118 2904 2119 2908
rect 2123 2904 2124 2908
rect 2118 2903 2124 2904
rect 2198 2908 2204 2909
rect 2198 2904 2199 2908
rect 2203 2904 2204 2908
rect 2198 2903 2204 2904
rect 2278 2908 2284 2909
rect 2278 2904 2279 2908
rect 2283 2904 2284 2908
rect 2278 2903 2284 2904
rect 2358 2908 2364 2909
rect 2358 2904 2359 2908
rect 2363 2904 2364 2908
rect 2358 2903 2364 2904
rect 2438 2908 2444 2909
rect 2438 2904 2439 2908
rect 2443 2904 2444 2908
rect 2438 2903 2444 2904
rect 2518 2908 2524 2909
rect 2518 2904 2519 2908
rect 2523 2904 2524 2908
rect 2518 2903 2524 2904
rect 2598 2908 2604 2909
rect 2598 2904 2599 2908
rect 2603 2904 2604 2908
rect 2598 2903 2604 2904
rect 2686 2908 2692 2909
rect 2686 2904 2687 2908
rect 2691 2904 2692 2908
rect 2686 2903 2692 2904
rect 2782 2908 2788 2909
rect 2782 2904 2783 2908
rect 2787 2904 2788 2908
rect 2782 2903 2788 2904
rect 2902 2908 2908 2909
rect 2902 2904 2903 2908
rect 2907 2904 2908 2908
rect 2902 2903 2908 2904
rect 3030 2908 3036 2909
rect 3030 2904 3031 2908
rect 3035 2904 3036 2908
rect 3030 2903 3036 2904
rect 3174 2908 3180 2909
rect 3174 2904 3175 2908
rect 3179 2904 3180 2908
rect 3174 2903 3180 2904
rect 3326 2908 3332 2909
rect 3326 2904 3327 2908
rect 3331 2904 3332 2908
rect 3326 2903 3332 2904
rect 3486 2908 3492 2909
rect 3486 2904 3487 2908
rect 3491 2904 3492 2908
rect 3590 2907 3591 2911
rect 3595 2907 3596 2911
rect 3590 2906 3596 2907
rect 3486 2903 3492 2904
rect 2120 2887 2122 2903
rect 2200 2887 2202 2903
rect 2280 2887 2282 2903
rect 2360 2887 2362 2903
rect 2440 2887 2442 2903
rect 2520 2887 2522 2903
rect 2600 2887 2602 2903
rect 2688 2887 2690 2903
rect 2784 2887 2786 2903
rect 2904 2887 2906 2903
rect 3032 2887 3034 2903
rect 3176 2887 3178 2903
rect 3328 2887 3330 2903
rect 3488 2887 3490 2903
rect 3592 2887 3594 2906
rect 1871 2886 1875 2887
rect 1694 2883 1700 2884
rect 1830 2885 1836 2886
rect 110 2880 116 2881
rect 1830 2881 1831 2885
rect 1835 2881 1836 2885
rect 1871 2881 1875 2882
rect 2047 2886 2051 2887
rect 2047 2881 2051 2882
rect 2119 2886 2123 2887
rect 2119 2881 2123 2882
rect 2135 2886 2139 2887
rect 2135 2881 2139 2882
rect 2199 2886 2203 2887
rect 2199 2881 2203 2882
rect 2239 2886 2243 2887
rect 2239 2881 2243 2882
rect 2279 2886 2283 2887
rect 2279 2881 2283 2882
rect 2343 2886 2347 2887
rect 2343 2881 2347 2882
rect 2359 2886 2363 2887
rect 2359 2881 2363 2882
rect 2439 2886 2443 2887
rect 2439 2881 2443 2882
rect 2463 2886 2467 2887
rect 2463 2881 2467 2882
rect 2519 2886 2523 2887
rect 2519 2881 2523 2882
rect 2591 2886 2595 2887
rect 2591 2881 2595 2882
rect 2599 2886 2603 2887
rect 2599 2881 2603 2882
rect 2687 2886 2691 2887
rect 2687 2881 2691 2882
rect 2727 2886 2731 2887
rect 2727 2881 2731 2882
rect 2783 2886 2787 2887
rect 2783 2881 2787 2882
rect 2879 2886 2883 2887
rect 2879 2881 2883 2882
rect 2903 2886 2907 2887
rect 2903 2881 2907 2882
rect 3031 2886 3035 2887
rect 3031 2881 3035 2882
rect 3175 2886 3179 2887
rect 3175 2881 3179 2882
rect 3191 2886 3195 2887
rect 3191 2881 3195 2882
rect 3327 2886 3331 2887
rect 3327 2881 3331 2882
rect 3359 2886 3363 2887
rect 3359 2881 3363 2882
rect 3487 2886 3491 2887
rect 3487 2881 3491 2882
rect 3503 2886 3507 2887
rect 3503 2881 3507 2882
rect 3591 2886 3595 2887
rect 3591 2881 3595 2882
rect 1830 2880 1836 2881
rect 110 2868 116 2869
rect 110 2864 111 2868
rect 115 2864 116 2868
rect 110 2863 116 2864
rect 1830 2868 1836 2869
rect 1830 2864 1831 2868
rect 1835 2864 1836 2868
rect 1830 2863 1836 2864
rect 112 2831 114 2863
rect 158 2850 164 2851
rect 158 2846 159 2850
rect 163 2846 164 2850
rect 158 2845 164 2846
rect 318 2850 324 2851
rect 318 2846 319 2850
rect 323 2846 324 2850
rect 318 2845 324 2846
rect 478 2850 484 2851
rect 478 2846 479 2850
rect 483 2846 484 2850
rect 478 2845 484 2846
rect 638 2850 644 2851
rect 638 2846 639 2850
rect 643 2846 644 2850
rect 638 2845 644 2846
rect 790 2850 796 2851
rect 790 2846 791 2850
rect 795 2846 796 2850
rect 790 2845 796 2846
rect 934 2850 940 2851
rect 934 2846 935 2850
rect 939 2846 940 2850
rect 934 2845 940 2846
rect 1062 2850 1068 2851
rect 1062 2846 1063 2850
rect 1067 2846 1068 2850
rect 1062 2845 1068 2846
rect 1182 2850 1188 2851
rect 1182 2846 1183 2850
rect 1187 2846 1188 2850
rect 1182 2845 1188 2846
rect 1294 2850 1300 2851
rect 1294 2846 1295 2850
rect 1299 2846 1300 2850
rect 1294 2845 1300 2846
rect 1398 2850 1404 2851
rect 1398 2846 1399 2850
rect 1403 2846 1404 2850
rect 1398 2845 1404 2846
rect 1494 2850 1500 2851
rect 1494 2846 1495 2850
rect 1499 2846 1500 2850
rect 1494 2845 1500 2846
rect 1598 2850 1604 2851
rect 1598 2846 1599 2850
rect 1603 2846 1604 2850
rect 1598 2845 1604 2846
rect 1702 2850 1708 2851
rect 1702 2846 1703 2850
rect 1707 2846 1708 2850
rect 1702 2845 1708 2846
rect 160 2831 162 2845
rect 320 2831 322 2845
rect 480 2831 482 2845
rect 640 2831 642 2845
rect 792 2831 794 2845
rect 936 2831 938 2845
rect 1064 2831 1066 2845
rect 1184 2831 1186 2845
rect 1296 2831 1298 2845
rect 1400 2831 1402 2845
rect 1496 2831 1498 2845
rect 1600 2831 1602 2845
rect 1704 2831 1706 2845
rect 1832 2831 1834 2863
rect 1872 2862 1874 2881
rect 2048 2865 2050 2881
rect 2136 2865 2138 2881
rect 2240 2865 2242 2881
rect 2344 2865 2346 2881
rect 2464 2865 2466 2881
rect 2592 2865 2594 2881
rect 2728 2865 2730 2881
rect 2880 2865 2882 2881
rect 3032 2865 3034 2881
rect 3192 2865 3194 2881
rect 3360 2865 3362 2881
rect 3504 2865 3506 2881
rect 2046 2864 2052 2865
rect 1870 2861 1876 2862
rect 1870 2857 1871 2861
rect 1875 2857 1876 2861
rect 2046 2860 2047 2864
rect 2051 2860 2052 2864
rect 2046 2859 2052 2860
rect 2134 2864 2140 2865
rect 2134 2860 2135 2864
rect 2139 2860 2140 2864
rect 2134 2859 2140 2860
rect 2238 2864 2244 2865
rect 2238 2860 2239 2864
rect 2243 2860 2244 2864
rect 2238 2859 2244 2860
rect 2342 2864 2348 2865
rect 2342 2860 2343 2864
rect 2347 2860 2348 2864
rect 2342 2859 2348 2860
rect 2462 2864 2468 2865
rect 2462 2860 2463 2864
rect 2467 2860 2468 2864
rect 2462 2859 2468 2860
rect 2590 2864 2596 2865
rect 2590 2860 2591 2864
rect 2595 2860 2596 2864
rect 2590 2859 2596 2860
rect 2726 2864 2732 2865
rect 2726 2860 2727 2864
rect 2731 2860 2732 2864
rect 2726 2859 2732 2860
rect 2878 2864 2884 2865
rect 2878 2860 2879 2864
rect 2883 2860 2884 2864
rect 2878 2859 2884 2860
rect 3030 2864 3036 2865
rect 3030 2860 3031 2864
rect 3035 2860 3036 2864
rect 3030 2859 3036 2860
rect 3190 2864 3196 2865
rect 3190 2860 3191 2864
rect 3195 2860 3196 2864
rect 3190 2859 3196 2860
rect 3358 2864 3364 2865
rect 3358 2860 3359 2864
rect 3363 2860 3364 2864
rect 3358 2859 3364 2860
rect 3502 2864 3508 2865
rect 3502 2860 3503 2864
rect 3507 2860 3508 2864
rect 3592 2862 3594 2881
rect 3502 2859 3508 2860
rect 3590 2861 3596 2862
rect 1870 2856 1876 2857
rect 3590 2857 3591 2861
rect 3595 2857 3596 2861
rect 3590 2856 3596 2857
rect 1870 2844 1876 2845
rect 1870 2840 1871 2844
rect 1875 2840 1876 2844
rect 1870 2839 1876 2840
rect 3590 2844 3596 2845
rect 3590 2840 3591 2844
rect 3595 2840 3596 2844
rect 3590 2839 3596 2840
rect 111 2830 115 2831
rect 111 2825 115 2826
rect 143 2830 147 2831
rect 143 2825 147 2826
rect 159 2830 163 2831
rect 159 2825 163 2826
rect 247 2830 251 2831
rect 247 2825 251 2826
rect 319 2830 323 2831
rect 319 2825 323 2826
rect 383 2830 387 2831
rect 383 2825 387 2826
rect 479 2830 483 2831
rect 479 2825 483 2826
rect 535 2830 539 2831
rect 535 2825 539 2826
rect 639 2830 643 2831
rect 639 2825 643 2826
rect 687 2830 691 2831
rect 687 2825 691 2826
rect 791 2830 795 2831
rect 791 2825 795 2826
rect 847 2830 851 2831
rect 847 2825 851 2826
rect 935 2830 939 2831
rect 935 2825 939 2826
rect 999 2830 1003 2831
rect 999 2825 1003 2826
rect 1063 2830 1067 2831
rect 1063 2825 1067 2826
rect 1143 2830 1147 2831
rect 1143 2825 1147 2826
rect 1183 2830 1187 2831
rect 1183 2825 1187 2826
rect 1279 2830 1283 2831
rect 1279 2825 1283 2826
rect 1295 2830 1299 2831
rect 1295 2825 1299 2826
rect 1399 2830 1403 2831
rect 1399 2825 1403 2826
rect 1407 2830 1411 2831
rect 1407 2825 1411 2826
rect 1495 2830 1499 2831
rect 1495 2825 1499 2826
rect 1527 2830 1531 2831
rect 1527 2825 1531 2826
rect 1599 2830 1603 2831
rect 1599 2825 1603 2826
rect 1647 2830 1651 2831
rect 1647 2825 1651 2826
rect 1703 2830 1707 2831
rect 1703 2825 1707 2826
rect 1751 2830 1755 2831
rect 1751 2825 1755 2826
rect 1831 2830 1835 2831
rect 1831 2825 1835 2826
rect 112 2797 114 2825
rect 144 2815 146 2825
rect 248 2815 250 2825
rect 384 2815 386 2825
rect 536 2815 538 2825
rect 688 2815 690 2825
rect 848 2815 850 2825
rect 1000 2815 1002 2825
rect 1144 2815 1146 2825
rect 1280 2815 1282 2825
rect 1408 2815 1410 2825
rect 1528 2815 1530 2825
rect 1648 2815 1650 2825
rect 1752 2815 1754 2825
rect 142 2814 148 2815
rect 142 2810 143 2814
rect 147 2810 148 2814
rect 142 2809 148 2810
rect 246 2814 252 2815
rect 246 2810 247 2814
rect 251 2810 252 2814
rect 246 2809 252 2810
rect 382 2814 388 2815
rect 382 2810 383 2814
rect 387 2810 388 2814
rect 382 2809 388 2810
rect 534 2814 540 2815
rect 534 2810 535 2814
rect 539 2810 540 2814
rect 534 2809 540 2810
rect 686 2814 692 2815
rect 686 2810 687 2814
rect 691 2810 692 2814
rect 686 2809 692 2810
rect 846 2814 852 2815
rect 846 2810 847 2814
rect 851 2810 852 2814
rect 846 2809 852 2810
rect 998 2814 1004 2815
rect 998 2810 999 2814
rect 1003 2810 1004 2814
rect 998 2809 1004 2810
rect 1142 2814 1148 2815
rect 1142 2810 1143 2814
rect 1147 2810 1148 2814
rect 1142 2809 1148 2810
rect 1278 2814 1284 2815
rect 1278 2810 1279 2814
rect 1283 2810 1284 2814
rect 1278 2809 1284 2810
rect 1406 2814 1412 2815
rect 1406 2810 1407 2814
rect 1411 2810 1412 2814
rect 1406 2809 1412 2810
rect 1526 2814 1532 2815
rect 1526 2810 1527 2814
rect 1531 2810 1532 2814
rect 1526 2809 1532 2810
rect 1646 2814 1652 2815
rect 1646 2810 1647 2814
rect 1651 2810 1652 2814
rect 1646 2809 1652 2810
rect 1750 2814 1756 2815
rect 1750 2810 1751 2814
rect 1755 2810 1756 2814
rect 1750 2809 1756 2810
rect 1832 2797 1834 2825
rect 1872 2799 1874 2839
rect 2054 2826 2060 2827
rect 2054 2822 2055 2826
rect 2059 2822 2060 2826
rect 2054 2821 2060 2822
rect 2142 2826 2148 2827
rect 2142 2822 2143 2826
rect 2147 2822 2148 2826
rect 2142 2821 2148 2822
rect 2246 2826 2252 2827
rect 2246 2822 2247 2826
rect 2251 2822 2252 2826
rect 2246 2821 2252 2822
rect 2350 2826 2356 2827
rect 2350 2822 2351 2826
rect 2355 2822 2356 2826
rect 2350 2821 2356 2822
rect 2470 2826 2476 2827
rect 2470 2822 2471 2826
rect 2475 2822 2476 2826
rect 2470 2821 2476 2822
rect 2598 2826 2604 2827
rect 2598 2822 2599 2826
rect 2603 2822 2604 2826
rect 2598 2821 2604 2822
rect 2734 2826 2740 2827
rect 2734 2822 2735 2826
rect 2739 2822 2740 2826
rect 2734 2821 2740 2822
rect 2886 2826 2892 2827
rect 2886 2822 2887 2826
rect 2891 2822 2892 2826
rect 2886 2821 2892 2822
rect 3038 2826 3044 2827
rect 3038 2822 3039 2826
rect 3043 2822 3044 2826
rect 3038 2821 3044 2822
rect 3198 2826 3204 2827
rect 3198 2822 3199 2826
rect 3203 2822 3204 2826
rect 3198 2821 3204 2822
rect 3366 2826 3372 2827
rect 3366 2822 3367 2826
rect 3371 2822 3372 2826
rect 3366 2821 3372 2822
rect 3510 2826 3516 2827
rect 3510 2822 3511 2826
rect 3515 2822 3516 2826
rect 3510 2821 3516 2822
rect 2056 2799 2058 2821
rect 2144 2799 2146 2821
rect 2248 2799 2250 2821
rect 2352 2799 2354 2821
rect 2472 2799 2474 2821
rect 2600 2799 2602 2821
rect 2736 2799 2738 2821
rect 2888 2799 2890 2821
rect 3040 2799 3042 2821
rect 3200 2799 3202 2821
rect 3368 2799 3370 2821
rect 3512 2799 3514 2821
rect 3592 2799 3594 2839
rect 1871 2798 1875 2799
rect 110 2796 116 2797
rect 110 2792 111 2796
rect 115 2792 116 2796
rect 110 2791 116 2792
rect 1830 2796 1836 2797
rect 1830 2792 1831 2796
rect 1835 2792 1836 2796
rect 1871 2793 1875 2794
rect 1903 2798 1907 2799
rect 1903 2793 1907 2794
rect 2015 2798 2019 2799
rect 2015 2793 2019 2794
rect 2055 2798 2059 2799
rect 2055 2793 2059 2794
rect 2143 2798 2147 2799
rect 2143 2793 2147 2794
rect 2167 2798 2171 2799
rect 2167 2793 2171 2794
rect 2247 2798 2251 2799
rect 2247 2793 2251 2794
rect 2327 2798 2331 2799
rect 2327 2793 2331 2794
rect 2351 2798 2355 2799
rect 2351 2793 2355 2794
rect 2471 2798 2475 2799
rect 2471 2793 2475 2794
rect 2487 2798 2491 2799
rect 2487 2793 2491 2794
rect 2599 2798 2603 2799
rect 2599 2793 2603 2794
rect 2639 2798 2643 2799
rect 2639 2793 2643 2794
rect 2735 2798 2739 2799
rect 2735 2793 2739 2794
rect 2791 2798 2795 2799
rect 2791 2793 2795 2794
rect 2887 2798 2891 2799
rect 2887 2793 2891 2794
rect 2943 2798 2947 2799
rect 2943 2793 2947 2794
rect 3039 2798 3043 2799
rect 3039 2793 3043 2794
rect 3087 2798 3091 2799
rect 3087 2793 3091 2794
rect 3199 2798 3203 2799
rect 3199 2793 3203 2794
rect 3231 2798 3235 2799
rect 3231 2793 3235 2794
rect 3367 2798 3371 2799
rect 3367 2793 3371 2794
rect 3383 2798 3387 2799
rect 3383 2793 3387 2794
rect 3511 2798 3515 2799
rect 3511 2793 3515 2794
rect 3591 2798 3595 2799
rect 3591 2793 3595 2794
rect 1830 2791 1836 2792
rect 110 2779 116 2780
rect 110 2775 111 2779
rect 115 2775 116 2779
rect 1830 2779 1836 2780
rect 110 2774 116 2775
rect 134 2776 140 2777
rect 112 2751 114 2774
rect 134 2772 135 2776
rect 139 2772 140 2776
rect 134 2771 140 2772
rect 238 2776 244 2777
rect 238 2772 239 2776
rect 243 2772 244 2776
rect 238 2771 244 2772
rect 374 2776 380 2777
rect 374 2772 375 2776
rect 379 2772 380 2776
rect 374 2771 380 2772
rect 526 2776 532 2777
rect 526 2772 527 2776
rect 531 2772 532 2776
rect 526 2771 532 2772
rect 678 2776 684 2777
rect 678 2772 679 2776
rect 683 2772 684 2776
rect 678 2771 684 2772
rect 838 2776 844 2777
rect 838 2772 839 2776
rect 843 2772 844 2776
rect 838 2771 844 2772
rect 990 2776 996 2777
rect 990 2772 991 2776
rect 995 2772 996 2776
rect 990 2771 996 2772
rect 1134 2776 1140 2777
rect 1134 2772 1135 2776
rect 1139 2772 1140 2776
rect 1134 2771 1140 2772
rect 1270 2776 1276 2777
rect 1270 2772 1271 2776
rect 1275 2772 1276 2776
rect 1270 2771 1276 2772
rect 1398 2776 1404 2777
rect 1398 2772 1399 2776
rect 1403 2772 1404 2776
rect 1398 2771 1404 2772
rect 1518 2776 1524 2777
rect 1518 2772 1519 2776
rect 1523 2772 1524 2776
rect 1518 2771 1524 2772
rect 1638 2776 1644 2777
rect 1638 2772 1639 2776
rect 1643 2772 1644 2776
rect 1638 2771 1644 2772
rect 1742 2776 1748 2777
rect 1742 2772 1743 2776
rect 1747 2772 1748 2776
rect 1830 2775 1831 2779
rect 1835 2775 1836 2779
rect 1830 2774 1836 2775
rect 1742 2771 1748 2772
rect 136 2751 138 2771
rect 240 2751 242 2771
rect 376 2751 378 2771
rect 528 2751 530 2771
rect 680 2751 682 2771
rect 840 2751 842 2771
rect 992 2751 994 2771
rect 1136 2751 1138 2771
rect 1272 2751 1274 2771
rect 1400 2751 1402 2771
rect 1520 2751 1522 2771
rect 1640 2751 1642 2771
rect 1744 2751 1746 2771
rect 1832 2751 1834 2774
rect 1872 2765 1874 2793
rect 1904 2783 1906 2793
rect 2016 2783 2018 2793
rect 2168 2783 2170 2793
rect 2328 2783 2330 2793
rect 2488 2783 2490 2793
rect 2640 2783 2642 2793
rect 2792 2783 2794 2793
rect 2944 2783 2946 2793
rect 3088 2783 3090 2793
rect 3232 2783 3234 2793
rect 3384 2783 3386 2793
rect 3512 2783 3514 2793
rect 1902 2782 1908 2783
rect 1902 2778 1903 2782
rect 1907 2778 1908 2782
rect 1902 2777 1908 2778
rect 2014 2782 2020 2783
rect 2014 2778 2015 2782
rect 2019 2778 2020 2782
rect 2014 2777 2020 2778
rect 2166 2782 2172 2783
rect 2166 2778 2167 2782
rect 2171 2778 2172 2782
rect 2166 2777 2172 2778
rect 2326 2782 2332 2783
rect 2326 2778 2327 2782
rect 2331 2778 2332 2782
rect 2326 2777 2332 2778
rect 2486 2782 2492 2783
rect 2486 2778 2487 2782
rect 2491 2778 2492 2782
rect 2486 2777 2492 2778
rect 2638 2782 2644 2783
rect 2638 2778 2639 2782
rect 2643 2778 2644 2782
rect 2638 2777 2644 2778
rect 2790 2782 2796 2783
rect 2790 2778 2791 2782
rect 2795 2778 2796 2782
rect 2790 2777 2796 2778
rect 2942 2782 2948 2783
rect 2942 2778 2943 2782
rect 2947 2778 2948 2782
rect 2942 2777 2948 2778
rect 3086 2782 3092 2783
rect 3086 2778 3087 2782
rect 3091 2778 3092 2782
rect 3086 2777 3092 2778
rect 3230 2782 3236 2783
rect 3230 2778 3231 2782
rect 3235 2778 3236 2782
rect 3230 2777 3236 2778
rect 3382 2782 3388 2783
rect 3382 2778 3383 2782
rect 3387 2778 3388 2782
rect 3382 2777 3388 2778
rect 3510 2782 3516 2783
rect 3510 2778 3511 2782
rect 3515 2778 3516 2782
rect 3510 2777 3516 2778
rect 3592 2765 3594 2793
rect 1870 2764 1876 2765
rect 1870 2760 1871 2764
rect 1875 2760 1876 2764
rect 1870 2759 1876 2760
rect 3590 2764 3596 2765
rect 3590 2760 3591 2764
rect 3595 2760 3596 2764
rect 3590 2759 3596 2760
rect 111 2750 115 2751
rect 111 2745 115 2746
rect 135 2750 139 2751
rect 135 2745 139 2746
rect 231 2750 235 2751
rect 231 2745 235 2746
rect 239 2750 243 2751
rect 239 2745 243 2746
rect 367 2750 371 2751
rect 367 2745 371 2746
rect 375 2750 379 2751
rect 375 2745 379 2746
rect 511 2750 515 2751
rect 511 2745 515 2746
rect 527 2750 531 2751
rect 527 2745 531 2746
rect 663 2750 667 2751
rect 663 2745 667 2746
rect 679 2750 683 2751
rect 679 2745 683 2746
rect 815 2750 819 2751
rect 815 2745 819 2746
rect 839 2750 843 2751
rect 839 2745 843 2746
rect 975 2750 979 2751
rect 975 2745 979 2746
rect 991 2750 995 2751
rect 991 2745 995 2746
rect 1135 2750 1139 2751
rect 1135 2745 1139 2746
rect 1271 2750 1275 2751
rect 1271 2745 1275 2746
rect 1287 2750 1291 2751
rect 1287 2745 1291 2746
rect 1399 2750 1403 2751
rect 1399 2745 1403 2746
rect 1447 2750 1451 2751
rect 1447 2745 1451 2746
rect 1519 2750 1523 2751
rect 1519 2745 1523 2746
rect 1607 2750 1611 2751
rect 1607 2745 1611 2746
rect 1639 2750 1643 2751
rect 1639 2745 1643 2746
rect 1743 2750 1747 2751
rect 1743 2745 1747 2746
rect 1831 2750 1835 2751
rect 1831 2745 1835 2746
rect 1870 2747 1876 2748
rect 112 2726 114 2745
rect 136 2729 138 2745
rect 232 2729 234 2745
rect 368 2729 370 2745
rect 512 2729 514 2745
rect 664 2729 666 2745
rect 816 2729 818 2745
rect 976 2729 978 2745
rect 1136 2729 1138 2745
rect 1288 2729 1290 2745
rect 1448 2729 1450 2745
rect 1608 2729 1610 2745
rect 1744 2729 1746 2745
rect 134 2728 140 2729
rect 110 2725 116 2726
rect 110 2721 111 2725
rect 115 2721 116 2725
rect 134 2724 135 2728
rect 139 2724 140 2728
rect 134 2723 140 2724
rect 230 2728 236 2729
rect 230 2724 231 2728
rect 235 2724 236 2728
rect 230 2723 236 2724
rect 366 2728 372 2729
rect 366 2724 367 2728
rect 371 2724 372 2728
rect 366 2723 372 2724
rect 510 2728 516 2729
rect 510 2724 511 2728
rect 515 2724 516 2728
rect 510 2723 516 2724
rect 662 2728 668 2729
rect 662 2724 663 2728
rect 667 2724 668 2728
rect 662 2723 668 2724
rect 814 2728 820 2729
rect 814 2724 815 2728
rect 819 2724 820 2728
rect 814 2723 820 2724
rect 974 2728 980 2729
rect 974 2724 975 2728
rect 979 2724 980 2728
rect 974 2723 980 2724
rect 1134 2728 1140 2729
rect 1134 2724 1135 2728
rect 1139 2724 1140 2728
rect 1134 2723 1140 2724
rect 1286 2728 1292 2729
rect 1286 2724 1287 2728
rect 1291 2724 1292 2728
rect 1286 2723 1292 2724
rect 1446 2728 1452 2729
rect 1446 2724 1447 2728
rect 1451 2724 1452 2728
rect 1446 2723 1452 2724
rect 1606 2728 1612 2729
rect 1606 2724 1607 2728
rect 1611 2724 1612 2728
rect 1606 2723 1612 2724
rect 1742 2728 1748 2729
rect 1742 2724 1743 2728
rect 1747 2724 1748 2728
rect 1832 2726 1834 2745
rect 1870 2743 1871 2747
rect 1875 2743 1876 2747
rect 3590 2747 3596 2748
rect 1870 2742 1876 2743
rect 1894 2744 1900 2745
rect 1742 2723 1748 2724
rect 1830 2725 1836 2726
rect 110 2720 116 2721
rect 1830 2721 1831 2725
rect 1835 2721 1836 2725
rect 1872 2723 1874 2742
rect 1894 2740 1895 2744
rect 1899 2740 1900 2744
rect 1894 2739 1900 2740
rect 2006 2744 2012 2745
rect 2006 2740 2007 2744
rect 2011 2740 2012 2744
rect 2006 2739 2012 2740
rect 2158 2744 2164 2745
rect 2158 2740 2159 2744
rect 2163 2740 2164 2744
rect 2158 2739 2164 2740
rect 2318 2744 2324 2745
rect 2318 2740 2319 2744
rect 2323 2740 2324 2744
rect 2318 2739 2324 2740
rect 2478 2744 2484 2745
rect 2478 2740 2479 2744
rect 2483 2740 2484 2744
rect 2478 2739 2484 2740
rect 2630 2744 2636 2745
rect 2630 2740 2631 2744
rect 2635 2740 2636 2744
rect 2630 2739 2636 2740
rect 2782 2744 2788 2745
rect 2782 2740 2783 2744
rect 2787 2740 2788 2744
rect 2782 2739 2788 2740
rect 2934 2744 2940 2745
rect 2934 2740 2935 2744
rect 2939 2740 2940 2744
rect 2934 2739 2940 2740
rect 3078 2744 3084 2745
rect 3078 2740 3079 2744
rect 3083 2740 3084 2744
rect 3078 2739 3084 2740
rect 3222 2744 3228 2745
rect 3222 2740 3223 2744
rect 3227 2740 3228 2744
rect 3222 2739 3228 2740
rect 3374 2744 3380 2745
rect 3374 2740 3375 2744
rect 3379 2740 3380 2744
rect 3374 2739 3380 2740
rect 3502 2744 3508 2745
rect 3502 2740 3503 2744
rect 3507 2740 3508 2744
rect 3590 2743 3591 2747
rect 3595 2743 3596 2747
rect 3590 2742 3596 2743
rect 3502 2739 3508 2740
rect 1896 2723 1898 2739
rect 2008 2723 2010 2739
rect 2160 2723 2162 2739
rect 2320 2723 2322 2739
rect 2480 2723 2482 2739
rect 2632 2723 2634 2739
rect 2784 2723 2786 2739
rect 2936 2723 2938 2739
rect 3080 2723 3082 2739
rect 3224 2723 3226 2739
rect 3376 2723 3378 2739
rect 3504 2723 3506 2739
rect 3592 2723 3594 2742
rect 1830 2720 1836 2721
rect 1871 2722 1875 2723
rect 1871 2717 1875 2718
rect 1895 2722 1899 2723
rect 1895 2717 1899 2718
rect 2007 2722 2011 2723
rect 2007 2717 2011 2718
rect 2103 2722 2107 2723
rect 2103 2717 2107 2718
rect 2159 2722 2163 2723
rect 2159 2717 2163 2718
rect 2319 2722 2323 2723
rect 2319 2717 2323 2718
rect 2327 2722 2331 2723
rect 2327 2717 2331 2718
rect 2479 2722 2483 2723
rect 2479 2717 2483 2718
rect 2535 2722 2539 2723
rect 2535 2717 2539 2718
rect 2631 2722 2635 2723
rect 2631 2717 2635 2718
rect 2735 2722 2739 2723
rect 2735 2717 2739 2718
rect 2783 2722 2787 2723
rect 2783 2717 2787 2718
rect 2911 2722 2915 2723
rect 2911 2717 2915 2718
rect 2935 2722 2939 2723
rect 2935 2717 2939 2718
rect 3071 2722 3075 2723
rect 3071 2717 3075 2718
rect 3079 2722 3083 2723
rect 3079 2717 3083 2718
rect 3223 2722 3227 2723
rect 3223 2717 3227 2718
rect 3375 2722 3379 2723
rect 3375 2717 3379 2718
rect 3503 2722 3507 2723
rect 3503 2717 3507 2718
rect 3591 2722 3595 2723
rect 3591 2717 3595 2718
rect 110 2708 116 2709
rect 110 2704 111 2708
rect 115 2704 116 2708
rect 110 2703 116 2704
rect 1830 2708 1836 2709
rect 1830 2704 1831 2708
rect 1835 2704 1836 2708
rect 1830 2703 1836 2704
rect 112 2667 114 2703
rect 142 2690 148 2691
rect 142 2686 143 2690
rect 147 2686 148 2690
rect 142 2685 148 2686
rect 238 2690 244 2691
rect 238 2686 239 2690
rect 243 2686 244 2690
rect 238 2685 244 2686
rect 374 2690 380 2691
rect 374 2686 375 2690
rect 379 2686 380 2690
rect 374 2685 380 2686
rect 518 2690 524 2691
rect 518 2686 519 2690
rect 523 2686 524 2690
rect 518 2685 524 2686
rect 670 2690 676 2691
rect 670 2686 671 2690
rect 675 2686 676 2690
rect 670 2685 676 2686
rect 822 2690 828 2691
rect 822 2686 823 2690
rect 827 2686 828 2690
rect 822 2685 828 2686
rect 982 2690 988 2691
rect 982 2686 983 2690
rect 987 2686 988 2690
rect 982 2685 988 2686
rect 1142 2690 1148 2691
rect 1142 2686 1143 2690
rect 1147 2686 1148 2690
rect 1142 2685 1148 2686
rect 1294 2690 1300 2691
rect 1294 2686 1295 2690
rect 1299 2686 1300 2690
rect 1294 2685 1300 2686
rect 1454 2690 1460 2691
rect 1454 2686 1455 2690
rect 1459 2686 1460 2690
rect 1454 2685 1460 2686
rect 1614 2690 1620 2691
rect 1614 2686 1615 2690
rect 1619 2686 1620 2690
rect 1614 2685 1620 2686
rect 1750 2690 1756 2691
rect 1750 2686 1751 2690
rect 1755 2686 1756 2690
rect 1750 2685 1756 2686
rect 144 2667 146 2685
rect 240 2667 242 2685
rect 376 2667 378 2685
rect 520 2667 522 2685
rect 672 2667 674 2685
rect 824 2667 826 2685
rect 984 2667 986 2685
rect 1144 2667 1146 2685
rect 1296 2667 1298 2685
rect 1456 2667 1458 2685
rect 1616 2667 1618 2685
rect 1752 2667 1754 2685
rect 1832 2667 1834 2703
rect 1872 2698 1874 2717
rect 1896 2701 1898 2717
rect 2104 2701 2106 2717
rect 2328 2701 2330 2717
rect 2536 2701 2538 2717
rect 2736 2701 2738 2717
rect 2912 2701 2914 2717
rect 3072 2701 3074 2717
rect 3224 2701 3226 2717
rect 3376 2701 3378 2717
rect 3504 2701 3506 2717
rect 1894 2700 1900 2701
rect 1870 2697 1876 2698
rect 1870 2693 1871 2697
rect 1875 2693 1876 2697
rect 1894 2696 1895 2700
rect 1899 2696 1900 2700
rect 1894 2695 1900 2696
rect 2102 2700 2108 2701
rect 2102 2696 2103 2700
rect 2107 2696 2108 2700
rect 2102 2695 2108 2696
rect 2326 2700 2332 2701
rect 2326 2696 2327 2700
rect 2331 2696 2332 2700
rect 2326 2695 2332 2696
rect 2534 2700 2540 2701
rect 2534 2696 2535 2700
rect 2539 2696 2540 2700
rect 2534 2695 2540 2696
rect 2734 2700 2740 2701
rect 2734 2696 2735 2700
rect 2739 2696 2740 2700
rect 2734 2695 2740 2696
rect 2910 2700 2916 2701
rect 2910 2696 2911 2700
rect 2915 2696 2916 2700
rect 2910 2695 2916 2696
rect 3070 2700 3076 2701
rect 3070 2696 3071 2700
rect 3075 2696 3076 2700
rect 3070 2695 3076 2696
rect 3222 2700 3228 2701
rect 3222 2696 3223 2700
rect 3227 2696 3228 2700
rect 3222 2695 3228 2696
rect 3374 2700 3380 2701
rect 3374 2696 3375 2700
rect 3379 2696 3380 2700
rect 3374 2695 3380 2696
rect 3502 2700 3508 2701
rect 3502 2696 3503 2700
rect 3507 2696 3508 2700
rect 3592 2698 3594 2717
rect 3502 2695 3508 2696
rect 3590 2697 3596 2698
rect 1870 2692 1876 2693
rect 3590 2693 3591 2697
rect 3595 2693 3596 2697
rect 3590 2692 3596 2693
rect 1870 2680 1876 2681
rect 1870 2676 1871 2680
rect 1875 2676 1876 2680
rect 1870 2675 1876 2676
rect 3590 2680 3596 2681
rect 3590 2676 3591 2680
rect 3595 2676 3596 2680
rect 3590 2675 3596 2676
rect 111 2666 115 2667
rect 111 2661 115 2662
rect 143 2666 147 2667
rect 143 2661 147 2662
rect 239 2666 243 2667
rect 239 2661 243 2662
rect 279 2666 283 2667
rect 279 2661 283 2662
rect 375 2666 379 2667
rect 375 2661 379 2662
rect 447 2666 451 2667
rect 447 2661 451 2662
rect 519 2666 523 2667
rect 519 2661 523 2662
rect 623 2666 627 2667
rect 623 2661 627 2662
rect 671 2666 675 2667
rect 671 2661 675 2662
rect 791 2666 795 2667
rect 791 2661 795 2662
rect 823 2666 827 2667
rect 823 2661 827 2662
rect 951 2666 955 2667
rect 951 2661 955 2662
rect 983 2666 987 2667
rect 983 2661 987 2662
rect 1103 2666 1107 2667
rect 1103 2661 1107 2662
rect 1143 2666 1147 2667
rect 1143 2661 1147 2662
rect 1247 2666 1251 2667
rect 1247 2661 1251 2662
rect 1295 2666 1299 2667
rect 1295 2661 1299 2662
rect 1399 2666 1403 2667
rect 1399 2661 1403 2662
rect 1455 2666 1459 2667
rect 1455 2661 1459 2662
rect 1551 2666 1555 2667
rect 1551 2661 1555 2662
rect 1615 2666 1619 2667
rect 1615 2661 1619 2662
rect 1751 2666 1755 2667
rect 1751 2661 1755 2662
rect 1831 2666 1835 2667
rect 1831 2661 1835 2662
rect 112 2633 114 2661
rect 144 2651 146 2661
rect 280 2651 282 2661
rect 448 2651 450 2661
rect 624 2651 626 2661
rect 792 2651 794 2661
rect 952 2651 954 2661
rect 1104 2651 1106 2661
rect 1248 2651 1250 2661
rect 1400 2651 1402 2661
rect 1552 2651 1554 2661
rect 142 2650 148 2651
rect 142 2646 143 2650
rect 147 2646 148 2650
rect 142 2645 148 2646
rect 278 2650 284 2651
rect 278 2646 279 2650
rect 283 2646 284 2650
rect 278 2645 284 2646
rect 446 2650 452 2651
rect 446 2646 447 2650
rect 451 2646 452 2650
rect 446 2645 452 2646
rect 622 2650 628 2651
rect 622 2646 623 2650
rect 627 2646 628 2650
rect 622 2645 628 2646
rect 790 2650 796 2651
rect 790 2646 791 2650
rect 795 2646 796 2650
rect 790 2645 796 2646
rect 950 2650 956 2651
rect 950 2646 951 2650
rect 955 2646 956 2650
rect 950 2645 956 2646
rect 1102 2650 1108 2651
rect 1102 2646 1103 2650
rect 1107 2646 1108 2650
rect 1102 2645 1108 2646
rect 1246 2650 1252 2651
rect 1246 2646 1247 2650
rect 1251 2646 1252 2650
rect 1246 2645 1252 2646
rect 1398 2650 1404 2651
rect 1398 2646 1399 2650
rect 1403 2646 1404 2650
rect 1398 2645 1404 2646
rect 1550 2650 1556 2651
rect 1550 2646 1551 2650
rect 1555 2646 1556 2650
rect 1550 2645 1556 2646
rect 1832 2633 1834 2661
rect 1872 2639 1874 2675
rect 1902 2662 1908 2663
rect 1902 2658 1903 2662
rect 1907 2658 1908 2662
rect 1902 2657 1908 2658
rect 2110 2662 2116 2663
rect 2110 2658 2111 2662
rect 2115 2658 2116 2662
rect 2110 2657 2116 2658
rect 2334 2662 2340 2663
rect 2334 2658 2335 2662
rect 2339 2658 2340 2662
rect 2334 2657 2340 2658
rect 2542 2662 2548 2663
rect 2542 2658 2543 2662
rect 2547 2658 2548 2662
rect 2542 2657 2548 2658
rect 2742 2662 2748 2663
rect 2742 2658 2743 2662
rect 2747 2658 2748 2662
rect 2742 2657 2748 2658
rect 2918 2662 2924 2663
rect 2918 2658 2919 2662
rect 2923 2658 2924 2662
rect 2918 2657 2924 2658
rect 3078 2662 3084 2663
rect 3078 2658 3079 2662
rect 3083 2658 3084 2662
rect 3078 2657 3084 2658
rect 3230 2662 3236 2663
rect 3230 2658 3231 2662
rect 3235 2658 3236 2662
rect 3230 2657 3236 2658
rect 3382 2662 3388 2663
rect 3382 2658 3383 2662
rect 3387 2658 3388 2662
rect 3382 2657 3388 2658
rect 3510 2662 3516 2663
rect 3510 2658 3511 2662
rect 3515 2658 3516 2662
rect 3510 2657 3516 2658
rect 1904 2639 1906 2657
rect 2112 2639 2114 2657
rect 2336 2639 2338 2657
rect 2544 2639 2546 2657
rect 2744 2639 2746 2657
rect 2920 2639 2922 2657
rect 3080 2639 3082 2657
rect 3232 2639 3234 2657
rect 3384 2639 3386 2657
rect 3512 2639 3514 2657
rect 3592 2639 3594 2675
rect 1871 2638 1875 2639
rect 1871 2633 1875 2634
rect 1903 2638 1907 2639
rect 1903 2633 1907 2634
rect 2055 2638 2059 2639
rect 2055 2633 2059 2634
rect 2111 2638 2115 2639
rect 2111 2633 2115 2634
rect 2263 2638 2267 2639
rect 2263 2633 2267 2634
rect 2335 2638 2339 2639
rect 2335 2633 2339 2634
rect 2495 2638 2499 2639
rect 2495 2633 2499 2634
rect 2543 2638 2547 2639
rect 2543 2633 2547 2634
rect 2743 2638 2747 2639
rect 2743 2633 2747 2634
rect 2751 2638 2755 2639
rect 2751 2633 2755 2634
rect 2919 2638 2923 2639
rect 2919 2633 2923 2634
rect 3015 2638 3019 2639
rect 3015 2633 3019 2634
rect 3079 2638 3083 2639
rect 3079 2633 3083 2634
rect 3231 2638 3235 2639
rect 3231 2633 3235 2634
rect 3287 2638 3291 2639
rect 3287 2633 3291 2634
rect 3383 2638 3387 2639
rect 3383 2633 3387 2634
rect 3511 2638 3515 2639
rect 3511 2633 3515 2634
rect 3591 2638 3595 2639
rect 3591 2633 3595 2634
rect 110 2632 116 2633
rect 110 2628 111 2632
rect 115 2628 116 2632
rect 110 2627 116 2628
rect 1830 2632 1836 2633
rect 1830 2628 1831 2632
rect 1835 2628 1836 2632
rect 1830 2627 1836 2628
rect 110 2615 116 2616
rect 110 2611 111 2615
rect 115 2611 116 2615
rect 1830 2615 1836 2616
rect 110 2610 116 2611
rect 134 2612 140 2613
rect 112 2587 114 2610
rect 134 2608 135 2612
rect 139 2608 140 2612
rect 134 2607 140 2608
rect 270 2612 276 2613
rect 270 2608 271 2612
rect 275 2608 276 2612
rect 270 2607 276 2608
rect 438 2612 444 2613
rect 438 2608 439 2612
rect 443 2608 444 2612
rect 438 2607 444 2608
rect 614 2612 620 2613
rect 614 2608 615 2612
rect 619 2608 620 2612
rect 614 2607 620 2608
rect 782 2612 788 2613
rect 782 2608 783 2612
rect 787 2608 788 2612
rect 782 2607 788 2608
rect 942 2612 948 2613
rect 942 2608 943 2612
rect 947 2608 948 2612
rect 942 2607 948 2608
rect 1094 2612 1100 2613
rect 1094 2608 1095 2612
rect 1099 2608 1100 2612
rect 1094 2607 1100 2608
rect 1238 2612 1244 2613
rect 1238 2608 1239 2612
rect 1243 2608 1244 2612
rect 1238 2607 1244 2608
rect 1390 2612 1396 2613
rect 1390 2608 1391 2612
rect 1395 2608 1396 2612
rect 1390 2607 1396 2608
rect 1542 2612 1548 2613
rect 1542 2608 1543 2612
rect 1547 2608 1548 2612
rect 1830 2611 1831 2615
rect 1835 2611 1836 2615
rect 1830 2610 1836 2611
rect 1542 2607 1548 2608
rect 136 2587 138 2607
rect 272 2587 274 2607
rect 440 2587 442 2607
rect 616 2587 618 2607
rect 784 2587 786 2607
rect 944 2587 946 2607
rect 1096 2587 1098 2607
rect 1240 2587 1242 2607
rect 1392 2587 1394 2607
rect 1544 2587 1546 2607
rect 1832 2587 1834 2610
rect 1872 2605 1874 2633
rect 1904 2623 1906 2633
rect 2056 2623 2058 2633
rect 2264 2623 2266 2633
rect 2496 2623 2498 2633
rect 2752 2623 2754 2633
rect 3016 2623 3018 2633
rect 3288 2623 3290 2633
rect 1902 2622 1908 2623
rect 1902 2618 1903 2622
rect 1907 2618 1908 2622
rect 1902 2617 1908 2618
rect 2054 2622 2060 2623
rect 2054 2618 2055 2622
rect 2059 2618 2060 2622
rect 2054 2617 2060 2618
rect 2262 2622 2268 2623
rect 2262 2618 2263 2622
rect 2267 2618 2268 2622
rect 2262 2617 2268 2618
rect 2494 2622 2500 2623
rect 2494 2618 2495 2622
rect 2499 2618 2500 2622
rect 2494 2617 2500 2618
rect 2750 2622 2756 2623
rect 2750 2618 2751 2622
rect 2755 2618 2756 2622
rect 2750 2617 2756 2618
rect 3014 2622 3020 2623
rect 3014 2618 3015 2622
rect 3019 2618 3020 2622
rect 3014 2617 3020 2618
rect 3286 2622 3292 2623
rect 3286 2618 3287 2622
rect 3291 2618 3292 2622
rect 3286 2617 3292 2618
rect 3592 2605 3594 2633
rect 1870 2604 1876 2605
rect 1870 2600 1871 2604
rect 1875 2600 1876 2604
rect 1870 2599 1876 2600
rect 3590 2604 3596 2605
rect 3590 2600 3591 2604
rect 3595 2600 3596 2604
rect 3590 2599 3596 2600
rect 1870 2587 1876 2588
rect 111 2586 115 2587
rect 111 2581 115 2582
rect 135 2586 139 2587
rect 135 2581 139 2582
rect 223 2586 227 2587
rect 223 2581 227 2582
rect 271 2586 275 2587
rect 271 2581 275 2582
rect 367 2586 371 2587
rect 367 2581 371 2582
rect 439 2586 443 2587
rect 439 2581 443 2582
rect 527 2586 531 2587
rect 527 2581 531 2582
rect 615 2586 619 2587
rect 615 2581 619 2582
rect 703 2586 707 2587
rect 703 2581 707 2582
rect 783 2586 787 2587
rect 783 2581 787 2582
rect 879 2586 883 2587
rect 879 2581 883 2582
rect 943 2586 947 2587
rect 943 2581 947 2582
rect 1047 2586 1051 2587
rect 1047 2581 1051 2582
rect 1095 2586 1099 2587
rect 1095 2581 1099 2582
rect 1207 2586 1211 2587
rect 1207 2581 1211 2582
rect 1239 2586 1243 2587
rect 1239 2581 1243 2582
rect 1359 2586 1363 2587
rect 1359 2581 1363 2582
rect 1391 2586 1395 2587
rect 1391 2581 1395 2582
rect 1511 2586 1515 2587
rect 1511 2581 1515 2582
rect 1543 2586 1547 2587
rect 1543 2581 1547 2582
rect 1671 2586 1675 2587
rect 1671 2581 1675 2582
rect 1831 2586 1835 2587
rect 1870 2583 1871 2587
rect 1875 2583 1876 2587
rect 3590 2587 3596 2588
rect 1870 2582 1876 2583
rect 1894 2584 1900 2585
rect 1831 2581 1835 2582
rect 112 2562 114 2581
rect 136 2565 138 2581
rect 224 2565 226 2581
rect 368 2565 370 2581
rect 528 2565 530 2581
rect 704 2565 706 2581
rect 880 2565 882 2581
rect 1048 2565 1050 2581
rect 1208 2565 1210 2581
rect 1360 2565 1362 2581
rect 1512 2565 1514 2581
rect 1672 2565 1674 2581
rect 134 2564 140 2565
rect 110 2561 116 2562
rect 110 2557 111 2561
rect 115 2557 116 2561
rect 134 2560 135 2564
rect 139 2560 140 2564
rect 134 2559 140 2560
rect 222 2564 228 2565
rect 222 2560 223 2564
rect 227 2560 228 2564
rect 222 2559 228 2560
rect 366 2564 372 2565
rect 366 2560 367 2564
rect 371 2560 372 2564
rect 366 2559 372 2560
rect 526 2564 532 2565
rect 526 2560 527 2564
rect 531 2560 532 2564
rect 526 2559 532 2560
rect 702 2564 708 2565
rect 702 2560 703 2564
rect 707 2560 708 2564
rect 702 2559 708 2560
rect 878 2564 884 2565
rect 878 2560 879 2564
rect 883 2560 884 2564
rect 878 2559 884 2560
rect 1046 2564 1052 2565
rect 1046 2560 1047 2564
rect 1051 2560 1052 2564
rect 1046 2559 1052 2560
rect 1206 2564 1212 2565
rect 1206 2560 1207 2564
rect 1211 2560 1212 2564
rect 1206 2559 1212 2560
rect 1358 2564 1364 2565
rect 1358 2560 1359 2564
rect 1363 2560 1364 2564
rect 1358 2559 1364 2560
rect 1510 2564 1516 2565
rect 1510 2560 1511 2564
rect 1515 2560 1516 2564
rect 1510 2559 1516 2560
rect 1670 2564 1676 2565
rect 1670 2560 1671 2564
rect 1675 2560 1676 2564
rect 1832 2562 1834 2581
rect 1872 2563 1874 2582
rect 1894 2580 1895 2584
rect 1899 2580 1900 2584
rect 1894 2579 1900 2580
rect 2046 2584 2052 2585
rect 2046 2580 2047 2584
rect 2051 2580 2052 2584
rect 2046 2579 2052 2580
rect 2254 2584 2260 2585
rect 2254 2580 2255 2584
rect 2259 2580 2260 2584
rect 2254 2579 2260 2580
rect 2486 2584 2492 2585
rect 2486 2580 2487 2584
rect 2491 2580 2492 2584
rect 2486 2579 2492 2580
rect 2742 2584 2748 2585
rect 2742 2580 2743 2584
rect 2747 2580 2748 2584
rect 2742 2579 2748 2580
rect 3006 2584 3012 2585
rect 3006 2580 3007 2584
rect 3011 2580 3012 2584
rect 3006 2579 3012 2580
rect 3278 2584 3284 2585
rect 3278 2580 3279 2584
rect 3283 2580 3284 2584
rect 3590 2583 3591 2587
rect 3595 2583 3596 2587
rect 3590 2582 3596 2583
rect 3278 2579 3284 2580
rect 1896 2563 1898 2579
rect 2048 2563 2050 2579
rect 2256 2563 2258 2579
rect 2488 2563 2490 2579
rect 2744 2563 2746 2579
rect 3008 2563 3010 2579
rect 3280 2563 3282 2579
rect 3592 2563 3594 2582
rect 1871 2562 1875 2563
rect 1670 2559 1676 2560
rect 1830 2561 1836 2562
rect 110 2556 116 2557
rect 1830 2557 1831 2561
rect 1835 2557 1836 2561
rect 1871 2557 1875 2558
rect 1895 2562 1899 2563
rect 1895 2557 1899 2558
rect 2007 2562 2011 2563
rect 2007 2557 2011 2558
rect 2047 2562 2051 2563
rect 2047 2557 2051 2558
rect 2159 2562 2163 2563
rect 2159 2557 2163 2558
rect 2255 2562 2259 2563
rect 2255 2557 2259 2558
rect 2319 2562 2323 2563
rect 2319 2557 2323 2558
rect 2471 2562 2475 2563
rect 2471 2557 2475 2558
rect 2487 2562 2491 2563
rect 2487 2557 2491 2558
rect 2623 2562 2627 2563
rect 2623 2557 2627 2558
rect 2743 2562 2747 2563
rect 2743 2557 2747 2558
rect 2759 2562 2763 2563
rect 2759 2557 2763 2558
rect 2887 2562 2891 2563
rect 2887 2557 2891 2558
rect 3007 2562 3011 2563
rect 3007 2557 3011 2558
rect 3119 2562 3123 2563
rect 3119 2557 3123 2558
rect 3223 2562 3227 2563
rect 3223 2557 3227 2558
rect 3279 2562 3283 2563
rect 3279 2557 3283 2558
rect 3319 2562 3323 2563
rect 3319 2557 3323 2558
rect 3423 2562 3427 2563
rect 3423 2557 3427 2558
rect 3503 2562 3507 2563
rect 3503 2557 3507 2558
rect 3591 2562 3595 2563
rect 3591 2557 3595 2558
rect 1830 2556 1836 2557
rect 110 2544 116 2545
rect 110 2540 111 2544
rect 115 2540 116 2544
rect 110 2539 116 2540
rect 1830 2544 1836 2545
rect 1830 2540 1831 2544
rect 1835 2540 1836 2544
rect 1830 2539 1836 2540
rect 112 2507 114 2539
rect 142 2526 148 2527
rect 142 2522 143 2526
rect 147 2522 148 2526
rect 142 2521 148 2522
rect 230 2526 236 2527
rect 230 2522 231 2526
rect 235 2522 236 2526
rect 230 2521 236 2522
rect 374 2526 380 2527
rect 374 2522 375 2526
rect 379 2522 380 2526
rect 374 2521 380 2522
rect 534 2526 540 2527
rect 534 2522 535 2526
rect 539 2522 540 2526
rect 534 2521 540 2522
rect 710 2526 716 2527
rect 710 2522 711 2526
rect 715 2522 716 2526
rect 710 2521 716 2522
rect 886 2526 892 2527
rect 886 2522 887 2526
rect 891 2522 892 2526
rect 886 2521 892 2522
rect 1054 2526 1060 2527
rect 1054 2522 1055 2526
rect 1059 2522 1060 2526
rect 1054 2521 1060 2522
rect 1214 2526 1220 2527
rect 1214 2522 1215 2526
rect 1219 2522 1220 2526
rect 1214 2521 1220 2522
rect 1366 2526 1372 2527
rect 1366 2522 1367 2526
rect 1371 2522 1372 2526
rect 1366 2521 1372 2522
rect 1518 2526 1524 2527
rect 1518 2522 1519 2526
rect 1523 2522 1524 2526
rect 1518 2521 1524 2522
rect 1678 2526 1684 2527
rect 1678 2522 1679 2526
rect 1683 2522 1684 2526
rect 1678 2521 1684 2522
rect 144 2507 146 2521
rect 232 2507 234 2521
rect 376 2507 378 2521
rect 536 2507 538 2521
rect 712 2507 714 2521
rect 888 2507 890 2521
rect 1056 2507 1058 2521
rect 1216 2507 1218 2521
rect 1368 2507 1370 2521
rect 1520 2507 1522 2521
rect 1680 2507 1682 2521
rect 1832 2507 1834 2539
rect 1872 2538 1874 2557
rect 1896 2541 1898 2557
rect 2008 2541 2010 2557
rect 2160 2541 2162 2557
rect 2320 2541 2322 2557
rect 2472 2541 2474 2557
rect 2624 2541 2626 2557
rect 2760 2541 2762 2557
rect 2888 2541 2890 2557
rect 3008 2541 3010 2557
rect 3120 2541 3122 2557
rect 3224 2541 3226 2557
rect 3320 2541 3322 2557
rect 3424 2541 3426 2557
rect 3504 2541 3506 2557
rect 1894 2540 1900 2541
rect 1870 2537 1876 2538
rect 1870 2533 1871 2537
rect 1875 2533 1876 2537
rect 1894 2536 1895 2540
rect 1899 2536 1900 2540
rect 1894 2535 1900 2536
rect 2006 2540 2012 2541
rect 2006 2536 2007 2540
rect 2011 2536 2012 2540
rect 2006 2535 2012 2536
rect 2158 2540 2164 2541
rect 2158 2536 2159 2540
rect 2163 2536 2164 2540
rect 2158 2535 2164 2536
rect 2318 2540 2324 2541
rect 2318 2536 2319 2540
rect 2323 2536 2324 2540
rect 2318 2535 2324 2536
rect 2470 2540 2476 2541
rect 2470 2536 2471 2540
rect 2475 2536 2476 2540
rect 2470 2535 2476 2536
rect 2622 2540 2628 2541
rect 2622 2536 2623 2540
rect 2627 2536 2628 2540
rect 2622 2535 2628 2536
rect 2758 2540 2764 2541
rect 2758 2536 2759 2540
rect 2763 2536 2764 2540
rect 2758 2535 2764 2536
rect 2886 2540 2892 2541
rect 2886 2536 2887 2540
rect 2891 2536 2892 2540
rect 2886 2535 2892 2536
rect 3006 2540 3012 2541
rect 3006 2536 3007 2540
rect 3011 2536 3012 2540
rect 3006 2535 3012 2536
rect 3118 2540 3124 2541
rect 3118 2536 3119 2540
rect 3123 2536 3124 2540
rect 3118 2535 3124 2536
rect 3222 2540 3228 2541
rect 3222 2536 3223 2540
rect 3227 2536 3228 2540
rect 3222 2535 3228 2536
rect 3318 2540 3324 2541
rect 3318 2536 3319 2540
rect 3323 2536 3324 2540
rect 3318 2535 3324 2536
rect 3422 2540 3428 2541
rect 3422 2536 3423 2540
rect 3427 2536 3428 2540
rect 3422 2535 3428 2536
rect 3502 2540 3508 2541
rect 3502 2536 3503 2540
rect 3507 2536 3508 2540
rect 3592 2538 3594 2557
rect 3502 2535 3508 2536
rect 3590 2537 3596 2538
rect 1870 2532 1876 2533
rect 3590 2533 3591 2537
rect 3595 2533 3596 2537
rect 3590 2532 3596 2533
rect 1870 2520 1876 2521
rect 1870 2516 1871 2520
rect 1875 2516 1876 2520
rect 1870 2515 1876 2516
rect 3590 2520 3596 2521
rect 3590 2516 3591 2520
rect 3595 2516 3596 2520
rect 3590 2515 3596 2516
rect 111 2506 115 2507
rect 111 2501 115 2502
rect 143 2506 147 2507
rect 143 2501 147 2502
rect 223 2506 227 2507
rect 223 2501 227 2502
rect 231 2506 235 2507
rect 231 2501 235 2502
rect 303 2506 307 2507
rect 303 2501 307 2502
rect 375 2506 379 2507
rect 375 2501 379 2502
rect 391 2506 395 2507
rect 391 2501 395 2502
rect 511 2506 515 2507
rect 511 2501 515 2502
rect 535 2506 539 2507
rect 535 2501 539 2502
rect 647 2506 651 2507
rect 647 2501 651 2502
rect 711 2506 715 2507
rect 711 2501 715 2502
rect 783 2506 787 2507
rect 783 2501 787 2502
rect 887 2506 891 2507
rect 887 2501 891 2502
rect 927 2506 931 2507
rect 927 2501 931 2502
rect 1055 2506 1059 2507
rect 1055 2501 1059 2502
rect 1063 2506 1067 2507
rect 1063 2501 1067 2502
rect 1191 2506 1195 2507
rect 1191 2501 1195 2502
rect 1215 2506 1219 2507
rect 1215 2501 1219 2502
rect 1311 2506 1315 2507
rect 1311 2501 1315 2502
rect 1367 2506 1371 2507
rect 1367 2501 1371 2502
rect 1431 2506 1435 2507
rect 1431 2501 1435 2502
rect 1519 2506 1523 2507
rect 1519 2501 1523 2502
rect 1551 2506 1555 2507
rect 1551 2501 1555 2502
rect 1671 2506 1675 2507
rect 1671 2501 1675 2502
rect 1679 2506 1683 2507
rect 1679 2501 1683 2502
rect 1831 2506 1835 2507
rect 1831 2501 1835 2502
rect 112 2473 114 2501
rect 144 2491 146 2501
rect 224 2491 226 2501
rect 304 2491 306 2501
rect 392 2491 394 2501
rect 512 2491 514 2501
rect 648 2491 650 2501
rect 784 2491 786 2501
rect 928 2491 930 2501
rect 1064 2491 1066 2501
rect 1192 2491 1194 2501
rect 1312 2491 1314 2501
rect 1432 2491 1434 2501
rect 1552 2491 1554 2501
rect 1672 2491 1674 2501
rect 142 2490 148 2491
rect 142 2486 143 2490
rect 147 2486 148 2490
rect 142 2485 148 2486
rect 222 2490 228 2491
rect 222 2486 223 2490
rect 227 2486 228 2490
rect 222 2485 228 2486
rect 302 2490 308 2491
rect 302 2486 303 2490
rect 307 2486 308 2490
rect 302 2485 308 2486
rect 390 2490 396 2491
rect 390 2486 391 2490
rect 395 2486 396 2490
rect 390 2485 396 2486
rect 510 2490 516 2491
rect 510 2486 511 2490
rect 515 2486 516 2490
rect 510 2485 516 2486
rect 646 2490 652 2491
rect 646 2486 647 2490
rect 651 2486 652 2490
rect 646 2485 652 2486
rect 782 2490 788 2491
rect 782 2486 783 2490
rect 787 2486 788 2490
rect 782 2485 788 2486
rect 926 2490 932 2491
rect 926 2486 927 2490
rect 931 2486 932 2490
rect 926 2485 932 2486
rect 1062 2490 1068 2491
rect 1062 2486 1063 2490
rect 1067 2486 1068 2490
rect 1062 2485 1068 2486
rect 1190 2490 1196 2491
rect 1190 2486 1191 2490
rect 1195 2486 1196 2490
rect 1190 2485 1196 2486
rect 1310 2490 1316 2491
rect 1310 2486 1311 2490
rect 1315 2486 1316 2490
rect 1310 2485 1316 2486
rect 1430 2490 1436 2491
rect 1430 2486 1431 2490
rect 1435 2486 1436 2490
rect 1430 2485 1436 2486
rect 1550 2490 1556 2491
rect 1550 2486 1551 2490
rect 1555 2486 1556 2490
rect 1550 2485 1556 2486
rect 1670 2490 1676 2491
rect 1670 2486 1671 2490
rect 1675 2486 1676 2490
rect 1670 2485 1676 2486
rect 1832 2473 1834 2501
rect 1872 2479 1874 2515
rect 1902 2502 1908 2503
rect 1902 2498 1903 2502
rect 1907 2498 1908 2502
rect 1902 2497 1908 2498
rect 2014 2502 2020 2503
rect 2014 2498 2015 2502
rect 2019 2498 2020 2502
rect 2014 2497 2020 2498
rect 2166 2502 2172 2503
rect 2166 2498 2167 2502
rect 2171 2498 2172 2502
rect 2166 2497 2172 2498
rect 2326 2502 2332 2503
rect 2326 2498 2327 2502
rect 2331 2498 2332 2502
rect 2326 2497 2332 2498
rect 2478 2502 2484 2503
rect 2478 2498 2479 2502
rect 2483 2498 2484 2502
rect 2478 2497 2484 2498
rect 2630 2502 2636 2503
rect 2630 2498 2631 2502
rect 2635 2498 2636 2502
rect 2630 2497 2636 2498
rect 2766 2502 2772 2503
rect 2766 2498 2767 2502
rect 2771 2498 2772 2502
rect 2766 2497 2772 2498
rect 2894 2502 2900 2503
rect 2894 2498 2895 2502
rect 2899 2498 2900 2502
rect 2894 2497 2900 2498
rect 3014 2502 3020 2503
rect 3014 2498 3015 2502
rect 3019 2498 3020 2502
rect 3014 2497 3020 2498
rect 3126 2502 3132 2503
rect 3126 2498 3127 2502
rect 3131 2498 3132 2502
rect 3126 2497 3132 2498
rect 3230 2502 3236 2503
rect 3230 2498 3231 2502
rect 3235 2498 3236 2502
rect 3230 2497 3236 2498
rect 3326 2502 3332 2503
rect 3326 2498 3327 2502
rect 3331 2498 3332 2502
rect 3326 2497 3332 2498
rect 3430 2502 3436 2503
rect 3430 2498 3431 2502
rect 3435 2498 3436 2502
rect 3430 2497 3436 2498
rect 3510 2502 3516 2503
rect 3510 2498 3511 2502
rect 3515 2498 3516 2502
rect 3510 2497 3516 2498
rect 1904 2479 1906 2497
rect 2016 2479 2018 2497
rect 2168 2479 2170 2497
rect 2328 2479 2330 2497
rect 2480 2479 2482 2497
rect 2632 2479 2634 2497
rect 2768 2479 2770 2497
rect 2896 2479 2898 2497
rect 3016 2479 3018 2497
rect 3128 2479 3130 2497
rect 3232 2479 3234 2497
rect 3328 2479 3330 2497
rect 3432 2479 3434 2497
rect 3512 2479 3514 2497
rect 3592 2479 3594 2515
rect 1871 2478 1875 2479
rect 1871 2473 1875 2474
rect 1903 2478 1907 2479
rect 1903 2473 1907 2474
rect 1999 2478 2003 2479
rect 1999 2473 2003 2474
rect 2015 2478 2019 2479
rect 2015 2473 2019 2474
rect 2127 2478 2131 2479
rect 2127 2473 2131 2474
rect 2167 2478 2171 2479
rect 2167 2473 2171 2474
rect 2263 2478 2267 2479
rect 2263 2473 2267 2474
rect 2327 2478 2331 2479
rect 2327 2473 2331 2474
rect 2407 2478 2411 2479
rect 2407 2473 2411 2474
rect 2479 2478 2483 2479
rect 2479 2473 2483 2474
rect 2551 2478 2555 2479
rect 2551 2473 2555 2474
rect 2631 2478 2635 2479
rect 2631 2473 2635 2474
rect 2703 2478 2707 2479
rect 2703 2473 2707 2474
rect 2767 2478 2771 2479
rect 2767 2473 2771 2474
rect 2863 2478 2867 2479
rect 2863 2473 2867 2474
rect 2895 2478 2899 2479
rect 2895 2473 2899 2474
rect 3015 2478 3019 2479
rect 3015 2473 3019 2474
rect 3023 2478 3027 2479
rect 3023 2473 3027 2474
rect 3127 2478 3131 2479
rect 3127 2473 3131 2474
rect 3191 2478 3195 2479
rect 3191 2473 3195 2474
rect 3231 2478 3235 2479
rect 3231 2473 3235 2474
rect 3327 2478 3331 2479
rect 3327 2473 3331 2474
rect 3359 2478 3363 2479
rect 3359 2473 3363 2474
rect 3431 2478 3435 2479
rect 3431 2473 3435 2474
rect 3511 2478 3515 2479
rect 3511 2473 3515 2474
rect 3591 2478 3595 2479
rect 3591 2473 3595 2474
rect 110 2472 116 2473
rect 110 2468 111 2472
rect 115 2468 116 2472
rect 110 2467 116 2468
rect 1830 2472 1836 2473
rect 1830 2468 1831 2472
rect 1835 2468 1836 2472
rect 1830 2467 1836 2468
rect 110 2455 116 2456
rect 110 2451 111 2455
rect 115 2451 116 2455
rect 1830 2455 1836 2456
rect 110 2450 116 2451
rect 134 2452 140 2453
rect 112 2419 114 2450
rect 134 2448 135 2452
rect 139 2448 140 2452
rect 134 2447 140 2448
rect 214 2452 220 2453
rect 214 2448 215 2452
rect 219 2448 220 2452
rect 214 2447 220 2448
rect 294 2452 300 2453
rect 294 2448 295 2452
rect 299 2448 300 2452
rect 294 2447 300 2448
rect 382 2452 388 2453
rect 382 2448 383 2452
rect 387 2448 388 2452
rect 382 2447 388 2448
rect 502 2452 508 2453
rect 502 2448 503 2452
rect 507 2448 508 2452
rect 502 2447 508 2448
rect 638 2452 644 2453
rect 638 2448 639 2452
rect 643 2448 644 2452
rect 638 2447 644 2448
rect 774 2452 780 2453
rect 774 2448 775 2452
rect 779 2448 780 2452
rect 774 2447 780 2448
rect 918 2452 924 2453
rect 918 2448 919 2452
rect 923 2448 924 2452
rect 918 2447 924 2448
rect 1054 2452 1060 2453
rect 1054 2448 1055 2452
rect 1059 2448 1060 2452
rect 1054 2447 1060 2448
rect 1182 2452 1188 2453
rect 1182 2448 1183 2452
rect 1187 2448 1188 2452
rect 1182 2447 1188 2448
rect 1302 2452 1308 2453
rect 1302 2448 1303 2452
rect 1307 2448 1308 2452
rect 1302 2447 1308 2448
rect 1422 2452 1428 2453
rect 1422 2448 1423 2452
rect 1427 2448 1428 2452
rect 1422 2447 1428 2448
rect 1542 2452 1548 2453
rect 1542 2448 1543 2452
rect 1547 2448 1548 2452
rect 1542 2447 1548 2448
rect 1662 2452 1668 2453
rect 1662 2448 1663 2452
rect 1667 2448 1668 2452
rect 1830 2451 1831 2455
rect 1835 2451 1836 2455
rect 1830 2450 1836 2451
rect 1662 2447 1668 2448
rect 136 2419 138 2447
rect 216 2419 218 2447
rect 296 2419 298 2447
rect 384 2419 386 2447
rect 504 2419 506 2447
rect 640 2419 642 2447
rect 776 2419 778 2447
rect 920 2419 922 2447
rect 1056 2419 1058 2447
rect 1184 2419 1186 2447
rect 1304 2419 1306 2447
rect 1424 2419 1426 2447
rect 1544 2419 1546 2447
rect 1664 2419 1666 2447
rect 1832 2419 1834 2450
rect 1872 2445 1874 2473
rect 2000 2463 2002 2473
rect 2128 2463 2130 2473
rect 2264 2463 2266 2473
rect 2408 2463 2410 2473
rect 2552 2463 2554 2473
rect 2704 2463 2706 2473
rect 2864 2463 2866 2473
rect 3024 2463 3026 2473
rect 3192 2463 3194 2473
rect 3360 2463 3362 2473
rect 3512 2463 3514 2473
rect 1998 2462 2004 2463
rect 1998 2458 1999 2462
rect 2003 2458 2004 2462
rect 1998 2457 2004 2458
rect 2126 2462 2132 2463
rect 2126 2458 2127 2462
rect 2131 2458 2132 2462
rect 2126 2457 2132 2458
rect 2262 2462 2268 2463
rect 2262 2458 2263 2462
rect 2267 2458 2268 2462
rect 2262 2457 2268 2458
rect 2406 2462 2412 2463
rect 2406 2458 2407 2462
rect 2411 2458 2412 2462
rect 2406 2457 2412 2458
rect 2550 2462 2556 2463
rect 2550 2458 2551 2462
rect 2555 2458 2556 2462
rect 2550 2457 2556 2458
rect 2702 2462 2708 2463
rect 2702 2458 2703 2462
rect 2707 2458 2708 2462
rect 2702 2457 2708 2458
rect 2862 2462 2868 2463
rect 2862 2458 2863 2462
rect 2867 2458 2868 2462
rect 2862 2457 2868 2458
rect 3022 2462 3028 2463
rect 3022 2458 3023 2462
rect 3027 2458 3028 2462
rect 3022 2457 3028 2458
rect 3190 2462 3196 2463
rect 3190 2458 3191 2462
rect 3195 2458 3196 2462
rect 3190 2457 3196 2458
rect 3358 2462 3364 2463
rect 3358 2458 3359 2462
rect 3363 2458 3364 2462
rect 3358 2457 3364 2458
rect 3510 2462 3516 2463
rect 3510 2458 3511 2462
rect 3515 2458 3516 2462
rect 3510 2457 3516 2458
rect 3592 2445 3594 2473
rect 1870 2444 1876 2445
rect 1870 2440 1871 2444
rect 1875 2440 1876 2444
rect 1870 2439 1876 2440
rect 3590 2444 3596 2445
rect 3590 2440 3591 2444
rect 3595 2440 3596 2444
rect 3590 2439 3596 2440
rect 1870 2427 1876 2428
rect 1870 2423 1871 2427
rect 1875 2423 1876 2427
rect 3590 2427 3596 2428
rect 1870 2422 1876 2423
rect 1990 2424 1996 2425
rect 111 2418 115 2419
rect 111 2413 115 2414
rect 135 2418 139 2419
rect 135 2413 139 2414
rect 215 2418 219 2419
rect 215 2413 219 2414
rect 295 2418 299 2419
rect 295 2413 299 2414
rect 383 2418 387 2419
rect 383 2413 387 2414
rect 503 2418 507 2419
rect 503 2413 507 2414
rect 639 2418 643 2419
rect 639 2413 643 2414
rect 775 2418 779 2419
rect 775 2413 779 2414
rect 919 2418 923 2419
rect 919 2413 923 2414
rect 1055 2418 1059 2419
rect 1055 2413 1059 2414
rect 1063 2418 1067 2419
rect 1063 2413 1067 2414
rect 1143 2418 1147 2419
rect 1143 2413 1147 2414
rect 1183 2418 1187 2419
rect 1183 2413 1187 2414
rect 1223 2418 1227 2419
rect 1223 2413 1227 2414
rect 1303 2418 1307 2419
rect 1303 2413 1307 2414
rect 1383 2418 1387 2419
rect 1383 2413 1387 2414
rect 1423 2418 1427 2419
rect 1423 2413 1427 2414
rect 1463 2418 1467 2419
rect 1463 2413 1467 2414
rect 1543 2418 1547 2419
rect 1543 2413 1547 2414
rect 1663 2418 1667 2419
rect 1663 2413 1667 2414
rect 1831 2418 1835 2419
rect 1831 2413 1835 2414
rect 112 2394 114 2413
rect 1064 2397 1066 2413
rect 1144 2397 1146 2413
rect 1224 2397 1226 2413
rect 1304 2397 1306 2413
rect 1384 2397 1386 2413
rect 1464 2397 1466 2413
rect 1062 2396 1068 2397
rect 110 2393 116 2394
rect 110 2389 111 2393
rect 115 2389 116 2393
rect 1062 2392 1063 2396
rect 1067 2392 1068 2396
rect 1062 2391 1068 2392
rect 1142 2396 1148 2397
rect 1142 2392 1143 2396
rect 1147 2392 1148 2396
rect 1142 2391 1148 2392
rect 1222 2396 1228 2397
rect 1222 2392 1223 2396
rect 1227 2392 1228 2396
rect 1222 2391 1228 2392
rect 1302 2396 1308 2397
rect 1302 2392 1303 2396
rect 1307 2392 1308 2396
rect 1302 2391 1308 2392
rect 1382 2396 1388 2397
rect 1382 2392 1383 2396
rect 1387 2392 1388 2396
rect 1382 2391 1388 2392
rect 1462 2396 1468 2397
rect 1462 2392 1463 2396
rect 1467 2392 1468 2396
rect 1832 2394 1834 2413
rect 1872 2399 1874 2422
rect 1990 2420 1991 2424
rect 1995 2420 1996 2424
rect 1990 2419 1996 2420
rect 2118 2424 2124 2425
rect 2118 2420 2119 2424
rect 2123 2420 2124 2424
rect 2118 2419 2124 2420
rect 2254 2424 2260 2425
rect 2254 2420 2255 2424
rect 2259 2420 2260 2424
rect 2254 2419 2260 2420
rect 2398 2424 2404 2425
rect 2398 2420 2399 2424
rect 2403 2420 2404 2424
rect 2398 2419 2404 2420
rect 2542 2424 2548 2425
rect 2542 2420 2543 2424
rect 2547 2420 2548 2424
rect 2542 2419 2548 2420
rect 2694 2424 2700 2425
rect 2694 2420 2695 2424
rect 2699 2420 2700 2424
rect 2694 2419 2700 2420
rect 2854 2424 2860 2425
rect 2854 2420 2855 2424
rect 2859 2420 2860 2424
rect 2854 2419 2860 2420
rect 3014 2424 3020 2425
rect 3014 2420 3015 2424
rect 3019 2420 3020 2424
rect 3014 2419 3020 2420
rect 3182 2424 3188 2425
rect 3182 2420 3183 2424
rect 3187 2420 3188 2424
rect 3182 2419 3188 2420
rect 3350 2424 3356 2425
rect 3350 2420 3351 2424
rect 3355 2420 3356 2424
rect 3350 2419 3356 2420
rect 3502 2424 3508 2425
rect 3502 2420 3503 2424
rect 3507 2420 3508 2424
rect 3590 2423 3591 2427
rect 3595 2423 3596 2427
rect 3590 2422 3596 2423
rect 3502 2419 3508 2420
rect 1992 2399 1994 2419
rect 2120 2399 2122 2419
rect 2256 2399 2258 2419
rect 2400 2399 2402 2419
rect 2544 2399 2546 2419
rect 2696 2399 2698 2419
rect 2856 2399 2858 2419
rect 3016 2399 3018 2419
rect 3184 2399 3186 2419
rect 3352 2399 3354 2419
rect 3504 2399 3506 2419
rect 3592 2399 3594 2422
rect 1871 2398 1875 2399
rect 1462 2391 1468 2392
rect 1830 2393 1836 2394
rect 1871 2393 1875 2394
rect 1991 2398 1995 2399
rect 1991 2393 1995 2394
rect 2119 2398 2123 2399
rect 2119 2393 2123 2394
rect 2143 2398 2147 2399
rect 2143 2393 2147 2394
rect 2239 2398 2243 2399
rect 2239 2393 2243 2394
rect 2255 2398 2259 2399
rect 2255 2393 2259 2394
rect 2343 2398 2347 2399
rect 2343 2393 2347 2394
rect 2399 2398 2403 2399
rect 2399 2393 2403 2394
rect 2455 2398 2459 2399
rect 2455 2393 2459 2394
rect 2543 2398 2547 2399
rect 2543 2393 2547 2394
rect 2575 2398 2579 2399
rect 2575 2393 2579 2394
rect 2695 2398 2699 2399
rect 2695 2393 2699 2394
rect 2703 2398 2707 2399
rect 2703 2393 2707 2394
rect 2847 2398 2851 2399
rect 2847 2393 2851 2394
rect 2855 2398 2859 2399
rect 2855 2393 2859 2394
rect 3007 2398 3011 2399
rect 3007 2393 3011 2394
rect 3015 2398 3019 2399
rect 3015 2393 3019 2394
rect 3175 2398 3179 2399
rect 3175 2393 3179 2394
rect 3183 2398 3187 2399
rect 3183 2393 3187 2394
rect 3351 2398 3355 2399
rect 3351 2393 3355 2394
rect 3503 2398 3507 2399
rect 3503 2393 3507 2394
rect 3591 2398 3595 2399
rect 3591 2393 3595 2394
rect 110 2388 116 2389
rect 1830 2389 1831 2393
rect 1835 2389 1836 2393
rect 1830 2388 1836 2389
rect 110 2376 116 2377
rect 110 2372 111 2376
rect 115 2372 116 2376
rect 110 2371 116 2372
rect 1830 2376 1836 2377
rect 1830 2372 1831 2376
rect 1835 2372 1836 2376
rect 1872 2374 1874 2393
rect 2144 2377 2146 2393
rect 2240 2377 2242 2393
rect 2344 2377 2346 2393
rect 2456 2377 2458 2393
rect 2576 2377 2578 2393
rect 2704 2377 2706 2393
rect 2848 2377 2850 2393
rect 3008 2377 3010 2393
rect 3176 2377 3178 2393
rect 3352 2377 3354 2393
rect 3504 2377 3506 2393
rect 2142 2376 2148 2377
rect 1830 2371 1836 2372
rect 1870 2373 1876 2374
rect 112 2335 114 2371
rect 1070 2358 1076 2359
rect 1070 2354 1071 2358
rect 1075 2354 1076 2358
rect 1070 2353 1076 2354
rect 1150 2358 1156 2359
rect 1150 2354 1151 2358
rect 1155 2354 1156 2358
rect 1150 2353 1156 2354
rect 1230 2358 1236 2359
rect 1230 2354 1231 2358
rect 1235 2354 1236 2358
rect 1230 2353 1236 2354
rect 1310 2358 1316 2359
rect 1310 2354 1311 2358
rect 1315 2354 1316 2358
rect 1310 2353 1316 2354
rect 1390 2358 1396 2359
rect 1390 2354 1391 2358
rect 1395 2354 1396 2358
rect 1390 2353 1396 2354
rect 1470 2358 1476 2359
rect 1470 2354 1471 2358
rect 1475 2354 1476 2358
rect 1470 2353 1476 2354
rect 1072 2335 1074 2353
rect 1152 2335 1154 2353
rect 1232 2335 1234 2353
rect 1312 2335 1314 2353
rect 1392 2335 1394 2353
rect 1472 2335 1474 2353
rect 1832 2335 1834 2371
rect 1870 2369 1871 2373
rect 1875 2369 1876 2373
rect 2142 2372 2143 2376
rect 2147 2372 2148 2376
rect 2142 2371 2148 2372
rect 2238 2376 2244 2377
rect 2238 2372 2239 2376
rect 2243 2372 2244 2376
rect 2238 2371 2244 2372
rect 2342 2376 2348 2377
rect 2342 2372 2343 2376
rect 2347 2372 2348 2376
rect 2342 2371 2348 2372
rect 2454 2376 2460 2377
rect 2454 2372 2455 2376
rect 2459 2372 2460 2376
rect 2454 2371 2460 2372
rect 2574 2376 2580 2377
rect 2574 2372 2575 2376
rect 2579 2372 2580 2376
rect 2574 2371 2580 2372
rect 2702 2376 2708 2377
rect 2702 2372 2703 2376
rect 2707 2372 2708 2376
rect 2702 2371 2708 2372
rect 2846 2376 2852 2377
rect 2846 2372 2847 2376
rect 2851 2372 2852 2376
rect 2846 2371 2852 2372
rect 3006 2376 3012 2377
rect 3006 2372 3007 2376
rect 3011 2372 3012 2376
rect 3006 2371 3012 2372
rect 3174 2376 3180 2377
rect 3174 2372 3175 2376
rect 3179 2372 3180 2376
rect 3174 2371 3180 2372
rect 3350 2376 3356 2377
rect 3350 2372 3351 2376
rect 3355 2372 3356 2376
rect 3350 2371 3356 2372
rect 3502 2376 3508 2377
rect 3502 2372 3503 2376
rect 3507 2372 3508 2376
rect 3592 2374 3594 2393
rect 3502 2371 3508 2372
rect 3590 2373 3596 2374
rect 1870 2368 1876 2369
rect 3590 2369 3591 2373
rect 3595 2369 3596 2373
rect 3590 2368 3596 2369
rect 1870 2356 1876 2357
rect 1870 2352 1871 2356
rect 1875 2352 1876 2356
rect 1870 2351 1876 2352
rect 3590 2356 3596 2357
rect 3590 2352 3591 2356
rect 3595 2352 3596 2356
rect 3590 2351 3596 2352
rect 111 2334 115 2335
rect 111 2329 115 2330
rect 359 2334 363 2335
rect 359 2329 363 2330
rect 439 2334 443 2335
rect 439 2329 443 2330
rect 519 2334 523 2335
rect 519 2329 523 2330
rect 599 2334 603 2335
rect 599 2329 603 2330
rect 679 2334 683 2335
rect 679 2329 683 2330
rect 759 2334 763 2335
rect 759 2329 763 2330
rect 839 2334 843 2335
rect 839 2329 843 2330
rect 919 2334 923 2335
rect 919 2329 923 2330
rect 999 2334 1003 2335
rect 999 2329 1003 2330
rect 1071 2334 1075 2335
rect 1071 2329 1075 2330
rect 1079 2334 1083 2335
rect 1079 2329 1083 2330
rect 1151 2334 1155 2335
rect 1151 2329 1155 2330
rect 1159 2334 1163 2335
rect 1159 2329 1163 2330
rect 1231 2334 1235 2335
rect 1231 2329 1235 2330
rect 1239 2334 1243 2335
rect 1239 2329 1243 2330
rect 1311 2334 1315 2335
rect 1311 2329 1315 2330
rect 1319 2334 1323 2335
rect 1319 2329 1323 2330
rect 1391 2334 1395 2335
rect 1391 2329 1395 2330
rect 1471 2334 1475 2335
rect 1471 2329 1475 2330
rect 1831 2334 1835 2335
rect 1831 2329 1835 2330
rect 112 2301 114 2329
rect 360 2319 362 2329
rect 440 2319 442 2329
rect 520 2319 522 2329
rect 600 2319 602 2329
rect 680 2319 682 2329
rect 760 2319 762 2329
rect 840 2319 842 2329
rect 920 2319 922 2329
rect 1000 2319 1002 2329
rect 1080 2319 1082 2329
rect 1160 2319 1162 2329
rect 1240 2319 1242 2329
rect 1320 2319 1322 2329
rect 358 2318 364 2319
rect 358 2314 359 2318
rect 363 2314 364 2318
rect 358 2313 364 2314
rect 438 2318 444 2319
rect 438 2314 439 2318
rect 443 2314 444 2318
rect 438 2313 444 2314
rect 518 2318 524 2319
rect 518 2314 519 2318
rect 523 2314 524 2318
rect 518 2313 524 2314
rect 598 2318 604 2319
rect 598 2314 599 2318
rect 603 2314 604 2318
rect 598 2313 604 2314
rect 678 2318 684 2319
rect 678 2314 679 2318
rect 683 2314 684 2318
rect 678 2313 684 2314
rect 758 2318 764 2319
rect 758 2314 759 2318
rect 763 2314 764 2318
rect 758 2313 764 2314
rect 838 2318 844 2319
rect 838 2314 839 2318
rect 843 2314 844 2318
rect 838 2313 844 2314
rect 918 2318 924 2319
rect 918 2314 919 2318
rect 923 2314 924 2318
rect 918 2313 924 2314
rect 998 2318 1004 2319
rect 998 2314 999 2318
rect 1003 2314 1004 2318
rect 998 2313 1004 2314
rect 1078 2318 1084 2319
rect 1078 2314 1079 2318
rect 1083 2314 1084 2318
rect 1078 2313 1084 2314
rect 1158 2318 1164 2319
rect 1158 2314 1159 2318
rect 1163 2314 1164 2318
rect 1158 2313 1164 2314
rect 1238 2318 1244 2319
rect 1238 2314 1239 2318
rect 1243 2314 1244 2318
rect 1238 2313 1244 2314
rect 1318 2318 1324 2319
rect 1318 2314 1319 2318
rect 1323 2314 1324 2318
rect 1318 2313 1324 2314
rect 1832 2301 1834 2329
rect 1872 2319 1874 2351
rect 2150 2338 2156 2339
rect 2150 2334 2151 2338
rect 2155 2334 2156 2338
rect 2150 2333 2156 2334
rect 2246 2338 2252 2339
rect 2246 2334 2247 2338
rect 2251 2334 2252 2338
rect 2246 2333 2252 2334
rect 2350 2338 2356 2339
rect 2350 2334 2351 2338
rect 2355 2334 2356 2338
rect 2350 2333 2356 2334
rect 2462 2338 2468 2339
rect 2462 2334 2463 2338
rect 2467 2334 2468 2338
rect 2462 2333 2468 2334
rect 2582 2338 2588 2339
rect 2582 2334 2583 2338
rect 2587 2334 2588 2338
rect 2582 2333 2588 2334
rect 2710 2338 2716 2339
rect 2710 2334 2711 2338
rect 2715 2334 2716 2338
rect 2710 2333 2716 2334
rect 2854 2338 2860 2339
rect 2854 2334 2855 2338
rect 2859 2334 2860 2338
rect 2854 2333 2860 2334
rect 3014 2338 3020 2339
rect 3014 2334 3015 2338
rect 3019 2334 3020 2338
rect 3014 2333 3020 2334
rect 3182 2338 3188 2339
rect 3182 2334 3183 2338
rect 3187 2334 3188 2338
rect 3182 2333 3188 2334
rect 3358 2338 3364 2339
rect 3358 2334 3359 2338
rect 3363 2334 3364 2338
rect 3358 2333 3364 2334
rect 3510 2338 3516 2339
rect 3510 2334 3511 2338
rect 3515 2334 3516 2338
rect 3510 2333 3516 2334
rect 2152 2319 2154 2333
rect 2248 2319 2250 2333
rect 2352 2319 2354 2333
rect 2464 2319 2466 2333
rect 2584 2319 2586 2333
rect 2712 2319 2714 2333
rect 2856 2319 2858 2333
rect 3016 2319 3018 2333
rect 3184 2319 3186 2333
rect 3360 2319 3362 2333
rect 3512 2319 3514 2333
rect 3592 2319 3594 2351
rect 1871 2318 1875 2319
rect 1871 2313 1875 2314
rect 2151 2318 2155 2319
rect 2151 2313 2155 2314
rect 2247 2318 2251 2319
rect 2247 2313 2251 2314
rect 2279 2318 2283 2319
rect 2279 2313 2283 2314
rect 2351 2318 2355 2319
rect 2351 2313 2355 2314
rect 2359 2318 2363 2319
rect 2359 2313 2363 2314
rect 2439 2318 2443 2319
rect 2439 2313 2443 2314
rect 2463 2318 2467 2319
rect 2463 2313 2467 2314
rect 2519 2318 2523 2319
rect 2519 2313 2523 2314
rect 2583 2318 2587 2319
rect 2583 2313 2587 2314
rect 2599 2318 2603 2319
rect 2599 2313 2603 2314
rect 2679 2318 2683 2319
rect 2679 2313 2683 2314
rect 2711 2318 2715 2319
rect 2711 2313 2715 2314
rect 2759 2318 2763 2319
rect 2759 2313 2763 2314
rect 2847 2318 2851 2319
rect 2847 2313 2851 2314
rect 2855 2318 2859 2319
rect 2855 2313 2859 2314
rect 2935 2318 2939 2319
rect 2935 2313 2939 2314
rect 3015 2318 3019 2319
rect 3015 2313 3019 2314
rect 3183 2318 3187 2319
rect 3183 2313 3187 2314
rect 3359 2318 3363 2319
rect 3359 2313 3363 2314
rect 3511 2318 3515 2319
rect 3511 2313 3515 2314
rect 3591 2318 3595 2319
rect 3591 2313 3595 2314
rect 110 2300 116 2301
rect 110 2296 111 2300
rect 115 2296 116 2300
rect 110 2295 116 2296
rect 1830 2300 1836 2301
rect 1830 2296 1831 2300
rect 1835 2296 1836 2300
rect 1830 2295 1836 2296
rect 1872 2285 1874 2313
rect 2280 2303 2282 2313
rect 2360 2303 2362 2313
rect 2440 2303 2442 2313
rect 2520 2303 2522 2313
rect 2600 2303 2602 2313
rect 2680 2303 2682 2313
rect 2760 2303 2762 2313
rect 2848 2303 2850 2313
rect 2936 2303 2938 2313
rect 2278 2302 2284 2303
rect 2278 2298 2279 2302
rect 2283 2298 2284 2302
rect 2278 2297 2284 2298
rect 2358 2302 2364 2303
rect 2358 2298 2359 2302
rect 2363 2298 2364 2302
rect 2358 2297 2364 2298
rect 2438 2302 2444 2303
rect 2438 2298 2439 2302
rect 2443 2298 2444 2302
rect 2438 2297 2444 2298
rect 2518 2302 2524 2303
rect 2518 2298 2519 2302
rect 2523 2298 2524 2302
rect 2518 2297 2524 2298
rect 2598 2302 2604 2303
rect 2598 2298 2599 2302
rect 2603 2298 2604 2302
rect 2598 2297 2604 2298
rect 2678 2302 2684 2303
rect 2678 2298 2679 2302
rect 2683 2298 2684 2302
rect 2678 2297 2684 2298
rect 2758 2302 2764 2303
rect 2758 2298 2759 2302
rect 2763 2298 2764 2302
rect 2758 2297 2764 2298
rect 2846 2302 2852 2303
rect 2846 2298 2847 2302
rect 2851 2298 2852 2302
rect 2846 2297 2852 2298
rect 2934 2302 2940 2303
rect 2934 2298 2935 2302
rect 2939 2298 2940 2302
rect 2934 2297 2940 2298
rect 3592 2285 3594 2313
rect 1870 2284 1876 2285
rect 110 2283 116 2284
rect 110 2279 111 2283
rect 115 2279 116 2283
rect 1830 2283 1836 2284
rect 110 2278 116 2279
rect 350 2280 356 2281
rect 112 2259 114 2278
rect 350 2276 351 2280
rect 355 2276 356 2280
rect 350 2275 356 2276
rect 430 2280 436 2281
rect 430 2276 431 2280
rect 435 2276 436 2280
rect 430 2275 436 2276
rect 510 2280 516 2281
rect 510 2276 511 2280
rect 515 2276 516 2280
rect 510 2275 516 2276
rect 590 2280 596 2281
rect 590 2276 591 2280
rect 595 2276 596 2280
rect 590 2275 596 2276
rect 670 2280 676 2281
rect 670 2276 671 2280
rect 675 2276 676 2280
rect 670 2275 676 2276
rect 750 2280 756 2281
rect 750 2276 751 2280
rect 755 2276 756 2280
rect 750 2275 756 2276
rect 830 2280 836 2281
rect 830 2276 831 2280
rect 835 2276 836 2280
rect 830 2275 836 2276
rect 910 2280 916 2281
rect 910 2276 911 2280
rect 915 2276 916 2280
rect 910 2275 916 2276
rect 990 2280 996 2281
rect 990 2276 991 2280
rect 995 2276 996 2280
rect 990 2275 996 2276
rect 1070 2280 1076 2281
rect 1070 2276 1071 2280
rect 1075 2276 1076 2280
rect 1070 2275 1076 2276
rect 1150 2280 1156 2281
rect 1150 2276 1151 2280
rect 1155 2276 1156 2280
rect 1150 2275 1156 2276
rect 1230 2280 1236 2281
rect 1230 2276 1231 2280
rect 1235 2276 1236 2280
rect 1230 2275 1236 2276
rect 1310 2280 1316 2281
rect 1310 2276 1311 2280
rect 1315 2276 1316 2280
rect 1830 2279 1831 2283
rect 1835 2279 1836 2283
rect 1870 2280 1871 2284
rect 1875 2280 1876 2284
rect 1870 2279 1876 2280
rect 3590 2284 3596 2285
rect 3590 2280 3591 2284
rect 3595 2280 3596 2284
rect 3590 2279 3596 2280
rect 1830 2278 1836 2279
rect 1310 2275 1316 2276
rect 352 2259 354 2275
rect 432 2259 434 2275
rect 512 2259 514 2275
rect 592 2259 594 2275
rect 672 2259 674 2275
rect 752 2259 754 2275
rect 832 2259 834 2275
rect 912 2259 914 2275
rect 992 2259 994 2275
rect 1072 2259 1074 2275
rect 1152 2259 1154 2275
rect 1232 2259 1234 2275
rect 1312 2259 1314 2275
rect 1832 2259 1834 2278
rect 1870 2267 1876 2268
rect 1870 2263 1871 2267
rect 1875 2263 1876 2267
rect 3590 2267 3596 2268
rect 1870 2262 1876 2263
rect 2270 2264 2276 2265
rect 111 2258 115 2259
rect 111 2253 115 2254
rect 351 2258 355 2259
rect 351 2253 355 2254
rect 375 2258 379 2259
rect 375 2253 379 2254
rect 431 2258 435 2259
rect 431 2253 435 2254
rect 455 2258 459 2259
rect 455 2253 459 2254
rect 511 2258 515 2259
rect 511 2253 515 2254
rect 535 2258 539 2259
rect 535 2253 539 2254
rect 591 2258 595 2259
rect 591 2253 595 2254
rect 615 2258 619 2259
rect 615 2253 619 2254
rect 671 2258 675 2259
rect 671 2253 675 2254
rect 695 2258 699 2259
rect 695 2253 699 2254
rect 751 2258 755 2259
rect 751 2253 755 2254
rect 775 2258 779 2259
rect 775 2253 779 2254
rect 831 2258 835 2259
rect 831 2253 835 2254
rect 855 2258 859 2259
rect 855 2253 859 2254
rect 911 2258 915 2259
rect 911 2253 915 2254
rect 935 2258 939 2259
rect 935 2253 939 2254
rect 991 2258 995 2259
rect 991 2253 995 2254
rect 1015 2258 1019 2259
rect 1015 2253 1019 2254
rect 1071 2258 1075 2259
rect 1071 2253 1075 2254
rect 1095 2258 1099 2259
rect 1095 2253 1099 2254
rect 1151 2258 1155 2259
rect 1151 2253 1155 2254
rect 1175 2258 1179 2259
rect 1175 2253 1179 2254
rect 1231 2258 1235 2259
rect 1231 2253 1235 2254
rect 1255 2258 1259 2259
rect 1255 2253 1259 2254
rect 1311 2258 1315 2259
rect 1311 2253 1315 2254
rect 1831 2258 1835 2259
rect 1831 2253 1835 2254
rect 112 2234 114 2253
rect 376 2237 378 2253
rect 456 2237 458 2253
rect 536 2237 538 2253
rect 616 2237 618 2253
rect 696 2237 698 2253
rect 776 2237 778 2253
rect 856 2237 858 2253
rect 936 2237 938 2253
rect 1016 2237 1018 2253
rect 1096 2237 1098 2253
rect 1176 2237 1178 2253
rect 1256 2237 1258 2253
rect 374 2236 380 2237
rect 110 2233 116 2234
rect 110 2229 111 2233
rect 115 2229 116 2233
rect 374 2232 375 2236
rect 379 2232 380 2236
rect 374 2231 380 2232
rect 454 2236 460 2237
rect 454 2232 455 2236
rect 459 2232 460 2236
rect 454 2231 460 2232
rect 534 2236 540 2237
rect 534 2232 535 2236
rect 539 2232 540 2236
rect 534 2231 540 2232
rect 614 2236 620 2237
rect 614 2232 615 2236
rect 619 2232 620 2236
rect 614 2231 620 2232
rect 694 2236 700 2237
rect 694 2232 695 2236
rect 699 2232 700 2236
rect 694 2231 700 2232
rect 774 2236 780 2237
rect 774 2232 775 2236
rect 779 2232 780 2236
rect 774 2231 780 2232
rect 854 2236 860 2237
rect 854 2232 855 2236
rect 859 2232 860 2236
rect 854 2231 860 2232
rect 934 2236 940 2237
rect 934 2232 935 2236
rect 939 2232 940 2236
rect 934 2231 940 2232
rect 1014 2236 1020 2237
rect 1014 2232 1015 2236
rect 1019 2232 1020 2236
rect 1014 2231 1020 2232
rect 1094 2236 1100 2237
rect 1094 2232 1095 2236
rect 1099 2232 1100 2236
rect 1094 2231 1100 2232
rect 1174 2236 1180 2237
rect 1174 2232 1175 2236
rect 1179 2232 1180 2236
rect 1174 2231 1180 2232
rect 1254 2236 1260 2237
rect 1254 2232 1255 2236
rect 1259 2232 1260 2236
rect 1832 2234 1834 2253
rect 1872 2243 1874 2262
rect 2270 2260 2271 2264
rect 2275 2260 2276 2264
rect 2270 2259 2276 2260
rect 2350 2264 2356 2265
rect 2350 2260 2351 2264
rect 2355 2260 2356 2264
rect 2350 2259 2356 2260
rect 2430 2264 2436 2265
rect 2430 2260 2431 2264
rect 2435 2260 2436 2264
rect 2430 2259 2436 2260
rect 2510 2264 2516 2265
rect 2510 2260 2511 2264
rect 2515 2260 2516 2264
rect 2510 2259 2516 2260
rect 2590 2264 2596 2265
rect 2590 2260 2591 2264
rect 2595 2260 2596 2264
rect 2590 2259 2596 2260
rect 2670 2264 2676 2265
rect 2670 2260 2671 2264
rect 2675 2260 2676 2264
rect 2670 2259 2676 2260
rect 2750 2264 2756 2265
rect 2750 2260 2751 2264
rect 2755 2260 2756 2264
rect 2750 2259 2756 2260
rect 2838 2264 2844 2265
rect 2838 2260 2839 2264
rect 2843 2260 2844 2264
rect 2838 2259 2844 2260
rect 2926 2264 2932 2265
rect 2926 2260 2927 2264
rect 2931 2260 2932 2264
rect 3590 2263 3591 2267
rect 3595 2263 3596 2267
rect 3590 2262 3596 2263
rect 2926 2259 2932 2260
rect 2272 2243 2274 2259
rect 2352 2243 2354 2259
rect 2432 2243 2434 2259
rect 2512 2243 2514 2259
rect 2592 2243 2594 2259
rect 2672 2243 2674 2259
rect 2752 2243 2754 2259
rect 2840 2243 2842 2259
rect 2928 2243 2930 2259
rect 3592 2243 3594 2262
rect 1871 2242 1875 2243
rect 1871 2237 1875 2238
rect 2271 2242 2275 2243
rect 2271 2237 2275 2238
rect 2311 2242 2315 2243
rect 2311 2237 2315 2238
rect 2351 2242 2355 2243
rect 2351 2237 2355 2238
rect 2399 2242 2403 2243
rect 2399 2237 2403 2238
rect 2431 2242 2435 2243
rect 2431 2237 2435 2238
rect 2495 2242 2499 2243
rect 2495 2237 2499 2238
rect 2511 2242 2515 2243
rect 2511 2237 2515 2238
rect 2591 2242 2595 2243
rect 2591 2237 2595 2238
rect 2599 2242 2603 2243
rect 2599 2237 2603 2238
rect 2671 2242 2675 2243
rect 2671 2237 2675 2238
rect 2719 2242 2723 2243
rect 2719 2237 2723 2238
rect 2751 2242 2755 2243
rect 2751 2237 2755 2238
rect 2839 2242 2843 2243
rect 2839 2237 2843 2238
rect 2855 2242 2859 2243
rect 2855 2237 2859 2238
rect 2927 2242 2931 2243
rect 2927 2237 2931 2238
rect 3007 2242 3011 2243
rect 3007 2237 3011 2238
rect 3175 2242 3179 2243
rect 3175 2237 3179 2238
rect 3351 2242 3355 2243
rect 3351 2237 3355 2238
rect 3503 2242 3507 2243
rect 3503 2237 3507 2238
rect 3591 2242 3595 2243
rect 3591 2237 3595 2238
rect 1254 2231 1260 2232
rect 1830 2233 1836 2234
rect 110 2228 116 2229
rect 1830 2229 1831 2233
rect 1835 2229 1836 2233
rect 1830 2228 1836 2229
rect 1872 2218 1874 2237
rect 2312 2221 2314 2237
rect 2400 2221 2402 2237
rect 2496 2221 2498 2237
rect 2600 2221 2602 2237
rect 2720 2221 2722 2237
rect 2856 2221 2858 2237
rect 3008 2221 3010 2237
rect 3176 2221 3178 2237
rect 3352 2221 3354 2237
rect 3504 2221 3506 2237
rect 2310 2220 2316 2221
rect 1870 2217 1876 2218
rect 110 2216 116 2217
rect 110 2212 111 2216
rect 115 2212 116 2216
rect 110 2211 116 2212
rect 1830 2216 1836 2217
rect 1830 2212 1831 2216
rect 1835 2212 1836 2216
rect 1870 2213 1871 2217
rect 1875 2213 1876 2217
rect 2310 2216 2311 2220
rect 2315 2216 2316 2220
rect 2310 2215 2316 2216
rect 2398 2220 2404 2221
rect 2398 2216 2399 2220
rect 2403 2216 2404 2220
rect 2398 2215 2404 2216
rect 2494 2220 2500 2221
rect 2494 2216 2495 2220
rect 2499 2216 2500 2220
rect 2494 2215 2500 2216
rect 2598 2220 2604 2221
rect 2598 2216 2599 2220
rect 2603 2216 2604 2220
rect 2598 2215 2604 2216
rect 2718 2220 2724 2221
rect 2718 2216 2719 2220
rect 2723 2216 2724 2220
rect 2718 2215 2724 2216
rect 2854 2220 2860 2221
rect 2854 2216 2855 2220
rect 2859 2216 2860 2220
rect 2854 2215 2860 2216
rect 3006 2220 3012 2221
rect 3006 2216 3007 2220
rect 3011 2216 3012 2220
rect 3006 2215 3012 2216
rect 3174 2220 3180 2221
rect 3174 2216 3175 2220
rect 3179 2216 3180 2220
rect 3174 2215 3180 2216
rect 3350 2220 3356 2221
rect 3350 2216 3351 2220
rect 3355 2216 3356 2220
rect 3350 2215 3356 2216
rect 3502 2220 3508 2221
rect 3502 2216 3503 2220
rect 3507 2216 3508 2220
rect 3592 2218 3594 2237
rect 3502 2215 3508 2216
rect 3590 2217 3596 2218
rect 1870 2212 1876 2213
rect 3590 2213 3591 2217
rect 3595 2213 3596 2217
rect 3590 2212 3596 2213
rect 1830 2211 1836 2212
rect 112 2171 114 2211
rect 382 2198 388 2199
rect 382 2194 383 2198
rect 387 2194 388 2198
rect 382 2193 388 2194
rect 462 2198 468 2199
rect 462 2194 463 2198
rect 467 2194 468 2198
rect 462 2193 468 2194
rect 542 2198 548 2199
rect 542 2194 543 2198
rect 547 2194 548 2198
rect 542 2193 548 2194
rect 622 2198 628 2199
rect 622 2194 623 2198
rect 627 2194 628 2198
rect 622 2193 628 2194
rect 702 2198 708 2199
rect 702 2194 703 2198
rect 707 2194 708 2198
rect 702 2193 708 2194
rect 782 2198 788 2199
rect 782 2194 783 2198
rect 787 2194 788 2198
rect 782 2193 788 2194
rect 862 2198 868 2199
rect 862 2194 863 2198
rect 867 2194 868 2198
rect 862 2193 868 2194
rect 942 2198 948 2199
rect 942 2194 943 2198
rect 947 2194 948 2198
rect 942 2193 948 2194
rect 1022 2198 1028 2199
rect 1022 2194 1023 2198
rect 1027 2194 1028 2198
rect 1022 2193 1028 2194
rect 1102 2198 1108 2199
rect 1102 2194 1103 2198
rect 1107 2194 1108 2198
rect 1102 2193 1108 2194
rect 1182 2198 1188 2199
rect 1182 2194 1183 2198
rect 1187 2194 1188 2198
rect 1182 2193 1188 2194
rect 1262 2198 1268 2199
rect 1262 2194 1263 2198
rect 1267 2194 1268 2198
rect 1262 2193 1268 2194
rect 384 2171 386 2193
rect 464 2171 466 2193
rect 544 2171 546 2193
rect 624 2171 626 2193
rect 704 2171 706 2193
rect 784 2171 786 2193
rect 864 2171 866 2193
rect 944 2171 946 2193
rect 1024 2171 1026 2193
rect 1104 2171 1106 2193
rect 1184 2171 1186 2193
rect 1264 2171 1266 2193
rect 1832 2171 1834 2211
rect 1870 2200 1876 2201
rect 1870 2196 1871 2200
rect 1875 2196 1876 2200
rect 1870 2195 1876 2196
rect 3590 2200 3596 2201
rect 3590 2196 3591 2200
rect 3595 2196 3596 2200
rect 3590 2195 3596 2196
rect 111 2170 115 2171
rect 111 2165 115 2166
rect 311 2170 315 2171
rect 311 2165 315 2166
rect 383 2170 387 2171
rect 383 2165 387 2166
rect 407 2170 411 2171
rect 407 2165 411 2166
rect 463 2170 467 2171
rect 463 2165 467 2166
rect 503 2170 507 2171
rect 503 2165 507 2166
rect 543 2170 547 2171
rect 543 2165 547 2166
rect 599 2170 603 2171
rect 599 2165 603 2166
rect 623 2170 627 2171
rect 623 2165 627 2166
rect 687 2170 691 2171
rect 687 2165 691 2166
rect 703 2170 707 2171
rect 703 2165 707 2166
rect 775 2170 779 2171
rect 775 2165 779 2166
rect 783 2170 787 2171
rect 783 2165 787 2166
rect 863 2170 867 2171
rect 863 2165 867 2166
rect 943 2170 947 2171
rect 943 2165 947 2166
rect 951 2170 955 2171
rect 951 2165 955 2166
rect 1023 2170 1027 2171
rect 1023 2165 1027 2166
rect 1039 2170 1043 2171
rect 1039 2165 1043 2166
rect 1103 2170 1107 2171
rect 1103 2165 1107 2166
rect 1127 2170 1131 2171
rect 1127 2165 1131 2166
rect 1183 2170 1187 2171
rect 1183 2165 1187 2166
rect 1223 2170 1227 2171
rect 1223 2165 1227 2166
rect 1263 2170 1267 2171
rect 1263 2165 1267 2166
rect 1831 2170 1835 2171
rect 1831 2165 1835 2166
rect 112 2137 114 2165
rect 312 2155 314 2165
rect 408 2155 410 2165
rect 504 2155 506 2165
rect 600 2155 602 2165
rect 688 2155 690 2165
rect 776 2155 778 2165
rect 864 2155 866 2165
rect 952 2155 954 2165
rect 1040 2155 1042 2165
rect 1128 2155 1130 2165
rect 1224 2155 1226 2165
rect 310 2154 316 2155
rect 310 2150 311 2154
rect 315 2150 316 2154
rect 310 2149 316 2150
rect 406 2154 412 2155
rect 406 2150 407 2154
rect 411 2150 412 2154
rect 406 2149 412 2150
rect 502 2154 508 2155
rect 502 2150 503 2154
rect 507 2150 508 2154
rect 502 2149 508 2150
rect 598 2154 604 2155
rect 598 2150 599 2154
rect 603 2150 604 2154
rect 598 2149 604 2150
rect 686 2154 692 2155
rect 686 2150 687 2154
rect 691 2150 692 2154
rect 686 2149 692 2150
rect 774 2154 780 2155
rect 774 2150 775 2154
rect 779 2150 780 2154
rect 774 2149 780 2150
rect 862 2154 868 2155
rect 862 2150 863 2154
rect 867 2150 868 2154
rect 862 2149 868 2150
rect 950 2154 956 2155
rect 950 2150 951 2154
rect 955 2150 956 2154
rect 950 2149 956 2150
rect 1038 2154 1044 2155
rect 1038 2150 1039 2154
rect 1043 2150 1044 2154
rect 1038 2149 1044 2150
rect 1126 2154 1132 2155
rect 1126 2150 1127 2154
rect 1131 2150 1132 2154
rect 1126 2149 1132 2150
rect 1222 2154 1228 2155
rect 1222 2150 1223 2154
rect 1227 2150 1228 2154
rect 1222 2149 1228 2150
rect 1832 2137 1834 2165
rect 1872 2163 1874 2195
rect 2318 2182 2324 2183
rect 2318 2178 2319 2182
rect 2323 2178 2324 2182
rect 2318 2177 2324 2178
rect 2406 2182 2412 2183
rect 2406 2178 2407 2182
rect 2411 2178 2412 2182
rect 2406 2177 2412 2178
rect 2502 2182 2508 2183
rect 2502 2178 2503 2182
rect 2507 2178 2508 2182
rect 2502 2177 2508 2178
rect 2606 2182 2612 2183
rect 2606 2178 2607 2182
rect 2611 2178 2612 2182
rect 2606 2177 2612 2178
rect 2726 2182 2732 2183
rect 2726 2178 2727 2182
rect 2731 2178 2732 2182
rect 2726 2177 2732 2178
rect 2862 2182 2868 2183
rect 2862 2178 2863 2182
rect 2867 2178 2868 2182
rect 2862 2177 2868 2178
rect 3014 2182 3020 2183
rect 3014 2178 3015 2182
rect 3019 2178 3020 2182
rect 3014 2177 3020 2178
rect 3182 2182 3188 2183
rect 3182 2178 3183 2182
rect 3187 2178 3188 2182
rect 3182 2177 3188 2178
rect 3358 2182 3364 2183
rect 3358 2178 3359 2182
rect 3363 2178 3364 2182
rect 3358 2177 3364 2178
rect 3510 2182 3516 2183
rect 3510 2178 3511 2182
rect 3515 2178 3516 2182
rect 3510 2177 3516 2178
rect 2320 2163 2322 2177
rect 2408 2163 2410 2177
rect 2504 2163 2506 2177
rect 2608 2163 2610 2177
rect 2728 2163 2730 2177
rect 2864 2163 2866 2177
rect 3016 2163 3018 2177
rect 3184 2163 3186 2177
rect 3360 2163 3362 2177
rect 3512 2163 3514 2177
rect 3592 2163 3594 2195
rect 1871 2162 1875 2163
rect 1871 2157 1875 2158
rect 1903 2162 1907 2163
rect 1903 2157 1907 2158
rect 1983 2162 1987 2163
rect 1983 2157 1987 2158
rect 2111 2162 2115 2163
rect 2111 2157 2115 2158
rect 2247 2162 2251 2163
rect 2247 2157 2251 2158
rect 2319 2162 2323 2163
rect 2319 2157 2323 2158
rect 2391 2162 2395 2163
rect 2391 2157 2395 2158
rect 2407 2162 2411 2163
rect 2407 2157 2411 2158
rect 2503 2162 2507 2163
rect 2503 2157 2507 2158
rect 2543 2162 2547 2163
rect 2543 2157 2547 2158
rect 2607 2162 2611 2163
rect 2607 2157 2611 2158
rect 2695 2162 2699 2163
rect 2695 2157 2699 2158
rect 2727 2162 2731 2163
rect 2727 2157 2731 2158
rect 2847 2162 2851 2163
rect 2847 2157 2851 2158
rect 2863 2162 2867 2163
rect 2863 2157 2867 2158
rect 3007 2162 3011 2163
rect 3007 2157 3011 2158
rect 3015 2162 3019 2163
rect 3015 2157 3019 2158
rect 3175 2162 3179 2163
rect 3175 2157 3179 2158
rect 3183 2162 3187 2163
rect 3183 2157 3187 2158
rect 3351 2162 3355 2163
rect 3351 2157 3355 2158
rect 3359 2162 3363 2163
rect 3359 2157 3363 2158
rect 3511 2162 3515 2163
rect 3511 2157 3515 2158
rect 3591 2162 3595 2163
rect 3591 2157 3595 2158
rect 110 2136 116 2137
rect 110 2132 111 2136
rect 115 2132 116 2136
rect 110 2131 116 2132
rect 1830 2136 1836 2137
rect 1830 2132 1831 2136
rect 1835 2132 1836 2136
rect 1830 2131 1836 2132
rect 1872 2129 1874 2157
rect 1904 2147 1906 2157
rect 1984 2147 1986 2157
rect 2112 2147 2114 2157
rect 2248 2147 2250 2157
rect 2392 2147 2394 2157
rect 2544 2147 2546 2157
rect 2696 2147 2698 2157
rect 2848 2147 2850 2157
rect 3008 2147 3010 2157
rect 3176 2147 3178 2157
rect 3352 2147 3354 2157
rect 3512 2147 3514 2157
rect 1902 2146 1908 2147
rect 1902 2142 1903 2146
rect 1907 2142 1908 2146
rect 1902 2141 1908 2142
rect 1982 2146 1988 2147
rect 1982 2142 1983 2146
rect 1987 2142 1988 2146
rect 1982 2141 1988 2142
rect 2110 2146 2116 2147
rect 2110 2142 2111 2146
rect 2115 2142 2116 2146
rect 2110 2141 2116 2142
rect 2246 2146 2252 2147
rect 2246 2142 2247 2146
rect 2251 2142 2252 2146
rect 2246 2141 2252 2142
rect 2390 2146 2396 2147
rect 2390 2142 2391 2146
rect 2395 2142 2396 2146
rect 2390 2141 2396 2142
rect 2542 2146 2548 2147
rect 2542 2142 2543 2146
rect 2547 2142 2548 2146
rect 2542 2141 2548 2142
rect 2694 2146 2700 2147
rect 2694 2142 2695 2146
rect 2699 2142 2700 2146
rect 2694 2141 2700 2142
rect 2846 2146 2852 2147
rect 2846 2142 2847 2146
rect 2851 2142 2852 2146
rect 2846 2141 2852 2142
rect 3006 2146 3012 2147
rect 3006 2142 3007 2146
rect 3011 2142 3012 2146
rect 3006 2141 3012 2142
rect 3174 2146 3180 2147
rect 3174 2142 3175 2146
rect 3179 2142 3180 2146
rect 3174 2141 3180 2142
rect 3350 2146 3356 2147
rect 3350 2142 3351 2146
rect 3355 2142 3356 2146
rect 3350 2141 3356 2142
rect 3510 2146 3516 2147
rect 3510 2142 3511 2146
rect 3515 2142 3516 2146
rect 3510 2141 3516 2142
rect 3592 2129 3594 2157
rect 1870 2128 1876 2129
rect 1870 2124 1871 2128
rect 1875 2124 1876 2128
rect 1870 2123 1876 2124
rect 3590 2128 3596 2129
rect 3590 2124 3591 2128
rect 3595 2124 3596 2128
rect 3590 2123 3596 2124
rect 110 2119 116 2120
rect 110 2115 111 2119
rect 115 2115 116 2119
rect 1830 2119 1836 2120
rect 110 2114 116 2115
rect 302 2116 308 2117
rect 112 2083 114 2114
rect 302 2112 303 2116
rect 307 2112 308 2116
rect 302 2111 308 2112
rect 398 2116 404 2117
rect 398 2112 399 2116
rect 403 2112 404 2116
rect 398 2111 404 2112
rect 494 2116 500 2117
rect 494 2112 495 2116
rect 499 2112 500 2116
rect 494 2111 500 2112
rect 590 2116 596 2117
rect 590 2112 591 2116
rect 595 2112 596 2116
rect 590 2111 596 2112
rect 678 2116 684 2117
rect 678 2112 679 2116
rect 683 2112 684 2116
rect 678 2111 684 2112
rect 766 2116 772 2117
rect 766 2112 767 2116
rect 771 2112 772 2116
rect 766 2111 772 2112
rect 854 2116 860 2117
rect 854 2112 855 2116
rect 859 2112 860 2116
rect 854 2111 860 2112
rect 942 2116 948 2117
rect 942 2112 943 2116
rect 947 2112 948 2116
rect 942 2111 948 2112
rect 1030 2116 1036 2117
rect 1030 2112 1031 2116
rect 1035 2112 1036 2116
rect 1030 2111 1036 2112
rect 1118 2116 1124 2117
rect 1118 2112 1119 2116
rect 1123 2112 1124 2116
rect 1118 2111 1124 2112
rect 1214 2116 1220 2117
rect 1214 2112 1215 2116
rect 1219 2112 1220 2116
rect 1830 2115 1831 2119
rect 1835 2115 1836 2119
rect 1830 2114 1836 2115
rect 1214 2111 1220 2112
rect 304 2083 306 2111
rect 400 2083 402 2111
rect 496 2083 498 2111
rect 592 2083 594 2111
rect 680 2083 682 2111
rect 768 2083 770 2111
rect 856 2083 858 2111
rect 944 2083 946 2111
rect 1032 2083 1034 2111
rect 1120 2083 1122 2111
rect 1216 2083 1218 2111
rect 1832 2083 1834 2114
rect 1870 2111 1876 2112
rect 1870 2107 1871 2111
rect 1875 2107 1876 2111
rect 3590 2111 3596 2112
rect 1870 2106 1876 2107
rect 1894 2108 1900 2109
rect 111 2082 115 2083
rect 111 2077 115 2078
rect 207 2082 211 2083
rect 207 2077 211 2078
rect 303 2082 307 2083
rect 303 2077 307 2078
rect 327 2082 331 2083
rect 327 2077 331 2078
rect 399 2082 403 2083
rect 399 2077 403 2078
rect 447 2082 451 2083
rect 447 2077 451 2078
rect 495 2082 499 2083
rect 495 2077 499 2078
rect 575 2082 579 2083
rect 575 2077 579 2078
rect 591 2082 595 2083
rect 591 2077 595 2078
rect 679 2082 683 2083
rect 679 2077 683 2078
rect 703 2082 707 2083
rect 703 2077 707 2078
rect 767 2082 771 2083
rect 767 2077 771 2078
rect 823 2082 827 2083
rect 823 2077 827 2078
rect 855 2082 859 2083
rect 855 2077 859 2078
rect 943 2082 947 2083
rect 943 2077 947 2078
rect 1031 2082 1035 2083
rect 1031 2077 1035 2078
rect 1063 2082 1067 2083
rect 1063 2077 1067 2078
rect 1119 2082 1123 2083
rect 1119 2077 1123 2078
rect 1175 2082 1179 2083
rect 1175 2077 1179 2078
rect 1215 2082 1219 2083
rect 1215 2077 1219 2078
rect 1279 2082 1283 2083
rect 1279 2077 1283 2078
rect 1375 2082 1379 2083
rect 1375 2077 1379 2078
rect 1471 2082 1475 2083
rect 1471 2077 1475 2078
rect 1567 2082 1571 2083
rect 1567 2077 1571 2078
rect 1663 2082 1667 2083
rect 1663 2077 1667 2078
rect 1743 2082 1747 2083
rect 1743 2077 1747 2078
rect 1831 2082 1835 2083
rect 1872 2079 1874 2106
rect 1894 2104 1895 2108
rect 1899 2104 1900 2108
rect 1894 2103 1900 2104
rect 1974 2108 1980 2109
rect 1974 2104 1975 2108
rect 1979 2104 1980 2108
rect 1974 2103 1980 2104
rect 2102 2108 2108 2109
rect 2102 2104 2103 2108
rect 2107 2104 2108 2108
rect 2102 2103 2108 2104
rect 2238 2108 2244 2109
rect 2238 2104 2239 2108
rect 2243 2104 2244 2108
rect 2238 2103 2244 2104
rect 2382 2108 2388 2109
rect 2382 2104 2383 2108
rect 2387 2104 2388 2108
rect 2382 2103 2388 2104
rect 2534 2108 2540 2109
rect 2534 2104 2535 2108
rect 2539 2104 2540 2108
rect 2534 2103 2540 2104
rect 2686 2108 2692 2109
rect 2686 2104 2687 2108
rect 2691 2104 2692 2108
rect 2686 2103 2692 2104
rect 2838 2108 2844 2109
rect 2838 2104 2839 2108
rect 2843 2104 2844 2108
rect 2838 2103 2844 2104
rect 2998 2108 3004 2109
rect 2998 2104 2999 2108
rect 3003 2104 3004 2108
rect 2998 2103 3004 2104
rect 3166 2108 3172 2109
rect 3166 2104 3167 2108
rect 3171 2104 3172 2108
rect 3166 2103 3172 2104
rect 3342 2108 3348 2109
rect 3342 2104 3343 2108
rect 3347 2104 3348 2108
rect 3342 2103 3348 2104
rect 3502 2108 3508 2109
rect 3502 2104 3503 2108
rect 3507 2104 3508 2108
rect 3590 2107 3591 2111
rect 3595 2107 3596 2111
rect 3590 2106 3596 2107
rect 3502 2103 3508 2104
rect 1896 2079 1898 2103
rect 1976 2079 1978 2103
rect 2104 2079 2106 2103
rect 2240 2079 2242 2103
rect 2384 2079 2386 2103
rect 2536 2079 2538 2103
rect 2688 2079 2690 2103
rect 2840 2079 2842 2103
rect 3000 2079 3002 2103
rect 3168 2079 3170 2103
rect 3344 2079 3346 2103
rect 3504 2079 3506 2103
rect 3592 2079 3594 2106
rect 1831 2077 1835 2078
rect 1871 2078 1875 2079
rect 112 2058 114 2077
rect 208 2061 210 2077
rect 328 2061 330 2077
rect 448 2061 450 2077
rect 576 2061 578 2077
rect 704 2061 706 2077
rect 824 2061 826 2077
rect 944 2061 946 2077
rect 1064 2061 1066 2077
rect 1176 2061 1178 2077
rect 1280 2061 1282 2077
rect 1376 2061 1378 2077
rect 1472 2061 1474 2077
rect 1568 2061 1570 2077
rect 1664 2061 1666 2077
rect 1744 2061 1746 2077
rect 206 2060 212 2061
rect 110 2057 116 2058
rect 110 2053 111 2057
rect 115 2053 116 2057
rect 206 2056 207 2060
rect 211 2056 212 2060
rect 206 2055 212 2056
rect 326 2060 332 2061
rect 326 2056 327 2060
rect 331 2056 332 2060
rect 326 2055 332 2056
rect 446 2060 452 2061
rect 446 2056 447 2060
rect 451 2056 452 2060
rect 446 2055 452 2056
rect 574 2060 580 2061
rect 574 2056 575 2060
rect 579 2056 580 2060
rect 574 2055 580 2056
rect 702 2060 708 2061
rect 702 2056 703 2060
rect 707 2056 708 2060
rect 702 2055 708 2056
rect 822 2060 828 2061
rect 822 2056 823 2060
rect 827 2056 828 2060
rect 822 2055 828 2056
rect 942 2060 948 2061
rect 942 2056 943 2060
rect 947 2056 948 2060
rect 942 2055 948 2056
rect 1062 2060 1068 2061
rect 1062 2056 1063 2060
rect 1067 2056 1068 2060
rect 1062 2055 1068 2056
rect 1174 2060 1180 2061
rect 1174 2056 1175 2060
rect 1179 2056 1180 2060
rect 1174 2055 1180 2056
rect 1278 2060 1284 2061
rect 1278 2056 1279 2060
rect 1283 2056 1284 2060
rect 1278 2055 1284 2056
rect 1374 2060 1380 2061
rect 1374 2056 1375 2060
rect 1379 2056 1380 2060
rect 1374 2055 1380 2056
rect 1470 2060 1476 2061
rect 1470 2056 1471 2060
rect 1475 2056 1476 2060
rect 1470 2055 1476 2056
rect 1566 2060 1572 2061
rect 1566 2056 1567 2060
rect 1571 2056 1572 2060
rect 1566 2055 1572 2056
rect 1662 2060 1668 2061
rect 1662 2056 1663 2060
rect 1667 2056 1668 2060
rect 1662 2055 1668 2056
rect 1742 2060 1748 2061
rect 1742 2056 1743 2060
rect 1747 2056 1748 2060
rect 1832 2058 1834 2077
rect 1871 2073 1875 2074
rect 1895 2078 1899 2079
rect 1895 2073 1899 2074
rect 1967 2078 1971 2079
rect 1967 2073 1971 2074
rect 1975 2078 1979 2079
rect 1975 2073 1979 2074
rect 2103 2078 2107 2079
rect 2103 2073 2107 2074
rect 2215 2078 2219 2079
rect 2215 2073 2219 2074
rect 2239 2078 2243 2079
rect 2239 2073 2243 2074
rect 2383 2078 2387 2079
rect 2383 2073 2387 2074
rect 2447 2078 2451 2079
rect 2447 2073 2451 2074
rect 2535 2078 2539 2079
rect 2535 2073 2539 2074
rect 2655 2078 2659 2079
rect 2655 2073 2659 2074
rect 2687 2078 2691 2079
rect 2687 2073 2691 2074
rect 2839 2078 2843 2079
rect 2839 2073 2843 2074
rect 2999 2078 3003 2079
rect 2999 2073 3003 2074
rect 3143 2078 3147 2079
rect 3143 2073 3147 2074
rect 3167 2078 3171 2079
rect 3167 2073 3171 2074
rect 3271 2078 3275 2079
rect 3271 2073 3275 2074
rect 3343 2078 3347 2079
rect 3343 2073 3347 2074
rect 3399 2078 3403 2079
rect 3399 2073 3403 2074
rect 3503 2078 3507 2079
rect 3503 2073 3507 2074
rect 3591 2078 3595 2079
rect 3591 2073 3595 2074
rect 1742 2055 1748 2056
rect 1830 2057 1836 2058
rect 110 2052 116 2053
rect 1830 2053 1831 2057
rect 1835 2053 1836 2057
rect 1872 2054 1874 2073
rect 1968 2057 1970 2073
rect 2216 2057 2218 2073
rect 2448 2057 2450 2073
rect 2656 2057 2658 2073
rect 2840 2057 2842 2073
rect 3000 2057 3002 2073
rect 3144 2057 3146 2073
rect 3272 2057 3274 2073
rect 3400 2057 3402 2073
rect 3504 2057 3506 2073
rect 1966 2056 1972 2057
rect 1830 2052 1836 2053
rect 1870 2053 1876 2054
rect 1870 2049 1871 2053
rect 1875 2049 1876 2053
rect 1966 2052 1967 2056
rect 1971 2052 1972 2056
rect 1966 2051 1972 2052
rect 2214 2056 2220 2057
rect 2214 2052 2215 2056
rect 2219 2052 2220 2056
rect 2214 2051 2220 2052
rect 2446 2056 2452 2057
rect 2446 2052 2447 2056
rect 2451 2052 2452 2056
rect 2446 2051 2452 2052
rect 2654 2056 2660 2057
rect 2654 2052 2655 2056
rect 2659 2052 2660 2056
rect 2654 2051 2660 2052
rect 2838 2056 2844 2057
rect 2838 2052 2839 2056
rect 2843 2052 2844 2056
rect 2838 2051 2844 2052
rect 2998 2056 3004 2057
rect 2998 2052 2999 2056
rect 3003 2052 3004 2056
rect 2998 2051 3004 2052
rect 3142 2056 3148 2057
rect 3142 2052 3143 2056
rect 3147 2052 3148 2056
rect 3142 2051 3148 2052
rect 3270 2056 3276 2057
rect 3270 2052 3271 2056
rect 3275 2052 3276 2056
rect 3270 2051 3276 2052
rect 3398 2056 3404 2057
rect 3398 2052 3399 2056
rect 3403 2052 3404 2056
rect 3398 2051 3404 2052
rect 3502 2056 3508 2057
rect 3502 2052 3503 2056
rect 3507 2052 3508 2056
rect 3592 2054 3594 2073
rect 3502 2051 3508 2052
rect 3590 2053 3596 2054
rect 1870 2048 1876 2049
rect 3590 2049 3591 2053
rect 3595 2049 3596 2053
rect 3590 2048 3596 2049
rect 110 2040 116 2041
rect 110 2036 111 2040
rect 115 2036 116 2040
rect 110 2035 116 2036
rect 1830 2040 1836 2041
rect 1830 2036 1831 2040
rect 1835 2036 1836 2040
rect 1830 2035 1836 2036
rect 1870 2036 1876 2037
rect 112 2003 114 2035
rect 214 2022 220 2023
rect 214 2018 215 2022
rect 219 2018 220 2022
rect 214 2017 220 2018
rect 334 2022 340 2023
rect 334 2018 335 2022
rect 339 2018 340 2022
rect 334 2017 340 2018
rect 454 2022 460 2023
rect 454 2018 455 2022
rect 459 2018 460 2022
rect 454 2017 460 2018
rect 582 2022 588 2023
rect 582 2018 583 2022
rect 587 2018 588 2022
rect 582 2017 588 2018
rect 710 2022 716 2023
rect 710 2018 711 2022
rect 715 2018 716 2022
rect 710 2017 716 2018
rect 830 2022 836 2023
rect 830 2018 831 2022
rect 835 2018 836 2022
rect 830 2017 836 2018
rect 950 2022 956 2023
rect 950 2018 951 2022
rect 955 2018 956 2022
rect 950 2017 956 2018
rect 1070 2022 1076 2023
rect 1070 2018 1071 2022
rect 1075 2018 1076 2022
rect 1070 2017 1076 2018
rect 1182 2022 1188 2023
rect 1182 2018 1183 2022
rect 1187 2018 1188 2022
rect 1182 2017 1188 2018
rect 1286 2022 1292 2023
rect 1286 2018 1287 2022
rect 1291 2018 1292 2022
rect 1286 2017 1292 2018
rect 1382 2022 1388 2023
rect 1382 2018 1383 2022
rect 1387 2018 1388 2022
rect 1382 2017 1388 2018
rect 1478 2022 1484 2023
rect 1478 2018 1479 2022
rect 1483 2018 1484 2022
rect 1478 2017 1484 2018
rect 1574 2022 1580 2023
rect 1574 2018 1575 2022
rect 1579 2018 1580 2022
rect 1574 2017 1580 2018
rect 1670 2022 1676 2023
rect 1670 2018 1671 2022
rect 1675 2018 1676 2022
rect 1670 2017 1676 2018
rect 1750 2022 1756 2023
rect 1750 2018 1751 2022
rect 1755 2018 1756 2022
rect 1750 2017 1756 2018
rect 216 2003 218 2017
rect 336 2003 338 2017
rect 456 2003 458 2017
rect 584 2003 586 2017
rect 712 2003 714 2017
rect 832 2003 834 2017
rect 952 2003 954 2017
rect 1072 2003 1074 2017
rect 1184 2003 1186 2017
rect 1288 2003 1290 2017
rect 1384 2003 1386 2017
rect 1480 2003 1482 2017
rect 1576 2003 1578 2017
rect 1672 2003 1674 2017
rect 1752 2003 1754 2017
rect 1832 2003 1834 2035
rect 1870 2032 1871 2036
rect 1875 2032 1876 2036
rect 1870 2031 1876 2032
rect 3590 2036 3596 2037
rect 3590 2032 3591 2036
rect 3595 2032 3596 2036
rect 3590 2031 3596 2032
rect 1872 2003 1874 2031
rect 1974 2018 1980 2019
rect 1974 2014 1975 2018
rect 1979 2014 1980 2018
rect 1974 2013 1980 2014
rect 2222 2018 2228 2019
rect 2222 2014 2223 2018
rect 2227 2014 2228 2018
rect 2222 2013 2228 2014
rect 2454 2018 2460 2019
rect 2454 2014 2455 2018
rect 2459 2014 2460 2018
rect 2454 2013 2460 2014
rect 2662 2018 2668 2019
rect 2662 2014 2663 2018
rect 2667 2014 2668 2018
rect 2662 2013 2668 2014
rect 2846 2018 2852 2019
rect 2846 2014 2847 2018
rect 2851 2014 2852 2018
rect 2846 2013 2852 2014
rect 3006 2018 3012 2019
rect 3006 2014 3007 2018
rect 3011 2014 3012 2018
rect 3006 2013 3012 2014
rect 3150 2018 3156 2019
rect 3150 2014 3151 2018
rect 3155 2014 3156 2018
rect 3150 2013 3156 2014
rect 3278 2018 3284 2019
rect 3278 2014 3279 2018
rect 3283 2014 3284 2018
rect 3278 2013 3284 2014
rect 3406 2018 3412 2019
rect 3406 2014 3407 2018
rect 3411 2014 3412 2018
rect 3406 2013 3412 2014
rect 3510 2018 3516 2019
rect 3510 2014 3511 2018
rect 3515 2014 3516 2018
rect 3510 2013 3516 2014
rect 1976 2003 1978 2013
rect 2224 2003 2226 2013
rect 2456 2003 2458 2013
rect 2664 2003 2666 2013
rect 2848 2003 2850 2013
rect 3008 2003 3010 2013
rect 3152 2003 3154 2013
rect 3280 2003 3282 2013
rect 3408 2003 3410 2013
rect 3512 2003 3514 2013
rect 3592 2003 3594 2031
rect 111 2002 115 2003
rect 111 1997 115 1998
rect 191 2002 195 2003
rect 191 1997 195 1998
rect 215 2002 219 2003
rect 215 1997 219 1998
rect 335 2002 339 2003
rect 335 1997 339 1998
rect 351 2002 355 2003
rect 351 1997 355 1998
rect 455 2002 459 2003
rect 455 1997 459 1998
rect 519 2002 523 2003
rect 519 1997 523 1998
rect 583 2002 587 2003
rect 583 1997 587 1998
rect 687 2002 691 2003
rect 687 1997 691 1998
rect 711 2002 715 2003
rect 711 1997 715 1998
rect 831 2002 835 2003
rect 831 1997 835 1998
rect 855 2002 859 2003
rect 855 1997 859 1998
rect 951 2002 955 2003
rect 951 1997 955 1998
rect 1015 2002 1019 2003
rect 1015 1997 1019 1998
rect 1071 2002 1075 2003
rect 1071 1997 1075 1998
rect 1167 2002 1171 2003
rect 1167 1997 1171 1998
rect 1183 2002 1187 2003
rect 1183 1997 1187 1998
rect 1287 2002 1291 2003
rect 1287 1997 1291 1998
rect 1311 2002 1315 2003
rect 1311 1997 1315 1998
rect 1383 2002 1387 2003
rect 1383 1997 1387 1998
rect 1447 2002 1451 2003
rect 1447 1997 1451 1998
rect 1479 2002 1483 2003
rect 1479 1997 1483 1998
rect 1575 2002 1579 2003
rect 1575 1997 1579 1998
rect 1583 2002 1587 2003
rect 1583 1997 1587 1998
rect 1671 2002 1675 2003
rect 1671 1997 1675 1998
rect 1719 2002 1723 2003
rect 1719 1997 1723 1998
rect 1751 2002 1755 2003
rect 1751 1997 1755 1998
rect 1831 2002 1835 2003
rect 1831 1997 1835 1998
rect 1871 2002 1875 2003
rect 1871 1997 1875 1998
rect 1959 2002 1963 2003
rect 1959 1997 1963 1998
rect 1975 2002 1979 2003
rect 1975 1997 1979 1998
rect 2079 2002 2083 2003
rect 2079 1997 2083 1998
rect 2199 2002 2203 2003
rect 2199 1997 2203 1998
rect 2223 2002 2227 2003
rect 2223 1997 2227 1998
rect 2319 2002 2323 2003
rect 2319 1997 2323 1998
rect 2447 2002 2451 2003
rect 2447 1997 2451 1998
rect 2455 2002 2459 2003
rect 2455 1997 2459 1998
rect 2583 2002 2587 2003
rect 2583 1997 2587 1998
rect 2663 2002 2667 2003
rect 2663 1997 2667 1998
rect 2743 2002 2747 2003
rect 2743 1997 2747 1998
rect 2847 2002 2851 2003
rect 2847 1997 2851 1998
rect 2919 2002 2923 2003
rect 2919 1997 2923 1998
rect 3007 2002 3011 2003
rect 3007 1997 3011 1998
rect 3119 2002 3123 2003
rect 3119 1997 3123 1998
rect 3151 2002 3155 2003
rect 3151 1997 3155 1998
rect 3279 2002 3283 2003
rect 3279 1997 3283 1998
rect 3327 2002 3331 2003
rect 3327 1997 3331 1998
rect 3407 2002 3411 2003
rect 3407 1997 3411 1998
rect 3511 2002 3515 2003
rect 3511 1997 3515 1998
rect 3591 2002 3595 2003
rect 3591 1997 3595 1998
rect 112 1969 114 1997
rect 192 1987 194 1997
rect 352 1987 354 1997
rect 520 1987 522 1997
rect 688 1987 690 1997
rect 856 1987 858 1997
rect 1016 1987 1018 1997
rect 1168 1987 1170 1997
rect 1312 1987 1314 1997
rect 1448 1987 1450 1997
rect 1584 1987 1586 1997
rect 1720 1987 1722 1997
rect 190 1986 196 1987
rect 190 1982 191 1986
rect 195 1982 196 1986
rect 190 1981 196 1982
rect 350 1986 356 1987
rect 350 1982 351 1986
rect 355 1982 356 1986
rect 350 1981 356 1982
rect 518 1986 524 1987
rect 518 1982 519 1986
rect 523 1982 524 1986
rect 518 1981 524 1982
rect 686 1986 692 1987
rect 686 1982 687 1986
rect 691 1982 692 1986
rect 686 1981 692 1982
rect 854 1986 860 1987
rect 854 1982 855 1986
rect 859 1982 860 1986
rect 854 1981 860 1982
rect 1014 1986 1020 1987
rect 1014 1982 1015 1986
rect 1019 1982 1020 1986
rect 1014 1981 1020 1982
rect 1166 1986 1172 1987
rect 1166 1982 1167 1986
rect 1171 1982 1172 1986
rect 1166 1981 1172 1982
rect 1310 1986 1316 1987
rect 1310 1982 1311 1986
rect 1315 1982 1316 1986
rect 1310 1981 1316 1982
rect 1446 1986 1452 1987
rect 1446 1982 1447 1986
rect 1451 1982 1452 1986
rect 1446 1981 1452 1982
rect 1582 1986 1588 1987
rect 1582 1982 1583 1986
rect 1587 1982 1588 1986
rect 1582 1981 1588 1982
rect 1718 1986 1724 1987
rect 1718 1982 1719 1986
rect 1723 1982 1724 1986
rect 1718 1981 1724 1982
rect 1832 1969 1834 1997
rect 1872 1969 1874 1997
rect 1960 1987 1962 1997
rect 2080 1987 2082 1997
rect 2200 1987 2202 1997
rect 2320 1987 2322 1997
rect 2448 1987 2450 1997
rect 2584 1987 2586 1997
rect 2744 1987 2746 1997
rect 2920 1987 2922 1997
rect 3120 1987 3122 1997
rect 3328 1987 3330 1997
rect 3512 1987 3514 1997
rect 1958 1986 1964 1987
rect 1958 1982 1959 1986
rect 1963 1982 1964 1986
rect 1958 1981 1964 1982
rect 2078 1986 2084 1987
rect 2078 1982 2079 1986
rect 2083 1982 2084 1986
rect 2078 1981 2084 1982
rect 2198 1986 2204 1987
rect 2198 1982 2199 1986
rect 2203 1982 2204 1986
rect 2198 1981 2204 1982
rect 2318 1986 2324 1987
rect 2318 1982 2319 1986
rect 2323 1982 2324 1986
rect 2318 1981 2324 1982
rect 2446 1986 2452 1987
rect 2446 1982 2447 1986
rect 2451 1982 2452 1986
rect 2446 1981 2452 1982
rect 2582 1986 2588 1987
rect 2582 1982 2583 1986
rect 2587 1982 2588 1986
rect 2582 1981 2588 1982
rect 2742 1986 2748 1987
rect 2742 1982 2743 1986
rect 2747 1982 2748 1986
rect 2742 1981 2748 1982
rect 2918 1986 2924 1987
rect 2918 1982 2919 1986
rect 2923 1982 2924 1986
rect 2918 1981 2924 1982
rect 3118 1986 3124 1987
rect 3118 1982 3119 1986
rect 3123 1982 3124 1986
rect 3118 1981 3124 1982
rect 3326 1986 3332 1987
rect 3326 1982 3327 1986
rect 3331 1982 3332 1986
rect 3326 1981 3332 1982
rect 3510 1986 3516 1987
rect 3510 1982 3511 1986
rect 3515 1982 3516 1986
rect 3510 1981 3516 1982
rect 3592 1969 3594 1997
rect 110 1968 116 1969
rect 110 1964 111 1968
rect 115 1964 116 1968
rect 110 1963 116 1964
rect 1830 1968 1836 1969
rect 1830 1964 1831 1968
rect 1835 1964 1836 1968
rect 1830 1963 1836 1964
rect 1870 1968 1876 1969
rect 1870 1964 1871 1968
rect 1875 1964 1876 1968
rect 1870 1963 1876 1964
rect 3590 1968 3596 1969
rect 3590 1964 3591 1968
rect 3595 1964 3596 1968
rect 3590 1963 3596 1964
rect 110 1951 116 1952
rect 110 1947 111 1951
rect 115 1947 116 1951
rect 1830 1951 1836 1952
rect 110 1946 116 1947
rect 182 1948 188 1949
rect 112 1923 114 1946
rect 182 1944 183 1948
rect 187 1944 188 1948
rect 182 1943 188 1944
rect 342 1948 348 1949
rect 342 1944 343 1948
rect 347 1944 348 1948
rect 342 1943 348 1944
rect 510 1948 516 1949
rect 510 1944 511 1948
rect 515 1944 516 1948
rect 510 1943 516 1944
rect 678 1948 684 1949
rect 678 1944 679 1948
rect 683 1944 684 1948
rect 678 1943 684 1944
rect 846 1948 852 1949
rect 846 1944 847 1948
rect 851 1944 852 1948
rect 846 1943 852 1944
rect 1006 1948 1012 1949
rect 1006 1944 1007 1948
rect 1011 1944 1012 1948
rect 1006 1943 1012 1944
rect 1158 1948 1164 1949
rect 1158 1944 1159 1948
rect 1163 1944 1164 1948
rect 1158 1943 1164 1944
rect 1302 1948 1308 1949
rect 1302 1944 1303 1948
rect 1307 1944 1308 1948
rect 1302 1943 1308 1944
rect 1438 1948 1444 1949
rect 1438 1944 1439 1948
rect 1443 1944 1444 1948
rect 1438 1943 1444 1944
rect 1574 1948 1580 1949
rect 1574 1944 1575 1948
rect 1579 1944 1580 1948
rect 1574 1943 1580 1944
rect 1710 1948 1716 1949
rect 1710 1944 1711 1948
rect 1715 1944 1716 1948
rect 1830 1947 1831 1951
rect 1835 1947 1836 1951
rect 1830 1946 1836 1947
rect 1870 1951 1876 1952
rect 1870 1947 1871 1951
rect 1875 1947 1876 1951
rect 3590 1951 3596 1952
rect 1870 1946 1876 1947
rect 1950 1948 1956 1949
rect 1710 1943 1716 1944
rect 184 1923 186 1943
rect 344 1923 346 1943
rect 512 1923 514 1943
rect 680 1923 682 1943
rect 848 1923 850 1943
rect 1008 1923 1010 1943
rect 1160 1923 1162 1943
rect 1304 1923 1306 1943
rect 1440 1923 1442 1943
rect 1576 1923 1578 1943
rect 1712 1923 1714 1943
rect 1832 1923 1834 1946
rect 111 1922 115 1923
rect 111 1917 115 1918
rect 135 1922 139 1923
rect 135 1917 139 1918
rect 183 1922 187 1923
rect 183 1917 187 1918
rect 239 1922 243 1923
rect 239 1917 243 1918
rect 343 1922 347 1923
rect 343 1917 347 1918
rect 375 1922 379 1923
rect 375 1917 379 1918
rect 511 1922 515 1923
rect 511 1917 515 1918
rect 527 1922 531 1923
rect 527 1917 531 1918
rect 679 1922 683 1923
rect 679 1917 683 1918
rect 687 1922 691 1923
rect 687 1917 691 1918
rect 847 1922 851 1923
rect 847 1917 851 1918
rect 1007 1922 1011 1923
rect 1007 1917 1011 1918
rect 1159 1922 1163 1923
rect 1159 1917 1163 1918
rect 1303 1922 1307 1923
rect 1303 1917 1307 1918
rect 1439 1922 1443 1923
rect 1439 1917 1443 1918
rect 1455 1922 1459 1923
rect 1455 1917 1459 1918
rect 1575 1922 1579 1923
rect 1575 1917 1579 1918
rect 1607 1922 1611 1923
rect 1607 1917 1611 1918
rect 1711 1922 1715 1923
rect 1711 1917 1715 1918
rect 1831 1922 1835 1923
rect 1872 1919 1874 1946
rect 1950 1944 1951 1948
rect 1955 1944 1956 1948
rect 1950 1943 1956 1944
rect 2070 1948 2076 1949
rect 2070 1944 2071 1948
rect 2075 1944 2076 1948
rect 2070 1943 2076 1944
rect 2190 1948 2196 1949
rect 2190 1944 2191 1948
rect 2195 1944 2196 1948
rect 2190 1943 2196 1944
rect 2310 1948 2316 1949
rect 2310 1944 2311 1948
rect 2315 1944 2316 1948
rect 2310 1943 2316 1944
rect 2438 1948 2444 1949
rect 2438 1944 2439 1948
rect 2443 1944 2444 1948
rect 2438 1943 2444 1944
rect 2574 1948 2580 1949
rect 2574 1944 2575 1948
rect 2579 1944 2580 1948
rect 2574 1943 2580 1944
rect 2734 1948 2740 1949
rect 2734 1944 2735 1948
rect 2739 1944 2740 1948
rect 2734 1943 2740 1944
rect 2910 1948 2916 1949
rect 2910 1944 2911 1948
rect 2915 1944 2916 1948
rect 2910 1943 2916 1944
rect 3110 1948 3116 1949
rect 3110 1944 3111 1948
rect 3115 1944 3116 1948
rect 3110 1943 3116 1944
rect 3318 1948 3324 1949
rect 3318 1944 3319 1948
rect 3323 1944 3324 1948
rect 3318 1943 3324 1944
rect 3502 1948 3508 1949
rect 3502 1944 3503 1948
rect 3507 1944 3508 1948
rect 3590 1947 3591 1951
rect 3595 1947 3596 1951
rect 3590 1946 3596 1947
rect 3502 1943 3508 1944
rect 1952 1919 1954 1943
rect 2072 1919 2074 1943
rect 2192 1919 2194 1943
rect 2312 1919 2314 1943
rect 2440 1919 2442 1943
rect 2576 1919 2578 1943
rect 2736 1919 2738 1943
rect 2912 1919 2914 1943
rect 3112 1919 3114 1943
rect 3320 1919 3322 1943
rect 3504 1919 3506 1943
rect 3592 1919 3594 1946
rect 1831 1917 1835 1918
rect 1871 1918 1875 1919
rect 112 1898 114 1917
rect 136 1901 138 1917
rect 240 1901 242 1917
rect 376 1901 378 1917
rect 528 1901 530 1917
rect 688 1901 690 1917
rect 848 1901 850 1917
rect 1008 1901 1010 1917
rect 1160 1901 1162 1917
rect 1304 1901 1306 1917
rect 1456 1901 1458 1917
rect 1608 1901 1610 1917
rect 134 1900 140 1901
rect 110 1897 116 1898
rect 110 1893 111 1897
rect 115 1893 116 1897
rect 134 1896 135 1900
rect 139 1896 140 1900
rect 134 1895 140 1896
rect 238 1900 244 1901
rect 238 1896 239 1900
rect 243 1896 244 1900
rect 238 1895 244 1896
rect 374 1900 380 1901
rect 374 1896 375 1900
rect 379 1896 380 1900
rect 374 1895 380 1896
rect 526 1900 532 1901
rect 526 1896 527 1900
rect 531 1896 532 1900
rect 526 1895 532 1896
rect 686 1900 692 1901
rect 686 1896 687 1900
rect 691 1896 692 1900
rect 686 1895 692 1896
rect 846 1900 852 1901
rect 846 1896 847 1900
rect 851 1896 852 1900
rect 846 1895 852 1896
rect 1006 1900 1012 1901
rect 1006 1896 1007 1900
rect 1011 1896 1012 1900
rect 1006 1895 1012 1896
rect 1158 1900 1164 1901
rect 1158 1896 1159 1900
rect 1163 1896 1164 1900
rect 1158 1895 1164 1896
rect 1302 1900 1308 1901
rect 1302 1896 1303 1900
rect 1307 1896 1308 1900
rect 1302 1895 1308 1896
rect 1454 1900 1460 1901
rect 1454 1896 1455 1900
rect 1459 1896 1460 1900
rect 1454 1895 1460 1896
rect 1606 1900 1612 1901
rect 1606 1896 1607 1900
rect 1611 1896 1612 1900
rect 1832 1898 1834 1917
rect 1871 1913 1875 1914
rect 1951 1918 1955 1919
rect 1951 1913 1955 1914
rect 2063 1918 2067 1919
rect 2063 1913 2067 1914
rect 2071 1918 2075 1919
rect 2071 1913 2075 1914
rect 2151 1918 2155 1919
rect 2151 1913 2155 1914
rect 2191 1918 2195 1919
rect 2191 1913 2195 1914
rect 2239 1918 2243 1919
rect 2239 1913 2243 1914
rect 2311 1918 2315 1919
rect 2311 1913 2315 1914
rect 2319 1918 2323 1919
rect 2319 1913 2323 1914
rect 2399 1918 2403 1919
rect 2399 1913 2403 1914
rect 2439 1918 2443 1919
rect 2439 1913 2443 1914
rect 2487 1918 2491 1919
rect 2487 1913 2491 1914
rect 2575 1918 2579 1919
rect 2575 1913 2579 1914
rect 2663 1918 2667 1919
rect 2663 1913 2667 1914
rect 2735 1918 2739 1919
rect 2735 1913 2739 1914
rect 2759 1918 2763 1919
rect 2759 1913 2763 1914
rect 2871 1918 2875 1919
rect 2871 1913 2875 1914
rect 2911 1918 2915 1919
rect 2911 1913 2915 1914
rect 2991 1918 2995 1919
rect 2991 1913 2995 1914
rect 3111 1918 3115 1919
rect 3111 1913 3115 1914
rect 3119 1918 3123 1919
rect 3119 1913 3123 1914
rect 3247 1918 3251 1919
rect 3247 1913 3251 1914
rect 3319 1918 3323 1919
rect 3319 1913 3323 1914
rect 3383 1918 3387 1919
rect 3383 1913 3387 1914
rect 3503 1918 3507 1919
rect 3503 1913 3507 1914
rect 3591 1918 3595 1919
rect 3591 1913 3595 1914
rect 1606 1895 1612 1896
rect 1830 1897 1836 1898
rect 110 1892 116 1893
rect 1830 1893 1831 1897
rect 1835 1893 1836 1897
rect 1872 1894 1874 1913
rect 2064 1897 2066 1913
rect 2152 1897 2154 1913
rect 2240 1897 2242 1913
rect 2320 1897 2322 1913
rect 2400 1897 2402 1913
rect 2488 1897 2490 1913
rect 2576 1897 2578 1913
rect 2664 1897 2666 1913
rect 2760 1897 2762 1913
rect 2872 1897 2874 1913
rect 2992 1897 2994 1913
rect 3120 1897 3122 1913
rect 3248 1897 3250 1913
rect 3384 1897 3386 1913
rect 3504 1897 3506 1913
rect 2062 1896 2068 1897
rect 1830 1892 1836 1893
rect 1870 1893 1876 1894
rect 1870 1889 1871 1893
rect 1875 1889 1876 1893
rect 2062 1892 2063 1896
rect 2067 1892 2068 1896
rect 2062 1891 2068 1892
rect 2150 1896 2156 1897
rect 2150 1892 2151 1896
rect 2155 1892 2156 1896
rect 2150 1891 2156 1892
rect 2238 1896 2244 1897
rect 2238 1892 2239 1896
rect 2243 1892 2244 1896
rect 2238 1891 2244 1892
rect 2318 1896 2324 1897
rect 2318 1892 2319 1896
rect 2323 1892 2324 1896
rect 2318 1891 2324 1892
rect 2398 1896 2404 1897
rect 2398 1892 2399 1896
rect 2403 1892 2404 1896
rect 2398 1891 2404 1892
rect 2486 1896 2492 1897
rect 2486 1892 2487 1896
rect 2491 1892 2492 1896
rect 2486 1891 2492 1892
rect 2574 1896 2580 1897
rect 2574 1892 2575 1896
rect 2579 1892 2580 1896
rect 2574 1891 2580 1892
rect 2662 1896 2668 1897
rect 2662 1892 2663 1896
rect 2667 1892 2668 1896
rect 2662 1891 2668 1892
rect 2758 1896 2764 1897
rect 2758 1892 2759 1896
rect 2763 1892 2764 1896
rect 2758 1891 2764 1892
rect 2870 1896 2876 1897
rect 2870 1892 2871 1896
rect 2875 1892 2876 1896
rect 2870 1891 2876 1892
rect 2990 1896 2996 1897
rect 2990 1892 2991 1896
rect 2995 1892 2996 1896
rect 2990 1891 2996 1892
rect 3118 1896 3124 1897
rect 3118 1892 3119 1896
rect 3123 1892 3124 1896
rect 3118 1891 3124 1892
rect 3246 1896 3252 1897
rect 3246 1892 3247 1896
rect 3251 1892 3252 1896
rect 3246 1891 3252 1892
rect 3382 1896 3388 1897
rect 3382 1892 3383 1896
rect 3387 1892 3388 1896
rect 3382 1891 3388 1892
rect 3502 1896 3508 1897
rect 3502 1892 3503 1896
rect 3507 1892 3508 1896
rect 3592 1894 3594 1913
rect 3502 1891 3508 1892
rect 3590 1893 3596 1894
rect 1870 1888 1876 1889
rect 3590 1889 3591 1893
rect 3595 1889 3596 1893
rect 3590 1888 3596 1889
rect 110 1880 116 1881
rect 110 1876 111 1880
rect 115 1876 116 1880
rect 110 1875 116 1876
rect 1830 1880 1836 1881
rect 1830 1876 1831 1880
rect 1835 1876 1836 1880
rect 1830 1875 1836 1876
rect 1870 1876 1876 1877
rect 112 1843 114 1875
rect 142 1862 148 1863
rect 142 1858 143 1862
rect 147 1858 148 1862
rect 142 1857 148 1858
rect 246 1862 252 1863
rect 246 1858 247 1862
rect 251 1858 252 1862
rect 246 1857 252 1858
rect 382 1862 388 1863
rect 382 1858 383 1862
rect 387 1858 388 1862
rect 382 1857 388 1858
rect 534 1862 540 1863
rect 534 1858 535 1862
rect 539 1858 540 1862
rect 534 1857 540 1858
rect 694 1862 700 1863
rect 694 1858 695 1862
rect 699 1858 700 1862
rect 694 1857 700 1858
rect 854 1862 860 1863
rect 854 1858 855 1862
rect 859 1858 860 1862
rect 854 1857 860 1858
rect 1014 1862 1020 1863
rect 1014 1858 1015 1862
rect 1019 1858 1020 1862
rect 1014 1857 1020 1858
rect 1166 1862 1172 1863
rect 1166 1858 1167 1862
rect 1171 1858 1172 1862
rect 1166 1857 1172 1858
rect 1310 1862 1316 1863
rect 1310 1858 1311 1862
rect 1315 1858 1316 1862
rect 1310 1857 1316 1858
rect 1462 1862 1468 1863
rect 1462 1858 1463 1862
rect 1467 1858 1468 1862
rect 1462 1857 1468 1858
rect 1614 1862 1620 1863
rect 1614 1858 1615 1862
rect 1619 1858 1620 1862
rect 1614 1857 1620 1858
rect 144 1843 146 1857
rect 248 1843 250 1857
rect 384 1843 386 1857
rect 536 1843 538 1857
rect 696 1843 698 1857
rect 856 1843 858 1857
rect 1016 1843 1018 1857
rect 1168 1843 1170 1857
rect 1312 1843 1314 1857
rect 1464 1843 1466 1857
rect 1616 1843 1618 1857
rect 1832 1843 1834 1875
rect 1870 1872 1871 1876
rect 1875 1872 1876 1876
rect 1870 1871 1876 1872
rect 3590 1876 3596 1877
rect 3590 1872 3591 1876
rect 3595 1872 3596 1876
rect 3590 1871 3596 1872
rect 111 1842 115 1843
rect 111 1837 115 1838
rect 143 1842 147 1843
rect 143 1837 147 1838
rect 247 1842 251 1843
rect 247 1837 251 1838
rect 287 1842 291 1843
rect 287 1837 291 1838
rect 383 1842 387 1843
rect 383 1837 387 1838
rect 471 1842 475 1843
rect 471 1837 475 1838
rect 535 1842 539 1843
rect 535 1837 539 1838
rect 663 1842 667 1843
rect 663 1837 667 1838
rect 695 1842 699 1843
rect 695 1837 699 1838
rect 847 1842 851 1843
rect 847 1837 851 1838
rect 855 1842 859 1843
rect 855 1837 859 1838
rect 1015 1842 1019 1843
rect 1015 1837 1019 1838
rect 1023 1842 1027 1843
rect 1023 1837 1027 1838
rect 1167 1842 1171 1843
rect 1167 1837 1171 1838
rect 1191 1842 1195 1843
rect 1191 1837 1195 1838
rect 1311 1842 1315 1843
rect 1311 1837 1315 1838
rect 1351 1842 1355 1843
rect 1351 1837 1355 1838
rect 1463 1842 1467 1843
rect 1463 1837 1467 1838
rect 1511 1842 1515 1843
rect 1511 1837 1515 1838
rect 1615 1842 1619 1843
rect 1615 1837 1619 1838
rect 1679 1842 1683 1843
rect 1679 1837 1683 1838
rect 1831 1842 1835 1843
rect 1831 1837 1835 1838
rect 112 1809 114 1837
rect 144 1827 146 1837
rect 288 1827 290 1837
rect 472 1827 474 1837
rect 664 1827 666 1837
rect 848 1827 850 1837
rect 1024 1827 1026 1837
rect 1192 1827 1194 1837
rect 1352 1827 1354 1837
rect 1512 1827 1514 1837
rect 1680 1827 1682 1837
rect 142 1826 148 1827
rect 142 1822 143 1826
rect 147 1822 148 1826
rect 142 1821 148 1822
rect 286 1826 292 1827
rect 286 1822 287 1826
rect 291 1822 292 1826
rect 286 1821 292 1822
rect 470 1826 476 1827
rect 470 1822 471 1826
rect 475 1822 476 1826
rect 470 1821 476 1822
rect 662 1826 668 1827
rect 662 1822 663 1826
rect 667 1822 668 1826
rect 662 1821 668 1822
rect 846 1826 852 1827
rect 846 1822 847 1826
rect 851 1822 852 1826
rect 846 1821 852 1822
rect 1022 1826 1028 1827
rect 1022 1822 1023 1826
rect 1027 1822 1028 1826
rect 1022 1821 1028 1822
rect 1190 1826 1196 1827
rect 1190 1822 1191 1826
rect 1195 1822 1196 1826
rect 1190 1821 1196 1822
rect 1350 1826 1356 1827
rect 1350 1822 1351 1826
rect 1355 1822 1356 1826
rect 1350 1821 1356 1822
rect 1510 1826 1516 1827
rect 1510 1822 1511 1826
rect 1515 1822 1516 1826
rect 1510 1821 1516 1822
rect 1678 1826 1684 1827
rect 1678 1822 1679 1826
rect 1683 1822 1684 1826
rect 1678 1821 1684 1822
rect 1832 1809 1834 1837
rect 1872 1827 1874 1871
rect 2070 1858 2076 1859
rect 2070 1854 2071 1858
rect 2075 1854 2076 1858
rect 2070 1853 2076 1854
rect 2158 1858 2164 1859
rect 2158 1854 2159 1858
rect 2163 1854 2164 1858
rect 2158 1853 2164 1854
rect 2246 1858 2252 1859
rect 2246 1854 2247 1858
rect 2251 1854 2252 1858
rect 2246 1853 2252 1854
rect 2326 1858 2332 1859
rect 2326 1854 2327 1858
rect 2331 1854 2332 1858
rect 2326 1853 2332 1854
rect 2406 1858 2412 1859
rect 2406 1854 2407 1858
rect 2411 1854 2412 1858
rect 2406 1853 2412 1854
rect 2494 1858 2500 1859
rect 2494 1854 2495 1858
rect 2499 1854 2500 1858
rect 2494 1853 2500 1854
rect 2582 1858 2588 1859
rect 2582 1854 2583 1858
rect 2587 1854 2588 1858
rect 2582 1853 2588 1854
rect 2670 1858 2676 1859
rect 2670 1854 2671 1858
rect 2675 1854 2676 1858
rect 2670 1853 2676 1854
rect 2766 1858 2772 1859
rect 2766 1854 2767 1858
rect 2771 1854 2772 1858
rect 2766 1853 2772 1854
rect 2878 1858 2884 1859
rect 2878 1854 2879 1858
rect 2883 1854 2884 1858
rect 2878 1853 2884 1854
rect 2998 1858 3004 1859
rect 2998 1854 2999 1858
rect 3003 1854 3004 1858
rect 2998 1853 3004 1854
rect 3126 1858 3132 1859
rect 3126 1854 3127 1858
rect 3131 1854 3132 1858
rect 3126 1853 3132 1854
rect 3254 1858 3260 1859
rect 3254 1854 3255 1858
rect 3259 1854 3260 1858
rect 3254 1853 3260 1854
rect 3390 1858 3396 1859
rect 3390 1854 3391 1858
rect 3395 1854 3396 1858
rect 3390 1853 3396 1854
rect 3510 1858 3516 1859
rect 3510 1854 3511 1858
rect 3515 1854 3516 1858
rect 3510 1853 3516 1854
rect 2072 1827 2074 1853
rect 2160 1827 2162 1853
rect 2248 1827 2250 1853
rect 2328 1827 2330 1853
rect 2408 1827 2410 1853
rect 2496 1827 2498 1853
rect 2584 1827 2586 1853
rect 2672 1827 2674 1853
rect 2768 1827 2770 1853
rect 2880 1827 2882 1853
rect 3000 1827 3002 1853
rect 3128 1827 3130 1853
rect 3256 1827 3258 1853
rect 3392 1827 3394 1853
rect 3512 1827 3514 1853
rect 3592 1827 3594 1871
rect 1871 1826 1875 1827
rect 1871 1821 1875 1822
rect 2071 1826 2075 1827
rect 2071 1821 2075 1822
rect 2095 1826 2099 1827
rect 2095 1821 2099 1822
rect 2159 1826 2163 1827
rect 2159 1821 2163 1822
rect 2239 1826 2243 1827
rect 2239 1821 2243 1822
rect 2247 1826 2251 1827
rect 2247 1821 2251 1822
rect 2327 1826 2331 1827
rect 2327 1821 2331 1822
rect 2399 1826 2403 1827
rect 2399 1821 2403 1822
rect 2407 1826 2411 1827
rect 2407 1821 2411 1822
rect 2495 1826 2499 1827
rect 2495 1821 2499 1822
rect 2559 1826 2563 1827
rect 2559 1821 2563 1822
rect 2583 1826 2587 1827
rect 2583 1821 2587 1822
rect 2671 1826 2675 1827
rect 2671 1821 2675 1822
rect 2719 1826 2723 1827
rect 2719 1821 2723 1822
rect 2767 1826 2771 1827
rect 2767 1821 2771 1822
rect 2879 1826 2883 1827
rect 2879 1821 2883 1822
rect 2999 1826 3003 1827
rect 2999 1821 3003 1822
rect 3031 1826 3035 1827
rect 3031 1821 3035 1822
rect 3127 1826 3131 1827
rect 3127 1821 3131 1822
rect 3175 1826 3179 1827
rect 3175 1821 3179 1822
rect 3255 1826 3259 1827
rect 3255 1821 3259 1822
rect 3319 1826 3323 1827
rect 3319 1821 3323 1822
rect 3391 1826 3395 1827
rect 3391 1821 3395 1822
rect 3471 1826 3475 1827
rect 3471 1821 3475 1822
rect 3511 1826 3515 1827
rect 3511 1821 3515 1822
rect 3591 1826 3595 1827
rect 3591 1821 3595 1822
rect 110 1808 116 1809
rect 110 1804 111 1808
rect 115 1804 116 1808
rect 110 1803 116 1804
rect 1830 1808 1836 1809
rect 1830 1804 1831 1808
rect 1835 1804 1836 1808
rect 1830 1803 1836 1804
rect 1872 1793 1874 1821
rect 2096 1811 2098 1821
rect 2240 1811 2242 1821
rect 2400 1811 2402 1821
rect 2560 1811 2562 1821
rect 2720 1811 2722 1821
rect 2880 1811 2882 1821
rect 3032 1811 3034 1821
rect 3176 1811 3178 1821
rect 3320 1811 3322 1821
rect 3472 1811 3474 1821
rect 2094 1810 2100 1811
rect 2094 1806 2095 1810
rect 2099 1806 2100 1810
rect 2094 1805 2100 1806
rect 2238 1810 2244 1811
rect 2238 1806 2239 1810
rect 2243 1806 2244 1810
rect 2238 1805 2244 1806
rect 2398 1810 2404 1811
rect 2398 1806 2399 1810
rect 2403 1806 2404 1810
rect 2398 1805 2404 1806
rect 2558 1810 2564 1811
rect 2558 1806 2559 1810
rect 2563 1806 2564 1810
rect 2558 1805 2564 1806
rect 2718 1810 2724 1811
rect 2718 1806 2719 1810
rect 2723 1806 2724 1810
rect 2718 1805 2724 1806
rect 2878 1810 2884 1811
rect 2878 1806 2879 1810
rect 2883 1806 2884 1810
rect 2878 1805 2884 1806
rect 3030 1810 3036 1811
rect 3030 1806 3031 1810
rect 3035 1806 3036 1810
rect 3030 1805 3036 1806
rect 3174 1810 3180 1811
rect 3174 1806 3175 1810
rect 3179 1806 3180 1810
rect 3174 1805 3180 1806
rect 3318 1810 3324 1811
rect 3318 1806 3319 1810
rect 3323 1806 3324 1810
rect 3318 1805 3324 1806
rect 3470 1810 3476 1811
rect 3470 1806 3471 1810
rect 3475 1806 3476 1810
rect 3470 1805 3476 1806
rect 3592 1793 3594 1821
rect 1870 1792 1876 1793
rect 110 1791 116 1792
rect 110 1787 111 1791
rect 115 1787 116 1791
rect 1830 1791 1836 1792
rect 110 1786 116 1787
rect 134 1788 140 1789
rect 112 1759 114 1786
rect 134 1784 135 1788
rect 139 1784 140 1788
rect 134 1783 140 1784
rect 278 1788 284 1789
rect 278 1784 279 1788
rect 283 1784 284 1788
rect 278 1783 284 1784
rect 462 1788 468 1789
rect 462 1784 463 1788
rect 467 1784 468 1788
rect 462 1783 468 1784
rect 654 1788 660 1789
rect 654 1784 655 1788
rect 659 1784 660 1788
rect 654 1783 660 1784
rect 838 1788 844 1789
rect 838 1784 839 1788
rect 843 1784 844 1788
rect 838 1783 844 1784
rect 1014 1788 1020 1789
rect 1014 1784 1015 1788
rect 1019 1784 1020 1788
rect 1014 1783 1020 1784
rect 1182 1788 1188 1789
rect 1182 1784 1183 1788
rect 1187 1784 1188 1788
rect 1182 1783 1188 1784
rect 1342 1788 1348 1789
rect 1342 1784 1343 1788
rect 1347 1784 1348 1788
rect 1342 1783 1348 1784
rect 1502 1788 1508 1789
rect 1502 1784 1503 1788
rect 1507 1784 1508 1788
rect 1502 1783 1508 1784
rect 1670 1788 1676 1789
rect 1670 1784 1671 1788
rect 1675 1784 1676 1788
rect 1830 1787 1831 1791
rect 1835 1787 1836 1791
rect 1870 1788 1871 1792
rect 1875 1788 1876 1792
rect 1870 1787 1876 1788
rect 3590 1792 3596 1793
rect 3590 1788 3591 1792
rect 3595 1788 3596 1792
rect 3590 1787 3596 1788
rect 1830 1786 1836 1787
rect 1670 1783 1676 1784
rect 136 1759 138 1783
rect 280 1759 282 1783
rect 464 1759 466 1783
rect 656 1759 658 1783
rect 840 1759 842 1783
rect 1016 1759 1018 1783
rect 1184 1759 1186 1783
rect 1344 1759 1346 1783
rect 1504 1759 1506 1783
rect 1672 1759 1674 1783
rect 1832 1759 1834 1786
rect 1870 1775 1876 1776
rect 1870 1771 1871 1775
rect 1875 1771 1876 1775
rect 3590 1775 3596 1776
rect 1870 1770 1876 1771
rect 2086 1772 2092 1773
rect 111 1758 115 1759
rect 111 1753 115 1754
rect 135 1758 139 1759
rect 135 1753 139 1754
rect 215 1758 219 1759
rect 215 1753 219 1754
rect 279 1758 283 1759
rect 279 1753 283 1754
rect 343 1758 347 1759
rect 343 1753 347 1754
rect 463 1758 467 1759
rect 463 1753 467 1754
rect 495 1758 499 1759
rect 495 1753 499 1754
rect 655 1758 659 1759
rect 655 1753 659 1754
rect 663 1758 667 1759
rect 663 1753 667 1754
rect 839 1758 843 1759
rect 839 1753 843 1754
rect 1007 1758 1011 1759
rect 1007 1753 1011 1754
rect 1015 1758 1019 1759
rect 1015 1753 1019 1754
rect 1167 1758 1171 1759
rect 1167 1753 1171 1754
rect 1183 1758 1187 1759
rect 1183 1753 1187 1754
rect 1319 1758 1323 1759
rect 1319 1753 1323 1754
rect 1343 1758 1347 1759
rect 1343 1753 1347 1754
rect 1463 1758 1467 1759
rect 1463 1753 1467 1754
rect 1503 1758 1507 1759
rect 1503 1753 1507 1754
rect 1607 1758 1611 1759
rect 1607 1753 1611 1754
rect 1671 1758 1675 1759
rect 1671 1753 1675 1754
rect 1743 1758 1747 1759
rect 1743 1753 1747 1754
rect 1831 1758 1835 1759
rect 1831 1753 1835 1754
rect 112 1734 114 1753
rect 136 1737 138 1753
rect 216 1737 218 1753
rect 344 1737 346 1753
rect 496 1737 498 1753
rect 664 1737 666 1753
rect 840 1737 842 1753
rect 1008 1737 1010 1753
rect 1168 1737 1170 1753
rect 1320 1737 1322 1753
rect 1464 1737 1466 1753
rect 1608 1737 1610 1753
rect 1744 1737 1746 1753
rect 134 1736 140 1737
rect 110 1733 116 1734
rect 110 1729 111 1733
rect 115 1729 116 1733
rect 134 1732 135 1736
rect 139 1732 140 1736
rect 134 1731 140 1732
rect 214 1736 220 1737
rect 214 1732 215 1736
rect 219 1732 220 1736
rect 214 1731 220 1732
rect 342 1736 348 1737
rect 342 1732 343 1736
rect 347 1732 348 1736
rect 342 1731 348 1732
rect 494 1736 500 1737
rect 494 1732 495 1736
rect 499 1732 500 1736
rect 494 1731 500 1732
rect 662 1736 668 1737
rect 662 1732 663 1736
rect 667 1732 668 1736
rect 662 1731 668 1732
rect 838 1736 844 1737
rect 838 1732 839 1736
rect 843 1732 844 1736
rect 838 1731 844 1732
rect 1006 1736 1012 1737
rect 1006 1732 1007 1736
rect 1011 1732 1012 1736
rect 1006 1731 1012 1732
rect 1166 1736 1172 1737
rect 1166 1732 1167 1736
rect 1171 1732 1172 1736
rect 1166 1731 1172 1732
rect 1318 1736 1324 1737
rect 1318 1732 1319 1736
rect 1323 1732 1324 1736
rect 1318 1731 1324 1732
rect 1462 1736 1468 1737
rect 1462 1732 1463 1736
rect 1467 1732 1468 1736
rect 1462 1731 1468 1732
rect 1606 1736 1612 1737
rect 1606 1732 1607 1736
rect 1611 1732 1612 1736
rect 1606 1731 1612 1732
rect 1742 1736 1748 1737
rect 1742 1732 1743 1736
rect 1747 1732 1748 1736
rect 1832 1734 1834 1753
rect 1872 1747 1874 1770
rect 2086 1768 2087 1772
rect 2091 1768 2092 1772
rect 2086 1767 2092 1768
rect 2230 1772 2236 1773
rect 2230 1768 2231 1772
rect 2235 1768 2236 1772
rect 2230 1767 2236 1768
rect 2390 1772 2396 1773
rect 2390 1768 2391 1772
rect 2395 1768 2396 1772
rect 2390 1767 2396 1768
rect 2550 1772 2556 1773
rect 2550 1768 2551 1772
rect 2555 1768 2556 1772
rect 2550 1767 2556 1768
rect 2710 1772 2716 1773
rect 2710 1768 2711 1772
rect 2715 1768 2716 1772
rect 2710 1767 2716 1768
rect 2870 1772 2876 1773
rect 2870 1768 2871 1772
rect 2875 1768 2876 1772
rect 2870 1767 2876 1768
rect 3022 1772 3028 1773
rect 3022 1768 3023 1772
rect 3027 1768 3028 1772
rect 3022 1767 3028 1768
rect 3166 1772 3172 1773
rect 3166 1768 3167 1772
rect 3171 1768 3172 1772
rect 3166 1767 3172 1768
rect 3310 1772 3316 1773
rect 3310 1768 3311 1772
rect 3315 1768 3316 1772
rect 3310 1767 3316 1768
rect 3462 1772 3468 1773
rect 3462 1768 3463 1772
rect 3467 1768 3468 1772
rect 3590 1771 3591 1775
rect 3595 1771 3596 1775
rect 3590 1770 3596 1771
rect 3462 1767 3468 1768
rect 2088 1747 2090 1767
rect 2232 1747 2234 1767
rect 2392 1747 2394 1767
rect 2552 1747 2554 1767
rect 2712 1747 2714 1767
rect 2872 1747 2874 1767
rect 3024 1747 3026 1767
rect 3168 1747 3170 1767
rect 3312 1747 3314 1767
rect 3464 1747 3466 1767
rect 3592 1747 3594 1770
rect 1871 1746 1875 1747
rect 1871 1741 1875 1742
rect 2087 1746 2091 1747
rect 2087 1741 2091 1742
rect 2103 1746 2107 1747
rect 2103 1741 2107 1742
rect 2231 1746 2235 1747
rect 2231 1741 2235 1742
rect 2239 1746 2243 1747
rect 2239 1741 2243 1742
rect 2383 1746 2387 1747
rect 2383 1741 2387 1742
rect 2391 1746 2395 1747
rect 2391 1741 2395 1742
rect 2527 1746 2531 1747
rect 2527 1741 2531 1742
rect 2551 1746 2555 1747
rect 2551 1741 2555 1742
rect 2663 1746 2667 1747
rect 2663 1741 2667 1742
rect 2711 1746 2715 1747
rect 2711 1741 2715 1742
rect 2799 1746 2803 1747
rect 2799 1741 2803 1742
rect 2871 1746 2875 1747
rect 2871 1741 2875 1742
rect 2927 1746 2931 1747
rect 2927 1741 2931 1742
rect 3023 1746 3027 1747
rect 3023 1741 3027 1742
rect 3047 1746 3051 1747
rect 3047 1741 3051 1742
rect 3159 1746 3163 1747
rect 3159 1741 3163 1742
rect 3167 1746 3171 1747
rect 3167 1741 3171 1742
rect 3271 1746 3275 1747
rect 3271 1741 3275 1742
rect 3311 1746 3315 1747
rect 3311 1741 3315 1742
rect 3391 1746 3395 1747
rect 3391 1741 3395 1742
rect 3463 1746 3467 1747
rect 3463 1741 3467 1742
rect 3503 1746 3507 1747
rect 3503 1741 3507 1742
rect 3591 1746 3595 1747
rect 3591 1741 3595 1742
rect 1742 1731 1748 1732
rect 1830 1733 1836 1734
rect 110 1728 116 1729
rect 1830 1729 1831 1733
rect 1835 1729 1836 1733
rect 1830 1728 1836 1729
rect 1872 1722 1874 1741
rect 2104 1725 2106 1741
rect 2240 1725 2242 1741
rect 2384 1725 2386 1741
rect 2528 1725 2530 1741
rect 2664 1725 2666 1741
rect 2800 1725 2802 1741
rect 2928 1725 2930 1741
rect 3048 1725 3050 1741
rect 3160 1725 3162 1741
rect 3272 1725 3274 1741
rect 3392 1725 3394 1741
rect 3504 1725 3506 1741
rect 2102 1724 2108 1725
rect 1870 1721 1876 1722
rect 1870 1717 1871 1721
rect 1875 1717 1876 1721
rect 2102 1720 2103 1724
rect 2107 1720 2108 1724
rect 2102 1719 2108 1720
rect 2238 1724 2244 1725
rect 2238 1720 2239 1724
rect 2243 1720 2244 1724
rect 2238 1719 2244 1720
rect 2382 1724 2388 1725
rect 2382 1720 2383 1724
rect 2387 1720 2388 1724
rect 2382 1719 2388 1720
rect 2526 1724 2532 1725
rect 2526 1720 2527 1724
rect 2531 1720 2532 1724
rect 2526 1719 2532 1720
rect 2662 1724 2668 1725
rect 2662 1720 2663 1724
rect 2667 1720 2668 1724
rect 2662 1719 2668 1720
rect 2798 1724 2804 1725
rect 2798 1720 2799 1724
rect 2803 1720 2804 1724
rect 2798 1719 2804 1720
rect 2926 1724 2932 1725
rect 2926 1720 2927 1724
rect 2931 1720 2932 1724
rect 2926 1719 2932 1720
rect 3046 1724 3052 1725
rect 3046 1720 3047 1724
rect 3051 1720 3052 1724
rect 3046 1719 3052 1720
rect 3158 1724 3164 1725
rect 3158 1720 3159 1724
rect 3163 1720 3164 1724
rect 3158 1719 3164 1720
rect 3270 1724 3276 1725
rect 3270 1720 3271 1724
rect 3275 1720 3276 1724
rect 3270 1719 3276 1720
rect 3390 1724 3396 1725
rect 3390 1720 3391 1724
rect 3395 1720 3396 1724
rect 3390 1719 3396 1720
rect 3502 1724 3508 1725
rect 3502 1720 3503 1724
rect 3507 1720 3508 1724
rect 3592 1722 3594 1741
rect 3502 1719 3508 1720
rect 3590 1721 3596 1722
rect 110 1716 116 1717
rect 110 1712 111 1716
rect 115 1712 116 1716
rect 110 1711 116 1712
rect 1830 1716 1836 1717
rect 1870 1716 1876 1717
rect 3590 1717 3591 1721
rect 3595 1717 3596 1721
rect 3590 1716 3596 1717
rect 1830 1712 1831 1716
rect 1835 1712 1836 1716
rect 1830 1711 1836 1712
rect 112 1679 114 1711
rect 142 1698 148 1699
rect 142 1694 143 1698
rect 147 1694 148 1698
rect 142 1693 148 1694
rect 222 1698 228 1699
rect 222 1694 223 1698
rect 227 1694 228 1698
rect 222 1693 228 1694
rect 350 1698 356 1699
rect 350 1694 351 1698
rect 355 1694 356 1698
rect 350 1693 356 1694
rect 502 1698 508 1699
rect 502 1694 503 1698
rect 507 1694 508 1698
rect 502 1693 508 1694
rect 670 1698 676 1699
rect 670 1694 671 1698
rect 675 1694 676 1698
rect 670 1693 676 1694
rect 846 1698 852 1699
rect 846 1694 847 1698
rect 851 1694 852 1698
rect 846 1693 852 1694
rect 1014 1698 1020 1699
rect 1014 1694 1015 1698
rect 1019 1694 1020 1698
rect 1014 1693 1020 1694
rect 1174 1698 1180 1699
rect 1174 1694 1175 1698
rect 1179 1694 1180 1698
rect 1174 1693 1180 1694
rect 1326 1698 1332 1699
rect 1326 1694 1327 1698
rect 1331 1694 1332 1698
rect 1326 1693 1332 1694
rect 1470 1698 1476 1699
rect 1470 1694 1471 1698
rect 1475 1694 1476 1698
rect 1470 1693 1476 1694
rect 1614 1698 1620 1699
rect 1614 1694 1615 1698
rect 1619 1694 1620 1698
rect 1614 1693 1620 1694
rect 1750 1698 1756 1699
rect 1750 1694 1751 1698
rect 1755 1694 1756 1698
rect 1750 1693 1756 1694
rect 144 1679 146 1693
rect 224 1679 226 1693
rect 352 1679 354 1693
rect 504 1679 506 1693
rect 672 1679 674 1693
rect 848 1679 850 1693
rect 1016 1679 1018 1693
rect 1176 1679 1178 1693
rect 1328 1679 1330 1693
rect 1472 1679 1474 1693
rect 1616 1679 1618 1693
rect 1752 1679 1754 1693
rect 1832 1679 1834 1711
rect 1870 1704 1876 1705
rect 1870 1700 1871 1704
rect 1875 1700 1876 1704
rect 1870 1699 1876 1700
rect 3590 1704 3596 1705
rect 3590 1700 3591 1704
rect 3595 1700 3596 1704
rect 3590 1699 3596 1700
rect 111 1678 115 1679
rect 111 1673 115 1674
rect 143 1678 147 1679
rect 143 1673 147 1674
rect 223 1678 227 1679
rect 223 1673 227 1674
rect 295 1678 299 1679
rect 295 1673 299 1674
rect 351 1678 355 1679
rect 351 1673 355 1674
rect 479 1678 483 1679
rect 479 1673 483 1674
rect 503 1678 507 1679
rect 503 1673 507 1674
rect 671 1678 675 1679
rect 671 1673 675 1674
rect 847 1678 851 1679
rect 847 1673 851 1674
rect 855 1678 859 1679
rect 855 1673 859 1674
rect 1015 1678 1019 1679
rect 1015 1673 1019 1674
rect 1031 1678 1035 1679
rect 1031 1673 1035 1674
rect 1175 1678 1179 1679
rect 1175 1673 1179 1674
rect 1199 1678 1203 1679
rect 1199 1673 1203 1674
rect 1327 1678 1331 1679
rect 1327 1673 1331 1674
rect 1359 1678 1363 1679
rect 1359 1673 1363 1674
rect 1471 1678 1475 1679
rect 1471 1673 1475 1674
rect 1519 1678 1523 1679
rect 1519 1673 1523 1674
rect 1615 1678 1619 1679
rect 1615 1673 1619 1674
rect 1679 1678 1683 1679
rect 1679 1673 1683 1674
rect 1751 1678 1755 1679
rect 1751 1673 1755 1674
rect 1831 1678 1835 1679
rect 1831 1673 1835 1674
rect 112 1645 114 1673
rect 144 1663 146 1673
rect 296 1663 298 1673
rect 480 1663 482 1673
rect 672 1663 674 1673
rect 856 1663 858 1673
rect 1032 1663 1034 1673
rect 1200 1663 1202 1673
rect 1360 1663 1362 1673
rect 1520 1663 1522 1673
rect 1680 1663 1682 1673
rect 142 1662 148 1663
rect 142 1658 143 1662
rect 147 1658 148 1662
rect 142 1657 148 1658
rect 294 1662 300 1663
rect 294 1658 295 1662
rect 299 1658 300 1662
rect 294 1657 300 1658
rect 478 1662 484 1663
rect 478 1658 479 1662
rect 483 1658 484 1662
rect 478 1657 484 1658
rect 670 1662 676 1663
rect 670 1658 671 1662
rect 675 1658 676 1662
rect 670 1657 676 1658
rect 854 1662 860 1663
rect 854 1658 855 1662
rect 859 1658 860 1662
rect 854 1657 860 1658
rect 1030 1662 1036 1663
rect 1030 1658 1031 1662
rect 1035 1658 1036 1662
rect 1030 1657 1036 1658
rect 1198 1662 1204 1663
rect 1198 1658 1199 1662
rect 1203 1658 1204 1662
rect 1198 1657 1204 1658
rect 1358 1662 1364 1663
rect 1358 1658 1359 1662
rect 1363 1658 1364 1662
rect 1358 1657 1364 1658
rect 1518 1662 1524 1663
rect 1518 1658 1519 1662
rect 1523 1658 1524 1662
rect 1518 1657 1524 1658
rect 1678 1662 1684 1663
rect 1678 1658 1679 1662
rect 1683 1658 1684 1662
rect 1678 1657 1684 1658
rect 1832 1645 1834 1673
rect 1872 1667 1874 1699
rect 2110 1686 2116 1687
rect 2110 1682 2111 1686
rect 2115 1682 2116 1686
rect 2110 1681 2116 1682
rect 2246 1686 2252 1687
rect 2246 1682 2247 1686
rect 2251 1682 2252 1686
rect 2246 1681 2252 1682
rect 2390 1686 2396 1687
rect 2390 1682 2391 1686
rect 2395 1682 2396 1686
rect 2390 1681 2396 1682
rect 2534 1686 2540 1687
rect 2534 1682 2535 1686
rect 2539 1682 2540 1686
rect 2534 1681 2540 1682
rect 2670 1686 2676 1687
rect 2670 1682 2671 1686
rect 2675 1682 2676 1686
rect 2670 1681 2676 1682
rect 2806 1686 2812 1687
rect 2806 1682 2807 1686
rect 2811 1682 2812 1686
rect 2806 1681 2812 1682
rect 2934 1686 2940 1687
rect 2934 1682 2935 1686
rect 2939 1682 2940 1686
rect 2934 1681 2940 1682
rect 3054 1686 3060 1687
rect 3054 1682 3055 1686
rect 3059 1682 3060 1686
rect 3054 1681 3060 1682
rect 3166 1686 3172 1687
rect 3166 1682 3167 1686
rect 3171 1682 3172 1686
rect 3166 1681 3172 1682
rect 3278 1686 3284 1687
rect 3278 1682 3279 1686
rect 3283 1682 3284 1686
rect 3278 1681 3284 1682
rect 3398 1686 3404 1687
rect 3398 1682 3399 1686
rect 3403 1682 3404 1686
rect 3398 1681 3404 1682
rect 3510 1686 3516 1687
rect 3510 1682 3511 1686
rect 3515 1682 3516 1686
rect 3510 1681 3516 1682
rect 2112 1667 2114 1681
rect 2248 1667 2250 1681
rect 2392 1667 2394 1681
rect 2536 1667 2538 1681
rect 2672 1667 2674 1681
rect 2808 1667 2810 1681
rect 2936 1667 2938 1681
rect 3056 1667 3058 1681
rect 3168 1667 3170 1681
rect 3280 1667 3282 1681
rect 3400 1667 3402 1681
rect 3512 1667 3514 1681
rect 3592 1667 3594 1699
rect 1871 1666 1875 1667
rect 1871 1661 1875 1662
rect 1967 1666 1971 1667
rect 1967 1661 1971 1662
rect 2087 1666 2091 1667
rect 2087 1661 2091 1662
rect 2111 1666 2115 1667
rect 2111 1661 2115 1662
rect 2215 1666 2219 1667
rect 2215 1661 2219 1662
rect 2247 1666 2251 1667
rect 2247 1661 2251 1662
rect 2351 1666 2355 1667
rect 2351 1661 2355 1662
rect 2391 1666 2395 1667
rect 2391 1661 2395 1662
rect 2495 1666 2499 1667
rect 2495 1661 2499 1662
rect 2535 1666 2539 1667
rect 2535 1661 2539 1662
rect 2639 1666 2643 1667
rect 2639 1661 2643 1662
rect 2671 1666 2675 1667
rect 2671 1661 2675 1662
rect 2783 1666 2787 1667
rect 2783 1661 2787 1662
rect 2807 1666 2811 1667
rect 2807 1661 2811 1662
rect 2927 1666 2931 1667
rect 2927 1661 2931 1662
rect 2935 1666 2939 1667
rect 2935 1661 2939 1662
rect 3055 1666 3059 1667
rect 3055 1661 3059 1662
rect 3071 1666 3075 1667
rect 3071 1661 3075 1662
rect 3167 1666 3171 1667
rect 3167 1661 3171 1662
rect 3223 1666 3227 1667
rect 3223 1661 3227 1662
rect 3279 1666 3283 1667
rect 3279 1661 3283 1662
rect 3375 1666 3379 1667
rect 3375 1661 3379 1662
rect 3399 1666 3403 1667
rect 3399 1661 3403 1662
rect 3511 1666 3515 1667
rect 3511 1661 3515 1662
rect 3591 1666 3595 1667
rect 3591 1661 3595 1662
rect 110 1644 116 1645
rect 110 1640 111 1644
rect 115 1640 116 1644
rect 110 1639 116 1640
rect 1830 1644 1836 1645
rect 1830 1640 1831 1644
rect 1835 1640 1836 1644
rect 1830 1639 1836 1640
rect 1872 1633 1874 1661
rect 1968 1651 1970 1661
rect 2088 1651 2090 1661
rect 2216 1651 2218 1661
rect 2352 1651 2354 1661
rect 2496 1651 2498 1661
rect 2640 1651 2642 1661
rect 2784 1651 2786 1661
rect 2928 1651 2930 1661
rect 3072 1651 3074 1661
rect 3224 1651 3226 1661
rect 3376 1651 3378 1661
rect 3512 1651 3514 1661
rect 1966 1650 1972 1651
rect 1966 1646 1967 1650
rect 1971 1646 1972 1650
rect 1966 1645 1972 1646
rect 2086 1650 2092 1651
rect 2086 1646 2087 1650
rect 2091 1646 2092 1650
rect 2086 1645 2092 1646
rect 2214 1650 2220 1651
rect 2214 1646 2215 1650
rect 2219 1646 2220 1650
rect 2214 1645 2220 1646
rect 2350 1650 2356 1651
rect 2350 1646 2351 1650
rect 2355 1646 2356 1650
rect 2350 1645 2356 1646
rect 2494 1650 2500 1651
rect 2494 1646 2495 1650
rect 2499 1646 2500 1650
rect 2494 1645 2500 1646
rect 2638 1650 2644 1651
rect 2638 1646 2639 1650
rect 2643 1646 2644 1650
rect 2638 1645 2644 1646
rect 2782 1650 2788 1651
rect 2782 1646 2783 1650
rect 2787 1646 2788 1650
rect 2782 1645 2788 1646
rect 2926 1650 2932 1651
rect 2926 1646 2927 1650
rect 2931 1646 2932 1650
rect 2926 1645 2932 1646
rect 3070 1650 3076 1651
rect 3070 1646 3071 1650
rect 3075 1646 3076 1650
rect 3070 1645 3076 1646
rect 3222 1650 3228 1651
rect 3222 1646 3223 1650
rect 3227 1646 3228 1650
rect 3222 1645 3228 1646
rect 3374 1650 3380 1651
rect 3374 1646 3375 1650
rect 3379 1646 3380 1650
rect 3374 1645 3380 1646
rect 3510 1650 3516 1651
rect 3510 1646 3511 1650
rect 3515 1646 3516 1650
rect 3510 1645 3516 1646
rect 3592 1633 3594 1661
rect 1870 1632 1876 1633
rect 1870 1628 1871 1632
rect 1875 1628 1876 1632
rect 110 1627 116 1628
rect 110 1623 111 1627
rect 115 1623 116 1627
rect 1830 1627 1836 1628
rect 1870 1627 1876 1628
rect 3590 1632 3596 1633
rect 3590 1628 3591 1632
rect 3595 1628 3596 1632
rect 3590 1627 3596 1628
rect 110 1622 116 1623
rect 134 1624 140 1625
rect 112 1603 114 1622
rect 134 1620 135 1624
rect 139 1620 140 1624
rect 134 1619 140 1620
rect 286 1624 292 1625
rect 286 1620 287 1624
rect 291 1620 292 1624
rect 286 1619 292 1620
rect 470 1624 476 1625
rect 470 1620 471 1624
rect 475 1620 476 1624
rect 470 1619 476 1620
rect 662 1624 668 1625
rect 662 1620 663 1624
rect 667 1620 668 1624
rect 662 1619 668 1620
rect 846 1624 852 1625
rect 846 1620 847 1624
rect 851 1620 852 1624
rect 846 1619 852 1620
rect 1022 1624 1028 1625
rect 1022 1620 1023 1624
rect 1027 1620 1028 1624
rect 1022 1619 1028 1620
rect 1190 1624 1196 1625
rect 1190 1620 1191 1624
rect 1195 1620 1196 1624
rect 1190 1619 1196 1620
rect 1350 1624 1356 1625
rect 1350 1620 1351 1624
rect 1355 1620 1356 1624
rect 1350 1619 1356 1620
rect 1510 1624 1516 1625
rect 1510 1620 1511 1624
rect 1515 1620 1516 1624
rect 1510 1619 1516 1620
rect 1670 1624 1676 1625
rect 1670 1620 1671 1624
rect 1675 1620 1676 1624
rect 1830 1623 1831 1627
rect 1835 1623 1836 1627
rect 1830 1622 1836 1623
rect 1670 1619 1676 1620
rect 136 1603 138 1619
rect 288 1603 290 1619
rect 472 1603 474 1619
rect 664 1603 666 1619
rect 848 1603 850 1619
rect 1024 1603 1026 1619
rect 1192 1603 1194 1619
rect 1352 1603 1354 1619
rect 1512 1603 1514 1619
rect 1672 1603 1674 1619
rect 1832 1603 1834 1622
rect 1870 1615 1876 1616
rect 1870 1611 1871 1615
rect 1875 1611 1876 1615
rect 3590 1615 3596 1616
rect 1870 1610 1876 1611
rect 1958 1612 1964 1613
rect 111 1602 115 1603
rect 111 1597 115 1598
rect 135 1602 139 1603
rect 135 1597 139 1598
rect 159 1602 163 1603
rect 159 1597 163 1598
rect 287 1602 291 1603
rect 287 1597 291 1598
rect 423 1602 427 1603
rect 423 1597 427 1598
rect 471 1602 475 1603
rect 471 1597 475 1598
rect 567 1602 571 1603
rect 567 1597 571 1598
rect 663 1602 667 1603
rect 663 1597 667 1598
rect 711 1602 715 1603
rect 711 1597 715 1598
rect 847 1602 851 1603
rect 847 1597 851 1598
rect 983 1602 987 1603
rect 983 1597 987 1598
rect 1023 1602 1027 1603
rect 1023 1597 1027 1598
rect 1119 1602 1123 1603
rect 1119 1597 1123 1598
rect 1191 1602 1195 1603
rect 1191 1597 1195 1598
rect 1247 1602 1251 1603
rect 1247 1597 1251 1598
rect 1351 1602 1355 1603
rect 1351 1597 1355 1598
rect 1375 1602 1379 1603
rect 1375 1597 1379 1598
rect 1511 1602 1515 1603
rect 1511 1597 1515 1598
rect 1671 1602 1675 1603
rect 1671 1597 1675 1598
rect 1831 1602 1835 1603
rect 1831 1597 1835 1598
rect 112 1578 114 1597
rect 160 1581 162 1597
rect 288 1581 290 1597
rect 424 1581 426 1597
rect 568 1581 570 1597
rect 712 1581 714 1597
rect 848 1581 850 1597
rect 984 1581 986 1597
rect 1120 1581 1122 1597
rect 1248 1581 1250 1597
rect 1376 1581 1378 1597
rect 1512 1581 1514 1597
rect 158 1580 164 1581
rect 110 1577 116 1578
rect 110 1573 111 1577
rect 115 1573 116 1577
rect 158 1576 159 1580
rect 163 1576 164 1580
rect 158 1575 164 1576
rect 286 1580 292 1581
rect 286 1576 287 1580
rect 291 1576 292 1580
rect 286 1575 292 1576
rect 422 1580 428 1581
rect 422 1576 423 1580
rect 427 1576 428 1580
rect 422 1575 428 1576
rect 566 1580 572 1581
rect 566 1576 567 1580
rect 571 1576 572 1580
rect 566 1575 572 1576
rect 710 1580 716 1581
rect 710 1576 711 1580
rect 715 1576 716 1580
rect 710 1575 716 1576
rect 846 1580 852 1581
rect 846 1576 847 1580
rect 851 1576 852 1580
rect 846 1575 852 1576
rect 982 1580 988 1581
rect 982 1576 983 1580
rect 987 1576 988 1580
rect 982 1575 988 1576
rect 1118 1580 1124 1581
rect 1118 1576 1119 1580
rect 1123 1576 1124 1580
rect 1118 1575 1124 1576
rect 1246 1580 1252 1581
rect 1246 1576 1247 1580
rect 1251 1576 1252 1580
rect 1246 1575 1252 1576
rect 1374 1580 1380 1581
rect 1374 1576 1375 1580
rect 1379 1576 1380 1580
rect 1374 1575 1380 1576
rect 1510 1580 1516 1581
rect 1510 1576 1511 1580
rect 1515 1576 1516 1580
rect 1832 1578 1834 1597
rect 1872 1583 1874 1610
rect 1958 1608 1959 1612
rect 1963 1608 1964 1612
rect 1958 1607 1964 1608
rect 2078 1612 2084 1613
rect 2078 1608 2079 1612
rect 2083 1608 2084 1612
rect 2078 1607 2084 1608
rect 2206 1612 2212 1613
rect 2206 1608 2207 1612
rect 2211 1608 2212 1612
rect 2206 1607 2212 1608
rect 2342 1612 2348 1613
rect 2342 1608 2343 1612
rect 2347 1608 2348 1612
rect 2342 1607 2348 1608
rect 2486 1612 2492 1613
rect 2486 1608 2487 1612
rect 2491 1608 2492 1612
rect 2486 1607 2492 1608
rect 2630 1612 2636 1613
rect 2630 1608 2631 1612
rect 2635 1608 2636 1612
rect 2630 1607 2636 1608
rect 2774 1612 2780 1613
rect 2774 1608 2775 1612
rect 2779 1608 2780 1612
rect 2774 1607 2780 1608
rect 2918 1612 2924 1613
rect 2918 1608 2919 1612
rect 2923 1608 2924 1612
rect 2918 1607 2924 1608
rect 3062 1612 3068 1613
rect 3062 1608 3063 1612
rect 3067 1608 3068 1612
rect 3062 1607 3068 1608
rect 3214 1612 3220 1613
rect 3214 1608 3215 1612
rect 3219 1608 3220 1612
rect 3214 1607 3220 1608
rect 3366 1612 3372 1613
rect 3366 1608 3367 1612
rect 3371 1608 3372 1612
rect 3366 1607 3372 1608
rect 3502 1612 3508 1613
rect 3502 1608 3503 1612
rect 3507 1608 3508 1612
rect 3590 1611 3591 1615
rect 3595 1611 3596 1615
rect 3590 1610 3596 1611
rect 3502 1607 3508 1608
rect 1960 1583 1962 1607
rect 2080 1583 2082 1607
rect 2208 1583 2210 1607
rect 2344 1583 2346 1607
rect 2488 1583 2490 1607
rect 2632 1583 2634 1607
rect 2776 1583 2778 1607
rect 2920 1583 2922 1607
rect 3064 1583 3066 1607
rect 3216 1583 3218 1607
rect 3368 1583 3370 1607
rect 3504 1583 3506 1607
rect 3592 1583 3594 1610
rect 1871 1582 1875 1583
rect 1510 1575 1516 1576
rect 1830 1577 1836 1578
rect 1871 1577 1875 1578
rect 1895 1582 1899 1583
rect 1895 1577 1899 1578
rect 1959 1582 1963 1583
rect 1959 1577 1963 1578
rect 2047 1582 2051 1583
rect 2047 1577 2051 1578
rect 2079 1582 2083 1583
rect 2079 1577 2083 1578
rect 2207 1582 2211 1583
rect 2207 1577 2211 1578
rect 2343 1582 2347 1583
rect 2343 1577 2347 1578
rect 2367 1582 2371 1583
rect 2367 1577 2371 1578
rect 2487 1582 2491 1583
rect 2487 1577 2491 1578
rect 2527 1582 2531 1583
rect 2527 1577 2531 1578
rect 2631 1582 2635 1583
rect 2631 1577 2635 1578
rect 2687 1582 2691 1583
rect 2687 1577 2691 1578
rect 2775 1582 2779 1583
rect 2775 1577 2779 1578
rect 2839 1582 2843 1583
rect 2839 1577 2843 1578
rect 2919 1582 2923 1583
rect 2919 1577 2923 1578
rect 2983 1582 2987 1583
rect 2983 1577 2987 1578
rect 3063 1582 3067 1583
rect 3063 1577 3067 1578
rect 3119 1582 3123 1583
rect 3119 1577 3123 1578
rect 3215 1582 3219 1583
rect 3215 1577 3219 1578
rect 3255 1582 3259 1583
rect 3255 1577 3259 1578
rect 3367 1582 3371 1583
rect 3367 1577 3371 1578
rect 3391 1582 3395 1583
rect 3391 1577 3395 1578
rect 3503 1582 3507 1583
rect 3503 1577 3507 1578
rect 3591 1582 3595 1583
rect 3591 1577 3595 1578
rect 110 1572 116 1573
rect 1830 1573 1831 1577
rect 1835 1573 1836 1577
rect 1830 1572 1836 1573
rect 110 1560 116 1561
rect 110 1556 111 1560
rect 115 1556 116 1560
rect 110 1555 116 1556
rect 1830 1560 1836 1561
rect 1830 1556 1831 1560
rect 1835 1556 1836 1560
rect 1872 1558 1874 1577
rect 1896 1561 1898 1577
rect 2048 1561 2050 1577
rect 2208 1561 2210 1577
rect 2368 1561 2370 1577
rect 2528 1561 2530 1577
rect 2688 1561 2690 1577
rect 2840 1561 2842 1577
rect 2984 1561 2986 1577
rect 3120 1561 3122 1577
rect 3256 1561 3258 1577
rect 3392 1561 3394 1577
rect 3504 1561 3506 1577
rect 1894 1560 1900 1561
rect 1830 1555 1836 1556
rect 1870 1557 1876 1558
rect 112 1523 114 1555
rect 166 1542 172 1543
rect 166 1538 167 1542
rect 171 1538 172 1542
rect 166 1537 172 1538
rect 294 1542 300 1543
rect 294 1538 295 1542
rect 299 1538 300 1542
rect 294 1537 300 1538
rect 430 1542 436 1543
rect 430 1538 431 1542
rect 435 1538 436 1542
rect 430 1537 436 1538
rect 574 1542 580 1543
rect 574 1538 575 1542
rect 579 1538 580 1542
rect 574 1537 580 1538
rect 718 1542 724 1543
rect 718 1538 719 1542
rect 723 1538 724 1542
rect 718 1537 724 1538
rect 854 1542 860 1543
rect 854 1538 855 1542
rect 859 1538 860 1542
rect 854 1537 860 1538
rect 990 1542 996 1543
rect 990 1538 991 1542
rect 995 1538 996 1542
rect 990 1537 996 1538
rect 1126 1542 1132 1543
rect 1126 1538 1127 1542
rect 1131 1538 1132 1542
rect 1126 1537 1132 1538
rect 1254 1542 1260 1543
rect 1254 1538 1255 1542
rect 1259 1538 1260 1542
rect 1254 1537 1260 1538
rect 1382 1542 1388 1543
rect 1382 1538 1383 1542
rect 1387 1538 1388 1542
rect 1382 1537 1388 1538
rect 1518 1542 1524 1543
rect 1518 1538 1519 1542
rect 1523 1538 1524 1542
rect 1518 1537 1524 1538
rect 168 1523 170 1537
rect 296 1523 298 1537
rect 432 1523 434 1537
rect 576 1523 578 1537
rect 720 1523 722 1537
rect 856 1523 858 1537
rect 992 1523 994 1537
rect 1128 1523 1130 1537
rect 1256 1523 1258 1537
rect 1384 1523 1386 1537
rect 1520 1523 1522 1537
rect 1832 1523 1834 1555
rect 1870 1553 1871 1557
rect 1875 1553 1876 1557
rect 1894 1556 1895 1560
rect 1899 1556 1900 1560
rect 1894 1555 1900 1556
rect 2046 1560 2052 1561
rect 2046 1556 2047 1560
rect 2051 1556 2052 1560
rect 2046 1555 2052 1556
rect 2206 1560 2212 1561
rect 2206 1556 2207 1560
rect 2211 1556 2212 1560
rect 2206 1555 2212 1556
rect 2366 1560 2372 1561
rect 2366 1556 2367 1560
rect 2371 1556 2372 1560
rect 2366 1555 2372 1556
rect 2526 1560 2532 1561
rect 2526 1556 2527 1560
rect 2531 1556 2532 1560
rect 2526 1555 2532 1556
rect 2686 1560 2692 1561
rect 2686 1556 2687 1560
rect 2691 1556 2692 1560
rect 2686 1555 2692 1556
rect 2838 1560 2844 1561
rect 2838 1556 2839 1560
rect 2843 1556 2844 1560
rect 2838 1555 2844 1556
rect 2982 1560 2988 1561
rect 2982 1556 2983 1560
rect 2987 1556 2988 1560
rect 2982 1555 2988 1556
rect 3118 1560 3124 1561
rect 3118 1556 3119 1560
rect 3123 1556 3124 1560
rect 3118 1555 3124 1556
rect 3254 1560 3260 1561
rect 3254 1556 3255 1560
rect 3259 1556 3260 1560
rect 3254 1555 3260 1556
rect 3390 1560 3396 1561
rect 3390 1556 3391 1560
rect 3395 1556 3396 1560
rect 3390 1555 3396 1556
rect 3502 1560 3508 1561
rect 3502 1556 3503 1560
rect 3507 1556 3508 1560
rect 3592 1558 3594 1577
rect 3502 1555 3508 1556
rect 3590 1557 3596 1558
rect 1870 1552 1876 1553
rect 3590 1553 3591 1557
rect 3595 1553 3596 1557
rect 3590 1552 3596 1553
rect 1870 1540 1876 1541
rect 1870 1536 1871 1540
rect 1875 1536 1876 1540
rect 1870 1535 1876 1536
rect 3590 1540 3596 1541
rect 3590 1536 3591 1540
rect 3595 1536 3596 1540
rect 3590 1535 3596 1536
rect 111 1522 115 1523
rect 111 1517 115 1518
rect 167 1522 171 1523
rect 167 1517 171 1518
rect 231 1522 235 1523
rect 231 1517 235 1518
rect 295 1522 299 1523
rect 295 1517 299 1518
rect 375 1522 379 1523
rect 375 1517 379 1518
rect 431 1522 435 1523
rect 431 1517 435 1518
rect 519 1522 523 1523
rect 519 1517 523 1518
rect 575 1522 579 1523
rect 575 1517 579 1518
rect 655 1522 659 1523
rect 655 1517 659 1518
rect 719 1522 723 1523
rect 719 1517 723 1518
rect 783 1522 787 1523
rect 783 1517 787 1518
rect 855 1522 859 1523
rect 855 1517 859 1518
rect 903 1522 907 1523
rect 903 1517 907 1518
rect 991 1522 995 1523
rect 991 1517 995 1518
rect 1015 1522 1019 1523
rect 1015 1517 1019 1518
rect 1119 1522 1123 1523
rect 1119 1517 1123 1518
rect 1127 1522 1131 1523
rect 1127 1517 1131 1518
rect 1215 1522 1219 1523
rect 1215 1517 1219 1518
rect 1255 1522 1259 1523
rect 1255 1517 1259 1518
rect 1319 1522 1323 1523
rect 1319 1517 1323 1518
rect 1383 1522 1387 1523
rect 1383 1517 1387 1518
rect 1423 1522 1427 1523
rect 1423 1517 1427 1518
rect 1519 1522 1523 1523
rect 1519 1517 1523 1518
rect 1831 1522 1835 1523
rect 1831 1517 1835 1518
rect 112 1489 114 1517
rect 232 1507 234 1517
rect 376 1507 378 1517
rect 520 1507 522 1517
rect 656 1507 658 1517
rect 784 1507 786 1517
rect 904 1507 906 1517
rect 1016 1507 1018 1517
rect 1120 1507 1122 1517
rect 1216 1507 1218 1517
rect 1320 1507 1322 1517
rect 1424 1507 1426 1517
rect 230 1506 236 1507
rect 230 1502 231 1506
rect 235 1502 236 1506
rect 230 1501 236 1502
rect 374 1506 380 1507
rect 374 1502 375 1506
rect 379 1502 380 1506
rect 374 1501 380 1502
rect 518 1506 524 1507
rect 518 1502 519 1506
rect 523 1502 524 1506
rect 518 1501 524 1502
rect 654 1506 660 1507
rect 654 1502 655 1506
rect 659 1502 660 1506
rect 654 1501 660 1502
rect 782 1506 788 1507
rect 782 1502 783 1506
rect 787 1502 788 1506
rect 782 1501 788 1502
rect 902 1506 908 1507
rect 902 1502 903 1506
rect 907 1502 908 1506
rect 902 1501 908 1502
rect 1014 1506 1020 1507
rect 1014 1502 1015 1506
rect 1019 1502 1020 1506
rect 1014 1501 1020 1502
rect 1118 1506 1124 1507
rect 1118 1502 1119 1506
rect 1123 1502 1124 1506
rect 1118 1501 1124 1502
rect 1214 1506 1220 1507
rect 1214 1502 1215 1506
rect 1219 1502 1220 1506
rect 1214 1501 1220 1502
rect 1318 1506 1324 1507
rect 1318 1502 1319 1506
rect 1323 1502 1324 1506
rect 1318 1501 1324 1502
rect 1422 1506 1428 1507
rect 1422 1502 1423 1506
rect 1427 1502 1428 1506
rect 1422 1501 1428 1502
rect 1832 1489 1834 1517
rect 1872 1499 1874 1535
rect 1902 1522 1908 1523
rect 1902 1518 1903 1522
rect 1907 1518 1908 1522
rect 1902 1517 1908 1518
rect 2054 1522 2060 1523
rect 2054 1518 2055 1522
rect 2059 1518 2060 1522
rect 2054 1517 2060 1518
rect 2214 1522 2220 1523
rect 2214 1518 2215 1522
rect 2219 1518 2220 1522
rect 2214 1517 2220 1518
rect 2374 1522 2380 1523
rect 2374 1518 2375 1522
rect 2379 1518 2380 1522
rect 2374 1517 2380 1518
rect 2534 1522 2540 1523
rect 2534 1518 2535 1522
rect 2539 1518 2540 1522
rect 2534 1517 2540 1518
rect 2694 1522 2700 1523
rect 2694 1518 2695 1522
rect 2699 1518 2700 1522
rect 2694 1517 2700 1518
rect 2846 1522 2852 1523
rect 2846 1518 2847 1522
rect 2851 1518 2852 1522
rect 2846 1517 2852 1518
rect 2990 1522 2996 1523
rect 2990 1518 2991 1522
rect 2995 1518 2996 1522
rect 2990 1517 2996 1518
rect 3126 1522 3132 1523
rect 3126 1518 3127 1522
rect 3131 1518 3132 1522
rect 3126 1517 3132 1518
rect 3262 1522 3268 1523
rect 3262 1518 3263 1522
rect 3267 1518 3268 1522
rect 3262 1517 3268 1518
rect 3398 1522 3404 1523
rect 3398 1518 3399 1522
rect 3403 1518 3404 1522
rect 3398 1517 3404 1518
rect 3510 1522 3516 1523
rect 3510 1518 3511 1522
rect 3515 1518 3516 1522
rect 3510 1517 3516 1518
rect 1904 1499 1906 1517
rect 2056 1499 2058 1517
rect 2216 1499 2218 1517
rect 2376 1499 2378 1517
rect 2536 1499 2538 1517
rect 2696 1499 2698 1517
rect 2848 1499 2850 1517
rect 2992 1499 2994 1517
rect 3128 1499 3130 1517
rect 3264 1499 3266 1517
rect 3400 1499 3402 1517
rect 3512 1499 3514 1517
rect 3592 1499 3594 1535
rect 1871 1498 1875 1499
rect 1871 1493 1875 1494
rect 1903 1498 1907 1499
rect 1903 1493 1907 1494
rect 2007 1498 2011 1499
rect 2007 1493 2011 1494
rect 2055 1498 2059 1499
rect 2055 1493 2059 1494
rect 2135 1498 2139 1499
rect 2135 1493 2139 1494
rect 2215 1498 2219 1499
rect 2215 1493 2219 1494
rect 2271 1498 2275 1499
rect 2271 1493 2275 1494
rect 2375 1498 2379 1499
rect 2375 1493 2379 1494
rect 2415 1498 2419 1499
rect 2415 1493 2419 1494
rect 2535 1498 2539 1499
rect 2535 1493 2539 1494
rect 2567 1498 2571 1499
rect 2567 1493 2571 1494
rect 2695 1498 2699 1499
rect 2695 1493 2699 1494
rect 2719 1498 2723 1499
rect 2719 1493 2723 1494
rect 2847 1498 2851 1499
rect 2847 1493 2851 1494
rect 2879 1498 2883 1499
rect 2879 1493 2883 1494
rect 2991 1498 2995 1499
rect 2991 1493 2995 1494
rect 3039 1498 3043 1499
rect 3039 1493 3043 1494
rect 3127 1498 3131 1499
rect 3127 1493 3131 1494
rect 3199 1498 3203 1499
rect 3199 1493 3203 1494
rect 3263 1498 3267 1499
rect 3263 1493 3267 1494
rect 3367 1498 3371 1499
rect 3367 1493 3371 1494
rect 3399 1498 3403 1499
rect 3399 1493 3403 1494
rect 3511 1498 3515 1499
rect 3511 1493 3515 1494
rect 3591 1498 3595 1499
rect 3591 1493 3595 1494
rect 110 1488 116 1489
rect 110 1484 111 1488
rect 115 1484 116 1488
rect 110 1483 116 1484
rect 1830 1488 1836 1489
rect 1830 1484 1831 1488
rect 1835 1484 1836 1488
rect 1830 1483 1836 1484
rect 110 1471 116 1472
rect 110 1467 111 1471
rect 115 1467 116 1471
rect 1830 1471 1836 1472
rect 110 1466 116 1467
rect 222 1468 228 1469
rect 112 1439 114 1466
rect 222 1464 223 1468
rect 227 1464 228 1468
rect 222 1463 228 1464
rect 366 1468 372 1469
rect 366 1464 367 1468
rect 371 1464 372 1468
rect 366 1463 372 1464
rect 510 1468 516 1469
rect 510 1464 511 1468
rect 515 1464 516 1468
rect 510 1463 516 1464
rect 646 1468 652 1469
rect 646 1464 647 1468
rect 651 1464 652 1468
rect 646 1463 652 1464
rect 774 1468 780 1469
rect 774 1464 775 1468
rect 779 1464 780 1468
rect 774 1463 780 1464
rect 894 1468 900 1469
rect 894 1464 895 1468
rect 899 1464 900 1468
rect 894 1463 900 1464
rect 1006 1468 1012 1469
rect 1006 1464 1007 1468
rect 1011 1464 1012 1468
rect 1006 1463 1012 1464
rect 1110 1468 1116 1469
rect 1110 1464 1111 1468
rect 1115 1464 1116 1468
rect 1110 1463 1116 1464
rect 1206 1468 1212 1469
rect 1206 1464 1207 1468
rect 1211 1464 1212 1468
rect 1206 1463 1212 1464
rect 1310 1468 1316 1469
rect 1310 1464 1311 1468
rect 1315 1464 1316 1468
rect 1310 1463 1316 1464
rect 1414 1468 1420 1469
rect 1414 1464 1415 1468
rect 1419 1464 1420 1468
rect 1830 1467 1831 1471
rect 1835 1467 1836 1471
rect 1830 1466 1836 1467
rect 1414 1463 1420 1464
rect 224 1439 226 1463
rect 368 1439 370 1463
rect 512 1439 514 1463
rect 648 1439 650 1463
rect 776 1439 778 1463
rect 896 1439 898 1463
rect 1008 1439 1010 1463
rect 1112 1439 1114 1463
rect 1208 1439 1210 1463
rect 1312 1439 1314 1463
rect 1416 1439 1418 1463
rect 1832 1439 1834 1466
rect 1872 1465 1874 1493
rect 1904 1483 1906 1493
rect 2008 1483 2010 1493
rect 2136 1483 2138 1493
rect 2272 1483 2274 1493
rect 2416 1483 2418 1493
rect 2568 1483 2570 1493
rect 2720 1483 2722 1493
rect 2880 1483 2882 1493
rect 3040 1483 3042 1493
rect 3200 1483 3202 1493
rect 3368 1483 3370 1493
rect 3512 1483 3514 1493
rect 1902 1482 1908 1483
rect 1902 1478 1903 1482
rect 1907 1478 1908 1482
rect 1902 1477 1908 1478
rect 2006 1482 2012 1483
rect 2006 1478 2007 1482
rect 2011 1478 2012 1482
rect 2006 1477 2012 1478
rect 2134 1482 2140 1483
rect 2134 1478 2135 1482
rect 2139 1478 2140 1482
rect 2134 1477 2140 1478
rect 2270 1482 2276 1483
rect 2270 1478 2271 1482
rect 2275 1478 2276 1482
rect 2270 1477 2276 1478
rect 2414 1482 2420 1483
rect 2414 1478 2415 1482
rect 2419 1478 2420 1482
rect 2414 1477 2420 1478
rect 2566 1482 2572 1483
rect 2566 1478 2567 1482
rect 2571 1478 2572 1482
rect 2566 1477 2572 1478
rect 2718 1482 2724 1483
rect 2718 1478 2719 1482
rect 2723 1478 2724 1482
rect 2718 1477 2724 1478
rect 2878 1482 2884 1483
rect 2878 1478 2879 1482
rect 2883 1478 2884 1482
rect 2878 1477 2884 1478
rect 3038 1482 3044 1483
rect 3038 1478 3039 1482
rect 3043 1478 3044 1482
rect 3038 1477 3044 1478
rect 3198 1482 3204 1483
rect 3198 1478 3199 1482
rect 3203 1478 3204 1482
rect 3198 1477 3204 1478
rect 3366 1482 3372 1483
rect 3366 1478 3367 1482
rect 3371 1478 3372 1482
rect 3366 1477 3372 1478
rect 3510 1482 3516 1483
rect 3510 1478 3511 1482
rect 3515 1478 3516 1482
rect 3510 1477 3516 1478
rect 3592 1465 3594 1493
rect 1870 1464 1876 1465
rect 1870 1460 1871 1464
rect 1875 1460 1876 1464
rect 1870 1459 1876 1460
rect 3590 1464 3596 1465
rect 3590 1460 3591 1464
rect 3595 1460 3596 1464
rect 3590 1459 3596 1460
rect 1870 1447 1876 1448
rect 1870 1443 1871 1447
rect 1875 1443 1876 1447
rect 3590 1447 3596 1448
rect 1870 1442 1876 1443
rect 1894 1444 1900 1445
rect 111 1438 115 1439
rect 111 1433 115 1434
rect 223 1438 227 1439
rect 223 1433 227 1434
rect 255 1438 259 1439
rect 255 1433 259 1434
rect 351 1438 355 1439
rect 351 1433 355 1434
rect 367 1438 371 1439
rect 367 1433 371 1434
rect 447 1438 451 1439
rect 447 1433 451 1434
rect 511 1438 515 1439
rect 511 1433 515 1434
rect 543 1438 547 1439
rect 543 1433 547 1434
rect 631 1438 635 1439
rect 631 1433 635 1434
rect 647 1438 651 1439
rect 647 1433 651 1434
rect 719 1438 723 1439
rect 719 1433 723 1434
rect 775 1438 779 1439
rect 775 1433 779 1434
rect 807 1438 811 1439
rect 807 1433 811 1434
rect 895 1438 899 1439
rect 895 1433 899 1434
rect 919 1438 923 1439
rect 919 1433 923 1434
rect 1007 1438 1011 1439
rect 1007 1433 1011 1434
rect 1047 1438 1051 1439
rect 1047 1433 1051 1434
rect 1111 1438 1115 1439
rect 1111 1433 1115 1434
rect 1207 1438 1211 1439
rect 1207 1433 1211 1434
rect 1311 1438 1315 1439
rect 1311 1433 1315 1434
rect 1383 1438 1387 1439
rect 1383 1433 1387 1434
rect 1415 1438 1419 1439
rect 1415 1433 1419 1434
rect 1575 1438 1579 1439
rect 1575 1433 1579 1434
rect 1743 1438 1747 1439
rect 1743 1433 1747 1434
rect 1831 1438 1835 1439
rect 1831 1433 1835 1434
rect 112 1414 114 1433
rect 256 1417 258 1433
rect 352 1417 354 1433
rect 448 1417 450 1433
rect 544 1417 546 1433
rect 632 1417 634 1433
rect 720 1417 722 1433
rect 808 1417 810 1433
rect 920 1417 922 1433
rect 1048 1417 1050 1433
rect 1208 1417 1210 1433
rect 1384 1417 1386 1433
rect 1576 1417 1578 1433
rect 1744 1417 1746 1433
rect 254 1416 260 1417
rect 110 1413 116 1414
rect 110 1409 111 1413
rect 115 1409 116 1413
rect 254 1412 255 1416
rect 259 1412 260 1416
rect 254 1411 260 1412
rect 350 1416 356 1417
rect 350 1412 351 1416
rect 355 1412 356 1416
rect 350 1411 356 1412
rect 446 1416 452 1417
rect 446 1412 447 1416
rect 451 1412 452 1416
rect 446 1411 452 1412
rect 542 1416 548 1417
rect 542 1412 543 1416
rect 547 1412 548 1416
rect 542 1411 548 1412
rect 630 1416 636 1417
rect 630 1412 631 1416
rect 635 1412 636 1416
rect 630 1411 636 1412
rect 718 1416 724 1417
rect 718 1412 719 1416
rect 723 1412 724 1416
rect 718 1411 724 1412
rect 806 1416 812 1417
rect 806 1412 807 1416
rect 811 1412 812 1416
rect 806 1411 812 1412
rect 918 1416 924 1417
rect 918 1412 919 1416
rect 923 1412 924 1416
rect 918 1411 924 1412
rect 1046 1416 1052 1417
rect 1046 1412 1047 1416
rect 1051 1412 1052 1416
rect 1046 1411 1052 1412
rect 1206 1416 1212 1417
rect 1206 1412 1207 1416
rect 1211 1412 1212 1416
rect 1206 1411 1212 1412
rect 1382 1416 1388 1417
rect 1382 1412 1383 1416
rect 1387 1412 1388 1416
rect 1382 1411 1388 1412
rect 1574 1416 1580 1417
rect 1574 1412 1575 1416
rect 1579 1412 1580 1416
rect 1574 1411 1580 1412
rect 1742 1416 1748 1417
rect 1742 1412 1743 1416
rect 1747 1412 1748 1416
rect 1832 1414 1834 1433
rect 1872 1423 1874 1442
rect 1894 1440 1895 1444
rect 1899 1440 1900 1444
rect 1894 1439 1900 1440
rect 1998 1444 2004 1445
rect 1998 1440 1999 1444
rect 2003 1440 2004 1444
rect 1998 1439 2004 1440
rect 2126 1444 2132 1445
rect 2126 1440 2127 1444
rect 2131 1440 2132 1444
rect 2126 1439 2132 1440
rect 2262 1444 2268 1445
rect 2262 1440 2263 1444
rect 2267 1440 2268 1444
rect 2262 1439 2268 1440
rect 2406 1444 2412 1445
rect 2406 1440 2407 1444
rect 2411 1440 2412 1444
rect 2406 1439 2412 1440
rect 2558 1444 2564 1445
rect 2558 1440 2559 1444
rect 2563 1440 2564 1444
rect 2558 1439 2564 1440
rect 2710 1444 2716 1445
rect 2710 1440 2711 1444
rect 2715 1440 2716 1444
rect 2710 1439 2716 1440
rect 2870 1444 2876 1445
rect 2870 1440 2871 1444
rect 2875 1440 2876 1444
rect 2870 1439 2876 1440
rect 3030 1444 3036 1445
rect 3030 1440 3031 1444
rect 3035 1440 3036 1444
rect 3030 1439 3036 1440
rect 3190 1444 3196 1445
rect 3190 1440 3191 1444
rect 3195 1440 3196 1444
rect 3190 1439 3196 1440
rect 3358 1444 3364 1445
rect 3358 1440 3359 1444
rect 3363 1440 3364 1444
rect 3358 1439 3364 1440
rect 3502 1444 3508 1445
rect 3502 1440 3503 1444
rect 3507 1440 3508 1444
rect 3590 1443 3591 1447
rect 3595 1443 3596 1447
rect 3590 1442 3596 1443
rect 3502 1439 3508 1440
rect 1896 1423 1898 1439
rect 2000 1423 2002 1439
rect 2128 1423 2130 1439
rect 2264 1423 2266 1439
rect 2408 1423 2410 1439
rect 2560 1423 2562 1439
rect 2712 1423 2714 1439
rect 2872 1423 2874 1439
rect 3032 1423 3034 1439
rect 3192 1423 3194 1439
rect 3360 1423 3362 1439
rect 3504 1423 3506 1439
rect 3592 1423 3594 1442
rect 1871 1422 1875 1423
rect 1871 1417 1875 1418
rect 1895 1422 1899 1423
rect 1895 1417 1899 1418
rect 1999 1422 2003 1423
rect 1999 1417 2003 1418
rect 2023 1422 2027 1423
rect 2023 1417 2027 1418
rect 2127 1422 2131 1423
rect 2127 1417 2131 1418
rect 2167 1422 2171 1423
rect 2167 1417 2171 1418
rect 2263 1422 2267 1423
rect 2263 1417 2267 1418
rect 2303 1422 2307 1423
rect 2303 1417 2307 1418
rect 2407 1422 2411 1423
rect 2407 1417 2411 1418
rect 2431 1422 2435 1423
rect 2431 1417 2435 1418
rect 2551 1422 2555 1423
rect 2551 1417 2555 1418
rect 2559 1422 2563 1423
rect 2559 1417 2563 1418
rect 2671 1422 2675 1423
rect 2671 1417 2675 1418
rect 2711 1422 2715 1423
rect 2711 1417 2715 1418
rect 2791 1422 2795 1423
rect 2791 1417 2795 1418
rect 2871 1422 2875 1423
rect 2871 1417 2875 1418
rect 2911 1422 2915 1423
rect 2911 1417 2915 1418
rect 3031 1422 3035 1423
rect 3031 1417 3035 1418
rect 3191 1422 3195 1423
rect 3191 1417 3195 1418
rect 3359 1422 3363 1423
rect 3359 1417 3363 1418
rect 3503 1422 3507 1423
rect 3503 1417 3507 1418
rect 3591 1422 3595 1423
rect 3591 1417 3595 1418
rect 1742 1411 1748 1412
rect 1830 1413 1836 1414
rect 110 1408 116 1409
rect 1830 1409 1831 1413
rect 1835 1409 1836 1413
rect 1830 1408 1836 1409
rect 1872 1398 1874 1417
rect 1896 1401 1898 1417
rect 2024 1401 2026 1417
rect 2168 1401 2170 1417
rect 2304 1401 2306 1417
rect 2432 1401 2434 1417
rect 2552 1401 2554 1417
rect 2672 1401 2674 1417
rect 2792 1401 2794 1417
rect 2912 1401 2914 1417
rect 1894 1400 1900 1401
rect 1870 1397 1876 1398
rect 110 1396 116 1397
rect 110 1392 111 1396
rect 115 1392 116 1396
rect 110 1391 116 1392
rect 1830 1396 1836 1397
rect 1830 1392 1831 1396
rect 1835 1392 1836 1396
rect 1870 1393 1871 1397
rect 1875 1393 1876 1397
rect 1894 1396 1895 1400
rect 1899 1396 1900 1400
rect 1894 1395 1900 1396
rect 2022 1400 2028 1401
rect 2022 1396 2023 1400
rect 2027 1396 2028 1400
rect 2022 1395 2028 1396
rect 2166 1400 2172 1401
rect 2166 1396 2167 1400
rect 2171 1396 2172 1400
rect 2166 1395 2172 1396
rect 2302 1400 2308 1401
rect 2302 1396 2303 1400
rect 2307 1396 2308 1400
rect 2302 1395 2308 1396
rect 2430 1400 2436 1401
rect 2430 1396 2431 1400
rect 2435 1396 2436 1400
rect 2430 1395 2436 1396
rect 2550 1400 2556 1401
rect 2550 1396 2551 1400
rect 2555 1396 2556 1400
rect 2550 1395 2556 1396
rect 2670 1400 2676 1401
rect 2670 1396 2671 1400
rect 2675 1396 2676 1400
rect 2670 1395 2676 1396
rect 2790 1400 2796 1401
rect 2790 1396 2791 1400
rect 2795 1396 2796 1400
rect 2790 1395 2796 1396
rect 2910 1400 2916 1401
rect 2910 1396 2911 1400
rect 2915 1396 2916 1400
rect 3592 1398 3594 1417
rect 2910 1395 2916 1396
rect 3590 1397 3596 1398
rect 1870 1392 1876 1393
rect 3590 1393 3591 1397
rect 3595 1393 3596 1397
rect 3590 1392 3596 1393
rect 1830 1391 1836 1392
rect 112 1363 114 1391
rect 262 1378 268 1379
rect 262 1374 263 1378
rect 267 1374 268 1378
rect 262 1373 268 1374
rect 358 1378 364 1379
rect 358 1374 359 1378
rect 363 1374 364 1378
rect 358 1373 364 1374
rect 454 1378 460 1379
rect 454 1374 455 1378
rect 459 1374 460 1378
rect 454 1373 460 1374
rect 550 1378 556 1379
rect 550 1374 551 1378
rect 555 1374 556 1378
rect 550 1373 556 1374
rect 638 1378 644 1379
rect 638 1374 639 1378
rect 643 1374 644 1378
rect 638 1373 644 1374
rect 726 1378 732 1379
rect 726 1374 727 1378
rect 731 1374 732 1378
rect 726 1373 732 1374
rect 814 1378 820 1379
rect 814 1374 815 1378
rect 819 1374 820 1378
rect 814 1373 820 1374
rect 926 1378 932 1379
rect 926 1374 927 1378
rect 931 1374 932 1378
rect 926 1373 932 1374
rect 1054 1378 1060 1379
rect 1054 1374 1055 1378
rect 1059 1374 1060 1378
rect 1054 1373 1060 1374
rect 1214 1378 1220 1379
rect 1214 1374 1215 1378
rect 1219 1374 1220 1378
rect 1214 1373 1220 1374
rect 1390 1378 1396 1379
rect 1390 1374 1391 1378
rect 1395 1374 1396 1378
rect 1390 1373 1396 1374
rect 1582 1378 1588 1379
rect 1582 1374 1583 1378
rect 1587 1374 1588 1378
rect 1582 1373 1588 1374
rect 1750 1378 1756 1379
rect 1750 1374 1751 1378
rect 1755 1374 1756 1378
rect 1750 1373 1756 1374
rect 264 1363 266 1373
rect 360 1363 362 1373
rect 456 1363 458 1373
rect 552 1363 554 1373
rect 640 1363 642 1373
rect 728 1363 730 1373
rect 816 1363 818 1373
rect 928 1363 930 1373
rect 1056 1363 1058 1373
rect 1216 1363 1218 1373
rect 1392 1363 1394 1373
rect 1584 1363 1586 1373
rect 1752 1363 1754 1373
rect 1832 1363 1834 1391
rect 1870 1380 1876 1381
rect 1870 1376 1871 1380
rect 1875 1376 1876 1380
rect 1870 1375 1876 1376
rect 3590 1380 3596 1381
rect 3590 1376 3591 1380
rect 3595 1376 3596 1380
rect 3590 1375 3596 1376
rect 111 1362 115 1363
rect 111 1357 115 1358
rect 263 1362 267 1363
rect 263 1357 267 1358
rect 359 1362 363 1363
rect 359 1357 363 1358
rect 455 1362 459 1363
rect 455 1357 459 1358
rect 471 1362 475 1363
rect 471 1357 475 1358
rect 551 1362 555 1363
rect 551 1357 555 1358
rect 591 1362 595 1363
rect 591 1357 595 1358
rect 639 1362 643 1363
rect 639 1357 643 1358
rect 727 1362 731 1363
rect 727 1357 731 1358
rect 815 1362 819 1363
rect 815 1357 819 1358
rect 863 1362 867 1363
rect 863 1357 867 1358
rect 927 1362 931 1363
rect 927 1357 931 1358
rect 1007 1362 1011 1363
rect 1007 1357 1011 1358
rect 1055 1362 1059 1363
rect 1055 1357 1059 1358
rect 1143 1362 1147 1363
rect 1143 1357 1147 1358
rect 1215 1362 1219 1363
rect 1215 1357 1219 1358
rect 1279 1362 1283 1363
rect 1279 1357 1283 1358
rect 1391 1362 1395 1363
rect 1391 1357 1395 1358
rect 1407 1362 1411 1363
rect 1407 1357 1411 1358
rect 1527 1362 1531 1363
rect 1527 1357 1531 1358
rect 1583 1362 1587 1363
rect 1583 1357 1587 1358
rect 1647 1362 1651 1363
rect 1647 1357 1651 1358
rect 1751 1362 1755 1363
rect 1751 1357 1755 1358
rect 1831 1362 1835 1363
rect 1831 1357 1835 1358
rect 112 1329 114 1357
rect 360 1347 362 1357
rect 472 1347 474 1357
rect 592 1347 594 1357
rect 728 1347 730 1357
rect 864 1347 866 1357
rect 1008 1347 1010 1357
rect 1144 1347 1146 1357
rect 1280 1347 1282 1357
rect 1408 1347 1410 1357
rect 1528 1347 1530 1357
rect 1648 1347 1650 1357
rect 1752 1347 1754 1357
rect 358 1346 364 1347
rect 358 1342 359 1346
rect 363 1342 364 1346
rect 358 1341 364 1342
rect 470 1346 476 1347
rect 470 1342 471 1346
rect 475 1342 476 1346
rect 470 1341 476 1342
rect 590 1346 596 1347
rect 590 1342 591 1346
rect 595 1342 596 1346
rect 590 1341 596 1342
rect 726 1346 732 1347
rect 726 1342 727 1346
rect 731 1342 732 1346
rect 726 1341 732 1342
rect 862 1346 868 1347
rect 862 1342 863 1346
rect 867 1342 868 1346
rect 862 1341 868 1342
rect 1006 1346 1012 1347
rect 1006 1342 1007 1346
rect 1011 1342 1012 1346
rect 1006 1341 1012 1342
rect 1142 1346 1148 1347
rect 1142 1342 1143 1346
rect 1147 1342 1148 1346
rect 1142 1341 1148 1342
rect 1278 1346 1284 1347
rect 1278 1342 1279 1346
rect 1283 1342 1284 1346
rect 1278 1341 1284 1342
rect 1406 1346 1412 1347
rect 1406 1342 1407 1346
rect 1411 1342 1412 1346
rect 1406 1341 1412 1342
rect 1526 1346 1532 1347
rect 1526 1342 1527 1346
rect 1531 1342 1532 1346
rect 1526 1341 1532 1342
rect 1646 1346 1652 1347
rect 1646 1342 1647 1346
rect 1651 1342 1652 1346
rect 1646 1341 1652 1342
rect 1750 1346 1756 1347
rect 1750 1342 1751 1346
rect 1755 1342 1756 1346
rect 1750 1341 1756 1342
rect 1832 1329 1834 1357
rect 1872 1339 1874 1375
rect 1902 1362 1908 1363
rect 1902 1358 1903 1362
rect 1907 1358 1908 1362
rect 1902 1357 1908 1358
rect 2030 1362 2036 1363
rect 2030 1358 2031 1362
rect 2035 1358 2036 1362
rect 2030 1357 2036 1358
rect 2174 1362 2180 1363
rect 2174 1358 2175 1362
rect 2179 1358 2180 1362
rect 2174 1357 2180 1358
rect 2310 1362 2316 1363
rect 2310 1358 2311 1362
rect 2315 1358 2316 1362
rect 2310 1357 2316 1358
rect 2438 1362 2444 1363
rect 2438 1358 2439 1362
rect 2443 1358 2444 1362
rect 2438 1357 2444 1358
rect 2558 1362 2564 1363
rect 2558 1358 2559 1362
rect 2563 1358 2564 1362
rect 2558 1357 2564 1358
rect 2678 1362 2684 1363
rect 2678 1358 2679 1362
rect 2683 1358 2684 1362
rect 2678 1357 2684 1358
rect 2798 1362 2804 1363
rect 2798 1358 2799 1362
rect 2803 1358 2804 1362
rect 2798 1357 2804 1358
rect 2918 1362 2924 1363
rect 2918 1358 2919 1362
rect 2923 1358 2924 1362
rect 2918 1357 2924 1358
rect 1904 1339 1906 1357
rect 2032 1339 2034 1357
rect 2176 1339 2178 1357
rect 2312 1339 2314 1357
rect 2440 1339 2442 1357
rect 2560 1339 2562 1357
rect 2680 1339 2682 1357
rect 2800 1339 2802 1357
rect 2920 1339 2922 1357
rect 3592 1339 3594 1375
rect 1871 1338 1875 1339
rect 1871 1333 1875 1334
rect 1903 1338 1907 1339
rect 1903 1333 1907 1334
rect 1927 1338 1931 1339
rect 1927 1333 1931 1334
rect 2031 1338 2035 1339
rect 2031 1333 2035 1334
rect 2047 1338 2051 1339
rect 2047 1333 2051 1334
rect 2175 1338 2179 1339
rect 2175 1333 2179 1334
rect 2183 1338 2187 1339
rect 2183 1333 2187 1334
rect 2311 1338 2315 1339
rect 2311 1333 2315 1334
rect 2319 1338 2323 1339
rect 2319 1333 2323 1334
rect 2439 1338 2443 1339
rect 2439 1333 2443 1334
rect 2455 1338 2459 1339
rect 2455 1333 2459 1334
rect 2559 1338 2563 1339
rect 2559 1333 2563 1334
rect 2591 1338 2595 1339
rect 2591 1333 2595 1334
rect 2679 1338 2683 1339
rect 2679 1333 2683 1334
rect 2719 1338 2723 1339
rect 2719 1333 2723 1334
rect 2799 1338 2803 1339
rect 2799 1333 2803 1334
rect 2839 1338 2843 1339
rect 2839 1333 2843 1334
rect 2919 1338 2923 1339
rect 2919 1333 2923 1334
rect 2951 1338 2955 1339
rect 2951 1333 2955 1334
rect 3063 1338 3067 1339
rect 3063 1333 3067 1334
rect 3183 1338 3187 1339
rect 3183 1333 3187 1334
rect 3591 1338 3595 1339
rect 3591 1333 3595 1334
rect 110 1328 116 1329
rect 110 1324 111 1328
rect 115 1324 116 1328
rect 110 1323 116 1324
rect 1830 1328 1836 1329
rect 1830 1324 1831 1328
rect 1835 1324 1836 1328
rect 1830 1323 1836 1324
rect 110 1311 116 1312
rect 110 1307 111 1311
rect 115 1307 116 1311
rect 1830 1311 1836 1312
rect 110 1306 116 1307
rect 350 1308 356 1309
rect 112 1283 114 1306
rect 350 1304 351 1308
rect 355 1304 356 1308
rect 350 1303 356 1304
rect 462 1308 468 1309
rect 462 1304 463 1308
rect 467 1304 468 1308
rect 462 1303 468 1304
rect 582 1308 588 1309
rect 582 1304 583 1308
rect 587 1304 588 1308
rect 582 1303 588 1304
rect 718 1308 724 1309
rect 718 1304 719 1308
rect 723 1304 724 1308
rect 718 1303 724 1304
rect 854 1308 860 1309
rect 854 1304 855 1308
rect 859 1304 860 1308
rect 854 1303 860 1304
rect 998 1308 1004 1309
rect 998 1304 999 1308
rect 1003 1304 1004 1308
rect 998 1303 1004 1304
rect 1134 1308 1140 1309
rect 1134 1304 1135 1308
rect 1139 1304 1140 1308
rect 1134 1303 1140 1304
rect 1270 1308 1276 1309
rect 1270 1304 1271 1308
rect 1275 1304 1276 1308
rect 1270 1303 1276 1304
rect 1398 1308 1404 1309
rect 1398 1304 1399 1308
rect 1403 1304 1404 1308
rect 1398 1303 1404 1304
rect 1518 1308 1524 1309
rect 1518 1304 1519 1308
rect 1523 1304 1524 1308
rect 1518 1303 1524 1304
rect 1638 1308 1644 1309
rect 1638 1304 1639 1308
rect 1643 1304 1644 1308
rect 1638 1303 1644 1304
rect 1742 1308 1748 1309
rect 1742 1304 1743 1308
rect 1747 1304 1748 1308
rect 1830 1307 1831 1311
rect 1835 1307 1836 1311
rect 1830 1306 1836 1307
rect 1742 1303 1748 1304
rect 352 1283 354 1303
rect 464 1283 466 1303
rect 584 1283 586 1303
rect 720 1283 722 1303
rect 856 1283 858 1303
rect 1000 1283 1002 1303
rect 1136 1283 1138 1303
rect 1272 1283 1274 1303
rect 1400 1283 1402 1303
rect 1520 1283 1522 1303
rect 1640 1283 1642 1303
rect 1744 1283 1746 1303
rect 1832 1283 1834 1306
rect 1872 1305 1874 1333
rect 1928 1323 1930 1333
rect 2048 1323 2050 1333
rect 2184 1323 2186 1333
rect 2320 1323 2322 1333
rect 2456 1323 2458 1333
rect 2592 1323 2594 1333
rect 2720 1323 2722 1333
rect 2840 1323 2842 1333
rect 2952 1323 2954 1333
rect 3064 1323 3066 1333
rect 3184 1323 3186 1333
rect 1926 1322 1932 1323
rect 1926 1318 1927 1322
rect 1931 1318 1932 1322
rect 1926 1317 1932 1318
rect 2046 1322 2052 1323
rect 2046 1318 2047 1322
rect 2051 1318 2052 1322
rect 2046 1317 2052 1318
rect 2182 1322 2188 1323
rect 2182 1318 2183 1322
rect 2187 1318 2188 1322
rect 2182 1317 2188 1318
rect 2318 1322 2324 1323
rect 2318 1318 2319 1322
rect 2323 1318 2324 1322
rect 2318 1317 2324 1318
rect 2454 1322 2460 1323
rect 2454 1318 2455 1322
rect 2459 1318 2460 1322
rect 2454 1317 2460 1318
rect 2590 1322 2596 1323
rect 2590 1318 2591 1322
rect 2595 1318 2596 1322
rect 2590 1317 2596 1318
rect 2718 1322 2724 1323
rect 2718 1318 2719 1322
rect 2723 1318 2724 1322
rect 2718 1317 2724 1318
rect 2838 1322 2844 1323
rect 2838 1318 2839 1322
rect 2843 1318 2844 1322
rect 2838 1317 2844 1318
rect 2950 1322 2956 1323
rect 2950 1318 2951 1322
rect 2955 1318 2956 1322
rect 2950 1317 2956 1318
rect 3062 1322 3068 1323
rect 3062 1318 3063 1322
rect 3067 1318 3068 1322
rect 3062 1317 3068 1318
rect 3182 1322 3188 1323
rect 3182 1318 3183 1322
rect 3187 1318 3188 1322
rect 3182 1317 3188 1318
rect 3592 1305 3594 1333
rect 1870 1304 1876 1305
rect 1870 1300 1871 1304
rect 1875 1300 1876 1304
rect 1870 1299 1876 1300
rect 3590 1304 3596 1305
rect 3590 1300 3591 1304
rect 3595 1300 3596 1304
rect 3590 1299 3596 1300
rect 1870 1287 1876 1288
rect 1870 1283 1871 1287
rect 1875 1283 1876 1287
rect 3590 1287 3596 1288
rect 111 1282 115 1283
rect 111 1277 115 1278
rect 311 1282 315 1283
rect 311 1277 315 1278
rect 351 1282 355 1283
rect 351 1277 355 1278
rect 415 1282 419 1283
rect 415 1277 419 1278
rect 463 1282 467 1283
rect 463 1277 467 1278
rect 535 1282 539 1283
rect 535 1277 539 1278
rect 583 1282 587 1283
rect 583 1277 587 1278
rect 671 1282 675 1283
rect 671 1277 675 1278
rect 719 1282 723 1283
rect 719 1277 723 1278
rect 815 1282 819 1283
rect 815 1277 819 1278
rect 855 1282 859 1283
rect 855 1277 859 1278
rect 959 1282 963 1283
rect 959 1277 963 1278
rect 999 1282 1003 1283
rect 999 1277 1003 1278
rect 1103 1282 1107 1283
rect 1103 1277 1107 1278
rect 1135 1282 1139 1283
rect 1135 1277 1139 1278
rect 1239 1282 1243 1283
rect 1239 1277 1243 1278
rect 1271 1282 1275 1283
rect 1271 1277 1275 1278
rect 1375 1282 1379 1283
rect 1375 1277 1379 1278
rect 1399 1282 1403 1283
rect 1399 1277 1403 1278
rect 1503 1282 1507 1283
rect 1503 1277 1507 1278
rect 1519 1282 1523 1283
rect 1519 1277 1523 1278
rect 1631 1282 1635 1283
rect 1631 1277 1635 1278
rect 1639 1282 1643 1283
rect 1639 1277 1643 1278
rect 1743 1282 1747 1283
rect 1743 1277 1747 1278
rect 1831 1282 1835 1283
rect 1870 1282 1876 1283
rect 1918 1284 1924 1285
rect 1831 1277 1835 1278
rect 112 1258 114 1277
rect 312 1261 314 1277
rect 416 1261 418 1277
rect 536 1261 538 1277
rect 672 1261 674 1277
rect 816 1261 818 1277
rect 960 1261 962 1277
rect 1104 1261 1106 1277
rect 1240 1261 1242 1277
rect 1376 1261 1378 1277
rect 1504 1261 1506 1277
rect 1632 1261 1634 1277
rect 1744 1261 1746 1277
rect 310 1260 316 1261
rect 110 1257 116 1258
rect 110 1253 111 1257
rect 115 1253 116 1257
rect 310 1256 311 1260
rect 315 1256 316 1260
rect 310 1255 316 1256
rect 414 1260 420 1261
rect 414 1256 415 1260
rect 419 1256 420 1260
rect 414 1255 420 1256
rect 534 1260 540 1261
rect 534 1256 535 1260
rect 539 1256 540 1260
rect 534 1255 540 1256
rect 670 1260 676 1261
rect 670 1256 671 1260
rect 675 1256 676 1260
rect 670 1255 676 1256
rect 814 1260 820 1261
rect 814 1256 815 1260
rect 819 1256 820 1260
rect 814 1255 820 1256
rect 958 1260 964 1261
rect 958 1256 959 1260
rect 963 1256 964 1260
rect 958 1255 964 1256
rect 1102 1260 1108 1261
rect 1102 1256 1103 1260
rect 1107 1256 1108 1260
rect 1102 1255 1108 1256
rect 1238 1260 1244 1261
rect 1238 1256 1239 1260
rect 1243 1256 1244 1260
rect 1238 1255 1244 1256
rect 1374 1260 1380 1261
rect 1374 1256 1375 1260
rect 1379 1256 1380 1260
rect 1374 1255 1380 1256
rect 1502 1260 1508 1261
rect 1502 1256 1503 1260
rect 1507 1256 1508 1260
rect 1502 1255 1508 1256
rect 1630 1260 1636 1261
rect 1630 1256 1631 1260
rect 1635 1256 1636 1260
rect 1630 1255 1636 1256
rect 1742 1260 1748 1261
rect 1742 1256 1743 1260
rect 1747 1256 1748 1260
rect 1832 1258 1834 1277
rect 1742 1255 1748 1256
rect 1830 1257 1836 1258
rect 110 1252 116 1253
rect 1830 1253 1831 1257
rect 1835 1253 1836 1257
rect 1872 1255 1874 1282
rect 1918 1280 1919 1284
rect 1923 1280 1924 1284
rect 1918 1279 1924 1280
rect 2038 1284 2044 1285
rect 2038 1280 2039 1284
rect 2043 1280 2044 1284
rect 2038 1279 2044 1280
rect 2174 1284 2180 1285
rect 2174 1280 2175 1284
rect 2179 1280 2180 1284
rect 2174 1279 2180 1280
rect 2310 1284 2316 1285
rect 2310 1280 2311 1284
rect 2315 1280 2316 1284
rect 2310 1279 2316 1280
rect 2446 1284 2452 1285
rect 2446 1280 2447 1284
rect 2451 1280 2452 1284
rect 2446 1279 2452 1280
rect 2582 1284 2588 1285
rect 2582 1280 2583 1284
rect 2587 1280 2588 1284
rect 2582 1279 2588 1280
rect 2710 1284 2716 1285
rect 2710 1280 2711 1284
rect 2715 1280 2716 1284
rect 2710 1279 2716 1280
rect 2830 1284 2836 1285
rect 2830 1280 2831 1284
rect 2835 1280 2836 1284
rect 2830 1279 2836 1280
rect 2942 1284 2948 1285
rect 2942 1280 2943 1284
rect 2947 1280 2948 1284
rect 2942 1279 2948 1280
rect 3054 1284 3060 1285
rect 3054 1280 3055 1284
rect 3059 1280 3060 1284
rect 3054 1279 3060 1280
rect 3174 1284 3180 1285
rect 3174 1280 3175 1284
rect 3179 1280 3180 1284
rect 3590 1283 3591 1287
rect 3595 1283 3596 1287
rect 3590 1282 3596 1283
rect 3174 1279 3180 1280
rect 1920 1255 1922 1279
rect 2040 1255 2042 1279
rect 2176 1255 2178 1279
rect 2312 1255 2314 1279
rect 2448 1255 2450 1279
rect 2584 1255 2586 1279
rect 2712 1255 2714 1279
rect 2832 1255 2834 1279
rect 2944 1255 2946 1279
rect 3056 1255 3058 1279
rect 3176 1255 3178 1279
rect 3592 1255 3594 1282
rect 1830 1252 1836 1253
rect 1871 1254 1875 1255
rect 1871 1249 1875 1250
rect 1895 1254 1899 1255
rect 1895 1249 1899 1250
rect 1919 1254 1923 1255
rect 1919 1249 1923 1250
rect 2039 1254 2043 1255
rect 2039 1249 2043 1250
rect 2071 1254 2075 1255
rect 2071 1249 2075 1250
rect 2175 1254 2179 1255
rect 2175 1249 2179 1250
rect 2271 1254 2275 1255
rect 2271 1249 2275 1250
rect 2311 1254 2315 1255
rect 2311 1249 2315 1250
rect 2447 1254 2451 1255
rect 2447 1249 2451 1250
rect 2471 1254 2475 1255
rect 2471 1249 2475 1250
rect 2583 1254 2587 1255
rect 2583 1249 2587 1250
rect 2663 1254 2667 1255
rect 2663 1249 2667 1250
rect 2711 1254 2715 1255
rect 2711 1249 2715 1250
rect 2831 1254 2835 1255
rect 2831 1249 2835 1250
rect 2847 1254 2851 1255
rect 2847 1249 2851 1250
rect 2943 1254 2947 1255
rect 2943 1249 2947 1250
rect 3023 1254 3027 1255
rect 3023 1249 3027 1250
rect 3055 1254 3059 1255
rect 3055 1249 3059 1250
rect 3175 1254 3179 1255
rect 3175 1249 3179 1250
rect 3191 1254 3195 1255
rect 3191 1249 3195 1250
rect 3359 1254 3363 1255
rect 3359 1249 3363 1250
rect 3503 1254 3507 1255
rect 3503 1249 3507 1250
rect 3591 1254 3595 1255
rect 3591 1249 3595 1250
rect 110 1240 116 1241
rect 110 1236 111 1240
rect 115 1236 116 1240
rect 110 1235 116 1236
rect 1830 1240 1836 1241
rect 1830 1236 1831 1240
rect 1835 1236 1836 1240
rect 1830 1235 1836 1236
rect 112 1207 114 1235
rect 318 1222 324 1223
rect 318 1218 319 1222
rect 323 1218 324 1222
rect 318 1217 324 1218
rect 422 1222 428 1223
rect 422 1218 423 1222
rect 427 1218 428 1222
rect 422 1217 428 1218
rect 542 1222 548 1223
rect 542 1218 543 1222
rect 547 1218 548 1222
rect 542 1217 548 1218
rect 678 1222 684 1223
rect 678 1218 679 1222
rect 683 1218 684 1222
rect 678 1217 684 1218
rect 822 1222 828 1223
rect 822 1218 823 1222
rect 827 1218 828 1222
rect 822 1217 828 1218
rect 966 1222 972 1223
rect 966 1218 967 1222
rect 971 1218 972 1222
rect 966 1217 972 1218
rect 1110 1222 1116 1223
rect 1110 1218 1111 1222
rect 1115 1218 1116 1222
rect 1110 1217 1116 1218
rect 1246 1222 1252 1223
rect 1246 1218 1247 1222
rect 1251 1218 1252 1222
rect 1246 1217 1252 1218
rect 1382 1222 1388 1223
rect 1382 1218 1383 1222
rect 1387 1218 1388 1222
rect 1382 1217 1388 1218
rect 1510 1222 1516 1223
rect 1510 1218 1511 1222
rect 1515 1218 1516 1222
rect 1510 1217 1516 1218
rect 1638 1222 1644 1223
rect 1638 1218 1639 1222
rect 1643 1218 1644 1222
rect 1638 1217 1644 1218
rect 1750 1222 1756 1223
rect 1750 1218 1751 1222
rect 1755 1218 1756 1222
rect 1750 1217 1756 1218
rect 320 1207 322 1217
rect 424 1207 426 1217
rect 544 1207 546 1217
rect 680 1207 682 1217
rect 824 1207 826 1217
rect 968 1207 970 1217
rect 1112 1207 1114 1217
rect 1248 1207 1250 1217
rect 1384 1207 1386 1217
rect 1512 1207 1514 1217
rect 1640 1207 1642 1217
rect 1752 1207 1754 1217
rect 1832 1207 1834 1235
rect 1872 1230 1874 1249
rect 1896 1233 1898 1249
rect 2072 1233 2074 1249
rect 2272 1233 2274 1249
rect 2472 1233 2474 1249
rect 2664 1233 2666 1249
rect 2848 1233 2850 1249
rect 3024 1233 3026 1249
rect 3192 1233 3194 1249
rect 3360 1233 3362 1249
rect 3504 1233 3506 1249
rect 1894 1232 1900 1233
rect 1870 1229 1876 1230
rect 1870 1225 1871 1229
rect 1875 1225 1876 1229
rect 1894 1228 1895 1232
rect 1899 1228 1900 1232
rect 1894 1227 1900 1228
rect 2070 1232 2076 1233
rect 2070 1228 2071 1232
rect 2075 1228 2076 1232
rect 2070 1227 2076 1228
rect 2270 1232 2276 1233
rect 2270 1228 2271 1232
rect 2275 1228 2276 1232
rect 2270 1227 2276 1228
rect 2470 1232 2476 1233
rect 2470 1228 2471 1232
rect 2475 1228 2476 1232
rect 2470 1227 2476 1228
rect 2662 1232 2668 1233
rect 2662 1228 2663 1232
rect 2667 1228 2668 1232
rect 2662 1227 2668 1228
rect 2846 1232 2852 1233
rect 2846 1228 2847 1232
rect 2851 1228 2852 1232
rect 2846 1227 2852 1228
rect 3022 1232 3028 1233
rect 3022 1228 3023 1232
rect 3027 1228 3028 1232
rect 3022 1227 3028 1228
rect 3190 1232 3196 1233
rect 3190 1228 3191 1232
rect 3195 1228 3196 1232
rect 3190 1227 3196 1228
rect 3358 1232 3364 1233
rect 3358 1228 3359 1232
rect 3363 1228 3364 1232
rect 3358 1227 3364 1228
rect 3502 1232 3508 1233
rect 3502 1228 3503 1232
rect 3507 1228 3508 1232
rect 3592 1230 3594 1249
rect 3502 1227 3508 1228
rect 3590 1229 3596 1230
rect 1870 1224 1876 1225
rect 3590 1225 3591 1229
rect 3595 1225 3596 1229
rect 3590 1224 3596 1225
rect 1870 1212 1876 1213
rect 1870 1208 1871 1212
rect 1875 1208 1876 1212
rect 1870 1207 1876 1208
rect 3590 1212 3596 1213
rect 3590 1208 3591 1212
rect 3595 1208 3596 1212
rect 3590 1207 3596 1208
rect 111 1206 115 1207
rect 111 1201 115 1202
rect 239 1206 243 1207
rect 239 1201 243 1202
rect 319 1206 323 1207
rect 319 1201 323 1202
rect 415 1206 419 1207
rect 415 1201 419 1202
rect 423 1206 427 1207
rect 423 1201 427 1202
rect 543 1206 547 1207
rect 543 1201 547 1202
rect 591 1206 595 1207
rect 591 1201 595 1202
rect 679 1206 683 1207
rect 679 1201 683 1202
rect 759 1206 763 1207
rect 759 1201 763 1202
rect 823 1206 827 1207
rect 823 1201 827 1202
rect 927 1206 931 1207
rect 927 1201 931 1202
rect 967 1206 971 1207
rect 967 1201 971 1202
rect 1079 1206 1083 1207
rect 1079 1201 1083 1202
rect 1111 1206 1115 1207
rect 1111 1201 1115 1202
rect 1223 1206 1227 1207
rect 1223 1201 1227 1202
rect 1247 1206 1251 1207
rect 1247 1201 1251 1202
rect 1367 1206 1371 1207
rect 1367 1201 1371 1202
rect 1383 1206 1387 1207
rect 1383 1201 1387 1202
rect 1503 1206 1507 1207
rect 1503 1201 1507 1202
rect 1511 1206 1515 1207
rect 1511 1201 1515 1202
rect 1639 1206 1643 1207
rect 1639 1201 1643 1202
rect 1751 1206 1755 1207
rect 1751 1201 1755 1202
rect 1831 1206 1835 1207
rect 1831 1201 1835 1202
rect 112 1173 114 1201
rect 240 1191 242 1201
rect 416 1191 418 1201
rect 592 1191 594 1201
rect 760 1191 762 1201
rect 928 1191 930 1201
rect 1080 1191 1082 1201
rect 1224 1191 1226 1201
rect 1368 1191 1370 1201
rect 1504 1191 1506 1201
rect 1640 1191 1642 1201
rect 1752 1191 1754 1201
rect 238 1190 244 1191
rect 238 1186 239 1190
rect 243 1186 244 1190
rect 238 1185 244 1186
rect 414 1190 420 1191
rect 414 1186 415 1190
rect 419 1186 420 1190
rect 414 1185 420 1186
rect 590 1190 596 1191
rect 590 1186 591 1190
rect 595 1186 596 1190
rect 590 1185 596 1186
rect 758 1190 764 1191
rect 758 1186 759 1190
rect 763 1186 764 1190
rect 758 1185 764 1186
rect 926 1190 932 1191
rect 926 1186 927 1190
rect 931 1186 932 1190
rect 926 1185 932 1186
rect 1078 1190 1084 1191
rect 1078 1186 1079 1190
rect 1083 1186 1084 1190
rect 1078 1185 1084 1186
rect 1222 1190 1228 1191
rect 1222 1186 1223 1190
rect 1227 1186 1228 1190
rect 1222 1185 1228 1186
rect 1366 1190 1372 1191
rect 1366 1186 1367 1190
rect 1371 1186 1372 1190
rect 1366 1185 1372 1186
rect 1502 1190 1508 1191
rect 1502 1186 1503 1190
rect 1507 1186 1508 1190
rect 1502 1185 1508 1186
rect 1638 1190 1644 1191
rect 1638 1186 1639 1190
rect 1643 1186 1644 1190
rect 1638 1185 1644 1186
rect 1750 1190 1756 1191
rect 1750 1186 1751 1190
rect 1755 1186 1756 1190
rect 1750 1185 1756 1186
rect 1832 1173 1834 1201
rect 1872 1175 1874 1207
rect 1902 1194 1908 1195
rect 1902 1190 1903 1194
rect 1907 1190 1908 1194
rect 1902 1189 1908 1190
rect 2078 1194 2084 1195
rect 2078 1190 2079 1194
rect 2083 1190 2084 1194
rect 2078 1189 2084 1190
rect 2278 1194 2284 1195
rect 2278 1190 2279 1194
rect 2283 1190 2284 1194
rect 2278 1189 2284 1190
rect 2478 1194 2484 1195
rect 2478 1190 2479 1194
rect 2483 1190 2484 1194
rect 2478 1189 2484 1190
rect 2670 1194 2676 1195
rect 2670 1190 2671 1194
rect 2675 1190 2676 1194
rect 2670 1189 2676 1190
rect 2854 1194 2860 1195
rect 2854 1190 2855 1194
rect 2859 1190 2860 1194
rect 2854 1189 2860 1190
rect 3030 1194 3036 1195
rect 3030 1190 3031 1194
rect 3035 1190 3036 1194
rect 3030 1189 3036 1190
rect 3198 1194 3204 1195
rect 3198 1190 3199 1194
rect 3203 1190 3204 1194
rect 3198 1189 3204 1190
rect 3366 1194 3372 1195
rect 3366 1190 3367 1194
rect 3371 1190 3372 1194
rect 3366 1189 3372 1190
rect 3510 1194 3516 1195
rect 3510 1190 3511 1194
rect 3515 1190 3516 1194
rect 3510 1189 3516 1190
rect 1904 1175 1906 1189
rect 2080 1175 2082 1189
rect 2280 1175 2282 1189
rect 2480 1175 2482 1189
rect 2672 1175 2674 1189
rect 2856 1175 2858 1189
rect 3032 1175 3034 1189
rect 3200 1175 3202 1189
rect 3368 1175 3370 1189
rect 3512 1175 3514 1189
rect 3592 1175 3594 1207
rect 1871 1174 1875 1175
rect 110 1172 116 1173
rect 110 1168 111 1172
rect 115 1168 116 1172
rect 110 1167 116 1168
rect 1830 1172 1836 1173
rect 1830 1168 1831 1172
rect 1835 1168 1836 1172
rect 1871 1169 1875 1170
rect 1903 1174 1907 1175
rect 1903 1169 1907 1170
rect 1983 1174 1987 1175
rect 1983 1169 1987 1170
rect 2079 1174 2083 1175
rect 2079 1169 2083 1170
rect 2087 1174 2091 1175
rect 2087 1169 2091 1170
rect 2215 1174 2219 1175
rect 2215 1169 2219 1170
rect 2279 1174 2283 1175
rect 2279 1169 2283 1170
rect 2367 1174 2371 1175
rect 2367 1169 2371 1170
rect 2479 1174 2483 1175
rect 2479 1169 2483 1170
rect 2527 1174 2531 1175
rect 2527 1169 2531 1170
rect 2671 1174 2675 1175
rect 2671 1169 2675 1170
rect 2687 1174 2691 1175
rect 2687 1169 2691 1170
rect 2839 1174 2843 1175
rect 2839 1169 2843 1170
rect 2855 1174 2859 1175
rect 2855 1169 2859 1170
rect 2983 1174 2987 1175
rect 2983 1169 2987 1170
rect 3031 1174 3035 1175
rect 3031 1169 3035 1170
rect 3127 1174 3131 1175
rect 3127 1169 3131 1170
rect 3199 1174 3203 1175
rect 3199 1169 3203 1170
rect 3263 1174 3267 1175
rect 3263 1169 3267 1170
rect 3367 1174 3371 1175
rect 3367 1169 3371 1170
rect 3399 1174 3403 1175
rect 3399 1169 3403 1170
rect 3511 1174 3515 1175
rect 3511 1169 3515 1170
rect 3591 1174 3595 1175
rect 3591 1169 3595 1170
rect 1830 1167 1836 1168
rect 110 1155 116 1156
rect 110 1151 111 1155
rect 115 1151 116 1155
rect 1830 1155 1836 1156
rect 110 1150 116 1151
rect 230 1152 236 1153
rect 112 1127 114 1150
rect 230 1148 231 1152
rect 235 1148 236 1152
rect 230 1147 236 1148
rect 406 1152 412 1153
rect 406 1148 407 1152
rect 411 1148 412 1152
rect 406 1147 412 1148
rect 582 1152 588 1153
rect 582 1148 583 1152
rect 587 1148 588 1152
rect 582 1147 588 1148
rect 750 1152 756 1153
rect 750 1148 751 1152
rect 755 1148 756 1152
rect 750 1147 756 1148
rect 918 1152 924 1153
rect 918 1148 919 1152
rect 923 1148 924 1152
rect 918 1147 924 1148
rect 1070 1152 1076 1153
rect 1070 1148 1071 1152
rect 1075 1148 1076 1152
rect 1070 1147 1076 1148
rect 1214 1152 1220 1153
rect 1214 1148 1215 1152
rect 1219 1148 1220 1152
rect 1214 1147 1220 1148
rect 1358 1152 1364 1153
rect 1358 1148 1359 1152
rect 1363 1148 1364 1152
rect 1358 1147 1364 1148
rect 1494 1152 1500 1153
rect 1494 1148 1495 1152
rect 1499 1148 1500 1152
rect 1494 1147 1500 1148
rect 1630 1152 1636 1153
rect 1630 1148 1631 1152
rect 1635 1148 1636 1152
rect 1630 1147 1636 1148
rect 1742 1152 1748 1153
rect 1742 1148 1743 1152
rect 1747 1148 1748 1152
rect 1830 1151 1831 1155
rect 1835 1151 1836 1155
rect 1830 1150 1836 1151
rect 1742 1147 1748 1148
rect 232 1127 234 1147
rect 408 1127 410 1147
rect 584 1127 586 1147
rect 752 1127 754 1147
rect 920 1127 922 1147
rect 1072 1127 1074 1147
rect 1216 1127 1218 1147
rect 1360 1127 1362 1147
rect 1496 1127 1498 1147
rect 1632 1127 1634 1147
rect 1744 1127 1746 1147
rect 1832 1127 1834 1150
rect 1872 1141 1874 1169
rect 1904 1159 1906 1169
rect 1984 1159 1986 1169
rect 2088 1159 2090 1169
rect 2216 1159 2218 1169
rect 2368 1159 2370 1169
rect 2528 1159 2530 1169
rect 2688 1159 2690 1169
rect 2840 1159 2842 1169
rect 2984 1159 2986 1169
rect 3128 1159 3130 1169
rect 3264 1159 3266 1169
rect 3400 1159 3402 1169
rect 3512 1159 3514 1169
rect 1902 1158 1908 1159
rect 1902 1154 1903 1158
rect 1907 1154 1908 1158
rect 1902 1153 1908 1154
rect 1982 1158 1988 1159
rect 1982 1154 1983 1158
rect 1987 1154 1988 1158
rect 1982 1153 1988 1154
rect 2086 1158 2092 1159
rect 2086 1154 2087 1158
rect 2091 1154 2092 1158
rect 2086 1153 2092 1154
rect 2214 1158 2220 1159
rect 2214 1154 2215 1158
rect 2219 1154 2220 1158
rect 2214 1153 2220 1154
rect 2366 1158 2372 1159
rect 2366 1154 2367 1158
rect 2371 1154 2372 1158
rect 2366 1153 2372 1154
rect 2526 1158 2532 1159
rect 2526 1154 2527 1158
rect 2531 1154 2532 1158
rect 2526 1153 2532 1154
rect 2686 1158 2692 1159
rect 2686 1154 2687 1158
rect 2691 1154 2692 1158
rect 2686 1153 2692 1154
rect 2838 1158 2844 1159
rect 2838 1154 2839 1158
rect 2843 1154 2844 1158
rect 2838 1153 2844 1154
rect 2982 1158 2988 1159
rect 2982 1154 2983 1158
rect 2987 1154 2988 1158
rect 2982 1153 2988 1154
rect 3126 1158 3132 1159
rect 3126 1154 3127 1158
rect 3131 1154 3132 1158
rect 3126 1153 3132 1154
rect 3262 1158 3268 1159
rect 3262 1154 3263 1158
rect 3267 1154 3268 1158
rect 3262 1153 3268 1154
rect 3398 1158 3404 1159
rect 3398 1154 3399 1158
rect 3403 1154 3404 1158
rect 3398 1153 3404 1154
rect 3510 1158 3516 1159
rect 3510 1154 3511 1158
rect 3515 1154 3516 1158
rect 3510 1153 3516 1154
rect 3592 1141 3594 1169
rect 1870 1140 1876 1141
rect 1870 1136 1871 1140
rect 1875 1136 1876 1140
rect 1870 1135 1876 1136
rect 3590 1140 3596 1141
rect 3590 1136 3591 1140
rect 3595 1136 3596 1140
rect 3590 1135 3596 1136
rect 111 1126 115 1127
rect 111 1121 115 1122
rect 143 1126 147 1127
rect 143 1121 147 1122
rect 231 1126 235 1127
rect 231 1121 235 1122
rect 279 1126 283 1127
rect 279 1121 283 1122
rect 407 1126 411 1127
rect 407 1121 411 1122
rect 423 1126 427 1127
rect 423 1121 427 1122
rect 567 1126 571 1127
rect 567 1121 571 1122
rect 583 1126 587 1127
rect 583 1121 587 1122
rect 711 1126 715 1127
rect 711 1121 715 1122
rect 751 1126 755 1127
rect 751 1121 755 1122
rect 847 1126 851 1127
rect 847 1121 851 1122
rect 919 1126 923 1127
rect 919 1121 923 1122
rect 975 1126 979 1127
rect 975 1121 979 1122
rect 1071 1126 1075 1127
rect 1071 1121 1075 1122
rect 1103 1126 1107 1127
rect 1103 1121 1107 1122
rect 1215 1126 1219 1127
rect 1215 1121 1219 1122
rect 1223 1126 1227 1127
rect 1223 1121 1227 1122
rect 1343 1126 1347 1127
rect 1343 1121 1347 1122
rect 1359 1126 1363 1127
rect 1359 1121 1363 1122
rect 1471 1126 1475 1127
rect 1471 1121 1475 1122
rect 1495 1126 1499 1127
rect 1495 1121 1499 1122
rect 1631 1126 1635 1127
rect 1631 1121 1635 1122
rect 1743 1126 1747 1127
rect 1743 1121 1747 1122
rect 1831 1126 1835 1127
rect 1831 1121 1835 1122
rect 1870 1123 1876 1124
rect 112 1102 114 1121
rect 144 1105 146 1121
rect 280 1105 282 1121
rect 424 1105 426 1121
rect 568 1105 570 1121
rect 712 1105 714 1121
rect 848 1105 850 1121
rect 976 1105 978 1121
rect 1104 1105 1106 1121
rect 1224 1105 1226 1121
rect 1344 1105 1346 1121
rect 1472 1105 1474 1121
rect 142 1104 148 1105
rect 110 1101 116 1102
rect 110 1097 111 1101
rect 115 1097 116 1101
rect 142 1100 143 1104
rect 147 1100 148 1104
rect 142 1099 148 1100
rect 278 1104 284 1105
rect 278 1100 279 1104
rect 283 1100 284 1104
rect 278 1099 284 1100
rect 422 1104 428 1105
rect 422 1100 423 1104
rect 427 1100 428 1104
rect 422 1099 428 1100
rect 566 1104 572 1105
rect 566 1100 567 1104
rect 571 1100 572 1104
rect 566 1099 572 1100
rect 710 1104 716 1105
rect 710 1100 711 1104
rect 715 1100 716 1104
rect 710 1099 716 1100
rect 846 1104 852 1105
rect 846 1100 847 1104
rect 851 1100 852 1104
rect 846 1099 852 1100
rect 974 1104 980 1105
rect 974 1100 975 1104
rect 979 1100 980 1104
rect 974 1099 980 1100
rect 1102 1104 1108 1105
rect 1102 1100 1103 1104
rect 1107 1100 1108 1104
rect 1102 1099 1108 1100
rect 1222 1104 1228 1105
rect 1222 1100 1223 1104
rect 1227 1100 1228 1104
rect 1222 1099 1228 1100
rect 1342 1104 1348 1105
rect 1342 1100 1343 1104
rect 1347 1100 1348 1104
rect 1342 1099 1348 1100
rect 1470 1104 1476 1105
rect 1470 1100 1471 1104
rect 1475 1100 1476 1104
rect 1832 1102 1834 1121
rect 1870 1119 1871 1123
rect 1875 1119 1876 1123
rect 3590 1123 3596 1124
rect 1870 1118 1876 1119
rect 1894 1120 1900 1121
rect 1470 1099 1476 1100
rect 1830 1101 1836 1102
rect 110 1096 116 1097
rect 1830 1097 1831 1101
rect 1835 1097 1836 1101
rect 1830 1096 1836 1097
rect 1872 1091 1874 1118
rect 1894 1116 1895 1120
rect 1899 1116 1900 1120
rect 1894 1115 1900 1116
rect 1974 1120 1980 1121
rect 1974 1116 1975 1120
rect 1979 1116 1980 1120
rect 1974 1115 1980 1116
rect 2078 1120 2084 1121
rect 2078 1116 2079 1120
rect 2083 1116 2084 1120
rect 2078 1115 2084 1116
rect 2206 1120 2212 1121
rect 2206 1116 2207 1120
rect 2211 1116 2212 1120
rect 2206 1115 2212 1116
rect 2358 1120 2364 1121
rect 2358 1116 2359 1120
rect 2363 1116 2364 1120
rect 2358 1115 2364 1116
rect 2518 1120 2524 1121
rect 2518 1116 2519 1120
rect 2523 1116 2524 1120
rect 2518 1115 2524 1116
rect 2678 1120 2684 1121
rect 2678 1116 2679 1120
rect 2683 1116 2684 1120
rect 2678 1115 2684 1116
rect 2830 1120 2836 1121
rect 2830 1116 2831 1120
rect 2835 1116 2836 1120
rect 2830 1115 2836 1116
rect 2974 1120 2980 1121
rect 2974 1116 2975 1120
rect 2979 1116 2980 1120
rect 2974 1115 2980 1116
rect 3118 1120 3124 1121
rect 3118 1116 3119 1120
rect 3123 1116 3124 1120
rect 3118 1115 3124 1116
rect 3254 1120 3260 1121
rect 3254 1116 3255 1120
rect 3259 1116 3260 1120
rect 3254 1115 3260 1116
rect 3390 1120 3396 1121
rect 3390 1116 3391 1120
rect 3395 1116 3396 1120
rect 3390 1115 3396 1116
rect 3502 1120 3508 1121
rect 3502 1116 3503 1120
rect 3507 1116 3508 1120
rect 3590 1119 3591 1123
rect 3595 1119 3596 1123
rect 3590 1118 3596 1119
rect 3502 1115 3508 1116
rect 1896 1091 1898 1115
rect 1976 1091 1978 1115
rect 2080 1091 2082 1115
rect 2208 1091 2210 1115
rect 2360 1091 2362 1115
rect 2520 1091 2522 1115
rect 2680 1091 2682 1115
rect 2832 1091 2834 1115
rect 2976 1091 2978 1115
rect 3120 1091 3122 1115
rect 3256 1091 3258 1115
rect 3392 1091 3394 1115
rect 3504 1091 3506 1115
rect 3592 1091 3594 1118
rect 1871 1090 1875 1091
rect 1871 1085 1875 1086
rect 1895 1090 1899 1091
rect 1895 1085 1899 1086
rect 1975 1090 1979 1091
rect 1975 1085 1979 1086
rect 2079 1090 2083 1091
rect 2079 1085 2083 1086
rect 2167 1090 2171 1091
rect 2167 1085 2171 1086
rect 2207 1090 2211 1091
rect 2207 1085 2211 1086
rect 2255 1090 2259 1091
rect 2255 1085 2259 1086
rect 2359 1090 2363 1091
rect 2359 1085 2363 1086
rect 2479 1090 2483 1091
rect 2479 1085 2483 1086
rect 2519 1090 2523 1091
rect 2519 1085 2523 1086
rect 2607 1090 2611 1091
rect 2607 1085 2611 1086
rect 2679 1090 2683 1091
rect 2679 1085 2683 1086
rect 2751 1090 2755 1091
rect 2751 1085 2755 1086
rect 2831 1090 2835 1091
rect 2831 1085 2835 1086
rect 2895 1090 2899 1091
rect 2895 1085 2899 1086
rect 2975 1090 2979 1091
rect 2975 1085 2979 1086
rect 3047 1090 3051 1091
rect 3047 1085 3051 1086
rect 3119 1090 3123 1091
rect 3119 1085 3123 1086
rect 3207 1090 3211 1091
rect 3207 1085 3211 1086
rect 3255 1090 3259 1091
rect 3255 1085 3259 1086
rect 3367 1090 3371 1091
rect 3367 1085 3371 1086
rect 3391 1090 3395 1091
rect 3391 1085 3395 1086
rect 3503 1090 3507 1091
rect 3503 1085 3507 1086
rect 3591 1090 3595 1091
rect 3591 1085 3595 1086
rect 110 1084 116 1085
rect 110 1080 111 1084
rect 115 1080 116 1084
rect 110 1079 116 1080
rect 1830 1084 1836 1085
rect 1830 1080 1831 1084
rect 1835 1080 1836 1084
rect 1830 1079 1836 1080
rect 112 1043 114 1079
rect 150 1066 156 1067
rect 150 1062 151 1066
rect 155 1062 156 1066
rect 150 1061 156 1062
rect 286 1066 292 1067
rect 286 1062 287 1066
rect 291 1062 292 1066
rect 286 1061 292 1062
rect 430 1066 436 1067
rect 430 1062 431 1066
rect 435 1062 436 1066
rect 430 1061 436 1062
rect 574 1066 580 1067
rect 574 1062 575 1066
rect 579 1062 580 1066
rect 574 1061 580 1062
rect 718 1066 724 1067
rect 718 1062 719 1066
rect 723 1062 724 1066
rect 718 1061 724 1062
rect 854 1066 860 1067
rect 854 1062 855 1066
rect 859 1062 860 1066
rect 854 1061 860 1062
rect 982 1066 988 1067
rect 982 1062 983 1066
rect 987 1062 988 1066
rect 982 1061 988 1062
rect 1110 1066 1116 1067
rect 1110 1062 1111 1066
rect 1115 1062 1116 1066
rect 1110 1061 1116 1062
rect 1230 1066 1236 1067
rect 1230 1062 1231 1066
rect 1235 1062 1236 1066
rect 1230 1061 1236 1062
rect 1350 1066 1356 1067
rect 1350 1062 1351 1066
rect 1355 1062 1356 1066
rect 1350 1061 1356 1062
rect 1478 1066 1484 1067
rect 1478 1062 1479 1066
rect 1483 1062 1484 1066
rect 1478 1061 1484 1062
rect 152 1043 154 1061
rect 288 1043 290 1061
rect 432 1043 434 1061
rect 576 1043 578 1061
rect 720 1043 722 1061
rect 856 1043 858 1061
rect 984 1043 986 1061
rect 1112 1043 1114 1061
rect 1232 1043 1234 1061
rect 1352 1043 1354 1061
rect 1480 1043 1482 1061
rect 1832 1043 1834 1079
rect 1872 1066 1874 1085
rect 2168 1069 2170 1085
rect 2256 1069 2258 1085
rect 2360 1069 2362 1085
rect 2480 1069 2482 1085
rect 2608 1069 2610 1085
rect 2752 1069 2754 1085
rect 2896 1069 2898 1085
rect 3048 1069 3050 1085
rect 3208 1069 3210 1085
rect 3368 1069 3370 1085
rect 3504 1069 3506 1085
rect 2166 1068 2172 1069
rect 1870 1065 1876 1066
rect 1870 1061 1871 1065
rect 1875 1061 1876 1065
rect 2166 1064 2167 1068
rect 2171 1064 2172 1068
rect 2166 1063 2172 1064
rect 2254 1068 2260 1069
rect 2254 1064 2255 1068
rect 2259 1064 2260 1068
rect 2254 1063 2260 1064
rect 2358 1068 2364 1069
rect 2358 1064 2359 1068
rect 2363 1064 2364 1068
rect 2358 1063 2364 1064
rect 2478 1068 2484 1069
rect 2478 1064 2479 1068
rect 2483 1064 2484 1068
rect 2478 1063 2484 1064
rect 2606 1068 2612 1069
rect 2606 1064 2607 1068
rect 2611 1064 2612 1068
rect 2606 1063 2612 1064
rect 2750 1068 2756 1069
rect 2750 1064 2751 1068
rect 2755 1064 2756 1068
rect 2750 1063 2756 1064
rect 2894 1068 2900 1069
rect 2894 1064 2895 1068
rect 2899 1064 2900 1068
rect 2894 1063 2900 1064
rect 3046 1068 3052 1069
rect 3046 1064 3047 1068
rect 3051 1064 3052 1068
rect 3046 1063 3052 1064
rect 3206 1068 3212 1069
rect 3206 1064 3207 1068
rect 3211 1064 3212 1068
rect 3206 1063 3212 1064
rect 3366 1068 3372 1069
rect 3366 1064 3367 1068
rect 3371 1064 3372 1068
rect 3366 1063 3372 1064
rect 3502 1068 3508 1069
rect 3502 1064 3503 1068
rect 3507 1064 3508 1068
rect 3592 1066 3594 1085
rect 3502 1063 3508 1064
rect 3590 1065 3596 1066
rect 1870 1060 1876 1061
rect 3590 1061 3591 1065
rect 3595 1061 3596 1065
rect 3590 1060 3596 1061
rect 1870 1048 1876 1049
rect 1870 1044 1871 1048
rect 1875 1044 1876 1048
rect 1870 1043 1876 1044
rect 3590 1048 3596 1049
rect 3590 1044 3591 1048
rect 3595 1044 3596 1048
rect 3590 1043 3596 1044
rect 111 1042 115 1043
rect 111 1037 115 1038
rect 143 1042 147 1043
rect 143 1037 147 1038
rect 151 1042 155 1043
rect 151 1037 155 1038
rect 263 1042 267 1043
rect 263 1037 267 1038
rect 287 1042 291 1043
rect 287 1037 291 1038
rect 407 1042 411 1043
rect 407 1037 411 1038
rect 431 1042 435 1043
rect 431 1037 435 1038
rect 551 1042 555 1043
rect 551 1037 555 1038
rect 575 1042 579 1043
rect 575 1037 579 1038
rect 687 1042 691 1043
rect 687 1037 691 1038
rect 719 1042 723 1043
rect 719 1037 723 1038
rect 807 1042 811 1043
rect 807 1037 811 1038
rect 855 1042 859 1043
rect 855 1037 859 1038
rect 927 1042 931 1043
rect 927 1037 931 1038
rect 983 1042 987 1043
rect 983 1037 987 1038
rect 1039 1042 1043 1043
rect 1039 1037 1043 1038
rect 1111 1042 1115 1043
rect 1111 1037 1115 1038
rect 1143 1042 1147 1043
rect 1143 1037 1147 1038
rect 1231 1042 1235 1043
rect 1231 1037 1235 1038
rect 1247 1042 1251 1043
rect 1247 1037 1251 1038
rect 1351 1042 1355 1043
rect 1351 1037 1355 1038
rect 1359 1042 1363 1043
rect 1359 1037 1363 1038
rect 1479 1042 1483 1043
rect 1479 1037 1483 1038
rect 1831 1042 1835 1043
rect 1831 1037 1835 1038
rect 112 1009 114 1037
rect 144 1027 146 1037
rect 264 1027 266 1037
rect 408 1027 410 1037
rect 552 1027 554 1037
rect 688 1027 690 1037
rect 808 1027 810 1037
rect 928 1027 930 1037
rect 1040 1027 1042 1037
rect 1144 1027 1146 1037
rect 1248 1027 1250 1037
rect 1360 1027 1362 1037
rect 142 1026 148 1027
rect 142 1022 143 1026
rect 147 1022 148 1026
rect 142 1021 148 1022
rect 262 1026 268 1027
rect 262 1022 263 1026
rect 267 1022 268 1026
rect 262 1021 268 1022
rect 406 1026 412 1027
rect 406 1022 407 1026
rect 411 1022 412 1026
rect 406 1021 412 1022
rect 550 1026 556 1027
rect 550 1022 551 1026
rect 555 1022 556 1026
rect 550 1021 556 1022
rect 686 1026 692 1027
rect 686 1022 687 1026
rect 691 1022 692 1026
rect 686 1021 692 1022
rect 806 1026 812 1027
rect 806 1022 807 1026
rect 811 1022 812 1026
rect 806 1021 812 1022
rect 926 1026 932 1027
rect 926 1022 927 1026
rect 931 1022 932 1026
rect 926 1021 932 1022
rect 1038 1026 1044 1027
rect 1038 1022 1039 1026
rect 1043 1022 1044 1026
rect 1038 1021 1044 1022
rect 1142 1026 1148 1027
rect 1142 1022 1143 1026
rect 1147 1022 1148 1026
rect 1142 1021 1148 1022
rect 1246 1026 1252 1027
rect 1246 1022 1247 1026
rect 1251 1022 1252 1026
rect 1246 1021 1252 1022
rect 1358 1026 1364 1027
rect 1358 1022 1359 1026
rect 1363 1022 1364 1026
rect 1358 1021 1364 1022
rect 1832 1009 1834 1037
rect 1872 1015 1874 1043
rect 2174 1030 2180 1031
rect 2174 1026 2175 1030
rect 2179 1026 2180 1030
rect 2174 1025 2180 1026
rect 2262 1030 2268 1031
rect 2262 1026 2263 1030
rect 2267 1026 2268 1030
rect 2262 1025 2268 1026
rect 2366 1030 2372 1031
rect 2366 1026 2367 1030
rect 2371 1026 2372 1030
rect 2366 1025 2372 1026
rect 2486 1030 2492 1031
rect 2486 1026 2487 1030
rect 2491 1026 2492 1030
rect 2486 1025 2492 1026
rect 2614 1030 2620 1031
rect 2614 1026 2615 1030
rect 2619 1026 2620 1030
rect 2614 1025 2620 1026
rect 2758 1030 2764 1031
rect 2758 1026 2759 1030
rect 2763 1026 2764 1030
rect 2758 1025 2764 1026
rect 2902 1030 2908 1031
rect 2902 1026 2903 1030
rect 2907 1026 2908 1030
rect 2902 1025 2908 1026
rect 3054 1030 3060 1031
rect 3054 1026 3055 1030
rect 3059 1026 3060 1030
rect 3054 1025 3060 1026
rect 3214 1030 3220 1031
rect 3214 1026 3215 1030
rect 3219 1026 3220 1030
rect 3214 1025 3220 1026
rect 3374 1030 3380 1031
rect 3374 1026 3375 1030
rect 3379 1026 3380 1030
rect 3374 1025 3380 1026
rect 3510 1030 3516 1031
rect 3510 1026 3511 1030
rect 3515 1026 3516 1030
rect 3510 1025 3516 1026
rect 2176 1015 2178 1025
rect 2264 1015 2266 1025
rect 2368 1015 2370 1025
rect 2488 1015 2490 1025
rect 2616 1015 2618 1025
rect 2760 1015 2762 1025
rect 2904 1015 2906 1025
rect 3056 1015 3058 1025
rect 3216 1015 3218 1025
rect 3376 1015 3378 1025
rect 3512 1015 3514 1025
rect 3592 1015 3594 1043
rect 1871 1014 1875 1015
rect 1871 1009 1875 1010
rect 2175 1014 2179 1015
rect 2175 1009 2179 1010
rect 2263 1014 2267 1015
rect 2263 1009 2267 1010
rect 2303 1014 2307 1015
rect 2303 1009 2307 1010
rect 2367 1014 2371 1015
rect 2367 1009 2371 1010
rect 2383 1014 2387 1015
rect 2383 1009 2387 1010
rect 2471 1014 2475 1015
rect 2471 1009 2475 1010
rect 2487 1014 2491 1015
rect 2487 1009 2491 1010
rect 2567 1014 2571 1015
rect 2567 1009 2571 1010
rect 2615 1014 2619 1015
rect 2615 1009 2619 1010
rect 2671 1014 2675 1015
rect 2671 1009 2675 1010
rect 2759 1014 2763 1015
rect 2759 1009 2763 1010
rect 2783 1014 2787 1015
rect 2783 1009 2787 1010
rect 2903 1014 2907 1015
rect 2903 1009 2907 1010
rect 2911 1014 2915 1015
rect 2911 1009 2915 1010
rect 3055 1014 3059 1015
rect 3055 1009 3059 1010
rect 3207 1014 3211 1015
rect 3207 1009 3211 1010
rect 3215 1014 3219 1015
rect 3215 1009 3219 1010
rect 3367 1014 3371 1015
rect 3367 1009 3371 1010
rect 3375 1014 3379 1015
rect 3375 1009 3379 1010
rect 3511 1014 3515 1015
rect 3511 1009 3515 1010
rect 3591 1014 3595 1015
rect 3591 1009 3595 1010
rect 110 1008 116 1009
rect 110 1004 111 1008
rect 115 1004 116 1008
rect 110 1003 116 1004
rect 1830 1008 1836 1009
rect 1830 1004 1831 1008
rect 1835 1004 1836 1008
rect 1830 1003 1836 1004
rect 110 991 116 992
rect 110 987 111 991
rect 115 987 116 991
rect 1830 991 1836 992
rect 110 986 116 987
rect 134 988 140 989
rect 112 959 114 986
rect 134 984 135 988
rect 139 984 140 988
rect 134 983 140 984
rect 254 988 260 989
rect 254 984 255 988
rect 259 984 260 988
rect 254 983 260 984
rect 398 988 404 989
rect 398 984 399 988
rect 403 984 404 988
rect 398 983 404 984
rect 542 988 548 989
rect 542 984 543 988
rect 547 984 548 988
rect 542 983 548 984
rect 678 988 684 989
rect 678 984 679 988
rect 683 984 684 988
rect 678 983 684 984
rect 798 988 804 989
rect 798 984 799 988
rect 803 984 804 988
rect 798 983 804 984
rect 918 988 924 989
rect 918 984 919 988
rect 923 984 924 988
rect 918 983 924 984
rect 1030 988 1036 989
rect 1030 984 1031 988
rect 1035 984 1036 988
rect 1030 983 1036 984
rect 1134 988 1140 989
rect 1134 984 1135 988
rect 1139 984 1140 988
rect 1134 983 1140 984
rect 1238 988 1244 989
rect 1238 984 1239 988
rect 1243 984 1244 988
rect 1238 983 1244 984
rect 1350 988 1356 989
rect 1350 984 1351 988
rect 1355 984 1356 988
rect 1830 987 1831 991
rect 1835 987 1836 991
rect 1830 986 1836 987
rect 1350 983 1356 984
rect 136 959 138 983
rect 256 959 258 983
rect 400 959 402 983
rect 544 959 546 983
rect 680 959 682 983
rect 800 959 802 983
rect 920 959 922 983
rect 1032 959 1034 983
rect 1136 959 1138 983
rect 1240 959 1242 983
rect 1352 959 1354 983
rect 1832 959 1834 986
rect 1872 981 1874 1009
rect 2304 999 2306 1009
rect 2384 999 2386 1009
rect 2472 999 2474 1009
rect 2568 999 2570 1009
rect 2672 999 2674 1009
rect 2784 999 2786 1009
rect 2912 999 2914 1009
rect 3056 999 3058 1009
rect 3208 999 3210 1009
rect 3368 999 3370 1009
rect 3512 999 3514 1009
rect 2302 998 2308 999
rect 2302 994 2303 998
rect 2307 994 2308 998
rect 2302 993 2308 994
rect 2382 998 2388 999
rect 2382 994 2383 998
rect 2387 994 2388 998
rect 2382 993 2388 994
rect 2470 998 2476 999
rect 2470 994 2471 998
rect 2475 994 2476 998
rect 2470 993 2476 994
rect 2566 998 2572 999
rect 2566 994 2567 998
rect 2571 994 2572 998
rect 2566 993 2572 994
rect 2670 998 2676 999
rect 2670 994 2671 998
rect 2675 994 2676 998
rect 2670 993 2676 994
rect 2782 998 2788 999
rect 2782 994 2783 998
rect 2787 994 2788 998
rect 2782 993 2788 994
rect 2910 998 2916 999
rect 2910 994 2911 998
rect 2915 994 2916 998
rect 2910 993 2916 994
rect 3054 998 3060 999
rect 3054 994 3055 998
rect 3059 994 3060 998
rect 3054 993 3060 994
rect 3206 998 3212 999
rect 3206 994 3207 998
rect 3211 994 3212 998
rect 3206 993 3212 994
rect 3366 998 3372 999
rect 3366 994 3367 998
rect 3371 994 3372 998
rect 3366 993 3372 994
rect 3510 998 3516 999
rect 3510 994 3511 998
rect 3515 994 3516 998
rect 3510 993 3516 994
rect 3592 981 3594 1009
rect 1870 980 1876 981
rect 1870 976 1871 980
rect 1875 976 1876 980
rect 1870 975 1876 976
rect 3590 980 3596 981
rect 3590 976 3591 980
rect 3595 976 3596 980
rect 3590 975 3596 976
rect 1870 963 1876 964
rect 1870 959 1871 963
rect 1875 959 1876 963
rect 3590 963 3596 964
rect 111 958 115 959
rect 111 953 115 954
rect 135 958 139 959
rect 135 953 139 954
rect 215 958 219 959
rect 215 953 219 954
rect 255 958 259 959
rect 255 953 259 954
rect 327 958 331 959
rect 327 953 331 954
rect 399 958 403 959
rect 399 953 403 954
rect 447 958 451 959
rect 447 953 451 954
rect 543 958 547 959
rect 543 953 547 954
rect 567 958 571 959
rect 567 953 571 954
rect 679 958 683 959
rect 679 953 683 954
rect 687 958 691 959
rect 687 953 691 954
rect 799 958 803 959
rect 799 953 803 954
rect 911 958 915 959
rect 911 953 915 954
rect 919 958 923 959
rect 919 953 923 954
rect 1015 958 1019 959
rect 1015 953 1019 954
rect 1031 958 1035 959
rect 1031 953 1035 954
rect 1119 958 1123 959
rect 1119 953 1123 954
rect 1135 958 1139 959
rect 1135 953 1139 954
rect 1223 958 1227 959
rect 1223 953 1227 954
rect 1239 958 1243 959
rect 1239 953 1243 954
rect 1327 958 1331 959
rect 1327 953 1331 954
rect 1351 958 1355 959
rect 1351 953 1355 954
rect 1831 958 1835 959
rect 1870 958 1876 959
rect 2294 960 2300 961
rect 1831 953 1835 954
rect 112 934 114 953
rect 136 937 138 953
rect 216 937 218 953
rect 328 937 330 953
rect 448 937 450 953
rect 568 937 570 953
rect 688 937 690 953
rect 800 937 802 953
rect 912 937 914 953
rect 1016 937 1018 953
rect 1120 937 1122 953
rect 1224 937 1226 953
rect 1328 937 1330 953
rect 134 936 140 937
rect 110 933 116 934
rect 110 929 111 933
rect 115 929 116 933
rect 134 932 135 936
rect 139 932 140 936
rect 134 931 140 932
rect 214 936 220 937
rect 214 932 215 936
rect 219 932 220 936
rect 214 931 220 932
rect 326 936 332 937
rect 326 932 327 936
rect 331 932 332 936
rect 326 931 332 932
rect 446 936 452 937
rect 446 932 447 936
rect 451 932 452 936
rect 446 931 452 932
rect 566 936 572 937
rect 566 932 567 936
rect 571 932 572 936
rect 566 931 572 932
rect 686 936 692 937
rect 686 932 687 936
rect 691 932 692 936
rect 686 931 692 932
rect 798 936 804 937
rect 798 932 799 936
rect 803 932 804 936
rect 798 931 804 932
rect 910 936 916 937
rect 910 932 911 936
rect 915 932 916 936
rect 910 931 916 932
rect 1014 936 1020 937
rect 1014 932 1015 936
rect 1019 932 1020 936
rect 1014 931 1020 932
rect 1118 936 1124 937
rect 1118 932 1119 936
rect 1123 932 1124 936
rect 1118 931 1124 932
rect 1222 936 1228 937
rect 1222 932 1223 936
rect 1227 932 1228 936
rect 1222 931 1228 932
rect 1326 936 1332 937
rect 1326 932 1327 936
rect 1331 932 1332 936
rect 1832 934 1834 953
rect 1326 931 1332 932
rect 1830 933 1836 934
rect 110 928 116 929
rect 1830 929 1831 933
rect 1835 929 1836 933
rect 1872 931 1874 958
rect 2294 956 2295 960
rect 2299 956 2300 960
rect 2294 955 2300 956
rect 2374 960 2380 961
rect 2374 956 2375 960
rect 2379 956 2380 960
rect 2374 955 2380 956
rect 2462 960 2468 961
rect 2462 956 2463 960
rect 2467 956 2468 960
rect 2462 955 2468 956
rect 2558 960 2564 961
rect 2558 956 2559 960
rect 2563 956 2564 960
rect 2558 955 2564 956
rect 2662 960 2668 961
rect 2662 956 2663 960
rect 2667 956 2668 960
rect 2662 955 2668 956
rect 2774 960 2780 961
rect 2774 956 2775 960
rect 2779 956 2780 960
rect 2774 955 2780 956
rect 2902 960 2908 961
rect 2902 956 2903 960
rect 2907 956 2908 960
rect 2902 955 2908 956
rect 3046 960 3052 961
rect 3046 956 3047 960
rect 3051 956 3052 960
rect 3046 955 3052 956
rect 3198 960 3204 961
rect 3198 956 3199 960
rect 3203 956 3204 960
rect 3198 955 3204 956
rect 3358 960 3364 961
rect 3358 956 3359 960
rect 3363 956 3364 960
rect 3358 955 3364 956
rect 3502 960 3508 961
rect 3502 956 3503 960
rect 3507 956 3508 960
rect 3590 959 3591 963
rect 3595 959 3596 963
rect 3590 958 3596 959
rect 3502 955 3508 956
rect 2296 931 2298 955
rect 2376 931 2378 955
rect 2464 931 2466 955
rect 2560 931 2562 955
rect 2664 931 2666 955
rect 2776 931 2778 955
rect 2904 931 2906 955
rect 3048 931 3050 955
rect 3200 931 3202 955
rect 3360 931 3362 955
rect 3504 931 3506 955
rect 3592 931 3594 958
rect 1830 928 1836 929
rect 1871 930 1875 931
rect 1871 925 1875 926
rect 2279 930 2283 931
rect 2279 925 2283 926
rect 2295 930 2299 931
rect 2295 925 2299 926
rect 2359 930 2363 931
rect 2359 925 2363 926
rect 2375 930 2379 931
rect 2375 925 2379 926
rect 2439 930 2443 931
rect 2439 925 2443 926
rect 2463 930 2467 931
rect 2463 925 2467 926
rect 2519 930 2523 931
rect 2519 925 2523 926
rect 2559 930 2563 931
rect 2559 925 2563 926
rect 2607 930 2611 931
rect 2607 925 2611 926
rect 2663 930 2667 931
rect 2663 925 2667 926
rect 2703 930 2707 931
rect 2703 925 2707 926
rect 2775 930 2779 931
rect 2775 925 2779 926
rect 2807 930 2811 931
rect 2807 925 2811 926
rect 2903 930 2907 931
rect 2903 925 2907 926
rect 2911 930 2915 931
rect 2911 925 2915 926
rect 3015 930 3019 931
rect 3015 925 3019 926
rect 3047 930 3051 931
rect 3047 925 3051 926
rect 3111 930 3115 931
rect 3111 925 3115 926
rect 3199 930 3203 931
rect 3199 925 3203 926
rect 3215 930 3219 931
rect 3215 925 3219 926
rect 3319 930 3323 931
rect 3319 925 3323 926
rect 3359 930 3363 931
rect 3359 925 3363 926
rect 3423 930 3427 931
rect 3423 925 3427 926
rect 3503 930 3507 931
rect 3503 925 3507 926
rect 3591 930 3595 931
rect 3591 925 3595 926
rect 110 916 116 917
rect 110 912 111 916
rect 115 912 116 916
rect 110 911 116 912
rect 1830 916 1836 917
rect 1830 912 1831 916
rect 1835 912 1836 916
rect 1830 911 1836 912
rect 112 875 114 911
rect 142 898 148 899
rect 142 894 143 898
rect 147 894 148 898
rect 142 893 148 894
rect 222 898 228 899
rect 222 894 223 898
rect 227 894 228 898
rect 222 893 228 894
rect 334 898 340 899
rect 334 894 335 898
rect 339 894 340 898
rect 334 893 340 894
rect 454 898 460 899
rect 454 894 455 898
rect 459 894 460 898
rect 454 893 460 894
rect 574 898 580 899
rect 574 894 575 898
rect 579 894 580 898
rect 574 893 580 894
rect 694 898 700 899
rect 694 894 695 898
rect 699 894 700 898
rect 694 893 700 894
rect 806 898 812 899
rect 806 894 807 898
rect 811 894 812 898
rect 806 893 812 894
rect 918 898 924 899
rect 918 894 919 898
rect 923 894 924 898
rect 918 893 924 894
rect 1022 898 1028 899
rect 1022 894 1023 898
rect 1027 894 1028 898
rect 1022 893 1028 894
rect 1126 898 1132 899
rect 1126 894 1127 898
rect 1131 894 1132 898
rect 1126 893 1132 894
rect 1230 898 1236 899
rect 1230 894 1231 898
rect 1235 894 1236 898
rect 1230 893 1236 894
rect 1334 898 1340 899
rect 1334 894 1335 898
rect 1339 894 1340 898
rect 1334 893 1340 894
rect 144 875 146 893
rect 224 875 226 893
rect 336 875 338 893
rect 456 875 458 893
rect 576 875 578 893
rect 696 875 698 893
rect 808 875 810 893
rect 920 875 922 893
rect 1024 875 1026 893
rect 1128 875 1130 893
rect 1232 875 1234 893
rect 1336 875 1338 893
rect 1832 875 1834 911
rect 1872 906 1874 925
rect 2280 909 2282 925
rect 2360 909 2362 925
rect 2440 909 2442 925
rect 2520 909 2522 925
rect 2608 909 2610 925
rect 2704 909 2706 925
rect 2808 909 2810 925
rect 2912 909 2914 925
rect 3016 909 3018 925
rect 3112 909 3114 925
rect 3216 909 3218 925
rect 3320 909 3322 925
rect 3424 909 3426 925
rect 3504 909 3506 925
rect 2278 908 2284 909
rect 1870 905 1876 906
rect 1870 901 1871 905
rect 1875 901 1876 905
rect 2278 904 2279 908
rect 2283 904 2284 908
rect 2278 903 2284 904
rect 2358 908 2364 909
rect 2358 904 2359 908
rect 2363 904 2364 908
rect 2358 903 2364 904
rect 2438 908 2444 909
rect 2438 904 2439 908
rect 2443 904 2444 908
rect 2438 903 2444 904
rect 2518 908 2524 909
rect 2518 904 2519 908
rect 2523 904 2524 908
rect 2518 903 2524 904
rect 2606 908 2612 909
rect 2606 904 2607 908
rect 2611 904 2612 908
rect 2606 903 2612 904
rect 2702 908 2708 909
rect 2702 904 2703 908
rect 2707 904 2708 908
rect 2702 903 2708 904
rect 2806 908 2812 909
rect 2806 904 2807 908
rect 2811 904 2812 908
rect 2806 903 2812 904
rect 2910 908 2916 909
rect 2910 904 2911 908
rect 2915 904 2916 908
rect 2910 903 2916 904
rect 3014 908 3020 909
rect 3014 904 3015 908
rect 3019 904 3020 908
rect 3014 903 3020 904
rect 3110 908 3116 909
rect 3110 904 3111 908
rect 3115 904 3116 908
rect 3110 903 3116 904
rect 3214 908 3220 909
rect 3214 904 3215 908
rect 3219 904 3220 908
rect 3214 903 3220 904
rect 3318 908 3324 909
rect 3318 904 3319 908
rect 3323 904 3324 908
rect 3318 903 3324 904
rect 3422 908 3428 909
rect 3422 904 3423 908
rect 3427 904 3428 908
rect 3422 903 3428 904
rect 3502 908 3508 909
rect 3502 904 3503 908
rect 3507 904 3508 908
rect 3592 906 3594 925
rect 3502 903 3508 904
rect 3590 905 3596 906
rect 1870 900 1876 901
rect 3590 901 3591 905
rect 3595 901 3596 905
rect 3590 900 3596 901
rect 1870 888 1876 889
rect 1870 884 1871 888
rect 1875 884 1876 888
rect 1870 883 1876 884
rect 3590 888 3596 889
rect 3590 884 3591 888
rect 3595 884 3596 888
rect 3590 883 3596 884
rect 111 874 115 875
rect 111 869 115 870
rect 143 874 147 875
rect 143 869 147 870
rect 223 874 227 875
rect 223 869 227 870
rect 255 874 259 875
rect 255 869 259 870
rect 335 874 339 875
rect 335 869 339 870
rect 399 874 403 875
rect 399 869 403 870
rect 455 874 459 875
rect 455 869 459 870
rect 559 874 563 875
rect 559 869 563 870
rect 575 874 579 875
rect 575 869 579 870
rect 695 874 699 875
rect 695 869 699 870
rect 719 874 723 875
rect 719 869 723 870
rect 807 874 811 875
rect 807 869 811 870
rect 871 874 875 875
rect 871 869 875 870
rect 919 874 923 875
rect 919 869 923 870
rect 1015 874 1019 875
rect 1015 869 1019 870
rect 1023 874 1027 875
rect 1023 869 1027 870
rect 1127 874 1131 875
rect 1127 869 1131 870
rect 1151 874 1155 875
rect 1151 869 1155 870
rect 1231 874 1235 875
rect 1231 869 1235 870
rect 1279 874 1283 875
rect 1279 869 1283 870
rect 1335 874 1339 875
rect 1335 869 1339 870
rect 1399 874 1403 875
rect 1399 869 1403 870
rect 1519 874 1523 875
rect 1519 869 1523 870
rect 1647 874 1651 875
rect 1647 869 1651 870
rect 1831 874 1835 875
rect 1831 869 1835 870
rect 112 841 114 869
rect 144 859 146 869
rect 256 859 258 869
rect 400 859 402 869
rect 560 859 562 869
rect 720 859 722 869
rect 872 859 874 869
rect 1016 859 1018 869
rect 1152 859 1154 869
rect 1280 859 1282 869
rect 1400 859 1402 869
rect 1520 859 1522 869
rect 1648 859 1650 869
rect 142 858 148 859
rect 142 854 143 858
rect 147 854 148 858
rect 142 853 148 854
rect 254 858 260 859
rect 254 854 255 858
rect 259 854 260 858
rect 254 853 260 854
rect 398 858 404 859
rect 398 854 399 858
rect 403 854 404 858
rect 398 853 404 854
rect 558 858 564 859
rect 558 854 559 858
rect 563 854 564 858
rect 558 853 564 854
rect 718 858 724 859
rect 718 854 719 858
rect 723 854 724 858
rect 718 853 724 854
rect 870 858 876 859
rect 870 854 871 858
rect 875 854 876 858
rect 870 853 876 854
rect 1014 858 1020 859
rect 1014 854 1015 858
rect 1019 854 1020 858
rect 1014 853 1020 854
rect 1150 858 1156 859
rect 1150 854 1151 858
rect 1155 854 1156 858
rect 1150 853 1156 854
rect 1278 858 1284 859
rect 1278 854 1279 858
rect 1283 854 1284 858
rect 1278 853 1284 854
rect 1398 858 1404 859
rect 1398 854 1399 858
rect 1403 854 1404 858
rect 1398 853 1404 854
rect 1518 858 1524 859
rect 1518 854 1519 858
rect 1523 854 1524 858
rect 1518 853 1524 854
rect 1646 858 1652 859
rect 1646 854 1647 858
rect 1651 854 1652 858
rect 1646 853 1652 854
rect 1832 841 1834 869
rect 1872 843 1874 883
rect 2286 870 2292 871
rect 2286 866 2287 870
rect 2291 866 2292 870
rect 2286 865 2292 866
rect 2366 870 2372 871
rect 2366 866 2367 870
rect 2371 866 2372 870
rect 2366 865 2372 866
rect 2446 870 2452 871
rect 2446 866 2447 870
rect 2451 866 2452 870
rect 2446 865 2452 866
rect 2526 870 2532 871
rect 2526 866 2527 870
rect 2531 866 2532 870
rect 2526 865 2532 866
rect 2614 870 2620 871
rect 2614 866 2615 870
rect 2619 866 2620 870
rect 2614 865 2620 866
rect 2710 870 2716 871
rect 2710 866 2711 870
rect 2715 866 2716 870
rect 2710 865 2716 866
rect 2814 870 2820 871
rect 2814 866 2815 870
rect 2819 866 2820 870
rect 2814 865 2820 866
rect 2918 870 2924 871
rect 2918 866 2919 870
rect 2923 866 2924 870
rect 2918 865 2924 866
rect 3022 870 3028 871
rect 3022 866 3023 870
rect 3027 866 3028 870
rect 3022 865 3028 866
rect 3118 870 3124 871
rect 3118 866 3119 870
rect 3123 866 3124 870
rect 3118 865 3124 866
rect 3222 870 3228 871
rect 3222 866 3223 870
rect 3227 866 3228 870
rect 3222 865 3228 866
rect 3326 870 3332 871
rect 3326 866 3327 870
rect 3331 866 3332 870
rect 3326 865 3332 866
rect 3430 870 3436 871
rect 3430 866 3431 870
rect 3435 866 3436 870
rect 3430 865 3436 866
rect 3510 870 3516 871
rect 3510 866 3511 870
rect 3515 866 3516 870
rect 3510 865 3516 866
rect 2288 843 2290 865
rect 2368 843 2370 865
rect 2448 843 2450 865
rect 2528 843 2530 865
rect 2616 843 2618 865
rect 2712 843 2714 865
rect 2816 843 2818 865
rect 2920 843 2922 865
rect 3024 843 3026 865
rect 3120 843 3122 865
rect 3224 843 3226 865
rect 3328 843 3330 865
rect 3432 843 3434 865
rect 3512 843 3514 865
rect 3592 843 3594 883
rect 1871 842 1875 843
rect 110 840 116 841
rect 110 836 111 840
rect 115 836 116 840
rect 110 835 116 836
rect 1830 840 1836 841
rect 1830 836 1831 840
rect 1835 836 1836 840
rect 1871 837 1875 838
rect 2167 842 2171 843
rect 2167 837 2171 838
rect 2247 842 2251 843
rect 2247 837 2251 838
rect 2287 842 2291 843
rect 2287 837 2291 838
rect 2327 842 2331 843
rect 2327 837 2331 838
rect 2367 842 2371 843
rect 2367 837 2371 838
rect 2423 842 2427 843
rect 2423 837 2427 838
rect 2447 842 2451 843
rect 2447 837 2451 838
rect 2527 842 2531 843
rect 2527 837 2531 838
rect 2535 842 2539 843
rect 2535 837 2539 838
rect 2615 842 2619 843
rect 2615 837 2619 838
rect 2655 842 2659 843
rect 2655 837 2659 838
rect 2711 842 2715 843
rect 2711 837 2715 838
rect 2783 842 2787 843
rect 2783 837 2787 838
rect 2815 842 2819 843
rect 2815 837 2819 838
rect 2911 842 2915 843
rect 2911 837 2915 838
rect 2919 842 2923 843
rect 2919 837 2923 838
rect 3023 842 3027 843
rect 3023 837 3027 838
rect 3039 842 3043 843
rect 3039 837 3043 838
rect 3119 842 3123 843
rect 3119 837 3123 838
rect 3159 842 3163 843
rect 3159 837 3163 838
rect 3223 842 3227 843
rect 3223 837 3227 838
rect 3279 842 3283 843
rect 3279 837 3283 838
rect 3327 842 3331 843
rect 3327 837 3331 838
rect 3407 842 3411 843
rect 3407 837 3411 838
rect 3431 842 3435 843
rect 3431 837 3435 838
rect 3511 842 3515 843
rect 3511 837 3515 838
rect 3591 842 3595 843
rect 3591 837 3595 838
rect 1830 835 1836 836
rect 110 823 116 824
rect 110 819 111 823
rect 115 819 116 823
rect 1830 823 1836 824
rect 110 818 116 819
rect 134 820 140 821
rect 112 787 114 818
rect 134 816 135 820
rect 139 816 140 820
rect 134 815 140 816
rect 246 820 252 821
rect 246 816 247 820
rect 251 816 252 820
rect 246 815 252 816
rect 390 820 396 821
rect 390 816 391 820
rect 395 816 396 820
rect 390 815 396 816
rect 550 820 556 821
rect 550 816 551 820
rect 555 816 556 820
rect 550 815 556 816
rect 710 820 716 821
rect 710 816 711 820
rect 715 816 716 820
rect 710 815 716 816
rect 862 820 868 821
rect 862 816 863 820
rect 867 816 868 820
rect 862 815 868 816
rect 1006 820 1012 821
rect 1006 816 1007 820
rect 1011 816 1012 820
rect 1006 815 1012 816
rect 1142 820 1148 821
rect 1142 816 1143 820
rect 1147 816 1148 820
rect 1142 815 1148 816
rect 1270 820 1276 821
rect 1270 816 1271 820
rect 1275 816 1276 820
rect 1270 815 1276 816
rect 1390 820 1396 821
rect 1390 816 1391 820
rect 1395 816 1396 820
rect 1390 815 1396 816
rect 1510 820 1516 821
rect 1510 816 1511 820
rect 1515 816 1516 820
rect 1510 815 1516 816
rect 1638 820 1644 821
rect 1638 816 1639 820
rect 1643 816 1644 820
rect 1830 819 1831 823
rect 1835 819 1836 823
rect 1830 818 1836 819
rect 1638 815 1644 816
rect 136 787 138 815
rect 248 787 250 815
rect 392 787 394 815
rect 552 787 554 815
rect 712 787 714 815
rect 864 787 866 815
rect 1008 787 1010 815
rect 1144 787 1146 815
rect 1272 787 1274 815
rect 1392 787 1394 815
rect 1512 787 1514 815
rect 1640 787 1642 815
rect 1832 787 1834 818
rect 1872 809 1874 837
rect 2168 827 2170 837
rect 2248 827 2250 837
rect 2328 827 2330 837
rect 2424 827 2426 837
rect 2536 827 2538 837
rect 2656 827 2658 837
rect 2784 827 2786 837
rect 2912 827 2914 837
rect 3040 827 3042 837
rect 3160 827 3162 837
rect 3280 827 3282 837
rect 3408 827 3410 837
rect 3512 827 3514 837
rect 2166 826 2172 827
rect 2166 822 2167 826
rect 2171 822 2172 826
rect 2166 821 2172 822
rect 2246 826 2252 827
rect 2246 822 2247 826
rect 2251 822 2252 826
rect 2246 821 2252 822
rect 2326 826 2332 827
rect 2326 822 2327 826
rect 2331 822 2332 826
rect 2326 821 2332 822
rect 2422 826 2428 827
rect 2422 822 2423 826
rect 2427 822 2428 826
rect 2422 821 2428 822
rect 2534 826 2540 827
rect 2534 822 2535 826
rect 2539 822 2540 826
rect 2534 821 2540 822
rect 2654 826 2660 827
rect 2654 822 2655 826
rect 2659 822 2660 826
rect 2654 821 2660 822
rect 2782 826 2788 827
rect 2782 822 2783 826
rect 2787 822 2788 826
rect 2782 821 2788 822
rect 2910 826 2916 827
rect 2910 822 2911 826
rect 2915 822 2916 826
rect 2910 821 2916 822
rect 3038 826 3044 827
rect 3038 822 3039 826
rect 3043 822 3044 826
rect 3038 821 3044 822
rect 3158 826 3164 827
rect 3158 822 3159 826
rect 3163 822 3164 826
rect 3158 821 3164 822
rect 3278 826 3284 827
rect 3278 822 3279 826
rect 3283 822 3284 826
rect 3278 821 3284 822
rect 3406 826 3412 827
rect 3406 822 3407 826
rect 3411 822 3412 826
rect 3406 821 3412 822
rect 3510 826 3516 827
rect 3510 822 3511 826
rect 3515 822 3516 826
rect 3510 821 3516 822
rect 3592 809 3594 837
rect 1870 808 1876 809
rect 1870 804 1871 808
rect 1875 804 1876 808
rect 1870 803 1876 804
rect 3590 808 3596 809
rect 3590 804 3591 808
rect 3595 804 3596 808
rect 3590 803 3596 804
rect 1870 791 1876 792
rect 1870 787 1871 791
rect 1875 787 1876 791
rect 3590 791 3596 792
rect 111 786 115 787
rect 111 781 115 782
rect 135 786 139 787
rect 135 781 139 782
rect 247 786 251 787
rect 247 781 251 782
rect 263 786 267 787
rect 263 781 267 782
rect 391 786 395 787
rect 391 781 395 782
rect 431 786 435 787
rect 431 781 435 782
rect 551 786 555 787
rect 551 781 555 782
rect 607 786 611 787
rect 607 781 611 782
rect 711 786 715 787
rect 711 781 715 782
rect 783 786 787 787
rect 783 781 787 782
rect 863 786 867 787
rect 863 781 867 782
rect 951 786 955 787
rect 951 781 955 782
rect 1007 786 1011 787
rect 1007 781 1011 782
rect 1103 786 1107 787
rect 1103 781 1107 782
rect 1143 786 1147 787
rect 1143 781 1147 782
rect 1247 786 1251 787
rect 1247 781 1251 782
rect 1271 786 1275 787
rect 1271 781 1275 782
rect 1383 786 1387 787
rect 1383 781 1387 782
rect 1391 786 1395 787
rect 1391 781 1395 782
rect 1511 786 1515 787
rect 1511 781 1515 782
rect 1639 786 1643 787
rect 1639 781 1643 782
rect 1743 786 1747 787
rect 1743 781 1747 782
rect 1831 786 1835 787
rect 1870 786 1876 787
rect 2158 788 2164 789
rect 1831 781 1835 782
rect 112 762 114 781
rect 136 765 138 781
rect 264 765 266 781
rect 432 765 434 781
rect 608 765 610 781
rect 784 765 786 781
rect 952 765 954 781
rect 1104 765 1106 781
rect 1248 765 1250 781
rect 1384 765 1386 781
rect 1512 765 1514 781
rect 1640 765 1642 781
rect 1744 765 1746 781
rect 134 764 140 765
rect 110 761 116 762
rect 110 757 111 761
rect 115 757 116 761
rect 134 760 135 764
rect 139 760 140 764
rect 134 759 140 760
rect 262 764 268 765
rect 262 760 263 764
rect 267 760 268 764
rect 262 759 268 760
rect 430 764 436 765
rect 430 760 431 764
rect 435 760 436 764
rect 430 759 436 760
rect 606 764 612 765
rect 606 760 607 764
rect 611 760 612 764
rect 606 759 612 760
rect 782 764 788 765
rect 782 760 783 764
rect 787 760 788 764
rect 782 759 788 760
rect 950 764 956 765
rect 950 760 951 764
rect 955 760 956 764
rect 950 759 956 760
rect 1102 764 1108 765
rect 1102 760 1103 764
rect 1107 760 1108 764
rect 1102 759 1108 760
rect 1246 764 1252 765
rect 1246 760 1247 764
rect 1251 760 1252 764
rect 1246 759 1252 760
rect 1382 764 1388 765
rect 1382 760 1383 764
rect 1387 760 1388 764
rect 1382 759 1388 760
rect 1510 764 1516 765
rect 1510 760 1511 764
rect 1515 760 1516 764
rect 1510 759 1516 760
rect 1638 764 1644 765
rect 1638 760 1639 764
rect 1643 760 1644 764
rect 1638 759 1644 760
rect 1742 764 1748 765
rect 1742 760 1743 764
rect 1747 760 1748 764
rect 1832 762 1834 781
rect 1742 759 1748 760
rect 1830 761 1836 762
rect 110 756 116 757
rect 1830 757 1831 761
rect 1835 757 1836 761
rect 1872 759 1874 786
rect 2158 784 2159 788
rect 2163 784 2164 788
rect 2158 783 2164 784
rect 2238 788 2244 789
rect 2238 784 2239 788
rect 2243 784 2244 788
rect 2238 783 2244 784
rect 2318 788 2324 789
rect 2318 784 2319 788
rect 2323 784 2324 788
rect 2318 783 2324 784
rect 2414 788 2420 789
rect 2414 784 2415 788
rect 2419 784 2420 788
rect 2414 783 2420 784
rect 2526 788 2532 789
rect 2526 784 2527 788
rect 2531 784 2532 788
rect 2526 783 2532 784
rect 2646 788 2652 789
rect 2646 784 2647 788
rect 2651 784 2652 788
rect 2646 783 2652 784
rect 2774 788 2780 789
rect 2774 784 2775 788
rect 2779 784 2780 788
rect 2774 783 2780 784
rect 2902 788 2908 789
rect 2902 784 2903 788
rect 2907 784 2908 788
rect 2902 783 2908 784
rect 3030 788 3036 789
rect 3030 784 3031 788
rect 3035 784 3036 788
rect 3030 783 3036 784
rect 3150 788 3156 789
rect 3150 784 3151 788
rect 3155 784 3156 788
rect 3150 783 3156 784
rect 3270 788 3276 789
rect 3270 784 3271 788
rect 3275 784 3276 788
rect 3270 783 3276 784
rect 3398 788 3404 789
rect 3398 784 3399 788
rect 3403 784 3404 788
rect 3398 783 3404 784
rect 3502 788 3508 789
rect 3502 784 3503 788
rect 3507 784 3508 788
rect 3590 787 3591 791
rect 3595 787 3596 791
rect 3590 786 3596 787
rect 3502 783 3508 784
rect 2160 759 2162 783
rect 2240 759 2242 783
rect 2320 759 2322 783
rect 2416 759 2418 783
rect 2528 759 2530 783
rect 2648 759 2650 783
rect 2776 759 2778 783
rect 2904 759 2906 783
rect 3032 759 3034 783
rect 3152 759 3154 783
rect 3272 759 3274 783
rect 3400 759 3402 783
rect 3504 759 3506 783
rect 3592 759 3594 786
rect 1830 756 1836 757
rect 1871 758 1875 759
rect 1871 753 1875 754
rect 1895 758 1899 759
rect 1895 753 1899 754
rect 1975 758 1979 759
rect 1975 753 1979 754
rect 2071 758 2075 759
rect 2071 753 2075 754
rect 2159 758 2163 759
rect 2159 753 2163 754
rect 2183 758 2187 759
rect 2183 753 2187 754
rect 2239 758 2243 759
rect 2239 753 2243 754
rect 2311 758 2315 759
rect 2311 753 2315 754
rect 2319 758 2323 759
rect 2319 753 2323 754
rect 2415 758 2419 759
rect 2415 753 2419 754
rect 2447 758 2451 759
rect 2447 753 2451 754
rect 2527 758 2531 759
rect 2527 753 2531 754
rect 2591 758 2595 759
rect 2591 753 2595 754
rect 2647 758 2651 759
rect 2647 753 2651 754
rect 2743 758 2747 759
rect 2743 753 2747 754
rect 2775 758 2779 759
rect 2775 753 2779 754
rect 2895 758 2899 759
rect 2895 753 2899 754
rect 2903 758 2907 759
rect 2903 753 2907 754
rect 3031 758 3035 759
rect 3031 753 3035 754
rect 3047 758 3051 759
rect 3047 753 3051 754
rect 3151 758 3155 759
rect 3151 753 3155 754
rect 3199 758 3203 759
rect 3199 753 3203 754
rect 3271 758 3275 759
rect 3271 753 3275 754
rect 3359 758 3363 759
rect 3359 753 3363 754
rect 3399 758 3403 759
rect 3399 753 3403 754
rect 3503 758 3507 759
rect 3503 753 3507 754
rect 3591 758 3595 759
rect 3591 753 3595 754
rect 110 744 116 745
rect 110 740 111 744
rect 115 740 116 744
rect 110 739 116 740
rect 1830 744 1836 745
rect 1830 740 1831 744
rect 1835 740 1836 744
rect 1830 739 1836 740
rect 112 699 114 739
rect 142 726 148 727
rect 142 722 143 726
rect 147 722 148 726
rect 142 721 148 722
rect 270 726 276 727
rect 270 722 271 726
rect 275 722 276 726
rect 270 721 276 722
rect 438 726 444 727
rect 438 722 439 726
rect 443 722 444 726
rect 438 721 444 722
rect 614 726 620 727
rect 614 722 615 726
rect 619 722 620 726
rect 614 721 620 722
rect 790 726 796 727
rect 790 722 791 726
rect 795 722 796 726
rect 790 721 796 722
rect 958 726 964 727
rect 958 722 959 726
rect 963 722 964 726
rect 958 721 964 722
rect 1110 726 1116 727
rect 1110 722 1111 726
rect 1115 722 1116 726
rect 1110 721 1116 722
rect 1254 726 1260 727
rect 1254 722 1255 726
rect 1259 722 1260 726
rect 1254 721 1260 722
rect 1390 726 1396 727
rect 1390 722 1391 726
rect 1395 722 1396 726
rect 1390 721 1396 722
rect 1518 726 1524 727
rect 1518 722 1519 726
rect 1523 722 1524 726
rect 1518 721 1524 722
rect 1646 726 1652 727
rect 1646 722 1647 726
rect 1651 722 1652 726
rect 1646 721 1652 722
rect 1750 726 1756 727
rect 1750 722 1751 726
rect 1755 722 1756 726
rect 1750 721 1756 722
rect 144 699 146 721
rect 272 699 274 721
rect 440 699 442 721
rect 616 699 618 721
rect 792 699 794 721
rect 960 699 962 721
rect 1112 699 1114 721
rect 1256 699 1258 721
rect 1392 699 1394 721
rect 1520 699 1522 721
rect 1648 699 1650 721
rect 1752 699 1754 721
rect 1832 699 1834 739
rect 1872 734 1874 753
rect 1896 737 1898 753
rect 1976 737 1978 753
rect 2072 737 2074 753
rect 2184 737 2186 753
rect 2312 737 2314 753
rect 2448 737 2450 753
rect 2592 737 2594 753
rect 2744 737 2746 753
rect 2896 737 2898 753
rect 3048 737 3050 753
rect 3200 737 3202 753
rect 3360 737 3362 753
rect 3504 737 3506 753
rect 1894 736 1900 737
rect 1870 733 1876 734
rect 1870 729 1871 733
rect 1875 729 1876 733
rect 1894 732 1895 736
rect 1899 732 1900 736
rect 1894 731 1900 732
rect 1974 736 1980 737
rect 1974 732 1975 736
rect 1979 732 1980 736
rect 1974 731 1980 732
rect 2070 736 2076 737
rect 2070 732 2071 736
rect 2075 732 2076 736
rect 2070 731 2076 732
rect 2182 736 2188 737
rect 2182 732 2183 736
rect 2187 732 2188 736
rect 2182 731 2188 732
rect 2310 736 2316 737
rect 2310 732 2311 736
rect 2315 732 2316 736
rect 2310 731 2316 732
rect 2446 736 2452 737
rect 2446 732 2447 736
rect 2451 732 2452 736
rect 2446 731 2452 732
rect 2590 736 2596 737
rect 2590 732 2591 736
rect 2595 732 2596 736
rect 2590 731 2596 732
rect 2742 736 2748 737
rect 2742 732 2743 736
rect 2747 732 2748 736
rect 2742 731 2748 732
rect 2894 736 2900 737
rect 2894 732 2895 736
rect 2899 732 2900 736
rect 2894 731 2900 732
rect 3046 736 3052 737
rect 3046 732 3047 736
rect 3051 732 3052 736
rect 3046 731 3052 732
rect 3198 736 3204 737
rect 3198 732 3199 736
rect 3203 732 3204 736
rect 3198 731 3204 732
rect 3358 736 3364 737
rect 3358 732 3359 736
rect 3363 732 3364 736
rect 3358 731 3364 732
rect 3502 736 3508 737
rect 3502 732 3503 736
rect 3507 732 3508 736
rect 3592 734 3594 753
rect 3502 731 3508 732
rect 3590 733 3596 734
rect 1870 728 1876 729
rect 3590 729 3591 733
rect 3595 729 3596 733
rect 3590 728 3596 729
rect 1870 716 1876 717
rect 1870 712 1871 716
rect 1875 712 1876 716
rect 1870 711 1876 712
rect 3590 716 3596 717
rect 3590 712 3591 716
rect 3595 712 3596 716
rect 3590 711 3596 712
rect 111 698 115 699
rect 111 693 115 694
rect 143 698 147 699
rect 143 693 147 694
rect 271 698 275 699
rect 271 693 275 694
rect 295 698 299 699
rect 295 693 299 694
rect 407 698 411 699
rect 407 693 411 694
rect 439 698 443 699
rect 439 693 443 694
rect 527 698 531 699
rect 527 693 531 694
rect 615 698 619 699
rect 615 693 619 694
rect 655 698 659 699
rect 655 693 659 694
rect 783 698 787 699
rect 783 693 787 694
rect 791 698 795 699
rect 791 693 795 694
rect 903 698 907 699
rect 903 693 907 694
rect 959 698 963 699
rect 959 693 963 694
rect 1023 698 1027 699
rect 1023 693 1027 694
rect 1111 698 1115 699
rect 1111 693 1115 694
rect 1135 698 1139 699
rect 1135 693 1139 694
rect 1247 698 1251 699
rect 1247 693 1251 694
rect 1255 698 1259 699
rect 1255 693 1259 694
rect 1351 698 1355 699
rect 1351 693 1355 694
rect 1391 698 1395 699
rect 1391 693 1395 694
rect 1455 698 1459 699
rect 1455 693 1459 694
rect 1519 698 1523 699
rect 1519 693 1523 694
rect 1559 698 1563 699
rect 1559 693 1563 694
rect 1647 698 1651 699
rect 1647 693 1651 694
rect 1663 698 1667 699
rect 1663 693 1667 694
rect 1751 698 1755 699
rect 1751 693 1755 694
rect 1831 698 1835 699
rect 1831 693 1835 694
rect 112 665 114 693
rect 296 683 298 693
rect 408 683 410 693
rect 528 683 530 693
rect 656 683 658 693
rect 784 683 786 693
rect 904 683 906 693
rect 1024 683 1026 693
rect 1136 683 1138 693
rect 1248 683 1250 693
rect 1352 683 1354 693
rect 1456 683 1458 693
rect 1560 683 1562 693
rect 1664 683 1666 693
rect 1752 683 1754 693
rect 294 682 300 683
rect 294 678 295 682
rect 299 678 300 682
rect 294 677 300 678
rect 406 682 412 683
rect 406 678 407 682
rect 411 678 412 682
rect 406 677 412 678
rect 526 682 532 683
rect 526 678 527 682
rect 531 678 532 682
rect 526 677 532 678
rect 654 682 660 683
rect 654 678 655 682
rect 659 678 660 682
rect 654 677 660 678
rect 782 682 788 683
rect 782 678 783 682
rect 787 678 788 682
rect 782 677 788 678
rect 902 682 908 683
rect 902 678 903 682
rect 907 678 908 682
rect 902 677 908 678
rect 1022 682 1028 683
rect 1022 678 1023 682
rect 1027 678 1028 682
rect 1022 677 1028 678
rect 1134 682 1140 683
rect 1134 678 1135 682
rect 1139 678 1140 682
rect 1134 677 1140 678
rect 1246 682 1252 683
rect 1246 678 1247 682
rect 1251 678 1252 682
rect 1246 677 1252 678
rect 1350 682 1356 683
rect 1350 678 1351 682
rect 1355 678 1356 682
rect 1350 677 1356 678
rect 1454 682 1460 683
rect 1454 678 1455 682
rect 1459 678 1460 682
rect 1454 677 1460 678
rect 1558 682 1564 683
rect 1558 678 1559 682
rect 1563 678 1564 682
rect 1558 677 1564 678
rect 1662 682 1668 683
rect 1662 678 1663 682
rect 1667 678 1668 682
rect 1662 677 1668 678
rect 1750 682 1756 683
rect 1750 678 1751 682
rect 1755 678 1756 682
rect 1750 677 1756 678
rect 1832 665 1834 693
rect 1872 679 1874 711
rect 1902 698 1908 699
rect 1902 694 1903 698
rect 1907 694 1908 698
rect 1902 693 1908 694
rect 1982 698 1988 699
rect 1982 694 1983 698
rect 1987 694 1988 698
rect 1982 693 1988 694
rect 2078 698 2084 699
rect 2078 694 2079 698
rect 2083 694 2084 698
rect 2078 693 2084 694
rect 2190 698 2196 699
rect 2190 694 2191 698
rect 2195 694 2196 698
rect 2190 693 2196 694
rect 2318 698 2324 699
rect 2318 694 2319 698
rect 2323 694 2324 698
rect 2318 693 2324 694
rect 2454 698 2460 699
rect 2454 694 2455 698
rect 2459 694 2460 698
rect 2454 693 2460 694
rect 2598 698 2604 699
rect 2598 694 2599 698
rect 2603 694 2604 698
rect 2598 693 2604 694
rect 2750 698 2756 699
rect 2750 694 2751 698
rect 2755 694 2756 698
rect 2750 693 2756 694
rect 2902 698 2908 699
rect 2902 694 2903 698
rect 2907 694 2908 698
rect 2902 693 2908 694
rect 3054 698 3060 699
rect 3054 694 3055 698
rect 3059 694 3060 698
rect 3054 693 3060 694
rect 3206 698 3212 699
rect 3206 694 3207 698
rect 3211 694 3212 698
rect 3206 693 3212 694
rect 3366 698 3372 699
rect 3366 694 3367 698
rect 3371 694 3372 698
rect 3366 693 3372 694
rect 3510 698 3516 699
rect 3510 694 3511 698
rect 3515 694 3516 698
rect 3510 693 3516 694
rect 1904 679 1906 693
rect 1984 679 1986 693
rect 2080 679 2082 693
rect 2192 679 2194 693
rect 2320 679 2322 693
rect 2456 679 2458 693
rect 2600 679 2602 693
rect 2752 679 2754 693
rect 2904 679 2906 693
rect 3056 679 3058 693
rect 3208 679 3210 693
rect 3368 679 3370 693
rect 3512 679 3514 693
rect 3592 679 3594 711
rect 1871 678 1875 679
rect 1871 673 1875 674
rect 1903 678 1907 679
rect 1903 673 1907 674
rect 1983 678 1987 679
rect 1983 673 1987 674
rect 2079 678 2083 679
rect 2079 673 2083 674
rect 2095 678 2099 679
rect 2095 673 2099 674
rect 2191 678 2195 679
rect 2191 673 2195 674
rect 2295 678 2299 679
rect 2295 673 2299 674
rect 2319 678 2323 679
rect 2319 673 2323 674
rect 2455 678 2459 679
rect 2455 673 2459 674
rect 2479 678 2483 679
rect 2479 673 2483 674
rect 2599 678 2603 679
rect 2599 673 2603 674
rect 2655 678 2659 679
rect 2655 673 2659 674
rect 2751 678 2755 679
rect 2751 673 2755 674
rect 2831 678 2835 679
rect 2831 673 2835 674
rect 2903 678 2907 679
rect 2903 673 2907 674
rect 3007 678 3011 679
rect 3007 673 3011 674
rect 3055 678 3059 679
rect 3055 673 3059 674
rect 3183 678 3187 679
rect 3183 673 3187 674
rect 3207 678 3211 679
rect 3207 673 3211 674
rect 3359 678 3363 679
rect 3359 673 3363 674
rect 3367 678 3371 679
rect 3367 673 3371 674
rect 3511 678 3515 679
rect 3511 673 3515 674
rect 3591 678 3595 679
rect 3591 673 3595 674
rect 110 664 116 665
rect 110 660 111 664
rect 115 660 116 664
rect 110 659 116 660
rect 1830 664 1836 665
rect 1830 660 1831 664
rect 1835 660 1836 664
rect 1830 659 1836 660
rect 110 647 116 648
rect 110 643 111 647
rect 115 643 116 647
rect 1830 647 1836 648
rect 110 642 116 643
rect 286 644 292 645
rect 112 619 114 642
rect 286 640 287 644
rect 291 640 292 644
rect 286 639 292 640
rect 398 644 404 645
rect 398 640 399 644
rect 403 640 404 644
rect 398 639 404 640
rect 518 644 524 645
rect 518 640 519 644
rect 523 640 524 644
rect 518 639 524 640
rect 646 644 652 645
rect 646 640 647 644
rect 651 640 652 644
rect 646 639 652 640
rect 774 644 780 645
rect 774 640 775 644
rect 779 640 780 644
rect 774 639 780 640
rect 894 644 900 645
rect 894 640 895 644
rect 899 640 900 644
rect 894 639 900 640
rect 1014 644 1020 645
rect 1014 640 1015 644
rect 1019 640 1020 644
rect 1014 639 1020 640
rect 1126 644 1132 645
rect 1126 640 1127 644
rect 1131 640 1132 644
rect 1126 639 1132 640
rect 1238 644 1244 645
rect 1238 640 1239 644
rect 1243 640 1244 644
rect 1238 639 1244 640
rect 1342 644 1348 645
rect 1342 640 1343 644
rect 1347 640 1348 644
rect 1342 639 1348 640
rect 1446 644 1452 645
rect 1446 640 1447 644
rect 1451 640 1452 644
rect 1446 639 1452 640
rect 1550 644 1556 645
rect 1550 640 1551 644
rect 1555 640 1556 644
rect 1550 639 1556 640
rect 1654 644 1660 645
rect 1654 640 1655 644
rect 1659 640 1660 644
rect 1654 639 1660 640
rect 1742 644 1748 645
rect 1742 640 1743 644
rect 1747 640 1748 644
rect 1830 643 1831 647
rect 1835 643 1836 647
rect 1872 645 1874 673
rect 1904 663 1906 673
rect 2096 663 2098 673
rect 2296 663 2298 673
rect 2480 663 2482 673
rect 2656 663 2658 673
rect 2832 663 2834 673
rect 3008 663 3010 673
rect 3184 663 3186 673
rect 3360 663 3362 673
rect 3512 663 3514 673
rect 1902 662 1908 663
rect 1902 658 1903 662
rect 1907 658 1908 662
rect 1902 657 1908 658
rect 2094 662 2100 663
rect 2094 658 2095 662
rect 2099 658 2100 662
rect 2094 657 2100 658
rect 2294 662 2300 663
rect 2294 658 2295 662
rect 2299 658 2300 662
rect 2294 657 2300 658
rect 2478 662 2484 663
rect 2478 658 2479 662
rect 2483 658 2484 662
rect 2478 657 2484 658
rect 2654 662 2660 663
rect 2654 658 2655 662
rect 2659 658 2660 662
rect 2654 657 2660 658
rect 2830 662 2836 663
rect 2830 658 2831 662
rect 2835 658 2836 662
rect 2830 657 2836 658
rect 3006 662 3012 663
rect 3006 658 3007 662
rect 3011 658 3012 662
rect 3006 657 3012 658
rect 3182 662 3188 663
rect 3182 658 3183 662
rect 3187 658 3188 662
rect 3182 657 3188 658
rect 3358 662 3364 663
rect 3358 658 3359 662
rect 3363 658 3364 662
rect 3358 657 3364 658
rect 3510 662 3516 663
rect 3510 658 3511 662
rect 3515 658 3516 662
rect 3510 657 3516 658
rect 3592 645 3594 673
rect 1830 642 1836 643
rect 1870 644 1876 645
rect 1742 639 1748 640
rect 288 619 290 639
rect 400 619 402 639
rect 520 619 522 639
rect 648 619 650 639
rect 776 619 778 639
rect 896 619 898 639
rect 1016 619 1018 639
rect 1128 619 1130 639
rect 1240 619 1242 639
rect 1344 619 1346 639
rect 1448 619 1450 639
rect 1552 619 1554 639
rect 1656 619 1658 639
rect 1744 619 1746 639
rect 1832 619 1834 642
rect 1870 640 1871 644
rect 1875 640 1876 644
rect 1870 639 1876 640
rect 3590 644 3596 645
rect 3590 640 3591 644
rect 3595 640 3596 644
rect 3590 639 3596 640
rect 1870 627 1876 628
rect 1870 623 1871 627
rect 1875 623 1876 627
rect 3590 627 3596 628
rect 1870 622 1876 623
rect 1894 624 1900 625
rect 111 618 115 619
rect 111 613 115 614
rect 287 618 291 619
rect 287 613 291 614
rect 311 618 315 619
rect 311 613 315 614
rect 391 618 395 619
rect 391 613 395 614
rect 399 618 403 619
rect 399 613 403 614
rect 471 618 475 619
rect 471 613 475 614
rect 519 618 523 619
rect 519 613 523 614
rect 559 618 563 619
rect 559 613 563 614
rect 647 618 651 619
rect 647 613 651 614
rect 735 618 739 619
rect 735 613 739 614
rect 775 618 779 619
rect 775 613 779 614
rect 823 618 827 619
rect 823 613 827 614
rect 895 618 899 619
rect 895 613 899 614
rect 911 618 915 619
rect 911 613 915 614
rect 999 618 1003 619
rect 999 613 1003 614
rect 1015 618 1019 619
rect 1015 613 1019 614
rect 1087 618 1091 619
rect 1087 613 1091 614
rect 1127 618 1131 619
rect 1127 613 1131 614
rect 1175 618 1179 619
rect 1175 613 1179 614
rect 1239 618 1243 619
rect 1239 613 1243 614
rect 1263 618 1267 619
rect 1263 613 1267 614
rect 1343 618 1347 619
rect 1343 613 1347 614
rect 1447 618 1451 619
rect 1447 613 1451 614
rect 1551 618 1555 619
rect 1551 613 1555 614
rect 1655 618 1659 619
rect 1655 613 1659 614
rect 1743 618 1747 619
rect 1743 613 1747 614
rect 1831 618 1835 619
rect 1831 613 1835 614
rect 112 594 114 613
rect 312 597 314 613
rect 392 597 394 613
rect 472 597 474 613
rect 560 597 562 613
rect 648 597 650 613
rect 736 597 738 613
rect 824 597 826 613
rect 912 597 914 613
rect 1000 597 1002 613
rect 1088 597 1090 613
rect 1176 597 1178 613
rect 1264 597 1266 613
rect 310 596 316 597
rect 110 593 116 594
rect 110 589 111 593
rect 115 589 116 593
rect 310 592 311 596
rect 315 592 316 596
rect 310 591 316 592
rect 390 596 396 597
rect 390 592 391 596
rect 395 592 396 596
rect 390 591 396 592
rect 470 596 476 597
rect 470 592 471 596
rect 475 592 476 596
rect 470 591 476 592
rect 558 596 564 597
rect 558 592 559 596
rect 563 592 564 596
rect 558 591 564 592
rect 646 596 652 597
rect 646 592 647 596
rect 651 592 652 596
rect 646 591 652 592
rect 734 596 740 597
rect 734 592 735 596
rect 739 592 740 596
rect 734 591 740 592
rect 822 596 828 597
rect 822 592 823 596
rect 827 592 828 596
rect 822 591 828 592
rect 910 596 916 597
rect 910 592 911 596
rect 915 592 916 596
rect 910 591 916 592
rect 998 596 1004 597
rect 998 592 999 596
rect 1003 592 1004 596
rect 998 591 1004 592
rect 1086 596 1092 597
rect 1086 592 1087 596
rect 1091 592 1092 596
rect 1086 591 1092 592
rect 1174 596 1180 597
rect 1174 592 1175 596
rect 1179 592 1180 596
rect 1174 591 1180 592
rect 1262 596 1268 597
rect 1262 592 1263 596
rect 1267 592 1268 596
rect 1832 594 1834 613
rect 1872 599 1874 622
rect 1894 620 1895 624
rect 1899 620 1900 624
rect 1894 619 1900 620
rect 2086 624 2092 625
rect 2086 620 2087 624
rect 2091 620 2092 624
rect 2086 619 2092 620
rect 2286 624 2292 625
rect 2286 620 2287 624
rect 2291 620 2292 624
rect 2286 619 2292 620
rect 2470 624 2476 625
rect 2470 620 2471 624
rect 2475 620 2476 624
rect 2470 619 2476 620
rect 2646 624 2652 625
rect 2646 620 2647 624
rect 2651 620 2652 624
rect 2646 619 2652 620
rect 2822 624 2828 625
rect 2822 620 2823 624
rect 2827 620 2828 624
rect 2822 619 2828 620
rect 2998 624 3004 625
rect 2998 620 2999 624
rect 3003 620 3004 624
rect 2998 619 3004 620
rect 3174 624 3180 625
rect 3174 620 3175 624
rect 3179 620 3180 624
rect 3174 619 3180 620
rect 3350 624 3356 625
rect 3350 620 3351 624
rect 3355 620 3356 624
rect 3350 619 3356 620
rect 3502 624 3508 625
rect 3502 620 3503 624
rect 3507 620 3508 624
rect 3590 623 3591 627
rect 3595 623 3596 627
rect 3590 622 3596 623
rect 3502 619 3508 620
rect 1896 599 1898 619
rect 2088 599 2090 619
rect 2288 599 2290 619
rect 2472 599 2474 619
rect 2648 599 2650 619
rect 2824 599 2826 619
rect 3000 599 3002 619
rect 3176 599 3178 619
rect 3352 599 3354 619
rect 3504 599 3506 619
rect 3592 599 3594 622
rect 1871 598 1875 599
rect 1262 591 1268 592
rect 1830 593 1836 594
rect 1871 593 1875 594
rect 1895 598 1899 599
rect 1895 593 1899 594
rect 1975 598 1979 599
rect 1975 593 1979 594
rect 2087 598 2091 599
rect 2087 593 2091 594
rect 2215 598 2219 599
rect 2215 593 2219 594
rect 2287 598 2291 599
rect 2287 593 2291 594
rect 2351 598 2355 599
rect 2351 593 2355 594
rect 2471 598 2475 599
rect 2471 593 2475 594
rect 2495 598 2499 599
rect 2495 593 2499 594
rect 2647 598 2651 599
rect 2647 593 2651 594
rect 2807 598 2811 599
rect 2807 593 2811 594
rect 2823 598 2827 599
rect 2823 593 2827 594
rect 2975 598 2979 599
rect 2975 593 2979 594
rect 2999 598 3003 599
rect 2999 593 3003 594
rect 3151 598 3155 599
rect 3151 593 3155 594
rect 3175 598 3179 599
rect 3175 593 3179 594
rect 3335 598 3339 599
rect 3335 593 3339 594
rect 3351 598 3355 599
rect 3351 593 3355 594
rect 3503 598 3507 599
rect 3503 593 3507 594
rect 3591 598 3595 599
rect 3591 593 3595 594
rect 110 588 116 589
rect 1830 589 1831 593
rect 1835 589 1836 593
rect 1830 588 1836 589
rect 110 576 116 577
rect 110 572 111 576
rect 115 572 116 576
rect 110 571 116 572
rect 1830 576 1836 577
rect 1830 572 1831 576
rect 1835 572 1836 576
rect 1872 574 1874 593
rect 1896 577 1898 593
rect 1976 577 1978 593
rect 2088 577 2090 593
rect 2216 577 2218 593
rect 2352 577 2354 593
rect 2496 577 2498 593
rect 2648 577 2650 593
rect 2808 577 2810 593
rect 2976 577 2978 593
rect 3152 577 3154 593
rect 3336 577 3338 593
rect 3504 577 3506 593
rect 1894 576 1900 577
rect 1830 571 1836 572
rect 1870 573 1876 574
rect 112 531 114 571
rect 318 558 324 559
rect 318 554 319 558
rect 323 554 324 558
rect 318 553 324 554
rect 398 558 404 559
rect 398 554 399 558
rect 403 554 404 558
rect 398 553 404 554
rect 478 558 484 559
rect 478 554 479 558
rect 483 554 484 558
rect 478 553 484 554
rect 566 558 572 559
rect 566 554 567 558
rect 571 554 572 558
rect 566 553 572 554
rect 654 558 660 559
rect 654 554 655 558
rect 659 554 660 558
rect 654 553 660 554
rect 742 558 748 559
rect 742 554 743 558
rect 747 554 748 558
rect 742 553 748 554
rect 830 558 836 559
rect 830 554 831 558
rect 835 554 836 558
rect 830 553 836 554
rect 918 558 924 559
rect 918 554 919 558
rect 923 554 924 558
rect 918 553 924 554
rect 1006 558 1012 559
rect 1006 554 1007 558
rect 1011 554 1012 558
rect 1006 553 1012 554
rect 1094 558 1100 559
rect 1094 554 1095 558
rect 1099 554 1100 558
rect 1094 553 1100 554
rect 1182 558 1188 559
rect 1182 554 1183 558
rect 1187 554 1188 558
rect 1182 553 1188 554
rect 1270 558 1276 559
rect 1270 554 1271 558
rect 1275 554 1276 558
rect 1270 553 1276 554
rect 320 531 322 553
rect 400 531 402 553
rect 480 531 482 553
rect 568 531 570 553
rect 656 531 658 553
rect 744 531 746 553
rect 832 531 834 553
rect 920 531 922 553
rect 1008 531 1010 553
rect 1096 531 1098 553
rect 1184 531 1186 553
rect 1272 531 1274 553
rect 1832 531 1834 571
rect 1870 569 1871 573
rect 1875 569 1876 573
rect 1894 572 1895 576
rect 1899 572 1900 576
rect 1894 571 1900 572
rect 1974 576 1980 577
rect 1974 572 1975 576
rect 1979 572 1980 576
rect 1974 571 1980 572
rect 2086 576 2092 577
rect 2086 572 2087 576
rect 2091 572 2092 576
rect 2086 571 2092 572
rect 2214 576 2220 577
rect 2214 572 2215 576
rect 2219 572 2220 576
rect 2214 571 2220 572
rect 2350 576 2356 577
rect 2350 572 2351 576
rect 2355 572 2356 576
rect 2350 571 2356 572
rect 2494 576 2500 577
rect 2494 572 2495 576
rect 2499 572 2500 576
rect 2494 571 2500 572
rect 2646 576 2652 577
rect 2646 572 2647 576
rect 2651 572 2652 576
rect 2646 571 2652 572
rect 2806 576 2812 577
rect 2806 572 2807 576
rect 2811 572 2812 576
rect 2806 571 2812 572
rect 2974 576 2980 577
rect 2974 572 2975 576
rect 2979 572 2980 576
rect 2974 571 2980 572
rect 3150 576 3156 577
rect 3150 572 3151 576
rect 3155 572 3156 576
rect 3150 571 3156 572
rect 3334 576 3340 577
rect 3334 572 3335 576
rect 3339 572 3340 576
rect 3334 571 3340 572
rect 3502 576 3508 577
rect 3502 572 3503 576
rect 3507 572 3508 576
rect 3592 574 3594 593
rect 3502 571 3508 572
rect 3590 573 3596 574
rect 1870 568 1876 569
rect 3590 569 3591 573
rect 3595 569 3596 573
rect 3590 568 3596 569
rect 1870 556 1876 557
rect 1870 552 1871 556
rect 1875 552 1876 556
rect 1870 551 1876 552
rect 3590 556 3596 557
rect 3590 552 3591 556
rect 3595 552 3596 556
rect 3590 551 3596 552
rect 111 530 115 531
rect 111 525 115 526
rect 239 530 243 531
rect 239 525 243 526
rect 319 530 323 531
rect 319 525 323 526
rect 343 530 347 531
rect 343 525 347 526
rect 399 530 403 531
rect 399 525 403 526
rect 439 530 443 531
rect 439 525 443 526
rect 479 530 483 531
rect 479 525 483 526
rect 535 530 539 531
rect 535 525 539 526
rect 567 530 571 531
rect 567 525 571 526
rect 631 530 635 531
rect 631 525 635 526
rect 655 530 659 531
rect 655 525 659 526
rect 719 530 723 531
rect 719 525 723 526
rect 743 530 747 531
rect 743 525 747 526
rect 807 530 811 531
rect 807 525 811 526
rect 831 530 835 531
rect 831 525 835 526
rect 895 530 899 531
rect 895 525 899 526
rect 919 530 923 531
rect 919 525 923 526
rect 983 530 987 531
rect 983 525 987 526
rect 1007 530 1011 531
rect 1007 525 1011 526
rect 1071 530 1075 531
rect 1071 525 1075 526
rect 1095 530 1099 531
rect 1095 525 1099 526
rect 1159 530 1163 531
rect 1159 525 1163 526
rect 1183 530 1187 531
rect 1183 525 1187 526
rect 1247 530 1251 531
rect 1247 525 1251 526
rect 1271 530 1275 531
rect 1271 525 1275 526
rect 1831 530 1835 531
rect 1831 525 1835 526
rect 112 497 114 525
rect 240 515 242 525
rect 344 515 346 525
rect 440 515 442 525
rect 536 515 538 525
rect 632 515 634 525
rect 720 515 722 525
rect 808 515 810 525
rect 896 515 898 525
rect 984 515 986 525
rect 1072 515 1074 525
rect 1160 515 1162 525
rect 1248 515 1250 525
rect 238 514 244 515
rect 238 510 239 514
rect 243 510 244 514
rect 238 509 244 510
rect 342 514 348 515
rect 342 510 343 514
rect 347 510 348 514
rect 342 509 348 510
rect 438 514 444 515
rect 438 510 439 514
rect 443 510 444 514
rect 438 509 444 510
rect 534 514 540 515
rect 534 510 535 514
rect 539 510 540 514
rect 534 509 540 510
rect 630 514 636 515
rect 630 510 631 514
rect 635 510 636 514
rect 630 509 636 510
rect 718 514 724 515
rect 718 510 719 514
rect 723 510 724 514
rect 718 509 724 510
rect 806 514 812 515
rect 806 510 807 514
rect 811 510 812 514
rect 806 509 812 510
rect 894 514 900 515
rect 894 510 895 514
rect 899 510 900 514
rect 894 509 900 510
rect 982 514 988 515
rect 982 510 983 514
rect 987 510 988 514
rect 982 509 988 510
rect 1070 514 1076 515
rect 1070 510 1071 514
rect 1075 510 1076 514
rect 1070 509 1076 510
rect 1158 514 1164 515
rect 1158 510 1159 514
rect 1163 510 1164 514
rect 1158 509 1164 510
rect 1246 514 1252 515
rect 1246 510 1247 514
rect 1251 510 1252 514
rect 1246 509 1252 510
rect 1832 497 1834 525
rect 1872 523 1874 551
rect 1902 538 1908 539
rect 1902 534 1903 538
rect 1907 534 1908 538
rect 1902 533 1908 534
rect 1982 538 1988 539
rect 1982 534 1983 538
rect 1987 534 1988 538
rect 1982 533 1988 534
rect 2094 538 2100 539
rect 2094 534 2095 538
rect 2099 534 2100 538
rect 2094 533 2100 534
rect 2222 538 2228 539
rect 2222 534 2223 538
rect 2227 534 2228 538
rect 2222 533 2228 534
rect 2358 538 2364 539
rect 2358 534 2359 538
rect 2363 534 2364 538
rect 2358 533 2364 534
rect 2502 538 2508 539
rect 2502 534 2503 538
rect 2507 534 2508 538
rect 2502 533 2508 534
rect 2654 538 2660 539
rect 2654 534 2655 538
rect 2659 534 2660 538
rect 2654 533 2660 534
rect 2814 538 2820 539
rect 2814 534 2815 538
rect 2819 534 2820 538
rect 2814 533 2820 534
rect 2982 538 2988 539
rect 2982 534 2983 538
rect 2987 534 2988 538
rect 2982 533 2988 534
rect 3158 538 3164 539
rect 3158 534 3159 538
rect 3163 534 3164 538
rect 3158 533 3164 534
rect 3342 538 3348 539
rect 3342 534 3343 538
rect 3347 534 3348 538
rect 3342 533 3348 534
rect 3510 538 3516 539
rect 3510 534 3511 538
rect 3515 534 3516 538
rect 3510 533 3516 534
rect 1904 523 1906 533
rect 1984 523 1986 533
rect 2096 523 2098 533
rect 2224 523 2226 533
rect 2360 523 2362 533
rect 2504 523 2506 533
rect 2656 523 2658 533
rect 2816 523 2818 533
rect 2984 523 2986 533
rect 3160 523 3162 533
rect 3344 523 3346 533
rect 3512 523 3514 533
rect 3592 523 3594 551
rect 1871 522 1875 523
rect 1871 517 1875 518
rect 1903 522 1907 523
rect 1903 517 1907 518
rect 1983 522 1987 523
rect 1983 517 1987 518
rect 2095 522 2099 523
rect 2095 517 2099 518
rect 2151 522 2155 523
rect 2151 517 2155 518
rect 2223 522 2227 523
rect 2223 517 2227 518
rect 2231 522 2235 523
rect 2231 517 2235 518
rect 2327 522 2331 523
rect 2327 517 2331 518
rect 2359 522 2363 523
rect 2359 517 2363 518
rect 2431 522 2435 523
rect 2431 517 2435 518
rect 2503 522 2507 523
rect 2503 517 2507 518
rect 2551 522 2555 523
rect 2551 517 2555 518
rect 2655 522 2659 523
rect 2655 517 2659 518
rect 2687 522 2691 523
rect 2687 517 2691 518
rect 2815 522 2819 523
rect 2815 517 2819 518
rect 2839 522 2843 523
rect 2839 517 2843 518
rect 2983 522 2987 523
rect 2983 517 2987 518
rect 2999 522 3003 523
rect 2999 517 3003 518
rect 3159 522 3163 523
rect 3159 517 3163 518
rect 3175 522 3179 523
rect 3175 517 3179 518
rect 3343 522 3347 523
rect 3343 517 3347 518
rect 3351 522 3355 523
rect 3351 517 3355 518
rect 3511 522 3515 523
rect 3511 517 3515 518
rect 3591 522 3595 523
rect 3591 517 3595 518
rect 110 496 116 497
rect 110 492 111 496
rect 115 492 116 496
rect 110 491 116 492
rect 1830 496 1836 497
rect 1830 492 1831 496
rect 1835 492 1836 496
rect 1830 491 1836 492
rect 1872 489 1874 517
rect 2152 507 2154 517
rect 2232 507 2234 517
rect 2328 507 2330 517
rect 2432 507 2434 517
rect 2552 507 2554 517
rect 2688 507 2690 517
rect 2840 507 2842 517
rect 3000 507 3002 517
rect 3176 507 3178 517
rect 3352 507 3354 517
rect 3512 507 3514 517
rect 2150 506 2156 507
rect 2150 502 2151 506
rect 2155 502 2156 506
rect 2150 501 2156 502
rect 2230 506 2236 507
rect 2230 502 2231 506
rect 2235 502 2236 506
rect 2230 501 2236 502
rect 2326 506 2332 507
rect 2326 502 2327 506
rect 2331 502 2332 506
rect 2326 501 2332 502
rect 2430 506 2436 507
rect 2430 502 2431 506
rect 2435 502 2436 506
rect 2430 501 2436 502
rect 2550 506 2556 507
rect 2550 502 2551 506
rect 2555 502 2556 506
rect 2550 501 2556 502
rect 2686 506 2692 507
rect 2686 502 2687 506
rect 2691 502 2692 506
rect 2686 501 2692 502
rect 2838 506 2844 507
rect 2838 502 2839 506
rect 2843 502 2844 506
rect 2838 501 2844 502
rect 2998 506 3004 507
rect 2998 502 2999 506
rect 3003 502 3004 506
rect 2998 501 3004 502
rect 3174 506 3180 507
rect 3174 502 3175 506
rect 3179 502 3180 506
rect 3174 501 3180 502
rect 3350 506 3356 507
rect 3350 502 3351 506
rect 3355 502 3356 506
rect 3350 501 3356 502
rect 3510 506 3516 507
rect 3510 502 3511 506
rect 3515 502 3516 506
rect 3510 501 3516 502
rect 3592 489 3594 517
rect 1870 488 1876 489
rect 1870 484 1871 488
rect 1875 484 1876 488
rect 1870 483 1876 484
rect 3590 488 3596 489
rect 3590 484 3591 488
rect 3595 484 3596 488
rect 3590 483 3596 484
rect 110 479 116 480
rect 110 475 111 479
rect 115 475 116 479
rect 1830 479 1836 480
rect 110 474 116 475
rect 230 476 236 477
rect 112 447 114 474
rect 230 472 231 476
rect 235 472 236 476
rect 230 471 236 472
rect 334 476 340 477
rect 334 472 335 476
rect 339 472 340 476
rect 334 471 340 472
rect 430 476 436 477
rect 430 472 431 476
rect 435 472 436 476
rect 430 471 436 472
rect 526 476 532 477
rect 526 472 527 476
rect 531 472 532 476
rect 526 471 532 472
rect 622 476 628 477
rect 622 472 623 476
rect 627 472 628 476
rect 622 471 628 472
rect 710 476 716 477
rect 710 472 711 476
rect 715 472 716 476
rect 710 471 716 472
rect 798 476 804 477
rect 798 472 799 476
rect 803 472 804 476
rect 798 471 804 472
rect 886 476 892 477
rect 886 472 887 476
rect 891 472 892 476
rect 886 471 892 472
rect 974 476 980 477
rect 974 472 975 476
rect 979 472 980 476
rect 974 471 980 472
rect 1062 476 1068 477
rect 1062 472 1063 476
rect 1067 472 1068 476
rect 1062 471 1068 472
rect 1150 476 1156 477
rect 1150 472 1151 476
rect 1155 472 1156 476
rect 1150 471 1156 472
rect 1238 476 1244 477
rect 1238 472 1239 476
rect 1243 472 1244 476
rect 1830 475 1831 479
rect 1835 475 1836 479
rect 1830 474 1836 475
rect 1238 471 1244 472
rect 232 447 234 471
rect 336 447 338 471
rect 432 447 434 471
rect 528 447 530 471
rect 624 447 626 471
rect 712 447 714 471
rect 800 447 802 471
rect 888 447 890 471
rect 976 447 978 471
rect 1064 447 1066 471
rect 1152 447 1154 471
rect 1240 447 1242 471
rect 1832 447 1834 474
rect 1870 471 1876 472
rect 1870 467 1871 471
rect 1875 467 1876 471
rect 3590 471 3596 472
rect 1870 466 1876 467
rect 2142 468 2148 469
rect 111 446 115 447
rect 111 441 115 442
rect 135 446 139 447
rect 135 441 139 442
rect 231 446 235 447
rect 231 441 235 442
rect 247 446 251 447
rect 247 441 251 442
rect 335 446 339 447
rect 335 441 339 442
rect 375 446 379 447
rect 375 441 379 442
rect 431 446 435 447
rect 431 441 435 442
rect 495 446 499 447
rect 495 441 499 442
rect 527 446 531 447
rect 527 441 531 442
rect 607 446 611 447
rect 607 441 611 442
rect 623 446 627 447
rect 623 441 627 442
rect 711 446 715 447
rect 711 441 715 442
rect 719 446 723 447
rect 719 441 723 442
rect 799 446 803 447
rect 799 441 803 442
rect 823 446 827 447
rect 823 441 827 442
rect 887 446 891 447
rect 887 441 891 442
rect 919 446 923 447
rect 919 441 923 442
rect 975 446 979 447
rect 975 441 979 442
rect 1007 446 1011 447
rect 1007 441 1011 442
rect 1063 446 1067 447
rect 1063 441 1067 442
rect 1103 446 1107 447
rect 1103 441 1107 442
rect 1151 446 1155 447
rect 1151 441 1155 442
rect 1199 446 1203 447
rect 1199 441 1203 442
rect 1239 446 1243 447
rect 1239 441 1243 442
rect 1295 446 1299 447
rect 1295 441 1299 442
rect 1831 446 1835 447
rect 1872 443 1874 466
rect 2142 464 2143 468
rect 2147 464 2148 468
rect 2142 463 2148 464
rect 2222 468 2228 469
rect 2222 464 2223 468
rect 2227 464 2228 468
rect 2222 463 2228 464
rect 2318 468 2324 469
rect 2318 464 2319 468
rect 2323 464 2324 468
rect 2318 463 2324 464
rect 2422 468 2428 469
rect 2422 464 2423 468
rect 2427 464 2428 468
rect 2422 463 2428 464
rect 2542 468 2548 469
rect 2542 464 2543 468
rect 2547 464 2548 468
rect 2542 463 2548 464
rect 2678 468 2684 469
rect 2678 464 2679 468
rect 2683 464 2684 468
rect 2678 463 2684 464
rect 2830 468 2836 469
rect 2830 464 2831 468
rect 2835 464 2836 468
rect 2830 463 2836 464
rect 2990 468 2996 469
rect 2990 464 2991 468
rect 2995 464 2996 468
rect 2990 463 2996 464
rect 3166 468 3172 469
rect 3166 464 3167 468
rect 3171 464 3172 468
rect 3166 463 3172 464
rect 3342 468 3348 469
rect 3342 464 3343 468
rect 3347 464 3348 468
rect 3342 463 3348 464
rect 3502 468 3508 469
rect 3502 464 3503 468
rect 3507 464 3508 468
rect 3590 467 3591 471
rect 3595 467 3596 471
rect 3590 466 3596 467
rect 3502 463 3508 464
rect 2144 443 2146 463
rect 2224 443 2226 463
rect 2320 443 2322 463
rect 2424 443 2426 463
rect 2544 443 2546 463
rect 2680 443 2682 463
rect 2832 443 2834 463
rect 2992 443 2994 463
rect 3168 443 3170 463
rect 3344 443 3346 463
rect 3504 443 3506 463
rect 3592 443 3594 466
rect 1831 441 1835 442
rect 1871 442 1875 443
rect 112 422 114 441
rect 136 425 138 441
rect 248 425 250 441
rect 376 425 378 441
rect 496 425 498 441
rect 608 425 610 441
rect 720 425 722 441
rect 824 425 826 441
rect 920 425 922 441
rect 1008 425 1010 441
rect 1104 425 1106 441
rect 1200 425 1202 441
rect 1296 425 1298 441
rect 134 424 140 425
rect 110 421 116 422
rect 110 417 111 421
rect 115 417 116 421
rect 134 420 135 424
rect 139 420 140 424
rect 134 419 140 420
rect 246 424 252 425
rect 246 420 247 424
rect 251 420 252 424
rect 246 419 252 420
rect 374 424 380 425
rect 374 420 375 424
rect 379 420 380 424
rect 374 419 380 420
rect 494 424 500 425
rect 494 420 495 424
rect 499 420 500 424
rect 494 419 500 420
rect 606 424 612 425
rect 606 420 607 424
rect 611 420 612 424
rect 606 419 612 420
rect 718 424 724 425
rect 718 420 719 424
rect 723 420 724 424
rect 718 419 724 420
rect 822 424 828 425
rect 822 420 823 424
rect 827 420 828 424
rect 822 419 828 420
rect 918 424 924 425
rect 918 420 919 424
rect 923 420 924 424
rect 918 419 924 420
rect 1006 424 1012 425
rect 1006 420 1007 424
rect 1011 420 1012 424
rect 1006 419 1012 420
rect 1102 424 1108 425
rect 1102 420 1103 424
rect 1107 420 1108 424
rect 1102 419 1108 420
rect 1198 424 1204 425
rect 1198 420 1199 424
rect 1203 420 1204 424
rect 1198 419 1204 420
rect 1294 424 1300 425
rect 1294 420 1295 424
rect 1299 420 1300 424
rect 1832 422 1834 441
rect 1871 437 1875 438
rect 2143 442 2147 443
rect 2143 437 2147 438
rect 2223 442 2227 443
rect 2223 437 2227 438
rect 2319 442 2323 443
rect 2319 437 2323 438
rect 2335 442 2339 443
rect 2335 437 2339 438
rect 2415 442 2419 443
rect 2415 437 2419 438
rect 2423 442 2427 443
rect 2423 437 2427 438
rect 2495 442 2499 443
rect 2495 437 2499 438
rect 2543 442 2547 443
rect 2543 437 2547 438
rect 2583 442 2587 443
rect 2583 437 2587 438
rect 2679 442 2683 443
rect 2679 437 2683 438
rect 2687 442 2691 443
rect 2687 437 2691 438
rect 2799 442 2803 443
rect 2799 437 2803 438
rect 2831 442 2835 443
rect 2831 437 2835 438
rect 2927 442 2931 443
rect 2927 437 2931 438
rect 2991 442 2995 443
rect 2991 437 2995 438
rect 3071 442 3075 443
rect 3071 437 3075 438
rect 3167 442 3171 443
rect 3167 437 3171 438
rect 3215 442 3219 443
rect 3215 437 3219 438
rect 3343 442 3347 443
rect 3343 437 3347 438
rect 3367 442 3371 443
rect 3367 437 3371 438
rect 3503 442 3507 443
rect 3503 437 3507 438
rect 3591 442 3595 443
rect 3591 437 3595 438
rect 1294 419 1300 420
rect 1830 421 1836 422
rect 110 416 116 417
rect 1830 417 1831 421
rect 1835 417 1836 421
rect 1872 418 1874 437
rect 2336 421 2338 437
rect 2416 421 2418 437
rect 2496 421 2498 437
rect 2584 421 2586 437
rect 2688 421 2690 437
rect 2800 421 2802 437
rect 2928 421 2930 437
rect 3072 421 3074 437
rect 3216 421 3218 437
rect 3368 421 3370 437
rect 3504 421 3506 437
rect 2334 420 2340 421
rect 1830 416 1836 417
rect 1870 417 1876 418
rect 1870 413 1871 417
rect 1875 413 1876 417
rect 2334 416 2335 420
rect 2339 416 2340 420
rect 2334 415 2340 416
rect 2414 420 2420 421
rect 2414 416 2415 420
rect 2419 416 2420 420
rect 2414 415 2420 416
rect 2494 420 2500 421
rect 2494 416 2495 420
rect 2499 416 2500 420
rect 2494 415 2500 416
rect 2582 420 2588 421
rect 2582 416 2583 420
rect 2587 416 2588 420
rect 2582 415 2588 416
rect 2686 420 2692 421
rect 2686 416 2687 420
rect 2691 416 2692 420
rect 2686 415 2692 416
rect 2798 420 2804 421
rect 2798 416 2799 420
rect 2803 416 2804 420
rect 2798 415 2804 416
rect 2926 420 2932 421
rect 2926 416 2927 420
rect 2931 416 2932 420
rect 2926 415 2932 416
rect 3070 420 3076 421
rect 3070 416 3071 420
rect 3075 416 3076 420
rect 3070 415 3076 416
rect 3214 420 3220 421
rect 3214 416 3215 420
rect 3219 416 3220 420
rect 3214 415 3220 416
rect 3366 420 3372 421
rect 3366 416 3367 420
rect 3371 416 3372 420
rect 3366 415 3372 416
rect 3502 420 3508 421
rect 3502 416 3503 420
rect 3507 416 3508 420
rect 3592 418 3594 437
rect 3502 415 3508 416
rect 3590 417 3596 418
rect 1870 412 1876 413
rect 3590 413 3591 417
rect 3595 413 3596 417
rect 3590 412 3596 413
rect 110 404 116 405
rect 110 400 111 404
rect 115 400 116 404
rect 110 399 116 400
rect 1830 404 1836 405
rect 1830 400 1831 404
rect 1835 400 1836 404
rect 1830 399 1836 400
rect 1870 400 1876 401
rect 112 359 114 399
rect 142 386 148 387
rect 142 382 143 386
rect 147 382 148 386
rect 142 381 148 382
rect 254 386 260 387
rect 254 382 255 386
rect 259 382 260 386
rect 254 381 260 382
rect 382 386 388 387
rect 382 382 383 386
rect 387 382 388 386
rect 382 381 388 382
rect 502 386 508 387
rect 502 382 503 386
rect 507 382 508 386
rect 502 381 508 382
rect 614 386 620 387
rect 614 382 615 386
rect 619 382 620 386
rect 614 381 620 382
rect 726 386 732 387
rect 726 382 727 386
rect 731 382 732 386
rect 726 381 732 382
rect 830 386 836 387
rect 830 382 831 386
rect 835 382 836 386
rect 830 381 836 382
rect 926 386 932 387
rect 926 382 927 386
rect 931 382 932 386
rect 926 381 932 382
rect 1014 386 1020 387
rect 1014 382 1015 386
rect 1019 382 1020 386
rect 1014 381 1020 382
rect 1110 386 1116 387
rect 1110 382 1111 386
rect 1115 382 1116 386
rect 1110 381 1116 382
rect 1206 386 1212 387
rect 1206 382 1207 386
rect 1211 382 1212 386
rect 1206 381 1212 382
rect 1302 386 1308 387
rect 1302 382 1303 386
rect 1307 382 1308 386
rect 1302 381 1308 382
rect 144 359 146 381
rect 256 359 258 381
rect 384 359 386 381
rect 504 359 506 381
rect 616 359 618 381
rect 728 359 730 381
rect 832 359 834 381
rect 928 359 930 381
rect 1016 359 1018 381
rect 1112 359 1114 381
rect 1208 359 1210 381
rect 1304 359 1306 381
rect 1832 359 1834 399
rect 1870 396 1871 400
rect 1875 396 1876 400
rect 1870 395 1876 396
rect 3590 400 3596 401
rect 3590 396 3591 400
rect 3595 396 3596 400
rect 3590 395 3596 396
rect 1872 359 1874 395
rect 2342 382 2348 383
rect 2342 378 2343 382
rect 2347 378 2348 382
rect 2342 377 2348 378
rect 2422 382 2428 383
rect 2422 378 2423 382
rect 2427 378 2428 382
rect 2422 377 2428 378
rect 2502 382 2508 383
rect 2502 378 2503 382
rect 2507 378 2508 382
rect 2502 377 2508 378
rect 2590 382 2596 383
rect 2590 378 2591 382
rect 2595 378 2596 382
rect 2590 377 2596 378
rect 2694 382 2700 383
rect 2694 378 2695 382
rect 2699 378 2700 382
rect 2694 377 2700 378
rect 2806 382 2812 383
rect 2806 378 2807 382
rect 2811 378 2812 382
rect 2806 377 2812 378
rect 2934 382 2940 383
rect 2934 378 2935 382
rect 2939 378 2940 382
rect 2934 377 2940 378
rect 3078 382 3084 383
rect 3078 378 3079 382
rect 3083 378 3084 382
rect 3078 377 3084 378
rect 3222 382 3228 383
rect 3222 378 3223 382
rect 3227 378 3228 382
rect 3222 377 3228 378
rect 3374 382 3380 383
rect 3374 378 3375 382
rect 3379 378 3380 382
rect 3374 377 3380 378
rect 3510 382 3516 383
rect 3510 378 3511 382
rect 3515 378 3516 382
rect 3510 377 3516 378
rect 2344 359 2346 377
rect 2424 359 2426 377
rect 2504 359 2506 377
rect 2592 359 2594 377
rect 2696 359 2698 377
rect 2808 359 2810 377
rect 2936 359 2938 377
rect 3080 359 3082 377
rect 3224 359 3226 377
rect 3376 359 3378 377
rect 3512 359 3514 377
rect 3592 359 3594 395
rect 111 358 115 359
rect 111 353 115 354
rect 143 358 147 359
rect 143 353 147 354
rect 247 358 251 359
rect 247 353 251 354
rect 255 358 259 359
rect 255 353 259 354
rect 375 358 379 359
rect 375 353 379 354
rect 383 358 387 359
rect 383 353 387 354
rect 503 358 507 359
rect 503 353 507 354
rect 511 358 515 359
rect 511 353 515 354
rect 615 358 619 359
rect 615 353 619 354
rect 647 358 651 359
rect 647 353 651 354
rect 727 358 731 359
rect 727 353 731 354
rect 775 358 779 359
rect 775 353 779 354
rect 831 358 835 359
rect 831 353 835 354
rect 895 358 899 359
rect 895 353 899 354
rect 927 358 931 359
rect 927 353 931 354
rect 1007 358 1011 359
rect 1007 353 1011 354
rect 1015 358 1019 359
rect 1015 353 1019 354
rect 1111 358 1115 359
rect 1111 353 1115 354
rect 1119 358 1123 359
rect 1119 353 1123 354
rect 1207 358 1211 359
rect 1207 353 1211 354
rect 1223 358 1227 359
rect 1223 353 1227 354
rect 1303 358 1307 359
rect 1303 353 1307 354
rect 1327 358 1331 359
rect 1327 353 1331 354
rect 1439 358 1443 359
rect 1439 353 1443 354
rect 1831 358 1835 359
rect 1831 353 1835 354
rect 1871 358 1875 359
rect 1871 353 1875 354
rect 2079 358 2083 359
rect 2079 353 2083 354
rect 2167 358 2171 359
rect 2167 353 2171 354
rect 2263 358 2267 359
rect 2263 353 2267 354
rect 2343 358 2347 359
rect 2343 353 2347 354
rect 2375 358 2379 359
rect 2375 353 2379 354
rect 2423 358 2427 359
rect 2423 353 2427 354
rect 2503 358 2507 359
rect 2503 353 2507 354
rect 2591 358 2595 359
rect 2591 353 2595 354
rect 2639 358 2643 359
rect 2639 353 2643 354
rect 2695 358 2699 359
rect 2695 353 2699 354
rect 2775 358 2779 359
rect 2775 353 2779 354
rect 2807 358 2811 359
rect 2807 353 2811 354
rect 2911 358 2915 359
rect 2911 353 2915 354
rect 2935 358 2939 359
rect 2935 353 2939 354
rect 3039 358 3043 359
rect 3039 353 3043 354
rect 3079 358 3083 359
rect 3079 353 3083 354
rect 3167 358 3171 359
rect 3167 353 3171 354
rect 3223 358 3227 359
rect 3223 353 3227 354
rect 3287 358 3291 359
rect 3287 353 3291 354
rect 3375 358 3379 359
rect 3375 353 3379 354
rect 3407 358 3411 359
rect 3407 353 3411 354
rect 3511 358 3515 359
rect 3511 353 3515 354
rect 3591 358 3595 359
rect 3591 353 3595 354
rect 112 325 114 353
rect 144 343 146 353
rect 248 343 250 353
rect 376 343 378 353
rect 512 343 514 353
rect 648 343 650 353
rect 776 343 778 353
rect 896 343 898 353
rect 1008 343 1010 353
rect 1120 343 1122 353
rect 1224 343 1226 353
rect 1328 343 1330 353
rect 1440 343 1442 353
rect 142 342 148 343
rect 142 338 143 342
rect 147 338 148 342
rect 142 337 148 338
rect 246 342 252 343
rect 246 338 247 342
rect 251 338 252 342
rect 246 337 252 338
rect 374 342 380 343
rect 374 338 375 342
rect 379 338 380 342
rect 374 337 380 338
rect 510 342 516 343
rect 510 338 511 342
rect 515 338 516 342
rect 510 337 516 338
rect 646 342 652 343
rect 646 338 647 342
rect 651 338 652 342
rect 646 337 652 338
rect 774 342 780 343
rect 774 338 775 342
rect 779 338 780 342
rect 774 337 780 338
rect 894 342 900 343
rect 894 338 895 342
rect 899 338 900 342
rect 894 337 900 338
rect 1006 342 1012 343
rect 1006 338 1007 342
rect 1011 338 1012 342
rect 1006 337 1012 338
rect 1118 342 1124 343
rect 1118 338 1119 342
rect 1123 338 1124 342
rect 1118 337 1124 338
rect 1222 342 1228 343
rect 1222 338 1223 342
rect 1227 338 1228 342
rect 1222 337 1228 338
rect 1326 342 1332 343
rect 1326 338 1327 342
rect 1331 338 1332 342
rect 1326 337 1332 338
rect 1438 342 1444 343
rect 1438 338 1439 342
rect 1443 338 1444 342
rect 1438 337 1444 338
rect 1832 325 1834 353
rect 1872 325 1874 353
rect 2080 343 2082 353
rect 2168 343 2170 353
rect 2264 343 2266 353
rect 2376 343 2378 353
rect 2504 343 2506 353
rect 2640 343 2642 353
rect 2776 343 2778 353
rect 2912 343 2914 353
rect 3040 343 3042 353
rect 3168 343 3170 353
rect 3288 343 3290 353
rect 3408 343 3410 353
rect 3512 343 3514 353
rect 2078 342 2084 343
rect 2078 338 2079 342
rect 2083 338 2084 342
rect 2078 337 2084 338
rect 2166 342 2172 343
rect 2166 338 2167 342
rect 2171 338 2172 342
rect 2166 337 2172 338
rect 2262 342 2268 343
rect 2262 338 2263 342
rect 2267 338 2268 342
rect 2262 337 2268 338
rect 2374 342 2380 343
rect 2374 338 2375 342
rect 2379 338 2380 342
rect 2374 337 2380 338
rect 2502 342 2508 343
rect 2502 338 2503 342
rect 2507 338 2508 342
rect 2502 337 2508 338
rect 2638 342 2644 343
rect 2638 338 2639 342
rect 2643 338 2644 342
rect 2638 337 2644 338
rect 2774 342 2780 343
rect 2774 338 2775 342
rect 2779 338 2780 342
rect 2774 337 2780 338
rect 2910 342 2916 343
rect 2910 338 2911 342
rect 2915 338 2916 342
rect 2910 337 2916 338
rect 3038 342 3044 343
rect 3038 338 3039 342
rect 3043 338 3044 342
rect 3038 337 3044 338
rect 3166 342 3172 343
rect 3166 338 3167 342
rect 3171 338 3172 342
rect 3166 337 3172 338
rect 3286 342 3292 343
rect 3286 338 3287 342
rect 3291 338 3292 342
rect 3286 337 3292 338
rect 3406 342 3412 343
rect 3406 338 3407 342
rect 3411 338 3412 342
rect 3406 337 3412 338
rect 3510 342 3516 343
rect 3510 338 3511 342
rect 3515 338 3516 342
rect 3510 337 3516 338
rect 3592 325 3594 353
rect 110 324 116 325
rect 110 320 111 324
rect 115 320 116 324
rect 110 319 116 320
rect 1830 324 1836 325
rect 1830 320 1831 324
rect 1835 320 1836 324
rect 1830 319 1836 320
rect 1870 324 1876 325
rect 1870 320 1871 324
rect 1875 320 1876 324
rect 1870 319 1876 320
rect 3590 324 3596 325
rect 3590 320 3591 324
rect 3595 320 3596 324
rect 3590 319 3596 320
rect 110 307 116 308
rect 110 303 111 307
rect 115 303 116 307
rect 1830 307 1836 308
rect 110 302 116 303
rect 134 304 140 305
rect 112 275 114 302
rect 134 300 135 304
rect 139 300 140 304
rect 134 299 140 300
rect 238 304 244 305
rect 238 300 239 304
rect 243 300 244 304
rect 238 299 244 300
rect 366 304 372 305
rect 366 300 367 304
rect 371 300 372 304
rect 366 299 372 300
rect 502 304 508 305
rect 502 300 503 304
rect 507 300 508 304
rect 502 299 508 300
rect 638 304 644 305
rect 638 300 639 304
rect 643 300 644 304
rect 638 299 644 300
rect 766 304 772 305
rect 766 300 767 304
rect 771 300 772 304
rect 766 299 772 300
rect 886 304 892 305
rect 886 300 887 304
rect 891 300 892 304
rect 886 299 892 300
rect 998 304 1004 305
rect 998 300 999 304
rect 1003 300 1004 304
rect 998 299 1004 300
rect 1110 304 1116 305
rect 1110 300 1111 304
rect 1115 300 1116 304
rect 1110 299 1116 300
rect 1214 304 1220 305
rect 1214 300 1215 304
rect 1219 300 1220 304
rect 1214 299 1220 300
rect 1318 304 1324 305
rect 1318 300 1319 304
rect 1323 300 1324 304
rect 1318 299 1324 300
rect 1430 304 1436 305
rect 1430 300 1431 304
rect 1435 300 1436 304
rect 1830 303 1831 307
rect 1835 303 1836 307
rect 1830 302 1836 303
rect 1870 307 1876 308
rect 1870 303 1871 307
rect 1875 303 1876 307
rect 3590 307 3596 308
rect 1870 302 1876 303
rect 2070 304 2076 305
rect 1430 299 1436 300
rect 136 275 138 299
rect 240 275 242 299
rect 368 275 370 299
rect 504 275 506 299
rect 640 275 642 299
rect 768 275 770 299
rect 888 275 890 299
rect 1000 275 1002 299
rect 1112 275 1114 299
rect 1216 275 1218 299
rect 1320 275 1322 299
rect 1432 275 1434 299
rect 1832 275 1834 302
rect 1872 275 1874 302
rect 2070 300 2071 304
rect 2075 300 2076 304
rect 2070 299 2076 300
rect 2158 304 2164 305
rect 2158 300 2159 304
rect 2163 300 2164 304
rect 2158 299 2164 300
rect 2254 304 2260 305
rect 2254 300 2255 304
rect 2259 300 2260 304
rect 2254 299 2260 300
rect 2366 304 2372 305
rect 2366 300 2367 304
rect 2371 300 2372 304
rect 2366 299 2372 300
rect 2494 304 2500 305
rect 2494 300 2495 304
rect 2499 300 2500 304
rect 2494 299 2500 300
rect 2630 304 2636 305
rect 2630 300 2631 304
rect 2635 300 2636 304
rect 2630 299 2636 300
rect 2766 304 2772 305
rect 2766 300 2767 304
rect 2771 300 2772 304
rect 2766 299 2772 300
rect 2902 304 2908 305
rect 2902 300 2903 304
rect 2907 300 2908 304
rect 2902 299 2908 300
rect 3030 304 3036 305
rect 3030 300 3031 304
rect 3035 300 3036 304
rect 3030 299 3036 300
rect 3158 304 3164 305
rect 3158 300 3159 304
rect 3163 300 3164 304
rect 3158 299 3164 300
rect 3278 304 3284 305
rect 3278 300 3279 304
rect 3283 300 3284 304
rect 3278 299 3284 300
rect 3398 304 3404 305
rect 3398 300 3399 304
rect 3403 300 3404 304
rect 3398 299 3404 300
rect 3502 304 3508 305
rect 3502 300 3503 304
rect 3507 300 3508 304
rect 3590 303 3591 307
rect 3595 303 3596 307
rect 3590 302 3596 303
rect 3502 299 3508 300
rect 2072 275 2074 299
rect 2160 275 2162 299
rect 2256 275 2258 299
rect 2368 275 2370 299
rect 2496 275 2498 299
rect 2632 275 2634 299
rect 2768 275 2770 299
rect 2904 275 2906 299
rect 3032 275 3034 299
rect 3160 275 3162 299
rect 3280 275 3282 299
rect 3400 275 3402 299
rect 3504 275 3506 299
rect 3592 275 3594 302
rect 111 274 115 275
rect 111 269 115 270
rect 135 274 139 275
rect 135 269 139 270
rect 223 274 227 275
rect 223 269 227 270
rect 239 274 243 275
rect 239 269 243 270
rect 335 274 339 275
rect 335 269 339 270
rect 367 274 371 275
rect 367 269 371 270
rect 463 274 467 275
rect 463 269 467 270
rect 503 274 507 275
rect 503 269 507 270
rect 599 274 603 275
rect 599 269 603 270
rect 639 274 643 275
rect 639 269 643 270
rect 735 274 739 275
rect 735 269 739 270
rect 767 274 771 275
rect 767 269 771 270
rect 871 274 875 275
rect 871 269 875 270
rect 887 274 891 275
rect 887 269 891 270
rect 999 274 1003 275
rect 999 269 1003 270
rect 1007 274 1011 275
rect 1007 269 1011 270
rect 1111 274 1115 275
rect 1111 269 1115 270
rect 1135 274 1139 275
rect 1135 269 1139 270
rect 1215 274 1219 275
rect 1215 269 1219 270
rect 1255 274 1259 275
rect 1255 269 1259 270
rect 1319 274 1323 275
rect 1319 269 1323 270
rect 1367 274 1371 275
rect 1367 269 1371 270
rect 1431 274 1435 275
rect 1431 269 1435 270
rect 1479 274 1483 275
rect 1479 269 1483 270
rect 1599 274 1603 275
rect 1599 269 1603 270
rect 1831 274 1835 275
rect 1831 269 1835 270
rect 1871 274 1875 275
rect 1871 269 1875 270
rect 1895 274 1899 275
rect 1895 269 1899 270
rect 1983 274 1987 275
rect 1983 269 1987 270
rect 2071 274 2075 275
rect 2071 269 2075 270
rect 2095 274 2099 275
rect 2095 269 2099 270
rect 2159 274 2163 275
rect 2159 269 2163 270
rect 2223 274 2227 275
rect 2223 269 2227 270
rect 2255 274 2259 275
rect 2255 269 2259 270
rect 2359 274 2363 275
rect 2359 269 2363 270
rect 2367 274 2371 275
rect 2367 269 2371 270
rect 2495 274 2499 275
rect 2495 269 2499 270
rect 2503 274 2507 275
rect 2503 269 2507 270
rect 2631 274 2635 275
rect 2631 269 2635 270
rect 2647 274 2651 275
rect 2647 269 2651 270
rect 2767 274 2771 275
rect 2767 269 2771 270
rect 2791 274 2795 275
rect 2791 269 2795 270
rect 2903 274 2907 275
rect 2903 269 2907 270
rect 2935 274 2939 275
rect 2935 269 2939 270
rect 3031 274 3035 275
rect 3031 269 3035 270
rect 3079 274 3083 275
rect 3079 269 3083 270
rect 3159 274 3163 275
rect 3159 269 3163 270
rect 3223 274 3227 275
rect 3223 269 3227 270
rect 3279 274 3283 275
rect 3279 269 3283 270
rect 3375 274 3379 275
rect 3375 269 3379 270
rect 3399 274 3403 275
rect 3399 269 3403 270
rect 3503 274 3507 275
rect 3503 269 3507 270
rect 3591 274 3595 275
rect 3591 269 3595 270
rect 112 250 114 269
rect 224 253 226 269
rect 336 253 338 269
rect 464 253 466 269
rect 600 253 602 269
rect 736 253 738 269
rect 872 253 874 269
rect 1008 253 1010 269
rect 1136 253 1138 269
rect 1256 253 1258 269
rect 1368 253 1370 269
rect 1480 253 1482 269
rect 1600 253 1602 269
rect 222 252 228 253
rect 110 249 116 250
rect 110 245 111 249
rect 115 245 116 249
rect 222 248 223 252
rect 227 248 228 252
rect 222 247 228 248
rect 334 252 340 253
rect 334 248 335 252
rect 339 248 340 252
rect 334 247 340 248
rect 462 252 468 253
rect 462 248 463 252
rect 467 248 468 252
rect 462 247 468 248
rect 598 252 604 253
rect 598 248 599 252
rect 603 248 604 252
rect 598 247 604 248
rect 734 252 740 253
rect 734 248 735 252
rect 739 248 740 252
rect 734 247 740 248
rect 870 252 876 253
rect 870 248 871 252
rect 875 248 876 252
rect 870 247 876 248
rect 1006 252 1012 253
rect 1006 248 1007 252
rect 1011 248 1012 252
rect 1006 247 1012 248
rect 1134 252 1140 253
rect 1134 248 1135 252
rect 1139 248 1140 252
rect 1134 247 1140 248
rect 1254 252 1260 253
rect 1254 248 1255 252
rect 1259 248 1260 252
rect 1254 247 1260 248
rect 1366 252 1372 253
rect 1366 248 1367 252
rect 1371 248 1372 252
rect 1366 247 1372 248
rect 1478 252 1484 253
rect 1478 248 1479 252
rect 1483 248 1484 252
rect 1478 247 1484 248
rect 1598 252 1604 253
rect 1598 248 1599 252
rect 1603 248 1604 252
rect 1832 250 1834 269
rect 1872 250 1874 269
rect 1896 253 1898 269
rect 1984 253 1986 269
rect 2096 253 2098 269
rect 2224 253 2226 269
rect 2360 253 2362 269
rect 2504 253 2506 269
rect 2648 253 2650 269
rect 2792 253 2794 269
rect 2936 253 2938 269
rect 3080 253 3082 269
rect 3224 253 3226 269
rect 3376 253 3378 269
rect 3504 253 3506 269
rect 1894 252 1900 253
rect 1598 247 1604 248
rect 1830 249 1836 250
rect 110 244 116 245
rect 1830 245 1831 249
rect 1835 245 1836 249
rect 1830 244 1836 245
rect 1870 249 1876 250
rect 1870 245 1871 249
rect 1875 245 1876 249
rect 1894 248 1895 252
rect 1899 248 1900 252
rect 1894 247 1900 248
rect 1982 252 1988 253
rect 1982 248 1983 252
rect 1987 248 1988 252
rect 1982 247 1988 248
rect 2094 252 2100 253
rect 2094 248 2095 252
rect 2099 248 2100 252
rect 2094 247 2100 248
rect 2222 252 2228 253
rect 2222 248 2223 252
rect 2227 248 2228 252
rect 2222 247 2228 248
rect 2358 252 2364 253
rect 2358 248 2359 252
rect 2363 248 2364 252
rect 2358 247 2364 248
rect 2502 252 2508 253
rect 2502 248 2503 252
rect 2507 248 2508 252
rect 2502 247 2508 248
rect 2646 252 2652 253
rect 2646 248 2647 252
rect 2651 248 2652 252
rect 2646 247 2652 248
rect 2790 252 2796 253
rect 2790 248 2791 252
rect 2795 248 2796 252
rect 2790 247 2796 248
rect 2934 252 2940 253
rect 2934 248 2935 252
rect 2939 248 2940 252
rect 2934 247 2940 248
rect 3078 252 3084 253
rect 3078 248 3079 252
rect 3083 248 3084 252
rect 3078 247 3084 248
rect 3222 252 3228 253
rect 3222 248 3223 252
rect 3227 248 3228 252
rect 3222 247 3228 248
rect 3374 252 3380 253
rect 3374 248 3375 252
rect 3379 248 3380 252
rect 3374 247 3380 248
rect 3502 252 3508 253
rect 3502 248 3503 252
rect 3507 248 3508 252
rect 3592 250 3594 269
rect 3502 247 3508 248
rect 3590 249 3596 250
rect 1870 244 1876 245
rect 3590 245 3591 249
rect 3595 245 3596 249
rect 3590 244 3596 245
rect 110 232 116 233
rect 110 228 111 232
rect 115 228 116 232
rect 110 227 116 228
rect 1830 232 1836 233
rect 1830 228 1831 232
rect 1835 228 1836 232
rect 1830 227 1836 228
rect 1870 232 1876 233
rect 1870 228 1871 232
rect 1875 228 1876 232
rect 1870 227 1876 228
rect 3590 232 3596 233
rect 3590 228 3591 232
rect 3595 228 3596 232
rect 3590 227 3596 228
rect 112 167 114 227
rect 230 214 236 215
rect 230 210 231 214
rect 235 210 236 214
rect 230 209 236 210
rect 342 214 348 215
rect 342 210 343 214
rect 347 210 348 214
rect 342 209 348 210
rect 470 214 476 215
rect 470 210 471 214
rect 475 210 476 214
rect 470 209 476 210
rect 606 214 612 215
rect 606 210 607 214
rect 611 210 612 214
rect 606 209 612 210
rect 742 214 748 215
rect 742 210 743 214
rect 747 210 748 214
rect 742 209 748 210
rect 878 214 884 215
rect 878 210 879 214
rect 883 210 884 214
rect 878 209 884 210
rect 1014 214 1020 215
rect 1014 210 1015 214
rect 1019 210 1020 214
rect 1014 209 1020 210
rect 1142 214 1148 215
rect 1142 210 1143 214
rect 1147 210 1148 214
rect 1142 209 1148 210
rect 1262 214 1268 215
rect 1262 210 1263 214
rect 1267 210 1268 214
rect 1262 209 1268 210
rect 1374 214 1380 215
rect 1374 210 1375 214
rect 1379 210 1380 214
rect 1374 209 1380 210
rect 1486 214 1492 215
rect 1486 210 1487 214
rect 1491 210 1492 214
rect 1486 209 1492 210
rect 1606 214 1612 215
rect 1606 210 1607 214
rect 1611 210 1612 214
rect 1606 209 1612 210
rect 232 167 234 209
rect 344 167 346 209
rect 472 167 474 209
rect 608 167 610 209
rect 744 167 746 209
rect 880 167 882 209
rect 1016 167 1018 209
rect 1144 167 1146 209
rect 1264 167 1266 209
rect 1376 167 1378 209
rect 1488 167 1490 209
rect 1608 167 1610 209
rect 1832 167 1834 227
rect 1872 187 1874 227
rect 1902 214 1908 215
rect 1902 210 1903 214
rect 1907 210 1908 214
rect 1902 209 1908 210
rect 1990 214 1996 215
rect 1990 210 1991 214
rect 1995 210 1996 214
rect 1990 209 1996 210
rect 2102 214 2108 215
rect 2102 210 2103 214
rect 2107 210 2108 214
rect 2102 209 2108 210
rect 2230 214 2236 215
rect 2230 210 2231 214
rect 2235 210 2236 214
rect 2230 209 2236 210
rect 2366 214 2372 215
rect 2366 210 2367 214
rect 2371 210 2372 214
rect 2366 209 2372 210
rect 2510 214 2516 215
rect 2510 210 2511 214
rect 2515 210 2516 214
rect 2510 209 2516 210
rect 2654 214 2660 215
rect 2654 210 2655 214
rect 2659 210 2660 214
rect 2654 209 2660 210
rect 2798 214 2804 215
rect 2798 210 2799 214
rect 2803 210 2804 214
rect 2798 209 2804 210
rect 2942 214 2948 215
rect 2942 210 2943 214
rect 2947 210 2948 214
rect 2942 209 2948 210
rect 3086 214 3092 215
rect 3086 210 3087 214
rect 3091 210 3092 214
rect 3086 209 3092 210
rect 3230 214 3236 215
rect 3230 210 3231 214
rect 3235 210 3236 214
rect 3230 209 3236 210
rect 3382 214 3388 215
rect 3382 210 3383 214
rect 3387 210 3388 214
rect 3382 209 3388 210
rect 3510 214 3516 215
rect 3510 210 3511 214
rect 3515 210 3516 214
rect 3510 209 3516 210
rect 1904 187 1906 209
rect 1992 187 1994 209
rect 2104 187 2106 209
rect 2232 187 2234 209
rect 2368 187 2370 209
rect 2512 187 2514 209
rect 2656 187 2658 209
rect 2800 187 2802 209
rect 2944 187 2946 209
rect 3088 187 3090 209
rect 3232 187 3234 209
rect 3384 187 3386 209
rect 3512 187 3514 209
rect 3592 187 3594 227
rect 1871 186 1875 187
rect 1871 181 1875 182
rect 1903 186 1907 187
rect 1903 181 1907 182
rect 1983 186 1987 187
rect 1983 181 1987 182
rect 1991 186 1995 187
rect 1991 181 1995 182
rect 2087 186 2091 187
rect 2087 181 2091 182
rect 2103 186 2107 187
rect 2103 181 2107 182
rect 2207 186 2211 187
rect 2207 181 2211 182
rect 2231 186 2235 187
rect 2231 181 2235 182
rect 2335 186 2339 187
rect 2335 181 2339 182
rect 2367 186 2371 187
rect 2367 181 2371 182
rect 2463 186 2467 187
rect 2463 181 2467 182
rect 2511 186 2515 187
rect 2511 181 2515 182
rect 2583 186 2587 187
rect 2583 181 2587 182
rect 2655 186 2659 187
rect 2655 181 2659 182
rect 2703 186 2707 187
rect 2703 181 2707 182
rect 2799 186 2803 187
rect 2799 181 2803 182
rect 2815 186 2819 187
rect 2815 181 2819 182
rect 2919 186 2923 187
rect 2919 181 2923 182
rect 2943 186 2947 187
rect 2943 181 2947 182
rect 3015 186 3019 187
rect 3015 181 3019 182
rect 3087 186 3091 187
rect 3087 181 3091 182
rect 3111 186 3115 187
rect 3111 181 3115 182
rect 3207 186 3211 187
rect 3207 181 3211 182
rect 3231 186 3235 187
rect 3231 181 3235 182
rect 3303 186 3307 187
rect 3303 181 3307 182
rect 3383 186 3387 187
rect 3383 181 3387 182
rect 3399 186 3403 187
rect 3399 181 3403 182
rect 3511 186 3515 187
rect 3511 181 3515 182
rect 3591 186 3595 187
rect 3591 181 3595 182
rect 111 166 115 167
rect 111 161 115 162
rect 159 166 163 167
rect 159 161 163 162
rect 231 166 235 167
rect 231 161 235 162
rect 239 166 243 167
rect 239 161 243 162
rect 319 166 323 167
rect 319 161 323 162
rect 343 166 347 167
rect 343 161 347 162
rect 399 166 403 167
rect 399 161 403 162
rect 471 166 475 167
rect 471 161 475 162
rect 479 166 483 167
rect 479 161 483 162
rect 559 166 563 167
rect 559 161 563 162
rect 607 166 611 167
rect 607 161 611 162
rect 647 166 651 167
rect 647 161 651 162
rect 735 166 739 167
rect 735 161 739 162
rect 743 166 747 167
rect 743 161 747 162
rect 823 166 827 167
rect 823 161 827 162
rect 879 166 883 167
rect 879 161 883 162
rect 911 166 915 167
rect 911 161 915 162
rect 999 166 1003 167
rect 999 161 1003 162
rect 1015 166 1019 167
rect 1015 161 1019 162
rect 1087 166 1091 167
rect 1087 161 1091 162
rect 1143 166 1147 167
rect 1143 161 1147 162
rect 1167 166 1171 167
rect 1167 161 1171 162
rect 1247 166 1251 167
rect 1247 161 1251 162
rect 1263 166 1267 167
rect 1263 161 1267 162
rect 1335 166 1339 167
rect 1335 161 1339 162
rect 1375 166 1379 167
rect 1375 161 1379 162
rect 1423 166 1427 167
rect 1423 161 1427 162
rect 1487 166 1491 167
rect 1487 161 1491 162
rect 1511 166 1515 167
rect 1511 161 1515 162
rect 1591 166 1595 167
rect 1591 161 1595 162
rect 1607 166 1611 167
rect 1607 161 1611 162
rect 1671 166 1675 167
rect 1671 161 1675 162
rect 1751 166 1755 167
rect 1751 161 1755 162
rect 1831 166 1835 167
rect 1831 161 1835 162
rect 112 133 114 161
rect 160 151 162 161
rect 240 151 242 161
rect 320 151 322 161
rect 400 151 402 161
rect 480 151 482 161
rect 560 151 562 161
rect 648 151 650 161
rect 736 151 738 161
rect 824 151 826 161
rect 912 151 914 161
rect 1000 151 1002 161
rect 1088 151 1090 161
rect 1168 151 1170 161
rect 1248 151 1250 161
rect 1336 151 1338 161
rect 1424 151 1426 161
rect 1512 151 1514 161
rect 1592 151 1594 161
rect 1672 151 1674 161
rect 1752 151 1754 161
rect 158 150 164 151
rect 158 146 159 150
rect 163 146 164 150
rect 158 145 164 146
rect 238 150 244 151
rect 238 146 239 150
rect 243 146 244 150
rect 238 145 244 146
rect 318 150 324 151
rect 318 146 319 150
rect 323 146 324 150
rect 318 145 324 146
rect 398 150 404 151
rect 398 146 399 150
rect 403 146 404 150
rect 398 145 404 146
rect 478 150 484 151
rect 478 146 479 150
rect 483 146 484 150
rect 478 145 484 146
rect 558 150 564 151
rect 558 146 559 150
rect 563 146 564 150
rect 558 145 564 146
rect 646 150 652 151
rect 646 146 647 150
rect 651 146 652 150
rect 646 145 652 146
rect 734 150 740 151
rect 734 146 735 150
rect 739 146 740 150
rect 734 145 740 146
rect 822 150 828 151
rect 822 146 823 150
rect 827 146 828 150
rect 822 145 828 146
rect 910 150 916 151
rect 910 146 911 150
rect 915 146 916 150
rect 910 145 916 146
rect 998 150 1004 151
rect 998 146 999 150
rect 1003 146 1004 150
rect 998 145 1004 146
rect 1086 150 1092 151
rect 1086 146 1087 150
rect 1091 146 1092 150
rect 1086 145 1092 146
rect 1166 150 1172 151
rect 1166 146 1167 150
rect 1171 146 1172 150
rect 1166 145 1172 146
rect 1246 150 1252 151
rect 1246 146 1247 150
rect 1251 146 1252 150
rect 1246 145 1252 146
rect 1334 150 1340 151
rect 1334 146 1335 150
rect 1339 146 1340 150
rect 1334 145 1340 146
rect 1422 150 1428 151
rect 1422 146 1423 150
rect 1427 146 1428 150
rect 1422 145 1428 146
rect 1510 150 1516 151
rect 1510 146 1511 150
rect 1515 146 1516 150
rect 1510 145 1516 146
rect 1590 150 1596 151
rect 1590 146 1591 150
rect 1595 146 1596 150
rect 1590 145 1596 146
rect 1670 150 1676 151
rect 1670 146 1671 150
rect 1675 146 1676 150
rect 1670 145 1676 146
rect 1750 150 1756 151
rect 1750 146 1751 150
rect 1755 146 1756 150
rect 1750 145 1756 146
rect 1832 133 1834 161
rect 1872 153 1874 181
rect 1904 171 1906 181
rect 1984 171 1986 181
rect 2088 171 2090 181
rect 2208 171 2210 181
rect 2336 171 2338 181
rect 2464 171 2466 181
rect 2584 171 2586 181
rect 2704 171 2706 181
rect 2816 171 2818 181
rect 2920 171 2922 181
rect 3016 171 3018 181
rect 3112 171 3114 181
rect 3208 171 3210 181
rect 3304 171 3306 181
rect 3400 171 3402 181
rect 1902 170 1908 171
rect 1902 166 1903 170
rect 1907 166 1908 170
rect 1902 165 1908 166
rect 1982 170 1988 171
rect 1982 166 1983 170
rect 1987 166 1988 170
rect 1982 165 1988 166
rect 2086 170 2092 171
rect 2086 166 2087 170
rect 2091 166 2092 170
rect 2086 165 2092 166
rect 2206 170 2212 171
rect 2206 166 2207 170
rect 2211 166 2212 170
rect 2206 165 2212 166
rect 2334 170 2340 171
rect 2334 166 2335 170
rect 2339 166 2340 170
rect 2334 165 2340 166
rect 2462 170 2468 171
rect 2462 166 2463 170
rect 2467 166 2468 170
rect 2462 165 2468 166
rect 2582 170 2588 171
rect 2582 166 2583 170
rect 2587 166 2588 170
rect 2582 165 2588 166
rect 2702 170 2708 171
rect 2702 166 2703 170
rect 2707 166 2708 170
rect 2702 165 2708 166
rect 2814 170 2820 171
rect 2814 166 2815 170
rect 2819 166 2820 170
rect 2814 165 2820 166
rect 2918 170 2924 171
rect 2918 166 2919 170
rect 2923 166 2924 170
rect 2918 165 2924 166
rect 3014 170 3020 171
rect 3014 166 3015 170
rect 3019 166 3020 170
rect 3014 165 3020 166
rect 3110 170 3116 171
rect 3110 166 3111 170
rect 3115 166 3116 170
rect 3110 165 3116 166
rect 3206 170 3212 171
rect 3206 166 3207 170
rect 3211 166 3212 170
rect 3206 165 3212 166
rect 3302 170 3308 171
rect 3302 166 3303 170
rect 3307 166 3308 170
rect 3302 165 3308 166
rect 3398 170 3404 171
rect 3398 166 3399 170
rect 3403 166 3404 170
rect 3398 165 3404 166
rect 3592 153 3594 181
rect 1870 152 1876 153
rect 1870 148 1871 152
rect 1875 148 1876 152
rect 1870 147 1876 148
rect 3590 152 3596 153
rect 3590 148 3591 152
rect 3595 148 3596 152
rect 3590 147 3596 148
rect 1870 135 1876 136
rect 110 132 116 133
rect 110 128 111 132
rect 115 128 116 132
rect 110 127 116 128
rect 1830 132 1836 133
rect 1830 128 1831 132
rect 1835 128 1836 132
rect 1870 131 1871 135
rect 1875 131 1876 135
rect 3590 135 3596 136
rect 1870 130 1876 131
rect 1894 132 1900 133
rect 1830 127 1836 128
rect 110 115 116 116
rect 110 111 111 115
rect 115 111 116 115
rect 1830 115 1836 116
rect 110 110 116 111
rect 150 112 156 113
rect 112 91 114 110
rect 150 108 151 112
rect 155 108 156 112
rect 150 107 156 108
rect 230 112 236 113
rect 230 108 231 112
rect 235 108 236 112
rect 230 107 236 108
rect 310 112 316 113
rect 310 108 311 112
rect 315 108 316 112
rect 310 107 316 108
rect 390 112 396 113
rect 390 108 391 112
rect 395 108 396 112
rect 390 107 396 108
rect 470 112 476 113
rect 470 108 471 112
rect 475 108 476 112
rect 470 107 476 108
rect 550 112 556 113
rect 550 108 551 112
rect 555 108 556 112
rect 550 107 556 108
rect 638 112 644 113
rect 638 108 639 112
rect 643 108 644 112
rect 638 107 644 108
rect 726 112 732 113
rect 726 108 727 112
rect 731 108 732 112
rect 726 107 732 108
rect 814 112 820 113
rect 814 108 815 112
rect 819 108 820 112
rect 814 107 820 108
rect 902 112 908 113
rect 902 108 903 112
rect 907 108 908 112
rect 902 107 908 108
rect 990 112 996 113
rect 990 108 991 112
rect 995 108 996 112
rect 990 107 996 108
rect 1078 112 1084 113
rect 1078 108 1079 112
rect 1083 108 1084 112
rect 1078 107 1084 108
rect 1158 112 1164 113
rect 1158 108 1159 112
rect 1163 108 1164 112
rect 1158 107 1164 108
rect 1238 112 1244 113
rect 1238 108 1239 112
rect 1243 108 1244 112
rect 1238 107 1244 108
rect 1326 112 1332 113
rect 1326 108 1327 112
rect 1331 108 1332 112
rect 1326 107 1332 108
rect 1414 112 1420 113
rect 1414 108 1415 112
rect 1419 108 1420 112
rect 1414 107 1420 108
rect 1502 112 1508 113
rect 1502 108 1503 112
rect 1507 108 1508 112
rect 1502 107 1508 108
rect 1582 112 1588 113
rect 1582 108 1583 112
rect 1587 108 1588 112
rect 1582 107 1588 108
rect 1662 112 1668 113
rect 1662 108 1663 112
rect 1667 108 1668 112
rect 1662 107 1668 108
rect 1742 112 1748 113
rect 1742 108 1743 112
rect 1747 108 1748 112
rect 1830 111 1831 115
rect 1835 111 1836 115
rect 1872 111 1874 130
rect 1894 128 1895 132
rect 1899 128 1900 132
rect 1894 127 1900 128
rect 1974 132 1980 133
rect 1974 128 1975 132
rect 1979 128 1980 132
rect 1974 127 1980 128
rect 2078 132 2084 133
rect 2078 128 2079 132
rect 2083 128 2084 132
rect 2078 127 2084 128
rect 2198 132 2204 133
rect 2198 128 2199 132
rect 2203 128 2204 132
rect 2198 127 2204 128
rect 2326 132 2332 133
rect 2326 128 2327 132
rect 2331 128 2332 132
rect 2326 127 2332 128
rect 2454 132 2460 133
rect 2454 128 2455 132
rect 2459 128 2460 132
rect 2454 127 2460 128
rect 2574 132 2580 133
rect 2574 128 2575 132
rect 2579 128 2580 132
rect 2574 127 2580 128
rect 2694 132 2700 133
rect 2694 128 2695 132
rect 2699 128 2700 132
rect 2694 127 2700 128
rect 2806 132 2812 133
rect 2806 128 2807 132
rect 2811 128 2812 132
rect 2806 127 2812 128
rect 2910 132 2916 133
rect 2910 128 2911 132
rect 2915 128 2916 132
rect 2910 127 2916 128
rect 3006 132 3012 133
rect 3006 128 3007 132
rect 3011 128 3012 132
rect 3006 127 3012 128
rect 3102 132 3108 133
rect 3102 128 3103 132
rect 3107 128 3108 132
rect 3102 127 3108 128
rect 3198 132 3204 133
rect 3198 128 3199 132
rect 3203 128 3204 132
rect 3198 127 3204 128
rect 3294 132 3300 133
rect 3294 128 3295 132
rect 3299 128 3300 132
rect 3294 127 3300 128
rect 3390 132 3396 133
rect 3390 128 3391 132
rect 3395 128 3396 132
rect 3590 131 3591 135
rect 3595 131 3596 135
rect 3590 130 3596 131
rect 3390 127 3396 128
rect 1896 111 1898 127
rect 1976 111 1978 127
rect 2080 111 2082 127
rect 2200 111 2202 127
rect 2328 111 2330 127
rect 2456 111 2458 127
rect 2576 111 2578 127
rect 2696 111 2698 127
rect 2808 111 2810 127
rect 2912 111 2914 127
rect 3008 111 3010 127
rect 3104 111 3106 127
rect 3200 111 3202 127
rect 3296 111 3298 127
rect 3392 111 3394 127
rect 3592 111 3594 130
rect 1830 110 1836 111
rect 1871 110 1875 111
rect 1742 107 1748 108
rect 152 91 154 107
rect 232 91 234 107
rect 312 91 314 107
rect 392 91 394 107
rect 472 91 474 107
rect 552 91 554 107
rect 640 91 642 107
rect 728 91 730 107
rect 816 91 818 107
rect 904 91 906 107
rect 992 91 994 107
rect 1080 91 1082 107
rect 1160 91 1162 107
rect 1240 91 1242 107
rect 1328 91 1330 107
rect 1416 91 1418 107
rect 1504 91 1506 107
rect 1584 91 1586 107
rect 1664 91 1666 107
rect 1744 91 1746 107
rect 1832 91 1834 110
rect 1871 105 1875 106
rect 1895 110 1899 111
rect 1895 105 1899 106
rect 1975 110 1979 111
rect 1975 105 1979 106
rect 2079 110 2083 111
rect 2079 105 2083 106
rect 2199 110 2203 111
rect 2199 105 2203 106
rect 2327 110 2331 111
rect 2327 105 2331 106
rect 2455 110 2459 111
rect 2455 105 2459 106
rect 2575 110 2579 111
rect 2575 105 2579 106
rect 2695 110 2699 111
rect 2695 105 2699 106
rect 2807 110 2811 111
rect 2807 105 2811 106
rect 2911 110 2915 111
rect 2911 105 2915 106
rect 3007 110 3011 111
rect 3007 105 3011 106
rect 3103 110 3107 111
rect 3103 105 3107 106
rect 3199 110 3203 111
rect 3199 105 3203 106
rect 3295 110 3299 111
rect 3295 105 3299 106
rect 3391 110 3395 111
rect 3391 105 3395 106
rect 3591 110 3595 111
rect 3591 105 3595 106
rect 111 90 115 91
rect 111 85 115 86
rect 151 90 155 91
rect 151 85 155 86
rect 231 90 235 91
rect 231 85 235 86
rect 311 90 315 91
rect 311 85 315 86
rect 391 90 395 91
rect 391 85 395 86
rect 471 90 475 91
rect 471 85 475 86
rect 551 90 555 91
rect 551 85 555 86
rect 639 90 643 91
rect 639 85 643 86
rect 727 90 731 91
rect 727 85 731 86
rect 815 90 819 91
rect 815 85 819 86
rect 903 90 907 91
rect 903 85 907 86
rect 991 90 995 91
rect 991 85 995 86
rect 1079 90 1083 91
rect 1079 85 1083 86
rect 1159 90 1163 91
rect 1159 85 1163 86
rect 1239 90 1243 91
rect 1239 85 1243 86
rect 1327 90 1331 91
rect 1327 85 1331 86
rect 1415 90 1419 91
rect 1415 85 1419 86
rect 1503 90 1507 91
rect 1503 85 1507 86
rect 1583 90 1587 91
rect 1583 85 1587 86
rect 1663 90 1667 91
rect 1663 85 1667 86
rect 1743 90 1747 91
rect 1743 85 1747 86
rect 1831 90 1835 91
rect 1831 85 1835 86
<< m4c >>
rect 1871 3666 1875 3670
rect 2151 3666 2155 3670
rect 2439 3666 2443 3670
rect 2727 3666 2731 3670
rect 3015 3666 3019 3670
rect 3591 3666 3595 3670
rect 111 3638 115 3642
rect 143 3638 147 3642
rect 239 3638 243 3642
rect 367 3638 371 3642
rect 503 3638 507 3642
rect 639 3638 643 3642
rect 775 3638 779 3642
rect 911 3638 915 3642
rect 1055 3638 1059 3642
rect 1199 3638 1203 3642
rect 1831 3638 1835 3642
rect 1871 3590 1875 3594
rect 1903 3590 1907 3594
rect 1983 3590 1987 3594
rect 2071 3590 2075 3594
rect 2159 3590 2163 3594
rect 2175 3590 2179 3594
rect 2295 3590 2299 3594
rect 2423 3590 2427 3594
rect 2447 3590 2451 3594
rect 2559 3590 2563 3594
rect 2695 3590 2699 3594
rect 2735 3590 2739 3594
rect 2831 3590 2835 3594
rect 2975 3590 2979 3594
rect 3023 3590 3027 3594
rect 3119 3590 3123 3594
rect 3263 3590 3267 3594
rect 3591 3590 3595 3594
rect 111 3562 115 3566
rect 135 3562 139 3566
rect 183 3562 187 3566
rect 231 3562 235 3566
rect 303 3562 307 3566
rect 359 3562 363 3566
rect 415 3562 419 3566
rect 495 3562 499 3566
rect 527 3562 531 3566
rect 631 3562 635 3566
rect 735 3562 739 3566
rect 767 3562 771 3566
rect 831 3562 835 3566
rect 903 3562 907 3566
rect 919 3562 923 3566
rect 1007 3562 1011 3566
rect 1047 3562 1051 3566
rect 1095 3562 1099 3566
rect 1183 3562 1187 3566
rect 1191 3562 1195 3566
rect 1271 3562 1275 3566
rect 1359 3562 1363 3566
rect 1447 3562 1451 3566
rect 1831 3562 1835 3566
rect 1871 3514 1875 3518
rect 1895 3514 1899 3518
rect 1967 3514 1971 3518
rect 1975 3514 1979 3518
rect 2063 3514 2067 3518
rect 2151 3514 2155 3518
rect 2167 3514 2171 3518
rect 2287 3514 2291 3518
rect 2335 3514 2339 3518
rect 2415 3514 2419 3518
rect 2511 3514 2515 3518
rect 2551 3514 2555 3518
rect 2671 3514 2675 3518
rect 2687 3514 2691 3518
rect 2823 3514 2827 3518
rect 2959 3514 2963 3518
rect 2967 3514 2971 3518
rect 3079 3514 3083 3518
rect 3111 3514 3115 3518
rect 3191 3514 3195 3518
rect 3255 3514 3259 3518
rect 3303 3514 3307 3518
rect 3415 3514 3419 3518
rect 3503 3514 3507 3518
rect 3591 3514 3595 3518
rect 111 3478 115 3482
rect 191 3478 195 3482
rect 231 3478 235 3482
rect 311 3478 315 3482
rect 367 3478 371 3482
rect 423 3478 427 3482
rect 503 3478 507 3482
rect 535 3478 539 3482
rect 623 3478 627 3482
rect 639 3478 643 3482
rect 735 3478 739 3482
rect 743 3478 747 3482
rect 839 3478 843 3482
rect 927 3478 931 3482
rect 943 3478 947 3482
rect 1015 3478 1019 3482
rect 1039 3478 1043 3482
rect 1103 3478 1107 3482
rect 1135 3478 1139 3482
rect 1191 3478 1195 3482
rect 1231 3478 1235 3482
rect 1279 3478 1283 3482
rect 1327 3478 1331 3482
rect 1367 3478 1371 3482
rect 1455 3478 1459 3482
rect 1831 3478 1835 3482
rect 1871 3438 1875 3442
rect 1975 3438 1979 3442
rect 2007 3438 2011 3442
rect 2127 3438 2131 3442
rect 2159 3438 2163 3442
rect 2255 3438 2259 3442
rect 2343 3438 2347 3442
rect 2391 3438 2395 3442
rect 2519 3438 2523 3442
rect 2535 3438 2539 3442
rect 2679 3438 2683 3442
rect 2831 3438 2835 3442
rect 2967 3438 2971 3442
rect 2999 3438 3003 3442
rect 3087 3438 3091 3442
rect 3167 3438 3171 3442
rect 3199 3438 3203 3442
rect 3311 3438 3315 3442
rect 3343 3438 3347 3442
rect 3423 3438 3427 3442
rect 3511 3438 3515 3442
rect 3591 3438 3595 3442
rect 111 3398 115 3402
rect 215 3398 219 3402
rect 223 3398 227 3402
rect 359 3398 363 3402
rect 367 3398 371 3402
rect 495 3398 499 3402
rect 511 3398 515 3402
rect 615 3398 619 3402
rect 647 3398 651 3402
rect 727 3398 731 3402
rect 775 3398 779 3402
rect 831 3398 835 3402
rect 895 3398 899 3402
rect 935 3398 939 3402
rect 1015 3398 1019 3402
rect 1031 3398 1035 3402
rect 1127 3398 1131 3402
rect 1223 3398 1227 3402
rect 1239 3398 1243 3402
rect 1319 3398 1323 3402
rect 1351 3398 1355 3402
rect 1831 3398 1835 3402
rect 1871 3362 1875 3366
rect 1999 3362 2003 3366
rect 2015 3362 2019 3366
rect 2119 3362 2123 3366
rect 2151 3362 2155 3366
rect 2247 3362 2251 3366
rect 2295 3362 2299 3366
rect 2383 3362 2387 3366
rect 2439 3362 2443 3366
rect 2527 3362 2531 3366
rect 2583 3362 2587 3366
rect 2671 3362 2675 3366
rect 2727 3362 2731 3366
rect 2823 3362 2827 3366
rect 2871 3362 2875 3366
rect 2991 3362 2995 3366
rect 3023 3362 3027 3366
rect 3159 3362 3163 3366
rect 3183 3362 3187 3366
rect 3335 3362 3339 3366
rect 3351 3362 3355 3366
rect 3503 3362 3507 3366
rect 3591 3362 3595 3366
rect 111 3318 115 3322
rect 207 3318 211 3322
rect 223 3318 227 3322
rect 367 3318 371 3322
rect 375 3318 379 3322
rect 519 3318 523 3322
rect 655 3318 659 3322
rect 671 3318 675 3322
rect 783 3318 787 3322
rect 815 3318 819 3322
rect 903 3318 907 3322
rect 951 3318 955 3322
rect 1023 3318 1027 3322
rect 1087 3318 1091 3322
rect 1135 3318 1139 3322
rect 1215 3318 1219 3322
rect 1247 3318 1251 3322
rect 1343 3318 1347 3322
rect 1359 3318 1363 3322
rect 1471 3318 1475 3322
rect 1831 3318 1835 3322
rect 1871 3286 1875 3290
rect 1927 3286 1931 3290
rect 2023 3286 2027 3290
rect 2063 3286 2067 3290
rect 2159 3286 2163 3290
rect 2191 3286 2195 3290
rect 2303 3286 2307 3290
rect 2319 3286 2323 3290
rect 2447 3286 2451 3290
rect 2591 3286 2595 3290
rect 2735 3286 2739 3290
rect 2743 3286 2747 3290
rect 2879 3286 2883 3290
rect 2919 3286 2923 3290
rect 3031 3286 3035 3290
rect 3111 3286 3115 3290
rect 3191 3286 3195 3290
rect 3311 3286 3315 3290
rect 3359 3286 3363 3290
rect 3511 3286 3515 3290
rect 3591 3286 3595 3290
rect 111 3242 115 3246
rect 135 3242 139 3246
rect 199 3242 203 3246
rect 271 3242 275 3246
rect 359 3242 363 3246
rect 415 3242 419 3246
rect 511 3242 515 3246
rect 575 3242 579 3246
rect 663 3242 667 3246
rect 735 3242 739 3246
rect 807 3242 811 3246
rect 895 3242 899 3246
rect 943 3242 947 3246
rect 1047 3242 1051 3246
rect 1079 3242 1083 3246
rect 1191 3242 1195 3246
rect 1207 3242 1211 3246
rect 1327 3242 1331 3246
rect 1335 3242 1339 3246
rect 1463 3242 1467 3246
rect 1607 3242 1611 3246
rect 1831 3242 1835 3246
rect 1871 3210 1875 3214
rect 1895 3210 1899 3214
rect 1919 3210 1923 3214
rect 2007 3210 2011 3214
rect 2055 3210 2059 3214
rect 2143 3210 2147 3214
rect 2183 3210 2187 3214
rect 2295 3210 2299 3214
rect 2311 3210 2315 3214
rect 2439 3210 2443 3214
rect 2455 3210 2459 3214
rect 2583 3210 2587 3214
rect 2623 3210 2627 3214
rect 2735 3210 2739 3214
rect 2799 3210 2803 3214
rect 2911 3210 2915 3214
rect 2975 3210 2979 3214
rect 3103 3210 3107 3214
rect 3151 3210 3155 3214
rect 3303 3210 3307 3214
rect 3327 3210 3331 3214
rect 3503 3210 3507 3214
rect 3591 3210 3595 3214
rect 111 3158 115 3162
rect 143 3158 147 3162
rect 175 3158 179 3162
rect 279 3158 283 3162
rect 319 3158 323 3162
rect 423 3158 427 3162
rect 463 3158 467 3162
rect 583 3158 587 3162
rect 607 3158 611 3162
rect 743 3158 747 3162
rect 871 3158 875 3162
rect 903 3158 907 3162
rect 991 3158 995 3162
rect 1055 3158 1059 3162
rect 1103 3158 1107 3162
rect 1199 3158 1203 3162
rect 1207 3158 1211 3162
rect 1311 3158 1315 3162
rect 1335 3158 1339 3162
rect 1407 3158 1411 3162
rect 1471 3158 1475 3162
rect 1495 3158 1499 3162
rect 1583 3158 1587 3162
rect 1615 3158 1619 3162
rect 1671 3158 1675 3162
rect 1751 3158 1755 3162
rect 1831 3158 1835 3162
rect 1871 3134 1875 3138
rect 1903 3134 1907 3138
rect 2015 3134 2019 3138
rect 2071 3134 2075 3138
rect 2151 3134 2155 3138
rect 2263 3134 2267 3138
rect 2303 3134 2307 3138
rect 2455 3134 2459 3138
rect 2463 3134 2467 3138
rect 2631 3134 2635 3138
rect 2647 3134 2651 3138
rect 2807 3134 2811 3138
rect 2831 3134 2835 3138
rect 2983 3134 2987 3138
rect 3015 3134 3019 3138
rect 3159 3134 3163 3138
rect 3199 3134 3203 3138
rect 3335 3134 3339 3138
rect 3391 3134 3395 3138
rect 3511 3134 3515 3138
rect 3591 3134 3595 3138
rect 111 3070 115 3074
rect 135 3070 139 3074
rect 167 3070 171 3074
rect 223 3070 227 3074
rect 311 3070 315 3074
rect 327 3070 331 3074
rect 439 3070 443 3074
rect 455 3070 459 3074
rect 551 3070 555 3074
rect 599 3070 603 3074
rect 663 3070 667 3074
rect 735 3070 739 3074
rect 863 3070 867 3074
rect 983 3070 987 3074
rect 1095 3070 1099 3074
rect 1199 3070 1203 3074
rect 1303 3070 1307 3074
rect 1399 3070 1403 3074
rect 1487 3070 1491 3074
rect 1575 3070 1579 3074
rect 1663 3070 1667 3074
rect 1743 3070 1747 3074
rect 1831 3070 1835 3074
rect 1871 3046 1875 3050
rect 1895 3046 1899 3050
rect 2063 3046 2067 3050
rect 2199 3046 2203 3050
rect 2255 3046 2259 3050
rect 2335 3046 2339 3050
rect 2447 3046 2451 3050
rect 2479 3046 2483 3050
rect 2623 3046 2627 3050
rect 2639 3046 2643 3050
rect 2767 3046 2771 3050
rect 2823 3046 2827 3050
rect 2903 3046 2907 3050
rect 3007 3046 3011 3050
rect 3039 3046 3043 3050
rect 3183 3046 3187 3050
rect 3191 3046 3195 3050
rect 3327 3046 3331 3050
rect 3383 3046 3387 3050
rect 3591 3046 3595 3050
rect 111 2982 115 2986
rect 143 2982 147 2986
rect 159 2982 163 2986
rect 231 2982 235 2986
rect 319 2982 323 2986
rect 335 2982 339 2986
rect 447 2982 451 2986
rect 487 2982 491 2986
rect 559 2982 563 2986
rect 647 2982 651 2986
rect 671 2982 675 2986
rect 799 2982 803 2986
rect 943 2982 947 2986
rect 1079 2982 1083 2986
rect 1199 2982 1203 2986
rect 1311 2982 1315 2986
rect 1423 2982 1427 2986
rect 1535 2982 1539 2986
rect 1647 2982 1651 2986
rect 1831 2982 1835 2986
rect 1871 2958 1875 2962
rect 2127 2958 2131 2962
rect 2207 2958 2211 2962
rect 2287 2958 2291 2962
rect 2343 2958 2347 2962
rect 2367 2958 2371 2962
rect 2447 2958 2451 2962
rect 2487 2958 2491 2962
rect 2527 2958 2531 2962
rect 2607 2958 2611 2962
rect 2631 2958 2635 2962
rect 2695 2958 2699 2962
rect 2775 2958 2779 2962
rect 2791 2958 2795 2962
rect 2911 2958 2915 2962
rect 3039 2958 3043 2962
rect 3047 2958 3051 2962
rect 3183 2958 3187 2962
rect 3191 2958 3195 2962
rect 3335 2958 3339 2962
rect 3495 2958 3499 2962
rect 3591 2958 3595 2962
rect 111 2906 115 2910
rect 151 2906 155 2910
rect 311 2906 315 2910
rect 471 2906 475 2910
rect 479 2906 483 2910
rect 631 2906 635 2910
rect 639 2906 643 2910
rect 783 2906 787 2910
rect 791 2906 795 2910
rect 927 2906 931 2910
rect 935 2906 939 2910
rect 1055 2906 1059 2910
rect 1071 2906 1075 2910
rect 1175 2906 1179 2910
rect 1191 2906 1195 2910
rect 1287 2906 1291 2910
rect 1303 2906 1307 2910
rect 1391 2906 1395 2910
rect 1415 2906 1419 2910
rect 1487 2906 1491 2910
rect 1527 2906 1531 2910
rect 1591 2906 1595 2910
rect 1639 2906 1643 2910
rect 1695 2906 1699 2910
rect 1831 2906 1835 2910
rect 1871 2882 1875 2886
rect 2047 2882 2051 2886
rect 2119 2882 2123 2886
rect 2135 2882 2139 2886
rect 2199 2882 2203 2886
rect 2239 2882 2243 2886
rect 2279 2882 2283 2886
rect 2343 2882 2347 2886
rect 2359 2882 2363 2886
rect 2439 2882 2443 2886
rect 2463 2882 2467 2886
rect 2519 2882 2523 2886
rect 2591 2882 2595 2886
rect 2599 2882 2603 2886
rect 2687 2882 2691 2886
rect 2727 2882 2731 2886
rect 2783 2882 2787 2886
rect 2879 2882 2883 2886
rect 2903 2882 2907 2886
rect 3031 2882 3035 2886
rect 3175 2882 3179 2886
rect 3191 2882 3195 2886
rect 3327 2882 3331 2886
rect 3359 2882 3363 2886
rect 3487 2882 3491 2886
rect 3503 2882 3507 2886
rect 3591 2882 3595 2886
rect 111 2826 115 2830
rect 143 2826 147 2830
rect 159 2826 163 2830
rect 247 2826 251 2830
rect 319 2826 323 2830
rect 383 2826 387 2830
rect 479 2826 483 2830
rect 535 2826 539 2830
rect 639 2826 643 2830
rect 687 2826 691 2830
rect 791 2826 795 2830
rect 847 2826 851 2830
rect 935 2826 939 2830
rect 999 2826 1003 2830
rect 1063 2826 1067 2830
rect 1143 2826 1147 2830
rect 1183 2826 1187 2830
rect 1279 2826 1283 2830
rect 1295 2826 1299 2830
rect 1399 2826 1403 2830
rect 1407 2826 1411 2830
rect 1495 2826 1499 2830
rect 1527 2826 1531 2830
rect 1599 2826 1603 2830
rect 1647 2826 1651 2830
rect 1703 2826 1707 2830
rect 1751 2826 1755 2830
rect 1831 2826 1835 2830
rect 1871 2794 1875 2798
rect 1903 2794 1907 2798
rect 2015 2794 2019 2798
rect 2055 2794 2059 2798
rect 2143 2794 2147 2798
rect 2167 2794 2171 2798
rect 2247 2794 2251 2798
rect 2327 2794 2331 2798
rect 2351 2794 2355 2798
rect 2471 2794 2475 2798
rect 2487 2794 2491 2798
rect 2599 2794 2603 2798
rect 2639 2794 2643 2798
rect 2735 2794 2739 2798
rect 2791 2794 2795 2798
rect 2887 2794 2891 2798
rect 2943 2794 2947 2798
rect 3039 2794 3043 2798
rect 3087 2794 3091 2798
rect 3199 2794 3203 2798
rect 3231 2794 3235 2798
rect 3367 2794 3371 2798
rect 3383 2794 3387 2798
rect 3511 2794 3515 2798
rect 3591 2794 3595 2798
rect 111 2746 115 2750
rect 135 2746 139 2750
rect 231 2746 235 2750
rect 239 2746 243 2750
rect 367 2746 371 2750
rect 375 2746 379 2750
rect 511 2746 515 2750
rect 527 2746 531 2750
rect 663 2746 667 2750
rect 679 2746 683 2750
rect 815 2746 819 2750
rect 839 2746 843 2750
rect 975 2746 979 2750
rect 991 2746 995 2750
rect 1135 2746 1139 2750
rect 1271 2746 1275 2750
rect 1287 2746 1291 2750
rect 1399 2746 1403 2750
rect 1447 2746 1451 2750
rect 1519 2746 1523 2750
rect 1607 2746 1611 2750
rect 1639 2746 1643 2750
rect 1743 2746 1747 2750
rect 1831 2746 1835 2750
rect 1871 2718 1875 2722
rect 1895 2718 1899 2722
rect 2007 2718 2011 2722
rect 2103 2718 2107 2722
rect 2159 2718 2163 2722
rect 2319 2718 2323 2722
rect 2327 2718 2331 2722
rect 2479 2718 2483 2722
rect 2535 2718 2539 2722
rect 2631 2718 2635 2722
rect 2735 2718 2739 2722
rect 2783 2718 2787 2722
rect 2911 2718 2915 2722
rect 2935 2718 2939 2722
rect 3071 2718 3075 2722
rect 3079 2718 3083 2722
rect 3223 2718 3227 2722
rect 3375 2718 3379 2722
rect 3503 2718 3507 2722
rect 3591 2718 3595 2722
rect 111 2662 115 2666
rect 143 2662 147 2666
rect 239 2662 243 2666
rect 279 2662 283 2666
rect 375 2662 379 2666
rect 447 2662 451 2666
rect 519 2662 523 2666
rect 623 2662 627 2666
rect 671 2662 675 2666
rect 791 2662 795 2666
rect 823 2662 827 2666
rect 951 2662 955 2666
rect 983 2662 987 2666
rect 1103 2662 1107 2666
rect 1143 2662 1147 2666
rect 1247 2662 1251 2666
rect 1295 2662 1299 2666
rect 1399 2662 1403 2666
rect 1455 2662 1459 2666
rect 1551 2662 1555 2666
rect 1615 2662 1619 2666
rect 1751 2662 1755 2666
rect 1831 2662 1835 2666
rect 1871 2634 1875 2638
rect 1903 2634 1907 2638
rect 2055 2634 2059 2638
rect 2111 2634 2115 2638
rect 2263 2634 2267 2638
rect 2335 2634 2339 2638
rect 2495 2634 2499 2638
rect 2543 2634 2547 2638
rect 2743 2634 2747 2638
rect 2751 2634 2755 2638
rect 2919 2634 2923 2638
rect 3015 2634 3019 2638
rect 3079 2634 3083 2638
rect 3231 2634 3235 2638
rect 3287 2634 3291 2638
rect 3383 2634 3387 2638
rect 3511 2634 3515 2638
rect 3591 2634 3595 2638
rect 111 2582 115 2586
rect 135 2582 139 2586
rect 223 2582 227 2586
rect 271 2582 275 2586
rect 367 2582 371 2586
rect 439 2582 443 2586
rect 527 2582 531 2586
rect 615 2582 619 2586
rect 703 2582 707 2586
rect 783 2582 787 2586
rect 879 2582 883 2586
rect 943 2582 947 2586
rect 1047 2582 1051 2586
rect 1095 2582 1099 2586
rect 1207 2582 1211 2586
rect 1239 2582 1243 2586
rect 1359 2582 1363 2586
rect 1391 2582 1395 2586
rect 1511 2582 1515 2586
rect 1543 2582 1547 2586
rect 1671 2582 1675 2586
rect 1831 2582 1835 2586
rect 1871 2558 1875 2562
rect 1895 2558 1899 2562
rect 2007 2558 2011 2562
rect 2047 2558 2051 2562
rect 2159 2558 2163 2562
rect 2255 2558 2259 2562
rect 2319 2558 2323 2562
rect 2471 2558 2475 2562
rect 2487 2558 2491 2562
rect 2623 2558 2627 2562
rect 2743 2558 2747 2562
rect 2759 2558 2763 2562
rect 2887 2558 2891 2562
rect 3007 2558 3011 2562
rect 3119 2558 3123 2562
rect 3223 2558 3227 2562
rect 3279 2558 3283 2562
rect 3319 2558 3323 2562
rect 3423 2558 3427 2562
rect 3503 2558 3507 2562
rect 3591 2558 3595 2562
rect 111 2502 115 2506
rect 143 2502 147 2506
rect 223 2502 227 2506
rect 231 2502 235 2506
rect 303 2502 307 2506
rect 375 2502 379 2506
rect 391 2502 395 2506
rect 511 2502 515 2506
rect 535 2502 539 2506
rect 647 2502 651 2506
rect 711 2502 715 2506
rect 783 2502 787 2506
rect 887 2502 891 2506
rect 927 2502 931 2506
rect 1055 2502 1059 2506
rect 1063 2502 1067 2506
rect 1191 2502 1195 2506
rect 1215 2502 1219 2506
rect 1311 2502 1315 2506
rect 1367 2502 1371 2506
rect 1431 2502 1435 2506
rect 1519 2502 1523 2506
rect 1551 2502 1555 2506
rect 1671 2502 1675 2506
rect 1679 2502 1683 2506
rect 1831 2502 1835 2506
rect 1871 2474 1875 2478
rect 1903 2474 1907 2478
rect 1999 2474 2003 2478
rect 2015 2474 2019 2478
rect 2127 2474 2131 2478
rect 2167 2474 2171 2478
rect 2263 2474 2267 2478
rect 2327 2474 2331 2478
rect 2407 2474 2411 2478
rect 2479 2474 2483 2478
rect 2551 2474 2555 2478
rect 2631 2474 2635 2478
rect 2703 2474 2707 2478
rect 2767 2474 2771 2478
rect 2863 2474 2867 2478
rect 2895 2474 2899 2478
rect 3015 2474 3019 2478
rect 3023 2474 3027 2478
rect 3127 2474 3131 2478
rect 3191 2474 3195 2478
rect 3231 2474 3235 2478
rect 3327 2474 3331 2478
rect 3359 2474 3363 2478
rect 3431 2474 3435 2478
rect 3511 2474 3515 2478
rect 3591 2474 3595 2478
rect 111 2414 115 2418
rect 135 2414 139 2418
rect 215 2414 219 2418
rect 295 2414 299 2418
rect 383 2414 387 2418
rect 503 2414 507 2418
rect 639 2414 643 2418
rect 775 2414 779 2418
rect 919 2414 923 2418
rect 1055 2414 1059 2418
rect 1063 2414 1067 2418
rect 1143 2414 1147 2418
rect 1183 2414 1187 2418
rect 1223 2414 1227 2418
rect 1303 2414 1307 2418
rect 1383 2414 1387 2418
rect 1423 2414 1427 2418
rect 1463 2414 1467 2418
rect 1543 2414 1547 2418
rect 1663 2414 1667 2418
rect 1831 2414 1835 2418
rect 1871 2394 1875 2398
rect 1991 2394 1995 2398
rect 2119 2394 2123 2398
rect 2143 2394 2147 2398
rect 2239 2394 2243 2398
rect 2255 2394 2259 2398
rect 2343 2394 2347 2398
rect 2399 2394 2403 2398
rect 2455 2394 2459 2398
rect 2543 2394 2547 2398
rect 2575 2394 2579 2398
rect 2695 2394 2699 2398
rect 2703 2394 2707 2398
rect 2847 2394 2851 2398
rect 2855 2394 2859 2398
rect 3007 2394 3011 2398
rect 3015 2394 3019 2398
rect 3175 2394 3179 2398
rect 3183 2394 3187 2398
rect 3351 2394 3355 2398
rect 3503 2394 3507 2398
rect 3591 2394 3595 2398
rect 111 2330 115 2334
rect 359 2330 363 2334
rect 439 2330 443 2334
rect 519 2330 523 2334
rect 599 2330 603 2334
rect 679 2330 683 2334
rect 759 2330 763 2334
rect 839 2330 843 2334
rect 919 2330 923 2334
rect 999 2330 1003 2334
rect 1071 2330 1075 2334
rect 1079 2330 1083 2334
rect 1151 2330 1155 2334
rect 1159 2330 1163 2334
rect 1231 2330 1235 2334
rect 1239 2330 1243 2334
rect 1311 2330 1315 2334
rect 1319 2330 1323 2334
rect 1391 2330 1395 2334
rect 1471 2330 1475 2334
rect 1831 2330 1835 2334
rect 1871 2314 1875 2318
rect 2151 2314 2155 2318
rect 2247 2314 2251 2318
rect 2279 2314 2283 2318
rect 2351 2314 2355 2318
rect 2359 2314 2363 2318
rect 2439 2314 2443 2318
rect 2463 2314 2467 2318
rect 2519 2314 2523 2318
rect 2583 2314 2587 2318
rect 2599 2314 2603 2318
rect 2679 2314 2683 2318
rect 2711 2314 2715 2318
rect 2759 2314 2763 2318
rect 2847 2314 2851 2318
rect 2855 2314 2859 2318
rect 2935 2314 2939 2318
rect 3015 2314 3019 2318
rect 3183 2314 3187 2318
rect 3359 2314 3363 2318
rect 3511 2314 3515 2318
rect 3591 2314 3595 2318
rect 111 2254 115 2258
rect 351 2254 355 2258
rect 375 2254 379 2258
rect 431 2254 435 2258
rect 455 2254 459 2258
rect 511 2254 515 2258
rect 535 2254 539 2258
rect 591 2254 595 2258
rect 615 2254 619 2258
rect 671 2254 675 2258
rect 695 2254 699 2258
rect 751 2254 755 2258
rect 775 2254 779 2258
rect 831 2254 835 2258
rect 855 2254 859 2258
rect 911 2254 915 2258
rect 935 2254 939 2258
rect 991 2254 995 2258
rect 1015 2254 1019 2258
rect 1071 2254 1075 2258
rect 1095 2254 1099 2258
rect 1151 2254 1155 2258
rect 1175 2254 1179 2258
rect 1231 2254 1235 2258
rect 1255 2254 1259 2258
rect 1311 2254 1315 2258
rect 1831 2254 1835 2258
rect 1871 2238 1875 2242
rect 2271 2238 2275 2242
rect 2311 2238 2315 2242
rect 2351 2238 2355 2242
rect 2399 2238 2403 2242
rect 2431 2238 2435 2242
rect 2495 2238 2499 2242
rect 2511 2238 2515 2242
rect 2591 2238 2595 2242
rect 2599 2238 2603 2242
rect 2671 2238 2675 2242
rect 2719 2238 2723 2242
rect 2751 2238 2755 2242
rect 2839 2238 2843 2242
rect 2855 2238 2859 2242
rect 2927 2238 2931 2242
rect 3007 2238 3011 2242
rect 3175 2238 3179 2242
rect 3351 2238 3355 2242
rect 3503 2238 3507 2242
rect 3591 2238 3595 2242
rect 111 2166 115 2170
rect 311 2166 315 2170
rect 383 2166 387 2170
rect 407 2166 411 2170
rect 463 2166 467 2170
rect 503 2166 507 2170
rect 543 2166 547 2170
rect 599 2166 603 2170
rect 623 2166 627 2170
rect 687 2166 691 2170
rect 703 2166 707 2170
rect 775 2166 779 2170
rect 783 2166 787 2170
rect 863 2166 867 2170
rect 943 2166 947 2170
rect 951 2166 955 2170
rect 1023 2166 1027 2170
rect 1039 2166 1043 2170
rect 1103 2166 1107 2170
rect 1127 2166 1131 2170
rect 1183 2166 1187 2170
rect 1223 2166 1227 2170
rect 1263 2166 1267 2170
rect 1831 2166 1835 2170
rect 1871 2158 1875 2162
rect 1903 2158 1907 2162
rect 1983 2158 1987 2162
rect 2111 2158 2115 2162
rect 2247 2158 2251 2162
rect 2319 2158 2323 2162
rect 2391 2158 2395 2162
rect 2407 2158 2411 2162
rect 2503 2158 2507 2162
rect 2543 2158 2547 2162
rect 2607 2158 2611 2162
rect 2695 2158 2699 2162
rect 2727 2158 2731 2162
rect 2847 2158 2851 2162
rect 2863 2158 2867 2162
rect 3007 2158 3011 2162
rect 3015 2158 3019 2162
rect 3175 2158 3179 2162
rect 3183 2158 3187 2162
rect 3351 2158 3355 2162
rect 3359 2158 3363 2162
rect 3511 2158 3515 2162
rect 3591 2158 3595 2162
rect 111 2078 115 2082
rect 207 2078 211 2082
rect 303 2078 307 2082
rect 327 2078 331 2082
rect 399 2078 403 2082
rect 447 2078 451 2082
rect 495 2078 499 2082
rect 575 2078 579 2082
rect 591 2078 595 2082
rect 679 2078 683 2082
rect 703 2078 707 2082
rect 767 2078 771 2082
rect 823 2078 827 2082
rect 855 2078 859 2082
rect 943 2078 947 2082
rect 1031 2078 1035 2082
rect 1063 2078 1067 2082
rect 1119 2078 1123 2082
rect 1175 2078 1179 2082
rect 1215 2078 1219 2082
rect 1279 2078 1283 2082
rect 1375 2078 1379 2082
rect 1471 2078 1475 2082
rect 1567 2078 1571 2082
rect 1663 2078 1667 2082
rect 1743 2078 1747 2082
rect 1831 2078 1835 2082
rect 1871 2074 1875 2078
rect 1895 2074 1899 2078
rect 1967 2074 1971 2078
rect 1975 2074 1979 2078
rect 2103 2074 2107 2078
rect 2215 2074 2219 2078
rect 2239 2074 2243 2078
rect 2383 2074 2387 2078
rect 2447 2074 2451 2078
rect 2535 2074 2539 2078
rect 2655 2074 2659 2078
rect 2687 2074 2691 2078
rect 2839 2074 2843 2078
rect 2999 2074 3003 2078
rect 3143 2074 3147 2078
rect 3167 2074 3171 2078
rect 3271 2074 3275 2078
rect 3343 2074 3347 2078
rect 3399 2074 3403 2078
rect 3503 2074 3507 2078
rect 3591 2074 3595 2078
rect 111 1998 115 2002
rect 191 1998 195 2002
rect 215 1998 219 2002
rect 335 1998 339 2002
rect 351 1998 355 2002
rect 455 1998 459 2002
rect 519 1998 523 2002
rect 583 1998 587 2002
rect 687 1998 691 2002
rect 711 1998 715 2002
rect 831 1998 835 2002
rect 855 1998 859 2002
rect 951 1998 955 2002
rect 1015 1998 1019 2002
rect 1071 1998 1075 2002
rect 1167 1998 1171 2002
rect 1183 1998 1187 2002
rect 1287 1998 1291 2002
rect 1311 1998 1315 2002
rect 1383 1998 1387 2002
rect 1447 1998 1451 2002
rect 1479 1998 1483 2002
rect 1575 1998 1579 2002
rect 1583 1998 1587 2002
rect 1671 1998 1675 2002
rect 1719 1998 1723 2002
rect 1751 1998 1755 2002
rect 1831 1998 1835 2002
rect 1871 1998 1875 2002
rect 1959 1998 1963 2002
rect 1975 1998 1979 2002
rect 2079 1998 2083 2002
rect 2199 1998 2203 2002
rect 2223 1998 2227 2002
rect 2319 1998 2323 2002
rect 2447 1998 2451 2002
rect 2455 1998 2459 2002
rect 2583 1998 2587 2002
rect 2663 1998 2667 2002
rect 2743 1998 2747 2002
rect 2847 1998 2851 2002
rect 2919 1998 2923 2002
rect 3007 1998 3011 2002
rect 3119 1998 3123 2002
rect 3151 1998 3155 2002
rect 3279 1998 3283 2002
rect 3327 1998 3331 2002
rect 3407 1998 3411 2002
rect 3511 1998 3515 2002
rect 3591 1998 3595 2002
rect 111 1918 115 1922
rect 135 1918 139 1922
rect 183 1918 187 1922
rect 239 1918 243 1922
rect 343 1918 347 1922
rect 375 1918 379 1922
rect 511 1918 515 1922
rect 527 1918 531 1922
rect 679 1918 683 1922
rect 687 1918 691 1922
rect 847 1918 851 1922
rect 1007 1918 1011 1922
rect 1159 1918 1163 1922
rect 1303 1918 1307 1922
rect 1439 1918 1443 1922
rect 1455 1918 1459 1922
rect 1575 1918 1579 1922
rect 1607 1918 1611 1922
rect 1711 1918 1715 1922
rect 1831 1918 1835 1922
rect 1871 1914 1875 1918
rect 1951 1914 1955 1918
rect 2063 1914 2067 1918
rect 2071 1914 2075 1918
rect 2151 1914 2155 1918
rect 2191 1914 2195 1918
rect 2239 1914 2243 1918
rect 2311 1914 2315 1918
rect 2319 1914 2323 1918
rect 2399 1914 2403 1918
rect 2439 1914 2443 1918
rect 2487 1914 2491 1918
rect 2575 1914 2579 1918
rect 2663 1914 2667 1918
rect 2735 1914 2739 1918
rect 2759 1914 2763 1918
rect 2871 1914 2875 1918
rect 2911 1914 2915 1918
rect 2991 1914 2995 1918
rect 3111 1914 3115 1918
rect 3119 1914 3123 1918
rect 3247 1914 3251 1918
rect 3319 1914 3323 1918
rect 3383 1914 3387 1918
rect 3503 1914 3507 1918
rect 3591 1914 3595 1918
rect 111 1838 115 1842
rect 143 1838 147 1842
rect 247 1838 251 1842
rect 287 1838 291 1842
rect 383 1838 387 1842
rect 471 1838 475 1842
rect 535 1838 539 1842
rect 663 1838 667 1842
rect 695 1838 699 1842
rect 847 1838 851 1842
rect 855 1838 859 1842
rect 1015 1838 1019 1842
rect 1023 1838 1027 1842
rect 1167 1838 1171 1842
rect 1191 1838 1195 1842
rect 1311 1838 1315 1842
rect 1351 1838 1355 1842
rect 1463 1838 1467 1842
rect 1511 1838 1515 1842
rect 1615 1838 1619 1842
rect 1679 1838 1683 1842
rect 1831 1838 1835 1842
rect 1871 1822 1875 1826
rect 2071 1822 2075 1826
rect 2095 1822 2099 1826
rect 2159 1822 2163 1826
rect 2239 1822 2243 1826
rect 2247 1822 2251 1826
rect 2327 1822 2331 1826
rect 2399 1822 2403 1826
rect 2407 1822 2411 1826
rect 2495 1822 2499 1826
rect 2559 1822 2563 1826
rect 2583 1822 2587 1826
rect 2671 1822 2675 1826
rect 2719 1822 2723 1826
rect 2767 1822 2771 1826
rect 2879 1822 2883 1826
rect 2999 1822 3003 1826
rect 3031 1822 3035 1826
rect 3127 1822 3131 1826
rect 3175 1822 3179 1826
rect 3255 1822 3259 1826
rect 3319 1822 3323 1826
rect 3391 1822 3395 1826
rect 3471 1822 3475 1826
rect 3511 1822 3515 1826
rect 3591 1822 3595 1826
rect 111 1754 115 1758
rect 135 1754 139 1758
rect 215 1754 219 1758
rect 279 1754 283 1758
rect 343 1754 347 1758
rect 463 1754 467 1758
rect 495 1754 499 1758
rect 655 1754 659 1758
rect 663 1754 667 1758
rect 839 1754 843 1758
rect 1007 1754 1011 1758
rect 1015 1754 1019 1758
rect 1167 1754 1171 1758
rect 1183 1754 1187 1758
rect 1319 1754 1323 1758
rect 1343 1754 1347 1758
rect 1463 1754 1467 1758
rect 1503 1754 1507 1758
rect 1607 1754 1611 1758
rect 1671 1754 1675 1758
rect 1743 1754 1747 1758
rect 1831 1754 1835 1758
rect 1871 1742 1875 1746
rect 2087 1742 2091 1746
rect 2103 1742 2107 1746
rect 2231 1742 2235 1746
rect 2239 1742 2243 1746
rect 2383 1742 2387 1746
rect 2391 1742 2395 1746
rect 2527 1742 2531 1746
rect 2551 1742 2555 1746
rect 2663 1742 2667 1746
rect 2711 1742 2715 1746
rect 2799 1742 2803 1746
rect 2871 1742 2875 1746
rect 2927 1742 2931 1746
rect 3023 1742 3027 1746
rect 3047 1742 3051 1746
rect 3159 1742 3163 1746
rect 3167 1742 3171 1746
rect 3271 1742 3275 1746
rect 3311 1742 3315 1746
rect 3391 1742 3395 1746
rect 3463 1742 3467 1746
rect 3503 1742 3507 1746
rect 3591 1742 3595 1746
rect 111 1674 115 1678
rect 143 1674 147 1678
rect 223 1674 227 1678
rect 295 1674 299 1678
rect 351 1674 355 1678
rect 479 1674 483 1678
rect 503 1674 507 1678
rect 671 1674 675 1678
rect 847 1674 851 1678
rect 855 1674 859 1678
rect 1015 1674 1019 1678
rect 1031 1674 1035 1678
rect 1175 1674 1179 1678
rect 1199 1674 1203 1678
rect 1327 1674 1331 1678
rect 1359 1674 1363 1678
rect 1471 1674 1475 1678
rect 1519 1674 1523 1678
rect 1615 1674 1619 1678
rect 1679 1674 1683 1678
rect 1751 1674 1755 1678
rect 1831 1674 1835 1678
rect 1871 1662 1875 1666
rect 1967 1662 1971 1666
rect 2087 1662 2091 1666
rect 2111 1662 2115 1666
rect 2215 1662 2219 1666
rect 2247 1662 2251 1666
rect 2351 1662 2355 1666
rect 2391 1662 2395 1666
rect 2495 1662 2499 1666
rect 2535 1662 2539 1666
rect 2639 1662 2643 1666
rect 2671 1662 2675 1666
rect 2783 1662 2787 1666
rect 2807 1662 2811 1666
rect 2927 1662 2931 1666
rect 2935 1662 2939 1666
rect 3055 1662 3059 1666
rect 3071 1662 3075 1666
rect 3167 1662 3171 1666
rect 3223 1662 3227 1666
rect 3279 1662 3283 1666
rect 3375 1662 3379 1666
rect 3399 1662 3403 1666
rect 3511 1662 3515 1666
rect 3591 1662 3595 1666
rect 111 1598 115 1602
rect 135 1598 139 1602
rect 159 1598 163 1602
rect 287 1598 291 1602
rect 423 1598 427 1602
rect 471 1598 475 1602
rect 567 1598 571 1602
rect 663 1598 667 1602
rect 711 1598 715 1602
rect 847 1598 851 1602
rect 983 1598 987 1602
rect 1023 1598 1027 1602
rect 1119 1598 1123 1602
rect 1191 1598 1195 1602
rect 1247 1598 1251 1602
rect 1351 1598 1355 1602
rect 1375 1598 1379 1602
rect 1511 1598 1515 1602
rect 1671 1598 1675 1602
rect 1831 1598 1835 1602
rect 1871 1578 1875 1582
rect 1895 1578 1899 1582
rect 1959 1578 1963 1582
rect 2047 1578 2051 1582
rect 2079 1578 2083 1582
rect 2207 1578 2211 1582
rect 2343 1578 2347 1582
rect 2367 1578 2371 1582
rect 2487 1578 2491 1582
rect 2527 1578 2531 1582
rect 2631 1578 2635 1582
rect 2687 1578 2691 1582
rect 2775 1578 2779 1582
rect 2839 1578 2843 1582
rect 2919 1578 2923 1582
rect 2983 1578 2987 1582
rect 3063 1578 3067 1582
rect 3119 1578 3123 1582
rect 3215 1578 3219 1582
rect 3255 1578 3259 1582
rect 3367 1578 3371 1582
rect 3391 1578 3395 1582
rect 3503 1578 3507 1582
rect 3591 1578 3595 1582
rect 111 1518 115 1522
rect 167 1518 171 1522
rect 231 1518 235 1522
rect 295 1518 299 1522
rect 375 1518 379 1522
rect 431 1518 435 1522
rect 519 1518 523 1522
rect 575 1518 579 1522
rect 655 1518 659 1522
rect 719 1518 723 1522
rect 783 1518 787 1522
rect 855 1518 859 1522
rect 903 1518 907 1522
rect 991 1518 995 1522
rect 1015 1518 1019 1522
rect 1119 1518 1123 1522
rect 1127 1518 1131 1522
rect 1215 1518 1219 1522
rect 1255 1518 1259 1522
rect 1319 1518 1323 1522
rect 1383 1518 1387 1522
rect 1423 1518 1427 1522
rect 1519 1518 1523 1522
rect 1831 1518 1835 1522
rect 1871 1494 1875 1498
rect 1903 1494 1907 1498
rect 2007 1494 2011 1498
rect 2055 1494 2059 1498
rect 2135 1494 2139 1498
rect 2215 1494 2219 1498
rect 2271 1494 2275 1498
rect 2375 1494 2379 1498
rect 2415 1494 2419 1498
rect 2535 1494 2539 1498
rect 2567 1494 2571 1498
rect 2695 1494 2699 1498
rect 2719 1494 2723 1498
rect 2847 1494 2851 1498
rect 2879 1494 2883 1498
rect 2991 1494 2995 1498
rect 3039 1494 3043 1498
rect 3127 1494 3131 1498
rect 3199 1494 3203 1498
rect 3263 1494 3267 1498
rect 3367 1494 3371 1498
rect 3399 1494 3403 1498
rect 3511 1494 3515 1498
rect 3591 1494 3595 1498
rect 111 1434 115 1438
rect 223 1434 227 1438
rect 255 1434 259 1438
rect 351 1434 355 1438
rect 367 1434 371 1438
rect 447 1434 451 1438
rect 511 1434 515 1438
rect 543 1434 547 1438
rect 631 1434 635 1438
rect 647 1434 651 1438
rect 719 1434 723 1438
rect 775 1434 779 1438
rect 807 1434 811 1438
rect 895 1434 899 1438
rect 919 1434 923 1438
rect 1007 1434 1011 1438
rect 1047 1434 1051 1438
rect 1111 1434 1115 1438
rect 1207 1434 1211 1438
rect 1311 1434 1315 1438
rect 1383 1434 1387 1438
rect 1415 1434 1419 1438
rect 1575 1434 1579 1438
rect 1743 1434 1747 1438
rect 1831 1434 1835 1438
rect 1871 1418 1875 1422
rect 1895 1418 1899 1422
rect 1999 1418 2003 1422
rect 2023 1418 2027 1422
rect 2127 1418 2131 1422
rect 2167 1418 2171 1422
rect 2263 1418 2267 1422
rect 2303 1418 2307 1422
rect 2407 1418 2411 1422
rect 2431 1418 2435 1422
rect 2551 1418 2555 1422
rect 2559 1418 2563 1422
rect 2671 1418 2675 1422
rect 2711 1418 2715 1422
rect 2791 1418 2795 1422
rect 2871 1418 2875 1422
rect 2911 1418 2915 1422
rect 3031 1418 3035 1422
rect 3191 1418 3195 1422
rect 3359 1418 3363 1422
rect 3503 1418 3507 1422
rect 3591 1418 3595 1422
rect 111 1358 115 1362
rect 263 1358 267 1362
rect 359 1358 363 1362
rect 455 1358 459 1362
rect 471 1358 475 1362
rect 551 1358 555 1362
rect 591 1358 595 1362
rect 639 1358 643 1362
rect 727 1358 731 1362
rect 815 1358 819 1362
rect 863 1358 867 1362
rect 927 1358 931 1362
rect 1007 1358 1011 1362
rect 1055 1358 1059 1362
rect 1143 1358 1147 1362
rect 1215 1358 1219 1362
rect 1279 1358 1283 1362
rect 1391 1358 1395 1362
rect 1407 1358 1411 1362
rect 1527 1358 1531 1362
rect 1583 1358 1587 1362
rect 1647 1358 1651 1362
rect 1751 1358 1755 1362
rect 1831 1358 1835 1362
rect 1871 1334 1875 1338
rect 1903 1334 1907 1338
rect 1927 1334 1931 1338
rect 2031 1334 2035 1338
rect 2047 1334 2051 1338
rect 2175 1334 2179 1338
rect 2183 1334 2187 1338
rect 2311 1334 2315 1338
rect 2319 1334 2323 1338
rect 2439 1334 2443 1338
rect 2455 1334 2459 1338
rect 2559 1334 2563 1338
rect 2591 1334 2595 1338
rect 2679 1334 2683 1338
rect 2719 1334 2723 1338
rect 2799 1334 2803 1338
rect 2839 1334 2843 1338
rect 2919 1334 2923 1338
rect 2951 1334 2955 1338
rect 3063 1334 3067 1338
rect 3183 1334 3187 1338
rect 3591 1334 3595 1338
rect 111 1278 115 1282
rect 311 1278 315 1282
rect 351 1278 355 1282
rect 415 1278 419 1282
rect 463 1278 467 1282
rect 535 1278 539 1282
rect 583 1278 587 1282
rect 671 1278 675 1282
rect 719 1278 723 1282
rect 815 1278 819 1282
rect 855 1278 859 1282
rect 959 1278 963 1282
rect 999 1278 1003 1282
rect 1103 1278 1107 1282
rect 1135 1278 1139 1282
rect 1239 1278 1243 1282
rect 1271 1278 1275 1282
rect 1375 1278 1379 1282
rect 1399 1278 1403 1282
rect 1503 1278 1507 1282
rect 1519 1278 1523 1282
rect 1631 1278 1635 1282
rect 1639 1278 1643 1282
rect 1743 1278 1747 1282
rect 1831 1278 1835 1282
rect 1871 1250 1875 1254
rect 1895 1250 1899 1254
rect 1919 1250 1923 1254
rect 2039 1250 2043 1254
rect 2071 1250 2075 1254
rect 2175 1250 2179 1254
rect 2271 1250 2275 1254
rect 2311 1250 2315 1254
rect 2447 1250 2451 1254
rect 2471 1250 2475 1254
rect 2583 1250 2587 1254
rect 2663 1250 2667 1254
rect 2711 1250 2715 1254
rect 2831 1250 2835 1254
rect 2847 1250 2851 1254
rect 2943 1250 2947 1254
rect 3023 1250 3027 1254
rect 3055 1250 3059 1254
rect 3175 1250 3179 1254
rect 3191 1250 3195 1254
rect 3359 1250 3363 1254
rect 3503 1250 3507 1254
rect 3591 1250 3595 1254
rect 111 1202 115 1206
rect 239 1202 243 1206
rect 319 1202 323 1206
rect 415 1202 419 1206
rect 423 1202 427 1206
rect 543 1202 547 1206
rect 591 1202 595 1206
rect 679 1202 683 1206
rect 759 1202 763 1206
rect 823 1202 827 1206
rect 927 1202 931 1206
rect 967 1202 971 1206
rect 1079 1202 1083 1206
rect 1111 1202 1115 1206
rect 1223 1202 1227 1206
rect 1247 1202 1251 1206
rect 1367 1202 1371 1206
rect 1383 1202 1387 1206
rect 1503 1202 1507 1206
rect 1511 1202 1515 1206
rect 1639 1202 1643 1206
rect 1751 1202 1755 1206
rect 1831 1202 1835 1206
rect 1871 1170 1875 1174
rect 1903 1170 1907 1174
rect 1983 1170 1987 1174
rect 2079 1170 2083 1174
rect 2087 1170 2091 1174
rect 2215 1170 2219 1174
rect 2279 1170 2283 1174
rect 2367 1170 2371 1174
rect 2479 1170 2483 1174
rect 2527 1170 2531 1174
rect 2671 1170 2675 1174
rect 2687 1170 2691 1174
rect 2839 1170 2843 1174
rect 2855 1170 2859 1174
rect 2983 1170 2987 1174
rect 3031 1170 3035 1174
rect 3127 1170 3131 1174
rect 3199 1170 3203 1174
rect 3263 1170 3267 1174
rect 3367 1170 3371 1174
rect 3399 1170 3403 1174
rect 3511 1170 3515 1174
rect 3591 1170 3595 1174
rect 111 1122 115 1126
rect 143 1122 147 1126
rect 231 1122 235 1126
rect 279 1122 283 1126
rect 407 1122 411 1126
rect 423 1122 427 1126
rect 567 1122 571 1126
rect 583 1122 587 1126
rect 711 1122 715 1126
rect 751 1122 755 1126
rect 847 1122 851 1126
rect 919 1122 923 1126
rect 975 1122 979 1126
rect 1071 1122 1075 1126
rect 1103 1122 1107 1126
rect 1215 1122 1219 1126
rect 1223 1122 1227 1126
rect 1343 1122 1347 1126
rect 1359 1122 1363 1126
rect 1471 1122 1475 1126
rect 1495 1122 1499 1126
rect 1631 1122 1635 1126
rect 1743 1122 1747 1126
rect 1831 1122 1835 1126
rect 1871 1086 1875 1090
rect 1895 1086 1899 1090
rect 1975 1086 1979 1090
rect 2079 1086 2083 1090
rect 2167 1086 2171 1090
rect 2207 1086 2211 1090
rect 2255 1086 2259 1090
rect 2359 1086 2363 1090
rect 2479 1086 2483 1090
rect 2519 1086 2523 1090
rect 2607 1086 2611 1090
rect 2679 1086 2683 1090
rect 2751 1086 2755 1090
rect 2831 1086 2835 1090
rect 2895 1086 2899 1090
rect 2975 1086 2979 1090
rect 3047 1086 3051 1090
rect 3119 1086 3123 1090
rect 3207 1086 3211 1090
rect 3255 1086 3259 1090
rect 3367 1086 3371 1090
rect 3391 1086 3395 1090
rect 3503 1086 3507 1090
rect 3591 1086 3595 1090
rect 111 1038 115 1042
rect 143 1038 147 1042
rect 151 1038 155 1042
rect 263 1038 267 1042
rect 287 1038 291 1042
rect 407 1038 411 1042
rect 431 1038 435 1042
rect 551 1038 555 1042
rect 575 1038 579 1042
rect 687 1038 691 1042
rect 719 1038 723 1042
rect 807 1038 811 1042
rect 855 1038 859 1042
rect 927 1038 931 1042
rect 983 1038 987 1042
rect 1039 1038 1043 1042
rect 1111 1038 1115 1042
rect 1143 1038 1147 1042
rect 1231 1038 1235 1042
rect 1247 1038 1251 1042
rect 1351 1038 1355 1042
rect 1359 1038 1363 1042
rect 1479 1038 1483 1042
rect 1831 1038 1835 1042
rect 1871 1010 1875 1014
rect 2175 1010 2179 1014
rect 2263 1010 2267 1014
rect 2303 1010 2307 1014
rect 2367 1010 2371 1014
rect 2383 1010 2387 1014
rect 2471 1010 2475 1014
rect 2487 1010 2491 1014
rect 2567 1010 2571 1014
rect 2615 1010 2619 1014
rect 2671 1010 2675 1014
rect 2759 1010 2763 1014
rect 2783 1010 2787 1014
rect 2903 1010 2907 1014
rect 2911 1010 2915 1014
rect 3055 1010 3059 1014
rect 3207 1010 3211 1014
rect 3215 1010 3219 1014
rect 3367 1010 3371 1014
rect 3375 1010 3379 1014
rect 3511 1010 3515 1014
rect 3591 1010 3595 1014
rect 111 954 115 958
rect 135 954 139 958
rect 215 954 219 958
rect 255 954 259 958
rect 327 954 331 958
rect 399 954 403 958
rect 447 954 451 958
rect 543 954 547 958
rect 567 954 571 958
rect 679 954 683 958
rect 687 954 691 958
rect 799 954 803 958
rect 911 954 915 958
rect 919 954 923 958
rect 1015 954 1019 958
rect 1031 954 1035 958
rect 1119 954 1123 958
rect 1135 954 1139 958
rect 1223 954 1227 958
rect 1239 954 1243 958
rect 1327 954 1331 958
rect 1351 954 1355 958
rect 1831 954 1835 958
rect 1871 926 1875 930
rect 2279 926 2283 930
rect 2295 926 2299 930
rect 2359 926 2363 930
rect 2375 926 2379 930
rect 2439 926 2443 930
rect 2463 926 2467 930
rect 2519 926 2523 930
rect 2559 926 2563 930
rect 2607 926 2611 930
rect 2663 926 2667 930
rect 2703 926 2707 930
rect 2775 926 2779 930
rect 2807 926 2811 930
rect 2903 926 2907 930
rect 2911 926 2915 930
rect 3015 926 3019 930
rect 3047 926 3051 930
rect 3111 926 3115 930
rect 3199 926 3203 930
rect 3215 926 3219 930
rect 3319 926 3323 930
rect 3359 926 3363 930
rect 3423 926 3427 930
rect 3503 926 3507 930
rect 3591 926 3595 930
rect 111 870 115 874
rect 143 870 147 874
rect 223 870 227 874
rect 255 870 259 874
rect 335 870 339 874
rect 399 870 403 874
rect 455 870 459 874
rect 559 870 563 874
rect 575 870 579 874
rect 695 870 699 874
rect 719 870 723 874
rect 807 870 811 874
rect 871 870 875 874
rect 919 870 923 874
rect 1015 870 1019 874
rect 1023 870 1027 874
rect 1127 870 1131 874
rect 1151 870 1155 874
rect 1231 870 1235 874
rect 1279 870 1283 874
rect 1335 870 1339 874
rect 1399 870 1403 874
rect 1519 870 1523 874
rect 1647 870 1651 874
rect 1831 870 1835 874
rect 1871 838 1875 842
rect 2167 838 2171 842
rect 2247 838 2251 842
rect 2287 838 2291 842
rect 2327 838 2331 842
rect 2367 838 2371 842
rect 2423 838 2427 842
rect 2447 838 2451 842
rect 2527 838 2531 842
rect 2535 838 2539 842
rect 2615 838 2619 842
rect 2655 838 2659 842
rect 2711 838 2715 842
rect 2783 838 2787 842
rect 2815 838 2819 842
rect 2911 838 2915 842
rect 2919 838 2923 842
rect 3023 838 3027 842
rect 3039 838 3043 842
rect 3119 838 3123 842
rect 3159 838 3163 842
rect 3223 838 3227 842
rect 3279 838 3283 842
rect 3327 838 3331 842
rect 3407 838 3411 842
rect 3431 838 3435 842
rect 3511 838 3515 842
rect 3591 838 3595 842
rect 111 782 115 786
rect 135 782 139 786
rect 247 782 251 786
rect 263 782 267 786
rect 391 782 395 786
rect 431 782 435 786
rect 551 782 555 786
rect 607 782 611 786
rect 711 782 715 786
rect 783 782 787 786
rect 863 782 867 786
rect 951 782 955 786
rect 1007 782 1011 786
rect 1103 782 1107 786
rect 1143 782 1147 786
rect 1247 782 1251 786
rect 1271 782 1275 786
rect 1383 782 1387 786
rect 1391 782 1395 786
rect 1511 782 1515 786
rect 1639 782 1643 786
rect 1743 782 1747 786
rect 1831 782 1835 786
rect 1871 754 1875 758
rect 1895 754 1899 758
rect 1975 754 1979 758
rect 2071 754 2075 758
rect 2159 754 2163 758
rect 2183 754 2187 758
rect 2239 754 2243 758
rect 2311 754 2315 758
rect 2319 754 2323 758
rect 2415 754 2419 758
rect 2447 754 2451 758
rect 2527 754 2531 758
rect 2591 754 2595 758
rect 2647 754 2651 758
rect 2743 754 2747 758
rect 2775 754 2779 758
rect 2895 754 2899 758
rect 2903 754 2907 758
rect 3031 754 3035 758
rect 3047 754 3051 758
rect 3151 754 3155 758
rect 3199 754 3203 758
rect 3271 754 3275 758
rect 3359 754 3363 758
rect 3399 754 3403 758
rect 3503 754 3507 758
rect 3591 754 3595 758
rect 111 694 115 698
rect 143 694 147 698
rect 271 694 275 698
rect 295 694 299 698
rect 407 694 411 698
rect 439 694 443 698
rect 527 694 531 698
rect 615 694 619 698
rect 655 694 659 698
rect 783 694 787 698
rect 791 694 795 698
rect 903 694 907 698
rect 959 694 963 698
rect 1023 694 1027 698
rect 1111 694 1115 698
rect 1135 694 1139 698
rect 1247 694 1251 698
rect 1255 694 1259 698
rect 1351 694 1355 698
rect 1391 694 1395 698
rect 1455 694 1459 698
rect 1519 694 1523 698
rect 1559 694 1563 698
rect 1647 694 1651 698
rect 1663 694 1667 698
rect 1751 694 1755 698
rect 1831 694 1835 698
rect 1871 674 1875 678
rect 1903 674 1907 678
rect 1983 674 1987 678
rect 2079 674 2083 678
rect 2095 674 2099 678
rect 2191 674 2195 678
rect 2295 674 2299 678
rect 2319 674 2323 678
rect 2455 674 2459 678
rect 2479 674 2483 678
rect 2599 674 2603 678
rect 2655 674 2659 678
rect 2751 674 2755 678
rect 2831 674 2835 678
rect 2903 674 2907 678
rect 3007 674 3011 678
rect 3055 674 3059 678
rect 3183 674 3187 678
rect 3207 674 3211 678
rect 3359 674 3363 678
rect 3367 674 3371 678
rect 3511 674 3515 678
rect 3591 674 3595 678
rect 111 614 115 618
rect 287 614 291 618
rect 311 614 315 618
rect 391 614 395 618
rect 399 614 403 618
rect 471 614 475 618
rect 519 614 523 618
rect 559 614 563 618
rect 647 614 651 618
rect 735 614 739 618
rect 775 614 779 618
rect 823 614 827 618
rect 895 614 899 618
rect 911 614 915 618
rect 999 614 1003 618
rect 1015 614 1019 618
rect 1087 614 1091 618
rect 1127 614 1131 618
rect 1175 614 1179 618
rect 1239 614 1243 618
rect 1263 614 1267 618
rect 1343 614 1347 618
rect 1447 614 1451 618
rect 1551 614 1555 618
rect 1655 614 1659 618
rect 1743 614 1747 618
rect 1831 614 1835 618
rect 1871 594 1875 598
rect 1895 594 1899 598
rect 1975 594 1979 598
rect 2087 594 2091 598
rect 2215 594 2219 598
rect 2287 594 2291 598
rect 2351 594 2355 598
rect 2471 594 2475 598
rect 2495 594 2499 598
rect 2647 594 2651 598
rect 2807 594 2811 598
rect 2823 594 2827 598
rect 2975 594 2979 598
rect 2999 594 3003 598
rect 3151 594 3155 598
rect 3175 594 3179 598
rect 3335 594 3339 598
rect 3351 594 3355 598
rect 3503 594 3507 598
rect 3591 594 3595 598
rect 111 526 115 530
rect 239 526 243 530
rect 319 526 323 530
rect 343 526 347 530
rect 399 526 403 530
rect 439 526 443 530
rect 479 526 483 530
rect 535 526 539 530
rect 567 526 571 530
rect 631 526 635 530
rect 655 526 659 530
rect 719 526 723 530
rect 743 526 747 530
rect 807 526 811 530
rect 831 526 835 530
rect 895 526 899 530
rect 919 526 923 530
rect 983 526 987 530
rect 1007 526 1011 530
rect 1071 526 1075 530
rect 1095 526 1099 530
rect 1159 526 1163 530
rect 1183 526 1187 530
rect 1247 526 1251 530
rect 1271 526 1275 530
rect 1831 526 1835 530
rect 1871 518 1875 522
rect 1903 518 1907 522
rect 1983 518 1987 522
rect 2095 518 2099 522
rect 2151 518 2155 522
rect 2223 518 2227 522
rect 2231 518 2235 522
rect 2327 518 2331 522
rect 2359 518 2363 522
rect 2431 518 2435 522
rect 2503 518 2507 522
rect 2551 518 2555 522
rect 2655 518 2659 522
rect 2687 518 2691 522
rect 2815 518 2819 522
rect 2839 518 2843 522
rect 2983 518 2987 522
rect 2999 518 3003 522
rect 3159 518 3163 522
rect 3175 518 3179 522
rect 3343 518 3347 522
rect 3351 518 3355 522
rect 3511 518 3515 522
rect 3591 518 3595 522
rect 111 442 115 446
rect 135 442 139 446
rect 231 442 235 446
rect 247 442 251 446
rect 335 442 339 446
rect 375 442 379 446
rect 431 442 435 446
rect 495 442 499 446
rect 527 442 531 446
rect 607 442 611 446
rect 623 442 627 446
rect 711 442 715 446
rect 719 442 723 446
rect 799 442 803 446
rect 823 442 827 446
rect 887 442 891 446
rect 919 442 923 446
rect 975 442 979 446
rect 1007 442 1011 446
rect 1063 442 1067 446
rect 1103 442 1107 446
rect 1151 442 1155 446
rect 1199 442 1203 446
rect 1239 442 1243 446
rect 1295 442 1299 446
rect 1831 442 1835 446
rect 1871 438 1875 442
rect 2143 438 2147 442
rect 2223 438 2227 442
rect 2319 438 2323 442
rect 2335 438 2339 442
rect 2415 438 2419 442
rect 2423 438 2427 442
rect 2495 438 2499 442
rect 2543 438 2547 442
rect 2583 438 2587 442
rect 2679 438 2683 442
rect 2687 438 2691 442
rect 2799 438 2803 442
rect 2831 438 2835 442
rect 2927 438 2931 442
rect 2991 438 2995 442
rect 3071 438 3075 442
rect 3167 438 3171 442
rect 3215 438 3219 442
rect 3343 438 3347 442
rect 3367 438 3371 442
rect 3503 438 3507 442
rect 3591 438 3595 442
rect 111 354 115 358
rect 143 354 147 358
rect 247 354 251 358
rect 255 354 259 358
rect 375 354 379 358
rect 383 354 387 358
rect 503 354 507 358
rect 511 354 515 358
rect 615 354 619 358
rect 647 354 651 358
rect 727 354 731 358
rect 775 354 779 358
rect 831 354 835 358
rect 895 354 899 358
rect 927 354 931 358
rect 1007 354 1011 358
rect 1015 354 1019 358
rect 1111 354 1115 358
rect 1119 354 1123 358
rect 1207 354 1211 358
rect 1223 354 1227 358
rect 1303 354 1307 358
rect 1327 354 1331 358
rect 1439 354 1443 358
rect 1831 354 1835 358
rect 1871 354 1875 358
rect 2079 354 2083 358
rect 2167 354 2171 358
rect 2263 354 2267 358
rect 2343 354 2347 358
rect 2375 354 2379 358
rect 2423 354 2427 358
rect 2503 354 2507 358
rect 2591 354 2595 358
rect 2639 354 2643 358
rect 2695 354 2699 358
rect 2775 354 2779 358
rect 2807 354 2811 358
rect 2911 354 2915 358
rect 2935 354 2939 358
rect 3039 354 3043 358
rect 3079 354 3083 358
rect 3167 354 3171 358
rect 3223 354 3227 358
rect 3287 354 3291 358
rect 3375 354 3379 358
rect 3407 354 3411 358
rect 3511 354 3515 358
rect 3591 354 3595 358
rect 111 270 115 274
rect 135 270 139 274
rect 223 270 227 274
rect 239 270 243 274
rect 335 270 339 274
rect 367 270 371 274
rect 463 270 467 274
rect 503 270 507 274
rect 599 270 603 274
rect 639 270 643 274
rect 735 270 739 274
rect 767 270 771 274
rect 871 270 875 274
rect 887 270 891 274
rect 999 270 1003 274
rect 1007 270 1011 274
rect 1111 270 1115 274
rect 1135 270 1139 274
rect 1215 270 1219 274
rect 1255 270 1259 274
rect 1319 270 1323 274
rect 1367 270 1371 274
rect 1431 270 1435 274
rect 1479 270 1483 274
rect 1599 270 1603 274
rect 1831 270 1835 274
rect 1871 270 1875 274
rect 1895 270 1899 274
rect 1983 270 1987 274
rect 2071 270 2075 274
rect 2095 270 2099 274
rect 2159 270 2163 274
rect 2223 270 2227 274
rect 2255 270 2259 274
rect 2359 270 2363 274
rect 2367 270 2371 274
rect 2495 270 2499 274
rect 2503 270 2507 274
rect 2631 270 2635 274
rect 2647 270 2651 274
rect 2767 270 2771 274
rect 2791 270 2795 274
rect 2903 270 2907 274
rect 2935 270 2939 274
rect 3031 270 3035 274
rect 3079 270 3083 274
rect 3159 270 3163 274
rect 3223 270 3227 274
rect 3279 270 3283 274
rect 3375 270 3379 274
rect 3399 270 3403 274
rect 3503 270 3507 274
rect 3591 270 3595 274
rect 1871 182 1875 186
rect 1903 182 1907 186
rect 1983 182 1987 186
rect 1991 182 1995 186
rect 2087 182 2091 186
rect 2103 182 2107 186
rect 2207 182 2211 186
rect 2231 182 2235 186
rect 2335 182 2339 186
rect 2367 182 2371 186
rect 2463 182 2467 186
rect 2511 182 2515 186
rect 2583 182 2587 186
rect 2655 182 2659 186
rect 2703 182 2707 186
rect 2799 182 2803 186
rect 2815 182 2819 186
rect 2919 182 2923 186
rect 2943 182 2947 186
rect 3015 182 3019 186
rect 3087 182 3091 186
rect 3111 182 3115 186
rect 3207 182 3211 186
rect 3231 182 3235 186
rect 3303 182 3307 186
rect 3383 182 3387 186
rect 3399 182 3403 186
rect 3511 182 3515 186
rect 3591 182 3595 186
rect 111 162 115 166
rect 159 162 163 166
rect 231 162 235 166
rect 239 162 243 166
rect 319 162 323 166
rect 343 162 347 166
rect 399 162 403 166
rect 471 162 475 166
rect 479 162 483 166
rect 559 162 563 166
rect 607 162 611 166
rect 647 162 651 166
rect 735 162 739 166
rect 743 162 747 166
rect 823 162 827 166
rect 879 162 883 166
rect 911 162 915 166
rect 999 162 1003 166
rect 1015 162 1019 166
rect 1087 162 1091 166
rect 1143 162 1147 166
rect 1167 162 1171 166
rect 1247 162 1251 166
rect 1263 162 1267 166
rect 1335 162 1339 166
rect 1375 162 1379 166
rect 1423 162 1427 166
rect 1487 162 1491 166
rect 1511 162 1515 166
rect 1591 162 1595 166
rect 1607 162 1611 166
rect 1671 162 1675 166
rect 1751 162 1755 166
rect 1831 162 1835 166
rect 1871 106 1875 110
rect 1895 106 1899 110
rect 1975 106 1979 110
rect 2079 106 2083 110
rect 2199 106 2203 110
rect 2327 106 2331 110
rect 2455 106 2459 110
rect 2575 106 2579 110
rect 2695 106 2699 110
rect 2807 106 2811 110
rect 2911 106 2915 110
rect 3007 106 3011 110
rect 3103 106 3107 110
rect 3199 106 3203 110
rect 3295 106 3299 110
rect 3391 106 3395 110
rect 3591 106 3595 110
rect 111 86 115 90
rect 151 86 155 90
rect 231 86 235 90
rect 311 86 315 90
rect 391 86 395 90
rect 471 86 475 90
rect 551 86 555 90
rect 639 86 643 90
rect 727 86 731 90
rect 815 86 819 90
rect 903 86 907 90
rect 991 86 995 90
rect 1079 86 1083 90
rect 1159 86 1163 90
rect 1239 86 1243 90
rect 1327 86 1331 90
rect 1415 86 1419 90
rect 1503 86 1507 90
rect 1583 86 1587 90
rect 1663 86 1667 90
rect 1743 86 1747 90
rect 1831 86 1835 90
<< m4 >>
rect 1842 3665 1843 3671
rect 1849 3670 3619 3671
rect 1849 3666 1871 3670
rect 1875 3666 2151 3670
rect 2155 3666 2439 3670
rect 2443 3666 2727 3670
rect 2731 3666 3015 3670
rect 3019 3666 3591 3670
rect 3595 3666 3619 3670
rect 1849 3665 3619 3666
rect 3625 3665 3626 3671
rect 96 3637 97 3643
rect 103 3642 1855 3643
rect 103 3638 111 3642
rect 115 3638 143 3642
rect 147 3638 239 3642
rect 243 3638 367 3642
rect 371 3638 503 3642
rect 507 3638 639 3642
rect 643 3638 775 3642
rect 779 3638 911 3642
rect 915 3638 1055 3642
rect 1059 3638 1199 3642
rect 1203 3638 1831 3642
rect 1835 3638 1855 3642
rect 103 3637 1855 3638
rect 1861 3637 1862 3643
rect 1854 3589 1855 3595
rect 1861 3594 3631 3595
rect 1861 3590 1871 3594
rect 1875 3590 1903 3594
rect 1907 3590 1983 3594
rect 1987 3590 2071 3594
rect 2075 3590 2159 3594
rect 2163 3590 2175 3594
rect 2179 3590 2295 3594
rect 2299 3590 2423 3594
rect 2427 3590 2447 3594
rect 2451 3590 2559 3594
rect 2563 3590 2695 3594
rect 2699 3590 2735 3594
rect 2739 3590 2831 3594
rect 2835 3590 2975 3594
rect 2979 3590 3023 3594
rect 3027 3590 3119 3594
rect 3123 3590 3263 3594
rect 3267 3590 3591 3594
rect 3595 3590 3631 3594
rect 1861 3589 3631 3590
rect 3637 3589 3638 3595
rect 84 3561 85 3567
rect 91 3566 1843 3567
rect 91 3562 111 3566
rect 115 3562 135 3566
rect 139 3562 183 3566
rect 187 3562 231 3566
rect 235 3562 303 3566
rect 307 3562 359 3566
rect 363 3562 415 3566
rect 419 3562 495 3566
rect 499 3562 527 3566
rect 531 3562 631 3566
rect 635 3562 735 3566
rect 739 3562 767 3566
rect 771 3562 831 3566
rect 835 3562 903 3566
rect 907 3562 919 3566
rect 923 3562 1007 3566
rect 1011 3562 1047 3566
rect 1051 3562 1095 3566
rect 1099 3562 1183 3566
rect 1187 3562 1191 3566
rect 1195 3562 1271 3566
rect 1275 3562 1359 3566
rect 1363 3562 1447 3566
rect 1451 3562 1831 3566
rect 1835 3562 1843 3566
rect 91 3561 1843 3562
rect 1849 3561 1850 3567
rect 1842 3513 1843 3519
rect 1849 3518 3619 3519
rect 1849 3514 1871 3518
rect 1875 3514 1895 3518
rect 1899 3514 1967 3518
rect 1971 3514 1975 3518
rect 1979 3514 2063 3518
rect 2067 3514 2151 3518
rect 2155 3514 2167 3518
rect 2171 3514 2287 3518
rect 2291 3514 2335 3518
rect 2339 3514 2415 3518
rect 2419 3514 2511 3518
rect 2515 3514 2551 3518
rect 2555 3514 2671 3518
rect 2675 3514 2687 3518
rect 2691 3514 2823 3518
rect 2827 3514 2959 3518
rect 2963 3514 2967 3518
rect 2971 3514 3079 3518
rect 3083 3514 3111 3518
rect 3115 3514 3191 3518
rect 3195 3514 3255 3518
rect 3259 3514 3303 3518
rect 3307 3514 3415 3518
rect 3419 3514 3503 3518
rect 3507 3514 3591 3518
rect 3595 3514 3619 3518
rect 1849 3513 3619 3514
rect 3625 3513 3626 3519
rect 96 3477 97 3483
rect 103 3482 1855 3483
rect 103 3478 111 3482
rect 115 3478 191 3482
rect 195 3478 231 3482
rect 235 3478 311 3482
rect 315 3478 367 3482
rect 371 3478 423 3482
rect 427 3478 503 3482
rect 507 3478 535 3482
rect 539 3478 623 3482
rect 627 3478 639 3482
rect 643 3478 735 3482
rect 739 3478 743 3482
rect 747 3478 839 3482
rect 843 3478 927 3482
rect 931 3478 943 3482
rect 947 3478 1015 3482
rect 1019 3478 1039 3482
rect 1043 3478 1103 3482
rect 1107 3478 1135 3482
rect 1139 3478 1191 3482
rect 1195 3478 1231 3482
rect 1235 3478 1279 3482
rect 1283 3478 1327 3482
rect 1331 3478 1367 3482
rect 1371 3478 1455 3482
rect 1459 3478 1831 3482
rect 1835 3478 1855 3482
rect 103 3477 1855 3478
rect 1861 3477 1862 3483
rect 1854 3437 1855 3443
rect 1861 3442 3631 3443
rect 1861 3438 1871 3442
rect 1875 3438 1975 3442
rect 1979 3438 2007 3442
rect 2011 3438 2127 3442
rect 2131 3438 2159 3442
rect 2163 3438 2255 3442
rect 2259 3438 2343 3442
rect 2347 3438 2391 3442
rect 2395 3438 2519 3442
rect 2523 3438 2535 3442
rect 2539 3438 2679 3442
rect 2683 3438 2831 3442
rect 2835 3438 2967 3442
rect 2971 3438 2999 3442
rect 3003 3438 3087 3442
rect 3091 3438 3167 3442
rect 3171 3438 3199 3442
rect 3203 3438 3311 3442
rect 3315 3438 3343 3442
rect 3347 3438 3423 3442
rect 3427 3438 3511 3442
rect 3515 3438 3591 3442
rect 3595 3438 3631 3442
rect 1861 3437 3631 3438
rect 3637 3437 3638 3443
rect 84 3397 85 3403
rect 91 3402 1843 3403
rect 91 3398 111 3402
rect 115 3398 215 3402
rect 219 3398 223 3402
rect 227 3398 359 3402
rect 363 3398 367 3402
rect 371 3398 495 3402
rect 499 3398 511 3402
rect 515 3398 615 3402
rect 619 3398 647 3402
rect 651 3398 727 3402
rect 731 3398 775 3402
rect 779 3398 831 3402
rect 835 3398 895 3402
rect 899 3398 935 3402
rect 939 3398 1015 3402
rect 1019 3398 1031 3402
rect 1035 3398 1127 3402
rect 1131 3398 1223 3402
rect 1227 3398 1239 3402
rect 1243 3398 1319 3402
rect 1323 3398 1351 3402
rect 1355 3398 1831 3402
rect 1835 3398 1843 3402
rect 91 3397 1843 3398
rect 1849 3397 1850 3403
rect 1842 3361 1843 3367
rect 1849 3366 3619 3367
rect 1849 3362 1871 3366
rect 1875 3362 1999 3366
rect 2003 3362 2015 3366
rect 2019 3362 2119 3366
rect 2123 3362 2151 3366
rect 2155 3362 2247 3366
rect 2251 3362 2295 3366
rect 2299 3362 2383 3366
rect 2387 3362 2439 3366
rect 2443 3362 2527 3366
rect 2531 3362 2583 3366
rect 2587 3362 2671 3366
rect 2675 3362 2727 3366
rect 2731 3362 2823 3366
rect 2827 3362 2871 3366
rect 2875 3362 2991 3366
rect 2995 3362 3023 3366
rect 3027 3362 3159 3366
rect 3163 3362 3183 3366
rect 3187 3362 3335 3366
rect 3339 3362 3351 3366
rect 3355 3362 3503 3366
rect 3507 3362 3591 3366
rect 3595 3362 3619 3366
rect 1849 3361 3619 3362
rect 3625 3361 3626 3367
rect 96 3317 97 3323
rect 103 3322 1855 3323
rect 103 3318 111 3322
rect 115 3318 207 3322
rect 211 3318 223 3322
rect 227 3318 367 3322
rect 371 3318 375 3322
rect 379 3318 519 3322
rect 523 3318 655 3322
rect 659 3318 671 3322
rect 675 3318 783 3322
rect 787 3318 815 3322
rect 819 3318 903 3322
rect 907 3318 951 3322
rect 955 3318 1023 3322
rect 1027 3318 1087 3322
rect 1091 3318 1135 3322
rect 1139 3318 1215 3322
rect 1219 3318 1247 3322
rect 1251 3318 1343 3322
rect 1347 3318 1359 3322
rect 1363 3318 1471 3322
rect 1475 3318 1831 3322
rect 1835 3318 1855 3322
rect 103 3317 1855 3318
rect 1861 3317 1862 3323
rect 1854 3285 1855 3291
rect 1861 3290 3631 3291
rect 1861 3286 1871 3290
rect 1875 3286 1927 3290
rect 1931 3286 2023 3290
rect 2027 3286 2063 3290
rect 2067 3286 2159 3290
rect 2163 3286 2191 3290
rect 2195 3286 2303 3290
rect 2307 3286 2319 3290
rect 2323 3286 2447 3290
rect 2451 3286 2591 3290
rect 2595 3286 2735 3290
rect 2739 3286 2743 3290
rect 2747 3286 2879 3290
rect 2883 3286 2919 3290
rect 2923 3286 3031 3290
rect 3035 3286 3111 3290
rect 3115 3286 3191 3290
rect 3195 3286 3311 3290
rect 3315 3286 3359 3290
rect 3363 3286 3511 3290
rect 3515 3286 3591 3290
rect 3595 3286 3631 3290
rect 1861 3285 3631 3286
rect 3637 3285 3638 3291
rect 84 3241 85 3247
rect 91 3246 1843 3247
rect 91 3242 111 3246
rect 115 3242 135 3246
rect 139 3242 199 3246
rect 203 3242 271 3246
rect 275 3242 359 3246
rect 363 3242 415 3246
rect 419 3242 511 3246
rect 515 3242 575 3246
rect 579 3242 663 3246
rect 667 3242 735 3246
rect 739 3242 807 3246
rect 811 3242 895 3246
rect 899 3242 943 3246
rect 947 3242 1047 3246
rect 1051 3242 1079 3246
rect 1083 3242 1191 3246
rect 1195 3242 1207 3246
rect 1211 3242 1327 3246
rect 1331 3242 1335 3246
rect 1339 3242 1463 3246
rect 1467 3242 1607 3246
rect 1611 3242 1831 3246
rect 1835 3242 1843 3246
rect 91 3241 1843 3242
rect 1849 3241 1850 3247
rect 1842 3209 1843 3215
rect 1849 3214 3619 3215
rect 1849 3210 1871 3214
rect 1875 3210 1895 3214
rect 1899 3210 1919 3214
rect 1923 3210 2007 3214
rect 2011 3210 2055 3214
rect 2059 3210 2143 3214
rect 2147 3210 2183 3214
rect 2187 3210 2295 3214
rect 2299 3210 2311 3214
rect 2315 3210 2439 3214
rect 2443 3210 2455 3214
rect 2459 3210 2583 3214
rect 2587 3210 2623 3214
rect 2627 3210 2735 3214
rect 2739 3210 2799 3214
rect 2803 3210 2911 3214
rect 2915 3210 2975 3214
rect 2979 3210 3103 3214
rect 3107 3210 3151 3214
rect 3155 3210 3303 3214
rect 3307 3210 3327 3214
rect 3331 3210 3503 3214
rect 3507 3210 3591 3214
rect 3595 3210 3619 3214
rect 1849 3209 3619 3210
rect 3625 3209 3626 3215
rect 96 3157 97 3163
rect 103 3162 1855 3163
rect 103 3158 111 3162
rect 115 3158 143 3162
rect 147 3158 175 3162
rect 179 3158 279 3162
rect 283 3158 319 3162
rect 323 3158 423 3162
rect 427 3158 463 3162
rect 467 3158 583 3162
rect 587 3158 607 3162
rect 611 3158 743 3162
rect 747 3158 871 3162
rect 875 3158 903 3162
rect 907 3158 991 3162
rect 995 3158 1055 3162
rect 1059 3158 1103 3162
rect 1107 3158 1199 3162
rect 1203 3158 1207 3162
rect 1211 3158 1311 3162
rect 1315 3158 1335 3162
rect 1339 3158 1407 3162
rect 1411 3158 1471 3162
rect 1475 3158 1495 3162
rect 1499 3158 1583 3162
rect 1587 3158 1615 3162
rect 1619 3158 1671 3162
rect 1675 3158 1751 3162
rect 1755 3158 1831 3162
rect 1835 3158 1855 3162
rect 103 3157 1855 3158
rect 1861 3157 1862 3163
rect 1854 3133 1855 3139
rect 1861 3138 3631 3139
rect 1861 3134 1871 3138
rect 1875 3134 1903 3138
rect 1907 3134 2015 3138
rect 2019 3134 2071 3138
rect 2075 3134 2151 3138
rect 2155 3134 2263 3138
rect 2267 3134 2303 3138
rect 2307 3134 2455 3138
rect 2459 3134 2463 3138
rect 2467 3134 2631 3138
rect 2635 3134 2647 3138
rect 2651 3134 2807 3138
rect 2811 3134 2831 3138
rect 2835 3134 2983 3138
rect 2987 3134 3015 3138
rect 3019 3134 3159 3138
rect 3163 3134 3199 3138
rect 3203 3134 3335 3138
rect 3339 3134 3391 3138
rect 3395 3134 3511 3138
rect 3515 3134 3591 3138
rect 3595 3134 3631 3138
rect 1861 3133 3631 3134
rect 3637 3133 3638 3139
rect 84 3069 85 3075
rect 91 3074 1843 3075
rect 91 3070 111 3074
rect 115 3070 135 3074
rect 139 3070 167 3074
rect 171 3070 223 3074
rect 227 3070 311 3074
rect 315 3070 327 3074
rect 331 3070 439 3074
rect 443 3070 455 3074
rect 459 3070 551 3074
rect 555 3070 599 3074
rect 603 3070 663 3074
rect 667 3070 735 3074
rect 739 3070 863 3074
rect 867 3070 983 3074
rect 987 3070 1095 3074
rect 1099 3070 1199 3074
rect 1203 3070 1303 3074
rect 1307 3070 1399 3074
rect 1403 3070 1487 3074
rect 1491 3070 1575 3074
rect 1579 3070 1663 3074
rect 1667 3070 1743 3074
rect 1747 3070 1831 3074
rect 1835 3070 1843 3074
rect 91 3069 1843 3070
rect 1849 3069 1850 3075
rect 1842 3045 1843 3051
rect 1849 3050 3619 3051
rect 1849 3046 1871 3050
rect 1875 3046 1895 3050
rect 1899 3046 2063 3050
rect 2067 3046 2199 3050
rect 2203 3046 2255 3050
rect 2259 3046 2335 3050
rect 2339 3046 2447 3050
rect 2451 3046 2479 3050
rect 2483 3046 2623 3050
rect 2627 3046 2639 3050
rect 2643 3046 2767 3050
rect 2771 3046 2823 3050
rect 2827 3046 2903 3050
rect 2907 3046 3007 3050
rect 3011 3046 3039 3050
rect 3043 3046 3183 3050
rect 3187 3046 3191 3050
rect 3195 3046 3327 3050
rect 3331 3046 3383 3050
rect 3387 3046 3591 3050
rect 3595 3046 3619 3050
rect 1849 3045 3619 3046
rect 3625 3045 3626 3051
rect 96 2981 97 2987
rect 103 2986 1855 2987
rect 103 2982 111 2986
rect 115 2982 143 2986
rect 147 2982 159 2986
rect 163 2982 231 2986
rect 235 2982 319 2986
rect 323 2982 335 2986
rect 339 2982 447 2986
rect 451 2982 487 2986
rect 491 2982 559 2986
rect 563 2982 647 2986
rect 651 2982 671 2986
rect 675 2982 799 2986
rect 803 2982 943 2986
rect 947 2982 1079 2986
rect 1083 2982 1199 2986
rect 1203 2982 1311 2986
rect 1315 2982 1423 2986
rect 1427 2982 1535 2986
rect 1539 2982 1647 2986
rect 1651 2982 1831 2986
rect 1835 2982 1855 2986
rect 103 2981 1855 2982
rect 1861 2981 1862 2987
rect 1854 2957 1855 2963
rect 1861 2962 3631 2963
rect 1861 2958 1871 2962
rect 1875 2958 2127 2962
rect 2131 2958 2207 2962
rect 2211 2958 2287 2962
rect 2291 2958 2343 2962
rect 2347 2958 2367 2962
rect 2371 2958 2447 2962
rect 2451 2958 2487 2962
rect 2491 2958 2527 2962
rect 2531 2958 2607 2962
rect 2611 2958 2631 2962
rect 2635 2958 2695 2962
rect 2699 2958 2775 2962
rect 2779 2958 2791 2962
rect 2795 2958 2911 2962
rect 2915 2958 3039 2962
rect 3043 2958 3047 2962
rect 3051 2958 3183 2962
rect 3187 2958 3191 2962
rect 3195 2958 3335 2962
rect 3339 2958 3495 2962
rect 3499 2958 3591 2962
rect 3595 2958 3631 2962
rect 1861 2957 3631 2958
rect 3637 2957 3638 2963
rect 84 2905 85 2911
rect 91 2910 1843 2911
rect 91 2906 111 2910
rect 115 2906 151 2910
rect 155 2906 311 2910
rect 315 2906 471 2910
rect 475 2906 479 2910
rect 483 2906 631 2910
rect 635 2906 639 2910
rect 643 2906 783 2910
rect 787 2906 791 2910
rect 795 2906 927 2910
rect 931 2906 935 2910
rect 939 2906 1055 2910
rect 1059 2906 1071 2910
rect 1075 2906 1175 2910
rect 1179 2906 1191 2910
rect 1195 2906 1287 2910
rect 1291 2906 1303 2910
rect 1307 2906 1391 2910
rect 1395 2906 1415 2910
rect 1419 2906 1487 2910
rect 1491 2906 1527 2910
rect 1531 2906 1591 2910
rect 1595 2906 1639 2910
rect 1643 2906 1695 2910
rect 1699 2906 1831 2910
rect 1835 2906 1843 2910
rect 91 2905 1843 2906
rect 1849 2905 1850 2911
rect 1842 2881 1843 2887
rect 1849 2886 3619 2887
rect 1849 2882 1871 2886
rect 1875 2882 2047 2886
rect 2051 2882 2119 2886
rect 2123 2882 2135 2886
rect 2139 2882 2199 2886
rect 2203 2882 2239 2886
rect 2243 2882 2279 2886
rect 2283 2882 2343 2886
rect 2347 2882 2359 2886
rect 2363 2882 2439 2886
rect 2443 2882 2463 2886
rect 2467 2882 2519 2886
rect 2523 2882 2591 2886
rect 2595 2882 2599 2886
rect 2603 2882 2687 2886
rect 2691 2882 2727 2886
rect 2731 2882 2783 2886
rect 2787 2882 2879 2886
rect 2883 2882 2903 2886
rect 2907 2882 3031 2886
rect 3035 2882 3175 2886
rect 3179 2882 3191 2886
rect 3195 2882 3327 2886
rect 3331 2882 3359 2886
rect 3363 2882 3487 2886
rect 3491 2882 3503 2886
rect 3507 2882 3591 2886
rect 3595 2882 3619 2886
rect 1849 2881 3619 2882
rect 3625 2881 3626 2887
rect 96 2825 97 2831
rect 103 2830 1855 2831
rect 103 2826 111 2830
rect 115 2826 143 2830
rect 147 2826 159 2830
rect 163 2826 247 2830
rect 251 2826 319 2830
rect 323 2826 383 2830
rect 387 2826 479 2830
rect 483 2826 535 2830
rect 539 2826 639 2830
rect 643 2826 687 2830
rect 691 2826 791 2830
rect 795 2826 847 2830
rect 851 2826 935 2830
rect 939 2826 999 2830
rect 1003 2826 1063 2830
rect 1067 2826 1143 2830
rect 1147 2826 1183 2830
rect 1187 2826 1279 2830
rect 1283 2826 1295 2830
rect 1299 2826 1399 2830
rect 1403 2826 1407 2830
rect 1411 2826 1495 2830
rect 1499 2826 1527 2830
rect 1531 2826 1599 2830
rect 1603 2826 1647 2830
rect 1651 2826 1703 2830
rect 1707 2826 1751 2830
rect 1755 2826 1831 2830
rect 1835 2826 1855 2830
rect 103 2825 1855 2826
rect 1861 2825 1862 2831
rect 1854 2793 1855 2799
rect 1861 2798 3631 2799
rect 1861 2794 1871 2798
rect 1875 2794 1903 2798
rect 1907 2794 2015 2798
rect 2019 2794 2055 2798
rect 2059 2794 2143 2798
rect 2147 2794 2167 2798
rect 2171 2794 2247 2798
rect 2251 2794 2327 2798
rect 2331 2794 2351 2798
rect 2355 2794 2471 2798
rect 2475 2794 2487 2798
rect 2491 2794 2599 2798
rect 2603 2794 2639 2798
rect 2643 2794 2735 2798
rect 2739 2794 2791 2798
rect 2795 2794 2887 2798
rect 2891 2794 2943 2798
rect 2947 2794 3039 2798
rect 3043 2794 3087 2798
rect 3091 2794 3199 2798
rect 3203 2794 3231 2798
rect 3235 2794 3367 2798
rect 3371 2794 3383 2798
rect 3387 2794 3511 2798
rect 3515 2794 3591 2798
rect 3595 2794 3631 2798
rect 1861 2793 3631 2794
rect 3637 2793 3638 2799
rect 84 2745 85 2751
rect 91 2750 1843 2751
rect 91 2746 111 2750
rect 115 2746 135 2750
rect 139 2746 231 2750
rect 235 2746 239 2750
rect 243 2746 367 2750
rect 371 2746 375 2750
rect 379 2746 511 2750
rect 515 2746 527 2750
rect 531 2746 663 2750
rect 667 2746 679 2750
rect 683 2746 815 2750
rect 819 2746 839 2750
rect 843 2746 975 2750
rect 979 2746 991 2750
rect 995 2746 1135 2750
rect 1139 2746 1271 2750
rect 1275 2746 1287 2750
rect 1291 2746 1399 2750
rect 1403 2746 1447 2750
rect 1451 2746 1519 2750
rect 1523 2746 1607 2750
rect 1611 2746 1639 2750
rect 1643 2746 1743 2750
rect 1747 2746 1831 2750
rect 1835 2746 1843 2750
rect 91 2745 1843 2746
rect 1849 2745 1850 2751
rect 1842 2717 1843 2723
rect 1849 2722 3619 2723
rect 1849 2718 1871 2722
rect 1875 2718 1895 2722
rect 1899 2718 2007 2722
rect 2011 2718 2103 2722
rect 2107 2718 2159 2722
rect 2163 2718 2319 2722
rect 2323 2718 2327 2722
rect 2331 2718 2479 2722
rect 2483 2718 2535 2722
rect 2539 2718 2631 2722
rect 2635 2718 2735 2722
rect 2739 2718 2783 2722
rect 2787 2718 2911 2722
rect 2915 2718 2935 2722
rect 2939 2718 3071 2722
rect 3075 2718 3079 2722
rect 3083 2718 3223 2722
rect 3227 2718 3375 2722
rect 3379 2718 3503 2722
rect 3507 2718 3591 2722
rect 3595 2718 3619 2722
rect 1849 2717 3619 2718
rect 3625 2717 3626 2723
rect 96 2661 97 2667
rect 103 2666 1855 2667
rect 103 2662 111 2666
rect 115 2662 143 2666
rect 147 2662 239 2666
rect 243 2662 279 2666
rect 283 2662 375 2666
rect 379 2662 447 2666
rect 451 2662 519 2666
rect 523 2662 623 2666
rect 627 2662 671 2666
rect 675 2662 791 2666
rect 795 2662 823 2666
rect 827 2662 951 2666
rect 955 2662 983 2666
rect 987 2662 1103 2666
rect 1107 2662 1143 2666
rect 1147 2662 1247 2666
rect 1251 2662 1295 2666
rect 1299 2662 1399 2666
rect 1403 2662 1455 2666
rect 1459 2662 1551 2666
rect 1555 2662 1615 2666
rect 1619 2662 1751 2666
rect 1755 2662 1831 2666
rect 1835 2662 1855 2666
rect 103 2661 1855 2662
rect 1861 2661 1862 2667
rect 1854 2633 1855 2639
rect 1861 2638 3631 2639
rect 1861 2634 1871 2638
rect 1875 2634 1903 2638
rect 1907 2634 2055 2638
rect 2059 2634 2111 2638
rect 2115 2634 2263 2638
rect 2267 2634 2335 2638
rect 2339 2634 2495 2638
rect 2499 2634 2543 2638
rect 2547 2634 2743 2638
rect 2747 2634 2751 2638
rect 2755 2634 2919 2638
rect 2923 2634 3015 2638
rect 3019 2634 3079 2638
rect 3083 2634 3231 2638
rect 3235 2634 3287 2638
rect 3291 2634 3383 2638
rect 3387 2634 3511 2638
rect 3515 2634 3591 2638
rect 3595 2634 3631 2638
rect 1861 2633 3631 2634
rect 3637 2633 3638 2639
rect 84 2581 85 2587
rect 91 2586 1843 2587
rect 91 2582 111 2586
rect 115 2582 135 2586
rect 139 2582 223 2586
rect 227 2582 271 2586
rect 275 2582 367 2586
rect 371 2582 439 2586
rect 443 2582 527 2586
rect 531 2582 615 2586
rect 619 2582 703 2586
rect 707 2582 783 2586
rect 787 2582 879 2586
rect 883 2582 943 2586
rect 947 2582 1047 2586
rect 1051 2582 1095 2586
rect 1099 2582 1207 2586
rect 1211 2582 1239 2586
rect 1243 2582 1359 2586
rect 1363 2582 1391 2586
rect 1395 2582 1511 2586
rect 1515 2582 1543 2586
rect 1547 2582 1671 2586
rect 1675 2582 1831 2586
rect 1835 2582 1843 2586
rect 91 2581 1843 2582
rect 1849 2581 1850 2587
rect 1842 2557 1843 2563
rect 1849 2562 3619 2563
rect 1849 2558 1871 2562
rect 1875 2558 1895 2562
rect 1899 2558 2007 2562
rect 2011 2558 2047 2562
rect 2051 2558 2159 2562
rect 2163 2558 2255 2562
rect 2259 2558 2319 2562
rect 2323 2558 2471 2562
rect 2475 2558 2487 2562
rect 2491 2558 2623 2562
rect 2627 2558 2743 2562
rect 2747 2558 2759 2562
rect 2763 2558 2887 2562
rect 2891 2558 3007 2562
rect 3011 2558 3119 2562
rect 3123 2558 3223 2562
rect 3227 2558 3279 2562
rect 3283 2558 3319 2562
rect 3323 2558 3423 2562
rect 3427 2558 3503 2562
rect 3507 2558 3591 2562
rect 3595 2558 3619 2562
rect 1849 2557 3619 2558
rect 3625 2557 3626 2563
rect 96 2501 97 2507
rect 103 2506 1855 2507
rect 103 2502 111 2506
rect 115 2502 143 2506
rect 147 2502 223 2506
rect 227 2502 231 2506
rect 235 2502 303 2506
rect 307 2502 375 2506
rect 379 2502 391 2506
rect 395 2502 511 2506
rect 515 2502 535 2506
rect 539 2502 647 2506
rect 651 2502 711 2506
rect 715 2502 783 2506
rect 787 2502 887 2506
rect 891 2502 927 2506
rect 931 2502 1055 2506
rect 1059 2502 1063 2506
rect 1067 2502 1191 2506
rect 1195 2502 1215 2506
rect 1219 2502 1311 2506
rect 1315 2502 1367 2506
rect 1371 2502 1431 2506
rect 1435 2502 1519 2506
rect 1523 2502 1551 2506
rect 1555 2502 1671 2506
rect 1675 2502 1679 2506
rect 1683 2502 1831 2506
rect 1835 2502 1855 2506
rect 103 2501 1855 2502
rect 1861 2501 1862 2507
rect 1854 2473 1855 2479
rect 1861 2478 3631 2479
rect 1861 2474 1871 2478
rect 1875 2474 1903 2478
rect 1907 2474 1999 2478
rect 2003 2474 2015 2478
rect 2019 2474 2127 2478
rect 2131 2474 2167 2478
rect 2171 2474 2263 2478
rect 2267 2474 2327 2478
rect 2331 2474 2407 2478
rect 2411 2474 2479 2478
rect 2483 2474 2551 2478
rect 2555 2474 2631 2478
rect 2635 2474 2703 2478
rect 2707 2474 2767 2478
rect 2771 2474 2863 2478
rect 2867 2474 2895 2478
rect 2899 2474 3015 2478
rect 3019 2474 3023 2478
rect 3027 2474 3127 2478
rect 3131 2474 3191 2478
rect 3195 2474 3231 2478
rect 3235 2474 3327 2478
rect 3331 2474 3359 2478
rect 3363 2474 3431 2478
rect 3435 2474 3511 2478
rect 3515 2474 3591 2478
rect 3595 2474 3631 2478
rect 1861 2473 3631 2474
rect 3637 2473 3638 2479
rect 84 2413 85 2419
rect 91 2418 1843 2419
rect 91 2414 111 2418
rect 115 2414 135 2418
rect 139 2414 215 2418
rect 219 2414 295 2418
rect 299 2414 383 2418
rect 387 2414 503 2418
rect 507 2414 639 2418
rect 643 2414 775 2418
rect 779 2414 919 2418
rect 923 2414 1055 2418
rect 1059 2414 1063 2418
rect 1067 2414 1143 2418
rect 1147 2414 1183 2418
rect 1187 2414 1223 2418
rect 1227 2414 1303 2418
rect 1307 2414 1383 2418
rect 1387 2414 1423 2418
rect 1427 2414 1463 2418
rect 1467 2414 1543 2418
rect 1547 2414 1663 2418
rect 1667 2414 1831 2418
rect 1835 2414 1843 2418
rect 91 2413 1843 2414
rect 1849 2413 1850 2419
rect 1842 2393 1843 2399
rect 1849 2398 3619 2399
rect 1849 2394 1871 2398
rect 1875 2394 1991 2398
rect 1995 2394 2119 2398
rect 2123 2394 2143 2398
rect 2147 2394 2239 2398
rect 2243 2394 2255 2398
rect 2259 2394 2343 2398
rect 2347 2394 2399 2398
rect 2403 2394 2455 2398
rect 2459 2394 2543 2398
rect 2547 2394 2575 2398
rect 2579 2394 2695 2398
rect 2699 2394 2703 2398
rect 2707 2394 2847 2398
rect 2851 2394 2855 2398
rect 2859 2394 3007 2398
rect 3011 2394 3015 2398
rect 3019 2394 3175 2398
rect 3179 2394 3183 2398
rect 3187 2394 3351 2398
rect 3355 2394 3503 2398
rect 3507 2394 3591 2398
rect 3595 2394 3619 2398
rect 1849 2393 3619 2394
rect 3625 2393 3626 2399
rect 96 2329 97 2335
rect 103 2334 1855 2335
rect 103 2330 111 2334
rect 115 2330 359 2334
rect 363 2330 439 2334
rect 443 2330 519 2334
rect 523 2330 599 2334
rect 603 2330 679 2334
rect 683 2330 759 2334
rect 763 2330 839 2334
rect 843 2330 919 2334
rect 923 2330 999 2334
rect 1003 2330 1071 2334
rect 1075 2330 1079 2334
rect 1083 2330 1151 2334
rect 1155 2330 1159 2334
rect 1163 2330 1231 2334
rect 1235 2330 1239 2334
rect 1243 2330 1311 2334
rect 1315 2330 1319 2334
rect 1323 2330 1391 2334
rect 1395 2330 1471 2334
rect 1475 2330 1831 2334
rect 1835 2330 1855 2334
rect 103 2329 1855 2330
rect 1861 2329 1862 2335
rect 1854 2313 1855 2319
rect 1861 2318 3631 2319
rect 1861 2314 1871 2318
rect 1875 2314 2151 2318
rect 2155 2314 2247 2318
rect 2251 2314 2279 2318
rect 2283 2314 2351 2318
rect 2355 2314 2359 2318
rect 2363 2314 2439 2318
rect 2443 2314 2463 2318
rect 2467 2314 2519 2318
rect 2523 2314 2583 2318
rect 2587 2314 2599 2318
rect 2603 2314 2679 2318
rect 2683 2314 2711 2318
rect 2715 2314 2759 2318
rect 2763 2314 2847 2318
rect 2851 2314 2855 2318
rect 2859 2314 2935 2318
rect 2939 2314 3015 2318
rect 3019 2314 3183 2318
rect 3187 2314 3359 2318
rect 3363 2314 3511 2318
rect 3515 2314 3591 2318
rect 3595 2314 3631 2318
rect 1861 2313 3631 2314
rect 3637 2313 3638 2319
rect 84 2253 85 2259
rect 91 2258 1843 2259
rect 91 2254 111 2258
rect 115 2254 351 2258
rect 355 2254 375 2258
rect 379 2254 431 2258
rect 435 2254 455 2258
rect 459 2254 511 2258
rect 515 2254 535 2258
rect 539 2254 591 2258
rect 595 2254 615 2258
rect 619 2254 671 2258
rect 675 2254 695 2258
rect 699 2254 751 2258
rect 755 2254 775 2258
rect 779 2254 831 2258
rect 835 2254 855 2258
rect 859 2254 911 2258
rect 915 2254 935 2258
rect 939 2254 991 2258
rect 995 2254 1015 2258
rect 1019 2254 1071 2258
rect 1075 2254 1095 2258
rect 1099 2254 1151 2258
rect 1155 2254 1175 2258
rect 1179 2254 1231 2258
rect 1235 2254 1255 2258
rect 1259 2254 1311 2258
rect 1315 2254 1831 2258
rect 1835 2254 1843 2258
rect 91 2253 1843 2254
rect 1849 2253 1850 2259
rect 1842 2237 1843 2243
rect 1849 2242 3619 2243
rect 1849 2238 1871 2242
rect 1875 2238 2271 2242
rect 2275 2238 2311 2242
rect 2315 2238 2351 2242
rect 2355 2238 2399 2242
rect 2403 2238 2431 2242
rect 2435 2238 2495 2242
rect 2499 2238 2511 2242
rect 2515 2238 2591 2242
rect 2595 2238 2599 2242
rect 2603 2238 2671 2242
rect 2675 2238 2719 2242
rect 2723 2238 2751 2242
rect 2755 2238 2839 2242
rect 2843 2238 2855 2242
rect 2859 2238 2927 2242
rect 2931 2238 3007 2242
rect 3011 2238 3175 2242
rect 3179 2238 3351 2242
rect 3355 2238 3503 2242
rect 3507 2238 3591 2242
rect 3595 2238 3619 2242
rect 1849 2237 3619 2238
rect 3625 2237 3626 2243
rect 96 2165 97 2171
rect 103 2170 1855 2171
rect 103 2166 111 2170
rect 115 2166 311 2170
rect 315 2166 383 2170
rect 387 2166 407 2170
rect 411 2166 463 2170
rect 467 2166 503 2170
rect 507 2166 543 2170
rect 547 2166 599 2170
rect 603 2166 623 2170
rect 627 2166 687 2170
rect 691 2166 703 2170
rect 707 2166 775 2170
rect 779 2166 783 2170
rect 787 2166 863 2170
rect 867 2166 943 2170
rect 947 2166 951 2170
rect 955 2166 1023 2170
rect 1027 2166 1039 2170
rect 1043 2166 1103 2170
rect 1107 2166 1127 2170
rect 1131 2166 1183 2170
rect 1187 2166 1223 2170
rect 1227 2166 1263 2170
rect 1267 2166 1831 2170
rect 1835 2166 1855 2170
rect 103 2165 1855 2166
rect 1861 2165 1862 2171
rect 1854 2163 1862 2165
rect 1854 2157 1855 2163
rect 1861 2162 3631 2163
rect 1861 2158 1871 2162
rect 1875 2158 1903 2162
rect 1907 2158 1983 2162
rect 1987 2158 2111 2162
rect 2115 2158 2247 2162
rect 2251 2158 2319 2162
rect 2323 2158 2391 2162
rect 2395 2158 2407 2162
rect 2411 2158 2503 2162
rect 2507 2158 2543 2162
rect 2547 2158 2607 2162
rect 2611 2158 2695 2162
rect 2699 2158 2727 2162
rect 2731 2158 2847 2162
rect 2851 2158 2863 2162
rect 2867 2158 3007 2162
rect 3011 2158 3015 2162
rect 3019 2158 3175 2162
rect 3179 2158 3183 2162
rect 3187 2158 3351 2162
rect 3355 2158 3359 2162
rect 3363 2158 3511 2162
rect 3515 2158 3591 2162
rect 3595 2158 3631 2162
rect 1861 2157 3631 2158
rect 3637 2157 3638 2163
rect 84 2077 85 2083
rect 91 2082 1843 2083
rect 91 2078 111 2082
rect 115 2078 207 2082
rect 211 2078 303 2082
rect 307 2078 327 2082
rect 331 2078 399 2082
rect 403 2078 447 2082
rect 451 2078 495 2082
rect 499 2078 575 2082
rect 579 2078 591 2082
rect 595 2078 679 2082
rect 683 2078 703 2082
rect 707 2078 767 2082
rect 771 2078 823 2082
rect 827 2078 855 2082
rect 859 2078 943 2082
rect 947 2078 1031 2082
rect 1035 2078 1063 2082
rect 1067 2078 1119 2082
rect 1123 2078 1175 2082
rect 1179 2078 1215 2082
rect 1219 2078 1279 2082
rect 1283 2078 1375 2082
rect 1379 2078 1471 2082
rect 1475 2078 1567 2082
rect 1571 2078 1663 2082
rect 1667 2078 1743 2082
rect 1747 2078 1831 2082
rect 1835 2078 1843 2082
rect 91 2077 1843 2078
rect 1849 2079 1850 2083
rect 1849 2078 3626 2079
rect 1849 2077 1871 2078
rect 1842 2074 1871 2077
rect 1875 2074 1895 2078
rect 1899 2074 1967 2078
rect 1971 2074 1975 2078
rect 1979 2074 2103 2078
rect 2107 2074 2215 2078
rect 2219 2074 2239 2078
rect 2243 2074 2383 2078
rect 2387 2074 2447 2078
rect 2451 2074 2535 2078
rect 2539 2074 2655 2078
rect 2659 2074 2687 2078
rect 2691 2074 2839 2078
rect 2843 2074 2999 2078
rect 3003 2074 3143 2078
rect 3147 2074 3167 2078
rect 3171 2074 3271 2078
rect 3275 2074 3343 2078
rect 3347 2074 3399 2078
rect 3403 2074 3503 2078
rect 3507 2074 3591 2078
rect 3595 2074 3626 2078
rect 1842 2073 3626 2074
rect 96 1997 97 2003
rect 103 2002 1855 2003
rect 103 1998 111 2002
rect 115 1998 191 2002
rect 195 1998 215 2002
rect 219 1998 335 2002
rect 339 1998 351 2002
rect 355 1998 455 2002
rect 459 1998 519 2002
rect 523 1998 583 2002
rect 587 1998 687 2002
rect 691 1998 711 2002
rect 715 1998 831 2002
rect 835 1998 855 2002
rect 859 1998 951 2002
rect 955 1998 1015 2002
rect 1019 1998 1071 2002
rect 1075 1998 1167 2002
rect 1171 1998 1183 2002
rect 1187 1998 1287 2002
rect 1291 1998 1311 2002
rect 1315 1998 1383 2002
rect 1387 1998 1447 2002
rect 1451 1998 1479 2002
rect 1483 1998 1575 2002
rect 1579 1998 1583 2002
rect 1587 1998 1671 2002
rect 1675 1998 1719 2002
rect 1723 1998 1751 2002
rect 1755 1998 1831 2002
rect 1835 1998 1855 2002
rect 103 1997 1855 1998
rect 1861 2002 3638 2003
rect 1861 1998 1871 2002
rect 1875 1998 1959 2002
rect 1963 1998 1975 2002
rect 1979 1998 2079 2002
rect 2083 1998 2199 2002
rect 2203 1998 2223 2002
rect 2227 1998 2319 2002
rect 2323 1998 2447 2002
rect 2451 1998 2455 2002
rect 2459 1998 2583 2002
rect 2587 1998 2663 2002
rect 2667 1998 2743 2002
rect 2747 1998 2847 2002
rect 2851 1998 2919 2002
rect 2923 1998 3007 2002
rect 3011 1998 3119 2002
rect 3123 1998 3151 2002
rect 3155 1998 3279 2002
rect 3283 1998 3327 2002
rect 3331 1998 3407 2002
rect 3411 1998 3511 2002
rect 3515 1998 3591 2002
rect 3595 1998 3638 2002
rect 1861 1997 3638 1998
rect 84 1917 85 1923
rect 91 1922 1843 1923
rect 91 1918 111 1922
rect 115 1918 135 1922
rect 139 1918 183 1922
rect 187 1918 239 1922
rect 243 1918 343 1922
rect 347 1918 375 1922
rect 379 1918 511 1922
rect 515 1918 527 1922
rect 531 1918 679 1922
rect 683 1918 687 1922
rect 691 1918 847 1922
rect 851 1918 1007 1922
rect 1011 1918 1159 1922
rect 1163 1918 1303 1922
rect 1307 1918 1439 1922
rect 1443 1918 1455 1922
rect 1459 1918 1575 1922
rect 1579 1918 1607 1922
rect 1611 1918 1711 1922
rect 1715 1918 1831 1922
rect 1835 1918 1843 1922
rect 91 1917 1843 1918
rect 1849 1919 1850 1923
rect 1849 1918 3626 1919
rect 1849 1917 1871 1918
rect 1842 1914 1871 1917
rect 1875 1914 1951 1918
rect 1955 1914 2063 1918
rect 2067 1914 2071 1918
rect 2075 1914 2151 1918
rect 2155 1914 2191 1918
rect 2195 1914 2239 1918
rect 2243 1914 2311 1918
rect 2315 1914 2319 1918
rect 2323 1914 2399 1918
rect 2403 1914 2439 1918
rect 2443 1914 2487 1918
rect 2491 1914 2575 1918
rect 2579 1914 2663 1918
rect 2667 1914 2735 1918
rect 2739 1914 2759 1918
rect 2763 1914 2871 1918
rect 2875 1914 2911 1918
rect 2915 1914 2991 1918
rect 2995 1914 3111 1918
rect 3115 1914 3119 1918
rect 3123 1914 3247 1918
rect 3251 1914 3319 1918
rect 3323 1914 3383 1918
rect 3387 1914 3503 1918
rect 3507 1914 3591 1918
rect 3595 1914 3626 1918
rect 1842 1913 3626 1914
rect 96 1837 97 1843
rect 103 1842 1855 1843
rect 103 1838 111 1842
rect 115 1838 143 1842
rect 147 1838 247 1842
rect 251 1838 287 1842
rect 291 1838 383 1842
rect 387 1838 471 1842
rect 475 1838 535 1842
rect 539 1838 663 1842
rect 667 1838 695 1842
rect 699 1838 847 1842
rect 851 1838 855 1842
rect 859 1838 1015 1842
rect 1019 1838 1023 1842
rect 1027 1838 1167 1842
rect 1171 1838 1191 1842
rect 1195 1838 1311 1842
rect 1315 1838 1351 1842
rect 1355 1838 1463 1842
rect 1467 1838 1511 1842
rect 1515 1838 1615 1842
rect 1619 1838 1679 1842
rect 1683 1838 1831 1842
rect 1835 1838 1855 1842
rect 103 1837 1855 1838
rect 1861 1837 1862 1843
rect 1854 1821 1855 1827
rect 1861 1826 3631 1827
rect 1861 1822 1871 1826
rect 1875 1822 2071 1826
rect 2075 1822 2095 1826
rect 2099 1822 2159 1826
rect 2163 1822 2239 1826
rect 2243 1822 2247 1826
rect 2251 1822 2327 1826
rect 2331 1822 2399 1826
rect 2403 1822 2407 1826
rect 2411 1822 2495 1826
rect 2499 1822 2559 1826
rect 2563 1822 2583 1826
rect 2587 1822 2671 1826
rect 2675 1822 2719 1826
rect 2723 1822 2767 1826
rect 2771 1822 2879 1826
rect 2883 1822 2999 1826
rect 3003 1822 3031 1826
rect 3035 1822 3127 1826
rect 3131 1822 3175 1826
rect 3179 1822 3255 1826
rect 3259 1822 3319 1826
rect 3323 1822 3391 1826
rect 3395 1822 3471 1826
rect 3475 1822 3511 1826
rect 3515 1822 3591 1826
rect 3595 1822 3631 1826
rect 1861 1821 3631 1822
rect 3637 1821 3638 1827
rect 84 1753 85 1759
rect 91 1758 1843 1759
rect 91 1754 111 1758
rect 115 1754 135 1758
rect 139 1754 215 1758
rect 219 1754 279 1758
rect 283 1754 343 1758
rect 347 1754 463 1758
rect 467 1754 495 1758
rect 499 1754 655 1758
rect 659 1754 663 1758
rect 667 1754 839 1758
rect 843 1754 1007 1758
rect 1011 1754 1015 1758
rect 1019 1754 1167 1758
rect 1171 1754 1183 1758
rect 1187 1754 1319 1758
rect 1323 1754 1343 1758
rect 1347 1754 1463 1758
rect 1467 1754 1503 1758
rect 1507 1754 1607 1758
rect 1611 1754 1671 1758
rect 1675 1754 1743 1758
rect 1747 1754 1831 1758
rect 1835 1754 1843 1758
rect 91 1753 1843 1754
rect 1849 1753 1850 1759
rect 1842 1741 1843 1747
rect 1849 1746 3619 1747
rect 1849 1742 1871 1746
rect 1875 1742 2087 1746
rect 2091 1742 2103 1746
rect 2107 1742 2231 1746
rect 2235 1742 2239 1746
rect 2243 1742 2383 1746
rect 2387 1742 2391 1746
rect 2395 1742 2527 1746
rect 2531 1742 2551 1746
rect 2555 1742 2663 1746
rect 2667 1742 2711 1746
rect 2715 1742 2799 1746
rect 2803 1742 2871 1746
rect 2875 1742 2927 1746
rect 2931 1742 3023 1746
rect 3027 1742 3047 1746
rect 3051 1742 3159 1746
rect 3163 1742 3167 1746
rect 3171 1742 3271 1746
rect 3275 1742 3311 1746
rect 3315 1742 3391 1746
rect 3395 1742 3463 1746
rect 3467 1742 3503 1746
rect 3507 1742 3591 1746
rect 3595 1742 3619 1746
rect 1849 1741 3619 1742
rect 3625 1741 3626 1747
rect 96 1673 97 1679
rect 103 1678 1855 1679
rect 103 1674 111 1678
rect 115 1674 143 1678
rect 147 1674 223 1678
rect 227 1674 295 1678
rect 299 1674 351 1678
rect 355 1674 479 1678
rect 483 1674 503 1678
rect 507 1674 671 1678
rect 675 1674 847 1678
rect 851 1674 855 1678
rect 859 1674 1015 1678
rect 1019 1674 1031 1678
rect 1035 1674 1175 1678
rect 1179 1674 1199 1678
rect 1203 1674 1327 1678
rect 1331 1674 1359 1678
rect 1363 1674 1471 1678
rect 1475 1674 1519 1678
rect 1523 1674 1615 1678
rect 1619 1674 1679 1678
rect 1683 1674 1751 1678
rect 1755 1674 1831 1678
rect 1835 1674 1855 1678
rect 103 1673 1855 1674
rect 1861 1673 1862 1679
rect 1854 1661 1855 1667
rect 1861 1666 3631 1667
rect 1861 1662 1871 1666
rect 1875 1662 1967 1666
rect 1971 1662 2087 1666
rect 2091 1662 2111 1666
rect 2115 1662 2215 1666
rect 2219 1662 2247 1666
rect 2251 1662 2351 1666
rect 2355 1662 2391 1666
rect 2395 1662 2495 1666
rect 2499 1662 2535 1666
rect 2539 1662 2639 1666
rect 2643 1662 2671 1666
rect 2675 1662 2783 1666
rect 2787 1662 2807 1666
rect 2811 1662 2927 1666
rect 2931 1662 2935 1666
rect 2939 1662 3055 1666
rect 3059 1662 3071 1666
rect 3075 1662 3167 1666
rect 3171 1662 3223 1666
rect 3227 1662 3279 1666
rect 3283 1662 3375 1666
rect 3379 1662 3399 1666
rect 3403 1662 3511 1666
rect 3515 1662 3591 1666
rect 3595 1662 3631 1666
rect 1861 1661 3631 1662
rect 3637 1661 3638 1667
rect 84 1597 85 1603
rect 91 1602 1843 1603
rect 91 1598 111 1602
rect 115 1598 135 1602
rect 139 1598 159 1602
rect 163 1598 287 1602
rect 291 1598 423 1602
rect 427 1598 471 1602
rect 475 1598 567 1602
rect 571 1598 663 1602
rect 667 1598 711 1602
rect 715 1598 847 1602
rect 851 1598 983 1602
rect 987 1598 1023 1602
rect 1027 1598 1119 1602
rect 1123 1598 1191 1602
rect 1195 1598 1247 1602
rect 1251 1598 1351 1602
rect 1355 1598 1375 1602
rect 1379 1598 1511 1602
rect 1515 1598 1671 1602
rect 1675 1598 1831 1602
rect 1835 1598 1843 1602
rect 91 1597 1843 1598
rect 1849 1597 1850 1603
rect 1842 1577 1843 1583
rect 1849 1582 3619 1583
rect 1849 1578 1871 1582
rect 1875 1578 1895 1582
rect 1899 1578 1959 1582
rect 1963 1578 2047 1582
rect 2051 1578 2079 1582
rect 2083 1578 2207 1582
rect 2211 1578 2343 1582
rect 2347 1578 2367 1582
rect 2371 1578 2487 1582
rect 2491 1578 2527 1582
rect 2531 1578 2631 1582
rect 2635 1578 2687 1582
rect 2691 1578 2775 1582
rect 2779 1578 2839 1582
rect 2843 1578 2919 1582
rect 2923 1578 2983 1582
rect 2987 1578 3063 1582
rect 3067 1578 3119 1582
rect 3123 1578 3215 1582
rect 3219 1578 3255 1582
rect 3259 1578 3367 1582
rect 3371 1578 3391 1582
rect 3395 1578 3503 1582
rect 3507 1578 3591 1582
rect 3595 1578 3619 1582
rect 1849 1577 3619 1578
rect 3625 1577 3626 1583
rect 96 1517 97 1523
rect 103 1522 1855 1523
rect 103 1518 111 1522
rect 115 1518 167 1522
rect 171 1518 231 1522
rect 235 1518 295 1522
rect 299 1518 375 1522
rect 379 1518 431 1522
rect 435 1518 519 1522
rect 523 1518 575 1522
rect 579 1518 655 1522
rect 659 1518 719 1522
rect 723 1518 783 1522
rect 787 1518 855 1522
rect 859 1518 903 1522
rect 907 1518 991 1522
rect 995 1518 1015 1522
rect 1019 1518 1119 1522
rect 1123 1518 1127 1522
rect 1131 1518 1215 1522
rect 1219 1518 1255 1522
rect 1259 1518 1319 1522
rect 1323 1518 1383 1522
rect 1387 1518 1423 1522
rect 1427 1518 1519 1522
rect 1523 1518 1831 1522
rect 1835 1518 1855 1522
rect 103 1517 1855 1518
rect 1861 1517 1862 1523
rect 1854 1493 1855 1499
rect 1861 1498 3631 1499
rect 1861 1494 1871 1498
rect 1875 1494 1903 1498
rect 1907 1494 2007 1498
rect 2011 1494 2055 1498
rect 2059 1494 2135 1498
rect 2139 1494 2215 1498
rect 2219 1494 2271 1498
rect 2275 1494 2375 1498
rect 2379 1494 2415 1498
rect 2419 1494 2535 1498
rect 2539 1494 2567 1498
rect 2571 1494 2695 1498
rect 2699 1494 2719 1498
rect 2723 1494 2847 1498
rect 2851 1494 2879 1498
rect 2883 1494 2991 1498
rect 2995 1494 3039 1498
rect 3043 1494 3127 1498
rect 3131 1494 3199 1498
rect 3203 1494 3263 1498
rect 3267 1494 3367 1498
rect 3371 1494 3399 1498
rect 3403 1494 3511 1498
rect 3515 1494 3591 1498
rect 3595 1494 3631 1498
rect 1861 1493 3631 1494
rect 3637 1493 3638 1499
rect 84 1433 85 1439
rect 91 1438 1843 1439
rect 91 1434 111 1438
rect 115 1434 223 1438
rect 227 1434 255 1438
rect 259 1434 351 1438
rect 355 1434 367 1438
rect 371 1434 447 1438
rect 451 1434 511 1438
rect 515 1434 543 1438
rect 547 1434 631 1438
rect 635 1434 647 1438
rect 651 1434 719 1438
rect 723 1434 775 1438
rect 779 1434 807 1438
rect 811 1434 895 1438
rect 899 1434 919 1438
rect 923 1434 1007 1438
rect 1011 1434 1047 1438
rect 1051 1434 1111 1438
rect 1115 1434 1207 1438
rect 1211 1434 1311 1438
rect 1315 1434 1383 1438
rect 1387 1434 1415 1438
rect 1419 1434 1575 1438
rect 1579 1434 1743 1438
rect 1747 1434 1831 1438
rect 1835 1434 1843 1438
rect 91 1433 1843 1434
rect 1849 1433 1850 1439
rect 1842 1417 1843 1423
rect 1849 1422 3619 1423
rect 1849 1418 1871 1422
rect 1875 1418 1895 1422
rect 1899 1418 1999 1422
rect 2003 1418 2023 1422
rect 2027 1418 2127 1422
rect 2131 1418 2167 1422
rect 2171 1418 2263 1422
rect 2267 1418 2303 1422
rect 2307 1418 2407 1422
rect 2411 1418 2431 1422
rect 2435 1418 2551 1422
rect 2555 1418 2559 1422
rect 2563 1418 2671 1422
rect 2675 1418 2711 1422
rect 2715 1418 2791 1422
rect 2795 1418 2871 1422
rect 2875 1418 2911 1422
rect 2915 1418 3031 1422
rect 3035 1418 3191 1422
rect 3195 1418 3359 1422
rect 3363 1418 3503 1422
rect 3507 1418 3591 1422
rect 3595 1418 3619 1422
rect 1849 1417 3619 1418
rect 3625 1417 3626 1423
rect 96 1357 97 1363
rect 103 1362 1855 1363
rect 103 1358 111 1362
rect 115 1358 263 1362
rect 267 1358 359 1362
rect 363 1358 455 1362
rect 459 1358 471 1362
rect 475 1358 551 1362
rect 555 1358 591 1362
rect 595 1358 639 1362
rect 643 1358 727 1362
rect 731 1358 815 1362
rect 819 1358 863 1362
rect 867 1358 927 1362
rect 931 1358 1007 1362
rect 1011 1358 1055 1362
rect 1059 1358 1143 1362
rect 1147 1358 1215 1362
rect 1219 1358 1279 1362
rect 1283 1358 1391 1362
rect 1395 1358 1407 1362
rect 1411 1358 1527 1362
rect 1531 1358 1583 1362
rect 1587 1358 1647 1362
rect 1651 1358 1751 1362
rect 1755 1358 1831 1362
rect 1835 1358 1855 1362
rect 103 1357 1855 1358
rect 1861 1357 1862 1363
rect 1854 1333 1855 1339
rect 1861 1338 3631 1339
rect 1861 1334 1871 1338
rect 1875 1334 1903 1338
rect 1907 1334 1927 1338
rect 1931 1334 2031 1338
rect 2035 1334 2047 1338
rect 2051 1334 2175 1338
rect 2179 1334 2183 1338
rect 2187 1334 2311 1338
rect 2315 1334 2319 1338
rect 2323 1334 2439 1338
rect 2443 1334 2455 1338
rect 2459 1334 2559 1338
rect 2563 1334 2591 1338
rect 2595 1334 2679 1338
rect 2683 1334 2719 1338
rect 2723 1334 2799 1338
rect 2803 1334 2839 1338
rect 2843 1334 2919 1338
rect 2923 1334 2951 1338
rect 2955 1334 3063 1338
rect 3067 1334 3183 1338
rect 3187 1334 3591 1338
rect 3595 1334 3631 1338
rect 1861 1333 3631 1334
rect 3637 1333 3638 1339
rect 84 1277 85 1283
rect 91 1282 1843 1283
rect 91 1278 111 1282
rect 115 1278 311 1282
rect 315 1278 351 1282
rect 355 1278 415 1282
rect 419 1278 463 1282
rect 467 1278 535 1282
rect 539 1278 583 1282
rect 587 1278 671 1282
rect 675 1278 719 1282
rect 723 1278 815 1282
rect 819 1278 855 1282
rect 859 1278 959 1282
rect 963 1278 999 1282
rect 1003 1278 1103 1282
rect 1107 1278 1135 1282
rect 1139 1278 1239 1282
rect 1243 1278 1271 1282
rect 1275 1278 1375 1282
rect 1379 1278 1399 1282
rect 1403 1278 1503 1282
rect 1507 1278 1519 1282
rect 1523 1278 1631 1282
rect 1635 1278 1639 1282
rect 1643 1278 1743 1282
rect 1747 1278 1831 1282
rect 1835 1278 1843 1282
rect 91 1277 1843 1278
rect 1849 1277 1850 1283
rect 1842 1249 1843 1255
rect 1849 1254 3619 1255
rect 1849 1250 1871 1254
rect 1875 1250 1895 1254
rect 1899 1250 1919 1254
rect 1923 1250 2039 1254
rect 2043 1250 2071 1254
rect 2075 1250 2175 1254
rect 2179 1250 2271 1254
rect 2275 1250 2311 1254
rect 2315 1250 2447 1254
rect 2451 1250 2471 1254
rect 2475 1250 2583 1254
rect 2587 1250 2663 1254
rect 2667 1250 2711 1254
rect 2715 1250 2831 1254
rect 2835 1250 2847 1254
rect 2851 1250 2943 1254
rect 2947 1250 3023 1254
rect 3027 1250 3055 1254
rect 3059 1250 3175 1254
rect 3179 1250 3191 1254
rect 3195 1250 3359 1254
rect 3363 1250 3503 1254
rect 3507 1250 3591 1254
rect 3595 1250 3619 1254
rect 1849 1249 3619 1250
rect 3625 1249 3626 1255
rect 96 1201 97 1207
rect 103 1206 1855 1207
rect 103 1202 111 1206
rect 115 1202 239 1206
rect 243 1202 319 1206
rect 323 1202 415 1206
rect 419 1202 423 1206
rect 427 1202 543 1206
rect 547 1202 591 1206
rect 595 1202 679 1206
rect 683 1202 759 1206
rect 763 1202 823 1206
rect 827 1202 927 1206
rect 931 1202 967 1206
rect 971 1202 1079 1206
rect 1083 1202 1111 1206
rect 1115 1202 1223 1206
rect 1227 1202 1247 1206
rect 1251 1202 1367 1206
rect 1371 1202 1383 1206
rect 1387 1202 1503 1206
rect 1507 1202 1511 1206
rect 1515 1202 1639 1206
rect 1643 1202 1751 1206
rect 1755 1202 1831 1206
rect 1835 1202 1855 1206
rect 103 1201 1855 1202
rect 1861 1201 1862 1207
rect 1854 1169 1855 1175
rect 1861 1174 3631 1175
rect 1861 1170 1871 1174
rect 1875 1170 1903 1174
rect 1907 1170 1983 1174
rect 1987 1170 2079 1174
rect 2083 1170 2087 1174
rect 2091 1170 2215 1174
rect 2219 1170 2279 1174
rect 2283 1170 2367 1174
rect 2371 1170 2479 1174
rect 2483 1170 2527 1174
rect 2531 1170 2671 1174
rect 2675 1170 2687 1174
rect 2691 1170 2839 1174
rect 2843 1170 2855 1174
rect 2859 1170 2983 1174
rect 2987 1170 3031 1174
rect 3035 1170 3127 1174
rect 3131 1170 3199 1174
rect 3203 1170 3263 1174
rect 3267 1170 3367 1174
rect 3371 1170 3399 1174
rect 3403 1170 3511 1174
rect 3515 1170 3591 1174
rect 3595 1170 3631 1174
rect 1861 1169 3631 1170
rect 3637 1169 3638 1175
rect 84 1121 85 1127
rect 91 1126 1843 1127
rect 91 1122 111 1126
rect 115 1122 143 1126
rect 147 1122 231 1126
rect 235 1122 279 1126
rect 283 1122 407 1126
rect 411 1122 423 1126
rect 427 1122 567 1126
rect 571 1122 583 1126
rect 587 1122 711 1126
rect 715 1122 751 1126
rect 755 1122 847 1126
rect 851 1122 919 1126
rect 923 1122 975 1126
rect 979 1122 1071 1126
rect 1075 1122 1103 1126
rect 1107 1122 1215 1126
rect 1219 1122 1223 1126
rect 1227 1122 1343 1126
rect 1347 1122 1359 1126
rect 1363 1122 1471 1126
rect 1475 1122 1495 1126
rect 1499 1122 1631 1126
rect 1635 1122 1743 1126
rect 1747 1122 1831 1126
rect 1835 1122 1843 1126
rect 91 1121 1843 1122
rect 1849 1121 1850 1127
rect 1842 1085 1843 1091
rect 1849 1090 3619 1091
rect 1849 1086 1871 1090
rect 1875 1086 1895 1090
rect 1899 1086 1975 1090
rect 1979 1086 2079 1090
rect 2083 1086 2167 1090
rect 2171 1086 2207 1090
rect 2211 1086 2255 1090
rect 2259 1086 2359 1090
rect 2363 1086 2479 1090
rect 2483 1086 2519 1090
rect 2523 1086 2607 1090
rect 2611 1086 2679 1090
rect 2683 1086 2751 1090
rect 2755 1086 2831 1090
rect 2835 1086 2895 1090
rect 2899 1086 2975 1090
rect 2979 1086 3047 1090
rect 3051 1086 3119 1090
rect 3123 1086 3207 1090
rect 3211 1086 3255 1090
rect 3259 1086 3367 1090
rect 3371 1086 3391 1090
rect 3395 1086 3503 1090
rect 3507 1086 3591 1090
rect 3595 1086 3619 1090
rect 1849 1085 3619 1086
rect 3625 1085 3626 1091
rect 96 1037 97 1043
rect 103 1042 1855 1043
rect 103 1038 111 1042
rect 115 1038 143 1042
rect 147 1038 151 1042
rect 155 1038 263 1042
rect 267 1038 287 1042
rect 291 1038 407 1042
rect 411 1038 431 1042
rect 435 1038 551 1042
rect 555 1038 575 1042
rect 579 1038 687 1042
rect 691 1038 719 1042
rect 723 1038 807 1042
rect 811 1038 855 1042
rect 859 1038 927 1042
rect 931 1038 983 1042
rect 987 1038 1039 1042
rect 1043 1038 1111 1042
rect 1115 1038 1143 1042
rect 1147 1038 1231 1042
rect 1235 1038 1247 1042
rect 1251 1038 1351 1042
rect 1355 1038 1359 1042
rect 1363 1038 1479 1042
rect 1483 1038 1831 1042
rect 1835 1038 1855 1042
rect 103 1037 1855 1038
rect 1861 1037 1862 1043
rect 1854 1009 1855 1015
rect 1861 1014 3631 1015
rect 1861 1010 1871 1014
rect 1875 1010 2175 1014
rect 2179 1010 2263 1014
rect 2267 1010 2303 1014
rect 2307 1010 2367 1014
rect 2371 1010 2383 1014
rect 2387 1010 2471 1014
rect 2475 1010 2487 1014
rect 2491 1010 2567 1014
rect 2571 1010 2615 1014
rect 2619 1010 2671 1014
rect 2675 1010 2759 1014
rect 2763 1010 2783 1014
rect 2787 1010 2903 1014
rect 2907 1010 2911 1014
rect 2915 1010 3055 1014
rect 3059 1010 3207 1014
rect 3211 1010 3215 1014
rect 3219 1010 3367 1014
rect 3371 1010 3375 1014
rect 3379 1010 3511 1014
rect 3515 1010 3591 1014
rect 3595 1010 3631 1014
rect 1861 1009 3631 1010
rect 3637 1009 3638 1015
rect 84 953 85 959
rect 91 958 1843 959
rect 91 954 111 958
rect 115 954 135 958
rect 139 954 215 958
rect 219 954 255 958
rect 259 954 327 958
rect 331 954 399 958
rect 403 954 447 958
rect 451 954 543 958
rect 547 954 567 958
rect 571 954 679 958
rect 683 954 687 958
rect 691 954 799 958
rect 803 954 911 958
rect 915 954 919 958
rect 923 954 1015 958
rect 1019 954 1031 958
rect 1035 954 1119 958
rect 1123 954 1135 958
rect 1139 954 1223 958
rect 1227 954 1239 958
rect 1243 954 1327 958
rect 1331 954 1351 958
rect 1355 954 1831 958
rect 1835 954 1843 958
rect 91 953 1843 954
rect 1849 953 1850 959
rect 1842 925 1843 931
rect 1849 930 3619 931
rect 1849 926 1871 930
rect 1875 926 2279 930
rect 2283 926 2295 930
rect 2299 926 2359 930
rect 2363 926 2375 930
rect 2379 926 2439 930
rect 2443 926 2463 930
rect 2467 926 2519 930
rect 2523 926 2559 930
rect 2563 926 2607 930
rect 2611 926 2663 930
rect 2667 926 2703 930
rect 2707 926 2775 930
rect 2779 926 2807 930
rect 2811 926 2903 930
rect 2907 926 2911 930
rect 2915 926 3015 930
rect 3019 926 3047 930
rect 3051 926 3111 930
rect 3115 926 3199 930
rect 3203 926 3215 930
rect 3219 926 3319 930
rect 3323 926 3359 930
rect 3363 926 3423 930
rect 3427 926 3503 930
rect 3507 926 3591 930
rect 3595 926 3619 930
rect 1849 925 3619 926
rect 3625 925 3626 931
rect 96 869 97 875
rect 103 874 1855 875
rect 103 870 111 874
rect 115 870 143 874
rect 147 870 223 874
rect 227 870 255 874
rect 259 870 335 874
rect 339 870 399 874
rect 403 870 455 874
rect 459 870 559 874
rect 563 870 575 874
rect 579 870 695 874
rect 699 870 719 874
rect 723 870 807 874
rect 811 870 871 874
rect 875 870 919 874
rect 923 870 1015 874
rect 1019 870 1023 874
rect 1027 870 1127 874
rect 1131 870 1151 874
rect 1155 870 1231 874
rect 1235 870 1279 874
rect 1283 870 1335 874
rect 1339 870 1399 874
rect 1403 870 1519 874
rect 1523 870 1647 874
rect 1651 870 1831 874
rect 1835 870 1855 874
rect 103 869 1855 870
rect 1861 869 1862 875
rect 1854 837 1855 843
rect 1861 842 3631 843
rect 1861 838 1871 842
rect 1875 838 2167 842
rect 2171 838 2247 842
rect 2251 838 2287 842
rect 2291 838 2327 842
rect 2331 838 2367 842
rect 2371 838 2423 842
rect 2427 838 2447 842
rect 2451 838 2527 842
rect 2531 838 2535 842
rect 2539 838 2615 842
rect 2619 838 2655 842
rect 2659 838 2711 842
rect 2715 838 2783 842
rect 2787 838 2815 842
rect 2819 838 2911 842
rect 2915 838 2919 842
rect 2923 838 3023 842
rect 3027 838 3039 842
rect 3043 838 3119 842
rect 3123 838 3159 842
rect 3163 838 3223 842
rect 3227 838 3279 842
rect 3283 838 3327 842
rect 3331 838 3407 842
rect 3411 838 3431 842
rect 3435 838 3511 842
rect 3515 838 3591 842
rect 3595 838 3631 842
rect 1861 837 3631 838
rect 3637 837 3638 843
rect 84 781 85 787
rect 91 786 1843 787
rect 91 782 111 786
rect 115 782 135 786
rect 139 782 247 786
rect 251 782 263 786
rect 267 782 391 786
rect 395 782 431 786
rect 435 782 551 786
rect 555 782 607 786
rect 611 782 711 786
rect 715 782 783 786
rect 787 782 863 786
rect 867 782 951 786
rect 955 782 1007 786
rect 1011 782 1103 786
rect 1107 782 1143 786
rect 1147 782 1247 786
rect 1251 782 1271 786
rect 1275 782 1383 786
rect 1387 782 1391 786
rect 1395 782 1511 786
rect 1515 782 1639 786
rect 1643 782 1743 786
rect 1747 782 1831 786
rect 1835 782 1843 786
rect 91 781 1843 782
rect 1849 781 1850 787
rect 1842 753 1843 759
rect 1849 758 3619 759
rect 1849 754 1871 758
rect 1875 754 1895 758
rect 1899 754 1975 758
rect 1979 754 2071 758
rect 2075 754 2159 758
rect 2163 754 2183 758
rect 2187 754 2239 758
rect 2243 754 2311 758
rect 2315 754 2319 758
rect 2323 754 2415 758
rect 2419 754 2447 758
rect 2451 754 2527 758
rect 2531 754 2591 758
rect 2595 754 2647 758
rect 2651 754 2743 758
rect 2747 754 2775 758
rect 2779 754 2895 758
rect 2899 754 2903 758
rect 2907 754 3031 758
rect 3035 754 3047 758
rect 3051 754 3151 758
rect 3155 754 3199 758
rect 3203 754 3271 758
rect 3275 754 3359 758
rect 3363 754 3399 758
rect 3403 754 3503 758
rect 3507 754 3591 758
rect 3595 754 3619 758
rect 1849 753 3619 754
rect 3625 753 3626 759
rect 96 693 97 699
rect 103 698 1855 699
rect 103 694 111 698
rect 115 694 143 698
rect 147 694 271 698
rect 275 694 295 698
rect 299 694 407 698
rect 411 694 439 698
rect 443 694 527 698
rect 531 694 615 698
rect 619 694 655 698
rect 659 694 783 698
rect 787 694 791 698
rect 795 694 903 698
rect 907 694 959 698
rect 963 694 1023 698
rect 1027 694 1111 698
rect 1115 694 1135 698
rect 1139 694 1247 698
rect 1251 694 1255 698
rect 1259 694 1351 698
rect 1355 694 1391 698
rect 1395 694 1455 698
rect 1459 694 1519 698
rect 1523 694 1559 698
rect 1563 694 1647 698
rect 1651 694 1663 698
rect 1667 694 1751 698
rect 1755 694 1831 698
rect 1835 694 1855 698
rect 103 693 1855 694
rect 1861 693 1862 699
rect 1854 673 1855 679
rect 1861 678 3631 679
rect 1861 674 1871 678
rect 1875 674 1903 678
rect 1907 674 1983 678
rect 1987 674 2079 678
rect 2083 674 2095 678
rect 2099 674 2191 678
rect 2195 674 2295 678
rect 2299 674 2319 678
rect 2323 674 2455 678
rect 2459 674 2479 678
rect 2483 674 2599 678
rect 2603 674 2655 678
rect 2659 674 2751 678
rect 2755 674 2831 678
rect 2835 674 2903 678
rect 2907 674 3007 678
rect 3011 674 3055 678
rect 3059 674 3183 678
rect 3187 674 3207 678
rect 3211 674 3359 678
rect 3363 674 3367 678
rect 3371 674 3511 678
rect 3515 674 3591 678
rect 3595 674 3631 678
rect 1861 673 3631 674
rect 3637 673 3638 679
rect 84 613 85 619
rect 91 618 1843 619
rect 91 614 111 618
rect 115 614 287 618
rect 291 614 311 618
rect 315 614 391 618
rect 395 614 399 618
rect 403 614 471 618
rect 475 614 519 618
rect 523 614 559 618
rect 563 614 647 618
rect 651 614 735 618
rect 739 614 775 618
rect 779 614 823 618
rect 827 614 895 618
rect 899 614 911 618
rect 915 614 999 618
rect 1003 614 1015 618
rect 1019 614 1087 618
rect 1091 614 1127 618
rect 1131 614 1175 618
rect 1179 614 1239 618
rect 1243 614 1263 618
rect 1267 614 1343 618
rect 1347 614 1447 618
rect 1451 614 1551 618
rect 1555 614 1655 618
rect 1659 614 1743 618
rect 1747 614 1831 618
rect 1835 614 1843 618
rect 91 613 1843 614
rect 1849 613 1850 619
rect 1842 593 1843 599
rect 1849 598 3619 599
rect 1849 594 1871 598
rect 1875 594 1895 598
rect 1899 594 1975 598
rect 1979 594 2087 598
rect 2091 594 2215 598
rect 2219 594 2287 598
rect 2291 594 2351 598
rect 2355 594 2471 598
rect 2475 594 2495 598
rect 2499 594 2647 598
rect 2651 594 2807 598
rect 2811 594 2823 598
rect 2827 594 2975 598
rect 2979 594 2999 598
rect 3003 594 3151 598
rect 3155 594 3175 598
rect 3179 594 3335 598
rect 3339 594 3351 598
rect 3355 594 3503 598
rect 3507 594 3591 598
rect 3595 594 3619 598
rect 1849 593 3619 594
rect 3625 593 3626 599
rect 96 525 97 531
rect 103 530 1855 531
rect 103 526 111 530
rect 115 526 239 530
rect 243 526 319 530
rect 323 526 343 530
rect 347 526 399 530
rect 403 526 439 530
rect 443 526 479 530
rect 483 526 535 530
rect 539 526 567 530
rect 571 526 631 530
rect 635 526 655 530
rect 659 526 719 530
rect 723 526 743 530
rect 747 526 807 530
rect 811 526 831 530
rect 835 526 895 530
rect 899 526 919 530
rect 923 526 983 530
rect 987 526 1007 530
rect 1011 526 1071 530
rect 1075 526 1095 530
rect 1099 526 1159 530
rect 1163 526 1183 530
rect 1187 526 1247 530
rect 1251 526 1271 530
rect 1275 526 1831 530
rect 1835 526 1855 530
rect 103 525 1855 526
rect 1861 525 1862 531
rect 1854 523 1862 525
rect 1854 517 1855 523
rect 1861 522 3631 523
rect 1861 518 1871 522
rect 1875 518 1903 522
rect 1907 518 1983 522
rect 1987 518 2095 522
rect 2099 518 2151 522
rect 2155 518 2223 522
rect 2227 518 2231 522
rect 2235 518 2327 522
rect 2331 518 2359 522
rect 2363 518 2431 522
rect 2435 518 2503 522
rect 2507 518 2551 522
rect 2555 518 2655 522
rect 2659 518 2687 522
rect 2691 518 2815 522
rect 2819 518 2839 522
rect 2843 518 2983 522
rect 2987 518 2999 522
rect 3003 518 3159 522
rect 3163 518 3175 522
rect 3179 518 3343 522
rect 3347 518 3351 522
rect 3355 518 3511 522
rect 3515 518 3591 522
rect 3595 518 3631 522
rect 1861 517 3631 518
rect 3637 517 3638 523
rect 84 441 85 447
rect 91 446 1843 447
rect 91 442 111 446
rect 115 442 135 446
rect 139 442 231 446
rect 235 442 247 446
rect 251 442 335 446
rect 339 442 375 446
rect 379 442 431 446
rect 435 442 495 446
rect 499 442 527 446
rect 531 442 607 446
rect 611 442 623 446
rect 627 442 711 446
rect 715 442 719 446
rect 723 442 799 446
rect 803 442 823 446
rect 827 442 887 446
rect 891 442 919 446
rect 923 442 975 446
rect 979 442 1007 446
rect 1011 442 1063 446
rect 1067 442 1103 446
rect 1107 442 1151 446
rect 1155 442 1199 446
rect 1203 442 1239 446
rect 1243 442 1295 446
rect 1299 442 1831 446
rect 1835 442 1843 446
rect 91 441 1843 442
rect 1849 443 1850 447
rect 1849 442 3626 443
rect 1849 441 1871 442
rect 1842 438 1871 441
rect 1875 438 2143 442
rect 2147 438 2223 442
rect 2227 438 2319 442
rect 2323 438 2335 442
rect 2339 438 2415 442
rect 2419 438 2423 442
rect 2427 438 2495 442
rect 2499 438 2543 442
rect 2547 438 2583 442
rect 2587 438 2679 442
rect 2683 438 2687 442
rect 2691 438 2799 442
rect 2803 438 2831 442
rect 2835 438 2927 442
rect 2931 438 2991 442
rect 2995 438 3071 442
rect 3075 438 3167 442
rect 3171 438 3215 442
rect 3219 438 3343 442
rect 3347 438 3367 442
rect 3371 438 3503 442
rect 3507 438 3591 442
rect 3595 438 3626 442
rect 1842 437 3626 438
rect 96 353 97 359
rect 103 358 1855 359
rect 103 354 111 358
rect 115 354 143 358
rect 147 354 247 358
rect 251 354 255 358
rect 259 354 375 358
rect 379 354 383 358
rect 387 354 503 358
rect 507 354 511 358
rect 515 354 615 358
rect 619 354 647 358
rect 651 354 727 358
rect 731 354 775 358
rect 779 354 831 358
rect 835 354 895 358
rect 899 354 927 358
rect 931 354 1007 358
rect 1011 354 1015 358
rect 1019 354 1111 358
rect 1115 354 1119 358
rect 1123 354 1207 358
rect 1211 354 1223 358
rect 1227 354 1303 358
rect 1307 354 1327 358
rect 1331 354 1439 358
rect 1443 354 1831 358
rect 1835 354 1855 358
rect 103 353 1855 354
rect 1861 358 3638 359
rect 1861 354 1871 358
rect 1875 354 2079 358
rect 2083 354 2167 358
rect 2171 354 2263 358
rect 2267 354 2343 358
rect 2347 354 2375 358
rect 2379 354 2423 358
rect 2427 354 2503 358
rect 2507 354 2591 358
rect 2595 354 2639 358
rect 2643 354 2695 358
rect 2699 354 2775 358
rect 2779 354 2807 358
rect 2811 354 2911 358
rect 2915 354 2935 358
rect 2939 354 3039 358
rect 3043 354 3079 358
rect 3083 354 3167 358
rect 3171 354 3223 358
rect 3227 354 3287 358
rect 3291 354 3375 358
rect 3379 354 3407 358
rect 3411 354 3511 358
rect 3515 354 3591 358
rect 3595 354 3638 358
rect 1861 353 3638 354
rect 84 269 85 275
rect 91 274 1843 275
rect 91 270 111 274
rect 115 270 135 274
rect 139 270 223 274
rect 227 270 239 274
rect 243 270 335 274
rect 339 270 367 274
rect 371 270 463 274
rect 467 270 503 274
rect 507 270 599 274
rect 603 270 639 274
rect 643 270 735 274
rect 739 270 767 274
rect 771 270 871 274
rect 875 270 887 274
rect 891 270 999 274
rect 1003 270 1007 274
rect 1011 270 1111 274
rect 1115 270 1135 274
rect 1139 270 1215 274
rect 1219 270 1255 274
rect 1259 270 1319 274
rect 1323 270 1367 274
rect 1371 270 1431 274
rect 1435 270 1479 274
rect 1483 270 1599 274
rect 1603 270 1831 274
rect 1835 270 1843 274
rect 91 269 1843 270
rect 1849 274 3626 275
rect 1849 270 1871 274
rect 1875 270 1895 274
rect 1899 270 1983 274
rect 1987 270 2071 274
rect 2075 270 2095 274
rect 2099 270 2159 274
rect 2163 270 2223 274
rect 2227 270 2255 274
rect 2259 270 2359 274
rect 2363 270 2367 274
rect 2371 270 2495 274
rect 2499 270 2503 274
rect 2507 270 2631 274
rect 2635 270 2647 274
rect 2651 270 2767 274
rect 2771 270 2791 274
rect 2795 270 2903 274
rect 2907 270 2935 274
rect 2939 270 3031 274
rect 3035 270 3079 274
rect 3083 270 3159 274
rect 3163 270 3223 274
rect 3227 270 3279 274
rect 3283 270 3375 274
rect 3379 270 3399 274
rect 3403 270 3503 274
rect 3507 270 3591 274
rect 3595 270 3626 274
rect 1849 269 3626 270
rect 1854 181 1855 187
rect 1861 186 3631 187
rect 1861 182 1871 186
rect 1875 182 1903 186
rect 1907 182 1983 186
rect 1987 182 1991 186
rect 1995 182 2087 186
rect 2091 182 2103 186
rect 2107 182 2207 186
rect 2211 182 2231 186
rect 2235 182 2335 186
rect 2339 182 2367 186
rect 2371 182 2463 186
rect 2467 182 2511 186
rect 2515 182 2583 186
rect 2587 182 2655 186
rect 2659 182 2703 186
rect 2707 182 2799 186
rect 2803 182 2815 186
rect 2819 182 2919 186
rect 2923 182 2943 186
rect 2947 182 3015 186
rect 3019 182 3087 186
rect 3091 182 3111 186
rect 3115 182 3207 186
rect 3211 182 3231 186
rect 3235 182 3303 186
rect 3307 182 3383 186
rect 3387 182 3399 186
rect 3403 182 3511 186
rect 3515 182 3591 186
rect 3595 182 3631 186
rect 1861 181 3631 182
rect 3637 181 3638 187
rect 96 161 97 167
rect 103 166 1855 167
rect 103 162 111 166
rect 115 162 159 166
rect 163 162 231 166
rect 235 162 239 166
rect 243 162 319 166
rect 323 162 343 166
rect 347 162 399 166
rect 403 162 471 166
rect 475 162 479 166
rect 483 162 559 166
rect 563 162 607 166
rect 611 162 647 166
rect 651 162 735 166
rect 739 162 743 166
rect 747 162 823 166
rect 827 162 879 166
rect 883 162 911 166
rect 915 162 999 166
rect 1003 162 1015 166
rect 1019 162 1087 166
rect 1091 162 1143 166
rect 1147 162 1167 166
rect 1171 162 1247 166
rect 1251 162 1263 166
rect 1267 162 1335 166
rect 1339 162 1375 166
rect 1379 162 1423 166
rect 1427 162 1487 166
rect 1491 162 1511 166
rect 1515 162 1591 166
rect 1595 162 1607 166
rect 1611 162 1671 166
rect 1675 162 1751 166
rect 1755 162 1831 166
rect 1835 162 1855 166
rect 103 161 1855 162
rect 1861 161 1862 167
rect 1842 105 1843 111
rect 1849 110 3619 111
rect 1849 106 1871 110
rect 1875 106 1895 110
rect 1899 106 1975 110
rect 1979 106 2079 110
rect 2083 106 2199 110
rect 2203 106 2327 110
rect 2331 106 2455 110
rect 2459 106 2575 110
rect 2579 106 2695 110
rect 2699 106 2807 110
rect 2811 106 2911 110
rect 2915 106 3007 110
rect 3011 106 3103 110
rect 3107 106 3199 110
rect 3203 106 3295 110
rect 3299 106 3391 110
rect 3395 106 3591 110
rect 3595 106 3619 110
rect 1849 105 3619 106
rect 3625 105 3626 111
rect 84 85 85 91
rect 91 90 1843 91
rect 91 86 111 90
rect 115 86 151 90
rect 155 86 231 90
rect 235 86 311 90
rect 315 86 391 90
rect 395 86 471 90
rect 475 86 551 90
rect 555 86 639 90
rect 643 86 727 90
rect 731 86 815 90
rect 819 86 903 90
rect 907 86 991 90
rect 995 86 1079 90
rect 1083 86 1159 90
rect 1163 86 1239 90
rect 1243 86 1327 90
rect 1331 86 1415 90
rect 1419 86 1503 90
rect 1507 86 1583 90
rect 1587 86 1663 90
rect 1667 86 1743 90
rect 1747 86 1831 90
rect 1835 86 1843 90
rect 91 85 1843 86
rect 1849 85 1850 91
<< m5c >>
rect 1843 3665 1849 3671
rect 3619 3665 3625 3671
rect 97 3637 103 3643
rect 1855 3637 1861 3643
rect 1855 3589 1861 3595
rect 3631 3589 3637 3595
rect 85 3561 91 3567
rect 1843 3561 1849 3567
rect 1843 3513 1849 3519
rect 3619 3513 3625 3519
rect 97 3477 103 3483
rect 1855 3477 1861 3483
rect 1855 3437 1861 3443
rect 3631 3437 3637 3443
rect 85 3397 91 3403
rect 1843 3397 1849 3403
rect 1843 3361 1849 3367
rect 3619 3361 3625 3367
rect 97 3317 103 3323
rect 1855 3317 1861 3323
rect 1855 3285 1861 3291
rect 3631 3285 3637 3291
rect 85 3241 91 3247
rect 1843 3241 1849 3247
rect 1843 3209 1849 3215
rect 3619 3209 3625 3215
rect 97 3157 103 3163
rect 1855 3157 1861 3163
rect 1855 3133 1861 3139
rect 3631 3133 3637 3139
rect 85 3069 91 3075
rect 1843 3069 1849 3075
rect 1843 3045 1849 3051
rect 3619 3045 3625 3051
rect 97 2981 103 2987
rect 1855 2981 1861 2987
rect 1855 2957 1861 2963
rect 3631 2957 3637 2963
rect 85 2905 91 2911
rect 1843 2905 1849 2911
rect 1843 2881 1849 2887
rect 3619 2881 3625 2887
rect 97 2825 103 2831
rect 1855 2825 1861 2831
rect 1855 2793 1861 2799
rect 3631 2793 3637 2799
rect 85 2745 91 2751
rect 1843 2745 1849 2751
rect 1843 2717 1849 2723
rect 3619 2717 3625 2723
rect 97 2661 103 2667
rect 1855 2661 1861 2667
rect 1855 2633 1861 2639
rect 3631 2633 3637 2639
rect 85 2581 91 2587
rect 1843 2581 1849 2587
rect 1843 2557 1849 2563
rect 3619 2557 3625 2563
rect 97 2501 103 2507
rect 1855 2501 1861 2507
rect 1855 2473 1861 2479
rect 3631 2473 3637 2479
rect 85 2413 91 2419
rect 1843 2413 1849 2419
rect 1843 2393 1849 2399
rect 3619 2393 3625 2399
rect 97 2329 103 2335
rect 1855 2329 1861 2335
rect 1855 2313 1861 2319
rect 3631 2313 3637 2319
rect 85 2253 91 2259
rect 1843 2253 1849 2259
rect 1843 2237 1849 2243
rect 3619 2237 3625 2243
rect 97 2165 103 2171
rect 1855 2165 1861 2171
rect 1855 2157 1861 2163
rect 3631 2157 3637 2163
rect 85 2077 91 2083
rect 1843 2077 1849 2083
rect 97 1997 103 2003
rect 1855 1997 1861 2003
rect 85 1917 91 1923
rect 1843 1917 1849 1923
rect 97 1837 103 1843
rect 1855 1837 1861 1843
rect 1855 1821 1861 1827
rect 3631 1821 3637 1827
rect 85 1753 91 1759
rect 1843 1753 1849 1759
rect 1843 1741 1849 1747
rect 3619 1741 3625 1747
rect 97 1673 103 1679
rect 1855 1673 1861 1679
rect 1855 1661 1861 1667
rect 3631 1661 3637 1667
rect 85 1597 91 1603
rect 1843 1597 1849 1603
rect 1843 1577 1849 1583
rect 3619 1577 3625 1583
rect 97 1517 103 1523
rect 1855 1517 1861 1523
rect 1855 1493 1861 1499
rect 3631 1493 3637 1499
rect 85 1433 91 1439
rect 1843 1433 1849 1439
rect 1843 1417 1849 1423
rect 3619 1417 3625 1423
rect 97 1357 103 1363
rect 1855 1357 1861 1363
rect 1855 1333 1861 1339
rect 3631 1333 3637 1339
rect 85 1277 91 1283
rect 1843 1277 1849 1283
rect 1843 1249 1849 1255
rect 3619 1249 3625 1255
rect 97 1201 103 1207
rect 1855 1201 1861 1207
rect 1855 1169 1861 1175
rect 3631 1169 3637 1175
rect 85 1121 91 1127
rect 1843 1121 1849 1127
rect 1843 1085 1849 1091
rect 3619 1085 3625 1091
rect 97 1037 103 1043
rect 1855 1037 1861 1043
rect 1855 1009 1861 1015
rect 3631 1009 3637 1015
rect 85 953 91 959
rect 1843 953 1849 959
rect 1843 925 1849 931
rect 3619 925 3625 931
rect 97 869 103 875
rect 1855 869 1861 875
rect 1855 837 1861 843
rect 3631 837 3637 843
rect 85 781 91 787
rect 1843 781 1849 787
rect 1843 753 1849 759
rect 3619 753 3625 759
rect 97 693 103 699
rect 1855 693 1861 699
rect 1855 673 1861 679
rect 3631 673 3637 679
rect 85 613 91 619
rect 1843 613 1849 619
rect 1843 593 1849 599
rect 3619 593 3625 599
rect 97 525 103 531
rect 1855 525 1861 531
rect 1855 517 1861 523
rect 3631 517 3637 523
rect 85 441 91 447
rect 1843 441 1849 447
rect 97 353 103 359
rect 1855 353 1861 359
rect 85 269 91 275
rect 1843 269 1849 275
rect 1855 181 1861 187
rect 3631 181 3637 187
rect 97 161 103 167
rect 1855 161 1861 167
rect 1843 105 1849 111
rect 3619 105 3625 111
rect 85 85 91 91
rect 1843 85 1849 91
<< m5 >>
rect 84 3567 92 3672
rect 84 3561 85 3567
rect 91 3561 92 3567
rect 84 3403 92 3561
rect 84 3397 85 3403
rect 91 3397 92 3403
rect 84 3247 92 3397
rect 84 3241 85 3247
rect 91 3241 92 3247
rect 84 3075 92 3241
rect 84 3069 85 3075
rect 91 3069 92 3075
rect 84 2911 92 3069
rect 84 2905 85 2911
rect 91 2905 92 2911
rect 84 2751 92 2905
rect 84 2745 85 2751
rect 91 2745 92 2751
rect 84 2587 92 2745
rect 84 2581 85 2587
rect 91 2581 92 2587
rect 84 2419 92 2581
rect 84 2413 85 2419
rect 91 2413 92 2419
rect 84 2259 92 2413
rect 84 2253 85 2259
rect 91 2253 92 2259
rect 84 2083 92 2253
rect 84 2077 85 2083
rect 91 2077 92 2083
rect 84 1923 92 2077
rect 84 1917 85 1923
rect 91 1917 92 1923
rect 84 1759 92 1917
rect 84 1753 85 1759
rect 91 1753 92 1759
rect 84 1603 92 1753
rect 84 1597 85 1603
rect 91 1597 92 1603
rect 84 1439 92 1597
rect 84 1433 85 1439
rect 91 1433 92 1439
rect 84 1283 92 1433
rect 84 1277 85 1283
rect 91 1277 92 1283
rect 84 1127 92 1277
rect 84 1121 85 1127
rect 91 1121 92 1127
rect 84 959 92 1121
rect 84 953 85 959
rect 91 953 92 959
rect 84 787 92 953
rect 84 781 85 787
rect 91 781 92 787
rect 84 619 92 781
rect 84 613 85 619
rect 91 613 92 619
rect 84 447 92 613
rect 84 441 85 447
rect 91 441 92 447
rect 84 275 92 441
rect 84 269 85 275
rect 91 269 92 275
rect 84 91 92 269
rect 84 85 85 91
rect 91 85 92 91
rect 84 72 92 85
rect 96 3643 104 3672
rect 96 3637 97 3643
rect 103 3637 104 3643
rect 96 3483 104 3637
rect 96 3477 97 3483
rect 103 3477 104 3483
rect 96 3323 104 3477
rect 96 3317 97 3323
rect 103 3317 104 3323
rect 96 3163 104 3317
rect 96 3157 97 3163
rect 103 3157 104 3163
rect 96 2987 104 3157
rect 96 2981 97 2987
rect 103 2981 104 2987
rect 96 2831 104 2981
rect 96 2825 97 2831
rect 103 2825 104 2831
rect 96 2667 104 2825
rect 96 2661 97 2667
rect 103 2661 104 2667
rect 96 2507 104 2661
rect 96 2501 97 2507
rect 103 2501 104 2507
rect 96 2335 104 2501
rect 96 2329 97 2335
rect 103 2329 104 2335
rect 96 2171 104 2329
rect 96 2165 97 2171
rect 103 2165 104 2171
rect 96 2003 104 2165
rect 96 1997 97 2003
rect 103 1997 104 2003
rect 96 1843 104 1997
rect 96 1837 97 1843
rect 103 1837 104 1843
rect 96 1679 104 1837
rect 96 1673 97 1679
rect 103 1673 104 1679
rect 96 1523 104 1673
rect 96 1517 97 1523
rect 103 1517 104 1523
rect 96 1363 104 1517
rect 96 1357 97 1363
rect 103 1357 104 1363
rect 96 1207 104 1357
rect 96 1201 97 1207
rect 103 1201 104 1207
rect 96 1043 104 1201
rect 96 1037 97 1043
rect 103 1037 104 1043
rect 96 875 104 1037
rect 96 869 97 875
rect 103 869 104 875
rect 96 699 104 869
rect 96 693 97 699
rect 103 693 104 699
rect 96 531 104 693
rect 96 525 97 531
rect 103 525 104 531
rect 96 359 104 525
rect 96 353 97 359
rect 103 353 104 359
rect 96 167 104 353
rect 96 161 97 167
rect 103 161 104 167
rect 96 72 104 161
rect 1842 3671 1850 3672
rect 1842 3665 1843 3671
rect 1849 3665 1850 3671
rect 1842 3567 1850 3665
rect 1842 3561 1843 3567
rect 1849 3561 1850 3567
rect 1842 3519 1850 3561
rect 1842 3513 1843 3519
rect 1849 3513 1850 3519
rect 1842 3403 1850 3513
rect 1842 3397 1843 3403
rect 1849 3397 1850 3403
rect 1842 3367 1850 3397
rect 1842 3361 1843 3367
rect 1849 3361 1850 3367
rect 1842 3247 1850 3361
rect 1842 3241 1843 3247
rect 1849 3241 1850 3247
rect 1842 3215 1850 3241
rect 1842 3209 1843 3215
rect 1849 3209 1850 3215
rect 1842 3075 1850 3209
rect 1842 3069 1843 3075
rect 1849 3069 1850 3075
rect 1842 3051 1850 3069
rect 1842 3045 1843 3051
rect 1849 3045 1850 3051
rect 1842 2911 1850 3045
rect 1842 2905 1843 2911
rect 1849 2905 1850 2911
rect 1842 2887 1850 2905
rect 1842 2881 1843 2887
rect 1849 2881 1850 2887
rect 1842 2751 1850 2881
rect 1842 2745 1843 2751
rect 1849 2745 1850 2751
rect 1842 2723 1850 2745
rect 1842 2717 1843 2723
rect 1849 2717 1850 2723
rect 1842 2587 1850 2717
rect 1842 2581 1843 2587
rect 1849 2581 1850 2587
rect 1842 2563 1850 2581
rect 1842 2557 1843 2563
rect 1849 2557 1850 2563
rect 1842 2419 1850 2557
rect 1842 2413 1843 2419
rect 1849 2413 1850 2419
rect 1842 2399 1850 2413
rect 1842 2393 1843 2399
rect 1849 2393 1850 2399
rect 1842 2259 1850 2393
rect 1842 2253 1843 2259
rect 1849 2253 1850 2259
rect 1842 2243 1850 2253
rect 1842 2237 1843 2243
rect 1849 2237 1850 2243
rect 1842 2083 1850 2237
rect 1842 2077 1843 2083
rect 1849 2077 1850 2083
rect 1842 1923 1850 2077
rect 1842 1917 1843 1923
rect 1849 1917 1850 1923
rect 1842 1759 1850 1917
rect 1842 1753 1843 1759
rect 1849 1753 1850 1759
rect 1842 1747 1850 1753
rect 1842 1741 1843 1747
rect 1849 1741 1850 1747
rect 1842 1603 1850 1741
rect 1842 1597 1843 1603
rect 1849 1597 1850 1603
rect 1842 1583 1850 1597
rect 1842 1577 1843 1583
rect 1849 1577 1850 1583
rect 1842 1439 1850 1577
rect 1842 1433 1843 1439
rect 1849 1433 1850 1439
rect 1842 1423 1850 1433
rect 1842 1417 1843 1423
rect 1849 1417 1850 1423
rect 1842 1283 1850 1417
rect 1842 1277 1843 1283
rect 1849 1277 1850 1283
rect 1842 1255 1850 1277
rect 1842 1249 1843 1255
rect 1849 1249 1850 1255
rect 1842 1127 1850 1249
rect 1842 1121 1843 1127
rect 1849 1121 1850 1127
rect 1842 1091 1850 1121
rect 1842 1085 1843 1091
rect 1849 1085 1850 1091
rect 1842 959 1850 1085
rect 1842 953 1843 959
rect 1849 953 1850 959
rect 1842 931 1850 953
rect 1842 925 1843 931
rect 1849 925 1850 931
rect 1842 787 1850 925
rect 1842 781 1843 787
rect 1849 781 1850 787
rect 1842 759 1850 781
rect 1842 753 1843 759
rect 1849 753 1850 759
rect 1842 619 1850 753
rect 1842 613 1843 619
rect 1849 613 1850 619
rect 1842 599 1850 613
rect 1842 593 1843 599
rect 1849 593 1850 599
rect 1842 447 1850 593
rect 1842 441 1843 447
rect 1849 441 1850 447
rect 1842 275 1850 441
rect 1842 269 1843 275
rect 1849 269 1850 275
rect 1842 111 1850 269
rect 1842 105 1843 111
rect 1849 105 1850 111
rect 1842 91 1850 105
rect 1842 85 1843 91
rect 1849 85 1850 91
rect 1842 72 1850 85
rect 1854 3643 1862 3672
rect 1854 3637 1855 3643
rect 1861 3637 1862 3643
rect 1854 3595 1862 3637
rect 1854 3589 1855 3595
rect 1861 3589 1862 3595
rect 1854 3483 1862 3589
rect 1854 3477 1855 3483
rect 1861 3477 1862 3483
rect 1854 3443 1862 3477
rect 1854 3437 1855 3443
rect 1861 3437 1862 3443
rect 1854 3323 1862 3437
rect 1854 3317 1855 3323
rect 1861 3317 1862 3323
rect 1854 3291 1862 3317
rect 1854 3285 1855 3291
rect 1861 3285 1862 3291
rect 1854 3163 1862 3285
rect 1854 3157 1855 3163
rect 1861 3157 1862 3163
rect 1854 3139 1862 3157
rect 1854 3133 1855 3139
rect 1861 3133 1862 3139
rect 1854 2987 1862 3133
rect 1854 2981 1855 2987
rect 1861 2981 1862 2987
rect 1854 2963 1862 2981
rect 1854 2957 1855 2963
rect 1861 2957 1862 2963
rect 1854 2831 1862 2957
rect 1854 2825 1855 2831
rect 1861 2825 1862 2831
rect 1854 2799 1862 2825
rect 1854 2793 1855 2799
rect 1861 2793 1862 2799
rect 1854 2667 1862 2793
rect 1854 2661 1855 2667
rect 1861 2661 1862 2667
rect 1854 2639 1862 2661
rect 1854 2633 1855 2639
rect 1861 2633 1862 2639
rect 1854 2507 1862 2633
rect 1854 2501 1855 2507
rect 1861 2501 1862 2507
rect 1854 2479 1862 2501
rect 1854 2473 1855 2479
rect 1861 2473 1862 2479
rect 1854 2335 1862 2473
rect 1854 2329 1855 2335
rect 1861 2329 1862 2335
rect 1854 2319 1862 2329
rect 1854 2313 1855 2319
rect 1861 2313 1862 2319
rect 1854 2171 1862 2313
rect 1854 2165 1855 2171
rect 1861 2165 1862 2171
rect 1854 2163 1862 2165
rect 1854 2157 1855 2163
rect 1861 2157 1862 2163
rect 1854 2003 1862 2157
rect 1854 1997 1855 2003
rect 1861 1997 1862 2003
rect 1854 1843 1862 1997
rect 1854 1837 1855 1843
rect 1861 1837 1862 1843
rect 1854 1827 1862 1837
rect 1854 1821 1855 1827
rect 1861 1821 1862 1827
rect 1854 1679 1862 1821
rect 1854 1673 1855 1679
rect 1861 1673 1862 1679
rect 1854 1667 1862 1673
rect 1854 1661 1855 1667
rect 1861 1661 1862 1667
rect 1854 1523 1862 1661
rect 1854 1517 1855 1523
rect 1861 1517 1862 1523
rect 1854 1499 1862 1517
rect 1854 1493 1855 1499
rect 1861 1493 1862 1499
rect 1854 1363 1862 1493
rect 1854 1357 1855 1363
rect 1861 1357 1862 1363
rect 1854 1339 1862 1357
rect 1854 1333 1855 1339
rect 1861 1333 1862 1339
rect 1854 1207 1862 1333
rect 1854 1201 1855 1207
rect 1861 1201 1862 1207
rect 1854 1175 1862 1201
rect 1854 1169 1855 1175
rect 1861 1169 1862 1175
rect 1854 1043 1862 1169
rect 1854 1037 1855 1043
rect 1861 1037 1862 1043
rect 1854 1015 1862 1037
rect 1854 1009 1855 1015
rect 1861 1009 1862 1015
rect 1854 875 1862 1009
rect 1854 869 1855 875
rect 1861 869 1862 875
rect 1854 843 1862 869
rect 1854 837 1855 843
rect 1861 837 1862 843
rect 1854 699 1862 837
rect 1854 693 1855 699
rect 1861 693 1862 699
rect 1854 679 1862 693
rect 1854 673 1855 679
rect 1861 673 1862 679
rect 1854 531 1862 673
rect 1854 525 1855 531
rect 1861 525 1862 531
rect 1854 523 1862 525
rect 1854 517 1855 523
rect 1861 517 1862 523
rect 1854 359 1862 517
rect 1854 353 1855 359
rect 1861 353 1862 359
rect 1854 187 1862 353
rect 1854 181 1855 187
rect 1861 181 1862 187
rect 1854 167 1862 181
rect 1854 161 1855 167
rect 1861 161 1862 167
rect 1854 72 1862 161
rect 3618 3671 3626 3672
rect 3618 3665 3619 3671
rect 3625 3665 3626 3671
rect 3618 3519 3626 3665
rect 3618 3513 3619 3519
rect 3625 3513 3626 3519
rect 3618 3367 3626 3513
rect 3618 3361 3619 3367
rect 3625 3361 3626 3367
rect 3618 3215 3626 3361
rect 3618 3209 3619 3215
rect 3625 3209 3626 3215
rect 3618 3051 3626 3209
rect 3618 3045 3619 3051
rect 3625 3045 3626 3051
rect 3618 2887 3626 3045
rect 3618 2881 3619 2887
rect 3625 2881 3626 2887
rect 3618 2723 3626 2881
rect 3618 2717 3619 2723
rect 3625 2717 3626 2723
rect 3618 2563 3626 2717
rect 3618 2557 3619 2563
rect 3625 2557 3626 2563
rect 3618 2399 3626 2557
rect 3618 2393 3619 2399
rect 3625 2393 3626 2399
rect 3618 2243 3626 2393
rect 3618 2237 3619 2243
rect 3625 2237 3626 2243
rect 3618 1747 3626 2237
rect 3618 1741 3619 1747
rect 3625 1741 3626 1747
rect 3618 1583 3626 1741
rect 3618 1577 3619 1583
rect 3625 1577 3626 1583
rect 3618 1423 3626 1577
rect 3618 1417 3619 1423
rect 3625 1417 3626 1423
rect 3618 1255 3626 1417
rect 3618 1249 3619 1255
rect 3625 1249 3626 1255
rect 3618 1091 3626 1249
rect 3618 1085 3619 1091
rect 3625 1085 3626 1091
rect 3618 931 3626 1085
rect 3618 925 3619 931
rect 3625 925 3626 931
rect 3618 759 3626 925
rect 3618 753 3619 759
rect 3625 753 3626 759
rect 3618 599 3626 753
rect 3618 593 3619 599
rect 3625 593 3626 599
rect 3618 111 3626 593
rect 3618 105 3619 111
rect 3625 105 3626 111
rect 3618 72 3626 105
rect 3630 3595 3638 3672
rect 3630 3589 3631 3595
rect 3637 3589 3638 3595
rect 3630 3443 3638 3589
rect 3630 3437 3631 3443
rect 3637 3437 3638 3443
rect 3630 3291 3638 3437
rect 3630 3285 3631 3291
rect 3637 3285 3638 3291
rect 3630 3139 3638 3285
rect 3630 3133 3631 3139
rect 3637 3133 3638 3139
rect 3630 2963 3638 3133
rect 3630 2957 3631 2963
rect 3637 2957 3638 2963
rect 3630 2799 3638 2957
rect 3630 2793 3631 2799
rect 3637 2793 3638 2799
rect 3630 2639 3638 2793
rect 3630 2633 3631 2639
rect 3637 2633 3638 2639
rect 3630 2479 3638 2633
rect 3630 2473 3631 2479
rect 3637 2473 3638 2479
rect 3630 2319 3638 2473
rect 3630 2313 3631 2319
rect 3637 2313 3638 2319
rect 3630 2163 3638 2313
rect 3630 2157 3631 2163
rect 3637 2157 3638 2163
rect 3630 1827 3638 2157
rect 3630 1821 3631 1827
rect 3637 1821 3638 1827
rect 3630 1667 3638 1821
rect 3630 1661 3631 1667
rect 3637 1661 3638 1667
rect 3630 1499 3638 1661
rect 3630 1493 3631 1499
rect 3637 1493 3638 1499
rect 3630 1339 3638 1493
rect 3630 1333 3631 1339
rect 3637 1333 3638 1339
rect 3630 1175 3638 1333
rect 3630 1169 3631 1175
rect 3637 1169 3638 1175
rect 3630 1015 3638 1169
rect 3630 1009 3631 1015
rect 3637 1009 3638 1015
rect 3630 843 3638 1009
rect 3630 837 3631 843
rect 3637 837 3638 843
rect 3630 679 3638 837
rect 3630 673 3631 679
rect 3637 673 3638 679
rect 3630 523 3638 673
rect 3630 517 3631 523
rect 3637 517 3638 523
rect 3630 187 3638 517
rect 3630 181 3631 187
rect 3637 181 3638 187
rect 3630 72 3638 181
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__173
timestamp 1731220559
transform 1 0 3584 0 -1 3648
box 7 3 12 24
use welltap_svt  __well_tap__172
timestamp 1731220559
transform 1 0 1864 0 -1 3648
box 7 3 12 24
use welltap_svt  __well_tap__171
timestamp 1731220559
transform 1 0 3584 0 1 3536
box 7 3 12 24
use welltap_svt  __well_tap__170
timestamp 1731220559
transform 1 0 1864 0 1 3536
box 7 3 12 24
use welltap_svt  __well_tap__169
timestamp 1731220559
transform 1 0 3584 0 -1 3496
box 7 3 12 24
use welltap_svt  __well_tap__168
timestamp 1731220559
transform 1 0 1864 0 -1 3496
box 7 3 12 24
use welltap_svt  __well_tap__167
timestamp 1731220559
transform 1 0 3584 0 1 3384
box 7 3 12 24
use welltap_svt  __well_tap__166
timestamp 1731220559
transform 1 0 1864 0 1 3384
box 7 3 12 24
use welltap_svt  __well_tap__165
timestamp 1731220559
transform 1 0 3584 0 -1 3344
box 7 3 12 24
use welltap_svt  __well_tap__164
timestamp 1731220559
transform 1 0 1864 0 -1 3344
box 7 3 12 24
use welltap_svt  __well_tap__163
timestamp 1731220559
transform 1 0 3584 0 1 3232
box 7 3 12 24
use welltap_svt  __well_tap__162
timestamp 1731220559
transform 1 0 1864 0 1 3232
box 7 3 12 24
use welltap_svt  __well_tap__161
timestamp 1731220559
transform 1 0 3584 0 -1 3192
box 7 3 12 24
use welltap_svt  __well_tap__160
timestamp 1731220559
transform 1 0 1864 0 -1 3192
box 7 3 12 24
use welltap_svt  __well_tap__159
timestamp 1731220559
transform 1 0 3584 0 1 3080
box 7 3 12 24
use welltap_svt  __well_tap__158
timestamp 1731220559
transform 1 0 1864 0 1 3080
box 7 3 12 24
use welltap_svt  __well_tap__157
timestamp 1731220559
transform 1 0 3584 0 -1 3028
box 7 3 12 24
use welltap_svt  __well_tap__156
timestamp 1731220559
transform 1 0 1864 0 -1 3028
box 7 3 12 24
use welltap_svt  __well_tap__155
timestamp 1731220559
transform 1 0 3584 0 1 2904
box 7 3 12 24
use welltap_svt  __well_tap__154
timestamp 1731220559
transform 1 0 1864 0 1 2904
box 7 3 12 24
use welltap_svt  __well_tap__153
timestamp 1731220559
transform 1 0 3584 0 -1 2864
box 7 3 12 24
use welltap_svt  __well_tap__152
timestamp 1731220559
transform 1 0 1864 0 -1 2864
box 7 3 12 24
use welltap_svt  __well_tap__151
timestamp 1731220559
transform 1 0 3584 0 1 2740
box 7 3 12 24
use welltap_svt  __well_tap__150
timestamp 1731220559
transform 1 0 1864 0 1 2740
box 7 3 12 24
use welltap_svt  __well_tap__149
timestamp 1731220559
transform 1 0 3584 0 -1 2700
box 7 3 12 24
use welltap_svt  __well_tap__148
timestamp 1731220559
transform 1 0 1864 0 -1 2700
box 7 3 12 24
use welltap_svt  __well_tap__147
timestamp 1731220559
transform 1 0 3584 0 1 2580
box 7 3 12 24
use welltap_svt  __well_tap__146
timestamp 1731220559
transform 1 0 1864 0 1 2580
box 7 3 12 24
use welltap_svt  __well_tap__145
timestamp 1731220559
transform 1 0 3584 0 -1 2540
box 7 3 12 24
use welltap_svt  __well_tap__144
timestamp 1731220559
transform 1 0 1864 0 -1 2540
box 7 3 12 24
use welltap_svt  __well_tap__143
timestamp 1731220559
transform 1 0 3584 0 1 2420
box 7 3 12 24
use welltap_svt  __well_tap__142
timestamp 1731220559
transform 1 0 1864 0 1 2420
box 7 3 12 24
use welltap_svt  __well_tap__141
timestamp 1731220559
transform 1 0 3584 0 -1 2376
box 7 3 12 24
use welltap_svt  __well_tap__140
timestamp 1731220559
transform 1 0 1864 0 -1 2376
box 7 3 12 24
use welltap_svt  __well_tap__139
timestamp 1731220559
transform 1 0 3584 0 1 2260
box 7 3 12 24
use welltap_svt  __well_tap__138
timestamp 1731220559
transform 1 0 1864 0 1 2260
box 7 3 12 24
use welltap_svt  __well_tap__137
timestamp 1731220559
transform 1 0 3584 0 -1 2220
box 7 3 12 24
use welltap_svt  __well_tap__136
timestamp 1731220559
transform 1 0 1864 0 -1 2220
box 7 3 12 24
use welltap_svt  __well_tap__135
timestamp 1731220559
transform 1 0 3584 0 1 2104
box 7 3 12 24
use welltap_svt  __well_tap__134
timestamp 1731220559
transform 1 0 1864 0 1 2104
box 7 3 12 24
use welltap_svt  __well_tap__133
timestamp 1731220559
transform 1 0 3584 0 -1 2056
box 7 3 12 24
use welltap_svt  __well_tap__132
timestamp 1731220559
transform 1 0 1864 0 -1 2056
box 7 3 12 24
use welltap_svt  __well_tap__131
timestamp 1731220559
transform 1 0 3584 0 1 1944
box 7 3 12 24
use welltap_svt  __well_tap__130
timestamp 1731220559
transform 1 0 1864 0 1 1944
box 7 3 12 24
use welltap_svt  __well_tap__129
timestamp 1731220559
transform 1 0 3584 0 -1 1896
box 7 3 12 24
use welltap_svt  __well_tap__128
timestamp 1731220559
transform 1 0 1864 0 -1 1896
box 7 3 12 24
use welltap_svt  __well_tap__127
timestamp 1731220559
transform 1 0 3584 0 1 1768
box 7 3 12 24
use welltap_svt  __well_tap__126
timestamp 1731220559
transform 1 0 1864 0 1 1768
box 7 3 12 24
use welltap_svt  __well_tap__125
timestamp 1731220559
transform 1 0 3584 0 -1 1724
box 7 3 12 24
use welltap_svt  __well_tap__124
timestamp 1731220559
transform 1 0 1864 0 -1 1724
box 7 3 12 24
use welltap_svt  __well_tap__123
timestamp 1731220559
transform 1 0 3584 0 1 1608
box 7 3 12 24
use welltap_svt  __well_tap__122
timestamp 1731220559
transform 1 0 1864 0 1 1608
box 7 3 12 24
use welltap_svt  __well_tap__121
timestamp 1731220559
transform 1 0 3584 0 -1 1560
box 7 3 12 24
use welltap_svt  __well_tap__120
timestamp 1731220559
transform 1 0 1864 0 -1 1560
box 7 3 12 24
use welltap_svt  __well_tap__119
timestamp 1731220559
transform 1 0 3584 0 1 1440
box 7 3 12 24
use welltap_svt  __well_tap__118
timestamp 1731220559
transform 1 0 1864 0 1 1440
box 7 3 12 24
use welltap_svt  __well_tap__117
timestamp 1731220559
transform 1 0 3584 0 -1 1400
box 7 3 12 24
use welltap_svt  __well_tap__116
timestamp 1731220559
transform 1 0 1864 0 -1 1400
box 7 3 12 24
use welltap_svt  __well_tap__115
timestamp 1731220559
transform 1 0 3584 0 1 1280
box 7 3 12 24
use welltap_svt  __well_tap__114
timestamp 1731220559
transform 1 0 1864 0 1 1280
box 7 3 12 24
use welltap_svt  __well_tap__113
timestamp 1731220559
transform 1 0 3584 0 -1 1232
box 7 3 12 24
use welltap_svt  __well_tap__112
timestamp 1731220559
transform 1 0 1864 0 -1 1232
box 7 3 12 24
use welltap_svt  __well_tap__111
timestamp 1731220559
transform 1 0 3584 0 1 1116
box 7 3 12 24
use welltap_svt  __well_tap__110
timestamp 1731220559
transform 1 0 1864 0 1 1116
box 7 3 12 24
use welltap_svt  __well_tap__109
timestamp 1731220559
transform 1 0 3584 0 -1 1068
box 7 3 12 24
use welltap_svt  __well_tap__108
timestamp 1731220559
transform 1 0 1864 0 -1 1068
box 7 3 12 24
use welltap_svt  __well_tap__107
timestamp 1731220559
transform 1 0 3584 0 1 956
box 7 3 12 24
use welltap_svt  __well_tap__106
timestamp 1731220559
transform 1 0 1864 0 1 956
box 7 3 12 24
use welltap_svt  __well_tap__105
timestamp 1731220559
transform 1 0 3584 0 -1 908
box 7 3 12 24
use welltap_svt  __well_tap__104
timestamp 1731220559
transform 1 0 1864 0 -1 908
box 7 3 12 24
use welltap_svt  __well_tap__103
timestamp 1731220559
transform 1 0 3584 0 1 784
box 7 3 12 24
use welltap_svt  __well_tap__102
timestamp 1731220559
transform 1 0 1864 0 1 784
box 7 3 12 24
use welltap_svt  __well_tap__101
timestamp 1731220559
transform 1 0 3584 0 -1 736
box 7 3 12 24
use welltap_svt  __well_tap__100
timestamp 1731220559
transform 1 0 1864 0 -1 736
box 7 3 12 24
use welltap_svt  __well_tap__99
timestamp 1731220559
transform 1 0 3584 0 1 620
box 7 3 12 24
use welltap_svt  __well_tap__98
timestamp 1731220559
transform 1 0 1864 0 1 620
box 7 3 12 24
use welltap_svt  __well_tap__97
timestamp 1731220559
transform 1 0 3584 0 -1 576
box 7 3 12 24
use welltap_svt  __well_tap__96
timestamp 1731220559
transform 1 0 1864 0 -1 576
box 7 3 12 24
use welltap_svt  __well_tap__95
timestamp 1731220559
transform 1 0 3584 0 1 464
box 7 3 12 24
use welltap_svt  __well_tap__94
timestamp 1731220559
transform 1 0 1864 0 1 464
box 7 3 12 24
use welltap_svt  __well_tap__93
timestamp 1731220559
transform 1 0 3584 0 -1 420
box 7 3 12 24
use welltap_svt  __well_tap__92
timestamp 1731220559
transform 1 0 1864 0 -1 420
box 7 3 12 24
use welltap_svt  __well_tap__91
timestamp 1731220559
transform 1 0 3584 0 1 300
box 7 3 12 24
use welltap_svt  __well_tap__90
timestamp 1731220559
transform 1 0 1864 0 1 300
box 7 3 12 24
use welltap_svt  __well_tap__89
timestamp 1731220559
transform 1 0 3584 0 -1 252
box 7 3 12 24
use welltap_svt  __well_tap__88
timestamp 1731220559
transform 1 0 1864 0 -1 252
box 7 3 12 24
use welltap_svt  __well_tap__87
timestamp 1731220559
transform 1 0 3584 0 1 128
box 7 3 12 24
use welltap_svt  __well_tap__86
timestamp 1731220559
transform 1 0 1864 0 1 128
box 7 3 12 24
use welltap_svt  __well_tap__85
timestamp 1731220559
transform 1 0 1824 0 1 3584
box 7 3 12 24
use welltap_svt  __well_tap__84
timestamp 1731220559
transform 1 0 104 0 1 3584
box 7 3 12 24
use welltap_svt  __well_tap__83
timestamp 1731220559
transform 1 0 1824 0 -1 3544
box 7 3 12 24
use welltap_svt  __well_tap__82
timestamp 1731220559
transform 1 0 104 0 -1 3544
box 7 3 12 24
use welltap_svt  __well_tap__81
timestamp 1731220559
transform 1 0 1824 0 1 3424
box 7 3 12 24
use welltap_svt  __well_tap__80
timestamp 1731220559
transform 1 0 104 0 1 3424
box 7 3 12 24
use welltap_svt  __well_tap__79
timestamp 1731220559
transform 1 0 1824 0 -1 3380
box 7 3 12 24
use welltap_svt  __well_tap__78
timestamp 1731220559
transform 1 0 104 0 -1 3380
box 7 3 12 24
use welltap_svt  __well_tap__77
timestamp 1731220559
transform 1 0 1824 0 1 3264
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220559
transform 1 0 104 0 1 3264
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220559
transform 1 0 1824 0 -1 3224
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220559
transform 1 0 104 0 -1 3224
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220559
transform 1 0 1824 0 1 3104
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220559
transform 1 0 104 0 1 3104
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220559
transform 1 0 1824 0 -1 3052
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220559
transform 1 0 104 0 -1 3052
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220559
transform 1 0 1824 0 1 2928
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220559
transform 1 0 104 0 1 2928
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220559
transform 1 0 1824 0 -1 2888
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220559
transform 1 0 104 0 -1 2888
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220559
transform 1 0 1824 0 1 2772
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220559
transform 1 0 104 0 1 2772
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220559
transform 1 0 1824 0 -1 2728
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220559
transform 1 0 104 0 -1 2728
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220559
transform 1 0 1824 0 1 2608
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220559
transform 1 0 104 0 1 2608
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220559
transform 1 0 1824 0 -1 2564
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220559
transform 1 0 104 0 -1 2564
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220559
transform 1 0 1824 0 1 2448
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220559
transform 1 0 104 0 1 2448
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220559
transform 1 0 1824 0 -1 2396
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220559
transform 1 0 104 0 -1 2396
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220559
transform 1 0 1824 0 1 2276
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220559
transform 1 0 104 0 1 2276
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220559
transform 1 0 1824 0 -1 2236
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220559
transform 1 0 104 0 -1 2236
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220559
transform 1 0 1824 0 1 2112
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220559
transform 1 0 104 0 1 2112
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220559
transform 1 0 1824 0 -1 2060
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220559
transform 1 0 104 0 -1 2060
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220559
transform 1 0 1824 0 1 1944
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220559
transform 1 0 104 0 1 1944
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220559
transform 1 0 1824 0 -1 1900
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220559
transform 1 0 104 0 -1 1900
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220559
transform 1 0 1824 0 1 1784
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220559
transform 1 0 104 0 1 1784
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220559
transform 1 0 1824 0 -1 1736
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220559
transform 1 0 104 0 -1 1736
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220559
transform 1 0 1824 0 1 1620
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220559
transform 1 0 104 0 1 1620
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220559
transform 1 0 1824 0 -1 1580
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220559
transform 1 0 104 0 -1 1580
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220559
transform 1 0 1824 0 1 1464
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220559
transform 1 0 104 0 1 1464
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220559
transform 1 0 1824 0 -1 1416
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220559
transform 1 0 104 0 -1 1416
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220559
transform 1 0 1824 0 1 1304
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220559
transform 1 0 104 0 1 1304
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220559
transform 1 0 1824 0 -1 1260
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220559
transform 1 0 104 0 -1 1260
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220559
transform 1 0 1824 0 1 1148
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220559
transform 1 0 104 0 1 1148
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220559
transform 1 0 1824 0 -1 1104
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220559
transform 1 0 104 0 -1 1104
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220559
transform 1 0 1824 0 1 984
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220559
transform 1 0 104 0 1 984
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220559
transform 1 0 1824 0 -1 936
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220559
transform 1 0 104 0 -1 936
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220559
transform 1 0 1824 0 1 816
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220559
transform 1 0 104 0 1 816
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220559
transform 1 0 1824 0 -1 764
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220559
transform 1 0 104 0 -1 764
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220559
transform 1 0 1824 0 1 640
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220559
transform 1 0 104 0 1 640
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220559
transform 1 0 1824 0 -1 596
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220559
transform 1 0 104 0 -1 596
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220559
transform 1 0 1824 0 1 472
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220559
transform 1 0 104 0 1 472
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220559
transform 1 0 1824 0 -1 424
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220559
transform 1 0 104 0 -1 424
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220559
transform 1 0 1824 0 1 300
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220559
transform 1 0 104 0 1 300
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220559
transform 1 0 1824 0 -1 252
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220559
transform 1 0 104 0 -1 252
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220559
transform 1 0 1824 0 1 108
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220559
transform 1 0 104 0 1 108
box 7 3 12 24
use _0_0std_0_0cells_0_0LATCHINV  tst_5999_6
timestamp 1731220559
transform 1 0 3496 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5998_6
timestamp 1731220559
transform 1 0 3496 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5997_6
timestamp 1731220559
transform 1 0 3392 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5996_6
timestamp 1731220559
transform 1 0 3496 0 -1 440
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5995_6
timestamp 1731220559
transform 1 0 3496 0 1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5994_6
timestamp 1731220559
transform 1 0 3496 0 -1 596
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5993_6
timestamp 1731220559
transform 1 0 3496 0 1 600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5992_6
timestamp 1731220559
transform 1 0 3496 0 -1 756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5991_6
timestamp 1731220559
transform 1 0 3496 0 1 764
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5990_6
timestamp 1731220559
transform 1 0 3416 0 -1 928
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5989_6
timestamp 1731220559
transform 1 0 3496 0 -1 928
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5988_6
timestamp 1731220559
transform 1 0 3496 0 1 936
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5987_6
timestamp 1731220559
transform 1 0 3496 0 -1 1088
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5986_6
timestamp 1731220559
transform 1 0 3496 0 1 1096
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5985_6
timestamp 1731220559
transform 1 0 3496 0 -1 1252
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5984_6
timestamp 1731220559
transform 1 0 3352 0 -1 1252
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5983_6
timestamp 1731220559
transform 1 0 3184 0 -1 1252
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5982_6
timestamp 1731220559
transform 1 0 3384 0 1 1096
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5981_6
timestamp 1731220559
transform 1 0 3248 0 1 1096
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5980_6
timestamp 1731220559
transform 1 0 3112 0 1 1096
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5979_6
timestamp 1731220559
transform 1 0 2968 0 1 1096
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5978_6
timestamp 1731220559
transform 1 0 3040 0 -1 1088
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5977_6
timestamp 1731220559
transform 1 0 3200 0 -1 1088
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5976_6
timestamp 1731220559
transform 1 0 3360 0 -1 1088
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5975_6
timestamp 1731220559
transform 1 0 3352 0 1 936
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5974_6
timestamp 1731220559
transform 1 0 3192 0 1 936
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5973_6
timestamp 1731220559
transform 1 0 3040 0 1 936
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5972_6
timestamp 1731220559
transform 1 0 3008 0 -1 928
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5971_6
timestamp 1731220559
transform 1 0 3104 0 -1 928
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5970_6
timestamp 1731220559
transform 1 0 3208 0 -1 928
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5969_6
timestamp 1731220559
transform 1 0 3312 0 -1 928
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5968_6
timestamp 1731220559
transform 1 0 3392 0 1 764
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5967_6
timestamp 1731220559
transform 1 0 3264 0 1 764
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5966_6
timestamp 1731220559
transform 1 0 3144 0 1 764
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5965_6
timestamp 1731220559
transform 1 0 3024 0 1 764
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5964_6
timestamp 1731220559
transform 1 0 3040 0 -1 756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5963_6
timestamp 1731220559
transform 1 0 3192 0 -1 756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5962_6
timestamp 1731220559
transform 1 0 3352 0 -1 756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5961_6
timestamp 1731220559
transform 1 0 3344 0 1 600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5960_6
timestamp 1731220559
transform 1 0 3168 0 1 600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5959_6
timestamp 1731220559
transform 1 0 2992 0 1 600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5958_6
timestamp 1731220559
transform 1 0 2816 0 1 600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5957_6
timestamp 1731220559
transform 1 0 2968 0 -1 596
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5956_6
timestamp 1731220559
transform 1 0 3144 0 -1 596
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5955_6
timestamp 1731220559
transform 1 0 3328 0 -1 596
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5954_6
timestamp 1731220559
transform 1 0 3336 0 1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5953_6
timestamp 1731220559
transform 1 0 3160 0 1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5952_6
timestamp 1731220559
transform 1 0 3208 0 -1 440
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5951_6
timestamp 1731220559
transform 1 0 3360 0 -1 440
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5950_6
timestamp 1731220559
transform 1 0 3272 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5949_6
timestamp 1731220559
transform 1 0 3152 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5948_6
timestamp 1731220559
transform 1 0 3024 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5947_6
timestamp 1731220559
transform 1 0 3072 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5946_6
timestamp 1731220559
transform 1 0 3216 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5945_6
timestamp 1731220559
transform 1 0 3368 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5944_6
timestamp 1731220559
transform 1 0 3384 0 1 108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5943_6
timestamp 1731220559
transform 1 0 3288 0 1 108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5942_6
timestamp 1731220559
transform 1 0 3192 0 1 108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5941_6
timestamp 1731220559
transform 1 0 3096 0 1 108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5940_6
timestamp 1731220559
transform 1 0 3000 0 1 108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5939_6
timestamp 1731220559
transform 1 0 2904 0 1 108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5938_6
timestamp 1731220559
transform 1 0 2800 0 1 108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5937_6
timestamp 1731220559
transform 1 0 2688 0 1 108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5936_6
timestamp 1731220559
transform 1 0 2568 0 1 108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5935_6
timestamp 1731220559
transform 1 0 2640 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5934_6
timestamp 1731220559
transform 1 0 2784 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5933_6
timestamp 1731220559
transform 1 0 2928 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5932_6
timestamp 1731220559
transform 1 0 2896 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5931_6
timestamp 1731220559
transform 1 0 2760 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5930_6
timestamp 1731220559
transform 1 0 2792 0 -1 440
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5929_6
timestamp 1731220559
transform 1 0 2920 0 -1 440
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5928_6
timestamp 1731220559
transform 1 0 3064 0 -1 440
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5927_6
timestamp 1731220559
transform 1 0 2984 0 1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5926_6
timestamp 1731220559
transform 1 0 2824 0 1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5925_6
timestamp 1731220559
transform 1 0 2800 0 -1 596
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5924_6
timestamp 1731220559
transform 1 0 2640 0 -1 596
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5923_6
timestamp 1731220559
transform 1 0 2640 0 1 600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5922_6
timestamp 1731220559
transform 1 0 2464 0 1 600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5921_6
timestamp 1731220559
transform 1 0 2584 0 -1 756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5920_6
timestamp 1731220559
transform 1 0 2736 0 -1 756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5919_6
timestamp 1731220559
transform 1 0 2888 0 -1 756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5918_6
timestamp 1731220559
transform 1 0 2768 0 1 764
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5917_6
timestamp 1731220559
transform 1 0 2896 0 1 764
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5916_6
timestamp 1731220559
transform 1 0 2904 0 -1 928
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5915_6
timestamp 1731220559
transform 1 0 2800 0 -1 928
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5914_6
timestamp 1731220559
transform 1 0 2896 0 1 936
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5913_6
timestamp 1731220559
transform 1 0 2768 0 1 936
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5912_6
timestamp 1731220559
transform 1 0 2744 0 -1 1088
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5911_6
timestamp 1731220559
transform 1 0 2888 0 -1 1088
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5910_6
timestamp 1731220559
transform 1 0 2824 0 1 1096
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5909_6
timestamp 1731220559
transform 1 0 2672 0 1 1096
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5908_6
timestamp 1731220559
transform 1 0 2656 0 -1 1252
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5907_6
timestamp 1731220559
transform 1 0 2464 0 -1 1252
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5906_6
timestamp 1731220559
transform 1 0 2840 0 -1 1252
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5905_6
timestamp 1731220559
transform 1 0 3016 0 -1 1252
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5904_6
timestamp 1731220559
transform 1 0 3168 0 1 1260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5903_6
timestamp 1731220559
transform 1 0 3048 0 1 1260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5902_6
timestamp 1731220559
transform 1 0 2936 0 1 1260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5901_6
timestamp 1731220559
transform 1 0 2824 0 1 1260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5900_6
timestamp 1731220559
transform 1 0 2704 0 1 1260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5899_6
timestamp 1731220559
transform 1 0 2576 0 1 1260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5898_6
timestamp 1731220559
transform 1 0 2904 0 -1 1420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5897_6
timestamp 1731220559
transform 1 0 2784 0 -1 1420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5896_6
timestamp 1731220559
transform 1 0 2664 0 -1 1420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5895_6
timestamp 1731220559
transform 1 0 2544 0 -1 1420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5894_6
timestamp 1731220559
transform 1 0 2424 0 -1 1420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5893_6
timestamp 1731220559
transform 1 0 2552 0 1 1420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5892_6
timestamp 1731220559
transform 1 0 2704 0 1 1420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5891_6
timestamp 1731220559
transform 1 0 2864 0 1 1420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5890_6
timestamp 1731220559
transform 1 0 3024 0 1 1420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5889_6
timestamp 1731220559
transform 1 0 2976 0 -1 1580
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5888_6
timestamp 1731220559
transform 1 0 2832 0 -1 1580
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5887_6
timestamp 1731220559
transform 1 0 2680 0 -1 1580
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5886_6
timestamp 1731220559
transform 1 0 2768 0 1 1588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5885_6
timestamp 1731220559
transform 1 0 2912 0 1 1588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5884_6
timestamp 1731220559
transform 1 0 3056 0 1 1588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5883_6
timestamp 1731220559
transform 1 0 3040 0 -1 1744
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5882_6
timestamp 1731220559
transform 1 0 2920 0 -1 1744
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5881_6
timestamp 1731220559
transform 1 0 2792 0 -1 1744
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5880_6
timestamp 1731220559
transform 1 0 2864 0 1 1748
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5879_6
timestamp 1731220559
transform 1 0 3016 0 1 1748
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5878_6
timestamp 1731220559
transform 1 0 3152 0 -1 1744
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5877_6
timestamp 1731220559
transform 1 0 3264 0 -1 1744
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5876_6
timestamp 1731220559
transform 1 0 3360 0 1 1588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5875_6
timestamp 1731220559
transform 1 0 3208 0 1 1588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5874_6
timestamp 1731220559
transform 1 0 3112 0 -1 1580
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5873_6
timestamp 1731220559
transform 1 0 3248 0 -1 1580
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5872_6
timestamp 1731220559
transform 1 0 3384 0 -1 1580
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5871_6
timestamp 1731220559
transform 1 0 3352 0 1 1420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5870_6
timestamp 1731220559
transform 1 0 3184 0 1 1420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5869_6
timestamp 1731220559
transform 1 0 3496 0 1 1420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5868_6
timestamp 1731220559
transform 1 0 3496 0 -1 1580
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5867_6
timestamp 1731220559
transform 1 0 3496 0 1 1588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5866_6
timestamp 1731220559
transform 1 0 3496 0 -1 1744
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5865_6
timestamp 1731220559
transform 1 0 3384 0 -1 1744
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5864_6
timestamp 1731220559
transform 1 0 3456 0 1 1748
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5863_6
timestamp 1731220559
transform 1 0 3304 0 1 1748
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5862_6
timestamp 1731220559
transform 1 0 3160 0 1 1748
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5861_6
timestamp 1731220559
transform 1 0 3240 0 -1 1916
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5860_6
timestamp 1731220559
transform 1 0 3112 0 -1 1916
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5859_6
timestamp 1731220559
transform 1 0 2984 0 -1 1916
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5858_6
timestamp 1731220559
transform 1 0 2864 0 -1 1916
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5857_6
timestamp 1731220559
transform 1 0 2752 0 -1 1916
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5856_6
timestamp 1731220559
transform 1 0 2656 0 -1 1916
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5855_6
timestamp 1731220559
transform 1 0 2568 0 -1 1916
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5854_6
timestamp 1731220559
transform 1 0 2480 0 -1 1916
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5853_6
timestamp 1731220559
transform 1 0 2392 0 -1 1916
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5852_6
timestamp 1731220559
transform 1 0 2312 0 -1 1916
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5851_6
timestamp 1731220559
transform 1 0 2432 0 1 1924
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5850_6
timestamp 1731220559
transform 1 0 2568 0 1 1924
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5849_6
timestamp 1731220559
transform 1 0 2728 0 1 1924
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5848_6
timestamp 1731220559
transform 1 0 2904 0 1 1924
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5847_6
timestamp 1731220559
transform 1 0 3312 0 1 1924
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5846_6
timestamp 1731220559
transform 1 0 3104 0 1 1924
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5845_6
timestamp 1731220559
transform 1 0 2992 0 -1 2076
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5844_6
timestamp 1731220559
transform 1 0 2832 0 -1 2076
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5843_6
timestamp 1731220559
transform 1 0 2648 0 -1 2076
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5842_6
timestamp 1731220559
transform 1 0 3136 0 -1 2076
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5841_6
timestamp 1731220559
transform 1 0 3264 0 -1 2076
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5840_6
timestamp 1731220559
transform 1 0 3336 0 1 2084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5839_6
timestamp 1731220559
transform 1 0 3160 0 1 2084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5838_6
timestamp 1731220559
transform 1 0 2992 0 1 2084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5837_6
timestamp 1731220559
transform 1 0 2832 0 1 2084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5836_6
timestamp 1731220559
transform 1 0 2680 0 1 2084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5835_6
timestamp 1731220559
transform 1 0 3168 0 -1 2240
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5834_6
timestamp 1731220559
transform 1 0 3000 0 -1 2240
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5833_6
timestamp 1731220559
transform 1 0 2848 0 -1 2240
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5832_6
timestamp 1731220559
transform 1 0 2712 0 -1 2240
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5831_6
timestamp 1731220559
transform 1 0 2592 0 -1 2240
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5830_6
timestamp 1731220559
transform 1 0 2584 0 1 2240
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5829_6
timestamp 1731220559
transform 1 0 2664 0 1 2240
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5828_6
timestamp 1731220559
transform 1 0 2920 0 1 2240
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5827_6
timestamp 1731220559
transform 1 0 2832 0 1 2240
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5826_6
timestamp 1731220559
transform 1 0 2744 0 1 2240
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5825_6
timestamp 1731220559
transform 1 0 2696 0 -1 2396
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5824_6
timestamp 1731220559
transform 1 0 2840 0 -1 2396
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5823_6
timestamp 1731220559
transform 1 0 3168 0 -1 2396
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5822_6
timestamp 1731220559
transform 1 0 3000 0 -1 2396
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5821_6
timestamp 1731220559
transform 1 0 2848 0 1 2400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5820_6
timestamp 1731220559
transform 1 0 2688 0 1 2400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5819_6
timestamp 1731220559
transform 1 0 3176 0 1 2400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5818_6
timestamp 1731220559
transform 1 0 3008 0 1 2400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5817_6
timestamp 1731220559
transform 1 0 3112 0 -1 2560
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5816_6
timestamp 1731220559
transform 1 0 2752 0 -1 2560
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5815_6
timestamp 1731220559
transform 1 0 2616 0 -1 2560
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5814_6
timestamp 1731220559
transform 1 0 2880 0 -1 2560
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5813_6
timestamp 1731220559
transform 1 0 3000 0 -1 2560
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5812_6
timestamp 1731220559
transform 1 0 3000 0 1 2560
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5811_6
timestamp 1731220559
transform 1 0 3272 0 1 2560
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5810_6
timestamp 1731220559
transform 1 0 3216 0 -1 2560
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5809_6
timestamp 1731220559
transform 1 0 3312 0 -1 2560
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5808_6
timestamp 1731220559
transform 1 0 3416 0 -1 2560
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5807_6
timestamp 1731220559
transform 1 0 3344 0 1 2400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5806_6
timestamp 1731220559
transform 1 0 3344 0 -1 2396
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5805_6
timestamp 1731220559
transform 1 0 3344 0 -1 2240
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5804_6
timestamp 1731220559
transform 1 0 3392 0 -1 2076
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5803_6
timestamp 1731220559
transform 1 0 3376 0 -1 1916
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5802_6
timestamp 1731220559
transform 1 0 3496 0 -1 1916
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5801_6
timestamp 1731220559
transform 1 0 3496 0 1 1924
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5800_6
timestamp 1731220559
transform 1 0 3496 0 -1 2076
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5799_6
timestamp 1731220559
transform 1 0 3496 0 1 2084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5798_6
timestamp 1731220559
transform 1 0 3496 0 -1 2240
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5797_6
timestamp 1731220559
transform 1 0 3496 0 -1 2396
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5796_6
timestamp 1731220559
transform 1 0 3496 0 1 2400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5795_6
timestamp 1731220559
transform 1 0 3496 0 -1 2560
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5794_6
timestamp 1731220559
transform 1 0 3496 0 -1 2720
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5793_6
timestamp 1731220559
transform 1 0 3496 0 1 2720
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5792_6
timestamp 1731220559
transform 1 0 3496 0 -1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5791_6
timestamp 1731220559
transform 1 0 3480 0 1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5790_6
timestamp 1731220559
transform 1 0 3352 0 -1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5789_6
timestamp 1731220559
transform 1 0 3368 0 1 2720
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5788_6
timestamp 1731220559
transform 1 0 3368 0 -1 2720
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5787_6
timestamp 1731220559
transform 1 0 3216 0 -1 2720
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5786_6
timestamp 1731220559
transform 1 0 3064 0 -1 2720
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5785_6
timestamp 1731220559
transform 1 0 2904 0 -1 2720
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5784_6
timestamp 1731220559
transform 1 0 2728 0 -1 2720
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5783_6
timestamp 1731220559
transform 1 0 3216 0 1 2720
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5782_6
timestamp 1731220559
transform 1 0 3072 0 1 2720
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5781_6
timestamp 1731220559
transform 1 0 2928 0 1 2720
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5780_6
timestamp 1731220559
transform 1 0 2776 0 1 2720
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5779_6
timestamp 1731220559
transform 1 0 2624 0 1 2720
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5778_6
timestamp 1731220559
transform 1 0 3024 0 -1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5777_6
timestamp 1731220559
transform 1 0 3184 0 -1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5776_6
timestamp 1731220559
transform 1 0 3320 0 1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5775_6
timestamp 1731220559
transform 1 0 3168 0 1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5774_6
timestamp 1731220559
transform 1 0 3032 0 -1 3048
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5773_6
timestamp 1731220559
transform 1 0 3176 0 -1 3048
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5772_6
timestamp 1731220559
transform 1 0 3320 0 -1 3048
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5771_6
timestamp 1731220559
transform 1 0 3184 0 1 3060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5770_6
timestamp 1731220559
transform 1 0 3000 0 1 3060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5769_6
timestamp 1731220559
transform 1 0 3376 0 1 3060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5768_6
timestamp 1731220559
transform 1 0 3320 0 -1 3212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5767_6
timestamp 1731220559
transform 1 0 3144 0 -1 3212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5766_6
timestamp 1731220559
transform 1 0 3496 0 -1 3212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5765_6
timestamp 1731220559
transform 1 0 3496 0 1 3212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5764_6
timestamp 1731220559
transform 1 0 3496 0 -1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5763_6
timestamp 1731220559
transform 1 0 3496 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5762_6
timestamp 1731220559
transform 1 0 3496 0 -1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5761_6
timestamp 1731220559
transform 1 0 3408 0 -1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5760_6
timestamp 1731220559
transform 1 0 3296 0 -1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5759_6
timestamp 1731220559
transform 1 0 3184 0 -1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5758_6
timestamp 1731220559
transform 1 0 3072 0 -1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5757_6
timestamp 1731220559
transform 1 0 2952 0 -1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5756_6
timestamp 1731220559
transform 1 0 2960 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5755_6
timestamp 1731220559
transform 1 0 3248 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5754_6
timestamp 1731220559
transform 1 0 3104 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5753_6
timestamp 1731220559
transform 1 0 3008 0 -1 3668
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5752_6
timestamp 1731220559
transform 1 0 2720 0 -1 3668
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5751_6
timestamp 1731220559
transform 1 0 2432 0 -1 3668
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5750_6
timestamp 1731220559
transform 1 0 2816 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5749_6
timestamp 1731220559
transform 1 0 2680 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5748_6
timestamp 1731220559
transform 1 0 2664 0 -1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5747_6
timestamp 1731220559
transform 1 0 2816 0 -1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5746_6
timestamp 1731220559
transform 1 0 2816 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5745_6
timestamp 1731220559
transform 1 0 2984 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5744_6
timestamp 1731220559
transform 1 0 3152 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5743_6
timestamp 1731220559
transform 1 0 3328 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5742_6
timestamp 1731220559
transform 1 0 3344 0 -1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5741_6
timestamp 1731220559
transform 1 0 3176 0 -1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5740_6
timestamp 1731220559
transform 1 0 3016 0 -1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5739_6
timestamp 1731220559
transform 1 0 2864 0 -1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5738_6
timestamp 1731220559
transform 1 0 2720 0 -1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5737_6
timestamp 1731220559
transform 1 0 3296 0 1 3212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5736_6
timestamp 1731220559
transform 1 0 3096 0 1 3212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5735_6
timestamp 1731220559
transform 1 0 2904 0 1 3212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5734_6
timestamp 1731220559
transform 1 0 2728 0 1 3212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5733_6
timestamp 1731220559
transform 1 0 2576 0 1 3212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5732_6
timestamp 1731220559
transform 1 0 2616 0 -1 3212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5731_6
timestamp 1731220559
transform 1 0 2792 0 -1 3212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5730_6
timestamp 1731220559
transform 1 0 2968 0 -1 3212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5729_6
timestamp 1731220559
transform 1 0 2816 0 1 3060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5728_6
timestamp 1731220559
transform 1 0 2632 0 1 3060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5727_6
timestamp 1731220559
transform 1 0 2616 0 -1 3048
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5726_6
timestamp 1731220559
transform 1 0 2760 0 -1 3048
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5725_6
timestamp 1731220559
transform 1 0 2896 0 -1 3048
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5724_6
timestamp 1731220559
transform 1 0 3024 0 1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5723_6
timestamp 1731220559
transform 1 0 2896 0 1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5722_6
timestamp 1731220559
transform 1 0 2872 0 -1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5721_6
timestamp 1731220559
transform 1 0 2720 0 -1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5720_6
timestamp 1731220559
transform 1 0 2584 0 -1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5719_6
timestamp 1731220559
transform 1 0 2776 0 1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5718_6
timestamp 1731220559
transform 1 0 2680 0 1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5717_6
timestamp 1731220559
transform 1 0 2592 0 1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5716_6
timestamp 1731220559
transform 1 0 2512 0 1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5715_6
timestamp 1731220559
transform 1 0 2432 0 1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5714_6
timestamp 1731220559
transform 1 0 2352 0 1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5713_6
timestamp 1731220559
transform 1 0 2272 0 1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5712_6
timestamp 1731220559
transform 1 0 2232 0 -1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5711_6
timestamp 1731220559
transform 1 0 2336 0 -1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5710_6
timestamp 1731220559
transform 1 0 2456 0 -1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5709_6
timestamp 1731220559
transform 1 0 2472 0 1 2720
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5708_6
timestamp 1731220559
transform 1 0 2000 0 1 2720
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5707_6
timestamp 1731220559
transform 1 0 1888 0 1 2720
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5706_6
timestamp 1731220559
transform 1 0 2096 0 -1 2720
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5705_6
timestamp 1731220559
transform 1 0 1888 0 -1 2720
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5704_6
timestamp 1731220559
transform 1 0 1736 0 -1 2748
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5703_6
timestamp 1731220559
transform 1 0 1600 0 -1 2748
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5702_6
timestamp 1731220559
transform 1 0 1736 0 1 2752
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5701_6
timestamp 1731220559
transform 1 0 1632 0 1 2752
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5700_6
timestamp 1731220559
transform 1 0 1512 0 1 2752
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5699_6
timestamp 1731220559
transform 1 0 1392 0 1 2752
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5698_6
timestamp 1731220559
transform 1 0 1688 0 -1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5697_6
timestamp 1731220559
transform 1 0 1584 0 -1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5696_6
timestamp 1731220559
transform 1 0 1480 0 -1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5695_6
timestamp 1731220559
transform 1 0 1384 0 -1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5694_6
timestamp 1731220559
transform 1 0 1632 0 1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5693_6
timestamp 1731220559
transform 1 0 1520 0 1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5692_6
timestamp 1731220559
transform 1 0 1408 0 1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5691_6
timestamp 1731220559
transform 1 0 1296 0 1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5690_6
timestamp 1731220559
transform 1 0 1184 0 1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5689_6
timestamp 1731220559
transform 1 0 1064 0 1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5688_6
timestamp 1731220559
transform 1 0 928 0 1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5687_6
timestamp 1731220559
transform 1 0 1280 0 -1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5686_6
timestamp 1731220559
transform 1 0 1168 0 -1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5685_6
timestamp 1731220559
transform 1 0 1048 0 -1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5684_6
timestamp 1731220559
transform 1 0 920 0 -1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5683_6
timestamp 1731220559
transform 1 0 984 0 1 2752
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5682_6
timestamp 1731220559
transform 1 0 1264 0 1 2752
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5681_6
timestamp 1731220559
transform 1 0 1128 0 1 2752
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5680_6
timestamp 1731220559
transform 1 0 1128 0 -1 2748
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5679_6
timestamp 1731220559
transform 1 0 968 0 -1 2748
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5678_6
timestamp 1731220559
transform 1 0 1280 0 -1 2748
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5677_6
timestamp 1731220559
transform 1 0 1440 0 -1 2748
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5676_6
timestamp 1731220559
transform 1 0 1536 0 1 2588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5675_6
timestamp 1731220559
transform 1 0 1384 0 1 2588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5674_6
timestamp 1731220559
transform 1 0 1232 0 1 2588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5673_6
timestamp 1731220559
transform 1 0 1088 0 1 2588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5672_6
timestamp 1731220559
transform 1 0 936 0 1 2588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5671_6
timestamp 1731220559
transform 1 0 1040 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5670_6
timestamp 1731220559
transform 1 0 1200 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5669_6
timestamp 1731220559
transform 1 0 1352 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5668_6
timestamp 1731220559
transform 1 0 1504 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5667_6
timestamp 1731220559
transform 1 0 1664 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5666_6
timestamp 1731220559
transform 1 0 1656 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5665_6
timestamp 1731220559
transform 1 0 1536 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5664_6
timestamp 1731220559
transform 1 0 1416 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5663_6
timestamp 1731220559
transform 1 0 1296 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5662_6
timestamp 1731220559
transform 1 0 1176 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5661_6
timestamp 1731220559
transform 1 0 1048 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5660_6
timestamp 1731220559
transform 1 0 1456 0 -1 2416
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5659_6
timestamp 1731220559
transform 1 0 1376 0 -1 2416
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5658_6
timestamp 1731220559
transform 1 0 1296 0 -1 2416
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5657_6
timestamp 1731220559
transform 1 0 1216 0 -1 2416
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5656_6
timestamp 1731220559
transform 1 0 1136 0 -1 2416
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5655_6
timestamp 1731220559
transform 1 0 1056 0 -1 2416
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5654_6
timestamp 1731220559
transform 1 0 1304 0 1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5653_6
timestamp 1731220559
transform 1 0 1224 0 1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5652_6
timestamp 1731220559
transform 1 0 1144 0 1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5651_6
timestamp 1731220559
transform 1 0 1064 0 1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5650_6
timestamp 1731220559
transform 1 0 984 0 1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5649_6
timestamp 1731220559
transform 1 0 1248 0 -1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5648_6
timestamp 1731220559
transform 1 0 1168 0 -1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5647_6
timestamp 1731220559
transform 1 0 1088 0 -1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5646_6
timestamp 1731220559
transform 1 0 1008 0 -1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5645_6
timestamp 1731220559
transform 1 0 928 0 -1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5644_6
timestamp 1731220559
transform 1 0 848 0 -1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5643_6
timestamp 1731220559
transform 1 0 848 0 1 2092
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5642_6
timestamp 1731220559
transform 1 0 936 0 1 2092
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5641_6
timestamp 1731220559
transform 1 0 1024 0 1 2092
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5640_6
timestamp 1731220559
transform 1 0 1112 0 1 2092
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5639_6
timestamp 1731220559
transform 1 0 1208 0 1 2092
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5638_6
timestamp 1731220559
transform 1 0 1168 0 -1 2080
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5637_6
timestamp 1731220559
transform 1 0 1056 0 -1 2080
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5636_6
timestamp 1731220559
transform 1 0 936 0 -1 2080
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5635_6
timestamp 1731220559
transform 1 0 1000 0 1 1924
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5634_6
timestamp 1731220559
transform 1 0 1152 0 1 1924
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5633_6
timestamp 1731220559
transform 1 0 1152 0 -1 1920
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5632_6
timestamp 1731220559
transform 1 0 1000 0 -1 1920
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5631_6
timestamp 1731220559
transform 1 0 1008 0 1 1764
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5630_6
timestamp 1731220559
transform 1 0 1160 0 -1 1756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5629_6
timestamp 1731220559
transform 1 0 1000 0 -1 1756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5628_6
timestamp 1731220559
transform 1 0 1016 0 1 1600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5627_6
timestamp 1731220559
transform 1 0 1112 0 -1 1600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5626_6
timestamp 1731220559
transform 1 0 976 0 -1 1600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5625_6
timestamp 1731220559
transform 1 0 1000 0 1 1444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5624_6
timestamp 1731220559
transform 1 0 888 0 1 1444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5623_6
timestamp 1731220559
transform 1 0 912 0 -1 1436
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5622_6
timestamp 1731220559
transform 1 0 848 0 1 1284
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5621_6
timestamp 1731220559
transform 1 0 992 0 1 1284
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5620_6
timestamp 1731220559
transform 1 0 1128 0 1 1284
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5619_6
timestamp 1731220559
transform 1 0 1096 0 -1 1280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5618_6
timestamp 1731220559
transform 1 0 952 0 -1 1280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5617_6
timestamp 1731220559
transform 1 0 808 0 -1 1280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5616_6
timestamp 1731220559
transform 1 0 744 0 1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5615_6
timestamp 1731220559
transform 1 0 912 0 1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5614_6
timestamp 1731220559
transform 1 0 840 0 -1 1124
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5613_6
timestamp 1731220559
transform 1 0 704 0 -1 1124
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5612_6
timestamp 1731220559
transform 1 0 560 0 -1 1124
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5611_6
timestamp 1731220559
transform 1 0 536 0 1 964
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5610_6
timestamp 1731220559
transform 1 0 672 0 1 964
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5609_6
timestamp 1731220559
transform 1 0 680 0 -1 956
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5608_6
timestamp 1731220559
transform 1 0 560 0 -1 956
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5607_6
timestamp 1731220559
transform 1 0 544 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5606_6
timestamp 1731220559
transform 1 0 704 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5605_6
timestamp 1731220559
transform 1 0 856 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5604_6
timestamp 1731220559
transform 1 0 776 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5603_6
timestamp 1731220559
transform 1 0 944 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5602_6
timestamp 1731220559
transform 1 0 888 0 1 620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5601_6
timestamp 1731220559
transform 1 0 768 0 1 620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5600_6
timestamp 1731220559
transform 1 0 640 0 1 620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5599_6
timestamp 1731220559
transform 1 0 728 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5598_6
timestamp 1731220559
transform 1 0 640 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5597_6
timestamp 1731220559
transform 1 0 520 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5596_6
timestamp 1731220559
transform 1 0 424 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5595_6
timestamp 1731220559
transform 1 0 488 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5594_6
timestamp 1731220559
transform 1 0 600 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5593_6
timestamp 1731220559
transform 1 0 712 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5592_6
timestamp 1731220559
transform 1 0 760 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5591_6
timestamp 1731220559
transform 1 0 632 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5590_6
timestamp 1731220559
transform 1 0 592 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5589_6
timestamp 1731220559
transform 1 0 728 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5588_6
timestamp 1731220559
transform 1 0 864 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5587_6
timestamp 1731220559
transform 1 0 808 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5586_6
timestamp 1731220559
transform 1 0 720 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5585_6
timestamp 1731220559
transform 1 0 632 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5584_6
timestamp 1731220559
transform 1 0 544 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5583_6
timestamp 1731220559
transform 1 0 464 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5582_6
timestamp 1731220559
transform 1 0 384 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5581_6
timestamp 1731220559
transform 1 0 304 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5580_6
timestamp 1731220559
transform 1 0 224 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5579_6
timestamp 1731220559
transform 1 0 144 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5578_6
timestamp 1731220559
transform 1 0 216 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5577_6
timestamp 1731220559
transform 1 0 328 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5576_6
timestamp 1731220559
transform 1 0 456 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5575_6
timestamp 1731220559
transform 1 0 496 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5574_6
timestamp 1731220559
transform 1 0 360 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5573_6
timestamp 1731220559
transform 1 0 232 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5572_6
timestamp 1731220559
transform 1 0 128 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5571_6
timestamp 1731220559
transform 1 0 128 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5570_6
timestamp 1731220559
transform 1 0 240 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5569_6
timestamp 1731220559
transform 1 0 368 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5568_6
timestamp 1731220559
transform 1 0 328 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5567_6
timestamp 1731220559
transform 1 0 224 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5566_6
timestamp 1731220559
transform 1 0 304 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5565_6
timestamp 1731220559
transform 1 0 384 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5564_6
timestamp 1731220559
transform 1 0 464 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5563_6
timestamp 1731220559
transform 1 0 552 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5562_6
timestamp 1731220559
transform 1 0 512 0 1 620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5561_6
timestamp 1731220559
transform 1 0 392 0 1 620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5560_6
timestamp 1731220559
transform 1 0 280 0 1 620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5559_6
timestamp 1731220559
transform 1 0 600 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5558_6
timestamp 1731220559
transform 1 0 424 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5557_6
timestamp 1731220559
transform 1 0 256 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5556_6
timestamp 1731220559
transform 1 0 128 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5555_6
timestamp 1731220559
transform 1 0 128 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5554_6
timestamp 1731220559
transform 1 0 240 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5553_6
timestamp 1731220559
transform 1 0 384 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5552_6
timestamp 1731220559
transform 1 0 440 0 -1 956
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5551_6
timestamp 1731220559
transform 1 0 320 0 -1 956
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5550_6
timestamp 1731220559
transform 1 0 208 0 -1 956
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5549_6
timestamp 1731220559
transform 1 0 128 0 -1 956
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5548_6
timestamp 1731220559
transform 1 0 128 0 1 964
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5547_6
timestamp 1731220559
transform 1 0 392 0 1 964
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5546_6
timestamp 1731220559
transform 1 0 248 0 1 964
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5545_6
timestamp 1731220559
transform 1 0 136 0 -1 1124
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5544_6
timestamp 1731220559
transform 1 0 272 0 -1 1124
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5543_6
timestamp 1731220559
transform 1 0 416 0 -1 1124
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5542_6
timestamp 1731220559
transform 1 0 576 0 1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5541_6
timestamp 1731220559
transform 1 0 400 0 1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5540_6
timestamp 1731220559
transform 1 0 224 0 1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5539_6
timestamp 1731220559
transform 1 0 304 0 -1 1280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5538_6
timestamp 1731220559
transform 1 0 408 0 -1 1280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5537_6
timestamp 1731220559
transform 1 0 528 0 -1 1280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5536_6
timestamp 1731220559
transform 1 0 664 0 -1 1280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5535_6
timestamp 1731220559
transform 1 0 712 0 1 1284
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5534_6
timestamp 1731220559
transform 1 0 576 0 1 1284
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5533_6
timestamp 1731220559
transform 1 0 456 0 1 1284
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5532_6
timestamp 1731220559
transform 1 0 344 0 1 1284
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5531_6
timestamp 1731220559
transform 1 0 248 0 -1 1436
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5530_6
timestamp 1731220559
transform 1 0 344 0 -1 1436
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5529_6
timestamp 1731220559
transform 1 0 440 0 -1 1436
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5528_6
timestamp 1731220559
transform 1 0 360 0 1 1444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5527_6
timestamp 1731220559
transform 1 0 216 0 1 1444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5526_6
timestamp 1731220559
transform 1 0 280 0 -1 1600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5525_6
timestamp 1731220559
transform 1 0 152 0 -1 1600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5524_6
timestamp 1731220559
transform 1 0 128 0 1 1600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5523_6
timestamp 1731220559
transform 1 0 280 0 1 1600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5522_6
timestamp 1731220559
transform 1 0 336 0 -1 1756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5521_6
timestamp 1731220559
transform 1 0 208 0 -1 1756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5520_6
timestamp 1731220559
transform 1 0 128 0 -1 1756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5519_6
timestamp 1731220559
transform 1 0 128 0 1 1764
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5518_6
timestamp 1731220559
transform 1 0 272 0 1 1764
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5517_6
timestamp 1731220559
transform 1 0 368 0 -1 1920
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5516_6
timestamp 1731220559
transform 1 0 232 0 -1 1920
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5515_6
timestamp 1731220559
transform 1 0 128 0 -1 1920
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5514_6
timestamp 1731220559
transform 1 0 176 0 1 1924
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5513_6
timestamp 1731220559
transform 1 0 336 0 1 1924
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5512_6
timestamp 1731220559
transform 1 0 440 0 -1 2080
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5511_6
timestamp 1731220559
transform 1 0 320 0 -1 2080
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5510_6
timestamp 1731220559
transform 1 0 200 0 -1 2080
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5509_6
timestamp 1731220559
transform 1 0 296 0 1 2092
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5508_6
timestamp 1731220559
transform 1 0 392 0 1 2092
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5507_6
timestamp 1731220559
transform 1 0 488 0 1 2092
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5506_6
timestamp 1731220559
transform 1 0 528 0 -1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5505_6
timestamp 1731220559
transform 1 0 448 0 -1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5504_6
timestamp 1731220559
transform 1 0 368 0 -1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5503_6
timestamp 1731220559
transform 1 0 344 0 1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5502_6
timestamp 1731220559
transform 1 0 424 0 1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5501_6
timestamp 1731220559
transform 1 0 504 0 1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5500_6
timestamp 1731220559
transform 1 0 584 0 1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5499_6
timestamp 1731220559
transform 1 0 664 0 1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5498_6
timestamp 1731220559
transform 1 0 744 0 1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5497_6
timestamp 1731220559
transform 1 0 904 0 1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5496_6
timestamp 1731220559
transform 1 0 824 0 1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5495_6
timestamp 1731220559
transform 1 0 768 0 -1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5494_6
timestamp 1731220559
transform 1 0 688 0 -1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5493_6
timestamp 1731220559
transform 1 0 608 0 -1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5492_6
timestamp 1731220559
transform 1 0 760 0 1 2092
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5491_6
timestamp 1731220559
transform 1 0 672 0 1 2092
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5490_6
timestamp 1731220559
transform 1 0 584 0 1 2092
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5489_6
timestamp 1731220559
transform 1 0 568 0 -1 2080
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5488_6
timestamp 1731220559
transform 1 0 696 0 -1 2080
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5487_6
timestamp 1731220559
transform 1 0 816 0 -1 2080
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5486_6
timestamp 1731220559
transform 1 0 840 0 1 1924
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5485_6
timestamp 1731220559
transform 1 0 672 0 1 1924
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5484_6
timestamp 1731220559
transform 1 0 504 0 1 1924
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5483_6
timestamp 1731220559
transform 1 0 520 0 -1 1920
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5482_6
timestamp 1731220559
transform 1 0 680 0 -1 1920
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5481_6
timestamp 1731220559
transform 1 0 840 0 -1 1920
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5480_6
timestamp 1731220559
transform 1 0 832 0 1 1764
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5479_6
timestamp 1731220559
transform 1 0 648 0 1 1764
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5478_6
timestamp 1731220559
transform 1 0 456 0 1 1764
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5477_6
timestamp 1731220559
transform 1 0 488 0 -1 1756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5476_6
timestamp 1731220559
transform 1 0 656 0 -1 1756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5475_6
timestamp 1731220559
transform 1 0 832 0 -1 1756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5474_6
timestamp 1731220559
transform 1 0 656 0 1 1600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5473_6
timestamp 1731220559
transform 1 0 464 0 1 1600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5472_6
timestamp 1731220559
transform 1 0 840 0 1 1600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5471_6
timestamp 1731220559
transform 1 0 840 0 -1 1600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5470_6
timestamp 1731220559
transform 1 0 704 0 -1 1600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5469_6
timestamp 1731220559
transform 1 0 560 0 -1 1600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5468_6
timestamp 1731220559
transform 1 0 416 0 -1 1600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5467_6
timestamp 1731220559
transform 1 0 504 0 1 1444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5466_6
timestamp 1731220559
transform 1 0 768 0 1 1444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5465_6
timestamp 1731220559
transform 1 0 640 0 1 1444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5464_6
timestamp 1731220559
transform 1 0 624 0 -1 1436
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5463_6
timestamp 1731220559
transform 1 0 536 0 -1 1436
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5462_6
timestamp 1731220559
transform 1 0 712 0 -1 1436
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5461_6
timestamp 1731220559
transform 1 0 800 0 -1 1436
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5460_6
timestamp 1731220559
transform 1 0 1040 0 -1 1436
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5459_6
timestamp 1731220559
transform 1 0 1200 0 -1 1436
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5458_6
timestamp 1731220559
transform 1 0 1568 0 -1 1436
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5457_6
timestamp 1731220559
transform 1 0 1376 0 -1 1436
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5456_6
timestamp 1731220559
transform 1 0 1304 0 1 1444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5455_6
timestamp 1731220559
transform 1 0 1200 0 1 1444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5454_6
timestamp 1731220559
transform 1 0 1104 0 1 1444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5453_6
timestamp 1731220559
transform 1 0 1408 0 1 1444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5452_6
timestamp 1731220559
transform 1 0 1504 0 -1 1600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5451_6
timestamp 1731220559
transform 1 0 1368 0 -1 1600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5450_6
timestamp 1731220559
transform 1 0 1240 0 -1 1600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5449_6
timestamp 1731220559
transform 1 0 1184 0 1 1600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5448_6
timestamp 1731220559
transform 1 0 1344 0 1 1600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5447_6
timestamp 1731220559
transform 1 0 1504 0 1 1600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5446_6
timestamp 1731220559
transform 1 0 1664 0 1 1600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5445_6
timestamp 1731220559
transform 1 0 1736 0 -1 1756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5444_6
timestamp 1731220559
transform 1 0 1600 0 -1 1756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5443_6
timestamp 1731220559
transform 1 0 1456 0 -1 1756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5442_6
timestamp 1731220559
transform 1 0 1312 0 -1 1756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5441_6
timestamp 1731220559
transform 1 0 1664 0 1 1764
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5440_6
timestamp 1731220559
transform 1 0 1496 0 1 1764
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5439_6
timestamp 1731220559
transform 1 0 1336 0 1 1764
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5438_6
timestamp 1731220559
transform 1 0 1176 0 1 1764
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5437_6
timestamp 1731220559
transform 1 0 1296 0 -1 1920
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5436_6
timestamp 1731220559
transform 1 0 1448 0 -1 1920
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5435_6
timestamp 1731220559
transform 1 0 1600 0 -1 1920
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5434_6
timestamp 1731220559
transform 1 0 1704 0 1 1924
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5433_6
timestamp 1731220559
transform 1 0 1568 0 1 1924
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5432_6
timestamp 1731220559
transform 1 0 1432 0 1 1924
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5431_6
timestamp 1731220559
transform 1 0 1296 0 1 1924
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5430_6
timestamp 1731220559
transform 1 0 1272 0 -1 2080
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5429_6
timestamp 1731220559
transform 1 0 1368 0 -1 2080
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5428_6
timestamp 1731220559
transform 1 0 1464 0 -1 2080
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5427_6
timestamp 1731220559
transform 1 0 1560 0 -1 2080
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5426_6
timestamp 1731220559
transform 1 0 1656 0 -1 2080
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5425_6
timestamp 1731220559
transform 1 0 1736 0 -1 2080
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5424_6
timestamp 1731220559
transform 1 0 1888 0 1 2084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5423_6
timestamp 1731220559
transform 1 0 1968 0 1 2084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5422_6
timestamp 1731220559
transform 1 0 2376 0 1 2084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5421_6
timestamp 1731220559
transform 1 0 2232 0 1 2084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5420_6
timestamp 1731220559
transform 1 0 2096 0 1 2084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5419_6
timestamp 1731220559
transform 1 0 1960 0 -1 2076
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5418_6
timestamp 1731220559
transform 1 0 1944 0 1 1924
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5417_6
timestamp 1731220559
transform 1 0 2064 0 1 1924
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5416_6
timestamp 1731220559
transform 1 0 2184 0 1 1924
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5415_6
timestamp 1731220559
transform 1 0 2144 0 -1 1916
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5414_6
timestamp 1731220559
transform 1 0 2056 0 -1 1916
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5413_6
timestamp 1731220559
transform 1 0 2080 0 1 1748
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5412_6
timestamp 1731220559
transform 1 0 2224 0 1 1748
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5411_6
timestamp 1731220559
transform 1 0 2384 0 1 1748
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5410_6
timestamp 1731220559
transform 1 0 2376 0 -1 1744
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5409_6
timestamp 1731220559
transform 1 0 2232 0 -1 1744
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5408_6
timestamp 1731220559
transform 1 0 2096 0 -1 1744
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5407_6
timestamp 1731220559
transform 1 0 2336 0 1 1588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5406_6
timestamp 1731220559
transform 1 0 2200 0 1 1588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5405_6
timestamp 1731220559
transform 1 0 2072 0 1 1588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5404_6
timestamp 1731220559
transform 1 0 1952 0 1 1588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5403_6
timestamp 1731220559
transform 1 0 1888 0 -1 1580
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5402_6
timestamp 1731220559
transform 1 0 2040 0 -1 1580
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5401_6
timestamp 1731220559
transform 1 0 2200 0 -1 1580
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5400_6
timestamp 1731220559
transform 1 0 2120 0 1 1420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5399_6
timestamp 1731220559
transform 1 0 1992 0 1 1420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5398_6
timestamp 1731220559
transform 1 0 1888 0 1 1420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5397_6
timestamp 1731220559
transform 1 0 1888 0 -1 1420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5396_6
timestamp 1731220559
transform 1 0 1736 0 -1 1436
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5395_6
timestamp 1731220559
transform 1 0 1736 0 1 1284
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5394_6
timestamp 1731220559
transform 1 0 1632 0 1 1284
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5393_6
timestamp 1731220559
transform 1 0 1512 0 1 1284
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5392_6
timestamp 1731220559
transform 1 0 1392 0 1 1284
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5391_6
timestamp 1731220559
transform 1 0 1264 0 1 1284
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5390_6
timestamp 1731220559
transform 1 0 1624 0 -1 1280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5389_6
timestamp 1731220559
transform 1 0 1496 0 -1 1280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5388_6
timestamp 1731220559
transform 1 0 1368 0 -1 1280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5387_6
timestamp 1731220559
transform 1 0 1232 0 -1 1280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5386_6
timestamp 1731220559
transform 1 0 1624 0 1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5385_6
timestamp 1731220559
transform 1 0 1488 0 1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5384_6
timestamp 1731220559
transform 1 0 1352 0 1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5383_6
timestamp 1731220559
transform 1 0 1208 0 1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5382_6
timestamp 1731220559
transform 1 0 1064 0 1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5381_6
timestamp 1731220559
transform 1 0 1464 0 -1 1124
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5380_6
timestamp 1731220559
transform 1 0 1336 0 -1 1124
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5379_6
timestamp 1731220559
transform 1 0 1216 0 -1 1124
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5378_6
timestamp 1731220559
transform 1 0 1096 0 -1 1124
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5377_6
timestamp 1731220559
transform 1 0 968 0 -1 1124
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5376_6
timestamp 1731220559
transform 1 0 1344 0 1 964
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5375_6
timestamp 1731220559
transform 1 0 1232 0 1 964
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5374_6
timestamp 1731220559
transform 1 0 1128 0 1 964
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5373_6
timestamp 1731220559
transform 1 0 1024 0 1 964
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5372_6
timestamp 1731220559
transform 1 0 912 0 1 964
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5371_6
timestamp 1731220559
transform 1 0 792 0 1 964
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5370_6
timestamp 1731220559
transform 1 0 792 0 -1 956
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5369_6
timestamp 1731220559
transform 1 0 904 0 -1 956
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5368_6
timestamp 1731220559
transform 1 0 1008 0 -1 956
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5367_6
timestamp 1731220559
transform 1 0 1112 0 -1 956
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5366_6
timestamp 1731220559
transform 1 0 1320 0 -1 956
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5365_6
timestamp 1731220559
transform 1 0 1216 0 -1 956
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5364_6
timestamp 1731220559
transform 1 0 1136 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5363_6
timestamp 1731220559
transform 1 0 1000 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5362_6
timestamp 1731220559
transform 1 0 1264 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5361_6
timestamp 1731220559
transform 1 0 1384 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5360_6
timestamp 1731220559
transform 1 0 1504 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5359_6
timestamp 1731220559
transform 1 0 1632 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5358_6
timestamp 1731220559
transform 1 0 1736 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5357_6
timestamp 1731220559
transform 1 0 1632 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5356_6
timestamp 1731220559
transform 1 0 1504 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5355_6
timestamp 1731220559
transform 1 0 1376 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5354_6
timestamp 1731220559
transform 1 0 1240 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5353_6
timestamp 1731220559
transform 1 0 1096 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5352_6
timestamp 1731220559
transform 1 0 1544 0 1 620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5351_6
timestamp 1731220559
transform 1 0 1440 0 1 620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5350_6
timestamp 1731220559
transform 1 0 1336 0 1 620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5349_6
timestamp 1731220559
transform 1 0 1232 0 1 620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5348_6
timestamp 1731220559
transform 1 0 1120 0 1 620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5347_6
timestamp 1731220559
transform 1 0 1008 0 1 620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5346_6
timestamp 1731220559
transform 1 0 1256 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5345_6
timestamp 1731220559
transform 1 0 1168 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5344_6
timestamp 1731220559
transform 1 0 1080 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5343_6
timestamp 1731220559
transform 1 0 992 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5342_6
timestamp 1731220559
transform 1 0 904 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5341_6
timestamp 1731220559
transform 1 0 816 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5340_6
timestamp 1731220559
transform 1 0 1232 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5339_6
timestamp 1731220559
transform 1 0 1144 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5338_6
timestamp 1731220559
transform 1 0 1056 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5337_6
timestamp 1731220559
transform 1 0 968 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5336_6
timestamp 1731220559
transform 1 0 880 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5335_6
timestamp 1731220559
transform 1 0 792 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5334_6
timestamp 1731220559
transform 1 0 704 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5333_6
timestamp 1731220559
transform 1 0 616 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5332_6
timestamp 1731220559
transform 1 0 816 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5331_6
timestamp 1731220559
transform 1 0 912 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5330_6
timestamp 1731220559
transform 1 0 1000 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5329_6
timestamp 1731220559
transform 1 0 1096 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5328_6
timestamp 1731220559
transform 1 0 1288 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5327_6
timestamp 1731220559
transform 1 0 1192 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5326_6
timestamp 1731220559
transform 1 0 1104 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5325_6
timestamp 1731220559
transform 1 0 992 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5324_6
timestamp 1731220559
transform 1 0 880 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5323_6
timestamp 1731220559
transform 1 0 1208 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5322_6
timestamp 1731220559
transform 1 0 1424 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5321_6
timestamp 1731220559
transform 1 0 1312 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5320_6
timestamp 1731220559
transform 1 0 1248 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5319_6
timestamp 1731220559
transform 1 0 1128 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5318_6
timestamp 1731220559
transform 1 0 1000 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5317_6
timestamp 1731220559
transform 1 0 1592 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5316_6
timestamp 1731220559
transform 1 0 1472 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5315_6
timestamp 1731220559
transform 1 0 1360 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5314_6
timestamp 1731220559
transform 1 0 1072 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5313_6
timestamp 1731220559
transform 1 0 984 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5312_6
timestamp 1731220559
transform 1 0 896 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5311_6
timestamp 1731220559
transform 1 0 1152 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5310_6
timestamp 1731220559
transform 1 0 1232 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5309_6
timestamp 1731220559
transform 1 0 1320 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5308_6
timestamp 1731220559
transform 1 0 1408 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5307_6
timestamp 1731220559
transform 1 0 1496 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5306_6
timestamp 1731220559
transform 1 0 1576 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5305_6
timestamp 1731220559
transform 1 0 1656 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5304_6
timestamp 1731220559
transform 1 0 1736 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5303_6
timestamp 1731220559
transform 1 0 1888 0 1 108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5302_6
timestamp 1731220559
transform 1 0 1968 0 1 108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5301_6
timestamp 1731220559
transform 1 0 2072 0 1 108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5300_6
timestamp 1731220559
transform 1 0 2448 0 1 108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5299_6
timestamp 1731220559
transform 1 0 2320 0 1 108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5298_6
timestamp 1731220559
transform 1 0 2192 0 1 108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5297_6
timestamp 1731220559
transform 1 0 2088 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5296_6
timestamp 1731220559
transform 1 0 1976 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5295_6
timestamp 1731220559
transform 1 0 1888 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5294_6
timestamp 1731220559
transform 1 0 2496 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5293_6
timestamp 1731220559
transform 1 0 2352 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5292_6
timestamp 1731220559
transform 1 0 2216 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5291_6
timestamp 1731220559
transform 1 0 2152 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5290_6
timestamp 1731220559
transform 1 0 2064 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5289_6
timestamp 1731220559
transform 1 0 2248 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5288_6
timestamp 1731220559
transform 1 0 2360 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5287_6
timestamp 1731220559
transform 1 0 2624 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5286_6
timestamp 1731220559
transform 1 0 2488 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5285_6
timestamp 1731220559
transform 1 0 2408 0 -1 440
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5284_6
timestamp 1731220559
transform 1 0 2328 0 -1 440
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5283_6
timestamp 1731220559
transform 1 0 2488 0 -1 440
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5282_6
timestamp 1731220559
transform 1 0 2576 0 -1 440
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5281_6
timestamp 1731220559
transform 1 0 2680 0 -1 440
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5280_6
timestamp 1731220559
transform 1 0 2672 0 1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5279_6
timestamp 1731220559
transform 1 0 2536 0 1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5278_6
timestamp 1731220559
transform 1 0 2416 0 1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5277_6
timestamp 1731220559
transform 1 0 2312 0 1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5276_6
timestamp 1731220559
transform 1 0 2216 0 1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5275_6
timestamp 1731220559
transform 1 0 2136 0 1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5274_6
timestamp 1731220559
transform 1 0 2488 0 -1 596
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5273_6
timestamp 1731220559
transform 1 0 2344 0 -1 596
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5272_6
timestamp 1731220559
transform 1 0 2208 0 -1 596
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5271_6
timestamp 1731220559
transform 1 0 2080 0 -1 596
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5270_6
timestamp 1731220559
transform 1 0 1968 0 -1 596
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5269_6
timestamp 1731220559
transform 1 0 1888 0 -1 596
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5268_6
timestamp 1731220559
transform 1 0 1888 0 1 600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5267_6
timestamp 1731220559
transform 1 0 1736 0 1 620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5266_6
timestamp 1731220559
transform 1 0 1648 0 1 620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5265_6
timestamp 1731220559
transform 1 0 2280 0 1 600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5264_6
timestamp 1731220559
transform 1 0 2080 0 1 600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5263_6
timestamp 1731220559
transform 1 0 2064 0 -1 756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5262_6
timestamp 1731220559
transform 1 0 1968 0 -1 756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5261_6
timestamp 1731220559
transform 1 0 1888 0 -1 756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5260_6
timestamp 1731220559
transform 1 0 2176 0 -1 756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5259_6
timestamp 1731220559
transform 1 0 2440 0 -1 756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5258_6
timestamp 1731220559
transform 1 0 2304 0 -1 756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5257_6
timestamp 1731220559
transform 1 0 2232 0 1 764
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5256_6
timestamp 1731220559
transform 1 0 2152 0 1 764
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5255_6
timestamp 1731220559
transform 1 0 2312 0 1 764
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5254_6
timestamp 1731220559
transform 1 0 2640 0 1 764
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5253_6
timestamp 1731220559
transform 1 0 2520 0 1 764
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5252_6
timestamp 1731220559
transform 1 0 2408 0 1 764
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5251_6
timestamp 1731220559
transform 1 0 2352 0 -1 928
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5250_6
timestamp 1731220559
transform 1 0 2272 0 -1 928
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5249_6
timestamp 1731220559
transform 1 0 2432 0 -1 928
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5248_6
timestamp 1731220559
transform 1 0 2512 0 -1 928
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5247_6
timestamp 1731220559
transform 1 0 2600 0 -1 928
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5246_6
timestamp 1731220559
transform 1 0 2696 0 -1 928
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5245_6
timestamp 1731220559
transform 1 0 2656 0 1 936
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5244_6
timestamp 1731220559
transform 1 0 2552 0 1 936
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5243_6
timestamp 1731220559
transform 1 0 2456 0 1 936
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5242_6
timestamp 1731220559
transform 1 0 2368 0 1 936
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5241_6
timestamp 1731220559
transform 1 0 2288 0 1 936
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5240_6
timestamp 1731220559
transform 1 0 2600 0 -1 1088
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5239_6
timestamp 1731220559
transform 1 0 2472 0 -1 1088
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5238_6
timestamp 1731220559
transform 1 0 2352 0 -1 1088
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5237_6
timestamp 1731220559
transform 1 0 2248 0 -1 1088
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5236_6
timestamp 1731220559
transform 1 0 2160 0 -1 1088
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5235_6
timestamp 1731220559
transform 1 0 2512 0 1 1096
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5234_6
timestamp 1731220559
transform 1 0 2352 0 1 1096
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5233_6
timestamp 1731220559
transform 1 0 2200 0 1 1096
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5232_6
timestamp 1731220559
transform 1 0 2072 0 1 1096
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5231_6
timestamp 1731220559
transform 1 0 1968 0 1 1096
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5230_6
timestamp 1731220559
transform 1 0 1888 0 1 1096
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5229_6
timestamp 1731220559
transform 1 0 1888 0 -1 1252
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5228_6
timestamp 1731220559
transform 1 0 1736 0 1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5227_6
timestamp 1731220559
transform 1 0 1736 0 -1 1280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5226_6
timestamp 1731220559
transform 1 0 2064 0 -1 1252
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5225_6
timestamp 1731220559
transform 1 0 2264 0 -1 1252
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5224_6
timestamp 1731220559
transform 1 0 2168 0 1 1260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5223_6
timestamp 1731220559
transform 1 0 2032 0 1 1260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5222_6
timestamp 1731220559
transform 1 0 1912 0 1 1260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5221_6
timestamp 1731220559
transform 1 0 2304 0 1 1260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5220_6
timestamp 1731220559
transform 1 0 2440 0 1 1260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5219_6
timestamp 1731220559
transform 1 0 2296 0 -1 1420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5218_6
timestamp 1731220559
transform 1 0 2160 0 -1 1420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5217_6
timestamp 1731220559
transform 1 0 2016 0 -1 1420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5216_6
timestamp 1731220559
transform 1 0 2256 0 1 1420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5215_6
timestamp 1731220559
transform 1 0 2400 0 1 1420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5214_6
timestamp 1731220559
transform 1 0 2360 0 -1 1580
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5213_6
timestamp 1731220559
transform 1 0 2520 0 -1 1580
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5212_6
timestamp 1731220559
transform 1 0 2480 0 1 1588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5211_6
timestamp 1731220559
transform 1 0 2624 0 1 1588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5210_6
timestamp 1731220559
transform 1 0 2520 0 -1 1744
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5209_6
timestamp 1731220559
transform 1 0 2656 0 -1 1744
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5208_6
timestamp 1731220559
transform 1 0 2704 0 1 1748
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5207_6
timestamp 1731220559
transform 1 0 2544 0 1 1748
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5206_6
timestamp 1731220559
transform 1 0 2232 0 -1 1916
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5205_6
timestamp 1731220559
transform 1 0 2304 0 1 1924
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5204_6
timestamp 1731220559
transform 1 0 2208 0 -1 2076
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5203_6
timestamp 1731220559
transform 1 0 2440 0 -1 2076
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5202_6
timestamp 1731220559
transform 1 0 2528 0 1 2084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5201_6
timestamp 1731220559
transform 1 0 2488 0 -1 2240
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5200_6
timestamp 1731220559
transform 1 0 2392 0 -1 2240
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5199_6
timestamp 1731220559
transform 1 0 2304 0 -1 2240
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5198_6
timestamp 1731220559
transform 1 0 2504 0 1 2240
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5197_6
timestamp 1731220559
transform 1 0 2424 0 1 2240
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5196_6
timestamp 1731220559
transform 1 0 2344 0 1 2240
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5195_6
timestamp 1731220559
transform 1 0 2264 0 1 2240
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5194_6
timestamp 1731220559
transform 1 0 2568 0 -1 2396
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5193_6
timestamp 1731220559
transform 1 0 2448 0 -1 2396
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5192_6
timestamp 1731220559
transform 1 0 2336 0 -1 2396
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5191_6
timestamp 1731220559
transform 1 0 2232 0 -1 2396
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5190_6
timestamp 1731220559
transform 1 0 2136 0 -1 2396
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5189_6
timestamp 1731220559
transform 1 0 2536 0 1 2400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5188_6
timestamp 1731220559
transform 1 0 2392 0 1 2400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5187_6
timestamp 1731220559
transform 1 0 2248 0 1 2400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5186_6
timestamp 1731220559
transform 1 0 2112 0 1 2400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5185_6
timestamp 1731220559
transform 1 0 1984 0 1 2400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5184_6
timestamp 1731220559
transform 1 0 2464 0 -1 2560
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5183_6
timestamp 1731220559
transform 1 0 2312 0 -1 2560
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5182_6
timestamp 1731220559
transform 1 0 2152 0 -1 2560
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5181_6
timestamp 1731220559
transform 1 0 2000 0 -1 2560
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5180_6
timestamp 1731220559
transform 1 0 1888 0 -1 2560
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5179_6
timestamp 1731220559
transform 1 0 2736 0 1 2560
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5178_6
timestamp 1731220559
transform 1 0 2480 0 1 2560
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5177_6
timestamp 1731220559
transform 1 0 2248 0 1 2560
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5176_6
timestamp 1731220559
transform 1 0 2040 0 1 2560
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5175_6
timestamp 1731220559
transform 1 0 1888 0 1 2560
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5174_6
timestamp 1731220559
transform 1 0 2528 0 -1 2720
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5173_6
timestamp 1731220559
transform 1 0 2320 0 -1 2720
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5172_6
timestamp 1731220559
transform 1 0 2312 0 1 2720
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5171_6
timestamp 1731220559
transform 1 0 2152 0 1 2720
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5170_6
timestamp 1731220559
transform 1 0 2128 0 -1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5169_6
timestamp 1731220559
transform 1 0 2040 0 -1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5168_6
timestamp 1731220559
transform 1 0 2112 0 1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5167_6
timestamp 1731220559
transform 1 0 2192 0 1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5166_6
timestamp 1731220559
transform 1 0 2192 0 -1 3048
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5165_6
timestamp 1731220559
transform 1 0 2472 0 -1 3048
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5164_6
timestamp 1731220559
transform 1 0 2328 0 -1 3048
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5163_6
timestamp 1731220559
transform 1 0 2248 0 1 3060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5162_6
timestamp 1731220559
transform 1 0 2056 0 1 3060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5161_6
timestamp 1731220559
transform 1 0 2440 0 1 3060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5160_6
timestamp 1731220559
transform 1 0 2448 0 -1 3212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5159_6
timestamp 1731220559
transform 1 0 2288 0 -1 3212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5158_6
timestamp 1731220559
transform 1 0 2304 0 1 3212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5157_6
timestamp 1731220559
transform 1 0 2432 0 1 3212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5156_6
timestamp 1731220559
transform 1 0 2432 0 -1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5155_6
timestamp 1731220559
transform 1 0 2576 0 -1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5154_6
timestamp 1731220559
transform 1 0 2664 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5153_6
timestamp 1731220559
transform 1 0 2520 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5152_6
timestamp 1731220559
transform 1 0 2376 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5151_6
timestamp 1731220559
transform 1 0 2328 0 -1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5150_6
timestamp 1731220559
transform 1 0 2504 0 -1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5149_6
timestamp 1731220559
transform 1 0 2544 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5148_6
timestamp 1731220559
transform 1 0 2408 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5147_6
timestamp 1731220559
transform 1 0 2280 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5146_6
timestamp 1731220559
transform 1 0 2144 0 -1 3668
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5145_6
timestamp 1731220559
transform 1 0 2160 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5144_6
timestamp 1731220559
transform 1 0 2056 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5143_6
timestamp 1731220559
transform 1 0 1968 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5142_6
timestamp 1731220559
transform 1 0 1888 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5141_6
timestamp 1731220559
transform 1 0 1960 0 -1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5140_6
timestamp 1731220559
transform 1 0 2144 0 -1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5139_6
timestamp 1731220559
transform 1 0 2112 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5138_6
timestamp 1731220559
transform 1 0 1992 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5137_6
timestamp 1731220559
transform 1 0 2240 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5136_6
timestamp 1731220559
transform 1 0 2288 0 -1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5135_6
timestamp 1731220559
transform 1 0 2144 0 -1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5134_6
timestamp 1731220559
transform 1 0 2008 0 -1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5133_6
timestamp 1731220559
transform 1 0 1912 0 1 3212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5132_6
timestamp 1731220559
transform 1 0 2048 0 1 3212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5131_6
timestamp 1731220559
transform 1 0 2176 0 1 3212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5130_6
timestamp 1731220559
transform 1 0 2136 0 -1 3212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5129_6
timestamp 1731220559
transform 1 0 2000 0 -1 3212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5128_6
timestamp 1731220559
transform 1 0 1888 0 -1 3212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5127_6
timestamp 1731220559
transform 1 0 1888 0 1 3060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5126_6
timestamp 1731220559
transform 1 0 1736 0 1 3084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5125_6
timestamp 1731220559
transform 1 0 1656 0 1 3084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5124_6
timestamp 1731220559
transform 1 0 1568 0 1 3084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5123_6
timestamp 1731220559
transform 1 0 1480 0 1 3084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5122_6
timestamp 1731220559
transform 1 0 1392 0 1 3084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5121_6
timestamp 1731220559
transform 1 0 1296 0 1 3084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5120_6
timestamp 1731220559
transform 1 0 1192 0 1 3084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5119_6
timestamp 1731220559
transform 1 0 1088 0 1 3084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5118_6
timestamp 1731220559
transform 1 0 976 0 1 3084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5117_6
timestamp 1731220559
transform 1 0 856 0 1 3084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5116_6
timestamp 1731220559
transform 1 0 1600 0 -1 3244
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5115_6
timestamp 1731220559
transform 1 0 1456 0 -1 3244
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5114_6
timestamp 1731220559
transform 1 0 1320 0 -1 3244
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5113_6
timestamp 1731220559
transform 1 0 1184 0 -1 3244
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5112_6
timestamp 1731220559
transform 1 0 1040 0 -1 3244
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5111_6
timestamp 1731220559
transform 1 0 1456 0 1 3244
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5110_6
timestamp 1731220559
transform 1 0 1328 0 1 3244
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5109_6
timestamp 1731220559
transform 1 0 1200 0 1 3244
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5108_6
timestamp 1731220559
transform 1 0 1072 0 1 3244
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5107_6
timestamp 1731220559
transform 1 0 936 0 1 3244
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5106_6
timestamp 1731220559
transform 1 0 1344 0 -1 3400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5105_6
timestamp 1731220559
transform 1 0 1232 0 -1 3400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5104_6
timestamp 1731220559
transform 1 0 1120 0 -1 3400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5103_6
timestamp 1731220559
transform 1 0 1008 0 -1 3400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5102_6
timestamp 1731220559
transform 1 0 888 0 -1 3400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5101_6
timestamp 1731220559
transform 1 0 1312 0 1 3404
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5100_6
timestamp 1731220559
transform 1 0 1216 0 1 3404
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_599_6
timestamp 1731220559
transform 1 0 1120 0 1 3404
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_598_6
timestamp 1731220559
transform 1 0 1024 0 1 3404
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_597_6
timestamp 1731220559
transform 1 0 928 0 1 3404
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_596_6
timestamp 1731220559
transform 1 0 1440 0 -1 3564
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_595_6
timestamp 1731220559
transform 1 0 1352 0 -1 3564
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_594_6
timestamp 1731220559
transform 1 0 1264 0 -1 3564
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_593_6
timestamp 1731220559
transform 1 0 1176 0 -1 3564
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_592_6
timestamp 1731220559
transform 1 0 1088 0 -1 3564
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_591_6
timestamp 1731220559
transform 1 0 1000 0 -1 3564
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_590_6
timestamp 1731220559
transform 1 0 1184 0 1 3564
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_589_6
timestamp 1731220559
transform 1 0 1040 0 1 3564
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_588_6
timestamp 1731220559
transform 1 0 896 0 1 3564
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_587_6
timestamp 1731220559
transform 1 0 760 0 1 3564
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_586_6
timestamp 1731220559
transform 1 0 912 0 -1 3564
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_585_6
timestamp 1731220559
transform 1 0 824 0 -1 3564
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_584_6
timestamp 1731220559
transform 1 0 728 0 -1 3564
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_583_6
timestamp 1731220559
transform 1 0 624 0 -1 3564
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_582_6
timestamp 1731220559
transform 1 0 520 0 -1 3564
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_581_6
timestamp 1731220559
transform 1 0 824 0 1 3404
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_580_6
timestamp 1731220559
transform 1 0 720 0 1 3404
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_579_6
timestamp 1731220559
transform 1 0 608 0 1 3404
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_578_6
timestamp 1731220559
transform 1 0 488 0 1 3404
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_577_6
timestamp 1731220559
transform 1 0 504 0 -1 3400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_576_6
timestamp 1731220559
transform 1 0 640 0 -1 3400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_575_6
timestamp 1731220559
transform 1 0 768 0 -1 3400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_574_6
timestamp 1731220559
transform 1 0 800 0 1 3244
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_573_6
timestamp 1731220559
transform 1 0 656 0 1 3244
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_572_6
timestamp 1731220559
transform 1 0 504 0 1 3244
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_571_6
timestamp 1731220559
transform 1 0 568 0 -1 3244
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_570_6
timestamp 1731220559
transform 1 0 728 0 -1 3244
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_569_6
timestamp 1731220559
transform 1 0 888 0 -1 3244
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_568_6
timestamp 1731220559
transform 1 0 728 0 1 3084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_567_6
timestamp 1731220559
transform 1 0 592 0 1 3084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_566_6
timestamp 1731220559
transform 1 0 448 0 1 3084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_565_6
timestamp 1731220559
transform 1 0 432 0 -1 3072
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_564_6
timestamp 1731220559
transform 1 0 544 0 -1 3072
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_563_6
timestamp 1731220559
transform 1 0 656 0 -1 3072
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_562_6
timestamp 1731220559
transform 1 0 784 0 1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_561_6
timestamp 1731220559
transform 1 0 632 0 1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_560_6
timestamp 1731220559
transform 1 0 472 0 1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_559_6
timestamp 1731220559
transform 1 0 464 0 -1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_558_6
timestamp 1731220559
transform 1 0 624 0 -1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_557_6
timestamp 1731220559
transform 1 0 776 0 -1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_556_6
timestamp 1731220559
transform 1 0 832 0 1 2752
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_555_6
timestamp 1731220559
transform 1 0 672 0 1 2752
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_554_6
timestamp 1731220559
transform 1 0 520 0 1 2752
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_553_6
timestamp 1731220559
transform 1 0 504 0 -1 2748
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_552_6
timestamp 1731220559
transform 1 0 656 0 -1 2748
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_551_6
timestamp 1731220559
transform 1 0 808 0 -1 2748
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_550_6
timestamp 1731220559
transform 1 0 776 0 1 2588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_549_6
timestamp 1731220559
transform 1 0 608 0 1 2588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_548_6
timestamp 1731220559
transform 1 0 520 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_547_6
timestamp 1731220559
transform 1 0 696 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_546_6
timestamp 1731220559
transform 1 0 872 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_545_6
timestamp 1731220559
transform 1 0 912 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_544_6
timestamp 1731220559
transform 1 0 768 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_543_6
timestamp 1731220559
transform 1 0 632 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_542_6
timestamp 1731220559
transform 1 0 496 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_541_6
timestamp 1731220559
transform 1 0 376 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_540_6
timestamp 1731220559
transform 1 0 288 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_539_6
timestamp 1731220559
transform 1 0 208 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_538_6
timestamp 1731220559
transform 1 0 128 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_537_6
timestamp 1731220559
transform 1 0 128 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_536_6
timestamp 1731220559
transform 1 0 216 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_535_6
timestamp 1731220559
transform 1 0 360 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_534_6
timestamp 1731220559
transform 1 0 432 0 1 2588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_533_6
timestamp 1731220559
transform 1 0 264 0 1 2588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_532_6
timestamp 1731220559
transform 1 0 128 0 1 2588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_531_6
timestamp 1731220559
transform 1 0 128 0 -1 2748
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_530_6
timestamp 1731220559
transform 1 0 224 0 -1 2748
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_529_6
timestamp 1731220559
transform 1 0 360 0 -1 2748
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_528_6
timestamp 1731220559
transform 1 0 368 0 1 2752
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_527_6
timestamp 1731220559
transform 1 0 232 0 1 2752
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_526_6
timestamp 1731220559
transform 1 0 128 0 1 2752
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_525_6
timestamp 1731220559
transform 1 0 144 0 -1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_524_6
timestamp 1731220559
transform 1 0 304 0 -1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_523_6
timestamp 1731220559
transform 1 0 304 0 1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_522_6
timestamp 1731220559
transform 1 0 144 0 1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_521_6
timestamp 1731220559
transform 1 0 128 0 -1 3072
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_520_6
timestamp 1731220559
transform 1 0 216 0 -1 3072
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_519_6
timestamp 1731220559
transform 1 0 320 0 -1 3072
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_518_6
timestamp 1731220559
transform 1 0 304 0 1 3084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_517_6
timestamp 1731220559
transform 1 0 160 0 1 3084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_516_6
timestamp 1731220559
transform 1 0 128 0 -1 3244
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_515_6
timestamp 1731220559
transform 1 0 408 0 -1 3244
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_514_6
timestamp 1731220559
transform 1 0 264 0 -1 3244
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_513_6
timestamp 1731220559
transform 1 0 192 0 1 3244
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_512_6
timestamp 1731220559
transform 1 0 352 0 1 3244
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_511_6
timestamp 1731220559
transform 1 0 360 0 -1 3400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_510_6
timestamp 1731220559
transform 1 0 208 0 -1 3400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_59_6
timestamp 1731220559
transform 1 0 216 0 1 3404
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_58_6
timestamp 1731220559
transform 1 0 352 0 1 3404
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_57_6
timestamp 1731220559
transform 1 0 296 0 -1 3564
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_56_6
timestamp 1731220559
transform 1 0 176 0 -1 3564
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_55_6
timestamp 1731220559
transform 1 0 408 0 -1 3564
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_54_6
timestamp 1731220559
transform 1 0 624 0 1 3564
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_53_6
timestamp 1731220559
transform 1 0 488 0 1 3564
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_52_6
timestamp 1731220559
transform 1 0 352 0 1 3564
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_51_6
timestamp 1731220559
transform 1 0 224 0 1 3564
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_50_6
timestamp 1731220559
transform 1 0 128 0 1 3564
box 8 4 70 72
<< end >>
