magic
tech sky130l
timestamp 1730254555
<< m1 >>
rect 8 72 12 76
rect 16 72 20 76
rect 24 72 28 76
rect 8 24 23 55
rect 8 4 12 8
<< labels >>
rlabel m1 s 8 72 12 76 6 in_50_6
port 1 nsew signal input
rlabel m1 s 8 4 12 8 6 out
port 2 nsew signal output
rlabel m1 s 16 72 20 76 6 Vdd
port 3 nsew power input
rlabel m1 s 24 72 28 76 6 GND
port 4 nsew ground input
<< properties >>
string LEFsite CoreSite
string LEFclass CORE
string FIXED_BBOX 0 0 32 80
string LEFsymmetry X Y
string LEFview TRUE
<< end >>
