magic
tech sky130l
timestamp 1729432489
<< ndiffusion >>
rect 8 10 13 12
rect 8 7 9 10
rect 12 7 13 10
rect 8 6 13 7
rect 15 10 20 12
rect 15 7 16 10
rect 19 7 20 10
rect 15 6 20 7
<< ndc >>
rect 9 7 12 10
rect 16 7 19 10
<< ntransistor >>
rect 13 6 15 12
<< pdiffusion >>
rect 8 28 13 29
rect 8 25 9 28
rect 12 25 13 28
rect 8 19 13 25
rect 15 28 20 29
rect 15 25 16 28
rect 19 25 20 28
rect 15 19 20 25
<< pdc >>
rect 9 25 12 28
rect 16 25 19 28
<< ptransistor >>
rect 13 19 15 29
<< polysilicon >>
rect 13 36 20 37
rect 13 33 16 36
rect 19 33 20 36
rect 13 32 20 33
rect 13 29 15 32
rect 13 12 15 19
rect 13 4 15 6
<< pc >>
rect 16 33 19 36
<< m1 >>
rect 16 36 20 37
rect 8 28 12 36
rect 8 25 9 28
rect 8 24 12 25
rect 19 33 20 36
rect 16 28 20 33
rect 19 25 20 28
rect 16 24 20 25
rect 8 10 12 11
rect 8 7 9 10
rect 8 4 12 7
rect 16 10 20 11
rect 19 7 20 10
rect 16 4 20 7
<< labels >>
rlabel ndiffusion 16 7 16 7 3 Y
rlabel pdiffusion 16 20 16 20 3 x
rlabel polysilicon 14 13 14 13 3 x
rlabel polysilicon 14 18 14 18 3 x
rlabel ndiffusion 9 7 9 7 3 GND
rlabel pdiffusion 9 20 9 20 3 Vdd
rlabel m1 9 33 9 33 3 Vdd
port 3 e
rlabel m1 9 5 9 5 2 GND
rlabel m1 19 5 19 5 8 Y
<< end >>
