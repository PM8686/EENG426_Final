magic
tech sky130l
timestamp 1731220617
<< m1 >>
rect 208 3619 212 3639
rect 296 3619 300 3639
rect 384 3619 388 3639
rect 472 3619 476 3639
rect 560 3619 564 3639
rect 648 3619 652 3639
rect 280 3511 284 3535
rect 456 3511 460 3535
rect 624 3511 628 3535
rect 928 3511 932 3535
rect 1064 3511 1068 3535
rect 1184 3511 1188 3535
rect 1304 3511 1308 3535
rect 1416 3511 1420 3535
rect 1520 3511 1524 3535
rect 1632 3511 1636 3535
rect 1720 3511 1724 3535
rect 240 3475 244 3495
rect 416 3475 420 3495
rect 584 3475 588 3495
rect 888 3475 892 3495
rect 1016 3475 1020 3495
rect 1272 3475 1276 3495
rect 1384 3475 1388 3495
rect 1600 3475 1604 3495
rect 1712 3475 1716 3495
rect 1808 3475 1812 3491
rect 1960 3471 1964 3491
rect 2056 3471 2060 3491
rect 2136 3471 2140 3491
rect 424 3375 428 3399
rect 632 3375 636 3399
rect 840 3375 844 3399
rect 1216 3375 1220 3399
rect 1392 3375 1396 3399
rect 1560 3375 1564 3399
rect 1720 3375 1724 3399
rect 2112 3371 2116 3395
rect 2248 3371 2252 3395
rect 2384 3371 2388 3395
rect 2648 3371 2652 3395
rect 2776 3371 2780 3395
rect 2912 3371 2916 3395
rect 3048 3371 3052 3395
rect 328 3331 332 3351
rect 472 3331 476 3351
rect 632 3331 636 3351
rect 800 3331 804 3351
rect 1096 3331 1100 3351
rect 1264 3331 1268 3351
rect 1416 3331 1420 3351
rect 1568 3331 1572 3351
rect 1960 3335 1964 3355
rect 2072 3335 2076 3355
rect 2216 3335 2220 3355
rect 2360 3335 2364 3355
rect 400 3227 404 3251
rect 1040 3227 1044 3251
rect 1184 3227 1188 3251
rect 1328 3227 1332 3251
rect 1480 3227 1484 3251
rect 2040 3235 2044 3259
rect 2168 3235 2172 3259
rect 2304 3235 2308 3259
rect 2448 3235 2452 3259
rect 2736 3235 2740 3259
rect 3024 3235 3028 3259
rect 3176 3235 3180 3259
rect 816 3179 820 3199
rect 968 3179 972 3199
rect 1104 3179 1108 3199
rect 1264 3179 1268 3199
rect 2072 3191 2076 3211
rect 2184 3191 2188 3211
rect 2312 3191 2316 3211
rect 2456 3191 2460 3211
rect 2744 3187 2748 3211
rect 2752 3131 2756 3211
rect 3192 3187 3196 3211
rect 256 3067 260 3091
rect 520 3067 524 3091
rect 640 3067 644 3091
rect 752 3067 756 3091
rect 960 3067 964 3091
rect 1064 3067 1068 3091
rect 1168 3067 1172 3091
rect 1264 3067 1268 3091
rect 2904 3087 2908 3171
rect 2912 3087 2916 3111
rect 3032 3087 3036 3111
rect 3264 3087 3268 3111
rect 3376 3087 3380 3111
rect 3472 3087 3476 3111
rect 664 3031 668 3051
rect 768 3031 772 3051
rect 864 3031 868 3051
rect 1056 3031 1060 3051
rect 2152 3047 2156 3067
rect 2296 3047 2300 3067
rect 2456 3047 2460 3067
rect 3048 3043 3052 3067
rect 3440 3047 3444 3067
rect 280 2919 284 2943
rect 776 2919 780 2943
rect 1184 2919 1188 2943
rect 1304 2919 1308 2943
rect 1712 2919 1716 2943
rect 2792 2935 2796 2959
rect 2896 2927 2900 2959
rect 3096 2935 3100 2959
rect 3192 2935 3196 2959
rect 3288 2935 3292 2959
rect 3384 2935 3388 2959
rect 3472 2915 3476 2959
rect 584 2883 588 2915
rect 624 2879 628 2903
rect 1480 2883 1484 2903
rect 1640 2883 1644 2903
rect 3056 2887 3060 2911
rect 648 2779 652 2803
rect 816 2779 820 2803
rect 1120 2779 1124 2803
rect 688 2735 692 2755
rect 696 2731 700 2763
rect 1264 2759 1268 2803
rect 1408 2779 1412 2803
rect 1552 2779 1556 2803
rect 1096 2735 1100 2755
rect 1360 2735 1364 2755
rect 1368 2731 1372 2763
rect 2744 2755 2748 2775
rect 2952 2755 2956 2775
rect 3064 2755 3068 2775
rect 3240 2755 3244 2775
rect 328 2631 332 2655
rect 456 2631 460 2655
rect 576 2631 580 2655
rect 928 2631 932 2655
rect 1040 2631 1044 2655
rect 1968 2655 1972 2679
rect 2144 2655 2148 2679
rect 2232 2655 2236 2679
rect 2320 2655 2324 2679
rect 2408 2655 2412 2679
rect 2496 2655 2500 2679
rect 2584 2655 2588 2679
rect 2672 2655 2676 2679
rect 2760 2655 2764 2679
rect 2848 2655 2852 2679
rect 2936 2655 2940 2679
rect 3024 2655 3028 2679
rect 3112 2655 3116 2679
rect 3200 2655 3204 2679
rect 3288 2655 3292 2679
rect 3384 2655 3388 2679
rect 1264 2631 1268 2655
rect 536 2591 540 2611
rect 624 2591 628 2611
rect 712 2591 716 2627
rect 888 2591 892 2611
rect 976 2591 980 2611
rect 1064 2591 1068 2611
rect 1240 2591 1244 2611
rect 1248 2587 1252 2619
rect 2224 2599 2228 2619
rect 2352 2599 2356 2619
rect 2488 2599 2492 2619
rect 2632 2599 2636 2619
rect 2928 2599 2932 2619
rect 752 2483 756 2507
rect 840 2483 844 2507
rect 1016 2483 1020 2507
rect 1104 2483 1108 2507
rect 1192 2483 1196 2507
rect 1280 2483 1284 2507
rect 2192 2499 2196 2523
rect 2304 2499 2308 2523
rect 2424 2499 2428 2523
rect 2552 2499 2556 2523
rect 424 2443 428 2463
rect 664 2439 668 2463
rect 1032 2443 1036 2463
rect 1280 2443 1284 2463
rect 1408 2443 1412 2463
rect 2152 2459 2156 2479
rect 2248 2459 2252 2479
rect 2352 2459 2356 2479
rect 2360 2455 2364 2487
rect 3472 2483 3476 2523
rect 2632 2459 2636 2479
rect 2776 2459 2780 2479
rect 2992 2459 2996 2479
rect 280 2323 284 2363
rect 1200 2339 1204 2363
rect 1368 2339 1372 2363
rect 1536 2339 1540 2363
rect 1704 2339 1708 2363
rect 2056 2355 2060 2379
rect 2176 2355 2180 2379
rect 2304 2355 2308 2379
rect 2440 2355 2444 2379
rect 2744 2355 2748 2379
rect 2920 2355 2924 2379
rect 3104 2355 3108 2379
rect 584 2299 588 2319
rect 776 2299 780 2319
rect 1504 2295 1508 2319
rect 1960 2311 1964 2331
rect 2088 2311 2092 2331
rect 2240 2311 2244 2331
rect 2392 2311 2396 2331
rect 2744 2311 2748 2331
rect 3032 2311 3036 2331
rect 3208 2311 3212 2331
rect 3360 2251 3364 2351
rect 3472 2335 3476 2379
rect 248 2191 252 2215
rect 400 2191 404 2215
rect 1008 2191 1012 2215
rect 1448 2191 1452 2215
rect 2016 2207 2020 2231
rect 2192 2207 2196 2231
rect 2376 2207 2380 2231
rect 2560 2207 2564 2231
rect 2904 2207 2908 2231
rect 3072 2207 3076 2231
rect 3232 2207 3236 2231
rect 280 2151 284 2171
rect 480 2151 484 2171
rect 584 2151 588 2171
rect 688 2151 692 2187
rect 792 2151 796 2171
rect 1120 2151 1124 2171
rect 1128 2147 1132 2179
rect 1880 2107 1884 2187
rect 1960 2167 1964 2187
rect 2136 2167 2140 2187
rect 2312 2167 2316 2187
rect 2496 2167 2500 2187
rect 2856 2167 2860 2187
rect 3000 2167 3004 2187
rect 3152 2167 3156 2187
rect 3296 2167 3300 2187
rect 408 2023 412 2083
rect 416 2043 420 2067
rect 600 2043 604 2067
rect 704 2043 708 2067
rect 920 2043 924 2067
rect 1024 2043 1028 2067
rect 1128 2043 1132 2067
rect 2368 2063 2372 2087
rect 2544 2063 2548 2087
rect 3032 2019 3036 2039
rect 288 1995 292 2019
rect 1216 1999 1220 2019
rect 512 1891 516 1915
rect 1256 1891 1260 1915
rect 1416 1891 1420 1915
rect 1576 1891 1580 1915
rect 2104 1915 2108 1939
rect 2192 1915 2196 1939
rect 2280 1915 2284 1939
rect 2376 1915 2380 1939
rect 1720 1891 1724 1915
rect 3472 1895 3476 1939
rect 2512 1867 2516 1891
rect 2712 1871 2716 1891
rect 3032 1871 3036 1891
rect 3224 1871 3228 1891
rect 616 1847 620 1867
rect 800 1847 804 1867
rect 1144 1847 1148 1867
rect 1480 1843 1484 1867
rect 1640 1843 1644 1867
rect 2432 1767 2436 1791
rect 2912 1767 2916 1791
rect 3040 1767 3044 1791
rect 3176 1767 3180 1791
rect 3312 1767 3316 1791
rect 256 1739 260 1763
rect 560 1739 564 1763
rect 712 1739 716 1763
rect 1416 1739 1420 1763
rect 2360 1723 2364 1743
rect 568 1647 572 1723
rect 800 1703 804 1723
rect 936 1703 940 1723
rect 1064 1703 1068 1723
rect 1248 1703 1252 1723
rect 2472 1723 2476 1743
rect 2600 1723 2604 1743
rect 3200 1723 3204 1743
rect 3328 1719 3332 1751
rect 256 1603 260 1627
rect 568 1603 572 1627
rect 1000 1603 1004 1627
rect 1272 1603 1276 1627
rect 1408 1603 1412 1627
rect 2240 1619 2244 1643
rect 2360 1619 2364 1643
rect 2496 1619 2500 1643
rect 2640 1619 2644 1643
rect 3472 1607 3476 1643
rect 2072 1583 2076 1603
rect 248 1563 252 1583
rect 600 1563 604 1583
rect 1080 1563 1084 1583
rect 1232 1563 1236 1583
rect 1376 1563 1380 1583
rect 1520 1563 1524 1583
rect 2168 1583 2172 1603
rect 2272 1583 2276 1603
rect 2400 1583 2404 1603
rect 2696 1579 2700 1603
rect 2848 1579 2852 1603
rect 3200 1579 3204 1603
rect 752 1459 756 1483
rect 928 1459 932 1483
rect 1248 1459 1252 1483
rect 1400 1459 1404 1483
rect 1552 1459 1556 1483
rect 1704 1459 1708 1483
rect 1968 1475 1972 1499
rect 2232 1475 2236 1499
rect 2376 1475 2380 1499
rect 2480 1459 2484 1499
rect 3048 1475 3052 1499
rect 456 1419 460 1439
rect 760 1419 764 1439
rect 1080 1415 1084 1439
rect 1376 1419 1380 1439
rect 1528 1419 1532 1439
rect 1808 1419 1812 1455
rect 1960 1435 1964 1455
rect 2104 1435 2108 1455
rect 2696 1435 2700 1455
rect 3200 1435 3204 1455
rect 3208 1431 3212 1463
rect 3264 1367 3268 1471
rect 432 1319 436 1343
rect 696 1319 700 1343
rect 1120 1319 1124 1343
rect 1272 1319 1276 1343
rect 1584 1319 1588 1343
rect 1720 1307 1724 1343
rect 2384 1311 2388 1347
rect 3056 1323 3060 1347
rect 3472 1311 3476 1347
rect 520 1283 524 1303
rect 608 1283 612 1303
rect 696 1283 700 1303
rect 784 1283 788 1303
rect 2208 1283 2212 1307
rect 3056 1287 3060 1307
rect 3232 1287 3236 1307
rect 624 1183 628 1207
rect 712 1163 716 1207
rect 888 1183 892 1207
rect 1088 1183 1092 1207
rect 1200 1183 1204 1207
rect 1328 1183 1332 1207
rect 1464 1183 1468 1207
rect 1720 1183 1724 1207
rect 2472 1167 2476 1203
rect 3472 1167 3476 1203
rect 424 1139 428 1159
rect 536 1139 540 1159
rect 1368 1139 1372 1159
rect 1376 1135 1380 1167
rect 1960 1143 1964 1163
rect 2080 1143 2084 1163
rect 2888 1143 2892 1163
rect 3232 1143 3236 1163
rect 280 1035 284 1059
rect 440 1035 444 1059
rect 776 1035 780 1059
rect 1096 1035 1100 1059
rect 1552 1035 1556 1059
rect 256 995 260 1015
rect 576 995 580 1015
rect 760 995 764 1015
rect 1128 995 1132 1015
rect 1296 995 1300 1015
rect 2168 995 2172 1015
rect 2296 995 2300 1015
rect 2704 995 2708 1031
rect 2904 995 2908 1015
rect 3056 995 3060 1015
rect 3232 995 3236 1015
rect 128 875 132 915
rect 456 891 460 975
rect 656 891 660 915
rect 848 891 852 915
rect 1216 891 1220 915
rect 1392 891 1396 915
rect 1568 891 1572 915
rect 1720 891 1724 915
rect 2120 875 2124 915
rect 224 851 228 871
rect 456 851 460 871
rect 568 851 572 871
rect 752 851 756 871
rect 1096 851 1100 871
rect 1280 851 1284 871
rect 1448 851 1452 871
rect 1616 851 1620 871
rect 2168 851 2172 871
rect 2256 851 2260 871
rect 2432 851 2436 871
rect 2552 851 2556 887
rect 2640 851 2644 871
rect 2776 851 2780 871
rect 2968 851 2972 871
rect 3160 851 3164 871
rect 264 751 268 775
rect 416 751 420 775
rect 576 751 580 775
rect 736 751 740 775
rect 1032 751 1036 775
rect 1176 751 1180 775
rect 1320 751 1324 775
rect 1472 751 1476 775
rect 2368 751 2372 775
rect 2776 751 2780 775
rect 2928 751 2932 775
rect 3104 751 3108 775
rect 3288 751 3292 775
rect 424 711 428 731
rect 512 711 516 731
rect 608 711 612 731
rect 704 711 708 731
rect 896 711 900 731
rect 992 711 996 731
rect 1096 711 1100 731
rect 1224 711 1228 731
rect 2336 711 2340 731
rect 2488 711 2492 731
rect 2768 711 2772 731
rect 2920 711 2924 731
rect 3064 711 3068 731
rect 560 607 564 631
rect 648 607 652 631
rect 736 607 740 631
rect 824 607 828 631
rect 912 595 916 631
rect 1176 607 1180 631
rect 2016 607 2020 631
rect 2192 607 2196 631
rect 3056 607 3060 631
rect 3344 607 3348 631
rect 568 571 572 591
rect 664 571 668 591
rect 1128 571 1132 591
rect 1264 571 1268 591
rect 1408 571 1412 591
rect 1416 567 1420 603
rect 2280 507 2284 591
rect 2416 571 2420 591
rect 2576 571 2580 603
rect 3472 595 3476 631
rect 2776 571 2780 591
rect 3128 571 3132 591
rect 1360 471 1364 495
rect 1696 471 1700 495
rect 2280 463 2284 487
rect 2840 463 2844 487
rect 3008 463 3012 487
rect 3168 451 3172 487
rect 216 427 220 447
rect 536 427 540 447
rect 712 427 716 447
rect 944 371 948 447
rect 1056 427 1060 447
rect 1272 427 1276 447
rect 1536 427 1540 447
rect 2312 427 2316 447
rect 2400 427 2404 447
rect 2496 427 2500 447
rect 2800 427 2804 447
rect 3256 427 3260 447
rect 3264 423 3268 439
rect 3472 371 3476 447
rect 256 327 260 351
rect 424 327 428 351
rect 600 327 604 351
rect 776 327 780 351
rect 1424 327 1428 351
rect 1584 327 1588 351
rect 2232 327 2236 351
rect 2320 327 2324 351
rect 2408 327 2412 351
rect 2496 327 2500 351
rect 3096 327 3100 351
rect 3296 327 3300 351
rect 464 287 468 307
rect 608 287 612 307
rect 768 287 772 307
rect 984 227 988 307
rect 1088 287 1092 307
rect 1608 283 1612 307
rect 2088 291 2092 311
rect 2184 291 2188 311
rect 2288 291 2292 311
rect 2600 291 2604 311
rect 2704 291 2708 311
rect 2808 291 2812 311
rect 2920 291 2924 311
rect 3472 235 3476 323
rect 496 183 500 207
rect 608 183 612 207
rect 728 183 732 207
rect 856 183 860 207
rect 1488 183 1492 207
rect 1616 183 1620 207
rect 1720 183 1724 207
rect 2760 191 2764 215
rect 2944 191 2948 215
rect 3120 191 3124 215
rect 3304 191 3308 215
rect 288 127 292 147
rect 376 127 380 147
rect 464 127 468 147
rect 552 127 556 147
rect 640 127 644 147
rect 728 127 732 147
rect 816 127 820 147
rect 904 127 908 147
rect 992 127 996 147
rect 1080 127 1084 147
rect 1256 127 1260 147
rect 1360 127 1364 147
rect 1464 127 1468 147
rect 1576 127 1580 147
rect 1584 123 1588 171
rect 1808 127 1812 143
rect 1960 123 1964 143
rect 2056 123 2060 143
rect 2136 123 2140 143
rect 2224 123 2228 143
rect 2336 123 2340 143
rect 2672 123 2676 143
rect 2784 123 2788 143
rect 2912 123 2916 143
rect 2992 123 2996 143
rect 3088 123 3092 143
rect 3184 123 3188 143
rect 3280 123 3284 143
rect 3376 123 3380 143
rect 3464 123 3468 143
<< m2c >>
rect 208 3639 212 3643
rect 240 3639 244 3643
rect 296 3639 300 3643
rect 328 3639 332 3643
rect 384 3639 388 3643
rect 416 3639 420 3643
rect 472 3639 476 3643
rect 504 3639 508 3643
rect 560 3639 564 3643
rect 592 3639 596 3643
rect 648 3639 652 3643
rect 680 3639 684 3643
rect 208 3615 212 3619
rect 296 3615 300 3619
rect 384 3615 388 3619
rect 472 3615 476 3619
rect 560 3615 564 3619
rect 648 3615 652 3619
rect 280 3535 284 3539
rect 456 3535 460 3539
rect 624 3535 628 3539
rect 928 3535 932 3539
rect 152 3507 156 3511
rect 280 3507 284 3511
rect 304 3507 308 3511
rect 456 3507 460 3511
rect 480 3507 484 3511
rect 624 3507 628 3511
rect 648 3507 652 3511
rect 808 3509 812 3513
rect 1064 3535 1068 3539
rect 1184 3535 1188 3539
rect 1304 3535 1308 3539
rect 1416 3535 1420 3539
rect 1520 3535 1524 3539
rect 1632 3535 1636 3539
rect 1720 3535 1724 3539
rect 928 3507 932 3511
rect 952 3507 956 3511
rect 1064 3507 1068 3511
rect 1088 3507 1092 3511
rect 1184 3507 1188 3511
rect 1208 3507 1212 3511
rect 1304 3507 1308 3511
rect 1328 3507 1332 3511
rect 1416 3507 1420 3511
rect 1440 3507 1444 3511
rect 1520 3507 1524 3511
rect 1544 3507 1548 3511
rect 1632 3507 1636 3511
rect 1656 3507 1660 3511
rect 1720 3507 1724 3511
rect 1744 3507 1748 3511
rect 160 3495 164 3499
rect 240 3495 244 3499
rect 336 3495 340 3499
rect 416 3495 420 3499
rect 504 3495 508 3499
rect 584 3495 588 3499
rect 664 3495 668 3499
rect 816 3495 820 3499
rect 888 3495 892 3499
rect 960 3495 964 3499
rect 1016 3495 1020 3499
rect 1096 3495 1100 3499
rect 1216 3495 1220 3499
rect 1272 3495 1276 3499
rect 1328 3495 1332 3499
rect 1384 3495 1388 3499
rect 1440 3495 1444 3499
rect 1544 3495 1548 3499
rect 1600 3495 1604 3499
rect 1656 3495 1660 3499
rect 1712 3495 1716 3499
rect 1744 3495 1748 3499
rect 240 3471 244 3475
rect 416 3471 420 3475
rect 584 3471 588 3475
rect 888 3471 892 3475
rect 1016 3471 1020 3475
rect 1272 3471 1276 3475
rect 1384 3471 1388 3475
rect 1600 3471 1604 3475
rect 1712 3471 1716 3475
rect 1808 3491 1812 3495
rect 1904 3491 1908 3495
rect 1960 3491 1964 3495
rect 1992 3491 1996 3495
rect 2056 3491 2060 3495
rect 2080 3491 2084 3495
rect 2136 3491 2140 3495
rect 2168 3491 2172 3495
rect 1808 3471 1812 3475
rect 1960 3467 1964 3471
rect 2056 3467 2060 3471
rect 2136 3467 2140 3471
rect 424 3399 428 3403
rect 632 3399 636 3403
rect 840 3399 844 3403
rect 1216 3399 1220 3403
rect 1392 3399 1396 3403
rect 1560 3399 1564 3403
rect 1720 3399 1724 3403
rect 2112 3395 2116 3399
rect 232 3371 236 3375
rect 424 3371 428 3375
rect 448 3371 452 3375
rect 632 3371 636 3375
rect 656 3371 660 3375
rect 840 3371 844 3375
rect 864 3371 868 3375
rect 1056 3371 1060 3375
rect 1216 3371 1220 3375
rect 1240 3371 1244 3375
rect 1392 3371 1396 3375
rect 1416 3371 1420 3375
rect 1560 3371 1564 3375
rect 1584 3371 1588 3375
rect 1720 3371 1724 3375
rect 1744 3371 1748 3375
rect 2248 3395 2252 3399
rect 2384 3395 2388 3399
rect 2648 3395 2652 3399
rect 2776 3395 2780 3399
rect 2912 3395 2916 3399
rect 3048 3395 3052 3399
rect 1904 3367 1908 3371
rect 2008 3367 2012 3371
rect 2112 3367 2116 3371
rect 2136 3367 2140 3371
rect 2248 3367 2252 3371
rect 2272 3367 2276 3371
rect 2384 3367 2388 3371
rect 2408 3367 2412 3371
rect 2544 3367 2548 3371
rect 2648 3367 2652 3371
rect 2672 3367 2676 3371
rect 2776 3367 2780 3371
rect 2800 3367 2804 3371
rect 2912 3367 2916 3371
rect 2936 3367 2940 3371
rect 3048 3367 3052 3371
rect 3072 3367 3076 3371
rect 1904 3355 1908 3359
rect 1960 3355 1964 3359
rect 2008 3355 2012 3359
rect 2072 3355 2076 3359
rect 2144 3355 2148 3359
rect 2216 3355 2220 3359
rect 2288 3355 2292 3359
rect 2360 3355 2364 3359
rect 2432 3355 2436 3359
rect 2568 3355 2572 3359
rect 2704 3355 2708 3359
rect 2840 3355 2844 3359
rect 2976 3355 2980 3359
rect 3112 3355 3116 3359
rect 248 3351 252 3355
rect 328 3351 332 3355
rect 392 3351 396 3355
rect 472 3351 476 3355
rect 552 3351 556 3355
rect 632 3351 636 3355
rect 720 3351 724 3355
rect 800 3351 804 3355
rect 880 3351 884 3355
rect 1040 3351 1044 3355
rect 1096 3351 1100 3355
rect 1192 3351 1196 3355
rect 1264 3351 1268 3355
rect 1344 3351 1348 3355
rect 1416 3351 1420 3355
rect 1496 3351 1500 3355
rect 1568 3351 1572 3355
rect 1648 3351 1652 3355
rect 328 3327 332 3331
rect 472 3327 476 3331
rect 632 3327 636 3331
rect 800 3327 804 3331
rect 1096 3327 1100 3331
rect 1264 3327 1268 3331
rect 1416 3327 1420 3331
rect 1960 3331 1964 3335
rect 2072 3331 2076 3335
rect 2216 3331 2220 3335
rect 2360 3331 2364 3335
rect 1568 3327 1572 3331
rect 2040 3259 2044 3263
rect 400 3251 404 3255
rect 1040 3251 1044 3255
rect 1184 3251 1188 3255
rect 1328 3251 1332 3255
rect 1480 3251 1484 3255
rect 2168 3259 2172 3263
rect 2304 3259 2308 3263
rect 2448 3259 2452 3263
rect 2736 3259 2740 3263
rect 3024 3259 3028 3263
rect 3176 3259 3180 3263
rect 1944 3231 1948 3235
rect 2040 3231 2044 3235
rect 2064 3231 2068 3235
rect 2168 3231 2172 3235
rect 2192 3231 2196 3235
rect 2304 3231 2308 3235
rect 2328 3231 2332 3235
rect 2448 3231 2452 3235
rect 2472 3231 2476 3235
rect 2616 3231 2620 3235
rect 2736 3231 2740 3235
rect 2760 3231 2764 3235
rect 2904 3231 2908 3235
rect 3024 3231 3028 3235
rect 3048 3231 3052 3235
rect 3176 3231 3180 3235
rect 3200 3231 3204 3235
rect 256 3223 260 3227
rect 400 3223 404 3227
rect 424 3223 428 3227
rect 592 3223 596 3227
rect 760 3223 764 3227
rect 912 3223 916 3227
rect 1040 3223 1044 3227
rect 1064 3223 1068 3227
rect 1184 3223 1188 3227
rect 1208 3223 1212 3227
rect 1328 3223 1332 3227
rect 1352 3223 1356 3227
rect 1480 3223 1484 3227
rect 1504 3223 1508 3227
rect 2016 3211 2020 3215
rect 2072 3211 2076 3215
rect 2128 3211 2132 3215
rect 2184 3211 2188 3215
rect 2248 3211 2252 3215
rect 2312 3211 2316 3215
rect 2384 3211 2388 3215
rect 2456 3211 2460 3215
rect 2528 3211 2532 3215
rect 2672 3211 2676 3215
rect 2744 3211 2748 3215
rect 184 3199 188 3203
rect 384 3199 388 3203
rect 568 3199 572 3203
rect 736 3199 740 3203
rect 816 3199 820 3203
rect 896 3199 900 3203
rect 968 3199 972 3203
rect 1048 3199 1052 3203
rect 1104 3199 1108 3203
rect 1200 3199 1204 3203
rect 1264 3199 1268 3203
rect 1360 3199 1364 3203
rect 816 3175 820 3179
rect 968 3175 972 3179
rect 1104 3175 1108 3179
rect 2072 3187 2076 3191
rect 2184 3187 2188 3191
rect 2312 3187 2316 3191
rect 2456 3187 2460 3191
rect 2744 3183 2748 3187
rect 2752 3211 2756 3215
rect 2824 3211 2828 3215
rect 2976 3211 2980 3215
rect 3128 3211 3132 3215
rect 3192 3211 3196 3215
rect 3288 3211 3292 3215
rect 1264 3175 1268 3179
rect 2560 3155 2564 3159
rect 3192 3183 3196 3187
rect 2752 3127 2756 3131
rect 2904 3171 2908 3175
rect 256 3091 260 3095
rect 520 3091 524 3095
rect 640 3091 644 3095
rect 752 3091 756 3095
rect 960 3091 964 3095
rect 1064 3091 1068 3095
rect 1168 3091 1172 3095
rect 1264 3091 1268 3095
rect 2072 3083 2076 3087
rect 2224 3083 2228 3087
rect 2376 3083 2380 3087
rect 2528 3083 2532 3087
rect 2672 3083 2676 3087
rect 2808 3083 2812 3087
rect 2904 3083 2908 3087
rect 2912 3111 2916 3115
rect 3032 3111 3036 3115
rect 3264 3111 3268 3115
rect 3376 3111 3380 3115
rect 3472 3111 3476 3115
rect 2912 3083 2916 3087
rect 2936 3083 2940 3087
rect 3032 3083 3036 3087
rect 3056 3083 3060 3087
rect 3176 3083 3180 3087
rect 3264 3083 3268 3087
rect 3288 3083 3292 3087
rect 3376 3083 3380 3087
rect 3400 3083 3404 3087
rect 3472 3083 3476 3087
rect 3496 3083 3500 3087
rect 1960 3067 1964 3071
rect 2088 3067 2092 3071
rect 2152 3067 2156 3071
rect 2224 3067 2228 3071
rect 2296 3067 2300 3071
rect 2376 3067 2380 3071
rect 2456 3067 2460 3071
rect 2536 3067 2540 3071
rect 2688 3067 2692 3071
rect 2840 3067 2844 3071
rect 2984 3067 2988 3071
rect 3048 3067 3052 3071
rect 3120 3067 3124 3071
rect 3248 3067 3252 3071
rect 3384 3067 3388 3071
rect 3440 3067 3444 3071
rect 3496 3067 3500 3071
rect 152 3063 156 3067
rect 256 3063 260 3067
rect 280 3063 284 3067
rect 416 3063 420 3067
rect 520 3063 524 3067
rect 544 3063 548 3067
rect 640 3063 644 3067
rect 664 3063 668 3067
rect 752 3063 756 3067
rect 776 3063 780 3067
rect 880 3063 884 3067
rect 960 3063 964 3067
rect 984 3063 988 3067
rect 1064 3063 1068 3067
rect 1088 3063 1092 3067
rect 1168 3063 1172 3067
rect 1192 3063 1196 3067
rect 1264 3063 1268 3067
rect 1296 3063 1300 3067
rect 152 3051 156 3055
rect 256 3051 260 3055
rect 376 3051 380 3055
rect 496 3051 500 3055
rect 608 3051 612 3055
rect 664 3051 668 3055
rect 712 3051 716 3055
rect 768 3051 772 3055
rect 808 3051 812 3055
rect 864 3051 868 3055
rect 904 3051 908 3055
rect 1000 3051 1004 3055
rect 1056 3051 1060 3055
rect 1096 3051 1100 3055
rect 1192 3051 1196 3055
rect 1296 3051 1300 3055
rect 664 3027 668 3031
rect 768 3027 772 3031
rect 864 3027 868 3031
rect 2152 3043 2156 3047
rect 2296 3043 2300 3047
rect 2456 3043 2460 3047
rect 3440 3043 3444 3047
rect 3048 3039 3052 3043
rect 1056 3027 1060 3031
rect 3528 3011 3532 3015
rect 184 2995 188 2999
rect 936 2995 940 2999
rect 2792 2959 2796 2963
rect 280 2943 284 2947
rect 776 2943 780 2947
rect 1184 2943 1188 2947
rect 1304 2943 1308 2947
rect 1712 2943 1716 2947
rect 2896 2959 2900 2963
rect 1904 2931 1908 2935
rect 1992 2931 1996 2935
rect 2080 2931 2084 2935
rect 2168 2931 2172 2935
rect 2256 2931 2260 2935
rect 2368 2931 2372 2935
rect 2480 2931 2484 2935
rect 2592 2931 2596 2935
rect 2704 2931 2708 2935
rect 2792 2931 2796 2935
rect 2816 2931 2820 2935
rect 3096 2959 3100 2963
rect 3192 2959 3196 2963
rect 3288 2959 3292 2963
rect 3384 2959 3388 2963
rect 3472 2959 3476 2963
rect 2920 2931 2924 2935
rect 3024 2931 3028 2935
rect 3096 2931 3100 2935
rect 3120 2931 3124 2935
rect 3192 2931 3196 2935
rect 3216 2931 3220 2935
rect 3288 2931 3292 2935
rect 3312 2931 3316 2935
rect 3384 2931 3388 2935
rect 3408 2931 3412 2935
rect 2896 2923 2900 2927
rect 152 2915 156 2919
rect 280 2915 284 2919
rect 304 2915 308 2919
rect 472 2915 476 2919
rect 584 2915 588 2919
rect 640 2915 644 2919
rect 776 2915 780 2919
rect 800 2915 804 2919
rect 944 2915 948 2919
rect 1080 2915 1084 2919
rect 1184 2915 1188 2919
rect 1208 2915 1212 2919
rect 1304 2915 1308 2919
rect 1328 2915 1332 2919
rect 1440 2915 1444 2919
rect 1544 2915 1548 2919
rect 1656 2915 1660 2919
rect 1712 2915 1716 2919
rect 1744 2915 1748 2919
rect 3496 2931 3500 2935
rect 152 2903 156 2907
rect 328 2903 332 2907
rect 528 2903 532 2907
rect 2904 2911 2908 2915
rect 3056 2911 3060 2915
rect 3208 2911 3212 2915
rect 3472 2911 3476 2915
rect 3496 2911 3500 2915
rect 584 2879 588 2883
rect 624 2903 628 2907
rect 720 2903 724 2907
rect 904 2903 908 2907
rect 1080 2903 1084 2907
rect 1248 2903 1252 2907
rect 1408 2903 1412 2907
rect 1480 2903 1484 2907
rect 1560 2903 1564 2907
rect 1640 2903 1644 2907
rect 1720 2903 1724 2907
rect 1480 2879 1484 2883
rect 3056 2883 3060 2887
rect 1640 2879 1644 2883
rect 624 2875 628 2879
rect 3528 2855 3532 2859
rect 184 2847 188 2851
rect 1280 2847 1284 2851
rect 648 2803 652 2807
rect 816 2803 820 2807
rect 1120 2803 1124 2807
rect 1264 2803 1268 2807
rect 176 2775 180 2779
rect 336 2775 340 2779
rect 504 2775 508 2779
rect 648 2775 652 2779
rect 672 2775 676 2779
rect 816 2775 820 2779
rect 840 2775 844 2779
rect 992 2775 996 2779
rect 1120 2775 1124 2779
rect 1144 2775 1148 2779
rect 696 2763 700 2767
rect 216 2755 220 2759
rect 344 2755 348 2759
rect 480 2755 484 2759
rect 616 2755 620 2759
rect 688 2755 692 2759
rect 688 2731 692 2735
rect 1408 2803 1412 2807
rect 1552 2803 1556 2807
rect 2848 2787 2852 2791
rect 2936 2787 2940 2791
rect 3024 2787 3028 2791
rect 3112 2787 3116 2791
rect 1288 2775 1292 2779
rect 1408 2775 1412 2779
rect 1432 2775 1436 2779
rect 1552 2775 1556 2779
rect 1576 2775 1580 2779
rect 2680 2775 2684 2779
rect 2744 2775 2748 2779
rect 2816 2775 2820 2779
rect 2952 2775 2956 2779
rect 2976 2775 2980 2779
rect 3064 2775 3068 2779
rect 3152 2775 3156 2779
rect 3240 2775 3244 2779
rect 3336 2775 3340 2779
rect 3496 2775 3500 2779
rect 1368 2763 1372 2767
rect 760 2755 764 2759
rect 896 2755 900 2759
rect 1032 2755 1036 2759
rect 1096 2755 1100 2759
rect 1160 2755 1164 2759
rect 1264 2755 1268 2759
rect 1296 2755 1300 2759
rect 1360 2755 1364 2759
rect 1096 2731 1100 2735
rect 1360 2731 1364 2735
rect 1432 2755 1436 2759
rect 2744 2751 2748 2755
rect 2952 2751 2956 2755
rect 3064 2751 3068 2755
rect 3240 2751 3244 2755
rect 696 2727 700 2731
rect 1368 2727 1372 2731
rect 3528 2719 3532 2723
rect 248 2699 252 2703
rect 1192 2699 1196 2703
rect 1968 2679 1972 2683
rect 328 2655 332 2659
rect 456 2655 460 2659
rect 576 2655 580 2659
rect 928 2655 932 2659
rect 1040 2655 1044 2659
rect 1264 2655 1268 2659
rect 2144 2679 2148 2683
rect 2232 2679 2236 2683
rect 2320 2679 2324 2683
rect 2408 2679 2412 2683
rect 2496 2679 2500 2683
rect 2584 2679 2588 2683
rect 2672 2679 2676 2683
rect 2760 2679 2764 2683
rect 2848 2679 2852 2683
rect 2936 2679 2940 2683
rect 3024 2679 3028 2683
rect 3112 2679 3116 2683
rect 3200 2679 3204 2683
rect 3288 2679 3292 2683
rect 3384 2679 3388 2683
rect 1904 2651 1908 2655
rect 1968 2651 1972 2655
rect 1992 2651 1996 2655
rect 2080 2651 2084 2655
rect 2144 2651 2148 2655
rect 2168 2651 2172 2655
rect 2232 2651 2236 2655
rect 2256 2651 2260 2655
rect 2320 2651 2324 2655
rect 2344 2651 2348 2655
rect 2408 2651 2412 2655
rect 2432 2651 2436 2655
rect 2496 2651 2500 2655
rect 2520 2651 2524 2655
rect 2584 2651 2588 2655
rect 2608 2651 2612 2655
rect 2672 2651 2676 2655
rect 2696 2651 2700 2655
rect 2760 2651 2764 2655
rect 2784 2651 2788 2655
rect 2848 2651 2852 2655
rect 2872 2651 2876 2655
rect 2936 2651 2940 2655
rect 2960 2651 2964 2655
rect 3024 2651 3028 2655
rect 3048 2651 3052 2655
rect 3112 2651 3116 2655
rect 3136 2651 3140 2655
rect 3200 2651 3204 2655
rect 3224 2651 3228 2655
rect 3288 2651 3292 2655
rect 3312 2651 3316 2655
rect 3384 2651 3388 2655
rect 3408 2651 3412 2655
rect 3496 2651 3500 2655
rect 232 2627 236 2631
rect 328 2627 332 2631
rect 352 2627 356 2631
rect 456 2627 460 2631
rect 480 2627 484 2631
rect 576 2627 580 2631
rect 600 2627 604 2631
rect 712 2627 716 2631
rect 720 2627 724 2631
rect 840 2627 844 2631
rect 928 2627 932 2631
rect 952 2627 956 2631
rect 1040 2627 1044 2631
rect 1064 2627 1068 2631
rect 1176 2627 1180 2631
rect 1264 2627 1268 2631
rect 1288 2627 1292 2631
rect 480 2611 484 2615
rect 536 2611 540 2615
rect 568 2611 572 2615
rect 624 2611 628 2615
rect 656 2611 660 2615
rect 536 2587 540 2591
rect 624 2587 628 2591
rect 1248 2619 1252 2623
rect 2168 2619 2172 2623
rect 2224 2619 2228 2623
rect 2288 2619 2292 2623
rect 2352 2619 2356 2623
rect 2424 2619 2428 2623
rect 2488 2619 2492 2623
rect 2560 2619 2564 2623
rect 2632 2619 2636 2623
rect 2704 2619 2708 2623
rect 2856 2619 2860 2623
rect 2928 2619 2932 2623
rect 3008 2619 3012 2623
rect 3168 2619 3172 2623
rect 744 2611 748 2615
rect 832 2611 836 2615
rect 888 2611 892 2615
rect 920 2611 924 2615
rect 976 2611 980 2615
rect 1008 2611 1012 2615
rect 1064 2611 1068 2615
rect 1096 2611 1100 2615
rect 1184 2611 1188 2615
rect 1240 2611 1244 2615
rect 712 2587 716 2591
rect 888 2587 892 2591
rect 976 2587 980 2591
rect 1064 2587 1068 2591
rect 1240 2587 1244 2591
rect 1272 2611 1276 2615
rect 2224 2595 2228 2599
rect 2352 2595 2356 2599
rect 2488 2595 2492 2599
rect 2632 2595 2636 2599
rect 2928 2595 2932 2599
rect 1248 2583 1252 2587
rect 3040 2563 3044 2567
rect 2192 2523 2196 2527
rect 752 2507 756 2511
rect 840 2507 844 2511
rect 1016 2507 1020 2511
rect 1104 2507 1108 2511
rect 1192 2507 1196 2511
rect 1280 2507 1284 2511
rect 2304 2523 2308 2527
rect 2424 2523 2428 2527
rect 2552 2523 2556 2527
rect 3472 2523 3476 2527
rect 2120 2495 2124 2499
rect 2192 2495 2196 2499
rect 2216 2495 2220 2499
rect 2304 2495 2308 2499
rect 2328 2495 2332 2499
rect 2424 2495 2428 2499
rect 2448 2495 2452 2499
rect 2552 2495 2556 2499
rect 2576 2495 2580 2499
rect 2712 2495 2716 2499
rect 2864 2495 2868 2499
rect 3016 2495 3020 2499
rect 3176 2495 3180 2499
rect 3344 2495 3348 2499
rect 2360 2487 2364 2491
rect 512 2479 516 2483
rect 600 2479 604 2483
rect 688 2479 692 2483
rect 752 2479 756 2483
rect 776 2479 780 2483
rect 840 2479 844 2483
rect 864 2479 868 2483
rect 952 2479 956 2483
rect 1016 2479 1020 2483
rect 1040 2479 1044 2483
rect 1104 2479 1108 2483
rect 1128 2479 1132 2483
rect 1192 2479 1196 2483
rect 1216 2479 1220 2483
rect 1280 2479 1284 2483
rect 1304 2479 1308 2483
rect 2096 2479 2100 2483
rect 2152 2479 2156 2483
rect 2192 2479 2196 2483
rect 2248 2479 2252 2483
rect 2296 2479 2300 2483
rect 2352 2479 2356 2483
rect 368 2463 372 2467
rect 424 2463 428 2467
rect 480 2463 484 2467
rect 600 2463 604 2467
rect 664 2463 668 2467
rect 728 2463 732 2467
rect 856 2463 860 2467
rect 976 2463 980 2467
rect 1032 2463 1036 2467
rect 1096 2463 1100 2467
rect 1216 2463 1220 2467
rect 1280 2463 1284 2467
rect 1344 2463 1348 2467
rect 1408 2463 1412 2467
rect 1472 2463 1476 2467
rect 424 2439 428 2443
rect 1032 2439 1036 2443
rect 1280 2439 1284 2443
rect 2152 2455 2156 2459
rect 2248 2455 2252 2459
rect 2352 2455 2356 2459
rect 3496 2495 3500 2499
rect 2416 2479 2420 2483
rect 2552 2479 2556 2483
rect 2632 2479 2636 2483
rect 2712 2479 2716 2483
rect 2776 2479 2780 2483
rect 2896 2479 2900 2483
rect 2992 2479 2996 2483
rect 3096 2479 3100 2483
rect 3304 2479 3308 2483
rect 3472 2479 3476 2483
rect 3496 2479 3500 2483
rect 2632 2455 2636 2459
rect 2776 2455 2780 2459
rect 2992 2455 2996 2459
rect 2360 2451 2364 2455
rect 1408 2439 1412 2443
rect 664 2435 668 2439
rect 3528 2423 3532 2427
rect 512 2407 516 2411
rect 2056 2379 2060 2383
rect 280 2363 284 2367
rect 152 2335 156 2339
rect 1200 2363 1204 2367
rect 1368 2363 1372 2367
rect 1536 2363 1540 2367
rect 1704 2363 1708 2367
rect 2176 2379 2180 2383
rect 2304 2379 2308 2383
rect 2440 2379 2444 2383
rect 2744 2379 2748 2383
rect 2920 2379 2924 2383
rect 3104 2379 3108 2383
rect 3472 2379 3476 2383
rect 1968 2351 1972 2355
rect 2056 2351 2060 2355
rect 2080 2351 2084 2355
rect 2176 2351 2180 2355
rect 2200 2351 2204 2355
rect 2304 2351 2308 2355
rect 2328 2351 2332 2355
rect 2440 2351 2444 2355
rect 2464 2351 2468 2355
rect 2608 2351 2612 2355
rect 2744 2351 2748 2355
rect 2768 2351 2772 2355
rect 2920 2351 2924 2355
rect 2944 2351 2948 2355
rect 3104 2351 3108 2355
rect 3128 2351 3132 2355
rect 3320 2351 3324 2355
rect 3360 2351 3364 2355
rect 304 2335 308 2339
rect 488 2335 492 2339
rect 680 2335 684 2339
rect 864 2335 868 2339
rect 1048 2335 1052 2339
rect 1200 2335 1204 2339
rect 1224 2335 1228 2339
rect 1368 2335 1372 2339
rect 1392 2335 1396 2339
rect 1536 2335 1540 2339
rect 1560 2335 1564 2339
rect 1704 2335 1708 2339
rect 1728 2335 1732 2339
rect 1904 2331 1908 2335
rect 1960 2331 1964 2335
rect 2016 2331 2020 2335
rect 2088 2331 2092 2335
rect 2168 2331 2172 2335
rect 2240 2331 2244 2335
rect 2320 2331 2324 2335
rect 2392 2331 2396 2335
rect 2472 2331 2476 2335
rect 2624 2331 2628 2335
rect 2744 2331 2748 2335
rect 2784 2331 2788 2335
rect 2952 2331 2956 2335
rect 3032 2331 3036 2335
rect 3120 2331 3124 2335
rect 3208 2331 3212 2335
rect 3296 2331 3300 2335
rect 152 2319 156 2323
rect 280 2319 284 2323
rect 304 2319 308 2323
rect 488 2319 492 2323
rect 584 2319 588 2323
rect 680 2319 684 2323
rect 776 2319 780 2323
rect 872 2319 876 2323
rect 1064 2319 1068 2323
rect 1240 2319 1244 2323
rect 1416 2319 1420 2323
rect 1504 2319 1508 2323
rect 1592 2319 1596 2323
rect 1744 2319 1748 2323
rect 584 2295 588 2299
rect 776 2295 780 2299
rect 1960 2307 1964 2311
rect 2088 2307 2092 2311
rect 2240 2307 2244 2311
rect 2392 2307 2396 2311
rect 2744 2307 2748 2311
rect 3032 2307 3036 2311
rect 3208 2307 3212 2311
rect 1504 2291 1508 2295
rect 184 2263 188 2267
rect 3496 2351 3500 2355
rect 3472 2331 3476 2335
rect 3480 2331 3484 2335
rect 3512 2275 3516 2279
rect 3360 2247 3364 2251
rect 2016 2231 2020 2235
rect 248 2215 252 2219
rect 400 2215 404 2219
rect 1008 2215 1012 2219
rect 1448 2215 1452 2219
rect 2192 2231 2196 2235
rect 2376 2231 2380 2235
rect 2560 2231 2564 2235
rect 2904 2231 2908 2235
rect 3072 2231 3076 2235
rect 3232 2231 3236 2235
rect 1904 2203 1908 2207
rect 2016 2203 2020 2207
rect 2040 2203 2044 2207
rect 2192 2203 2196 2207
rect 2216 2203 2220 2207
rect 2376 2203 2380 2207
rect 2400 2203 2404 2207
rect 2560 2203 2564 2207
rect 2584 2203 2588 2207
rect 2760 2203 2764 2207
rect 2904 2203 2908 2207
rect 2928 2203 2932 2207
rect 3072 2203 3076 2207
rect 3096 2203 3100 2207
rect 3232 2203 3236 2207
rect 3256 2203 3260 2207
rect 3424 2203 3428 2207
rect 152 2187 156 2191
rect 248 2187 252 2191
rect 272 2187 276 2191
rect 400 2187 404 2191
rect 424 2187 428 2191
rect 576 2187 580 2191
rect 688 2187 692 2191
rect 736 2187 740 2191
rect 888 2187 892 2191
rect 1008 2187 1012 2191
rect 1032 2187 1036 2191
rect 1176 2187 1180 2191
rect 1320 2187 1324 2191
rect 1448 2187 1452 2191
rect 1472 2187 1476 2191
rect 1880 2187 1884 2191
rect 1904 2187 1908 2191
rect 1960 2187 1964 2191
rect 2048 2187 2052 2191
rect 2136 2187 2140 2191
rect 2224 2187 2228 2191
rect 2312 2187 2316 2191
rect 2408 2187 2412 2191
rect 2496 2187 2500 2191
rect 2592 2187 2596 2191
rect 2768 2187 2772 2191
rect 2856 2187 2860 2191
rect 2928 2187 2932 2191
rect 3000 2187 3004 2191
rect 3080 2187 3084 2191
rect 3152 2187 3156 2191
rect 3224 2187 3228 2191
rect 3296 2187 3300 2191
rect 3368 2187 3372 2191
rect 3496 2187 3500 2191
rect 224 2171 228 2175
rect 280 2171 284 2175
rect 320 2171 324 2175
rect 424 2171 428 2175
rect 480 2171 484 2175
rect 528 2171 532 2175
rect 584 2171 588 2175
rect 632 2171 636 2175
rect 280 2147 284 2151
rect 480 2147 484 2151
rect 584 2147 588 2151
rect 1128 2179 1132 2183
rect 736 2171 740 2175
rect 792 2171 796 2175
rect 840 2171 844 2175
rect 952 2171 956 2175
rect 1064 2171 1068 2175
rect 1120 2171 1124 2175
rect 688 2147 692 2151
rect 792 2147 796 2151
rect 1120 2147 1124 2151
rect 1176 2171 1180 2175
rect 1128 2143 1132 2147
rect 352 2115 356 2119
rect 872 2115 876 2119
rect 1960 2163 1964 2167
rect 2136 2163 2140 2167
rect 2312 2163 2316 2167
rect 2496 2163 2500 2167
rect 2856 2163 2860 2167
rect 3000 2163 3004 2167
rect 3152 2163 3156 2167
rect 3296 2163 3300 2167
rect 3528 2131 3532 2135
rect 1880 2103 1884 2107
rect 2368 2087 2372 2091
rect 408 2083 412 2087
rect 336 2039 340 2043
rect 416 2067 420 2071
rect 600 2067 604 2071
rect 704 2067 708 2071
rect 920 2067 924 2071
rect 1024 2067 1028 2071
rect 1128 2067 1132 2071
rect 2544 2087 2548 2091
rect 1904 2059 1908 2063
rect 2040 2059 2044 2063
rect 2216 2059 2220 2063
rect 2368 2059 2372 2063
rect 2392 2059 2396 2063
rect 2544 2059 2548 2063
rect 2568 2059 2572 2063
rect 2736 2059 2740 2063
rect 2896 2059 2900 2063
rect 3048 2059 3052 2063
rect 3192 2059 3196 2063
rect 3336 2059 3340 2063
rect 3488 2059 3492 2063
rect 416 2039 420 2043
rect 440 2039 444 2043
rect 544 2039 548 2043
rect 600 2039 604 2043
rect 648 2039 652 2043
rect 704 2039 708 2043
rect 752 2039 756 2043
rect 848 2039 852 2043
rect 920 2039 924 2043
rect 944 2039 948 2043
rect 1024 2039 1028 2043
rect 1048 2039 1052 2043
rect 1128 2039 1132 2043
rect 1152 2039 1156 2043
rect 1256 2039 1260 2043
rect 1904 2039 1908 2043
rect 2024 2039 2028 2043
rect 2160 2039 2164 2043
rect 2304 2039 2308 2043
rect 2448 2039 2452 2043
rect 2600 2039 2604 2043
rect 2768 2039 2772 2043
rect 2944 2039 2948 2043
rect 3032 2039 3036 2043
rect 3128 2039 3132 2043
rect 3320 2039 3324 2043
rect 3496 2039 3500 2043
rect 224 2019 228 2023
rect 288 2019 292 2023
rect 400 2019 404 2023
rect 408 2019 412 2023
rect 568 2019 572 2023
rect 728 2019 732 2023
rect 872 2019 876 2023
rect 1008 2019 1012 2023
rect 1136 2019 1140 2023
rect 1216 2019 1220 2023
rect 1256 2019 1260 2023
rect 1376 2019 1380 2023
rect 1504 2019 1508 2023
rect 3032 2015 3036 2019
rect 1216 1995 1220 1999
rect 288 1991 292 1995
rect 3528 1983 3532 1987
rect 2104 1939 2108 1943
rect 512 1915 516 1919
rect 1256 1915 1260 1919
rect 1416 1915 1420 1919
rect 1576 1915 1580 1919
rect 1720 1915 1724 1919
rect 2192 1939 2196 1943
rect 2280 1939 2284 1943
rect 2376 1939 2380 1943
rect 3472 1939 3476 1943
rect 2040 1911 2044 1915
rect 2104 1911 2108 1915
rect 2128 1911 2132 1915
rect 2192 1911 2196 1915
rect 2216 1911 2220 1915
rect 2280 1911 2284 1915
rect 2304 1911 2308 1915
rect 2376 1911 2380 1915
rect 2400 1911 2404 1915
rect 2520 1911 2524 1915
rect 2672 1911 2676 1915
rect 2856 1911 2860 1915
rect 3064 1911 3068 1915
rect 3288 1911 3292 1915
rect 3496 1911 3500 1915
rect 2184 1891 2188 1895
rect 2272 1891 2276 1895
rect 2360 1891 2364 1895
rect 2448 1891 2452 1895
rect 2512 1891 2516 1895
rect 2536 1891 2540 1895
rect 2648 1891 2652 1895
rect 2712 1891 2716 1895
rect 2784 1891 2788 1895
rect 2944 1891 2948 1895
rect 3032 1891 3036 1895
rect 3128 1891 3132 1895
rect 3224 1891 3228 1895
rect 3320 1891 3324 1895
rect 3472 1891 3476 1895
rect 3496 1891 3500 1895
rect 152 1887 156 1891
rect 328 1887 332 1891
rect 512 1887 516 1891
rect 536 1887 540 1891
rect 736 1887 740 1891
rect 928 1887 932 1891
rect 1112 1887 1116 1891
rect 1256 1887 1260 1891
rect 1280 1887 1284 1891
rect 1416 1887 1420 1891
rect 1440 1887 1444 1891
rect 1576 1887 1580 1891
rect 1600 1887 1604 1891
rect 1720 1887 1724 1891
rect 1744 1887 1748 1891
rect 152 1867 156 1871
rect 320 1867 324 1871
rect 520 1867 524 1871
rect 616 1867 620 1871
rect 712 1867 716 1871
rect 800 1867 804 1871
rect 896 1867 900 1871
rect 1072 1867 1076 1871
rect 1144 1867 1148 1871
rect 1240 1867 1244 1871
rect 1400 1867 1404 1871
rect 1480 1867 1484 1871
rect 1560 1867 1564 1871
rect 1640 1867 1644 1871
rect 1720 1867 1724 1871
rect 2712 1867 2716 1871
rect 3032 1867 3036 1871
rect 3224 1867 3228 1871
rect 616 1843 620 1847
rect 800 1843 804 1847
rect 1144 1843 1148 1847
rect 1480 1839 1484 1843
rect 2512 1863 2516 1867
rect 1640 1839 1644 1843
rect 3528 1835 3532 1839
rect 184 1811 188 1815
rect 2432 1791 2436 1795
rect 2912 1791 2916 1795
rect 3040 1791 3044 1795
rect 3176 1791 3180 1795
rect 3312 1791 3316 1795
rect 256 1763 260 1767
rect 560 1763 564 1767
rect 712 1763 716 1767
rect 1416 1763 1420 1767
rect 2336 1763 2340 1767
rect 2432 1763 2436 1767
rect 2456 1763 2460 1767
rect 2576 1763 2580 1767
rect 2696 1763 2700 1767
rect 2816 1763 2820 1767
rect 2912 1763 2916 1767
rect 2936 1763 2940 1767
rect 3040 1763 3044 1767
rect 3064 1763 3068 1767
rect 3176 1763 3180 1767
rect 3200 1763 3204 1767
rect 3312 1763 3316 1767
rect 3336 1763 3340 1767
rect 3480 1763 3484 1767
rect 3328 1751 3332 1755
rect 2304 1743 2308 1747
rect 2360 1743 2364 1747
rect 2416 1743 2420 1747
rect 2472 1743 2476 1747
rect 2536 1743 2540 1747
rect 2600 1743 2604 1747
rect 2664 1743 2668 1747
rect 2784 1743 2788 1747
rect 2904 1743 2908 1747
rect 3024 1743 3028 1747
rect 3144 1743 3148 1747
rect 3200 1743 3204 1747
rect 3264 1743 3268 1747
rect 152 1735 156 1739
rect 256 1735 260 1739
rect 280 1735 284 1739
rect 432 1735 436 1739
rect 560 1735 564 1739
rect 584 1735 588 1739
rect 712 1735 716 1739
rect 736 1735 740 1739
rect 880 1735 884 1739
rect 1024 1735 1028 1739
rect 1160 1735 1164 1739
rect 1296 1735 1300 1739
rect 1416 1735 1420 1739
rect 1440 1735 1444 1739
rect 152 1723 156 1727
rect 288 1723 292 1727
rect 440 1723 444 1727
rect 568 1723 572 1727
rect 592 1723 596 1727
rect 736 1723 740 1727
rect 800 1723 804 1727
rect 872 1723 876 1727
rect 936 1723 940 1727
rect 1000 1723 1004 1727
rect 1064 1723 1068 1727
rect 1136 1723 1140 1727
rect 1248 1723 1252 1727
rect 1272 1723 1276 1727
rect 184 1667 188 1671
rect 800 1699 804 1703
rect 936 1699 940 1703
rect 1064 1699 1068 1703
rect 2360 1719 2364 1723
rect 2472 1719 2476 1723
rect 2600 1719 2604 1723
rect 3200 1719 3204 1723
rect 3392 1743 3396 1747
rect 3496 1743 3500 1747
rect 3328 1715 3332 1719
rect 1248 1699 1252 1703
rect 3528 1687 3532 1691
rect 568 1643 572 1647
rect 2240 1643 2244 1647
rect 256 1627 260 1631
rect 568 1627 572 1631
rect 1000 1627 1004 1631
rect 1272 1627 1276 1631
rect 1408 1627 1412 1631
rect 2360 1643 2364 1647
rect 2496 1643 2500 1647
rect 2640 1643 2644 1647
rect 3472 1643 3476 1647
rect 2160 1615 2164 1619
rect 2240 1615 2244 1619
rect 2264 1615 2268 1619
rect 2360 1615 2364 1619
rect 2384 1615 2388 1619
rect 2496 1615 2500 1619
rect 2520 1615 2524 1619
rect 2640 1615 2644 1619
rect 2664 1615 2668 1619
rect 2824 1615 2828 1619
rect 2992 1615 2996 1619
rect 3160 1615 3164 1619
rect 3336 1615 3340 1619
rect 3496 1615 3500 1619
rect 2016 1603 2020 1607
rect 2072 1603 2076 1607
rect 2112 1603 2116 1607
rect 2168 1603 2172 1607
rect 2216 1603 2220 1607
rect 2272 1603 2276 1607
rect 2336 1603 2340 1607
rect 2400 1603 2404 1607
rect 2472 1603 2476 1607
rect 2616 1603 2620 1607
rect 2696 1603 2700 1607
rect 2776 1603 2780 1607
rect 2848 1603 2852 1607
rect 2952 1603 2956 1607
rect 3136 1603 3140 1607
rect 3200 1603 3204 1607
rect 3328 1603 3332 1607
rect 3472 1603 3476 1607
rect 3496 1603 3500 1607
rect 152 1599 156 1603
rect 256 1599 260 1603
rect 280 1599 284 1603
rect 440 1599 444 1603
rect 568 1599 572 1603
rect 592 1599 596 1603
rect 744 1599 748 1603
rect 888 1599 892 1603
rect 1000 1599 1004 1603
rect 1024 1599 1028 1603
rect 1160 1599 1164 1603
rect 1272 1599 1276 1603
rect 1296 1599 1300 1603
rect 1408 1599 1412 1603
rect 1432 1599 1436 1603
rect 176 1583 180 1587
rect 248 1583 252 1587
rect 344 1583 348 1587
rect 520 1583 524 1587
rect 600 1583 604 1587
rect 688 1583 692 1587
rect 856 1583 860 1587
rect 1008 1583 1012 1587
rect 1080 1583 1084 1587
rect 1160 1583 1164 1587
rect 1232 1583 1236 1587
rect 1304 1583 1308 1587
rect 1376 1583 1380 1587
rect 1448 1583 1452 1587
rect 1520 1583 1524 1587
rect 1592 1583 1596 1587
rect 248 1559 252 1563
rect 600 1559 604 1563
rect 1080 1559 1084 1563
rect 1232 1559 1236 1563
rect 1376 1559 1380 1563
rect 2072 1579 2076 1583
rect 2168 1579 2172 1583
rect 2272 1579 2276 1583
rect 2400 1579 2404 1583
rect 2696 1575 2700 1579
rect 2848 1575 2852 1579
rect 3200 1575 3204 1579
rect 1520 1559 1524 1563
rect 1968 1499 1972 1503
rect 752 1483 756 1487
rect 928 1483 932 1487
rect 1248 1483 1252 1487
rect 1400 1483 1404 1487
rect 1552 1483 1556 1487
rect 1704 1483 1708 1487
rect 2232 1499 2236 1503
rect 2376 1499 2380 1503
rect 2480 1499 2484 1503
rect 1904 1471 1908 1475
rect 1968 1471 1972 1475
rect 1992 1471 1996 1475
rect 2120 1471 2124 1475
rect 2232 1471 2236 1475
rect 2256 1471 2260 1475
rect 2376 1471 2380 1475
rect 2400 1471 2404 1475
rect 3048 1499 3052 1503
rect 2560 1471 2564 1475
rect 2728 1471 2732 1475
rect 2896 1471 2900 1475
rect 3048 1471 3052 1475
rect 3072 1471 3076 1475
rect 3256 1471 3260 1475
rect 3264 1471 3268 1475
rect 3448 1471 3452 1475
rect 3208 1463 3212 1467
rect 232 1455 236 1459
rect 408 1455 412 1459
rect 592 1455 596 1459
rect 752 1455 756 1459
rect 776 1455 780 1459
rect 928 1455 932 1459
rect 952 1455 956 1459
rect 1112 1455 1116 1459
rect 1248 1455 1252 1459
rect 1272 1455 1276 1459
rect 1400 1455 1404 1459
rect 1424 1455 1428 1459
rect 1552 1455 1556 1459
rect 1576 1455 1580 1459
rect 1704 1455 1708 1459
rect 1728 1455 1732 1459
rect 1808 1455 1812 1459
rect 1904 1455 1908 1459
rect 1960 1455 1964 1459
rect 2032 1455 2036 1459
rect 2104 1455 2108 1459
rect 2184 1455 2188 1459
rect 2328 1455 2332 1459
rect 2472 1455 2476 1459
rect 2480 1455 2484 1459
rect 2624 1455 2628 1459
rect 2696 1455 2700 1459
rect 2776 1455 2780 1459
rect 2944 1455 2948 1459
rect 3112 1455 3116 1459
rect 3200 1455 3204 1459
rect 264 1439 268 1443
rect 392 1439 396 1443
rect 456 1439 460 1443
rect 528 1439 532 1443
rect 680 1439 684 1443
rect 760 1439 764 1443
rect 840 1439 844 1443
rect 1000 1439 1004 1443
rect 1080 1439 1084 1443
rect 1152 1439 1156 1443
rect 1304 1439 1308 1443
rect 1376 1439 1380 1443
rect 1456 1439 1460 1443
rect 1528 1439 1532 1443
rect 1608 1439 1612 1443
rect 1744 1439 1748 1443
rect 456 1415 460 1419
rect 760 1415 764 1419
rect 1376 1415 1380 1419
rect 1528 1415 1532 1419
rect 1960 1431 1964 1435
rect 2104 1431 2108 1435
rect 2696 1431 2700 1435
rect 3200 1431 3204 1435
rect 3208 1427 3212 1431
rect 1808 1415 1812 1419
rect 1080 1411 1084 1415
rect 560 1383 564 1387
rect 3288 1455 3292 1459
rect 3472 1455 3476 1459
rect 3504 1399 3508 1403
rect 3264 1363 3268 1367
rect 2384 1347 2388 1351
rect 432 1343 436 1347
rect 696 1343 700 1347
rect 368 1315 372 1319
rect 432 1315 436 1319
rect 456 1315 460 1319
rect 544 1317 548 1321
rect 1120 1343 1124 1347
rect 1272 1343 1276 1347
rect 1584 1343 1588 1347
rect 1720 1343 1724 1347
rect 640 1315 644 1319
rect 696 1315 700 1319
rect 744 1315 748 1319
rect 864 1315 868 1319
rect 1000 1315 1004 1319
rect 1120 1315 1124 1319
rect 1144 1315 1148 1319
rect 1272 1315 1276 1319
rect 1296 1315 1300 1319
rect 1448 1315 1452 1319
rect 1584 1315 1588 1319
rect 1608 1315 1612 1319
rect 1904 1319 1908 1323
rect 2160 1319 2164 1323
rect 1744 1315 1748 1319
rect 3056 1347 3060 1351
rect 3472 1347 3476 1351
rect 2408 1319 2412 1323
rect 2640 1319 2644 1323
rect 2864 1319 2868 1323
rect 3056 1319 3060 1323
rect 3080 1319 3084 1323
rect 3288 1319 3292 1323
rect 3496 1319 3500 1323
rect 1936 1307 1940 1311
rect 2120 1307 2124 1311
rect 2208 1307 2212 1311
rect 2296 1307 2300 1311
rect 2384 1307 2388 1311
rect 2464 1307 2468 1311
rect 2632 1307 2636 1311
rect 2800 1307 2804 1311
rect 2968 1307 2972 1311
rect 3056 1307 3060 1311
rect 3144 1307 3148 1311
rect 3232 1307 3236 1311
rect 3328 1307 3332 1311
rect 3472 1307 3476 1311
rect 3496 1307 3500 1311
rect 464 1303 468 1307
rect 520 1303 524 1307
rect 552 1303 556 1307
rect 608 1303 612 1307
rect 640 1303 644 1307
rect 696 1303 700 1307
rect 728 1303 732 1307
rect 784 1303 788 1307
rect 840 1303 844 1307
rect 976 1303 980 1307
rect 1144 1303 1148 1307
rect 1336 1303 1340 1307
rect 1544 1303 1548 1307
rect 1720 1303 1724 1307
rect 1744 1303 1748 1307
rect 520 1279 524 1283
rect 608 1279 612 1283
rect 696 1279 700 1283
rect 784 1279 788 1283
rect 3056 1283 3060 1287
rect 3232 1283 3236 1287
rect 2208 1279 2212 1283
rect 2496 1251 2500 1255
rect 3360 1251 3364 1255
rect 3528 1251 3532 1255
rect 624 1207 628 1211
rect 712 1207 716 1211
rect 560 1179 564 1183
rect 624 1179 628 1183
rect 648 1179 652 1183
rect 888 1207 892 1211
rect 736 1179 740 1183
rect 824 1181 828 1185
rect 1088 1207 1092 1211
rect 1200 1207 1204 1211
rect 1328 1207 1332 1211
rect 1464 1207 1468 1211
rect 1720 1207 1724 1211
rect 2472 1203 2476 1207
rect 888 1179 892 1183
rect 912 1179 916 1183
rect 1008 1179 1012 1183
rect 1088 1179 1092 1183
rect 1112 1179 1116 1183
rect 1200 1179 1204 1183
rect 1224 1179 1228 1183
rect 1328 1179 1332 1183
rect 1352 1179 1356 1183
rect 1464 1179 1468 1183
rect 1488 1179 1492 1183
rect 1624 1179 1628 1183
rect 1720 1179 1724 1183
rect 1744 1179 1748 1183
rect 2160 1175 2164 1179
rect 2336 1175 2340 1179
rect 1376 1167 1380 1171
rect 3472 1203 3476 1207
rect 2504 1175 2508 1179
rect 2672 1175 2676 1179
rect 2840 1175 2844 1179
rect 3008 1175 3012 1179
rect 3176 1175 3180 1179
rect 3344 1175 3348 1179
rect 3496 1175 3500 1179
rect 368 1159 372 1163
rect 424 1159 428 1163
rect 480 1159 484 1163
rect 536 1159 540 1163
rect 600 1159 604 1163
rect 712 1159 716 1163
rect 720 1159 724 1163
rect 840 1159 844 1163
rect 960 1159 964 1163
rect 1072 1159 1076 1163
rect 1192 1159 1196 1163
rect 1312 1159 1316 1163
rect 1368 1159 1372 1163
rect 424 1135 428 1139
rect 536 1135 540 1139
rect 1368 1135 1372 1139
rect 1904 1163 1908 1167
rect 1960 1163 1964 1167
rect 2016 1163 2020 1167
rect 2080 1163 2084 1167
rect 2152 1163 2156 1167
rect 2304 1163 2308 1167
rect 2464 1163 2468 1167
rect 2472 1163 2476 1167
rect 2632 1163 2636 1167
rect 2800 1163 2804 1167
rect 2888 1163 2892 1167
rect 2976 1163 2980 1167
rect 3152 1163 3156 1167
rect 3232 1163 3236 1167
rect 3336 1163 3340 1167
rect 3472 1163 3476 1167
rect 3496 1163 3500 1167
rect 1432 1159 1436 1163
rect 1960 1139 1964 1143
rect 2080 1139 2084 1143
rect 2888 1139 2892 1143
rect 3232 1139 3236 1143
rect 1376 1131 1380 1135
rect 3368 1107 3372 1111
rect 3528 1107 3532 1111
rect 632 1103 636 1107
rect 280 1059 284 1063
rect 440 1059 444 1063
rect 776 1059 780 1063
rect 1096 1059 1100 1063
rect 1552 1059 1556 1063
rect 160 1031 164 1035
rect 280 1031 284 1035
rect 304 1031 308 1035
rect 440 1031 444 1035
rect 464 1031 468 1035
rect 632 1031 636 1035
rect 776 1031 780 1035
rect 800 1031 804 1035
rect 960 1031 964 1035
rect 1096 1031 1100 1035
rect 1120 1031 1124 1035
rect 1272 1031 1276 1035
rect 1424 1031 1428 1035
rect 1552 1031 1556 1035
rect 1576 1031 1580 1035
rect 1912 1031 1916 1035
rect 2064 1031 2068 1035
rect 2232 1031 2236 1035
rect 2408 1031 2412 1035
rect 2584 1031 2588 1035
rect 2704 1031 2708 1035
rect 2752 1031 2756 1035
rect 2912 1031 2916 1035
rect 3064 1031 3068 1035
rect 3216 1031 3220 1035
rect 3368 1031 3372 1035
rect 3496 1031 3500 1035
rect 152 1015 156 1019
rect 256 1015 260 1019
rect 296 1015 300 1019
rect 480 1015 484 1019
rect 576 1015 580 1019
rect 672 1015 676 1019
rect 760 1015 764 1019
rect 856 1015 860 1019
rect 1040 1015 1044 1019
rect 1128 1015 1132 1019
rect 1216 1015 1220 1019
rect 1296 1015 1300 1019
rect 1384 1015 1388 1019
rect 1552 1015 1556 1019
rect 1720 1015 1724 1019
rect 1984 1015 1988 1019
rect 2104 1015 2108 1019
rect 2168 1015 2172 1019
rect 2232 1015 2236 1019
rect 2296 1015 2300 1019
rect 2368 1015 2372 1019
rect 2504 1015 2508 1019
rect 2648 1015 2652 1019
rect 256 991 260 995
rect 576 991 580 995
rect 760 991 764 995
rect 1128 991 1132 995
rect 1296 991 1300 995
rect 2168 991 2172 995
rect 2296 991 2300 995
rect 2800 1015 2804 1019
rect 2904 1015 2908 1019
rect 2968 1015 2972 1019
rect 3056 1015 3060 1019
rect 3144 1015 3148 1019
rect 3232 1015 3236 1019
rect 3320 1015 3324 1019
rect 3496 1015 3500 1019
rect 2704 991 2708 995
rect 2904 991 2908 995
rect 3056 991 3060 995
rect 3232 991 3236 995
rect 456 975 460 979
rect 128 915 132 919
rect 2536 959 2540 963
rect 656 915 660 919
rect 848 915 852 919
rect 1216 915 1220 919
rect 1392 915 1396 919
rect 1568 915 1572 919
rect 1720 915 1724 919
rect 2120 915 2124 919
rect 152 887 156 891
rect 304 887 308 891
rect 456 887 460 891
rect 488 887 492 891
rect 656 887 660 891
rect 680 887 684 891
rect 848 887 852 891
rect 872 887 876 891
rect 1064 887 1068 891
rect 1216 887 1220 891
rect 1240 887 1244 891
rect 1392 887 1396 891
rect 1416 887 1420 891
rect 1568 887 1572 891
rect 1592 887 1596 891
rect 1720 887 1724 891
rect 1744 887 1748 891
rect 2160 887 2164 891
rect 2248 887 2252 891
rect 2336 887 2340 891
rect 2424 887 2428 891
rect 2520 887 2524 891
rect 2552 887 2556 891
rect 2632 887 2636 891
rect 2768 887 2772 891
rect 2920 887 2924 891
rect 3096 887 3100 891
rect 3280 887 3284 891
rect 3472 887 3476 891
rect 128 871 132 875
rect 152 871 156 875
rect 224 871 228 875
rect 296 871 300 875
rect 456 871 460 875
rect 480 871 484 875
rect 568 871 572 875
rect 664 871 668 875
rect 752 871 756 875
rect 848 871 852 875
rect 1032 871 1036 875
rect 1096 871 1100 875
rect 1200 871 1204 875
rect 1280 871 1284 875
rect 1368 871 1372 875
rect 1448 871 1452 875
rect 1536 871 1540 875
rect 1616 871 1620 875
rect 1704 871 1708 875
rect 2112 871 2116 875
rect 2120 871 2124 875
rect 2168 871 2172 875
rect 2200 871 2204 875
rect 2256 871 2260 875
rect 2288 871 2292 875
rect 2376 871 2380 875
rect 2432 871 2436 875
rect 2464 871 2468 875
rect 224 847 228 851
rect 456 847 460 851
rect 568 847 572 851
rect 752 847 756 851
rect 1096 847 1100 851
rect 1280 847 1284 851
rect 1448 847 1452 851
rect 1616 847 1620 851
rect 2168 847 2172 851
rect 2256 847 2260 851
rect 2432 847 2436 851
rect 2576 871 2580 875
rect 2640 871 2644 875
rect 2712 871 2716 875
rect 2776 871 2780 875
rect 2880 871 2884 875
rect 2968 871 2972 875
rect 3064 871 3068 875
rect 3160 871 3164 875
rect 3264 871 3268 875
rect 3472 871 3476 875
rect 2552 847 2556 851
rect 2640 847 2644 851
rect 2776 847 2780 851
rect 2968 847 2972 851
rect 3160 847 3164 851
rect 2320 815 2324 819
rect 3504 815 3508 819
rect 264 775 268 779
rect 416 775 420 779
rect 576 775 580 779
rect 736 775 740 779
rect 1032 775 1036 779
rect 1176 775 1180 779
rect 1320 775 1324 779
rect 1472 775 1476 779
rect 2368 775 2372 779
rect 2776 775 2780 779
rect 2928 775 2932 779
rect 3104 775 3108 779
rect 3288 775 3292 779
rect 152 747 156 751
rect 264 747 268 751
rect 288 747 292 751
rect 416 747 420 751
rect 440 747 444 751
rect 576 747 580 751
rect 600 747 604 751
rect 736 747 740 751
rect 760 747 764 751
rect 912 747 916 751
rect 1032 747 1036 751
rect 1056 747 1060 751
rect 1176 747 1180 751
rect 1200 747 1204 751
rect 1320 747 1324 751
rect 1344 747 1348 751
rect 1472 747 1476 751
rect 1496 747 1500 751
rect 2216 747 2220 751
rect 2304 747 2308 751
rect 2368 747 2372 751
rect 2392 747 2396 751
rect 2480 747 2484 751
rect 2568 747 2572 751
rect 2672 747 2676 751
rect 2776 747 2780 751
rect 2800 747 2804 751
rect 2928 747 2932 751
rect 2952 747 2956 751
rect 3104 747 3108 751
rect 3128 747 3132 751
rect 3288 747 3292 751
rect 3312 747 3316 751
rect 3496 747 3500 751
rect 368 731 372 735
rect 424 731 428 735
rect 456 731 460 735
rect 512 731 516 735
rect 552 731 556 735
rect 608 731 612 735
rect 648 731 652 735
rect 704 731 708 735
rect 744 731 748 735
rect 840 731 844 735
rect 896 731 900 735
rect 936 731 940 735
rect 992 731 996 735
rect 1040 731 1044 735
rect 1096 731 1100 735
rect 1144 731 1148 735
rect 1224 731 1228 735
rect 1248 731 1252 735
rect 1952 731 1956 735
rect 2112 731 2116 735
rect 2264 731 2268 735
rect 2336 731 2340 735
rect 2416 731 2420 735
rect 2488 731 2492 735
rect 2560 731 2564 735
rect 2704 731 2708 735
rect 2768 731 2772 735
rect 2848 731 2852 735
rect 2920 731 2924 735
rect 2992 731 2996 735
rect 3064 731 3068 735
rect 3144 731 3148 735
rect 3296 731 3300 735
rect 3448 731 3452 735
rect 424 707 428 711
rect 512 707 516 711
rect 608 707 612 711
rect 704 707 708 711
rect 896 707 900 711
rect 992 707 996 711
rect 1096 707 1100 711
rect 1224 707 1228 711
rect 2336 707 2340 711
rect 2488 707 2492 711
rect 2768 707 2772 711
rect 2920 707 2924 711
rect 3064 707 3068 711
rect 560 631 564 635
rect 648 631 652 635
rect 736 631 740 635
rect 824 631 828 635
rect 912 631 916 635
rect 496 603 500 607
rect 560 603 564 607
rect 584 603 588 607
rect 648 603 652 607
rect 672 603 676 607
rect 736 603 740 607
rect 760 603 764 607
rect 824 603 828 607
rect 848 603 852 607
rect 1176 631 1180 635
rect 2016 631 2020 635
rect 2192 631 2196 635
rect 3056 631 3060 635
rect 3344 631 3348 635
rect 3472 631 3476 635
rect 936 603 940 607
rect 1024 603 1028 607
rect 1112 603 1116 607
rect 1176 603 1180 607
rect 1200 603 1204 607
rect 1288 603 1292 607
rect 1416 603 1420 607
rect 1904 603 1908 607
rect 2016 603 2020 607
rect 2040 603 2044 607
rect 2192 603 2196 607
rect 2216 603 2220 607
rect 2400 603 2404 607
rect 2576 603 2580 607
rect 2584 603 2588 607
rect 2760 603 2764 607
rect 2928 603 2932 607
rect 3056 603 3060 607
rect 3080 603 3084 607
rect 3224 603 3228 607
rect 3344 603 3348 607
rect 3368 603 3372 607
rect 512 591 516 595
rect 568 591 572 595
rect 608 591 612 595
rect 664 591 668 595
rect 712 591 716 595
rect 824 591 828 595
rect 912 591 916 595
rect 944 591 948 595
rect 1072 591 1076 595
rect 1128 591 1132 595
rect 1200 591 1204 595
rect 1264 591 1268 595
rect 1336 591 1340 595
rect 1408 591 1412 595
rect 568 567 572 571
rect 664 567 668 571
rect 1128 567 1132 571
rect 1264 567 1268 571
rect 1408 567 1412 571
rect 1480 591 1484 595
rect 1624 591 1628 595
rect 1744 591 1748 595
rect 1904 591 1908 595
rect 2096 591 2100 595
rect 2280 591 2284 595
rect 2312 591 2316 595
rect 2416 591 2420 595
rect 2520 591 2524 595
rect 1416 563 1420 567
rect 2416 567 2420 571
rect 3496 603 3500 607
rect 2712 591 2716 595
rect 2776 591 2780 595
rect 2888 591 2892 595
rect 3048 591 3052 595
rect 3128 591 3132 595
rect 3208 591 3212 595
rect 3360 591 3364 595
rect 3472 591 3476 595
rect 3496 591 3500 595
rect 2576 567 2580 571
rect 2776 567 2780 571
rect 3128 567 3132 571
rect 2280 503 2284 507
rect 1360 495 1364 499
rect 1696 495 1700 499
rect 2280 487 2284 491
rect 176 467 180 471
rect 320 467 324 471
rect 480 467 484 471
rect 648 467 652 471
rect 816 467 820 471
rect 976 467 980 471
rect 1120 467 1124 471
rect 1256 467 1260 471
rect 1360 467 1364 471
rect 1384 467 1388 471
rect 1512 467 1516 471
rect 1640 467 1644 471
rect 1696 467 1700 471
rect 1744 467 1748 471
rect 2840 487 2844 491
rect 3008 487 3012 491
rect 3168 487 3172 491
rect 2096 459 2100 463
rect 2280 459 2284 463
rect 2304 459 2308 463
rect 2504 459 2508 463
rect 2688 459 2692 463
rect 2840 459 2844 463
rect 2864 459 2868 463
rect 3008 459 3012 463
rect 3032 459 3036 463
rect 3192 459 3196 463
rect 3352 459 3356 463
rect 3496 459 3500 463
rect 152 447 156 451
rect 216 447 220 451
rect 280 447 284 451
rect 448 447 452 451
rect 536 447 540 451
rect 624 447 628 451
rect 712 447 716 451
rect 800 447 804 451
rect 944 447 948 451
rect 976 447 980 451
rect 1056 447 1060 451
rect 1136 447 1140 451
rect 1272 447 1276 451
rect 1296 447 1300 451
rect 1456 447 1460 451
rect 1536 447 1540 451
rect 1616 447 1620 451
rect 2256 447 2260 451
rect 2312 447 2316 451
rect 2344 447 2348 451
rect 2400 447 2404 451
rect 2440 447 2444 451
rect 2496 447 2500 451
rect 2536 447 2540 451
rect 2632 447 2636 451
rect 2744 447 2748 451
rect 2800 447 2804 451
rect 2872 447 2876 451
rect 3016 447 3020 451
rect 3168 447 3172 451
rect 3176 447 3180 451
rect 3256 447 3260 451
rect 3344 447 3348 451
rect 3472 447 3476 451
rect 3496 447 3500 451
rect 216 423 220 427
rect 536 423 540 427
rect 712 423 716 427
rect 1056 423 1060 427
rect 1272 423 1276 427
rect 1536 423 1540 427
rect 2312 423 2316 427
rect 2400 423 2404 427
rect 2496 423 2500 427
rect 2800 423 2804 427
rect 3256 423 3260 427
rect 3264 439 3268 443
rect 3264 419 3268 423
rect 944 367 948 371
rect 3472 367 3476 371
rect 256 351 260 355
rect 424 351 428 355
rect 600 351 604 355
rect 776 351 780 355
rect 1424 351 1428 355
rect 1584 351 1588 355
rect 2232 351 2236 355
rect 2320 351 2324 355
rect 2408 351 2412 355
rect 2496 351 2500 355
rect 3096 351 3100 355
rect 3296 351 3300 355
rect 152 323 156 327
rect 256 323 260 327
rect 280 323 284 327
rect 424 323 428 327
rect 448 323 452 327
rect 600 323 604 327
rect 624 323 628 327
rect 776 323 780 327
rect 800 323 804 327
rect 968 323 972 327
rect 1128 323 1132 327
rect 1288 323 1292 327
rect 1424 323 1428 327
rect 1448 323 1452 327
rect 1584 323 1588 327
rect 1608 323 1612 327
rect 2168 323 2172 327
rect 2232 323 2236 327
rect 2256 323 2260 327
rect 2320 323 2324 327
rect 2344 323 2348 327
rect 2408 323 2412 327
rect 2432 323 2436 327
rect 2496 323 2500 327
rect 2520 323 2524 327
rect 2632 323 2636 327
rect 2768 323 2772 327
rect 2936 323 2940 327
rect 3096 323 3100 327
rect 3120 323 3124 327
rect 3296 323 3300 327
rect 3320 323 3324 327
rect 3472 323 3476 327
rect 3496 323 3500 327
rect 2032 311 2036 315
rect 2088 311 2092 315
rect 2128 311 2132 315
rect 2184 311 2188 315
rect 2232 311 2236 315
rect 2288 311 2292 315
rect 2336 311 2340 315
rect 2440 311 2444 315
rect 2544 311 2548 315
rect 2600 311 2604 315
rect 2648 311 2652 315
rect 2704 311 2708 315
rect 2752 311 2756 315
rect 2808 311 2812 315
rect 2864 311 2868 315
rect 2920 311 2924 315
rect 2976 311 2980 315
rect 272 307 276 311
rect 400 307 404 311
rect 464 307 468 311
rect 536 307 540 311
rect 608 307 612 311
rect 688 307 692 311
rect 768 307 772 311
rect 848 307 852 311
rect 984 307 988 311
rect 1016 307 1020 311
rect 1088 307 1092 311
rect 1184 307 1188 311
rect 1352 307 1356 311
rect 1520 307 1524 311
rect 1608 307 1612 311
rect 1696 307 1700 311
rect 464 283 468 287
rect 608 283 612 287
rect 768 283 772 287
rect 1088 283 1092 287
rect 2088 287 2092 291
rect 2184 287 2188 291
rect 2288 287 2292 291
rect 2600 287 2604 291
rect 2704 287 2708 291
rect 2808 287 2812 291
rect 2920 287 2924 291
rect 1608 279 1612 283
rect 3472 231 3476 235
rect 984 223 988 227
rect 2760 215 2764 219
rect 496 207 500 211
rect 608 207 612 211
rect 728 207 732 211
rect 856 207 860 211
rect 1488 207 1492 211
rect 1616 207 1620 211
rect 1720 207 1724 211
rect 2944 215 2948 219
rect 3120 215 3124 219
rect 3304 215 3308 219
rect 1976 187 1980 191
rect 2192 187 2196 191
rect 2400 187 2404 191
rect 2600 187 2604 191
rect 2760 187 2764 191
rect 2784 187 2788 191
rect 2944 187 2948 191
rect 2968 187 2972 191
rect 3120 187 3124 191
rect 3144 187 3148 191
rect 3304 187 3308 191
rect 3328 187 3332 191
rect 3496 187 3500 191
rect 416 179 420 183
rect 496 179 500 183
rect 520 179 524 183
rect 608 179 612 183
rect 632 179 636 183
rect 728 179 732 183
rect 752 179 756 183
rect 856 179 860 183
rect 880 179 884 183
rect 1008 179 1012 183
rect 1136 179 1140 183
rect 1264 179 1268 183
rect 1392 179 1396 183
rect 1488 179 1492 183
rect 1512 179 1516 183
rect 1616 179 1620 183
rect 1640 179 1644 183
rect 1720 179 1724 183
rect 1744 179 1748 183
rect 1584 171 1588 175
rect 232 147 236 151
rect 288 147 292 151
rect 320 147 324 151
rect 376 147 380 151
rect 408 147 412 151
rect 464 147 468 151
rect 496 147 500 151
rect 552 147 556 151
rect 584 147 588 151
rect 640 147 644 151
rect 672 147 676 151
rect 728 147 732 151
rect 760 147 764 151
rect 816 147 820 151
rect 848 147 852 151
rect 904 147 908 151
rect 936 147 940 151
rect 992 147 996 151
rect 1024 147 1028 151
rect 1080 147 1084 151
rect 1112 147 1116 151
rect 1200 147 1204 151
rect 1256 147 1260 151
rect 1304 147 1308 151
rect 1360 147 1364 151
rect 1408 147 1412 151
rect 1464 147 1468 151
rect 1520 147 1524 151
rect 1576 147 1580 151
rect 288 123 292 127
rect 376 123 380 127
rect 464 123 468 127
rect 552 123 556 127
rect 640 123 644 127
rect 728 123 732 127
rect 816 123 820 127
rect 904 123 908 127
rect 992 123 996 127
rect 1080 123 1084 127
rect 1256 123 1260 127
rect 1360 123 1364 127
rect 1464 123 1468 127
rect 1576 123 1580 127
rect 1640 147 1644 151
rect 1744 147 1748 151
rect 1808 143 1812 147
rect 1904 143 1908 147
rect 1960 143 1964 147
rect 1992 143 1996 147
rect 2056 143 2060 147
rect 2080 143 2084 147
rect 2136 143 2140 147
rect 2168 143 2172 147
rect 2224 143 2228 147
rect 2280 143 2284 147
rect 2336 143 2340 147
rect 2392 143 2396 147
rect 2504 143 2508 147
rect 2616 143 2620 147
rect 2672 143 2676 147
rect 2728 143 2732 147
rect 2784 143 2788 147
rect 2832 143 2836 147
rect 2912 143 2916 147
rect 2936 143 2940 147
rect 2992 143 2996 147
rect 3032 143 3036 147
rect 3088 143 3092 147
rect 3128 143 3132 147
rect 3184 143 3188 147
rect 3224 143 3228 147
rect 3280 143 3284 147
rect 3320 143 3324 147
rect 3376 143 3380 147
rect 3408 143 3412 147
rect 3464 143 3468 147
rect 3496 143 3500 147
rect 1808 123 1812 127
rect 1584 119 1588 123
rect 1960 119 1964 123
rect 2056 119 2060 123
rect 2136 119 2140 123
rect 2224 119 2228 123
rect 2336 119 2340 123
rect 2672 119 2676 123
rect 2784 119 2788 123
rect 2912 119 2916 123
rect 2992 119 2996 123
rect 3088 119 3092 123
rect 3184 119 3188 123
rect 3280 119 3284 123
rect 3376 119 3380 123
rect 3464 119 3468 123
<< m2 >>
rect 207 3643 213 3644
rect 207 3639 208 3643
rect 212 3642 213 3643
rect 239 3643 245 3644
rect 239 3642 240 3643
rect 212 3640 240 3642
rect 212 3639 213 3640
rect 207 3638 213 3639
rect 239 3639 240 3640
rect 244 3639 245 3643
rect 239 3638 245 3639
rect 295 3643 301 3644
rect 295 3639 296 3643
rect 300 3642 301 3643
rect 327 3643 333 3644
rect 327 3642 328 3643
rect 300 3640 328 3642
rect 300 3639 301 3640
rect 295 3638 301 3639
rect 327 3639 328 3640
rect 332 3639 333 3643
rect 327 3638 333 3639
rect 383 3643 389 3644
rect 383 3639 384 3643
rect 388 3642 389 3643
rect 415 3643 421 3644
rect 415 3642 416 3643
rect 388 3640 416 3642
rect 388 3639 389 3640
rect 383 3638 389 3639
rect 415 3639 416 3640
rect 420 3639 421 3643
rect 415 3638 421 3639
rect 471 3643 477 3644
rect 471 3639 472 3643
rect 476 3642 477 3643
rect 503 3643 509 3644
rect 503 3642 504 3643
rect 476 3640 504 3642
rect 476 3639 477 3640
rect 471 3638 477 3639
rect 503 3639 504 3640
rect 508 3639 509 3643
rect 503 3638 509 3639
rect 559 3643 565 3644
rect 559 3639 560 3643
rect 564 3642 565 3643
rect 591 3643 597 3644
rect 591 3642 592 3643
rect 564 3640 592 3642
rect 564 3639 565 3640
rect 559 3638 565 3639
rect 591 3639 592 3640
rect 596 3639 597 3643
rect 591 3638 597 3639
rect 647 3643 653 3644
rect 647 3639 648 3643
rect 652 3642 653 3643
rect 679 3643 685 3644
rect 679 3642 680 3643
rect 652 3640 680 3642
rect 652 3639 653 3640
rect 647 3638 653 3639
rect 679 3639 680 3640
rect 684 3639 685 3643
rect 679 3638 685 3639
rect 142 3633 148 3634
rect 142 3629 143 3633
rect 147 3629 148 3633
rect 142 3628 148 3629
rect 230 3633 236 3634
rect 230 3629 231 3633
rect 235 3629 236 3633
rect 230 3628 236 3629
rect 318 3633 324 3634
rect 318 3629 319 3633
rect 323 3629 324 3633
rect 318 3628 324 3629
rect 406 3633 412 3634
rect 406 3629 407 3633
rect 411 3629 412 3633
rect 406 3628 412 3629
rect 494 3633 500 3634
rect 494 3629 495 3633
rect 499 3629 500 3633
rect 494 3628 500 3629
rect 582 3633 588 3634
rect 582 3629 583 3633
rect 587 3629 588 3633
rect 582 3628 588 3629
rect 670 3633 676 3634
rect 670 3629 671 3633
rect 675 3629 676 3633
rect 670 3628 676 3629
rect 110 3620 116 3621
rect 1822 3620 1828 3621
rect 110 3616 111 3620
rect 115 3616 116 3620
rect 207 3619 213 3620
rect 207 3618 208 3619
rect 197 3616 208 3618
rect 110 3615 116 3616
rect 207 3615 208 3616
rect 212 3615 213 3619
rect 295 3619 301 3620
rect 295 3618 296 3619
rect 285 3616 296 3618
rect 207 3614 213 3615
rect 295 3615 296 3616
rect 300 3615 301 3619
rect 383 3619 389 3620
rect 383 3618 384 3619
rect 373 3616 384 3618
rect 295 3614 301 3615
rect 383 3615 384 3616
rect 388 3615 389 3619
rect 471 3619 477 3620
rect 471 3618 472 3619
rect 461 3616 472 3618
rect 383 3614 389 3615
rect 471 3615 472 3616
rect 476 3615 477 3619
rect 559 3619 565 3620
rect 559 3618 560 3619
rect 549 3616 560 3618
rect 471 3614 477 3615
rect 559 3615 560 3616
rect 564 3615 565 3619
rect 647 3619 653 3620
rect 647 3618 648 3619
rect 637 3616 648 3618
rect 559 3614 565 3615
rect 647 3615 648 3616
rect 652 3615 653 3619
rect 1822 3616 1823 3620
rect 1827 3616 1828 3620
rect 1822 3615 1828 3616
rect 647 3614 653 3615
rect 110 3603 116 3604
rect 110 3599 111 3603
rect 115 3599 116 3603
rect 110 3598 116 3599
rect 650 3603 656 3604
rect 650 3599 651 3603
rect 655 3602 656 3603
rect 1822 3603 1828 3604
rect 655 3600 681 3602
rect 655 3599 656 3600
rect 650 3598 656 3599
rect 1822 3599 1823 3603
rect 1827 3599 1828 3603
rect 1822 3598 1828 3599
rect 134 3593 140 3594
rect 134 3589 135 3593
rect 139 3589 140 3593
rect 134 3588 140 3589
rect 222 3593 228 3594
rect 222 3589 223 3593
rect 227 3589 228 3593
rect 222 3588 228 3589
rect 310 3593 316 3594
rect 310 3589 311 3593
rect 315 3589 316 3593
rect 310 3588 316 3589
rect 398 3593 404 3594
rect 398 3589 399 3593
rect 403 3589 404 3593
rect 398 3588 404 3589
rect 486 3593 492 3594
rect 486 3589 487 3593
rect 491 3589 492 3593
rect 486 3588 492 3589
rect 574 3593 580 3594
rect 574 3589 575 3593
rect 579 3589 580 3593
rect 574 3588 580 3589
rect 662 3593 668 3594
rect 662 3589 663 3593
rect 667 3589 668 3593
rect 662 3588 668 3589
rect 1546 3571 1552 3572
rect 1546 3567 1547 3571
rect 1551 3570 1552 3571
rect 1551 3568 1710 3570
rect 1551 3567 1552 3568
rect 1546 3566 1552 3567
rect 134 3563 140 3564
rect 134 3559 135 3563
rect 139 3559 140 3563
rect 134 3558 140 3559
rect 286 3563 292 3564
rect 286 3559 287 3563
rect 291 3559 292 3563
rect 286 3558 292 3559
rect 462 3563 468 3564
rect 462 3559 463 3563
rect 467 3559 468 3563
rect 462 3558 468 3559
rect 630 3563 636 3564
rect 630 3559 631 3563
rect 635 3559 636 3563
rect 630 3558 636 3559
rect 790 3563 796 3564
rect 790 3559 791 3563
rect 795 3559 796 3563
rect 790 3558 796 3559
rect 934 3563 940 3564
rect 934 3559 935 3563
rect 939 3559 940 3563
rect 934 3558 940 3559
rect 1070 3563 1076 3564
rect 1070 3559 1071 3563
rect 1075 3559 1076 3563
rect 1070 3558 1076 3559
rect 1190 3563 1196 3564
rect 1190 3559 1191 3563
rect 1195 3559 1196 3563
rect 1190 3558 1196 3559
rect 1310 3563 1316 3564
rect 1310 3559 1311 3563
rect 1315 3559 1316 3563
rect 1310 3558 1316 3559
rect 1422 3563 1428 3564
rect 1422 3559 1423 3563
rect 1427 3559 1428 3563
rect 1422 3558 1428 3559
rect 1526 3563 1532 3564
rect 1526 3559 1527 3563
rect 1531 3559 1532 3563
rect 1526 3558 1532 3559
rect 1638 3563 1644 3564
rect 1638 3559 1639 3563
rect 1643 3559 1644 3563
rect 1638 3558 1644 3559
rect 558 3555 564 3556
rect 110 3553 116 3554
rect 110 3549 111 3553
rect 115 3549 116 3553
rect 558 3551 559 3555
rect 563 3554 564 3555
rect 1708 3554 1710 3568
rect 1726 3563 1732 3564
rect 1726 3559 1727 3563
rect 1731 3559 1732 3563
rect 1726 3558 1732 3559
rect 563 3552 649 3554
rect 1708 3552 1745 3554
rect 1822 3553 1828 3554
rect 563 3551 564 3552
rect 558 3550 564 3551
rect 110 3548 116 3549
rect 1822 3549 1823 3553
rect 1827 3549 1828 3553
rect 1822 3548 1828 3549
rect 279 3539 285 3540
rect 279 3538 280 3539
rect 110 3536 116 3537
rect 197 3536 280 3538
rect 110 3532 111 3536
rect 115 3532 116 3536
rect 279 3535 280 3536
rect 284 3535 285 3539
rect 455 3539 461 3540
rect 455 3538 456 3539
rect 349 3536 456 3538
rect 279 3534 285 3535
rect 455 3535 456 3536
rect 460 3535 461 3539
rect 623 3539 629 3540
rect 623 3538 624 3539
rect 525 3536 624 3538
rect 455 3534 461 3535
rect 623 3535 624 3536
rect 628 3535 629 3539
rect 927 3539 933 3540
rect 927 3538 928 3539
rect 853 3536 928 3538
rect 623 3534 629 3535
rect 927 3535 928 3536
rect 932 3535 933 3539
rect 1063 3539 1069 3540
rect 1063 3538 1064 3539
rect 997 3536 1064 3538
rect 927 3534 933 3535
rect 1063 3535 1064 3536
rect 1068 3535 1069 3539
rect 1183 3539 1189 3540
rect 1183 3538 1184 3539
rect 1133 3536 1184 3538
rect 1063 3534 1069 3535
rect 1183 3535 1184 3536
rect 1188 3535 1189 3539
rect 1303 3539 1309 3540
rect 1303 3538 1304 3539
rect 1253 3536 1304 3538
rect 1183 3534 1189 3535
rect 1303 3535 1304 3536
rect 1308 3535 1309 3539
rect 1415 3539 1421 3540
rect 1415 3538 1416 3539
rect 1373 3536 1416 3538
rect 1303 3534 1309 3535
rect 1415 3535 1416 3536
rect 1420 3535 1421 3539
rect 1519 3539 1525 3540
rect 1519 3538 1520 3539
rect 1485 3536 1520 3538
rect 1415 3534 1421 3535
rect 1519 3535 1520 3536
rect 1524 3535 1525 3539
rect 1631 3539 1637 3540
rect 1631 3538 1632 3539
rect 1589 3536 1632 3538
rect 1519 3534 1525 3535
rect 1631 3535 1632 3536
rect 1636 3535 1637 3539
rect 1719 3539 1725 3540
rect 1719 3538 1720 3539
rect 1701 3536 1720 3538
rect 1631 3534 1637 3535
rect 1719 3535 1720 3536
rect 1724 3535 1725 3539
rect 1719 3534 1725 3535
rect 1822 3536 1828 3537
rect 110 3531 116 3532
rect 1822 3532 1823 3536
rect 1827 3532 1828 3536
rect 1822 3531 1828 3532
rect 142 3523 148 3524
rect 142 3519 143 3523
rect 147 3519 148 3523
rect 142 3518 148 3519
rect 294 3523 300 3524
rect 294 3519 295 3523
rect 299 3519 300 3523
rect 294 3518 300 3519
rect 470 3523 476 3524
rect 470 3519 471 3523
rect 475 3519 476 3523
rect 470 3518 476 3519
rect 638 3523 644 3524
rect 638 3519 639 3523
rect 643 3519 644 3523
rect 638 3518 644 3519
rect 798 3523 804 3524
rect 798 3519 799 3523
rect 803 3519 804 3523
rect 798 3518 804 3519
rect 942 3523 948 3524
rect 942 3519 943 3523
rect 947 3519 948 3523
rect 942 3518 948 3519
rect 1078 3523 1084 3524
rect 1078 3519 1079 3523
rect 1083 3519 1084 3523
rect 1078 3518 1084 3519
rect 1198 3523 1204 3524
rect 1198 3519 1199 3523
rect 1203 3519 1204 3523
rect 1198 3518 1204 3519
rect 1318 3523 1324 3524
rect 1318 3519 1319 3523
rect 1323 3519 1324 3523
rect 1318 3518 1324 3519
rect 1430 3523 1436 3524
rect 1430 3519 1431 3523
rect 1435 3519 1436 3523
rect 1430 3518 1436 3519
rect 1534 3523 1540 3524
rect 1534 3519 1535 3523
rect 1539 3519 1540 3523
rect 1534 3518 1540 3519
rect 1646 3523 1652 3524
rect 1646 3519 1647 3523
rect 1651 3519 1652 3523
rect 1646 3518 1652 3519
rect 1734 3523 1740 3524
rect 1734 3519 1735 3523
rect 1739 3519 1740 3523
rect 1734 3518 1740 3519
rect 806 3515 812 3516
rect 151 3511 157 3512
rect 151 3507 152 3511
rect 156 3510 157 3511
rect 166 3511 172 3512
rect 166 3510 167 3511
rect 156 3508 167 3510
rect 156 3507 157 3508
rect 151 3506 157 3507
rect 166 3507 167 3508
rect 171 3507 172 3511
rect 166 3506 172 3507
rect 279 3511 285 3512
rect 279 3507 280 3511
rect 284 3510 285 3511
rect 303 3511 309 3512
rect 303 3510 304 3511
rect 284 3508 304 3510
rect 284 3507 285 3508
rect 279 3506 285 3507
rect 303 3507 304 3508
rect 308 3507 309 3511
rect 303 3506 309 3507
rect 455 3511 461 3512
rect 455 3507 456 3511
rect 460 3510 461 3511
rect 479 3511 485 3512
rect 479 3510 480 3511
rect 460 3508 480 3510
rect 460 3507 461 3508
rect 455 3506 461 3507
rect 479 3507 480 3508
rect 484 3507 485 3511
rect 479 3506 485 3507
rect 623 3511 629 3512
rect 623 3507 624 3511
rect 628 3510 629 3511
rect 647 3511 653 3512
rect 647 3510 648 3511
rect 628 3508 648 3510
rect 628 3507 629 3508
rect 623 3506 629 3507
rect 647 3507 648 3508
rect 652 3507 653 3511
rect 806 3511 807 3515
rect 811 3514 812 3515
rect 811 3513 813 3514
rect 806 3510 808 3511
rect 807 3509 808 3510
rect 812 3509 813 3513
rect 807 3508 813 3509
rect 927 3511 933 3512
rect 647 3506 653 3507
rect 927 3507 928 3511
rect 932 3510 933 3511
rect 951 3511 957 3512
rect 951 3510 952 3511
rect 932 3508 952 3510
rect 932 3507 933 3508
rect 927 3506 933 3507
rect 951 3507 952 3508
rect 956 3507 957 3511
rect 951 3506 957 3507
rect 1063 3511 1069 3512
rect 1063 3507 1064 3511
rect 1068 3510 1069 3511
rect 1087 3511 1093 3512
rect 1087 3510 1088 3511
rect 1068 3508 1088 3510
rect 1068 3507 1069 3508
rect 1063 3506 1069 3507
rect 1087 3507 1088 3508
rect 1092 3507 1093 3511
rect 1087 3506 1093 3507
rect 1183 3511 1189 3512
rect 1183 3507 1184 3511
rect 1188 3510 1189 3511
rect 1207 3511 1213 3512
rect 1207 3510 1208 3511
rect 1188 3508 1208 3510
rect 1188 3507 1189 3508
rect 1183 3506 1189 3507
rect 1207 3507 1208 3508
rect 1212 3507 1213 3511
rect 1207 3506 1213 3507
rect 1303 3511 1309 3512
rect 1303 3507 1304 3511
rect 1308 3510 1309 3511
rect 1327 3511 1333 3512
rect 1327 3510 1328 3511
rect 1308 3508 1328 3510
rect 1308 3507 1309 3508
rect 1303 3506 1309 3507
rect 1327 3507 1328 3508
rect 1332 3507 1333 3511
rect 1327 3506 1333 3507
rect 1415 3511 1421 3512
rect 1415 3507 1416 3511
rect 1420 3510 1421 3511
rect 1439 3511 1445 3512
rect 1439 3510 1440 3511
rect 1420 3508 1440 3510
rect 1420 3507 1421 3508
rect 1415 3506 1421 3507
rect 1439 3507 1440 3508
rect 1444 3507 1445 3511
rect 1439 3506 1445 3507
rect 1519 3511 1525 3512
rect 1519 3507 1520 3511
rect 1524 3510 1525 3511
rect 1543 3511 1549 3512
rect 1543 3510 1544 3511
rect 1524 3508 1544 3510
rect 1524 3507 1525 3508
rect 1519 3506 1525 3507
rect 1543 3507 1544 3508
rect 1548 3507 1549 3511
rect 1543 3506 1549 3507
rect 1631 3511 1637 3512
rect 1631 3507 1632 3511
rect 1636 3510 1637 3511
rect 1655 3511 1661 3512
rect 1655 3510 1656 3511
rect 1636 3508 1656 3510
rect 1636 3507 1637 3508
rect 1631 3506 1637 3507
rect 1655 3507 1656 3508
rect 1660 3507 1661 3511
rect 1655 3506 1661 3507
rect 1719 3511 1725 3512
rect 1719 3507 1720 3511
rect 1724 3510 1725 3511
rect 1743 3511 1749 3512
rect 1743 3510 1744 3511
rect 1724 3508 1744 3510
rect 1724 3507 1725 3508
rect 1719 3506 1725 3507
rect 1743 3507 1744 3508
rect 1748 3507 1749 3511
rect 1743 3506 1749 3507
rect 158 3499 165 3500
rect 158 3495 159 3499
rect 164 3495 165 3499
rect 158 3494 165 3495
rect 239 3499 245 3500
rect 239 3495 240 3499
rect 244 3498 245 3499
rect 335 3499 341 3500
rect 335 3498 336 3499
rect 244 3496 336 3498
rect 244 3495 245 3496
rect 239 3494 245 3495
rect 335 3495 336 3496
rect 340 3495 341 3499
rect 335 3494 341 3495
rect 415 3499 421 3500
rect 415 3495 416 3499
rect 420 3498 421 3499
rect 503 3499 509 3500
rect 503 3498 504 3499
rect 420 3496 504 3498
rect 420 3495 421 3496
rect 415 3494 421 3495
rect 503 3495 504 3496
rect 508 3495 509 3499
rect 503 3494 509 3495
rect 583 3499 589 3500
rect 583 3495 584 3499
rect 588 3498 589 3499
rect 663 3499 669 3500
rect 663 3498 664 3499
rect 588 3496 664 3498
rect 588 3495 589 3496
rect 583 3494 589 3495
rect 663 3495 664 3496
rect 668 3495 669 3499
rect 663 3494 669 3495
rect 815 3499 821 3500
rect 815 3495 816 3499
rect 820 3498 821 3499
rect 878 3499 884 3500
rect 878 3498 879 3499
rect 820 3496 879 3498
rect 820 3495 821 3496
rect 815 3494 821 3495
rect 878 3495 879 3496
rect 883 3495 884 3499
rect 878 3494 884 3495
rect 887 3499 893 3500
rect 887 3495 888 3499
rect 892 3498 893 3499
rect 959 3499 965 3500
rect 959 3498 960 3499
rect 892 3496 960 3498
rect 892 3495 893 3496
rect 887 3494 893 3495
rect 959 3495 960 3496
rect 964 3495 965 3499
rect 959 3494 965 3495
rect 1015 3499 1021 3500
rect 1015 3495 1016 3499
rect 1020 3498 1021 3499
rect 1095 3499 1101 3500
rect 1095 3498 1096 3499
rect 1020 3496 1096 3498
rect 1020 3495 1021 3496
rect 1015 3494 1021 3495
rect 1095 3495 1096 3496
rect 1100 3495 1101 3499
rect 1095 3494 1101 3495
rect 1146 3499 1152 3500
rect 1146 3495 1147 3499
rect 1151 3498 1152 3499
rect 1215 3499 1221 3500
rect 1215 3498 1216 3499
rect 1151 3496 1216 3498
rect 1151 3495 1152 3496
rect 1146 3494 1152 3495
rect 1215 3495 1216 3496
rect 1220 3495 1221 3499
rect 1215 3494 1221 3495
rect 1271 3499 1277 3500
rect 1271 3495 1272 3499
rect 1276 3498 1277 3499
rect 1327 3499 1333 3500
rect 1327 3498 1328 3499
rect 1276 3496 1328 3498
rect 1276 3495 1277 3496
rect 1271 3494 1277 3495
rect 1327 3495 1328 3496
rect 1332 3495 1333 3499
rect 1327 3494 1333 3495
rect 1383 3499 1389 3500
rect 1383 3495 1384 3499
rect 1388 3498 1389 3499
rect 1439 3499 1445 3500
rect 1439 3498 1440 3499
rect 1388 3496 1440 3498
rect 1388 3495 1389 3496
rect 1383 3494 1389 3495
rect 1439 3495 1440 3496
rect 1444 3495 1445 3499
rect 1439 3494 1445 3495
rect 1543 3499 1552 3500
rect 1543 3495 1544 3499
rect 1551 3495 1552 3499
rect 1543 3494 1552 3495
rect 1599 3499 1605 3500
rect 1599 3495 1600 3499
rect 1604 3498 1605 3499
rect 1655 3499 1661 3500
rect 1655 3498 1656 3499
rect 1604 3496 1656 3498
rect 1604 3495 1605 3496
rect 1599 3494 1605 3495
rect 1655 3495 1656 3496
rect 1660 3495 1661 3499
rect 1655 3494 1661 3495
rect 1711 3499 1717 3500
rect 1711 3495 1712 3499
rect 1716 3498 1717 3499
rect 1743 3499 1749 3500
rect 1743 3498 1744 3499
rect 1716 3496 1744 3498
rect 1716 3495 1717 3496
rect 1711 3494 1717 3495
rect 1743 3495 1744 3496
rect 1748 3495 1749 3499
rect 1743 3494 1749 3495
rect 1807 3495 1813 3496
rect 1807 3491 1808 3495
rect 1812 3494 1813 3495
rect 1903 3495 1909 3496
rect 1903 3494 1904 3495
rect 1812 3492 1904 3494
rect 1812 3491 1813 3492
rect 1807 3490 1813 3491
rect 1903 3491 1904 3492
rect 1908 3491 1909 3495
rect 1903 3490 1909 3491
rect 1959 3495 1965 3496
rect 1959 3491 1960 3495
rect 1964 3494 1965 3495
rect 1991 3495 1997 3496
rect 1991 3494 1992 3495
rect 1964 3492 1992 3494
rect 1964 3491 1965 3492
rect 1959 3490 1965 3491
rect 1991 3491 1992 3492
rect 1996 3491 1997 3495
rect 1991 3490 1997 3491
rect 2055 3495 2061 3496
rect 2055 3491 2056 3495
rect 2060 3494 2061 3495
rect 2079 3495 2085 3496
rect 2079 3494 2080 3495
rect 2060 3492 2080 3494
rect 2060 3491 2061 3492
rect 2055 3490 2061 3491
rect 2079 3491 2080 3492
rect 2084 3491 2085 3495
rect 2079 3490 2085 3491
rect 2135 3495 2141 3496
rect 2135 3491 2136 3495
rect 2140 3494 2141 3495
rect 2167 3495 2173 3496
rect 2167 3494 2168 3495
rect 2140 3492 2168 3494
rect 2140 3491 2141 3492
rect 2135 3490 2141 3491
rect 2167 3491 2168 3492
rect 2172 3491 2173 3495
rect 2167 3490 2173 3491
rect 150 3489 156 3490
rect 150 3485 151 3489
rect 155 3485 156 3489
rect 150 3484 156 3485
rect 326 3489 332 3490
rect 326 3485 327 3489
rect 331 3485 332 3489
rect 326 3484 332 3485
rect 494 3489 500 3490
rect 494 3485 495 3489
rect 499 3485 500 3489
rect 494 3484 500 3485
rect 654 3489 660 3490
rect 654 3485 655 3489
rect 659 3485 660 3489
rect 654 3484 660 3485
rect 806 3489 812 3490
rect 806 3485 807 3489
rect 811 3485 812 3489
rect 806 3484 812 3485
rect 950 3489 956 3490
rect 950 3485 951 3489
rect 955 3485 956 3489
rect 950 3484 956 3485
rect 1086 3489 1092 3490
rect 1086 3485 1087 3489
rect 1091 3485 1092 3489
rect 1086 3484 1092 3485
rect 1206 3489 1212 3490
rect 1206 3485 1207 3489
rect 1211 3485 1212 3489
rect 1206 3484 1212 3485
rect 1318 3489 1324 3490
rect 1318 3485 1319 3489
rect 1323 3485 1324 3489
rect 1318 3484 1324 3485
rect 1430 3489 1436 3490
rect 1430 3485 1431 3489
rect 1435 3485 1436 3489
rect 1430 3484 1436 3485
rect 1534 3489 1540 3490
rect 1534 3485 1535 3489
rect 1539 3485 1540 3489
rect 1534 3484 1540 3485
rect 1646 3489 1652 3490
rect 1646 3485 1647 3489
rect 1651 3485 1652 3489
rect 1646 3484 1652 3485
rect 1734 3489 1740 3490
rect 1734 3485 1735 3489
rect 1739 3485 1740 3489
rect 1734 3484 1740 3485
rect 1894 3485 1900 3486
rect 1894 3481 1895 3485
rect 1899 3481 1900 3485
rect 1894 3480 1900 3481
rect 1982 3485 1988 3486
rect 1982 3481 1983 3485
rect 1987 3481 1988 3485
rect 1982 3480 1988 3481
rect 2070 3485 2076 3486
rect 2070 3481 2071 3485
rect 2075 3481 2076 3485
rect 2070 3480 2076 3481
rect 2158 3485 2164 3486
rect 2158 3481 2159 3485
rect 2163 3481 2164 3485
rect 2158 3480 2164 3481
rect 110 3476 116 3477
rect 1822 3476 1828 3477
rect 110 3472 111 3476
rect 115 3472 116 3476
rect 239 3475 245 3476
rect 239 3474 240 3475
rect 205 3472 240 3474
rect 110 3471 116 3472
rect 239 3471 240 3472
rect 244 3471 245 3475
rect 415 3475 421 3476
rect 415 3474 416 3475
rect 381 3472 416 3474
rect 239 3470 245 3471
rect 415 3471 416 3472
rect 420 3471 421 3475
rect 583 3475 589 3476
rect 583 3474 584 3475
rect 549 3472 584 3474
rect 415 3470 421 3471
rect 583 3471 584 3472
rect 588 3471 589 3475
rect 887 3475 893 3476
rect 887 3474 888 3475
rect 861 3472 888 3474
rect 583 3470 589 3471
rect 887 3471 888 3472
rect 892 3471 893 3475
rect 1015 3475 1021 3476
rect 1015 3474 1016 3475
rect 1005 3472 1016 3474
rect 887 3470 893 3471
rect 1015 3471 1016 3472
rect 1020 3471 1021 3475
rect 1146 3475 1152 3476
rect 1146 3474 1147 3475
rect 1141 3472 1147 3474
rect 1015 3470 1021 3471
rect 1146 3471 1147 3472
rect 1151 3471 1152 3475
rect 1271 3475 1277 3476
rect 1271 3474 1272 3475
rect 1261 3472 1272 3474
rect 1146 3470 1152 3471
rect 1271 3471 1272 3472
rect 1276 3471 1277 3475
rect 1383 3475 1389 3476
rect 1383 3474 1384 3475
rect 1373 3472 1384 3474
rect 1271 3470 1277 3471
rect 1383 3471 1384 3472
rect 1388 3471 1389 3475
rect 1599 3475 1605 3476
rect 1599 3474 1600 3475
rect 1589 3472 1600 3474
rect 1383 3470 1389 3471
rect 1394 3471 1400 3472
rect 1394 3467 1395 3471
rect 1399 3470 1400 3471
rect 1599 3471 1600 3472
rect 1604 3471 1605 3475
rect 1711 3475 1717 3476
rect 1711 3474 1712 3475
rect 1701 3472 1712 3474
rect 1599 3470 1605 3471
rect 1711 3471 1712 3472
rect 1716 3471 1717 3475
rect 1807 3475 1813 3476
rect 1807 3474 1808 3475
rect 1789 3472 1808 3474
rect 1711 3470 1717 3471
rect 1807 3471 1808 3472
rect 1812 3471 1813 3475
rect 1822 3472 1823 3476
rect 1827 3472 1828 3476
rect 1822 3471 1828 3472
rect 1862 3472 1868 3473
rect 3574 3472 3580 3473
rect 1807 3470 1813 3471
rect 1399 3468 1449 3470
rect 1862 3468 1863 3472
rect 1867 3468 1868 3472
rect 1959 3471 1965 3472
rect 1959 3470 1960 3471
rect 1949 3468 1960 3470
rect 1399 3467 1400 3468
rect 1862 3467 1868 3468
rect 1959 3467 1960 3468
rect 1964 3467 1965 3471
rect 2055 3471 2061 3472
rect 2055 3470 2056 3471
rect 2037 3468 2056 3470
rect 1394 3466 1400 3467
rect 1959 3466 1965 3467
rect 2055 3467 2056 3468
rect 2060 3467 2061 3471
rect 2135 3471 2141 3472
rect 2135 3470 2136 3471
rect 2125 3468 2136 3470
rect 2055 3466 2061 3467
rect 2135 3467 2136 3468
rect 2140 3467 2141 3471
rect 3574 3468 3575 3472
rect 3579 3468 3580 3472
rect 3574 3467 3580 3468
rect 2135 3466 2141 3467
rect 110 3459 116 3460
rect 110 3455 111 3459
rect 115 3455 116 3459
rect 110 3454 116 3455
rect 562 3459 568 3460
rect 562 3455 563 3459
rect 567 3458 568 3459
rect 1822 3459 1828 3460
rect 567 3456 665 3458
rect 567 3455 568 3456
rect 562 3454 568 3455
rect 1822 3455 1823 3459
rect 1827 3455 1828 3459
rect 1822 3454 1828 3455
rect 1862 3455 1868 3456
rect 1862 3451 1863 3455
rect 1867 3451 1868 3455
rect 1862 3450 1868 3451
rect 2138 3455 2144 3456
rect 2138 3451 2139 3455
rect 2143 3454 2144 3455
rect 3574 3455 3580 3456
rect 2143 3452 2169 3454
rect 2143 3451 2144 3452
rect 2138 3450 2144 3451
rect 3574 3451 3575 3455
rect 3579 3451 3580 3455
rect 3574 3450 3580 3451
rect 142 3449 148 3450
rect 142 3445 143 3449
rect 147 3445 148 3449
rect 142 3444 148 3445
rect 318 3449 324 3450
rect 318 3445 319 3449
rect 323 3445 324 3449
rect 318 3444 324 3445
rect 486 3449 492 3450
rect 486 3445 487 3449
rect 491 3445 492 3449
rect 486 3444 492 3445
rect 646 3449 652 3450
rect 646 3445 647 3449
rect 651 3445 652 3449
rect 646 3444 652 3445
rect 798 3449 804 3450
rect 798 3445 799 3449
rect 803 3445 804 3449
rect 798 3444 804 3445
rect 942 3449 948 3450
rect 942 3445 943 3449
rect 947 3445 948 3449
rect 942 3444 948 3445
rect 1078 3449 1084 3450
rect 1078 3445 1079 3449
rect 1083 3445 1084 3449
rect 1078 3444 1084 3445
rect 1198 3449 1204 3450
rect 1198 3445 1199 3449
rect 1203 3445 1204 3449
rect 1198 3444 1204 3445
rect 1310 3449 1316 3450
rect 1310 3445 1311 3449
rect 1315 3445 1316 3449
rect 1310 3444 1316 3445
rect 1422 3449 1428 3450
rect 1422 3445 1423 3449
rect 1427 3445 1428 3449
rect 1422 3444 1428 3445
rect 1526 3449 1532 3450
rect 1526 3445 1527 3449
rect 1531 3445 1532 3449
rect 1526 3444 1532 3445
rect 1638 3449 1644 3450
rect 1638 3445 1639 3449
rect 1643 3445 1644 3449
rect 1638 3444 1644 3445
rect 1726 3449 1732 3450
rect 1726 3445 1727 3449
rect 1731 3445 1732 3449
rect 1726 3444 1732 3445
rect 1886 3445 1892 3446
rect 1886 3441 1887 3445
rect 1891 3441 1892 3445
rect 1886 3440 1892 3441
rect 1974 3445 1980 3446
rect 1974 3441 1975 3445
rect 1979 3441 1980 3445
rect 1974 3440 1980 3441
rect 2062 3445 2068 3446
rect 2062 3441 2063 3445
rect 2067 3441 2068 3445
rect 2062 3440 2068 3441
rect 2150 3445 2156 3446
rect 2150 3441 2151 3445
rect 2155 3441 2156 3445
rect 2150 3440 2156 3441
rect 1914 3439 1920 3440
rect 1914 3435 1915 3439
rect 1919 3438 1920 3439
rect 1919 3436 2001 3438
rect 1919 3435 1920 3436
rect 1914 3434 1920 3435
rect 1999 3430 2001 3436
rect 2138 3431 2144 3432
rect 2138 3430 2139 3431
rect 1999 3428 2139 3430
rect 214 3427 220 3428
rect 214 3423 215 3427
rect 219 3423 220 3427
rect 214 3422 220 3423
rect 430 3427 436 3428
rect 430 3423 431 3427
rect 435 3423 436 3427
rect 430 3422 436 3423
rect 638 3427 644 3428
rect 638 3423 639 3427
rect 643 3423 644 3427
rect 638 3422 644 3423
rect 846 3427 852 3428
rect 846 3423 847 3427
rect 851 3423 852 3427
rect 846 3422 852 3423
rect 1038 3427 1044 3428
rect 1038 3423 1039 3427
rect 1043 3423 1044 3427
rect 1038 3422 1044 3423
rect 1222 3427 1228 3428
rect 1222 3423 1223 3427
rect 1227 3423 1228 3427
rect 1222 3422 1228 3423
rect 1398 3427 1404 3428
rect 1398 3423 1399 3427
rect 1403 3423 1404 3427
rect 1398 3422 1404 3423
rect 1566 3427 1572 3428
rect 1566 3423 1567 3427
rect 1571 3423 1572 3427
rect 1566 3422 1572 3423
rect 1726 3427 1732 3428
rect 1726 3423 1727 3427
rect 1731 3423 1732 3427
rect 2138 3427 2139 3428
rect 2143 3427 2144 3431
rect 2138 3426 2144 3427
rect 1726 3422 1732 3423
rect 1886 3423 1892 3424
rect 738 3419 744 3420
rect 110 3417 116 3418
rect 110 3413 111 3417
rect 115 3413 116 3417
rect 738 3415 739 3419
rect 743 3418 744 3419
rect 1646 3419 1652 3420
rect 743 3416 865 3418
rect 743 3415 744 3416
rect 738 3414 744 3415
rect 1646 3415 1647 3419
rect 1651 3418 1652 3419
rect 1886 3419 1887 3423
rect 1891 3419 1892 3423
rect 1886 3418 1892 3419
rect 1990 3423 1996 3424
rect 1990 3419 1991 3423
rect 1995 3419 1996 3423
rect 1990 3418 1996 3419
rect 2118 3423 2124 3424
rect 2118 3419 2119 3423
rect 2123 3419 2124 3423
rect 2118 3418 2124 3419
rect 2254 3423 2260 3424
rect 2254 3419 2255 3423
rect 2259 3419 2260 3423
rect 2254 3418 2260 3419
rect 2390 3423 2396 3424
rect 2390 3419 2391 3423
rect 2395 3419 2396 3423
rect 2390 3418 2396 3419
rect 2526 3423 2532 3424
rect 2526 3419 2527 3423
rect 2531 3419 2532 3423
rect 2526 3418 2532 3419
rect 2654 3423 2660 3424
rect 2654 3419 2655 3423
rect 2659 3419 2660 3423
rect 2654 3418 2660 3419
rect 2782 3423 2788 3424
rect 2782 3419 2783 3423
rect 2787 3419 2788 3423
rect 2782 3418 2788 3419
rect 2918 3423 2924 3424
rect 2918 3419 2919 3423
rect 2923 3419 2924 3423
rect 2918 3418 2924 3419
rect 3054 3423 3060 3424
rect 3054 3419 3055 3423
rect 3059 3419 3060 3423
rect 3054 3418 3060 3419
rect 1651 3416 1745 3418
rect 1822 3417 1828 3418
rect 1651 3415 1652 3416
rect 1646 3414 1652 3415
rect 110 3412 116 3413
rect 1822 3413 1823 3417
rect 1827 3413 1828 3417
rect 2322 3415 2328 3416
rect 1822 3412 1828 3413
rect 1862 3413 1868 3414
rect 1862 3409 1863 3413
rect 1867 3409 1868 3413
rect 2322 3411 2323 3415
rect 2327 3414 2328 3415
rect 2327 3412 2409 3414
rect 3574 3413 3580 3414
rect 2327 3411 2328 3412
rect 2322 3410 2328 3411
rect 1862 3408 1868 3409
rect 3574 3409 3575 3413
rect 3579 3409 3580 3413
rect 3574 3408 3580 3409
rect 423 3403 429 3404
rect 423 3402 424 3403
rect 110 3400 116 3401
rect 277 3400 424 3402
rect 110 3396 111 3400
rect 115 3396 116 3400
rect 423 3399 424 3400
rect 428 3399 429 3403
rect 631 3403 637 3404
rect 631 3402 632 3403
rect 493 3400 632 3402
rect 423 3398 429 3399
rect 631 3399 632 3400
rect 636 3399 637 3403
rect 839 3403 845 3404
rect 839 3402 840 3403
rect 701 3400 840 3402
rect 631 3398 637 3399
rect 839 3399 840 3400
rect 844 3399 845 3403
rect 1215 3403 1221 3404
rect 1215 3402 1216 3403
rect 1101 3400 1216 3402
rect 839 3398 845 3399
rect 1215 3399 1216 3400
rect 1220 3399 1221 3403
rect 1391 3403 1397 3404
rect 1391 3402 1392 3403
rect 1285 3400 1392 3402
rect 1215 3398 1221 3399
rect 1391 3399 1392 3400
rect 1396 3399 1397 3403
rect 1559 3403 1565 3404
rect 1559 3402 1560 3403
rect 1461 3400 1560 3402
rect 1391 3398 1397 3399
rect 1559 3399 1560 3400
rect 1564 3399 1565 3403
rect 1719 3403 1725 3404
rect 1719 3402 1720 3403
rect 1629 3400 1720 3402
rect 1559 3398 1565 3399
rect 1719 3399 1720 3400
rect 1724 3399 1725 3403
rect 1719 3398 1725 3399
rect 1822 3400 1828 3401
rect 110 3395 116 3396
rect 1822 3396 1823 3400
rect 1827 3396 1828 3400
rect 1954 3399 1960 3400
rect 1954 3398 1955 3399
rect 1822 3395 1828 3396
rect 1862 3396 1868 3397
rect 1949 3396 1955 3398
rect 1862 3392 1863 3396
rect 1867 3392 1868 3396
rect 1954 3395 1955 3396
rect 1959 3395 1960 3399
rect 2111 3399 2117 3400
rect 2111 3398 2112 3399
rect 2053 3396 2112 3398
rect 1954 3394 1960 3395
rect 2111 3395 2112 3396
rect 2116 3395 2117 3399
rect 2247 3399 2253 3400
rect 2247 3398 2248 3399
rect 2181 3396 2248 3398
rect 2111 3394 2117 3395
rect 2247 3395 2248 3396
rect 2252 3395 2253 3399
rect 2383 3399 2389 3400
rect 2383 3398 2384 3399
rect 2317 3396 2384 3398
rect 2247 3394 2253 3395
rect 2383 3395 2384 3396
rect 2388 3395 2389 3399
rect 2647 3399 2653 3400
rect 2647 3398 2648 3399
rect 2589 3396 2648 3398
rect 2383 3394 2389 3395
rect 2647 3395 2648 3396
rect 2652 3395 2653 3399
rect 2775 3399 2781 3400
rect 2775 3398 2776 3399
rect 2717 3396 2776 3398
rect 2647 3394 2653 3395
rect 2775 3395 2776 3396
rect 2780 3395 2781 3399
rect 2911 3399 2917 3400
rect 2911 3398 2912 3399
rect 2845 3396 2912 3398
rect 2775 3394 2781 3395
rect 2911 3395 2912 3396
rect 2916 3395 2917 3399
rect 3047 3399 3053 3400
rect 3047 3398 3048 3399
rect 2981 3396 3048 3398
rect 2911 3394 2917 3395
rect 3047 3395 3048 3396
rect 3052 3395 3053 3399
rect 3122 3399 3128 3400
rect 3122 3398 3123 3399
rect 3117 3396 3123 3398
rect 3047 3394 3053 3395
rect 3122 3395 3123 3396
rect 3127 3395 3128 3399
rect 3122 3394 3128 3395
rect 3574 3396 3580 3397
rect 1862 3391 1868 3392
rect 3574 3392 3575 3396
rect 3579 3392 3580 3396
rect 3574 3391 3580 3392
rect 222 3387 228 3388
rect 222 3383 223 3387
rect 227 3383 228 3387
rect 222 3382 228 3383
rect 438 3387 444 3388
rect 438 3383 439 3387
rect 443 3383 444 3387
rect 438 3382 444 3383
rect 646 3387 652 3388
rect 646 3383 647 3387
rect 651 3383 652 3387
rect 646 3382 652 3383
rect 854 3387 860 3388
rect 854 3383 855 3387
rect 859 3383 860 3387
rect 854 3382 860 3383
rect 1046 3387 1052 3388
rect 1046 3383 1047 3387
rect 1051 3383 1052 3387
rect 1046 3382 1052 3383
rect 1230 3387 1236 3388
rect 1230 3383 1231 3387
rect 1235 3383 1236 3387
rect 1230 3382 1236 3383
rect 1406 3387 1412 3388
rect 1406 3383 1407 3387
rect 1411 3383 1412 3387
rect 1406 3382 1412 3383
rect 1574 3387 1580 3388
rect 1574 3383 1575 3387
rect 1579 3383 1580 3387
rect 1574 3382 1580 3383
rect 1734 3387 1740 3388
rect 1734 3383 1735 3387
rect 1739 3383 1740 3387
rect 1734 3382 1740 3383
rect 1894 3383 1900 3384
rect 1894 3379 1895 3383
rect 1899 3379 1900 3383
rect 1894 3378 1900 3379
rect 1998 3383 2004 3384
rect 1998 3379 1999 3383
rect 2003 3379 2004 3383
rect 1998 3378 2004 3379
rect 2126 3383 2132 3384
rect 2126 3379 2127 3383
rect 2131 3379 2132 3383
rect 2126 3378 2132 3379
rect 2262 3383 2268 3384
rect 2262 3379 2263 3383
rect 2267 3379 2268 3383
rect 2262 3378 2268 3379
rect 2398 3383 2404 3384
rect 2398 3379 2399 3383
rect 2403 3379 2404 3383
rect 2398 3378 2404 3379
rect 2534 3383 2540 3384
rect 2534 3379 2535 3383
rect 2539 3379 2540 3383
rect 2534 3378 2540 3379
rect 2662 3383 2668 3384
rect 2662 3379 2663 3383
rect 2667 3379 2668 3383
rect 2662 3378 2668 3379
rect 2790 3383 2796 3384
rect 2790 3379 2791 3383
rect 2795 3379 2796 3383
rect 2790 3378 2796 3379
rect 2926 3383 2932 3384
rect 2926 3379 2927 3383
rect 2931 3379 2932 3383
rect 2926 3378 2932 3379
rect 3062 3383 3068 3384
rect 3062 3379 3063 3383
rect 3067 3379 3068 3383
rect 3062 3378 3068 3379
rect 231 3375 240 3376
rect 231 3371 232 3375
rect 239 3371 240 3375
rect 231 3370 240 3371
rect 423 3375 429 3376
rect 423 3371 424 3375
rect 428 3374 429 3375
rect 447 3375 453 3376
rect 447 3374 448 3375
rect 428 3372 448 3374
rect 428 3371 429 3372
rect 423 3370 429 3371
rect 447 3371 448 3372
rect 452 3371 453 3375
rect 447 3370 453 3371
rect 631 3375 637 3376
rect 631 3371 632 3375
rect 636 3374 637 3375
rect 655 3375 661 3376
rect 655 3374 656 3375
rect 636 3372 656 3374
rect 636 3371 637 3372
rect 631 3370 637 3371
rect 655 3371 656 3372
rect 660 3371 661 3375
rect 655 3370 661 3371
rect 839 3375 845 3376
rect 839 3371 840 3375
rect 844 3374 845 3375
rect 863 3375 869 3376
rect 863 3374 864 3375
rect 844 3372 864 3374
rect 844 3371 845 3372
rect 839 3370 845 3371
rect 863 3371 864 3372
rect 868 3371 869 3375
rect 863 3370 869 3371
rect 1055 3375 1061 3376
rect 1055 3371 1056 3375
rect 1060 3374 1061 3375
rect 1206 3375 1212 3376
rect 1206 3374 1207 3375
rect 1060 3372 1207 3374
rect 1060 3371 1061 3372
rect 1055 3370 1061 3371
rect 1206 3371 1207 3372
rect 1211 3371 1212 3375
rect 1206 3370 1212 3371
rect 1215 3375 1221 3376
rect 1215 3371 1216 3375
rect 1220 3374 1221 3375
rect 1239 3375 1245 3376
rect 1239 3374 1240 3375
rect 1220 3372 1240 3374
rect 1220 3371 1221 3372
rect 1215 3370 1221 3371
rect 1239 3371 1240 3372
rect 1244 3371 1245 3375
rect 1239 3370 1245 3371
rect 1391 3375 1397 3376
rect 1391 3371 1392 3375
rect 1396 3374 1397 3375
rect 1415 3375 1421 3376
rect 1415 3374 1416 3375
rect 1396 3372 1416 3374
rect 1396 3371 1397 3372
rect 1391 3370 1397 3371
rect 1415 3371 1416 3372
rect 1420 3371 1421 3375
rect 1415 3370 1421 3371
rect 1559 3375 1565 3376
rect 1559 3371 1560 3375
rect 1564 3374 1565 3375
rect 1583 3375 1589 3376
rect 1583 3374 1584 3375
rect 1564 3372 1584 3374
rect 1564 3371 1565 3372
rect 1559 3370 1565 3371
rect 1583 3371 1584 3372
rect 1588 3371 1589 3375
rect 1583 3370 1589 3371
rect 1719 3375 1725 3376
rect 1719 3371 1720 3375
rect 1724 3374 1725 3375
rect 1743 3375 1749 3376
rect 1743 3374 1744 3375
rect 1724 3372 1744 3374
rect 1724 3371 1725 3372
rect 1719 3370 1725 3371
rect 1743 3371 1744 3372
rect 1748 3371 1749 3375
rect 1743 3370 1749 3371
rect 1903 3371 1909 3372
rect 1903 3367 1904 3371
rect 1908 3370 1909 3371
rect 1914 3371 1920 3372
rect 1914 3370 1915 3371
rect 1908 3368 1915 3370
rect 1908 3367 1909 3368
rect 1903 3366 1909 3367
rect 1914 3367 1915 3368
rect 1919 3367 1920 3371
rect 1914 3366 1920 3367
rect 1954 3371 1960 3372
rect 1954 3367 1955 3371
rect 1959 3370 1960 3371
rect 2007 3371 2013 3372
rect 2007 3370 2008 3371
rect 1959 3368 2008 3370
rect 1959 3367 1960 3368
rect 1954 3366 1960 3367
rect 2007 3367 2008 3368
rect 2012 3367 2013 3371
rect 2007 3366 2013 3367
rect 2111 3371 2117 3372
rect 2111 3367 2112 3371
rect 2116 3370 2117 3371
rect 2135 3371 2141 3372
rect 2135 3370 2136 3371
rect 2116 3368 2136 3370
rect 2116 3367 2117 3368
rect 2111 3366 2117 3367
rect 2135 3367 2136 3368
rect 2140 3367 2141 3371
rect 2135 3366 2141 3367
rect 2247 3371 2253 3372
rect 2247 3367 2248 3371
rect 2252 3370 2253 3371
rect 2271 3371 2277 3372
rect 2271 3370 2272 3371
rect 2252 3368 2272 3370
rect 2252 3367 2253 3368
rect 2247 3366 2253 3367
rect 2271 3367 2272 3368
rect 2276 3367 2277 3371
rect 2271 3366 2277 3367
rect 2383 3371 2389 3372
rect 2383 3367 2384 3371
rect 2388 3370 2389 3371
rect 2407 3371 2413 3372
rect 2407 3370 2408 3371
rect 2388 3368 2408 3370
rect 2388 3367 2389 3368
rect 2383 3366 2389 3367
rect 2407 3367 2408 3368
rect 2412 3367 2413 3371
rect 2407 3366 2413 3367
rect 2543 3371 2552 3372
rect 2543 3367 2544 3371
rect 2551 3367 2552 3371
rect 2543 3366 2552 3367
rect 2647 3371 2653 3372
rect 2647 3367 2648 3371
rect 2652 3370 2653 3371
rect 2671 3371 2677 3372
rect 2671 3370 2672 3371
rect 2652 3368 2672 3370
rect 2652 3367 2653 3368
rect 2647 3366 2653 3367
rect 2671 3367 2672 3368
rect 2676 3367 2677 3371
rect 2671 3366 2677 3367
rect 2775 3371 2781 3372
rect 2775 3367 2776 3371
rect 2780 3370 2781 3371
rect 2799 3371 2805 3372
rect 2799 3370 2800 3371
rect 2780 3368 2800 3370
rect 2780 3367 2781 3368
rect 2775 3366 2781 3367
rect 2799 3367 2800 3368
rect 2804 3367 2805 3371
rect 2799 3366 2805 3367
rect 2911 3371 2917 3372
rect 2911 3367 2912 3371
rect 2916 3370 2917 3371
rect 2935 3371 2941 3372
rect 2935 3370 2936 3371
rect 2916 3368 2936 3370
rect 2916 3367 2917 3368
rect 2911 3366 2917 3367
rect 2935 3367 2936 3368
rect 2940 3367 2941 3371
rect 2935 3366 2941 3367
rect 3047 3371 3053 3372
rect 3047 3367 3048 3371
rect 3052 3370 3053 3371
rect 3071 3371 3077 3372
rect 3071 3370 3072 3371
rect 3052 3368 3072 3370
rect 3052 3367 3053 3368
rect 3047 3366 3053 3367
rect 3071 3367 3072 3368
rect 3076 3367 3077 3371
rect 3071 3366 3077 3367
rect 738 3363 744 3364
rect 738 3362 739 3363
rect 284 3360 739 3362
rect 247 3355 253 3356
rect 247 3351 248 3355
rect 252 3354 253 3355
rect 284 3354 286 3360
rect 738 3359 739 3360
rect 743 3359 744 3363
rect 738 3358 744 3359
rect 1903 3359 1912 3360
rect 252 3352 286 3354
rect 327 3355 333 3356
rect 252 3351 253 3352
rect 247 3350 253 3351
rect 327 3351 328 3355
rect 332 3354 333 3355
rect 391 3355 397 3356
rect 391 3354 392 3355
rect 332 3352 392 3354
rect 332 3351 333 3352
rect 327 3350 333 3351
rect 391 3351 392 3352
rect 396 3351 397 3355
rect 391 3350 397 3351
rect 471 3355 477 3356
rect 471 3351 472 3355
rect 476 3354 477 3355
rect 551 3355 557 3356
rect 551 3354 552 3355
rect 476 3352 552 3354
rect 476 3351 477 3352
rect 471 3350 477 3351
rect 551 3351 552 3352
rect 556 3351 557 3355
rect 551 3350 557 3351
rect 631 3355 637 3356
rect 631 3351 632 3355
rect 636 3354 637 3355
rect 719 3355 725 3356
rect 719 3354 720 3355
rect 636 3352 720 3354
rect 636 3351 637 3352
rect 631 3350 637 3351
rect 719 3351 720 3352
rect 724 3351 725 3355
rect 719 3350 725 3351
rect 799 3355 805 3356
rect 799 3351 800 3355
rect 804 3354 805 3355
rect 879 3355 885 3356
rect 879 3354 880 3355
rect 804 3352 880 3354
rect 804 3351 805 3352
rect 799 3350 805 3351
rect 879 3351 880 3352
rect 884 3351 885 3355
rect 879 3350 885 3351
rect 1039 3355 1045 3356
rect 1039 3351 1040 3355
rect 1044 3354 1045 3355
rect 1086 3355 1092 3356
rect 1086 3354 1087 3355
rect 1044 3352 1087 3354
rect 1044 3351 1045 3352
rect 1039 3350 1045 3351
rect 1086 3351 1087 3352
rect 1091 3351 1092 3355
rect 1086 3350 1092 3351
rect 1095 3355 1101 3356
rect 1095 3351 1096 3355
rect 1100 3354 1101 3355
rect 1191 3355 1197 3356
rect 1191 3354 1192 3355
rect 1100 3352 1192 3354
rect 1100 3351 1101 3352
rect 1095 3350 1101 3351
rect 1191 3351 1192 3352
rect 1196 3351 1197 3355
rect 1191 3350 1197 3351
rect 1263 3355 1269 3356
rect 1263 3351 1264 3355
rect 1268 3354 1269 3355
rect 1343 3355 1349 3356
rect 1343 3354 1344 3355
rect 1268 3352 1344 3354
rect 1268 3351 1269 3352
rect 1263 3350 1269 3351
rect 1343 3351 1344 3352
rect 1348 3351 1349 3355
rect 1343 3350 1349 3351
rect 1415 3355 1421 3356
rect 1415 3351 1416 3355
rect 1420 3354 1421 3355
rect 1495 3355 1501 3356
rect 1495 3354 1496 3355
rect 1420 3352 1496 3354
rect 1420 3351 1421 3352
rect 1415 3350 1421 3351
rect 1495 3351 1496 3352
rect 1500 3351 1501 3355
rect 1495 3350 1501 3351
rect 1567 3355 1573 3356
rect 1567 3351 1568 3355
rect 1572 3354 1573 3355
rect 1647 3355 1653 3356
rect 1647 3354 1648 3355
rect 1572 3352 1648 3354
rect 1572 3351 1573 3352
rect 1567 3350 1573 3351
rect 1647 3351 1648 3352
rect 1652 3351 1653 3355
rect 1903 3355 1904 3359
rect 1911 3355 1912 3359
rect 1903 3354 1912 3355
rect 1959 3359 1965 3360
rect 1959 3355 1960 3359
rect 1964 3358 1965 3359
rect 2007 3359 2013 3360
rect 2007 3358 2008 3359
rect 1964 3356 2008 3358
rect 1964 3355 1965 3356
rect 1959 3354 1965 3355
rect 2007 3355 2008 3356
rect 2012 3355 2013 3359
rect 2007 3354 2013 3355
rect 2071 3359 2077 3360
rect 2071 3355 2072 3359
rect 2076 3358 2077 3359
rect 2143 3359 2149 3360
rect 2143 3358 2144 3359
rect 2076 3356 2144 3358
rect 2076 3355 2077 3356
rect 2071 3354 2077 3355
rect 2143 3355 2144 3356
rect 2148 3355 2149 3359
rect 2143 3354 2149 3355
rect 2215 3359 2221 3360
rect 2215 3355 2216 3359
rect 2220 3358 2221 3359
rect 2287 3359 2293 3360
rect 2287 3358 2288 3359
rect 2220 3356 2288 3358
rect 2220 3355 2221 3356
rect 2215 3354 2221 3355
rect 2287 3355 2288 3356
rect 2292 3355 2293 3359
rect 2287 3354 2293 3355
rect 2359 3359 2365 3360
rect 2359 3355 2360 3359
rect 2364 3358 2365 3359
rect 2431 3359 2437 3360
rect 2431 3358 2432 3359
rect 2364 3356 2432 3358
rect 2364 3355 2365 3356
rect 2359 3354 2365 3355
rect 2431 3355 2432 3356
rect 2436 3355 2437 3359
rect 2431 3354 2437 3355
rect 2567 3359 2573 3360
rect 2567 3355 2568 3359
rect 2572 3358 2573 3359
rect 2626 3359 2632 3360
rect 2626 3358 2627 3359
rect 2572 3356 2627 3358
rect 2572 3355 2573 3356
rect 2567 3354 2573 3355
rect 2626 3355 2627 3356
rect 2631 3355 2632 3359
rect 2626 3354 2632 3355
rect 2703 3359 2712 3360
rect 2703 3355 2704 3359
rect 2711 3355 2712 3359
rect 2703 3354 2712 3355
rect 2839 3359 2845 3360
rect 2839 3355 2840 3359
rect 2844 3358 2845 3359
rect 2898 3359 2904 3360
rect 2898 3358 2899 3359
rect 2844 3356 2899 3358
rect 2844 3355 2845 3356
rect 2839 3354 2845 3355
rect 2898 3355 2899 3356
rect 2903 3355 2904 3359
rect 2898 3354 2904 3355
rect 2975 3359 2981 3360
rect 2975 3355 2976 3359
rect 2980 3358 2981 3359
rect 3034 3359 3040 3360
rect 3034 3358 3035 3359
rect 2980 3356 3035 3358
rect 2980 3355 2981 3356
rect 2975 3354 2981 3355
rect 3034 3355 3035 3356
rect 3039 3355 3040 3359
rect 3034 3354 3040 3355
rect 3111 3359 3117 3360
rect 3111 3355 3112 3359
rect 3116 3358 3117 3359
rect 3122 3359 3128 3360
rect 3122 3358 3123 3359
rect 3116 3356 3123 3358
rect 3116 3355 3117 3356
rect 3111 3354 3117 3355
rect 3122 3355 3123 3356
rect 3127 3355 3128 3359
rect 3122 3354 3128 3355
rect 1647 3350 1653 3351
rect 1894 3349 1900 3350
rect 238 3345 244 3346
rect 238 3341 239 3345
rect 243 3341 244 3345
rect 238 3340 244 3341
rect 382 3345 388 3346
rect 382 3341 383 3345
rect 387 3341 388 3345
rect 382 3340 388 3341
rect 542 3345 548 3346
rect 542 3341 543 3345
rect 547 3341 548 3345
rect 542 3340 548 3341
rect 710 3345 716 3346
rect 710 3341 711 3345
rect 715 3341 716 3345
rect 710 3340 716 3341
rect 870 3345 876 3346
rect 870 3341 871 3345
rect 875 3341 876 3345
rect 870 3340 876 3341
rect 1030 3345 1036 3346
rect 1030 3341 1031 3345
rect 1035 3341 1036 3345
rect 1030 3340 1036 3341
rect 1182 3345 1188 3346
rect 1182 3341 1183 3345
rect 1187 3341 1188 3345
rect 1182 3340 1188 3341
rect 1334 3345 1340 3346
rect 1334 3341 1335 3345
rect 1339 3341 1340 3345
rect 1334 3340 1340 3341
rect 1486 3345 1492 3346
rect 1486 3341 1487 3345
rect 1491 3341 1492 3345
rect 1486 3340 1492 3341
rect 1638 3345 1644 3346
rect 1638 3341 1639 3345
rect 1643 3341 1644 3345
rect 1894 3345 1895 3349
rect 1899 3345 1900 3349
rect 1894 3344 1900 3345
rect 1998 3349 2004 3350
rect 1998 3345 1999 3349
rect 2003 3345 2004 3349
rect 1998 3344 2004 3345
rect 2134 3349 2140 3350
rect 2134 3345 2135 3349
rect 2139 3345 2140 3349
rect 2134 3344 2140 3345
rect 2278 3349 2284 3350
rect 2278 3345 2279 3349
rect 2283 3345 2284 3349
rect 2278 3344 2284 3345
rect 2422 3349 2428 3350
rect 2422 3345 2423 3349
rect 2427 3345 2428 3349
rect 2422 3344 2428 3345
rect 2558 3349 2564 3350
rect 2558 3345 2559 3349
rect 2563 3345 2564 3349
rect 2558 3344 2564 3345
rect 2694 3349 2700 3350
rect 2694 3345 2695 3349
rect 2699 3345 2700 3349
rect 2694 3344 2700 3345
rect 2830 3349 2836 3350
rect 2830 3345 2831 3349
rect 2835 3345 2836 3349
rect 2830 3344 2836 3345
rect 2966 3349 2972 3350
rect 2966 3345 2967 3349
rect 2971 3345 2972 3349
rect 2966 3344 2972 3345
rect 3102 3349 3108 3350
rect 3102 3345 3103 3349
rect 3107 3345 3108 3349
rect 3102 3344 3108 3345
rect 1638 3340 1644 3341
rect 1862 3336 1868 3337
rect 3574 3336 3580 3337
rect 110 3332 116 3333
rect 1822 3332 1828 3333
rect 110 3328 111 3332
rect 115 3328 116 3332
rect 327 3331 333 3332
rect 327 3330 328 3331
rect 293 3328 328 3330
rect 110 3327 116 3328
rect 327 3327 328 3328
rect 332 3327 333 3331
rect 471 3331 477 3332
rect 471 3330 472 3331
rect 437 3328 472 3330
rect 327 3326 333 3327
rect 471 3327 472 3328
rect 476 3327 477 3331
rect 631 3331 637 3332
rect 631 3330 632 3331
rect 597 3328 632 3330
rect 471 3326 477 3327
rect 631 3327 632 3328
rect 636 3327 637 3331
rect 799 3331 805 3332
rect 799 3330 800 3331
rect 765 3328 800 3330
rect 631 3326 637 3327
rect 799 3327 800 3328
rect 804 3327 805 3331
rect 1095 3331 1101 3332
rect 1095 3330 1096 3331
rect 1085 3328 1096 3330
rect 799 3326 805 3327
rect 1095 3327 1096 3328
rect 1100 3327 1101 3331
rect 1263 3331 1269 3332
rect 1263 3330 1264 3331
rect 1237 3328 1264 3330
rect 1095 3326 1101 3327
rect 1263 3327 1264 3328
rect 1268 3327 1269 3331
rect 1415 3331 1421 3332
rect 1415 3330 1416 3331
rect 1389 3328 1416 3330
rect 1263 3326 1269 3327
rect 1415 3327 1416 3328
rect 1420 3327 1421 3331
rect 1567 3331 1573 3332
rect 1567 3330 1568 3331
rect 1541 3328 1568 3330
rect 1415 3326 1421 3327
rect 1567 3327 1568 3328
rect 1572 3327 1573 3331
rect 1822 3328 1823 3332
rect 1827 3328 1828 3332
rect 1862 3332 1863 3336
rect 1867 3332 1868 3336
rect 1959 3335 1965 3336
rect 1959 3334 1960 3335
rect 1949 3332 1960 3334
rect 1862 3331 1868 3332
rect 1959 3331 1960 3332
rect 1964 3331 1965 3335
rect 2071 3335 2077 3336
rect 2071 3334 2072 3335
rect 2053 3332 2072 3334
rect 1959 3330 1965 3331
rect 2071 3331 2072 3332
rect 2076 3331 2077 3335
rect 2215 3335 2221 3336
rect 2215 3334 2216 3335
rect 2189 3332 2216 3334
rect 2071 3330 2077 3331
rect 2215 3331 2216 3332
rect 2220 3331 2221 3335
rect 2359 3335 2365 3336
rect 2359 3334 2360 3335
rect 2333 3332 2360 3334
rect 2215 3330 2221 3331
rect 2359 3331 2360 3332
rect 2364 3331 2365 3335
rect 3574 3332 3575 3336
rect 3579 3332 3580 3336
rect 2359 3330 2365 3331
rect 2546 3331 2552 3332
rect 1567 3326 1573 3327
rect 1582 3327 1588 3328
rect 1822 3327 1828 3328
rect 2546 3327 2547 3331
rect 2551 3330 2552 3331
rect 2626 3331 2632 3332
rect 2551 3328 2577 3330
rect 2551 3327 2552 3328
rect 1582 3323 1583 3327
rect 1587 3326 1588 3327
rect 2546 3326 2552 3327
rect 2626 3327 2627 3331
rect 2631 3330 2632 3331
rect 2898 3331 2904 3332
rect 2631 3328 2713 3330
rect 2631 3327 2632 3328
rect 2626 3326 2632 3327
rect 2898 3327 2899 3331
rect 2903 3330 2904 3331
rect 3034 3331 3040 3332
rect 3574 3331 3580 3332
rect 2903 3328 2985 3330
rect 2903 3327 2904 3328
rect 2898 3326 2904 3327
rect 3034 3327 3035 3331
rect 3039 3330 3040 3331
rect 3039 3328 3121 3330
rect 3039 3327 3040 3328
rect 3034 3326 3040 3327
rect 1587 3324 1657 3326
rect 1587 3323 1588 3324
rect 1582 3322 1588 3323
rect 1862 3319 1868 3320
rect 110 3315 116 3316
rect 110 3311 111 3315
rect 115 3311 116 3315
rect 110 3310 116 3311
rect 778 3315 784 3316
rect 778 3311 779 3315
rect 783 3314 784 3315
rect 1822 3315 1828 3316
rect 783 3312 881 3314
rect 783 3311 784 3312
rect 778 3310 784 3311
rect 1822 3311 1823 3315
rect 1827 3311 1828 3315
rect 1862 3315 1863 3319
rect 1867 3315 1868 3319
rect 1862 3314 1868 3315
rect 2358 3319 2364 3320
rect 2358 3315 2359 3319
rect 2363 3318 2364 3319
rect 2902 3319 2908 3320
rect 2902 3318 2903 3319
rect 2363 3316 2433 3318
rect 2881 3316 2903 3318
rect 2363 3315 2364 3316
rect 2358 3314 2364 3315
rect 2902 3315 2903 3316
rect 2907 3315 2908 3319
rect 2902 3314 2908 3315
rect 3574 3319 3580 3320
rect 3574 3315 3575 3319
rect 3579 3315 3580 3319
rect 3574 3314 3580 3315
rect 1822 3310 1828 3311
rect 1886 3309 1892 3310
rect 230 3305 236 3306
rect 230 3301 231 3305
rect 235 3301 236 3305
rect 230 3300 236 3301
rect 374 3305 380 3306
rect 374 3301 375 3305
rect 379 3301 380 3305
rect 374 3300 380 3301
rect 534 3305 540 3306
rect 534 3301 535 3305
rect 539 3301 540 3305
rect 534 3300 540 3301
rect 702 3305 708 3306
rect 702 3301 703 3305
rect 707 3301 708 3305
rect 702 3300 708 3301
rect 862 3305 868 3306
rect 862 3301 863 3305
rect 867 3301 868 3305
rect 862 3300 868 3301
rect 1022 3305 1028 3306
rect 1022 3301 1023 3305
rect 1027 3301 1028 3305
rect 1022 3300 1028 3301
rect 1174 3305 1180 3306
rect 1174 3301 1175 3305
rect 1179 3301 1180 3305
rect 1174 3300 1180 3301
rect 1326 3305 1332 3306
rect 1326 3301 1327 3305
rect 1331 3301 1332 3305
rect 1326 3300 1332 3301
rect 1478 3305 1484 3306
rect 1478 3301 1479 3305
rect 1483 3301 1484 3305
rect 1478 3300 1484 3301
rect 1630 3305 1636 3306
rect 1630 3301 1631 3305
rect 1635 3301 1636 3305
rect 1886 3305 1887 3309
rect 1891 3305 1892 3309
rect 1886 3304 1892 3305
rect 1990 3309 1996 3310
rect 1990 3305 1991 3309
rect 1995 3305 1996 3309
rect 1990 3304 1996 3305
rect 2126 3309 2132 3310
rect 2126 3305 2127 3309
rect 2131 3305 2132 3309
rect 2126 3304 2132 3305
rect 2270 3309 2276 3310
rect 2270 3305 2271 3309
rect 2275 3305 2276 3309
rect 2270 3304 2276 3305
rect 2414 3309 2420 3310
rect 2414 3305 2415 3309
rect 2419 3305 2420 3309
rect 2414 3304 2420 3305
rect 2550 3309 2556 3310
rect 2550 3305 2551 3309
rect 2555 3305 2556 3309
rect 2550 3304 2556 3305
rect 2686 3309 2692 3310
rect 2686 3305 2687 3309
rect 2691 3305 2692 3309
rect 2686 3304 2692 3305
rect 2822 3309 2828 3310
rect 2822 3305 2823 3309
rect 2827 3305 2828 3309
rect 2822 3304 2828 3305
rect 2958 3309 2964 3310
rect 2958 3305 2959 3309
rect 2963 3305 2964 3309
rect 2958 3304 2964 3305
rect 3094 3309 3100 3310
rect 3094 3305 3095 3309
rect 3099 3305 3100 3309
rect 3094 3304 3100 3305
rect 1630 3300 1636 3301
rect 1086 3287 1092 3288
rect 1086 3283 1087 3287
rect 1091 3286 1092 3287
rect 1926 3287 1932 3288
rect 1091 3284 1406 3286
rect 1091 3283 1092 3284
rect 1086 3282 1092 3283
rect 238 3279 244 3280
rect 238 3275 239 3279
rect 243 3275 244 3279
rect 238 3274 244 3275
rect 406 3279 412 3280
rect 406 3275 407 3279
rect 411 3275 412 3279
rect 406 3274 412 3275
rect 574 3279 580 3280
rect 574 3275 575 3279
rect 579 3275 580 3279
rect 574 3274 580 3275
rect 742 3279 748 3280
rect 742 3275 743 3279
rect 747 3275 748 3279
rect 742 3274 748 3275
rect 894 3279 900 3280
rect 894 3275 895 3279
rect 899 3275 900 3279
rect 894 3274 900 3275
rect 1046 3279 1052 3280
rect 1046 3275 1047 3279
rect 1051 3275 1052 3279
rect 1046 3274 1052 3275
rect 1190 3279 1196 3280
rect 1190 3275 1191 3279
rect 1195 3275 1196 3279
rect 1190 3274 1196 3275
rect 1334 3279 1340 3280
rect 1334 3275 1335 3279
rect 1339 3275 1340 3279
rect 1334 3274 1340 3275
rect 498 3271 504 3272
rect 110 3269 116 3270
rect 110 3265 111 3269
rect 115 3265 116 3269
rect 498 3267 499 3271
rect 503 3270 504 3271
rect 1404 3270 1406 3284
rect 1926 3283 1927 3287
rect 1931 3283 1932 3287
rect 1926 3282 1932 3283
rect 2046 3287 2052 3288
rect 2046 3283 2047 3287
rect 2051 3283 2052 3287
rect 2046 3282 2052 3283
rect 2174 3287 2180 3288
rect 2174 3283 2175 3287
rect 2179 3283 2180 3287
rect 2174 3282 2180 3283
rect 2310 3287 2316 3288
rect 2310 3283 2311 3287
rect 2315 3283 2316 3287
rect 2310 3282 2316 3283
rect 2454 3287 2460 3288
rect 2454 3283 2455 3287
rect 2459 3283 2460 3287
rect 2454 3282 2460 3283
rect 2598 3287 2604 3288
rect 2598 3283 2599 3287
rect 2603 3283 2604 3287
rect 2598 3282 2604 3283
rect 2742 3287 2748 3288
rect 2742 3283 2743 3287
rect 2747 3283 2748 3287
rect 2742 3282 2748 3283
rect 2886 3287 2892 3288
rect 2886 3283 2887 3287
rect 2891 3283 2892 3287
rect 2886 3282 2892 3283
rect 3030 3287 3036 3288
rect 3030 3283 3031 3287
rect 3035 3283 3036 3287
rect 3030 3282 3036 3283
rect 3182 3287 3188 3288
rect 3182 3283 3183 3287
rect 3187 3283 3188 3287
rect 3182 3282 3188 3283
rect 1486 3279 1492 3280
rect 1486 3275 1487 3279
rect 1491 3275 1492 3279
rect 2382 3279 2388 3280
rect 1486 3274 1492 3275
rect 1862 3277 1868 3278
rect 1862 3273 1863 3277
rect 1867 3273 1868 3277
rect 2382 3275 2383 3279
rect 2387 3278 2388 3279
rect 2706 3279 2712 3280
rect 2387 3276 2473 3278
rect 2387 3275 2388 3276
rect 2382 3274 2388 3275
rect 2706 3275 2707 3279
rect 2711 3278 2712 3279
rect 2711 3276 2761 3278
rect 3574 3277 3580 3278
rect 2711 3275 2712 3276
rect 2706 3274 2712 3275
rect 1862 3272 1868 3273
rect 3574 3273 3575 3277
rect 3579 3273 3580 3277
rect 3574 3272 3580 3273
rect 503 3268 593 3270
rect 1404 3268 1505 3270
rect 1822 3269 1828 3270
rect 503 3267 504 3268
rect 498 3266 504 3267
rect 110 3264 116 3265
rect 1822 3265 1823 3269
rect 1827 3265 1828 3269
rect 1822 3264 1828 3265
rect 2039 3263 2045 3264
rect 2039 3262 2040 3263
rect 1862 3260 1868 3261
rect 1989 3260 2040 3262
rect 1862 3256 1863 3260
rect 1867 3256 1868 3260
rect 2039 3259 2040 3260
rect 2044 3259 2045 3263
rect 2167 3263 2173 3264
rect 2167 3262 2168 3263
rect 2109 3260 2168 3262
rect 2039 3258 2045 3259
rect 2167 3259 2168 3260
rect 2172 3259 2173 3263
rect 2303 3263 2309 3264
rect 2303 3262 2304 3263
rect 2237 3260 2304 3262
rect 2167 3258 2173 3259
rect 2303 3259 2304 3260
rect 2308 3259 2309 3263
rect 2447 3263 2453 3264
rect 2447 3262 2448 3263
rect 2373 3260 2448 3262
rect 2303 3258 2309 3259
rect 2447 3259 2448 3260
rect 2452 3259 2453 3263
rect 2735 3263 2741 3264
rect 2735 3262 2736 3263
rect 2661 3260 2736 3262
rect 2447 3258 2453 3259
rect 2735 3259 2736 3260
rect 2740 3259 2741 3263
rect 3023 3263 3029 3264
rect 3023 3262 3024 3263
rect 2949 3260 3024 3262
rect 2735 3258 2741 3259
rect 3023 3259 3024 3260
rect 3028 3259 3029 3263
rect 3175 3263 3181 3264
rect 3175 3262 3176 3263
rect 3093 3260 3176 3262
rect 3023 3258 3029 3259
rect 3175 3259 3176 3260
rect 3180 3259 3181 3263
rect 3286 3263 3292 3264
rect 3286 3262 3287 3263
rect 3245 3260 3287 3262
rect 3175 3258 3181 3259
rect 3286 3259 3287 3260
rect 3291 3259 3292 3263
rect 3286 3258 3292 3259
rect 3574 3260 3580 3261
rect 399 3255 405 3256
rect 399 3254 400 3255
rect 110 3252 116 3253
rect 301 3252 400 3254
rect 110 3248 111 3252
rect 115 3248 116 3252
rect 399 3251 400 3252
rect 404 3251 405 3255
rect 566 3255 572 3256
rect 566 3254 567 3255
rect 469 3252 567 3254
rect 399 3250 405 3251
rect 566 3251 567 3252
rect 571 3251 572 3255
rect 566 3250 572 3251
rect 642 3255 648 3256
rect 642 3251 643 3255
rect 647 3254 648 3255
rect 1039 3255 1045 3256
rect 1039 3254 1040 3255
rect 647 3252 769 3254
rect 957 3252 1040 3254
rect 647 3251 648 3252
rect 642 3250 648 3251
rect 1039 3251 1040 3252
rect 1044 3251 1045 3255
rect 1183 3255 1189 3256
rect 1183 3254 1184 3255
rect 1109 3252 1184 3254
rect 1039 3250 1045 3251
rect 1183 3251 1184 3252
rect 1188 3251 1189 3255
rect 1327 3255 1333 3256
rect 1327 3254 1328 3255
rect 1253 3252 1328 3254
rect 1183 3250 1189 3251
rect 1327 3251 1328 3252
rect 1332 3251 1333 3255
rect 1479 3255 1485 3256
rect 1862 3255 1868 3256
rect 3574 3256 3575 3260
rect 3579 3256 3580 3260
rect 3574 3255 3580 3256
rect 1479 3254 1480 3255
rect 1397 3252 1480 3254
rect 1327 3250 1333 3251
rect 1479 3251 1480 3252
rect 1484 3251 1485 3255
rect 1479 3250 1485 3251
rect 1822 3252 1828 3253
rect 110 3247 116 3248
rect 1822 3248 1823 3252
rect 1827 3248 1828 3252
rect 1822 3247 1828 3248
rect 1934 3247 1940 3248
rect 1934 3243 1935 3247
rect 1939 3243 1940 3247
rect 1934 3242 1940 3243
rect 2054 3247 2060 3248
rect 2054 3243 2055 3247
rect 2059 3243 2060 3247
rect 2054 3242 2060 3243
rect 2182 3247 2188 3248
rect 2182 3243 2183 3247
rect 2187 3243 2188 3247
rect 2182 3242 2188 3243
rect 2318 3247 2324 3248
rect 2318 3243 2319 3247
rect 2323 3243 2324 3247
rect 2318 3242 2324 3243
rect 2462 3247 2468 3248
rect 2462 3243 2463 3247
rect 2467 3243 2468 3247
rect 2462 3242 2468 3243
rect 2606 3247 2612 3248
rect 2606 3243 2607 3247
rect 2611 3243 2612 3247
rect 2606 3242 2612 3243
rect 2750 3247 2756 3248
rect 2750 3243 2751 3247
rect 2755 3243 2756 3247
rect 2750 3242 2756 3243
rect 2894 3247 2900 3248
rect 2894 3243 2895 3247
rect 2899 3243 2900 3247
rect 2894 3242 2900 3243
rect 3038 3247 3044 3248
rect 3038 3243 3039 3247
rect 3043 3243 3044 3247
rect 3038 3242 3044 3243
rect 3190 3247 3196 3248
rect 3190 3243 3191 3247
rect 3195 3243 3196 3247
rect 3190 3242 3196 3243
rect 246 3239 252 3240
rect 246 3235 247 3239
rect 251 3235 252 3239
rect 246 3234 252 3235
rect 414 3239 420 3240
rect 414 3235 415 3239
rect 419 3235 420 3239
rect 414 3234 420 3235
rect 582 3239 588 3240
rect 582 3235 583 3239
rect 587 3235 588 3239
rect 582 3234 588 3235
rect 750 3239 756 3240
rect 750 3235 751 3239
rect 755 3235 756 3239
rect 750 3234 756 3235
rect 902 3239 908 3240
rect 902 3235 903 3239
rect 907 3235 908 3239
rect 902 3234 908 3235
rect 1054 3239 1060 3240
rect 1054 3235 1055 3239
rect 1059 3235 1060 3239
rect 1054 3234 1060 3235
rect 1198 3239 1204 3240
rect 1198 3235 1199 3239
rect 1203 3235 1204 3239
rect 1198 3234 1204 3235
rect 1342 3239 1348 3240
rect 1342 3235 1343 3239
rect 1347 3235 1348 3239
rect 1342 3234 1348 3235
rect 1494 3239 1500 3240
rect 1494 3235 1495 3239
rect 1499 3235 1500 3239
rect 1494 3234 1500 3235
rect 1943 3235 1952 3236
rect 1943 3231 1944 3235
rect 1951 3231 1952 3235
rect 1943 3230 1952 3231
rect 2039 3235 2045 3236
rect 2039 3231 2040 3235
rect 2044 3234 2045 3235
rect 2063 3235 2069 3236
rect 2063 3234 2064 3235
rect 2044 3232 2064 3234
rect 2044 3231 2045 3232
rect 2039 3230 2045 3231
rect 2063 3231 2064 3232
rect 2068 3231 2069 3235
rect 2063 3230 2069 3231
rect 2167 3235 2173 3236
rect 2167 3231 2168 3235
rect 2172 3234 2173 3235
rect 2191 3235 2197 3236
rect 2191 3234 2192 3235
rect 2172 3232 2192 3234
rect 2172 3231 2173 3232
rect 2167 3230 2173 3231
rect 2191 3231 2192 3232
rect 2196 3231 2197 3235
rect 2191 3230 2197 3231
rect 2303 3235 2309 3236
rect 2303 3231 2304 3235
rect 2308 3234 2309 3235
rect 2327 3235 2333 3236
rect 2327 3234 2328 3235
rect 2308 3232 2328 3234
rect 2308 3231 2309 3232
rect 2303 3230 2309 3231
rect 2327 3231 2328 3232
rect 2332 3231 2333 3235
rect 2327 3230 2333 3231
rect 2447 3235 2453 3236
rect 2447 3231 2448 3235
rect 2452 3234 2453 3235
rect 2471 3235 2477 3236
rect 2471 3234 2472 3235
rect 2452 3232 2472 3234
rect 2452 3231 2453 3232
rect 2447 3230 2453 3231
rect 2471 3231 2472 3232
rect 2476 3231 2477 3235
rect 2471 3230 2477 3231
rect 2615 3235 2624 3236
rect 2615 3231 2616 3235
rect 2623 3231 2624 3235
rect 2615 3230 2624 3231
rect 2735 3235 2741 3236
rect 2735 3231 2736 3235
rect 2740 3234 2741 3235
rect 2759 3235 2765 3236
rect 2759 3234 2760 3235
rect 2740 3232 2760 3234
rect 2740 3231 2741 3232
rect 2735 3230 2741 3231
rect 2759 3231 2760 3232
rect 2764 3231 2765 3235
rect 2759 3230 2765 3231
rect 2902 3235 2909 3236
rect 2902 3231 2903 3235
rect 2908 3231 2909 3235
rect 2902 3230 2909 3231
rect 3023 3235 3029 3236
rect 3023 3231 3024 3235
rect 3028 3234 3029 3235
rect 3047 3235 3053 3236
rect 3047 3234 3048 3235
rect 3028 3232 3048 3234
rect 3028 3231 3029 3232
rect 3023 3230 3029 3231
rect 3047 3231 3048 3232
rect 3052 3231 3053 3235
rect 3047 3230 3053 3231
rect 3175 3235 3181 3236
rect 3175 3231 3176 3235
rect 3180 3234 3181 3235
rect 3199 3235 3205 3236
rect 3199 3234 3200 3235
rect 3180 3232 3200 3234
rect 3180 3231 3181 3232
rect 3175 3230 3181 3231
rect 3199 3231 3200 3232
rect 3204 3231 3205 3235
rect 3199 3230 3205 3231
rect 255 3227 264 3228
rect 255 3223 256 3227
rect 263 3223 264 3227
rect 255 3222 264 3223
rect 399 3227 405 3228
rect 399 3223 400 3227
rect 404 3226 405 3227
rect 423 3227 429 3228
rect 423 3226 424 3227
rect 404 3224 424 3226
rect 404 3223 405 3224
rect 399 3222 405 3223
rect 423 3223 424 3224
rect 428 3223 429 3227
rect 423 3222 429 3223
rect 591 3227 597 3228
rect 591 3223 592 3227
rect 596 3226 597 3227
rect 642 3227 648 3228
rect 642 3226 643 3227
rect 596 3224 643 3226
rect 596 3223 597 3224
rect 591 3222 597 3223
rect 642 3223 643 3224
rect 647 3223 648 3227
rect 642 3222 648 3223
rect 759 3227 765 3228
rect 759 3223 760 3227
rect 764 3226 765 3227
rect 778 3227 784 3228
rect 778 3226 779 3227
rect 764 3224 779 3226
rect 764 3223 765 3224
rect 759 3222 765 3223
rect 778 3223 779 3224
rect 783 3223 784 3227
rect 778 3222 784 3223
rect 911 3227 917 3228
rect 911 3223 912 3227
rect 916 3226 917 3227
rect 1030 3227 1036 3228
rect 1030 3226 1031 3227
rect 916 3224 1031 3226
rect 916 3223 917 3224
rect 911 3222 917 3223
rect 1030 3223 1031 3224
rect 1035 3223 1036 3227
rect 1030 3222 1036 3223
rect 1039 3227 1045 3228
rect 1039 3223 1040 3227
rect 1044 3226 1045 3227
rect 1063 3227 1069 3228
rect 1063 3226 1064 3227
rect 1044 3224 1064 3226
rect 1044 3223 1045 3224
rect 1039 3222 1045 3223
rect 1063 3223 1064 3224
rect 1068 3223 1069 3227
rect 1063 3222 1069 3223
rect 1183 3227 1189 3228
rect 1183 3223 1184 3227
rect 1188 3226 1189 3227
rect 1207 3227 1213 3228
rect 1207 3226 1208 3227
rect 1188 3224 1208 3226
rect 1188 3223 1189 3224
rect 1183 3222 1189 3223
rect 1207 3223 1208 3224
rect 1212 3223 1213 3227
rect 1207 3222 1213 3223
rect 1327 3227 1333 3228
rect 1327 3223 1328 3227
rect 1332 3226 1333 3227
rect 1351 3227 1357 3228
rect 1351 3226 1352 3227
rect 1332 3224 1352 3226
rect 1332 3223 1333 3224
rect 1327 3222 1333 3223
rect 1351 3223 1352 3224
rect 1356 3223 1357 3227
rect 1351 3222 1357 3223
rect 1479 3227 1485 3228
rect 1479 3223 1480 3227
rect 1484 3226 1485 3227
rect 1503 3227 1509 3228
rect 1503 3226 1504 3227
rect 1484 3224 1504 3226
rect 1484 3223 1485 3224
rect 1479 3222 1485 3223
rect 1503 3223 1504 3224
rect 1508 3223 1509 3227
rect 1503 3222 1509 3223
rect 2382 3223 2388 3224
rect 2382 3222 2383 3223
rect 2064 3220 2383 3222
rect 2015 3215 2021 3216
rect 2015 3211 2016 3215
rect 2020 3214 2021 3215
rect 2064 3214 2066 3220
rect 2382 3219 2383 3220
rect 2387 3219 2388 3223
rect 2382 3218 2388 3219
rect 2020 3212 2066 3214
rect 2071 3215 2077 3216
rect 2020 3211 2021 3212
rect 2015 3210 2021 3211
rect 2071 3211 2072 3215
rect 2076 3214 2077 3215
rect 2127 3215 2133 3216
rect 2127 3214 2128 3215
rect 2076 3212 2128 3214
rect 2076 3211 2077 3212
rect 2071 3210 2077 3211
rect 2127 3211 2128 3212
rect 2132 3211 2133 3215
rect 2127 3210 2133 3211
rect 2183 3215 2189 3216
rect 2183 3211 2184 3215
rect 2188 3214 2189 3215
rect 2247 3215 2253 3216
rect 2247 3214 2248 3215
rect 2188 3212 2248 3214
rect 2188 3211 2189 3212
rect 2183 3210 2189 3211
rect 2247 3211 2248 3212
rect 2252 3211 2253 3215
rect 2247 3210 2253 3211
rect 2311 3215 2317 3216
rect 2311 3211 2312 3215
rect 2316 3214 2317 3215
rect 2383 3215 2389 3216
rect 2383 3214 2384 3215
rect 2316 3212 2384 3214
rect 2316 3211 2317 3212
rect 2311 3210 2317 3211
rect 2383 3211 2384 3212
rect 2388 3211 2389 3215
rect 2383 3210 2389 3211
rect 2455 3215 2461 3216
rect 2455 3211 2456 3215
rect 2460 3214 2461 3215
rect 2527 3215 2533 3216
rect 2527 3214 2528 3215
rect 2460 3212 2528 3214
rect 2460 3211 2461 3212
rect 2455 3210 2461 3211
rect 2527 3211 2528 3212
rect 2532 3211 2533 3215
rect 2527 3210 2533 3211
rect 2671 3215 2677 3216
rect 2671 3211 2672 3215
rect 2676 3214 2677 3215
rect 2743 3215 2749 3216
rect 2743 3214 2744 3215
rect 2676 3212 2744 3214
rect 2676 3211 2677 3212
rect 2671 3210 2677 3211
rect 2743 3211 2744 3212
rect 2748 3211 2749 3215
rect 2743 3210 2749 3211
rect 2751 3215 2757 3216
rect 2751 3211 2752 3215
rect 2756 3214 2757 3215
rect 2823 3215 2829 3216
rect 2823 3214 2824 3215
rect 2756 3212 2824 3214
rect 2756 3211 2757 3212
rect 2751 3210 2757 3211
rect 2823 3211 2824 3212
rect 2828 3211 2829 3215
rect 2823 3210 2829 3211
rect 2975 3215 2981 3216
rect 2975 3211 2976 3215
rect 2980 3214 2981 3215
rect 3046 3215 3052 3216
rect 3046 3214 3047 3215
rect 2980 3212 3047 3214
rect 2980 3211 2981 3212
rect 2975 3210 2981 3211
rect 3046 3211 3047 3212
rect 3051 3211 3052 3215
rect 3046 3210 3052 3211
rect 3127 3215 3133 3216
rect 3127 3211 3128 3215
rect 3132 3214 3133 3215
rect 3191 3215 3197 3216
rect 3191 3214 3192 3215
rect 3132 3212 3192 3214
rect 3132 3211 3133 3212
rect 3127 3210 3133 3211
rect 3191 3211 3192 3212
rect 3196 3211 3197 3215
rect 3191 3210 3197 3211
rect 3286 3215 3293 3216
rect 3286 3211 3287 3215
rect 3292 3211 3293 3215
rect 3286 3210 3293 3211
rect 2006 3205 2012 3206
rect 183 3203 189 3204
rect 183 3199 184 3203
rect 188 3202 189 3203
rect 258 3203 264 3204
rect 258 3202 259 3203
rect 188 3200 259 3202
rect 188 3199 189 3200
rect 183 3198 189 3199
rect 258 3199 259 3200
rect 263 3199 264 3203
rect 258 3198 264 3199
rect 383 3203 389 3204
rect 383 3199 384 3203
rect 388 3202 389 3203
rect 478 3203 484 3204
rect 478 3202 479 3203
rect 388 3200 479 3202
rect 388 3199 389 3200
rect 383 3198 389 3199
rect 478 3199 479 3200
rect 483 3199 484 3203
rect 478 3198 484 3199
rect 566 3203 573 3204
rect 566 3199 567 3203
rect 572 3199 573 3203
rect 566 3198 573 3199
rect 735 3203 741 3204
rect 735 3199 736 3203
rect 740 3202 741 3203
rect 806 3203 812 3204
rect 806 3202 807 3203
rect 740 3200 807 3202
rect 740 3199 741 3200
rect 735 3198 741 3199
rect 806 3199 807 3200
rect 811 3199 812 3203
rect 806 3198 812 3199
rect 815 3203 821 3204
rect 815 3199 816 3203
rect 820 3202 821 3203
rect 895 3203 901 3204
rect 895 3202 896 3203
rect 820 3200 896 3202
rect 820 3199 821 3200
rect 815 3198 821 3199
rect 895 3199 896 3200
rect 900 3199 901 3203
rect 895 3198 901 3199
rect 967 3203 973 3204
rect 967 3199 968 3203
rect 972 3202 973 3203
rect 1047 3203 1053 3204
rect 1047 3202 1048 3203
rect 972 3200 1048 3202
rect 972 3199 973 3200
rect 967 3198 973 3199
rect 1047 3199 1048 3200
rect 1052 3199 1053 3203
rect 1047 3198 1053 3199
rect 1103 3203 1109 3204
rect 1103 3199 1104 3203
rect 1108 3202 1109 3203
rect 1199 3203 1205 3204
rect 1199 3202 1200 3203
rect 1108 3200 1200 3202
rect 1108 3199 1109 3200
rect 1103 3198 1109 3199
rect 1199 3199 1200 3200
rect 1204 3199 1205 3203
rect 1199 3198 1205 3199
rect 1263 3203 1269 3204
rect 1263 3199 1264 3203
rect 1268 3202 1269 3203
rect 1359 3203 1365 3204
rect 1359 3202 1360 3203
rect 1268 3200 1360 3202
rect 1268 3199 1269 3200
rect 1263 3198 1269 3199
rect 1359 3199 1360 3200
rect 1364 3199 1365 3203
rect 2006 3201 2007 3205
rect 2011 3201 2012 3205
rect 2006 3200 2012 3201
rect 2118 3205 2124 3206
rect 2118 3201 2119 3205
rect 2123 3201 2124 3205
rect 2118 3200 2124 3201
rect 2238 3205 2244 3206
rect 2238 3201 2239 3205
rect 2243 3201 2244 3205
rect 2238 3200 2244 3201
rect 2374 3205 2380 3206
rect 2374 3201 2375 3205
rect 2379 3201 2380 3205
rect 2374 3200 2380 3201
rect 2518 3205 2524 3206
rect 2518 3201 2519 3205
rect 2523 3201 2524 3205
rect 2518 3200 2524 3201
rect 2662 3205 2668 3206
rect 2662 3201 2663 3205
rect 2667 3201 2668 3205
rect 2662 3200 2668 3201
rect 2814 3205 2820 3206
rect 2814 3201 2815 3205
rect 2819 3201 2820 3205
rect 2814 3200 2820 3201
rect 2966 3205 2972 3206
rect 2966 3201 2967 3205
rect 2971 3201 2972 3205
rect 2966 3200 2972 3201
rect 3118 3205 3124 3206
rect 3118 3201 3119 3205
rect 3123 3201 3124 3205
rect 3118 3200 3124 3201
rect 3278 3205 3284 3206
rect 3278 3201 3279 3205
rect 3283 3201 3284 3205
rect 3278 3200 3284 3201
rect 1359 3198 1365 3199
rect 174 3193 180 3194
rect 174 3189 175 3193
rect 179 3189 180 3193
rect 174 3188 180 3189
rect 374 3193 380 3194
rect 374 3189 375 3193
rect 379 3189 380 3193
rect 374 3188 380 3189
rect 558 3193 564 3194
rect 558 3189 559 3193
rect 563 3189 564 3193
rect 558 3188 564 3189
rect 726 3193 732 3194
rect 726 3189 727 3193
rect 731 3189 732 3193
rect 726 3188 732 3189
rect 886 3193 892 3194
rect 886 3189 887 3193
rect 891 3189 892 3193
rect 886 3188 892 3189
rect 1038 3193 1044 3194
rect 1038 3189 1039 3193
rect 1043 3189 1044 3193
rect 1038 3188 1044 3189
rect 1190 3193 1196 3194
rect 1190 3189 1191 3193
rect 1195 3189 1196 3193
rect 1190 3188 1196 3189
rect 1350 3193 1356 3194
rect 1350 3189 1351 3193
rect 1355 3189 1356 3193
rect 1350 3188 1356 3189
rect 1862 3192 1868 3193
rect 3574 3192 3580 3193
rect 1862 3188 1863 3192
rect 1867 3188 1868 3192
rect 2071 3191 2077 3192
rect 2071 3190 2072 3191
rect 2061 3188 2072 3190
rect 1862 3187 1868 3188
rect 2071 3187 2072 3188
rect 2076 3187 2077 3191
rect 2183 3191 2189 3192
rect 2183 3190 2184 3191
rect 2173 3188 2184 3190
rect 2071 3186 2077 3187
rect 2183 3187 2184 3188
rect 2188 3187 2189 3191
rect 2311 3191 2317 3192
rect 2311 3190 2312 3191
rect 2293 3188 2312 3190
rect 2183 3186 2189 3187
rect 2311 3187 2312 3188
rect 2316 3187 2317 3191
rect 2455 3191 2461 3192
rect 2455 3190 2456 3191
rect 2429 3188 2456 3190
rect 2311 3186 2317 3187
rect 2455 3187 2456 3188
rect 2460 3187 2461 3191
rect 3574 3188 3575 3192
rect 3579 3188 3580 3192
rect 2455 3186 2461 3187
rect 2618 3187 2624 3188
rect 2618 3183 2619 3187
rect 2623 3186 2624 3187
rect 2743 3187 2749 3188
rect 2623 3184 2681 3186
rect 2623 3183 2624 3184
rect 2618 3182 2624 3183
rect 2743 3183 2744 3187
rect 2748 3186 2749 3187
rect 3046 3187 3052 3188
rect 2748 3184 2833 3186
rect 2748 3183 2749 3184
rect 2743 3182 2749 3183
rect 3046 3183 3047 3187
rect 3051 3186 3052 3187
rect 3191 3187 3197 3188
rect 3574 3187 3580 3188
rect 3051 3184 3137 3186
rect 3051 3183 3052 3184
rect 3046 3182 3052 3183
rect 3191 3183 3192 3187
rect 3196 3186 3197 3187
rect 3196 3184 3297 3186
rect 3196 3183 3197 3184
rect 3191 3182 3197 3183
rect 110 3180 116 3181
rect 1822 3180 1828 3181
rect 110 3176 111 3180
rect 115 3176 116 3180
rect 815 3179 821 3180
rect 815 3178 816 3179
rect 781 3176 816 3178
rect 110 3175 116 3176
rect 258 3175 264 3176
rect 258 3171 259 3175
rect 263 3174 264 3175
rect 478 3175 484 3176
rect 263 3172 393 3174
rect 263 3171 264 3172
rect 258 3170 264 3171
rect 478 3171 479 3175
rect 483 3174 484 3175
rect 815 3175 816 3176
rect 820 3175 821 3179
rect 967 3179 973 3180
rect 967 3178 968 3179
rect 941 3176 968 3178
rect 815 3174 821 3175
rect 967 3175 968 3176
rect 972 3175 973 3179
rect 1103 3179 1109 3180
rect 1103 3178 1104 3179
rect 1093 3176 1104 3178
rect 967 3174 973 3175
rect 1103 3175 1104 3176
rect 1108 3175 1109 3179
rect 1263 3179 1269 3180
rect 1263 3178 1264 3179
rect 1245 3176 1264 3178
rect 1103 3174 1109 3175
rect 1263 3175 1264 3176
rect 1268 3175 1269 3179
rect 1822 3176 1823 3180
rect 1827 3176 1828 3180
rect 1263 3174 1269 3175
rect 1278 3175 1284 3176
rect 1822 3175 1828 3176
rect 1862 3175 1868 3176
rect 483 3172 577 3174
rect 483 3171 484 3172
rect 478 3170 484 3171
rect 1278 3171 1279 3175
rect 1283 3174 1284 3175
rect 1283 3172 1369 3174
rect 1283 3171 1284 3172
rect 1278 3170 1284 3171
rect 1862 3171 1863 3175
rect 1867 3171 1868 3175
rect 1862 3170 1868 3171
rect 2903 3175 2909 3176
rect 2903 3171 2904 3175
rect 2908 3174 2909 3175
rect 3574 3175 3580 3176
rect 2908 3172 2977 3174
rect 2908 3171 2909 3172
rect 2903 3170 2909 3171
rect 3574 3171 3575 3175
rect 3579 3171 3580 3175
rect 3574 3170 3580 3171
rect 1998 3165 2004 3166
rect 110 3163 116 3164
rect 110 3159 111 3163
rect 115 3159 116 3163
rect 110 3158 116 3159
rect 154 3163 160 3164
rect 154 3159 155 3163
rect 159 3162 160 3163
rect 1822 3163 1828 3164
rect 159 3160 185 3162
rect 159 3159 160 3160
rect 154 3158 160 3159
rect 1822 3159 1823 3163
rect 1827 3159 1828 3163
rect 1998 3161 1999 3165
rect 2003 3161 2004 3165
rect 1998 3160 2004 3161
rect 2110 3165 2116 3166
rect 2110 3161 2111 3165
rect 2115 3161 2116 3165
rect 2110 3160 2116 3161
rect 2230 3165 2236 3166
rect 2230 3161 2231 3165
rect 2235 3161 2236 3165
rect 2230 3160 2236 3161
rect 2366 3165 2372 3166
rect 2366 3161 2367 3165
rect 2371 3161 2372 3165
rect 2366 3160 2372 3161
rect 2510 3165 2516 3166
rect 2510 3161 2511 3165
rect 2515 3161 2516 3165
rect 2510 3160 2516 3161
rect 2654 3165 2660 3166
rect 2654 3161 2655 3165
rect 2659 3161 2660 3165
rect 2654 3160 2660 3161
rect 2806 3165 2812 3166
rect 2806 3161 2807 3165
rect 2811 3161 2812 3165
rect 2806 3160 2812 3161
rect 2958 3165 2964 3166
rect 2958 3161 2959 3165
rect 2963 3161 2964 3165
rect 2958 3160 2964 3161
rect 3110 3165 3116 3166
rect 3110 3161 3111 3165
rect 3115 3161 3116 3165
rect 3110 3160 3116 3161
rect 3270 3165 3276 3166
rect 3270 3161 3271 3165
rect 3275 3161 3276 3165
rect 3270 3160 3276 3161
rect 1822 3158 1828 3159
rect 2530 3159 2536 3160
rect 2530 3155 2531 3159
rect 2535 3158 2536 3159
rect 2559 3159 2565 3160
rect 2559 3158 2560 3159
rect 2535 3156 2560 3158
rect 2535 3155 2536 3156
rect 2530 3154 2536 3155
rect 2559 3155 2560 3156
rect 2564 3155 2565 3159
rect 2559 3154 2565 3155
rect 166 3153 172 3154
rect 166 3149 167 3153
rect 171 3149 172 3153
rect 166 3148 172 3149
rect 366 3153 372 3154
rect 366 3149 367 3153
rect 371 3149 372 3153
rect 366 3148 372 3149
rect 550 3153 556 3154
rect 550 3149 551 3153
rect 555 3149 556 3153
rect 550 3148 556 3149
rect 718 3153 724 3154
rect 718 3149 719 3153
rect 723 3149 724 3153
rect 718 3148 724 3149
rect 878 3153 884 3154
rect 878 3149 879 3153
rect 883 3149 884 3153
rect 878 3148 884 3149
rect 1030 3153 1036 3154
rect 1030 3149 1031 3153
rect 1035 3149 1036 3153
rect 1030 3148 1036 3149
rect 1182 3153 1188 3154
rect 1182 3149 1183 3153
rect 1187 3149 1188 3153
rect 1182 3148 1188 3149
rect 1342 3153 1348 3154
rect 1342 3149 1343 3153
rect 1347 3149 1348 3153
rect 1342 3148 1348 3149
rect 2054 3139 2060 3140
rect 2054 3135 2055 3139
rect 2059 3135 2060 3139
rect 2054 3134 2060 3135
rect 2206 3139 2212 3140
rect 2206 3135 2207 3139
rect 2211 3135 2212 3139
rect 2206 3134 2212 3135
rect 2358 3139 2364 3140
rect 2358 3135 2359 3139
rect 2363 3135 2364 3139
rect 2358 3134 2364 3135
rect 2510 3139 2516 3140
rect 2510 3135 2511 3139
rect 2515 3135 2516 3139
rect 2510 3134 2516 3135
rect 2654 3139 2660 3140
rect 2654 3135 2655 3139
rect 2659 3135 2660 3139
rect 2654 3134 2660 3135
rect 2790 3139 2796 3140
rect 2790 3135 2791 3139
rect 2795 3135 2796 3139
rect 2790 3134 2796 3135
rect 2918 3139 2924 3140
rect 2918 3135 2919 3139
rect 2923 3135 2924 3139
rect 2918 3134 2924 3135
rect 3038 3139 3044 3140
rect 3038 3135 3039 3139
rect 3043 3135 3044 3139
rect 3038 3134 3044 3135
rect 3158 3139 3164 3140
rect 3158 3135 3159 3139
rect 3163 3135 3164 3139
rect 3158 3134 3164 3135
rect 3270 3139 3276 3140
rect 3270 3135 3271 3139
rect 3275 3135 3276 3139
rect 3270 3134 3276 3135
rect 3382 3139 3388 3140
rect 3382 3135 3383 3139
rect 3387 3135 3388 3139
rect 3382 3134 3388 3135
rect 3478 3139 3484 3140
rect 3478 3135 3479 3139
rect 3483 3135 3484 3139
rect 3478 3134 3484 3135
rect 2751 3131 2757 3132
rect 2751 3130 2752 3131
rect 1862 3129 1868 3130
rect 610 3127 616 3128
rect 610 3123 611 3127
rect 615 3126 616 3127
rect 615 3124 718 3126
rect 1862 3125 1863 3129
rect 1867 3125 1868 3129
rect 2713 3128 2752 3130
rect 2751 3127 2752 3128
rect 2756 3127 2757 3131
rect 2751 3126 2757 3127
rect 3450 3131 3456 3132
rect 3450 3127 3451 3131
rect 3455 3130 3456 3131
rect 3455 3128 3497 3130
rect 3574 3129 3580 3130
rect 3455 3127 3456 3128
rect 3450 3126 3456 3127
rect 1862 3124 1868 3125
rect 3574 3125 3575 3129
rect 3579 3125 3580 3129
rect 3574 3124 3580 3125
rect 615 3123 616 3124
rect 610 3122 616 3123
rect 134 3119 140 3120
rect 134 3115 135 3119
rect 139 3115 140 3119
rect 134 3114 140 3115
rect 262 3119 268 3120
rect 262 3115 263 3119
rect 267 3115 268 3119
rect 262 3114 268 3115
rect 398 3119 404 3120
rect 398 3115 399 3119
rect 403 3115 404 3119
rect 398 3114 404 3115
rect 526 3119 532 3120
rect 526 3115 527 3119
rect 531 3115 532 3119
rect 526 3114 532 3115
rect 646 3119 652 3120
rect 646 3115 647 3119
rect 651 3115 652 3119
rect 646 3114 652 3115
rect 254 3111 260 3112
rect 110 3109 116 3110
rect 110 3105 111 3109
rect 115 3105 116 3109
rect 254 3107 255 3111
rect 259 3110 260 3111
rect 716 3110 718 3124
rect 758 3119 764 3120
rect 758 3115 759 3119
rect 763 3115 764 3119
rect 758 3114 764 3115
rect 862 3119 868 3120
rect 862 3115 863 3119
rect 867 3115 868 3119
rect 862 3114 868 3115
rect 966 3119 972 3120
rect 966 3115 967 3119
rect 971 3115 972 3119
rect 966 3114 972 3115
rect 1070 3119 1076 3120
rect 1070 3115 1071 3119
rect 1075 3115 1076 3119
rect 1070 3114 1076 3115
rect 1174 3119 1180 3120
rect 1174 3115 1175 3119
rect 1179 3115 1180 3119
rect 1174 3114 1180 3115
rect 1278 3119 1284 3120
rect 1278 3115 1279 3119
rect 1283 3115 1284 3119
rect 1278 3114 1284 3115
rect 1962 3115 1968 3116
rect 1862 3112 1868 3113
rect 1242 3111 1248 3112
rect 259 3108 281 3110
rect 716 3108 777 3110
rect 259 3107 260 3108
rect 254 3106 260 3107
rect 1242 3107 1243 3111
rect 1247 3110 1248 3111
rect 1247 3108 1297 3110
rect 1822 3109 1828 3110
rect 1247 3107 1248 3108
rect 1242 3106 1248 3107
rect 110 3104 116 3105
rect 1822 3105 1823 3109
rect 1827 3105 1828 3109
rect 1862 3108 1863 3112
rect 1867 3108 1868 3112
rect 1962 3111 1963 3115
rect 1967 3114 1968 3115
rect 2122 3115 2128 3116
rect 1967 3112 2081 3114
rect 1967 3111 1968 3112
rect 1962 3110 1968 3111
rect 2122 3111 2123 3115
rect 2127 3114 2128 3115
rect 2274 3115 2280 3116
rect 2127 3112 2233 3114
rect 2127 3111 2128 3112
rect 2122 3110 2128 3111
rect 2274 3111 2275 3115
rect 2279 3114 2280 3115
rect 2426 3115 2432 3116
rect 2279 3112 2385 3114
rect 2279 3111 2280 3112
rect 2274 3110 2280 3111
rect 2426 3111 2427 3115
rect 2431 3114 2432 3115
rect 2911 3115 2917 3116
rect 2911 3114 2912 3115
rect 2431 3112 2537 3114
rect 2853 3112 2912 3114
rect 2431 3111 2432 3112
rect 2426 3110 2432 3111
rect 2911 3111 2912 3112
rect 2916 3111 2917 3115
rect 3031 3115 3037 3116
rect 3031 3114 3032 3115
rect 2981 3112 3032 3114
rect 2911 3110 2917 3111
rect 3031 3111 3032 3112
rect 3036 3111 3037 3115
rect 3118 3115 3124 3116
rect 3118 3114 3119 3115
rect 3101 3112 3119 3114
rect 3031 3110 3037 3111
rect 3118 3111 3119 3112
rect 3123 3111 3124 3115
rect 3263 3115 3269 3116
rect 3263 3114 3264 3115
rect 3221 3112 3264 3114
rect 3118 3110 3124 3111
rect 3263 3111 3264 3112
rect 3268 3111 3269 3115
rect 3375 3115 3381 3116
rect 3375 3114 3376 3115
rect 3333 3112 3376 3114
rect 3263 3110 3269 3111
rect 3375 3111 3376 3112
rect 3380 3111 3381 3115
rect 3471 3115 3477 3116
rect 3471 3114 3472 3115
rect 3445 3112 3472 3114
rect 3375 3110 3381 3111
rect 3471 3111 3472 3112
rect 3476 3111 3477 3115
rect 3471 3110 3477 3111
rect 3574 3112 3580 3113
rect 1862 3107 1868 3108
rect 3574 3108 3575 3112
rect 3579 3108 3580 3112
rect 3574 3107 3580 3108
rect 1822 3104 1828 3105
rect 2062 3099 2068 3100
rect 255 3095 261 3096
rect 255 3094 256 3095
rect 110 3092 116 3093
rect 197 3092 256 3094
rect 110 3088 111 3092
rect 115 3088 116 3092
rect 255 3091 256 3092
rect 260 3091 261 3095
rect 519 3095 525 3096
rect 519 3094 520 3095
rect 461 3092 520 3094
rect 255 3090 261 3091
rect 519 3091 520 3092
rect 524 3091 525 3095
rect 639 3095 645 3096
rect 639 3094 640 3095
rect 589 3092 640 3094
rect 519 3090 525 3091
rect 639 3091 640 3092
rect 644 3091 645 3095
rect 751 3095 757 3096
rect 751 3094 752 3095
rect 709 3092 752 3094
rect 639 3090 645 3091
rect 751 3091 752 3092
rect 756 3091 757 3095
rect 959 3095 965 3096
rect 959 3094 960 3095
rect 925 3092 960 3094
rect 751 3090 757 3091
rect 959 3091 960 3092
rect 964 3091 965 3095
rect 1063 3095 1069 3096
rect 1063 3094 1064 3095
rect 1029 3092 1064 3094
rect 959 3090 965 3091
rect 1063 3091 1064 3092
rect 1068 3091 1069 3095
rect 1167 3095 1173 3096
rect 1167 3094 1168 3095
rect 1133 3092 1168 3094
rect 1063 3090 1069 3091
rect 1167 3091 1168 3092
rect 1172 3091 1173 3095
rect 1263 3095 1269 3096
rect 1263 3094 1264 3095
rect 1237 3092 1264 3094
rect 1167 3090 1173 3091
rect 1263 3091 1264 3092
rect 1268 3091 1269 3095
rect 2062 3095 2063 3099
rect 2067 3095 2068 3099
rect 2062 3094 2068 3095
rect 2214 3099 2220 3100
rect 2214 3095 2215 3099
rect 2219 3095 2220 3099
rect 2214 3094 2220 3095
rect 2366 3099 2372 3100
rect 2366 3095 2367 3099
rect 2371 3095 2372 3099
rect 2366 3094 2372 3095
rect 2518 3099 2524 3100
rect 2518 3095 2519 3099
rect 2523 3095 2524 3099
rect 2518 3094 2524 3095
rect 2662 3099 2668 3100
rect 2662 3095 2663 3099
rect 2667 3095 2668 3099
rect 2662 3094 2668 3095
rect 2798 3099 2804 3100
rect 2798 3095 2799 3099
rect 2803 3095 2804 3099
rect 2798 3094 2804 3095
rect 2926 3099 2932 3100
rect 2926 3095 2927 3099
rect 2931 3095 2932 3099
rect 2926 3094 2932 3095
rect 3046 3099 3052 3100
rect 3046 3095 3047 3099
rect 3051 3095 3052 3099
rect 3046 3094 3052 3095
rect 3166 3099 3172 3100
rect 3166 3095 3167 3099
rect 3171 3095 3172 3099
rect 3166 3094 3172 3095
rect 3278 3099 3284 3100
rect 3278 3095 3279 3099
rect 3283 3095 3284 3099
rect 3278 3094 3284 3095
rect 3390 3099 3396 3100
rect 3390 3095 3391 3099
rect 3395 3095 3396 3099
rect 3390 3094 3396 3095
rect 3486 3099 3492 3100
rect 3486 3095 3487 3099
rect 3491 3095 3492 3099
rect 3486 3094 3492 3095
rect 1263 3090 1269 3091
rect 1822 3092 1828 3093
rect 110 3087 116 3088
rect 1822 3088 1823 3092
rect 1827 3088 1828 3092
rect 1822 3087 1828 3088
rect 2071 3087 2077 3088
rect 2071 3083 2072 3087
rect 2076 3086 2077 3087
rect 2122 3087 2128 3088
rect 2122 3086 2123 3087
rect 2076 3084 2123 3086
rect 2076 3083 2077 3084
rect 2071 3082 2077 3083
rect 2122 3083 2123 3084
rect 2127 3083 2128 3087
rect 2122 3082 2128 3083
rect 2223 3087 2229 3088
rect 2223 3083 2224 3087
rect 2228 3086 2229 3087
rect 2274 3087 2280 3088
rect 2274 3086 2275 3087
rect 2228 3084 2275 3086
rect 2228 3083 2229 3084
rect 2223 3082 2229 3083
rect 2274 3083 2275 3084
rect 2279 3083 2280 3087
rect 2274 3082 2280 3083
rect 2375 3087 2381 3088
rect 2375 3083 2376 3087
rect 2380 3086 2381 3087
rect 2426 3087 2432 3088
rect 2426 3086 2427 3087
rect 2380 3084 2427 3086
rect 2380 3083 2381 3084
rect 2375 3082 2381 3083
rect 2426 3083 2427 3084
rect 2431 3083 2432 3087
rect 2426 3082 2432 3083
rect 2527 3087 2536 3088
rect 2527 3083 2528 3087
rect 2535 3083 2536 3087
rect 2527 3082 2536 3083
rect 2670 3087 2677 3088
rect 2670 3083 2671 3087
rect 2676 3083 2677 3087
rect 2670 3082 2677 3083
rect 2807 3087 2813 3088
rect 2807 3083 2808 3087
rect 2812 3086 2813 3087
rect 2903 3087 2909 3088
rect 2903 3086 2904 3087
rect 2812 3084 2904 3086
rect 2812 3083 2813 3084
rect 2807 3082 2813 3083
rect 2903 3083 2904 3084
rect 2908 3083 2909 3087
rect 2903 3082 2909 3083
rect 2911 3087 2917 3088
rect 2911 3083 2912 3087
rect 2916 3086 2917 3087
rect 2935 3087 2941 3088
rect 2935 3086 2936 3087
rect 2916 3084 2936 3086
rect 2916 3083 2917 3084
rect 2911 3082 2917 3083
rect 2935 3083 2936 3084
rect 2940 3083 2941 3087
rect 2935 3082 2941 3083
rect 3031 3087 3037 3088
rect 3031 3083 3032 3087
rect 3036 3086 3037 3087
rect 3055 3087 3061 3088
rect 3055 3086 3056 3087
rect 3036 3084 3056 3086
rect 3036 3083 3037 3084
rect 3031 3082 3037 3083
rect 3055 3083 3056 3084
rect 3060 3083 3061 3087
rect 3055 3082 3061 3083
rect 3175 3087 3184 3088
rect 3175 3083 3176 3087
rect 3183 3083 3184 3087
rect 3175 3082 3184 3083
rect 3263 3087 3269 3088
rect 3263 3083 3264 3087
rect 3268 3086 3269 3087
rect 3287 3087 3293 3088
rect 3287 3086 3288 3087
rect 3268 3084 3288 3086
rect 3268 3083 3269 3084
rect 3263 3082 3269 3083
rect 3287 3083 3288 3084
rect 3292 3083 3293 3087
rect 3287 3082 3293 3083
rect 3375 3087 3381 3088
rect 3375 3083 3376 3087
rect 3380 3086 3381 3087
rect 3399 3087 3405 3088
rect 3399 3086 3400 3087
rect 3380 3084 3400 3086
rect 3380 3083 3381 3084
rect 3375 3082 3381 3083
rect 3399 3083 3400 3084
rect 3404 3083 3405 3087
rect 3399 3082 3405 3083
rect 3471 3087 3477 3088
rect 3471 3083 3472 3087
rect 3476 3086 3477 3087
rect 3495 3087 3501 3088
rect 3495 3086 3496 3087
rect 3476 3084 3496 3086
rect 3476 3083 3477 3084
rect 3471 3082 3477 3083
rect 3495 3083 3496 3084
rect 3500 3083 3501 3087
rect 3495 3082 3501 3083
rect 142 3079 148 3080
rect 142 3075 143 3079
rect 147 3075 148 3079
rect 142 3074 148 3075
rect 270 3079 276 3080
rect 270 3075 271 3079
rect 275 3075 276 3079
rect 270 3074 276 3075
rect 406 3079 412 3080
rect 406 3075 407 3079
rect 411 3075 412 3079
rect 406 3074 412 3075
rect 534 3079 540 3080
rect 534 3075 535 3079
rect 539 3075 540 3079
rect 534 3074 540 3075
rect 654 3079 660 3080
rect 654 3075 655 3079
rect 659 3075 660 3079
rect 654 3074 660 3075
rect 766 3079 772 3080
rect 766 3075 767 3079
rect 771 3075 772 3079
rect 766 3074 772 3075
rect 870 3079 876 3080
rect 870 3075 871 3079
rect 875 3075 876 3079
rect 870 3074 876 3075
rect 974 3079 980 3080
rect 974 3075 975 3079
rect 979 3075 980 3079
rect 974 3074 980 3075
rect 1078 3079 1084 3080
rect 1078 3075 1079 3079
rect 1083 3075 1084 3079
rect 1078 3074 1084 3075
rect 1182 3079 1188 3080
rect 1182 3075 1183 3079
rect 1187 3075 1188 3079
rect 1182 3074 1188 3075
rect 1286 3079 1292 3080
rect 1286 3075 1287 3079
rect 1291 3075 1292 3079
rect 3450 3079 3456 3080
rect 3450 3078 3451 3079
rect 1286 3074 1292 3075
rect 3432 3076 3451 3078
rect 1959 3071 1968 3072
rect 151 3067 160 3068
rect 151 3063 152 3067
rect 159 3063 160 3067
rect 151 3062 160 3063
rect 255 3067 261 3068
rect 255 3063 256 3067
rect 260 3066 261 3067
rect 279 3067 285 3068
rect 279 3066 280 3067
rect 260 3064 280 3066
rect 260 3063 261 3064
rect 255 3062 261 3063
rect 279 3063 280 3064
rect 284 3063 285 3067
rect 279 3062 285 3063
rect 415 3067 421 3068
rect 415 3063 416 3067
rect 420 3066 421 3067
rect 426 3067 432 3068
rect 426 3066 427 3067
rect 420 3064 427 3066
rect 420 3063 421 3064
rect 415 3062 421 3063
rect 426 3063 427 3064
rect 431 3063 432 3067
rect 426 3062 432 3063
rect 519 3067 525 3068
rect 519 3063 520 3067
rect 524 3066 525 3067
rect 543 3067 549 3068
rect 543 3066 544 3067
rect 524 3064 544 3066
rect 524 3063 525 3064
rect 519 3062 525 3063
rect 543 3063 544 3064
rect 548 3063 549 3067
rect 543 3062 549 3063
rect 639 3067 645 3068
rect 639 3063 640 3067
rect 644 3066 645 3067
rect 663 3067 669 3068
rect 663 3066 664 3067
rect 644 3064 664 3066
rect 644 3063 645 3064
rect 639 3062 645 3063
rect 663 3063 664 3064
rect 668 3063 669 3067
rect 663 3062 669 3063
rect 751 3067 757 3068
rect 751 3063 752 3067
rect 756 3066 757 3067
rect 775 3067 781 3068
rect 775 3066 776 3067
rect 756 3064 776 3066
rect 756 3063 757 3064
rect 751 3062 757 3063
rect 775 3063 776 3064
rect 780 3063 781 3067
rect 775 3062 781 3063
rect 879 3067 885 3068
rect 879 3063 880 3067
rect 884 3066 885 3067
rect 950 3067 956 3068
rect 950 3066 951 3067
rect 884 3064 951 3066
rect 884 3063 885 3064
rect 879 3062 885 3063
rect 950 3063 951 3064
rect 955 3063 956 3067
rect 950 3062 956 3063
rect 959 3067 965 3068
rect 959 3063 960 3067
rect 964 3066 965 3067
rect 983 3067 989 3068
rect 983 3066 984 3067
rect 964 3064 984 3066
rect 964 3063 965 3064
rect 959 3062 965 3063
rect 983 3063 984 3064
rect 988 3063 989 3067
rect 983 3062 989 3063
rect 1063 3067 1069 3068
rect 1063 3063 1064 3067
rect 1068 3066 1069 3067
rect 1087 3067 1093 3068
rect 1087 3066 1088 3067
rect 1068 3064 1088 3066
rect 1068 3063 1069 3064
rect 1063 3062 1069 3063
rect 1087 3063 1088 3064
rect 1092 3063 1093 3067
rect 1087 3062 1093 3063
rect 1167 3067 1173 3068
rect 1167 3063 1168 3067
rect 1172 3066 1173 3067
rect 1191 3067 1197 3068
rect 1191 3066 1192 3067
rect 1172 3064 1192 3066
rect 1172 3063 1173 3064
rect 1167 3062 1173 3063
rect 1191 3063 1192 3064
rect 1196 3063 1197 3067
rect 1191 3062 1197 3063
rect 1263 3067 1269 3068
rect 1263 3063 1264 3067
rect 1268 3066 1269 3067
rect 1295 3067 1301 3068
rect 1295 3066 1296 3067
rect 1268 3064 1296 3066
rect 1268 3063 1269 3064
rect 1263 3062 1269 3063
rect 1295 3063 1296 3064
rect 1300 3063 1301 3067
rect 1959 3067 1960 3071
rect 1967 3067 1968 3071
rect 1959 3066 1968 3067
rect 2042 3071 2048 3072
rect 2042 3067 2043 3071
rect 2047 3070 2048 3071
rect 2087 3071 2093 3072
rect 2087 3070 2088 3071
rect 2047 3068 2088 3070
rect 2047 3067 2048 3068
rect 2042 3066 2048 3067
rect 2087 3067 2088 3068
rect 2092 3067 2093 3071
rect 2087 3066 2093 3067
rect 2151 3071 2157 3072
rect 2151 3067 2152 3071
rect 2156 3070 2157 3071
rect 2223 3071 2229 3072
rect 2223 3070 2224 3071
rect 2156 3068 2224 3070
rect 2156 3067 2157 3068
rect 2151 3066 2157 3067
rect 2223 3067 2224 3068
rect 2228 3067 2229 3071
rect 2223 3066 2229 3067
rect 2295 3071 2301 3072
rect 2295 3067 2296 3071
rect 2300 3070 2301 3071
rect 2375 3071 2381 3072
rect 2375 3070 2376 3071
rect 2300 3068 2376 3070
rect 2300 3067 2301 3068
rect 2295 3066 2301 3067
rect 2375 3067 2376 3068
rect 2380 3067 2381 3071
rect 2375 3066 2381 3067
rect 2455 3071 2461 3072
rect 2455 3067 2456 3071
rect 2460 3070 2461 3071
rect 2535 3071 2541 3072
rect 2535 3070 2536 3071
rect 2460 3068 2536 3070
rect 2460 3067 2461 3068
rect 2455 3066 2461 3067
rect 2535 3067 2536 3068
rect 2540 3067 2541 3071
rect 2535 3066 2541 3067
rect 2687 3071 2693 3072
rect 2687 3067 2688 3071
rect 2692 3070 2693 3071
rect 2766 3071 2772 3072
rect 2766 3070 2767 3071
rect 2692 3068 2767 3070
rect 2692 3067 2693 3068
rect 2687 3066 2693 3067
rect 2766 3067 2767 3068
rect 2771 3067 2772 3071
rect 2766 3066 2772 3067
rect 2839 3071 2845 3072
rect 2839 3067 2840 3071
rect 2844 3070 2845 3071
rect 2866 3071 2872 3072
rect 2866 3070 2867 3071
rect 2844 3068 2867 3070
rect 2844 3067 2845 3068
rect 2839 3066 2845 3067
rect 2866 3067 2867 3068
rect 2871 3067 2872 3071
rect 2866 3066 2872 3067
rect 2983 3071 2989 3072
rect 2983 3067 2984 3071
rect 2988 3070 2989 3071
rect 3047 3071 3053 3072
rect 3047 3070 3048 3071
rect 2988 3068 3048 3070
rect 2988 3067 2989 3068
rect 2983 3066 2989 3067
rect 3047 3067 3048 3068
rect 3052 3067 3053 3071
rect 3047 3066 3053 3067
rect 3118 3071 3125 3072
rect 3118 3067 3119 3071
rect 3124 3067 3125 3071
rect 3118 3066 3125 3067
rect 3247 3071 3253 3072
rect 3247 3067 3248 3071
rect 3252 3070 3253 3071
rect 3358 3071 3364 3072
rect 3358 3070 3359 3071
rect 3252 3068 3359 3070
rect 3252 3067 3253 3068
rect 3247 3066 3253 3067
rect 3358 3067 3359 3068
rect 3363 3067 3364 3071
rect 3358 3066 3364 3067
rect 3383 3071 3389 3072
rect 3383 3067 3384 3071
rect 3388 3070 3389 3071
rect 3432 3070 3434 3076
rect 3450 3075 3451 3076
rect 3455 3075 3456 3079
rect 3450 3074 3456 3075
rect 3388 3068 3434 3070
rect 3439 3071 3445 3072
rect 3388 3067 3389 3068
rect 3383 3066 3389 3067
rect 3439 3067 3440 3071
rect 3444 3070 3445 3071
rect 3495 3071 3501 3072
rect 3495 3070 3496 3071
rect 3444 3068 3496 3070
rect 3444 3067 3445 3068
rect 3439 3066 3445 3067
rect 3495 3067 3496 3068
rect 3500 3067 3501 3071
rect 3495 3066 3501 3067
rect 1295 3062 1301 3063
rect 1950 3061 1956 3062
rect 1950 3057 1951 3061
rect 1955 3057 1956 3061
rect 1950 3056 1956 3057
rect 2078 3061 2084 3062
rect 2078 3057 2079 3061
rect 2083 3057 2084 3061
rect 2078 3056 2084 3057
rect 2214 3061 2220 3062
rect 2214 3057 2215 3061
rect 2219 3057 2220 3061
rect 2214 3056 2220 3057
rect 2366 3061 2372 3062
rect 2366 3057 2367 3061
rect 2371 3057 2372 3061
rect 2366 3056 2372 3057
rect 2526 3061 2532 3062
rect 2526 3057 2527 3061
rect 2531 3057 2532 3061
rect 2526 3056 2532 3057
rect 2678 3061 2684 3062
rect 2678 3057 2679 3061
rect 2683 3057 2684 3061
rect 2678 3056 2684 3057
rect 2830 3061 2836 3062
rect 2830 3057 2831 3061
rect 2835 3057 2836 3061
rect 2830 3056 2836 3057
rect 2974 3061 2980 3062
rect 2974 3057 2975 3061
rect 2979 3057 2980 3061
rect 2974 3056 2980 3057
rect 3110 3061 3116 3062
rect 3110 3057 3111 3061
rect 3115 3057 3116 3061
rect 3110 3056 3116 3057
rect 3238 3061 3244 3062
rect 3238 3057 3239 3061
rect 3243 3057 3244 3061
rect 3238 3056 3244 3057
rect 3374 3061 3380 3062
rect 3374 3057 3375 3061
rect 3379 3057 3380 3061
rect 3374 3056 3380 3057
rect 3486 3061 3492 3062
rect 3486 3057 3487 3061
rect 3491 3057 3492 3061
rect 3486 3056 3492 3057
rect 151 3055 157 3056
rect 151 3051 152 3055
rect 156 3054 157 3055
rect 210 3055 216 3056
rect 210 3054 211 3055
rect 156 3052 211 3054
rect 156 3051 157 3052
rect 151 3050 157 3051
rect 210 3051 211 3052
rect 215 3051 216 3055
rect 210 3050 216 3051
rect 254 3055 261 3056
rect 254 3051 255 3055
rect 260 3051 261 3055
rect 254 3050 261 3051
rect 375 3055 381 3056
rect 375 3051 376 3055
rect 380 3054 381 3055
rect 438 3055 444 3056
rect 438 3054 439 3055
rect 380 3052 439 3054
rect 380 3051 381 3052
rect 375 3050 381 3051
rect 438 3051 439 3052
rect 443 3051 444 3055
rect 438 3050 444 3051
rect 495 3055 501 3056
rect 495 3051 496 3055
rect 500 3054 501 3055
rect 522 3055 528 3056
rect 522 3054 523 3055
rect 500 3052 523 3054
rect 500 3051 501 3052
rect 495 3050 501 3051
rect 522 3051 523 3052
rect 527 3051 528 3055
rect 522 3050 528 3051
rect 607 3055 616 3056
rect 607 3051 608 3055
rect 615 3051 616 3055
rect 607 3050 616 3051
rect 663 3055 669 3056
rect 663 3051 664 3055
rect 668 3054 669 3055
rect 711 3055 717 3056
rect 711 3054 712 3055
rect 668 3052 712 3054
rect 668 3051 669 3052
rect 663 3050 669 3051
rect 711 3051 712 3052
rect 716 3051 717 3055
rect 711 3050 717 3051
rect 767 3055 773 3056
rect 767 3051 768 3055
rect 772 3054 773 3055
rect 807 3055 813 3056
rect 807 3054 808 3055
rect 772 3052 808 3054
rect 772 3051 773 3052
rect 767 3050 773 3051
rect 807 3051 808 3052
rect 812 3051 813 3055
rect 807 3050 813 3051
rect 863 3055 869 3056
rect 863 3051 864 3055
rect 868 3054 869 3055
rect 903 3055 909 3056
rect 903 3054 904 3055
rect 868 3052 904 3054
rect 868 3051 869 3052
rect 863 3050 869 3051
rect 903 3051 904 3052
rect 908 3051 909 3055
rect 903 3050 909 3051
rect 998 3055 1005 3056
rect 998 3051 999 3055
rect 1004 3051 1005 3055
rect 998 3050 1005 3051
rect 1055 3055 1061 3056
rect 1055 3051 1056 3055
rect 1060 3054 1061 3055
rect 1095 3055 1101 3056
rect 1095 3054 1096 3055
rect 1060 3052 1096 3054
rect 1060 3051 1061 3052
rect 1055 3050 1061 3051
rect 1095 3051 1096 3052
rect 1100 3051 1101 3055
rect 1095 3050 1101 3051
rect 1146 3055 1152 3056
rect 1146 3051 1147 3055
rect 1151 3054 1152 3055
rect 1191 3055 1197 3056
rect 1191 3054 1192 3055
rect 1151 3052 1192 3054
rect 1151 3051 1152 3052
rect 1146 3050 1152 3051
rect 1191 3051 1192 3052
rect 1196 3051 1197 3055
rect 1191 3050 1197 3051
rect 1242 3055 1248 3056
rect 1242 3051 1243 3055
rect 1247 3054 1248 3055
rect 1295 3055 1301 3056
rect 1295 3054 1296 3055
rect 1247 3052 1296 3054
rect 1247 3051 1248 3052
rect 1242 3050 1248 3051
rect 1295 3051 1296 3052
rect 1300 3051 1301 3055
rect 1295 3050 1301 3051
rect 1862 3048 1868 3049
rect 3574 3048 3580 3049
rect 142 3045 148 3046
rect 142 3041 143 3045
rect 147 3041 148 3045
rect 142 3040 148 3041
rect 246 3045 252 3046
rect 246 3041 247 3045
rect 251 3041 252 3045
rect 246 3040 252 3041
rect 366 3045 372 3046
rect 366 3041 367 3045
rect 371 3041 372 3045
rect 366 3040 372 3041
rect 486 3045 492 3046
rect 486 3041 487 3045
rect 491 3041 492 3045
rect 486 3040 492 3041
rect 598 3045 604 3046
rect 598 3041 599 3045
rect 603 3041 604 3045
rect 598 3040 604 3041
rect 702 3045 708 3046
rect 702 3041 703 3045
rect 707 3041 708 3045
rect 702 3040 708 3041
rect 798 3045 804 3046
rect 798 3041 799 3045
rect 803 3041 804 3045
rect 798 3040 804 3041
rect 894 3045 900 3046
rect 894 3041 895 3045
rect 899 3041 900 3045
rect 894 3040 900 3041
rect 990 3045 996 3046
rect 990 3041 991 3045
rect 995 3041 996 3045
rect 990 3040 996 3041
rect 1086 3045 1092 3046
rect 1086 3041 1087 3045
rect 1091 3041 1092 3045
rect 1086 3040 1092 3041
rect 1182 3045 1188 3046
rect 1182 3041 1183 3045
rect 1187 3041 1188 3045
rect 1182 3040 1188 3041
rect 1286 3045 1292 3046
rect 1286 3041 1287 3045
rect 1291 3041 1292 3045
rect 1862 3044 1863 3048
rect 1867 3044 1868 3048
rect 2042 3047 2048 3048
rect 2042 3046 2043 3047
rect 2005 3044 2043 3046
rect 1862 3043 1868 3044
rect 2042 3043 2043 3044
rect 2047 3043 2048 3047
rect 2151 3047 2157 3048
rect 2151 3046 2152 3047
rect 2133 3044 2152 3046
rect 2042 3042 2048 3043
rect 2151 3043 2152 3044
rect 2156 3043 2157 3047
rect 2295 3047 2301 3048
rect 2295 3046 2296 3047
rect 2269 3044 2296 3046
rect 2151 3042 2157 3043
rect 2295 3043 2296 3044
rect 2300 3043 2301 3047
rect 2455 3047 2461 3048
rect 2455 3046 2456 3047
rect 2421 3044 2456 3046
rect 2295 3042 2301 3043
rect 2455 3043 2456 3044
rect 2460 3043 2461 3047
rect 3439 3047 3445 3048
rect 3439 3046 3440 3047
rect 3429 3044 3440 3046
rect 2455 3042 2461 3043
rect 2670 3043 2676 3044
rect 1286 3040 1292 3041
rect 2670 3039 2671 3043
rect 2675 3042 2676 3043
rect 2766 3043 2772 3044
rect 2675 3040 2697 3042
rect 2675 3039 2676 3040
rect 2670 3038 2676 3039
rect 2766 3039 2767 3043
rect 2771 3042 2772 3043
rect 3047 3043 3053 3044
rect 2771 3040 2849 3042
rect 2771 3039 2772 3040
rect 2766 3038 2772 3039
rect 3047 3039 3048 3043
rect 3052 3042 3053 3043
rect 3178 3043 3184 3044
rect 3052 3040 3129 3042
rect 3052 3039 3053 3040
rect 3047 3038 3053 3039
rect 3178 3039 3179 3043
rect 3183 3042 3184 3043
rect 3439 3043 3440 3044
rect 3444 3043 3445 3047
rect 3574 3044 3575 3048
rect 3579 3044 3580 3048
rect 3574 3043 3580 3044
rect 3439 3042 3445 3043
rect 3183 3040 3257 3042
rect 3183 3039 3184 3040
rect 3178 3038 3184 3039
rect 110 3032 116 3033
rect 1822 3032 1828 3033
rect 110 3028 111 3032
rect 115 3028 116 3032
rect 426 3031 432 3032
rect 426 3030 427 3031
rect 421 3028 427 3030
rect 110 3027 116 3028
rect 210 3027 216 3028
rect 210 3023 211 3027
rect 215 3026 216 3027
rect 426 3027 427 3028
rect 431 3027 432 3031
rect 663 3031 669 3032
rect 663 3030 664 3031
rect 653 3028 664 3030
rect 426 3026 432 3027
rect 438 3027 444 3028
rect 215 3024 265 3026
rect 215 3023 216 3024
rect 210 3022 216 3023
rect 438 3023 439 3027
rect 443 3026 444 3027
rect 663 3027 664 3028
rect 668 3027 669 3031
rect 767 3031 773 3032
rect 767 3030 768 3031
rect 757 3028 768 3030
rect 663 3026 669 3027
rect 767 3027 768 3028
rect 772 3027 773 3031
rect 863 3031 869 3032
rect 863 3030 864 3031
rect 853 3028 864 3030
rect 767 3026 773 3027
rect 863 3027 864 3028
rect 868 3027 869 3031
rect 1055 3031 1061 3032
rect 1055 3030 1056 3031
rect 1045 3028 1056 3030
rect 863 3026 869 3027
rect 1055 3027 1056 3028
rect 1060 3027 1061 3031
rect 1146 3031 1152 3032
rect 1146 3030 1147 3031
rect 1141 3028 1147 3030
rect 1055 3026 1061 3027
rect 1146 3027 1147 3028
rect 1151 3027 1152 3031
rect 1242 3031 1248 3032
rect 1242 3030 1243 3031
rect 1237 3028 1243 3030
rect 1146 3026 1152 3027
rect 1242 3027 1243 3028
rect 1247 3027 1248 3031
rect 1822 3028 1823 3032
rect 1827 3028 1828 3032
rect 1242 3026 1248 3027
rect 1250 3027 1256 3028
rect 1822 3027 1828 3028
rect 1862 3031 1868 3032
rect 1862 3027 1863 3031
rect 1867 3027 1868 3031
rect 2594 3031 2600 3032
rect 2594 3030 2595 3031
rect 2577 3028 2595 3030
rect 443 3024 505 3026
rect 443 3023 444 3024
rect 438 3022 444 3023
rect 1250 3023 1251 3027
rect 1255 3026 1256 3027
rect 1862 3026 1868 3027
rect 2594 3027 2595 3028
rect 2599 3027 2600 3031
rect 3574 3031 3580 3032
rect 2594 3026 2600 3027
rect 2913 3028 2985 3030
rect 1255 3024 1305 3026
rect 1255 3023 1256 3024
rect 1250 3022 1256 3023
rect 1942 3021 1948 3022
rect 1942 3017 1943 3021
rect 1947 3017 1948 3021
rect 1942 3016 1948 3017
rect 2070 3021 2076 3022
rect 2070 3017 2071 3021
rect 2075 3017 2076 3021
rect 2070 3016 2076 3017
rect 2206 3021 2212 3022
rect 2206 3017 2207 3021
rect 2211 3017 2212 3021
rect 2206 3016 2212 3017
rect 2358 3021 2364 3022
rect 2358 3017 2359 3021
rect 2363 3017 2364 3021
rect 2358 3016 2364 3017
rect 2518 3021 2524 3022
rect 2518 3017 2519 3021
rect 2523 3017 2524 3021
rect 2518 3016 2524 3017
rect 2670 3021 2676 3022
rect 2670 3017 2671 3021
rect 2675 3017 2676 3021
rect 2670 3016 2676 3017
rect 2822 3021 2828 3022
rect 2822 3017 2823 3021
rect 2827 3017 2828 3021
rect 2822 3016 2828 3017
rect 110 3015 116 3016
rect 110 3011 111 3015
rect 115 3011 116 3015
rect 110 3010 116 3011
rect 1822 3015 1828 3016
rect 1822 3011 1823 3015
rect 1827 3011 1828 3015
rect 1822 3010 1828 3011
rect 2706 3015 2712 3016
rect 2706 3011 2707 3015
rect 2711 3014 2712 3015
rect 2913 3014 2915 3028
rect 3574 3027 3575 3031
rect 3579 3027 3580 3031
rect 3574 3026 3580 3027
rect 2966 3021 2972 3022
rect 2966 3017 2967 3021
rect 2971 3017 2972 3021
rect 2966 3016 2972 3017
rect 3102 3021 3108 3022
rect 3102 3017 3103 3021
rect 3107 3017 3108 3021
rect 3102 3016 3108 3017
rect 3230 3021 3236 3022
rect 3230 3017 3231 3021
rect 3235 3017 3236 3021
rect 3230 3016 3236 3017
rect 3366 3021 3372 3022
rect 3366 3017 3367 3021
rect 3371 3017 3372 3021
rect 3366 3016 3372 3017
rect 3478 3021 3484 3022
rect 3478 3017 3479 3021
rect 3483 3017 3484 3021
rect 3478 3016 3484 3017
rect 2711 3012 2915 3014
rect 3498 3015 3504 3016
rect 2711 3011 2712 3012
rect 2706 3010 2712 3011
rect 3498 3011 3499 3015
rect 3503 3014 3504 3015
rect 3527 3015 3533 3016
rect 3527 3014 3528 3015
rect 3503 3012 3528 3014
rect 3503 3011 3504 3012
rect 3498 3010 3504 3011
rect 3527 3011 3528 3012
rect 3532 3011 3533 3015
rect 3527 3010 3533 3011
rect 134 3005 140 3006
rect 134 3001 135 3005
rect 139 3001 140 3005
rect 134 3000 140 3001
rect 238 3005 244 3006
rect 238 3001 239 3005
rect 243 3001 244 3005
rect 238 3000 244 3001
rect 358 3005 364 3006
rect 358 3001 359 3005
rect 363 3001 364 3005
rect 358 3000 364 3001
rect 478 3005 484 3006
rect 478 3001 479 3005
rect 483 3001 484 3005
rect 478 3000 484 3001
rect 590 3005 596 3006
rect 590 3001 591 3005
rect 595 3001 596 3005
rect 590 3000 596 3001
rect 694 3005 700 3006
rect 694 3001 695 3005
rect 699 3001 700 3005
rect 694 3000 700 3001
rect 790 3005 796 3006
rect 790 3001 791 3005
rect 795 3001 796 3005
rect 790 3000 796 3001
rect 886 3005 892 3006
rect 886 3001 887 3005
rect 891 3001 892 3005
rect 886 3000 892 3001
rect 982 3005 988 3006
rect 982 3001 983 3005
rect 987 3001 988 3005
rect 982 3000 988 3001
rect 1078 3005 1084 3006
rect 1078 3001 1079 3005
rect 1083 3001 1084 3005
rect 1078 3000 1084 3001
rect 1174 3005 1180 3006
rect 1174 3001 1175 3005
rect 1179 3001 1180 3005
rect 1174 3000 1180 3001
rect 1278 3005 1284 3006
rect 1278 3001 1279 3005
rect 1283 3001 1284 3005
rect 1278 3000 1284 3001
rect 154 2999 160 3000
rect 154 2995 155 2999
rect 159 2998 160 2999
rect 183 2999 189 3000
rect 183 2998 184 2999
rect 159 2996 184 2998
rect 159 2995 160 2996
rect 154 2994 160 2995
rect 183 2995 184 2996
rect 188 2995 189 2999
rect 183 2994 189 2995
rect 935 2999 941 3000
rect 935 2995 936 2999
rect 940 2998 941 2999
rect 946 2999 952 3000
rect 946 2998 947 2999
rect 940 2996 947 2998
rect 940 2995 941 2996
rect 935 2994 941 2995
rect 946 2995 947 2996
rect 951 2995 952 2999
rect 946 2994 952 2995
rect 1886 2987 1892 2988
rect 1886 2983 1887 2987
rect 1891 2983 1892 2987
rect 1886 2982 1892 2983
rect 1974 2987 1980 2988
rect 1974 2983 1975 2987
rect 1979 2983 1980 2987
rect 1974 2982 1980 2983
rect 2062 2987 2068 2988
rect 2062 2983 2063 2987
rect 2067 2983 2068 2987
rect 2062 2982 2068 2983
rect 2150 2987 2156 2988
rect 2150 2983 2151 2987
rect 2155 2983 2156 2987
rect 2150 2982 2156 2983
rect 2238 2987 2244 2988
rect 2238 2983 2239 2987
rect 2243 2983 2244 2987
rect 2238 2982 2244 2983
rect 2350 2987 2356 2988
rect 2350 2983 2351 2987
rect 2355 2983 2356 2987
rect 2350 2982 2356 2983
rect 2462 2987 2468 2988
rect 2462 2983 2463 2987
rect 2467 2983 2468 2987
rect 2462 2982 2468 2983
rect 2574 2987 2580 2988
rect 2574 2983 2575 2987
rect 2579 2983 2580 2987
rect 2574 2982 2580 2983
rect 2686 2987 2692 2988
rect 2686 2983 2687 2987
rect 2691 2983 2692 2987
rect 2686 2982 2692 2983
rect 2798 2987 2804 2988
rect 2798 2983 2799 2987
rect 2803 2983 2804 2987
rect 2798 2982 2804 2983
rect 2902 2987 2908 2988
rect 2902 2983 2903 2987
rect 2907 2983 2908 2987
rect 2902 2982 2908 2983
rect 3006 2987 3012 2988
rect 3006 2983 3007 2987
rect 3011 2983 3012 2987
rect 3006 2982 3012 2983
rect 3102 2987 3108 2988
rect 3102 2983 3103 2987
rect 3107 2983 3108 2987
rect 3102 2982 3108 2983
rect 3198 2987 3204 2988
rect 3198 2983 3199 2987
rect 3203 2983 3204 2987
rect 3198 2982 3204 2983
rect 3294 2987 3300 2988
rect 3294 2983 3295 2987
rect 3299 2983 3300 2987
rect 3294 2982 3300 2983
rect 3390 2987 3396 2988
rect 3390 2983 3391 2987
rect 3395 2983 3396 2987
rect 3390 2982 3396 2983
rect 3478 2987 3484 2988
rect 3478 2983 3479 2987
rect 3483 2983 3484 2987
rect 3478 2982 3484 2983
rect 2866 2979 2872 2980
rect 1862 2977 1868 2978
rect 1862 2973 1863 2977
rect 1867 2973 1868 2977
rect 2866 2975 2867 2979
rect 2871 2978 2872 2979
rect 3362 2979 3368 2980
rect 2871 2976 2921 2978
rect 2871 2975 2872 2976
rect 2866 2974 2872 2975
rect 3362 2975 3363 2979
rect 3367 2978 3368 2979
rect 3367 2976 3409 2978
rect 3574 2977 3580 2978
rect 3367 2975 3368 2976
rect 3362 2974 3368 2975
rect 1862 2972 1868 2973
rect 3574 2973 3575 2977
rect 3579 2973 3580 2977
rect 3574 2972 3580 2973
rect 134 2971 140 2972
rect 134 2967 135 2971
rect 139 2967 140 2971
rect 134 2966 140 2967
rect 286 2971 292 2972
rect 286 2967 287 2971
rect 291 2967 292 2971
rect 286 2966 292 2967
rect 454 2971 460 2972
rect 454 2967 455 2971
rect 459 2967 460 2971
rect 454 2966 460 2967
rect 622 2971 628 2972
rect 622 2967 623 2971
rect 627 2967 628 2971
rect 622 2966 628 2967
rect 782 2971 788 2972
rect 782 2967 783 2971
rect 787 2967 788 2971
rect 782 2966 788 2967
rect 926 2971 932 2972
rect 926 2967 927 2971
rect 931 2967 932 2971
rect 926 2966 932 2967
rect 1062 2971 1068 2972
rect 1062 2967 1063 2971
rect 1067 2967 1068 2971
rect 1062 2966 1068 2967
rect 1190 2971 1196 2972
rect 1190 2967 1191 2971
rect 1195 2967 1196 2971
rect 1190 2966 1196 2967
rect 1310 2971 1316 2972
rect 1310 2967 1311 2971
rect 1315 2967 1316 2971
rect 1310 2966 1316 2967
rect 1422 2971 1428 2972
rect 1422 2967 1423 2971
rect 1427 2967 1428 2971
rect 1422 2966 1428 2967
rect 1526 2971 1532 2972
rect 1526 2967 1527 2971
rect 1531 2967 1532 2971
rect 1526 2966 1532 2967
rect 1638 2971 1644 2972
rect 1638 2967 1639 2971
rect 1643 2967 1644 2971
rect 1638 2966 1644 2967
rect 1726 2971 1732 2972
rect 1726 2967 1727 2971
rect 1731 2967 1732 2971
rect 1726 2966 1732 2967
rect 522 2963 528 2964
rect 522 2962 523 2963
rect 110 2961 116 2962
rect 110 2957 111 2961
rect 115 2957 116 2961
rect 513 2960 523 2962
rect 522 2959 523 2960
rect 527 2959 528 2963
rect 522 2958 528 2959
rect 690 2963 696 2964
rect 690 2959 691 2963
rect 695 2962 696 2963
rect 998 2963 1004 2964
rect 998 2962 999 2963
rect 695 2960 801 2962
rect 985 2960 999 2962
rect 695 2959 696 2960
rect 690 2958 696 2959
rect 998 2959 999 2960
rect 1003 2959 1004 2963
rect 1870 2963 1876 2964
rect 998 2958 1004 2959
rect 1822 2961 1828 2962
rect 110 2956 116 2957
rect 1822 2957 1823 2961
rect 1827 2957 1828 2961
rect 1822 2956 1828 2957
rect 1862 2960 1868 2961
rect 1862 2956 1863 2960
rect 1867 2956 1868 2960
rect 1870 2959 1871 2963
rect 1875 2962 1876 2963
rect 1954 2963 1960 2964
rect 1875 2960 1913 2962
rect 1875 2959 1876 2960
rect 1870 2958 1876 2959
rect 1954 2959 1955 2963
rect 1959 2962 1960 2963
rect 2042 2963 2048 2964
rect 1959 2960 2001 2962
rect 1959 2959 1960 2960
rect 1954 2958 1960 2959
rect 2042 2959 2043 2963
rect 2047 2962 2048 2963
rect 2130 2963 2136 2964
rect 2047 2960 2089 2962
rect 2047 2959 2048 2960
rect 2042 2958 2048 2959
rect 2130 2959 2131 2963
rect 2135 2962 2136 2963
rect 2218 2963 2224 2964
rect 2135 2960 2177 2962
rect 2135 2959 2136 2960
rect 2130 2958 2136 2959
rect 2218 2959 2219 2963
rect 2223 2962 2224 2963
rect 2306 2963 2312 2964
rect 2223 2960 2265 2962
rect 2223 2959 2224 2960
rect 2218 2958 2224 2959
rect 2306 2959 2307 2963
rect 2311 2962 2312 2963
rect 2418 2963 2424 2964
rect 2311 2960 2377 2962
rect 2311 2959 2312 2960
rect 2306 2958 2312 2959
rect 2418 2959 2419 2963
rect 2423 2962 2424 2963
rect 2530 2963 2536 2964
rect 2423 2960 2489 2962
rect 2423 2959 2424 2960
rect 2418 2958 2424 2959
rect 2530 2959 2531 2963
rect 2535 2962 2536 2963
rect 2791 2963 2797 2964
rect 2791 2962 2792 2963
rect 2535 2960 2601 2962
rect 2749 2960 2792 2962
rect 2535 2959 2536 2960
rect 2530 2958 2536 2959
rect 2791 2959 2792 2960
rect 2796 2959 2797 2963
rect 2895 2963 2901 2964
rect 2895 2962 2896 2963
rect 2861 2960 2896 2962
rect 2791 2958 2797 2959
rect 2895 2959 2896 2960
rect 2900 2959 2901 2963
rect 3095 2963 3101 2964
rect 3095 2962 3096 2963
rect 3069 2960 3096 2962
rect 2895 2958 2901 2959
rect 3095 2959 3096 2960
rect 3100 2959 3101 2963
rect 3191 2963 3197 2964
rect 3191 2962 3192 2963
rect 3165 2960 3192 2962
rect 3095 2958 3101 2959
rect 3191 2959 3192 2960
rect 3196 2959 3197 2963
rect 3287 2963 3293 2964
rect 3287 2962 3288 2963
rect 3261 2960 3288 2962
rect 3191 2958 3197 2959
rect 3287 2959 3288 2960
rect 3292 2959 3293 2963
rect 3383 2963 3389 2964
rect 3383 2962 3384 2963
rect 3357 2960 3384 2962
rect 3287 2958 3293 2959
rect 3383 2959 3384 2960
rect 3388 2959 3389 2963
rect 3383 2958 3389 2959
rect 3471 2963 3477 2964
rect 3471 2959 3472 2963
rect 3476 2962 3477 2963
rect 3476 2960 3505 2962
rect 3574 2960 3580 2961
rect 3476 2959 3477 2960
rect 3471 2958 3477 2959
rect 1862 2955 1868 2956
rect 3574 2956 3575 2960
rect 3579 2956 3580 2960
rect 3574 2955 3580 2956
rect 279 2947 285 2948
rect 279 2946 280 2947
rect 110 2944 116 2945
rect 197 2944 280 2946
rect 110 2940 111 2944
rect 115 2940 116 2944
rect 279 2943 280 2944
rect 284 2943 285 2947
rect 354 2947 360 2948
rect 354 2946 355 2947
rect 349 2944 355 2946
rect 279 2942 285 2943
rect 354 2943 355 2944
rect 359 2943 360 2947
rect 775 2947 781 2948
rect 775 2946 776 2947
rect 685 2944 776 2946
rect 354 2942 360 2943
rect 775 2943 776 2944
rect 780 2943 781 2947
rect 1183 2947 1189 2948
rect 1183 2946 1184 2947
rect 1125 2944 1184 2946
rect 775 2942 781 2943
rect 1183 2943 1184 2944
rect 1188 2943 1189 2947
rect 1303 2947 1309 2948
rect 1303 2946 1304 2947
rect 1253 2944 1304 2946
rect 1183 2942 1189 2943
rect 1303 2943 1304 2944
rect 1308 2943 1309 2947
rect 1406 2947 1412 2948
rect 1406 2946 1407 2947
rect 1373 2944 1407 2946
rect 1303 2942 1309 2943
rect 1406 2943 1407 2944
rect 1411 2943 1412 2947
rect 1406 2942 1412 2943
rect 1414 2947 1420 2948
rect 1414 2943 1415 2947
rect 1419 2946 1420 2947
rect 1490 2947 1496 2948
rect 1419 2944 1449 2946
rect 1419 2943 1420 2944
rect 1414 2942 1420 2943
rect 1490 2943 1491 2947
rect 1495 2946 1496 2947
rect 1594 2947 1600 2948
rect 1495 2944 1553 2946
rect 1495 2943 1496 2944
rect 1490 2942 1496 2943
rect 1594 2943 1595 2947
rect 1599 2946 1600 2947
rect 1711 2947 1717 2948
rect 1599 2944 1665 2946
rect 1599 2943 1600 2944
rect 1594 2942 1600 2943
rect 1711 2943 1712 2947
rect 1716 2946 1717 2947
rect 1894 2947 1900 2948
rect 1716 2944 1753 2946
rect 1822 2944 1828 2945
rect 1716 2943 1717 2944
rect 1711 2942 1717 2943
rect 110 2939 116 2940
rect 1822 2940 1823 2944
rect 1827 2940 1828 2944
rect 1894 2943 1895 2947
rect 1899 2943 1900 2947
rect 1894 2942 1900 2943
rect 1982 2947 1988 2948
rect 1982 2943 1983 2947
rect 1987 2943 1988 2947
rect 1982 2942 1988 2943
rect 2070 2947 2076 2948
rect 2070 2943 2071 2947
rect 2075 2943 2076 2947
rect 2070 2942 2076 2943
rect 2158 2947 2164 2948
rect 2158 2943 2159 2947
rect 2163 2943 2164 2947
rect 2158 2942 2164 2943
rect 2246 2947 2252 2948
rect 2246 2943 2247 2947
rect 2251 2943 2252 2947
rect 2246 2942 2252 2943
rect 2358 2947 2364 2948
rect 2358 2943 2359 2947
rect 2363 2943 2364 2947
rect 2358 2942 2364 2943
rect 2470 2947 2476 2948
rect 2470 2943 2471 2947
rect 2475 2943 2476 2947
rect 2470 2942 2476 2943
rect 2582 2947 2588 2948
rect 2582 2943 2583 2947
rect 2587 2943 2588 2947
rect 2582 2942 2588 2943
rect 2694 2947 2700 2948
rect 2694 2943 2695 2947
rect 2699 2943 2700 2947
rect 2694 2942 2700 2943
rect 2806 2947 2812 2948
rect 2806 2943 2807 2947
rect 2811 2943 2812 2947
rect 2806 2942 2812 2943
rect 2910 2947 2916 2948
rect 2910 2943 2911 2947
rect 2915 2943 2916 2947
rect 2910 2942 2916 2943
rect 3014 2947 3020 2948
rect 3014 2943 3015 2947
rect 3019 2943 3020 2947
rect 3014 2942 3020 2943
rect 3110 2947 3116 2948
rect 3110 2943 3111 2947
rect 3115 2943 3116 2947
rect 3110 2942 3116 2943
rect 3206 2947 3212 2948
rect 3206 2943 3207 2947
rect 3211 2943 3212 2947
rect 3206 2942 3212 2943
rect 3302 2947 3308 2948
rect 3302 2943 3303 2947
rect 3307 2943 3308 2947
rect 3302 2942 3308 2943
rect 3398 2947 3404 2948
rect 3398 2943 3399 2947
rect 3403 2943 3404 2947
rect 3398 2942 3404 2943
rect 3486 2947 3492 2948
rect 3486 2943 3487 2947
rect 3491 2943 3492 2947
rect 3486 2942 3492 2943
rect 1822 2939 1828 2940
rect 1903 2935 1909 2936
rect 142 2931 148 2932
rect 142 2927 143 2931
rect 147 2927 148 2931
rect 142 2926 148 2927
rect 294 2931 300 2932
rect 294 2927 295 2931
rect 299 2927 300 2931
rect 294 2926 300 2927
rect 462 2931 468 2932
rect 462 2927 463 2931
rect 467 2927 468 2931
rect 462 2926 468 2927
rect 630 2931 636 2932
rect 630 2927 631 2931
rect 635 2927 636 2931
rect 630 2926 636 2927
rect 790 2931 796 2932
rect 790 2927 791 2931
rect 795 2927 796 2931
rect 790 2926 796 2927
rect 934 2931 940 2932
rect 934 2927 935 2931
rect 939 2927 940 2931
rect 934 2926 940 2927
rect 1070 2931 1076 2932
rect 1070 2927 1071 2931
rect 1075 2927 1076 2931
rect 1070 2926 1076 2927
rect 1198 2931 1204 2932
rect 1198 2927 1199 2931
rect 1203 2927 1204 2931
rect 1198 2926 1204 2927
rect 1318 2931 1324 2932
rect 1318 2927 1319 2931
rect 1323 2927 1324 2931
rect 1318 2926 1324 2927
rect 1430 2931 1436 2932
rect 1430 2927 1431 2931
rect 1435 2927 1436 2931
rect 1430 2926 1436 2927
rect 1534 2931 1540 2932
rect 1534 2927 1535 2931
rect 1539 2927 1540 2931
rect 1534 2926 1540 2927
rect 1646 2931 1652 2932
rect 1646 2927 1647 2931
rect 1651 2927 1652 2931
rect 1646 2926 1652 2927
rect 1734 2931 1740 2932
rect 1734 2927 1735 2931
rect 1739 2927 1740 2931
rect 1903 2931 1904 2935
rect 1908 2934 1909 2935
rect 1954 2935 1960 2936
rect 1954 2934 1955 2935
rect 1908 2932 1955 2934
rect 1908 2931 1909 2932
rect 1903 2930 1909 2931
rect 1954 2931 1955 2932
rect 1959 2931 1960 2935
rect 1954 2930 1960 2931
rect 1991 2935 1997 2936
rect 1991 2931 1992 2935
rect 1996 2934 1997 2935
rect 2042 2935 2048 2936
rect 2042 2934 2043 2935
rect 1996 2932 2043 2934
rect 1996 2931 1997 2932
rect 1991 2930 1997 2931
rect 2042 2931 2043 2932
rect 2047 2931 2048 2935
rect 2042 2930 2048 2931
rect 2079 2935 2085 2936
rect 2079 2931 2080 2935
rect 2084 2934 2085 2935
rect 2130 2935 2136 2936
rect 2130 2934 2131 2935
rect 2084 2932 2131 2934
rect 2084 2931 2085 2932
rect 2079 2930 2085 2931
rect 2130 2931 2131 2932
rect 2135 2931 2136 2935
rect 2130 2930 2136 2931
rect 2167 2935 2173 2936
rect 2167 2931 2168 2935
rect 2172 2934 2173 2935
rect 2218 2935 2224 2936
rect 2218 2934 2219 2935
rect 2172 2932 2219 2934
rect 2172 2931 2173 2932
rect 2167 2930 2173 2931
rect 2218 2931 2219 2932
rect 2223 2931 2224 2935
rect 2218 2930 2224 2931
rect 2255 2935 2261 2936
rect 2255 2931 2256 2935
rect 2260 2934 2261 2935
rect 2306 2935 2312 2936
rect 2306 2934 2307 2935
rect 2260 2932 2307 2934
rect 2260 2931 2261 2932
rect 2255 2930 2261 2931
rect 2306 2931 2307 2932
rect 2311 2931 2312 2935
rect 2306 2930 2312 2931
rect 2367 2935 2373 2936
rect 2367 2931 2368 2935
rect 2372 2934 2373 2935
rect 2418 2935 2424 2936
rect 2418 2934 2419 2935
rect 2372 2932 2419 2934
rect 2372 2931 2373 2932
rect 2367 2930 2373 2931
rect 2418 2931 2419 2932
rect 2423 2931 2424 2935
rect 2418 2930 2424 2931
rect 2479 2935 2485 2936
rect 2479 2931 2480 2935
rect 2484 2934 2485 2935
rect 2530 2935 2536 2936
rect 2530 2934 2531 2935
rect 2484 2932 2531 2934
rect 2484 2931 2485 2932
rect 2479 2930 2485 2931
rect 2530 2931 2531 2932
rect 2535 2931 2536 2935
rect 2530 2930 2536 2931
rect 2591 2935 2600 2936
rect 2591 2931 2592 2935
rect 2599 2931 2600 2935
rect 2591 2930 2600 2931
rect 2703 2935 2712 2936
rect 2703 2931 2704 2935
rect 2711 2931 2712 2935
rect 2703 2930 2712 2931
rect 2791 2935 2797 2936
rect 2791 2931 2792 2935
rect 2796 2934 2797 2935
rect 2815 2935 2821 2936
rect 2815 2934 2816 2935
rect 2796 2932 2816 2934
rect 2796 2931 2797 2932
rect 2791 2930 2797 2931
rect 2815 2931 2816 2932
rect 2820 2931 2821 2935
rect 2815 2930 2821 2931
rect 2919 2935 2925 2936
rect 2919 2931 2920 2935
rect 2924 2934 2925 2935
rect 2954 2935 2960 2936
rect 2954 2934 2955 2935
rect 2924 2932 2955 2934
rect 2924 2931 2925 2932
rect 2919 2930 2925 2931
rect 2954 2931 2955 2932
rect 2959 2931 2960 2935
rect 3023 2935 3029 2936
rect 3023 2934 3024 2935
rect 2954 2930 2960 2931
rect 2964 2932 3024 2934
rect 1734 2926 1740 2927
rect 2895 2927 2901 2928
rect 2895 2923 2896 2927
rect 2900 2926 2901 2927
rect 2964 2926 2966 2932
rect 3023 2931 3024 2932
rect 3028 2931 3029 2935
rect 3023 2930 3029 2931
rect 3095 2935 3101 2936
rect 3095 2931 3096 2935
rect 3100 2934 3101 2935
rect 3119 2935 3125 2936
rect 3119 2934 3120 2935
rect 3100 2932 3120 2934
rect 3100 2931 3101 2932
rect 3095 2930 3101 2931
rect 3119 2931 3120 2932
rect 3124 2931 3125 2935
rect 3119 2930 3125 2931
rect 3191 2935 3197 2936
rect 3191 2931 3192 2935
rect 3196 2934 3197 2935
rect 3215 2935 3221 2936
rect 3215 2934 3216 2935
rect 3196 2932 3216 2934
rect 3196 2931 3197 2932
rect 3191 2930 3197 2931
rect 3215 2931 3216 2932
rect 3220 2931 3221 2935
rect 3215 2930 3221 2931
rect 3287 2935 3293 2936
rect 3287 2931 3288 2935
rect 3292 2934 3293 2935
rect 3311 2935 3317 2936
rect 3311 2934 3312 2935
rect 3292 2932 3312 2934
rect 3292 2931 3293 2932
rect 3287 2930 3293 2931
rect 3311 2931 3312 2932
rect 3316 2931 3317 2935
rect 3311 2930 3317 2931
rect 3383 2935 3389 2936
rect 3383 2931 3384 2935
rect 3388 2934 3389 2935
rect 3407 2935 3413 2936
rect 3407 2934 3408 2935
rect 3388 2932 3408 2934
rect 3388 2931 3389 2932
rect 3383 2930 3389 2931
rect 3407 2931 3408 2932
rect 3412 2931 3413 2935
rect 3407 2930 3413 2931
rect 3495 2935 3504 2936
rect 3495 2931 3496 2935
rect 3503 2931 3504 2935
rect 3495 2930 3504 2931
rect 2900 2924 2966 2926
rect 2900 2923 2901 2924
rect 2895 2922 2901 2923
rect 151 2919 160 2920
rect 151 2915 152 2919
rect 159 2915 160 2919
rect 151 2914 160 2915
rect 279 2919 285 2920
rect 279 2915 280 2919
rect 284 2918 285 2919
rect 303 2919 309 2920
rect 303 2918 304 2919
rect 284 2916 304 2918
rect 284 2915 285 2916
rect 279 2914 285 2915
rect 303 2915 304 2916
rect 308 2915 309 2919
rect 303 2914 309 2915
rect 471 2919 480 2920
rect 471 2915 472 2919
rect 479 2915 480 2919
rect 471 2914 480 2915
rect 583 2919 589 2920
rect 583 2915 584 2919
rect 588 2918 589 2919
rect 639 2919 645 2920
rect 639 2918 640 2919
rect 588 2916 640 2918
rect 588 2915 589 2916
rect 583 2914 589 2915
rect 639 2915 640 2916
rect 644 2915 645 2919
rect 639 2914 645 2915
rect 775 2919 781 2920
rect 775 2915 776 2919
rect 780 2918 781 2919
rect 799 2919 805 2920
rect 799 2918 800 2919
rect 780 2916 800 2918
rect 780 2915 781 2916
rect 775 2914 781 2915
rect 799 2915 800 2916
rect 804 2915 805 2919
rect 799 2914 805 2915
rect 943 2919 952 2920
rect 943 2915 944 2919
rect 951 2915 952 2919
rect 943 2914 952 2915
rect 1079 2919 1085 2920
rect 1079 2915 1080 2919
rect 1084 2918 1085 2919
rect 1118 2919 1124 2920
rect 1118 2918 1119 2919
rect 1084 2916 1119 2918
rect 1084 2915 1085 2916
rect 1079 2914 1085 2915
rect 1118 2915 1119 2916
rect 1123 2915 1124 2919
rect 1118 2914 1124 2915
rect 1183 2919 1189 2920
rect 1183 2915 1184 2919
rect 1188 2918 1189 2919
rect 1207 2919 1213 2920
rect 1207 2918 1208 2919
rect 1188 2916 1208 2918
rect 1188 2915 1189 2916
rect 1183 2914 1189 2915
rect 1207 2915 1208 2916
rect 1212 2915 1213 2919
rect 1207 2914 1213 2915
rect 1303 2919 1309 2920
rect 1303 2915 1304 2919
rect 1308 2918 1309 2919
rect 1327 2919 1333 2920
rect 1327 2918 1328 2919
rect 1308 2916 1328 2918
rect 1308 2915 1309 2916
rect 1303 2914 1309 2915
rect 1327 2915 1328 2916
rect 1332 2915 1333 2919
rect 1327 2914 1333 2915
rect 1439 2919 1445 2920
rect 1439 2915 1440 2919
rect 1444 2918 1445 2919
rect 1490 2919 1496 2920
rect 1490 2918 1491 2919
rect 1444 2916 1491 2918
rect 1444 2915 1445 2916
rect 1439 2914 1445 2915
rect 1490 2915 1491 2916
rect 1495 2915 1496 2919
rect 1490 2914 1496 2915
rect 1543 2919 1549 2920
rect 1543 2915 1544 2919
rect 1548 2918 1549 2919
rect 1594 2919 1600 2920
rect 1594 2918 1595 2919
rect 1548 2916 1595 2918
rect 1548 2915 1549 2916
rect 1543 2914 1549 2915
rect 1594 2915 1595 2916
rect 1599 2915 1600 2919
rect 1594 2914 1600 2915
rect 1655 2919 1661 2920
rect 1655 2915 1656 2919
rect 1660 2918 1661 2919
rect 1711 2919 1717 2920
rect 1711 2918 1712 2919
rect 1660 2916 1712 2918
rect 1660 2915 1661 2916
rect 1655 2914 1661 2915
rect 1711 2915 1712 2916
rect 1716 2915 1717 2919
rect 1711 2914 1717 2915
rect 1743 2919 1749 2920
rect 1743 2915 1744 2919
rect 1748 2918 1749 2919
rect 1870 2919 1876 2920
rect 1870 2918 1871 2919
rect 1748 2916 1871 2918
rect 1748 2915 1749 2916
rect 1743 2914 1749 2915
rect 1870 2915 1871 2916
rect 1875 2915 1876 2919
rect 1870 2914 1876 2915
rect 2903 2915 2909 2916
rect 2903 2911 2904 2915
rect 2908 2914 2909 2915
rect 3055 2915 3061 2916
rect 3055 2914 3056 2915
rect 2908 2912 3056 2914
rect 2908 2911 2909 2912
rect 2903 2910 2909 2911
rect 3055 2911 3056 2912
rect 3060 2911 3061 2915
rect 3055 2910 3061 2911
rect 3162 2915 3168 2916
rect 3162 2911 3163 2915
rect 3167 2914 3168 2915
rect 3207 2915 3213 2916
rect 3207 2914 3208 2915
rect 3167 2912 3208 2914
rect 3167 2911 3168 2912
rect 3162 2910 3168 2911
rect 3207 2911 3208 2912
rect 3212 2911 3213 2915
rect 3207 2910 3213 2911
rect 3471 2915 3477 2916
rect 3471 2911 3472 2915
rect 3476 2914 3477 2915
rect 3495 2915 3501 2916
rect 3495 2914 3496 2915
rect 3476 2912 3496 2914
rect 3476 2911 3477 2912
rect 3471 2910 3477 2911
rect 3495 2911 3496 2912
rect 3500 2911 3501 2915
rect 3495 2910 3501 2911
rect 151 2907 157 2908
rect 151 2903 152 2907
rect 156 2906 157 2907
rect 234 2907 240 2908
rect 234 2906 235 2907
rect 156 2904 235 2906
rect 156 2903 157 2904
rect 151 2902 157 2903
rect 234 2903 235 2904
rect 239 2903 240 2907
rect 234 2902 240 2903
rect 327 2907 333 2908
rect 327 2903 328 2907
rect 332 2906 333 2907
rect 354 2907 360 2908
rect 354 2906 355 2907
rect 332 2904 355 2906
rect 332 2903 333 2904
rect 327 2902 333 2903
rect 354 2903 355 2904
rect 359 2903 360 2907
rect 354 2902 360 2903
rect 527 2907 533 2908
rect 527 2903 528 2907
rect 532 2906 533 2907
rect 623 2907 629 2908
rect 623 2906 624 2907
rect 532 2904 624 2906
rect 532 2903 533 2904
rect 527 2902 533 2903
rect 623 2903 624 2904
rect 628 2903 629 2907
rect 623 2902 629 2903
rect 719 2907 725 2908
rect 719 2903 720 2907
rect 724 2906 725 2907
rect 778 2907 784 2908
rect 778 2906 779 2907
rect 724 2904 779 2906
rect 724 2903 725 2904
rect 719 2902 725 2903
rect 778 2903 779 2904
rect 783 2903 784 2907
rect 778 2902 784 2903
rect 902 2907 909 2908
rect 902 2903 903 2907
rect 908 2903 909 2907
rect 902 2902 909 2903
rect 1079 2907 1085 2908
rect 1079 2903 1080 2907
rect 1084 2906 1085 2907
rect 1118 2907 1124 2908
rect 1118 2906 1119 2907
rect 1084 2904 1119 2906
rect 1084 2903 1085 2904
rect 1079 2902 1085 2903
rect 1118 2903 1119 2904
rect 1123 2903 1124 2907
rect 1118 2902 1124 2903
rect 1162 2907 1168 2908
rect 1162 2903 1163 2907
rect 1167 2906 1168 2907
rect 1247 2907 1253 2908
rect 1247 2906 1248 2907
rect 1167 2904 1248 2906
rect 1167 2903 1168 2904
rect 1162 2902 1168 2903
rect 1247 2903 1248 2904
rect 1252 2903 1253 2907
rect 1247 2902 1253 2903
rect 1406 2907 1413 2908
rect 1406 2903 1407 2907
rect 1412 2903 1413 2907
rect 1406 2902 1413 2903
rect 1479 2907 1485 2908
rect 1479 2903 1480 2907
rect 1484 2906 1485 2907
rect 1559 2907 1565 2908
rect 1559 2906 1560 2907
rect 1484 2904 1560 2906
rect 1484 2903 1485 2904
rect 1479 2902 1485 2903
rect 1559 2903 1560 2904
rect 1564 2903 1565 2907
rect 1559 2902 1565 2903
rect 1639 2907 1645 2908
rect 1639 2903 1640 2907
rect 1644 2906 1645 2907
rect 1719 2907 1725 2908
rect 1719 2906 1720 2907
rect 1644 2904 1720 2906
rect 1644 2903 1645 2904
rect 1639 2902 1645 2903
rect 1719 2903 1720 2904
rect 1724 2903 1725 2907
rect 1719 2902 1725 2903
rect 2894 2905 2900 2906
rect 2894 2901 2895 2905
rect 2899 2901 2900 2905
rect 2894 2900 2900 2901
rect 3198 2905 3204 2906
rect 3198 2901 3199 2905
rect 3203 2901 3204 2905
rect 3198 2900 3204 2901
rect 3486 2905 3492 2906
rect 3486 2901 3487 2905
rect 3491 2901 3492 2905
rect 3486 2900 3492 2901
rect 142 2897 148 2898
rect 142 2893 143 2897
rect 147 2893 148 2897
rect 142 2892 148 2893
rect 318 2897 324 2898
rect 318 2893 319 2897
rect 323 2893 324 2897
rect 318 2892 324 2893
rect 518 2897 524 2898
rect 518 2893 519 2897
rect 523 2893 524 2897
rect 518 2892 524 2893
rect 710 2897 716 2898
rect 710 2893 711 2897
rect 715 2893 716 2897
rect 710 2892 716 2893
rect 894 2897 900 2898
rect 894 2893 895 2897
rect 899 2893 900 2897
rect 894 2892 900 2893
rect 1070 2897 1076 2898
rect 1070 2893 1071 2897
rect 1075 2893 1076 2897
rect 1070 2892 1076 2893
rect 1238 2897 1244 2898
rect 1238 2893 1239 2897
rect 1243 2893 1244 2897
rect 1238 2892 1244 2893
rect 1398 2897 1404 2898
rect 1398 2893 1399 2897
rect 1403 2893 1404 2897
rect 1398 2892 1404 2893
rect 1550 2897 1556 2898
rect 1550 2893 1551 2897
rect 1555 2893 1556 2897
rect 1550 2892 1556 2893
rect 1710 2897 1716 2898
rect 1710 2893 1711 2897
rect 1715 2893 1716 2897
rect 1710 2892 1716 2893
rect 1862 2892 1868 2893
rect 3574 2892 3580 2893
rect 1862 2888 1863 2892
rect 1867 2888 1868 2892
rect 2954 2891 2960 2892
rect 2954 2890 2955 2891
rect 2949 2888 2955 2890
rect 1862 2887 1868 2888
rect 2954 2887 2955 2888
rect 2959 2887 2960 2891
rect 3574 2888 3575 2892
rect 3579 2888 3580 2892
rect 2954 2886 2960 2887
rect 3055 2887 3061 2888
rect 3574 2887 3580 2888
rect 110 2884 116 2885
rect 1822 2884 1828 2885
rect 110 2880 111 2884
rect 115 2880 116 2884
rect 583 2883 589 2884
rect 583 2882 584 2883
rect 573 2880 584 2882
rect 110 2879 116 2880
rect 234 2879 240 2880
rect 234 2875 235 2879
rect 239 2878 240 2879
rect 583 2879 584 2880
rect 588 2879 589 2883
rect 1162 2883 1168 2884
rect 1162 2882 1163 2883
rect 1125 2880 1163 2882
rect 583 2878 589 2879
rect 623 2879 629 2880
rect 239 2876 337 2878
rect 239 2875 240 2876
rect 234 2874 240 2875
rect 623 2875 624 2879
rect 628 2878 629 2879
rect 778 2879 784 2880
rect 628 2876 729 2878
rect 628 2875 629 2876
rect 623 2874 629 2875
rect 778 2875 779 2879
rect 783 2878 784 2879
rect 1162 2879 1163 2880
rect 1167 2879 1168 2883
rect 1479 2883 1485 2884
rect 1479 2882 1480 2883
rect 1453 2880 1480 2882
rect 1162 2878 1168 2879
rect 1479 2879 1480 2880
rect 1484 2879 1485 2883
rect 1639 2883 1645 2884
rect 1639 2882 1640 2883
rect 1605 2880 1640 2882
rect 1479 2878 1485 2879
rect 1639 2879 1640 2880
rect 1644 2879 1645 2883
rect 1822 2880 1823 2884
rect 1827 2880 1828 2884
rect 3055 2883 3056 2887
rect 3060 2886 3061 2887
rect 3060 2884 3217 2886
rect 3060 2883 3061 2884
rect 3055 2882 3061 2883
rect 1639 2878 1645 2879
rect 1650 2879 1656 2880
rect 1822 2879 1828 2880
rect 783 2876 913 2878
rect 783 2875 784 2876
rect 778 2874 784 2875
rect 1650 2875 1651 2879
rect 1655 2878 1656 2879
rect 1655 2876 1729 2878
rect 1655 2875 1656 2876
rect 1650 2874 1656 2875
rect 1862 2875 1868 2876
rect 1862 2871 1863 2875
rect 1867 2871 1868 2875
rect 1862 2870 1868 2871
rect 3574 2875 3580 2876
rect 3574 2871 3575 2875
rect 3579 2871 3580 2875
rect 3574 2870 3580 2871
rect 110 2867 116 2868
rect 110 2863 111 2867
rect 115 2863 116 2867
rect 110 2862 116 2863
rect 1822 2867 1828 2868
rect 1822 2863 1823 2867
rect 1827 2863 1828 2867
rect 1822 2862 1828 2863
rect 2886 2865 2892 2866
rect 2886 2861 2887 2865
rect 2891 2861 2892 2865
rect 2886 2860 2892 2861
rect 3190 2865 3196 2866
rect 3190 2861 3191 2865
rect 3195 2861 3196 2865
rect 3190 2860 3196 2861
rect 3478 2865 3484 2866
rect 3478 2861 3479 2865
rect 3483 2861 3484 2865
rect 3478 2860 3484 2861
rect 3498 2859 3504 2860
rect 134 2857 140 2858
rect 134 2853 135 2857
rect 139 2853 140 2857
rect 134 2852 140 2853
rect 310 2857 316 2858
rect 310 2853 311 2857
rect 315 2853 316 2857
rect 310 2852 316 2853
rect 510 2857 516 2858
rect 510 2853 511 2857
rect 515 2853 516 2857
rect 510 2852 516 2853
rect 702 2857 708 2858
rect 702 2853 703 2857
rect 707 2853 708 2857
rect 702 2852 708 2853
rect 886 2857 892 2858
rect 886 2853 887 2857
rect 891 2853 892 2857
rect 886 2852 892 2853
rect 1062 2857 1068 2858
rect 1062 2853 1063 2857
rect 1067 2853 1068 2857
rect 1062 2852 1068 2853
rect 1230 2857 1236 2858
rect 1230 2853 1231 2857
rect 1235 2853 1236 2857
rect 1230 2852 1236 2853
rect 1390 2857 1396 2858
rect 1390 2853 1391 2857
rect 1395 2853 1396 2857
rect 1390 2852 1396 2853
rect 1542 2857 1548 2858
rect 1542 2853 1543 2857
rect 1547 2853 1548 2857
rect 1542 2852 1548 2853
rect 1702 2857 1708 2858
rect 1702 2853 1703 2857
rect 1707 2853 1708 2857
rect 3498 2855 3499 2859
rect 3503 2858 3504 2859
rect 3527 2859 3533 2860
rect 3527 2858 3528 2859
rect 3503 2856 3528 2858
rect 3503 2855 3504 2856
rect 3498 2854 3504 2855
rect 3527 2855 3528 2856
rect 3532 2855 3533 2859
rect 3527 2854 3533 2855
rect 1702 2852 1708 2853
rect 178 2851 189 2852
rect 178 2847 179 2851
rect 183 2847 184 2851
rect 188 2847 189 2851
rect 178 2846 189 2847
rect 1279 2851 1285 2852
rect 1279 2847 1280 2851
rect 1284 2850 1285 2851
rect 1290 2851 1296 2852
rect 1290 2850 1291 2851
rect 1284 2848 1291 2850
rect 1284 2847 1285 2848
rect 1279 2846 1285 2847
rect 1290 2847 1291 2848
rect 1295 2847 1296 2851
rect 1290 2846 1296 2847
rect 2830 2843 2836 2844
rect 2830 2839 2831 2843
rect 2835 2839 2836 2843
rect 2830 2838 2836 2839
rect 2918 2843 2924 2844
rect 2918 2839 2919 2843
rect 2923 2839 2924 2843
rect 2918 2838 2924 2839
rect 3006 2843 3012 2844
rect 3006 2839 3007 2843
rect 3011 2839 3012 2843
rect 3006 2838 3012 2839
rect 3094 2843 3100 2844
rect 3094 2839 3095 2843
rect 3099 2839 3100 2843
rect 3094 2838 3100 2839
rect 3162 2835 3168 2836
rect 3162 2834 3163 2835
rect 1862 2833 1868 2834
rect 158 2831 164 2832
rect 158 2827 159 2831
rect 163 2827 164 2831
rect 158 2826 164 2827
rect 318 2831 324 2832
rect 318 2827 319 2831
rect 323 2827 324 2831
rect 318 2826 324 2827
rect 486 2831 492 2832
rect 486 2827 487 2831
rect 491 2827 492 2831
rect 486 2826 492 2827
rect 654 2831 660 2832
rect 654 2827 655 2831
rect 659 2827 660 2831
rect 654 2826 660 2827
rect 822 2831 828 2832
rect 822 2827 823 2831
rect 827 2827 828 2831
rect 822 2826 828 2827
rect 974 2831 980 2832
rect 974 2827 975 2831
rect 979 2827 980 2831
rect 974 2826 980 2827
rect 1126 2831 1132 2832
rect 1126 2827 1127 2831
rect 1131 2827 1132 2831
rect 1126 2826 1132 2827
rect 1270 2831 1276 2832
rect 1270 2827 1271 2831
rect 1275 2827 1276 2831
rect 1270 2826 1276 2827
rect 1414 2831 1420 2832
rect 1414 2827 1415 2831
rect 1419 2827 1420 2831
rect 1414 2826 1420 2827
rect 1558 2831 1564 2832
rect 1558 2827 1559 2831
rect 1563 2827 1564 2831
rect 1862 2829 1863 2833
rect 1867 2829 1868 2833
rect 3153 2832 3163 2834
rect 3162 2831 3163 2832
rect 3167 2831 3168 2835
rect 3162 2830 3168 2831
rect 3574 2833 3580 2834
rect 1862 2828 1868 2829
rect 3574 2829 3575 2833
rect 3579 2829 3580 2833
rect 3574 2828 3580 2829
rect 1558 2826 1564 2827
rect 902 2823 908 2824
rect 902 2822 903 2823
rect 110 2821 116 2822
rect 110 2817 111 2821
rect 115 2817 116 2821
rect 881 2820 903 2822
rect 902 2819 903 2820
rect 907 2819 908 2823
rect 902 2818 908 2819
rect 1482 2823 1488 2824
rect 1482 2819 1483 2823
rect 1487 2822 1488 2823
rect 1487 2820 1577 2822
rect 1822 2821 1828 2822
rect 1487 2819 1488 2820
rect 1482 2818 1488 2819
rect 110 2816 116 2817
rect 1822 2817 1823 2821
rect 1827 2817 1828 2821
rect 2898 2819 2904 2820
rect 2898 2818 2899 2819
rect 1822 2816 1828 2817
rect 1862 2816 1868 2817
rect 2893 2816 2899 2818
rect 1862 2812 1863 2816
rect 1867 2812 1868 2816
rect 2898 2815 2899 2816
rect 2903 2815 2904 2819
rect 2986 2819 2992 2820
rect 2986 2818 2987 2819
rect 2981 2816 2987 2818
rect 2898 2814 2904 2815
rect 2986 2815 2987 2816
rect 2991 2815 2992 2819
rect 3074 2819 3080 2820
rect 3074 2818 3075 2819
rect 3069 2816 3075 2818
rect 2986 2814 2992 2815
rect 3074 2815 3075 2816
rect 3079 2815 3080 2819
rect 3074 2814 3080 2815
rect 3574 2816 3580 2817
rect 1862 2811 1868 2812
rect 3574 2812 3575 2816
rect 3579 2812 3580 2816
rect 3574 2811 3580 2812
rect 250 2807 256 2808
rect 250 2806 251 2807
rect 110 2804 116 2805
rect 221 2804 251 2806
rect 110 2800 111 2804
rect 115 2800 116 2804
rect 250 2803 251 2804
rect 255 2803 256 2807
rect 386 2807 392 2808
rect 386 2806 387 2807
rect 381 2804 387 2806
rect 250 2802 256 2803
rect 386 2803 387 2804
rect 391 2803 392 2807
rect 647 2807 653 2808
rect 647 2806 648 2807
rect 549 2804 648 2806
rect 386 2802 392 2803
rect 647 2803 648 2804
rect 652 2803 653 2807
rect 815 2807 821 2808
rect 815 2806 816 2807
rect 717 2804 816 2806
rect 647 2802 653 2803
rect 815 2803 816 2804
rect 820 2803 821 2807
rect 1119 2807 1125 2808
rect 1119 2806 1120 2807
rect 1037 2804 1120 2806
rect 815 2802 821 2803
rect 1119 2803 1120 2804
rect 1124 2803 1125 2807
rect 1263 2807 1269 2808
rect 1263 2806 1264 2807
rect 1189 2804 1264 2806
rect 1119 2802 1125 2803
rect 1263 2803 1264 2804
rect 1268 2803 1269 2807
rect 1407 2807 1413 2808
rect 1407 2806 1408 2807
rect 1333 2804 1408 2806
rect 1263 2802 1269 2803
rect 1407 2803 1408 2804
rect 1412 2803 1413 2807
rect 1551 2807 1557 2808
rect 1551 2806 1552 2807
rect 1477 2804 1552 2806
rect 1407 2802 1413 2803
rect 1551 2803 1552 2804
rect 1556 2803 1557 2807
rect 1551 2802 1557 2803
rect 1822 2804 1828 2805
rect 110 2799 116 2800
rect 1822 2800 1823 2804
rect 1827 2800 1828 2804
rect 1822 2799 1828 2800
rect 2838 2803 2844 2804
rect 2838 2799 2839 2803
rect 2843 2799 2844 2803
rect 2838 2798 2844 2799
rect 2926 2803 2932 2804
rect 2926 2799 2927 2803
rect 2931 2799 2932 2803
rect 2926 2798 2932 2799
rect 3014 2803 3020 2804
rect 3014 2799 3015 2803
rect 3019 2799 3020 2803
rect 3014 2798 3020 2799
rect 3102 2803 3108 2804
rect 3102 2799 3103 2803
rect 3107 2799 3108 2803
rect 3102 2798 3108 2799
rect 166 2791 172 2792
rect 166 2787 167 2791
rect 171 2787 172 2791
rect 166 2786 172 2787
rect 326 2791 332 2792
rect 326 2787 327 2791
rect 331 2787 332 2791
rect 326 2786 332 2787
rect 494 2791 500 2792
rect 494 2787 495 2791
rect 499 2787 500 2791
rect 494 2786 500 2787
rect 662 2791 668 2792
rect 662 2787 663 2791
rect 667 2787 668 2791
rect 662 2786 668 2787
rect 830 2791 836 2792
rect 830 2787 831 2791
rect 835 2787 836 2791
rect 830 2786 836 2787
rect 982 2791 988 2792
rect 982 2787 983 2791
rect 987 2787 988 2791
rect 982 2786 988 2787
rect 1134 2791 1140 2792
rect 1134 2787 1135 2791
rect 1139 2787 1140 2791
rect 1134 2786 1140 2787
rect 1278 2791 1284 2792
rect 1278 2787 1279 2791
rect 1283 2787 1284 2791
rect 1278 2786 1284 2787
rect 1422 2791 1428 2792
rect 1422 2787 1423 2791
rect 1427 2787 1428 2791
rect 1422 2786 1428 2787
rect 1566 2791 1572 2792
rect 1566 2787 1567 2791
rect 1571 2787 1572 2791
rect 1566 2786 1572 2787
rect 2847 2791 2856 2792
rect 2847 2787 2848 2791
rect 2855 2787 2856 2791
rect 2847 2786 2856 2787
rect 2898 2791 2904 2792
rect 2898 2787 2899 2791
rect 2903 2790 2904 2791
rect 2935 2791 2941 2792
rect 2935 2790 2936 2791
rect 2903 2788 2936 2790
rect 2903 2787 2904 2788
rect 2898 2786 2904 2787
rect 2935 2787 2936 2788
rect 2940 2787 2941 2791
rect 2935 2786 2941 2787
rect 2986 2791 2992 2792
rect 2986 2787 2987 2791
rect 2991 2790 2992 2791
rect 3023 2791 3029 2792
rect 3023 2790 3024 2791
rect 2991 2788 3024 2790
rect 2991 2787 2992 2788
rect 2986 2786 2992 2787
rect 3023 2787 3024 2788
rect 3028 2787 3029 2791
rect 3023 2786 3029 2787
rect 3074 2791 3080 2792
rect 3074 2787 3075 2791
rect 3079 2790 3080 2791
rect 3111 2791 3117 2792
rect 3111 2790 3112 2791
rect 3079 2788 3112 2790
rect 3079 2787 3080 2788
rect 3074 2786 3080 2787
rect 3111 2787 3112 2788
rect 3116 2787 3117 2791
rect 3111 2786 3117 2787
rect 175 2779 184 2780
rect 175 2775 176 2779
rect 183 2775 184 2779
rect 175 2774 184 2775
rect 250 2779 256 2780
rect 250 2775 251 2779
rect 255 2778 256 2779
rect 335 2779 341 2780
rect 335 2778 336 2779
rect 255 2776 336 2778
rect 255 2775 256 2776
rect 250 2774 256 2775
rect 335 2775 336 2776
rect 340 2775 341 2779
rect 335 2774 341 2775
rect 503 2779 509 2780
rect 503 2775 504 2779
rect 508 2778 509 2779
rect 530 2779 536 2780
rect 530 2778 531 2779
rect 508 2776 531 2778
rect 508 2775 509 2776
rect 503 2774 509 2775
rect 530 2775 531 2776
rect 535 2775 536 2779
rect 530 2774 536 2775
rect 647 2779 653 2780
rect 647 2775 648 2779
rect 652 2778 653 2779
rect 671 2779 677 2780
rect 671 2778 672 2779
rect 652 2776 672 2778
rect 652 2775 653 2776
rect 647 2774 653 2775
rect 671 2775 672 2776
rect 676 2775 677 2779
rect 671 2774 677 2775
rect 815 2779 821 2780
rect 815 2775 816 2779
rect 820 2778 821 2779
rect 839 2779 845 2780
rect 839 2778 840 2779
rect 820 2776 840 2778
rect 820 2775 821 2776
rect 815 2774 821 2775
rect 839 2775 840 2776
rect 844 2775 845 2779
rect 839 2774 845 2775
rect 991 2779 1000 2780
rect 991 2775 992 2779
rect 999 2775 1000 2779
rect 991 2774 1000 2775
rect 1119 2779 1125 2780
rect 1119 2775 1120 2779
rect 1124 2778 1125 2779
rect 1143 2779 1149 2780
rect 1143 2778 1144 2779
rect 1124 2776 1144 2778
rect 1124 2775 1125 2776
rect 1119 2774 1125 2775
rect 1143 2775 1144 2776
rect 1148 2775 1149 2779
rect 1143 2774 1149 2775
rect 1287 2779 1296 2780
rect 1287 2775 1288 2779
rect 1295 2775 1296 2779
rect 1287 2774 1296 2775
rect 1407 2779 1413 2780
rect 1407 2775 1408 2779
rect 1412 2778 1413 2779
rect 1431 2779 1437 2780
rect 1431 2778 1432 2779
rect 1412 2776 1432 2778
rect 1412 2775 1413 2776
rect 1407 2774 1413 2775
rect 1431 2775 1432 2776
rect 1436 2775 1437 2779
rect 1431 2774 1437 2775
rect 1551 2779 1557 2780
rect 1551 2775 1552 2779
rect 1556 2778 1557 2779
rect 1575 2779 1581 2780
rect 1575 2778 1576 2779
rect 1556 2776 1576 2778
rect 1556 2775 1557 2776
rect 1551 2774 1557 2775
rect 1575 2775 1576 2776
rect 1580 2775 1581 2779
rect 1575 2774 1581 2775
rect 2679 2779 2685 2780
rect 2679 2775 2680 2779
rect 2684 2778 2685 2779
rect 2734 2779 2740 2780
rect 2734 2778 2735 2779
rect 2684 2776 2735 2778
rect 2684 2775 2685 2776
rect 2679 2774 2685 2775
rect 2734 2775 2735 2776
rect 2739 2775 2740 2779
rect 2734 2774 2740 2775
rect 2743 2779 2749 2780
rect 2743 2775 2744 2779
rect 2748 2778 2749 2779
rect 2815 2779 2821 2780
rect 2815 2778 2816 2779
rect 2748 2776 2816 2778
rect 2748 2775 2749 2776
rect 2743 2774 2749 2775
rect 2815 2775 2816 2776
rect 2820 2775 2821 2779
rect 2815 2774 2821 2775
rect 2951 2779 2957 2780
rect 2951 2775 2952 2779
rect 2956 2778 2957 2779
rect 2975 2779 2981 2780
rect 2975 2778 2976 2779
rect 2956 2776 2976 2778
rect 2956 2775 2957 2776
rect 2951 2774 2957 2775
rect 2975 2775 2976 2776
rect 2980 2775 2981 2779
rect 2975 2774 2981 2775
rect 3063 2779 3069 2780
rect 3063 2775 3064 2779
rect 3068 2778 3069 2779
rect 3151 2779 3157 2780
rect 3151 2778 3152 2779
rect 3068 2776 3152 2778
rect 3068 2775 3069 2776
rect 3063 2774 3069 2775
rect 3151 2775 3152 2776
rect 3156 2775 3157 2779
rect 3151 2774 3157 2775
rect 3239 2779 3245 2780
rect 3239 2775 3240 2779
rect 3244 2778 3245 2779
rect 3335 2779 3341 2780
rect 3335 2778 3336 2779
rect 3244 2776 3336 2778
rect 3244 2775 3245 2776
rect 3239 2774 3245 2775
rect 3335 2775 3336 2776
rect 3340 2775 3341 2779
rect 3335 2774 3341 2775
rect 3495 2779 3504 2780
rect 3495 2775 3496 2779
rect 3503 2775 3504 2779
rect 3495 2774 3504 2775
rect 2670 2769 2676 2770
rect 695 2767 701 2768
rect 695 2766 696 2767
rect 608 2764 696 2766
rect 215 2759 221 2760
rect 215 2755 216 2759
rect 220 2758 221 2759
rect 302 2759 308 2760
rect 302 2758 303 2759
rect 220 2756 303 2758
rect 220 2755 221 2756
rect 215 2754 221 2755
rect 302 2755 303 2756
rect 307 2755 308 2759
rect 302 2754 308 2755
rect 343 2759 349 2760
rect 343 2755 344 2759
rect 348 2758 349 2759
rect 386 2759 392 2760
rect 386 2758 387 2759
rect 348 2756 387 2758
rect 348 2755 349 2756
rect 343 2754 349 2755
rect 386 2755 387 2756
rect 391 2755 392 2759
rect 386 2754 392 2755
rect 479 2759 485 2760
rect 479 2755 480 2759
rect 484 2758 485 2759
rect 608 2758 610 2764
rect 695 2763 696 2764
rect 700 2763 701 2767
rect 1367 2767 1373 2768
rect 1367 2766 1368 2767
rect 695 2762 701 2763
rect 1024 2764 1368 2766
rect 484 2756 610 2758
rect 615 2759 621 2760
rect 484 2755 485 2756
rect 479 2754 485 2755
rect 615 2755 616 2759
rect 620 2758 621 2759
rect 650 2759 656 2760
rect 650 2758 651 2759
rect 620 2756 651 2758
rect 620 2755 621 2756
rect 615 2754 621 2755
rect 650 2755 651 2756
rect 655 2755 656 2759
rect 650 2754 656 2755
rect 687 2759 693 2760
rect 687 2755 688 2759
rect 692 2758 693 2759
rect 759 2759 765 2760
rect 759 2758 760 2759
rect 692 2756 760 2758
rect 692 2755 693 2756
rect 687 2754 693 2755
rect 759 2755 760 2756
rect 764 2755 765 2759
rect 759 2754 765 2755
rect 895 2759 901 2760
rect 895 2755 896 2759
rect 900 2758 901 2759
rect 1024 2758 1026 2764
rect 1367 2763 1368 2764
rect 1372 2763 1373 2767
rect 2670 2765 2671 2769
rect 2675 2765 2676 2769
rect 2670 2764 2676 2765
rect 2806 2769 2812 2770
rect 2806 2765 2807 2769
rect 2811 2765 2812 2769
rect 2806 2764 2812 2765
rect 2966 2769 2972 2770
rect 2966 2765 2967 2769
rect 2971 2765 2972 2769
rect 2966 2764 2972 2765
rect 3142 2769 3148 2770
rect 3142 2765 3143 2769
rect 3147 2765 3148 2769
rect 3142 2764 3148 2765
rect 3326 2769 3332 2770
rect 3326 2765 3327 2769
rect 3331 2765 3332 2769
rect 3326 2764 3332 2765
rect 3486 2769 3492 2770
rect 3486 2765 3487 2769
rect 3491 2765 3492 2769
rect 3486 2764 3492 2765
rect 1367 2762 1373 2763
rect 900 2756 1026 2758
rect 1031 2759 1037 2760
rect 900 2755 901 2756
rect 895 2754 901 2755
rect 1031 2755 1032 2759
rect 1036 2755 1037 2759
rect 1031 2754 1037 2755
rect 1095 2759 1101 2760
rect 1095 2755 1096 2759
rect 1100 2758 1101 2759
rect 1159 2759 1165 2760
rect 1159 2758 1160 2759
rect 1100 2756 1160 2758
rect 1100 2755 1101 2756
rect 1095 2754 1101 2755
rect 1159 2755 1160 2756
rect 1164 2755 1165 2759
rect 1159 2754 1165 2755
rect 1263 2759 1269 2760
rect 1263 2755 1264 2759
rect 1268 2758 1269 2759
rect 1295 2759 1301 2760
rect 1295 2758 1296 2759
rect 1268 2756 1296 2758
rect 1268 2755 1269 2756
rect 1263 2754 1269 2755
rect 1295 2755 1296 2756
rect 1300 2755 1301 2759
rect 1295 2754 1301 2755
rect 1359 2759 1365 2760
rect 1359 2755 1360 2759
rect 1364 2758 1365 2759
rect 1431 2759 1437 2760
rect 1431 2758 1432 2759
rect 1364 2756 1432 2758
rect 1364 2755 1365 2756
rect 1359 2754 1365 2755
rect 1431 2755 1432 2756
rect 1436 2755 1437 2759
rect 1431 2754 1437 2755
rect 1862 2756 1868 2757
rect 3574 2756 3580 2757
rect 940 2752 1034 2754
rect 1862 2752 1863 2756
rect 1867 2752 1868 2756
rect 2743 2755 2749 2756
rect 2743 2754 2744 2755
rect 2725 2752 2744 2754
rect 206 2749 212 2750
rect 206 2745 207 2749
rect 211 2745 212 2749
rect 206 2744 212 2745
rect 334 2749 340 2750
rect 334 2745 335 2749
rect 339 2745 340 2749
rect 334 2744 340 2745
rect 470 2749 476 2750
rect 470 2745 471 2749
rect 475 2745 476 2749
rect 470 2744 476 2745
rect 606 2749 612 2750
rect 606 2745 607 2749
rect 611 2745 612 2749
rect 606 2744 612 2745
rect 750 2749 756 2750
rect 750 2745 751 2749
rect 755 2745 756 2749
rect 750 2744 756 2745
rect 886 2749 892 2750
rect 886 2745 887 2749
rect 891 2745 892 2749
rect 886 2744 892 2745
rect 110 2736 116 2737
rect 110 2732 111 2736
rect 115 2732 116 2736
rect 530 2735 536 2736
rect 530 2734 531 2735
rect 525 2732 531 2734
rect 110 2731 116 2732
rect 302 2731 308 2732
rect 302 2727 303 2731
rect 307 2730 308 2731
rect 530 2731 531 2732
rect 535 2731 536 2735
rect 687 2735 693 2736
rect 687 2734 688 2735
rect 661 2732 688 2734
rect 530 2730 536 2731
rect 687 2731 688 2732
rect 692 2731 693 2735
rect 940 2733 942 2752
rect 1862 2751 1868 2752
rect 2743 2751 2744 2752
rect 2748 2751 2749 2755
rect 2951 2755 2957 2756
rect 2951 2754 2952 2755
rect 2861 2752 2952 2754
rect 2743 2750 2749 2751
rect 2951 2751 2952 2752
rect 2956 2751 2957 2755
rect 3063 2755 3069 2756
rect 3063 2754 3064 2755
rect 3021 2752 3064 2754
rect 2951 2750 2957 2751
rect 3063 2751 3064 2752
rect 3068 2751 3069 2755
rect 3239 2755 3245 2756
rect 3239 2754 3240 2755
rect 3197 2752 3240 2754
rect 3063 2750 3069 2751
rect 3239 2751 3240 2752
rect 3244 2751 3245 2755
rect 3574 2752 3575 2756
rect 3579 2752 3580 2756
rect 3239 2750 3245 2751
rect 3258 2751 3264 2752
rect 3574 2751 3580 2752
rect 1022 2749 1028 2750
rect 1022 2745 1023 2749
rect 1027 2745 1028 2749
rect 1022 2744 1028 2745
rect 1150 2749 1156 2750
rect 1150 2745 1151 2749
rect 1155 2745 1156 2749
rect 1150 2744 1156 2745
rect 1286 2749 1292 2750
rect 1286 2745 1287 2749
rect 1291 2745 1292 2749
rect 1286 2744 1292 2745
rect 1422 2749 1428 2750
rect 1422 2745 1423 2749
rect 1427 2745 1428 2749
rect 3258 2747 3259 2751
rect 3263 2750 3264 2751
rect 3263 2748 3345 2750
rect 3263 2747 3264 2748
rect 3258 2746 3264 2747
rect 1422 2744 1428 2745
rect 1862 2739 1868 2740
rect 1822 2736 1828 2737
rect 1095 2735 1101 2736
rect 1095 2734 1096 2735
rect 1077 2732 1096 2734
rect 687 2730 693 2731
rect 695 2731 701 2732
rect 307 2728 353 2730
rect 307 2727 308 2728
rect 302 2726 308 2727
rect 695 2727 696 2731
rect 700 2730 701 2731
rect 1095 2731 1096 2732
rect 1100 2731 1101 2735
rect 1359 2735 1365 2736
rect 1359 2734 1360 2735
rect 1341 2732 1360 2734
rect 1095 2730 1101 2731
rect 1359 2731 1360 2732
rect 1364 2731 1365 2735
rect 1822 2732 1823 2736
rect 1827 2732 1828 2736
rect 1862 2735 1863 2739
rect 1867 2735 1868 2739
rect 1862 2734 1868 2735
rect 3574 2739 3580 2740
rect 3574 2735 3575 2739
rect 3579 2735 3580 2739
rect 3574 2734 3580 2735
rect 1359 2730 1365 2731
rect 1367 2731 1373 2732
rect 1822 2731 1828 2732
rect 700 2728 769 2730
rect 700 2727 701 2728
rect 695 2726 701 2727
rect 1367 2727 1368 2731
rect 1372 2730 1373 2731
rect 1372 2728 1441 2730
rect 2662 2729 2668 2730
rect 1372 2727 1373 2728
rect 1367 2726 1373 2727
rect 2662 2725 2663 2729
rect 2667 2725 2668 2729
rect 2662 2724 2668 2725
rect 2798 2729 2804 2730
rect 2798 2725 2799 2729
rect 2803 2725 2804 2729
rect 2798 2724 2804 2725
rect 2958 2729 2964 2730
rect 2958 2725 2959 2729
rect 2963 2725 2964 2729
rect 2958 2724 2964 2725
rect 3134 2729 3140 2730
rect 3134 2725 3135 2729
rect 3139 2725 3140 2729
rect 3134 2724 3140 2725
rect 3318 2729 3324 2730
rect 3318 2725 3319 2729
rect 3323 2725 3324 2729
rect 3318 2724 3324 2725
rect 3478 2729 3484 2730
rect 3478 2725 3479 2729
rect 3483 2725 3484 2729
rect 3478 2724 3484 2725
rect 3498 2723 3504 2724
rect 110 2719 116 2720
rect 110 2715 111 2719
rect 115 2715 116 2719
rect 110 2714 116 2715
rect 1822 2719 1828 2720
rect 1822 2715 1823 2719
rect 1827 2715 1828 2719
rect 3498 2719 3499 2723
rect 3503 2722 3504 2723
rect 3527 2723 3533 2724
rect 3527 2722 3528 2723
rect 3503 2720 3528 2722
rect 3503 2719 3504 2720
rect 3498 2718 3504 2719
rect 3527 2719 3528 2720
rect 3532 2719 3533 2723
rect 3527 2718 3533 2719
rect 1822 2714 1828 2715
rect 198 2709 204 2710
rect 198 2705 199 2709
rect 203 2705 204 2709
rect 198 2704 204 2705
rect 326 2709 332 2710
rect 326 2705 327 2709
rect 331 2705 332 2709
rect 326 2704 332 2705
rect 462 2709 468 2710
rect 462 2705 463 2709
rect 467 2705 468 2709
rect 462 2704 468 2705
rect 598 2709 604 2710
rect 598 2705 599 2709
rect 603 2705 604 2709
rect 598 2704 604 2705
rect 742 2709 748 2710
rect 742 2705 743 2709
rect 747 2705 748 2709
rect 742 2704 748 2705
rect 878 2709 884 2710
rect 878 2705 879 2709
rect 883 2705 884 2709
rect 878 2704 884 2705
rect 1014 2709 1020 2710
rect 1014 2705 1015 2709
rect 1019 2705 1020 2709
rect 1014 2704 1020 2705
rect 1142 2709 1148 2710
rect 1142 2705 1143 2709
rect 1147 2705 1148 2709
rect 1142 2704 1148 2705
rect 1278 2709 1284 2710
rect 1278 2705 1279 2709
rect 1283 2705 1284 2709
rect 1278 2704 1284 2705
rect 1414 2709 1420 2710
rect 1414 2705 1415 2709
rect 1419 2705 1420 2709
rect 1414 2704 1420 2705
rect 1886 2707 1892 2708
rect 234 2703 240 2704
rect 234 2699 235 2703
rect 239 2702 240 2703
rect 247 2703 253 2704
rect 247 2702 248 2703
rect 239 2700 248 2702
rect 239 2699 240 2700
rect 234 2698 240 2699
rect 247 2699 248 2700
rect 252 2699 253 2703
rect 247 2698 253 2699
rect 1178 2703 1184 2704
rect 1178 2699 1179 2703
rect 1183 2702 1184 2703
rect 1191 2703 1197 2704
rect 1191 2702 1192 2703
rect 1183 2700 1192 2702
rect 1183 2699 1184 2700
rect 1178 2698 1184 2699
rect 1191 2699 1192 2700
rect 1196 2699 1197 2703
rect 1886 2703 1887 2707
rect 1891 2703 1892 2707
rect 1886 2702 1892 2703
rect 1974 2707 1980 2708
rect 1974 2703 1975 2707
rect 1979 2703 1980 2707
rect 1974 2702 1980 2703
rect 2062 2707 2068 2708
rect 2062 2703 2063 2707
rect 2067 2703 2068 2707
rect 2062 2702 2068 2703
rect 2150 2707 2156 2708
rect 2150 2703 2151 2707
rect 2155 2703 2156 2707
rect 2150 2702 2156 2703
rect 2238 2707 2244 2708
rect 2238 2703 2239 2707
rect 2243 2703 2244 2707
rect 2238 2702 2244 2703
rect 2326 2707 2332 2708
rect 2326 2703 2327 2707
rect 2331 2703 2332 2707
rect 2326 2702 2332 2703
rect 2414 2707 2420 2708
rect 2414 2703 2415 2707
rect 2419 2703 2420 2707
rect 2414 2702 2420 2703
rect 2502 2707 2508 2708
rect 2502 2703 2503 2707
rect 2507 2703 2508 2707
rect 2502 2702 2508 2703
rect 2590 2707 2596 2708
rect 2590 2703 2591 2707
rect 2595 2703 2596 2707
rect 2590 2702 2596 2703
rect 2678 2707 2684 2708
rect 2678 2703 2679 2707
rect 2683 2703 2684 2707
rect 2678 2702 2684 2703
rect 2766 2707 2772 2708
rect 2766 2703 2767 2707
rect 2771 2703 2772 2707
rect 2766 2702 2772 2703
rect 2854 2707 2860 2708
rect 2854 2703 2855 2707
rect 2859 2703 2860 2707
rect 2854 2702 2860 2703
rect 2942 2707 2948 2708
rect 2942 2703 2943 2707
rect 2947 2703 2948 2707
rect 2942 2702 2948 2703
rect 3030 2707 3036 2708
rect 3030 2703 3031 2707
rect 3035 2703 3036 2707
rect 3030 2702 3036 2703
rect 3118 2707 3124 2708
rect 3118 2703 3119 2707
rect 3123 2703 3124 2707
rect 3118 2702 3124 2703
rect 3206 2707 3212 2708
rect 3206 2703 3207 2707
rect 3211 2703 3212 2707
rect 3206 2702 3212 2703
rect 3294 2707 3300 2708
rect 3294 2703 3295 2707
rect 3299 2703 3300 2707
rect 3294 2702 3300 2703
rect 3390 2707 3396 2708
rect 3390 2703 3391 2707
rect 3395 2703 3396 2707
rect 3390 2702 3396 2703
rect 3478 2707 3484 2708
rect 3478 2703 3479 2707
rect 3483 2703 3484 2707
rect 3478 2702 3484 2703
rect 1191 2698 1197 2699
rect 3362 2699 3368 2700
rect 1862 2697 1868 2698
rect 1862 2693 1863 2697
rect 1867 2693 1868 2697
rect 3362 2695 3363 2699
rect 3367 2698 3368 2699
rect 3367 2696 3409 2698
rect 3574 2697 3580 2698
rect 3367 2695 3368 2696
rect 3362 2694 3368 2695
rect 1862 2692 1868 2693
rect 3574 2693 3575 2697
rect 3579 2693 3580 2697
rect 3574 2692 3580 2693
rect 214 2683 220 2684
rect 214 2679 215 2683
rect 219 2679 220 2683
rect 214 2678 220 2679
rect 334 2683 340 2684
rect 334 2679 335 2683
rect 339 2679 340 2683
rect 334 2678 340 2679
rect 462 2683 468 2684
rect 462 2679 463 2683
rect 467 2679 468 2683
rect 462 2678 468 2679
rect 582 2683 588 2684
rect 582 2679 583 2683
rect 587 2679 588 2683
rect 582 2678 588 2679
rect 702 2683 708 2684
rect 702 2679 703 2683
rect 707 2679 708 2683
rect 702 2678 708 2679
rect 822 2683 828 2684
rect 822 2679 823 2683
rect 827 2679 828 2683
rect 822 2678 828 2679
rect 934 2683 940 2684
rect 934 2679 935 2683
rect 939 2679 940 2683
rect 934 2678 940 2679
rect 1046 2683 1052 2684
rect 1046 2679 1047 2683
rect 1051 2679 1052 2683
rect 1046 2678 1052 2679
rect 1158 2683 1164 2684
rect 1158 2679 1159 2683
rect 1163 2679 1164 2683
rect 1158 2678 1164 2679
rect 1270 2683 1276 2684
rect 1270 2679 1271 2683
rect 1275 2679 1276 2683
rect 1967 2683 1973 2684
rect 1967 2682 1968 2683
rect 1270 2678 1276 2679
rect 1862 2680 1868 2681
rect 1949 2680 1968 2682
rect 1862 2676 1863 2680
rect 1867 2676 1868 2680
rect 1967 2679 1968 2680
rect 1972 2679 1973 2683
rect 2042 2683 2048 2684
rect 2042 2682 2043 2683
rect 2037 2680 2043 2682
rect 1967 2678 1973 2679
rect 2042 2679 2043 2680
rect 2047 2679 2048 2683
rect 2143 2683 2149 2684
rect 2143 2682 2144 2683
rect 2125 2680 2144 2682
rect 2042 2678 2048 2679
rect 2143 2679 2144 2680
rect 2148 2679 2149 2683
rect 2231 2683 2237 2684
rect 2231 2682 2232 2683
rect 2213 2680 2232 2682
rect 2143 2678 2149 2679
rect 2231 2679 2232 2680
rect 2236 2679 2237 2683
rect 2319 2683 2325 2684
rect 2319 2682 2320 2683
rect 2301 2680 2320 2682
rect 2231 2678 2237 2679
rect 2319 2679 2320 2680
rect 2324 2679 2325 2683
rect 2407 2683 2413 2684
rect 2407 2682 2408 2683
rect 2389 2680 2408 2682
rect 2319 2678 2325 2679
rect 2407 2679 2408 2680
rect 2412 2679 2413 2683
rect 2495 2683 2501 2684
rect 2495 2682 2496 2683
rect 2477 2680 2496 2682
rect 2407 2678 2413 2679
rect 2495 2679 2496 2680
rect 2500 2679 2501 2683
rect 2583 2683 2589 2684
rect 2583 2682 2584 2683
rect 2565 2680 2584 2682
rect 2495 2678 2501 2679
rect 2583 2679 2584 2680
rect 2588 2679 2589 2683
rect 2671 2683 2677 2684
rect 2671 2682 2672 2683
rect 2653 2680 2672 2682
rect 2583 2678 2589 2679
rect 2671 2679 2672 2680
rect 2676 2679 2677 2683
rect 2759 2683 2765 2684
rect 2759 2682 2760 2683
rect 2741 2680 2760 2682
rect 2671 2678 2677 2679
rect 2759 2679 2760 2680
rect 2764 2679 2765 2683
rect 2847 2683 2853 2684
rect 2847 2682 2848 2683
rect 2829 2680 2848 2682
rect 2759 2678 2765 2679
rect 2847 2679 2848 2680
rect 2852 2679 2853 2683
rect 2935 2683 2941 2684
rect 2935 2682 2936 2683
rect 2917 2680 2936 2682
rect 2847 2678 2853 2679
rect 2935 2679 2936 2680
rect 2940 2679 2941 2683
rect 3023 2683 3029 2684
rect 3023 2682 3024 2683
rect 3005 2680 3024 2682
rect 2935 2678 2941 2679
rect 3023 2679 3024 2680
rect 3028 2679 3029 2683
rect 3111 2683 3117 2684
rect 3111 2682 3112 2683
rect 3093 2680 3112 2682
rect 3023 2678 3029 2679
rect 3111 2679 3112 2680
rect 3116 2679 3117 2683
rect 3199 2683 3205 2684
rect 3199 2682 3200 2683
rect 3181 2680 3200 2682
rect 3111 2678 3117 2679
rect 3199 2679 3200 2680
rect 3204 2679 3205 2683
rect 3287 2683 3293 2684
rect 3287 2682 3288 2683
rect 3269 2680 3288 2682
rect 3199 2678 3205 2679
rect 3287 2679 3288 2680
rect 3292 2679 3293 2683
rect 3383 2683 3389 2684
rect 3383 2682 3384 2683
rect 3357 2680 3384 2682
rect 3287 2678 3293 2679
rect 3383 2679 3384 2680
rect 3388 2679 3389 2683
rect 3383 2678 3389 2679
rect 3470 2683 3476 2684
rect 3470 2679 3471 2683
rect 3475 2682 3476 2683
rect 3475 2680 3505 2682
rect 3574 2680 3580 2681
rect 3475 2679 3476 2680
rect 3470 2678 3476 2679
rect 650 2675 656 2676
rect 650 2674 651 2675
rect 110 2673 116 2674
rect 110 2669 111 2673
rect 115 2669 116 2673
rect 641 2672 651 2674
rect 650 2671 651 2672
rect 655 2671 656 2675
rect 650 2670 656 2671
rect 1226 2675 1232 2676
rect 1862 2675 1868 2676
rect 3574 2676 3575 2680
rect 3579 2676 3580 2680
rect 3574 2675 3580 2676
rect 1226 2671 1227 2675
rect 1231 2674 1232 2675
rect 1231 2672 1289 2674
rect 1822 2673 1828 2674
rect 1231 2671 1232 2672
rect 1226 2670 1232 2671
rect 110 2668 116 2669
rect 1822 2669 1823 2673
rect 1827 2669 1828 2673
rect 1822 2668 1828 2669
rect 1894 2667 1900 2668
rect 1894 2663 1895 2667
rect 1899 2663 1900 2667
rect 1894 2662 1900 2663
rect 1982 2667 1988 2668
rect 1982 2663 1983 2667
rect 1987 2663 1988 2667
rect 1982 2662 1988 2663
rect 2070 2667 2076 2668
rect 2070 2663 2071 2667
rect 2075 2663 2076 2667
rect 2070 2662 2076 2663
rect 2158 2667 2164 2668
rect 2158 2663 2159 2667
rect 2163 2663 2164 2667
rect 2158 2662 2164 2663
rect 2246 2667 2252 2668
rect 2246 2663 2247 2667
rect 2251 2663 2252 2667
rect 2246 2662 2252 2663
rect 2334 2667 2340 2668
rect 2334 2663 2335 2667
rect 2339 2663 2340 2667
rect 2334 2662 2340 2663
rect 2422 2667 2428 2668
rect 2422 2663 2423 2667
rect 2427 2663 2428 2667
rect 2422 2662 2428 2663
rect 2510 2667 2516 2668
rect 2510 2663 2511 2667
rect 2515 2663 2516 2667
rect 2510 2662 2516 2663
rect 2598 2667 2604 2668
rect 2598 2663 2599 2667
rect 2603 2663 2604 2667
rect 2598 2662 2604 2663
rect 2686 2667 2692 2668
rect 2686 2663 2687 2667
rect 2691 2663 2692 2667
rect 2686 2662 2692 2663
rect 2774 2667 2780 2668
rect 2774 2663 2775 2667
rect 2779 2663 2780 2667
rect 2774 2662 2780 2663
rect 2862 2667 2868 2668
rect 2862 2663 2863 2667
rect 2867 2663 2868 2667
rect 2862 2662 2868 2663
rect 2950 2667 2956 2668
rect 2950 2663 2951 2667
rect 2955 2663 2956 2667
rect 2950 2662 2956 2663
rect 3038 2667 3044 2668
rect 3038 2663 3039 2667
rect 3043 2663 3044 2667
rect 3038 2662 3044 2663
rect 3126 2667 3132 2668
rect 3126 2663 3127 2667
rect 3131 2663 3132 2667
rect 3126 2662 3132 2663
rect 3214 2667 3220 2668
rect 3214 2663 3215 2667
rect 3219 2663 3220 2667
rect 3214 2662 3220 2663
rect 3302 2667 3308 2668
rect 3302 2663 3303 2667
rect 3307 2663 3308 2667
rect 3302 2662 3308 2663
rect 3398 2667 3404 2668
rect 3398 2663 3399 2667
rect 3403 2663 3404 2667
rect 3398 2662 3404 2663
rect 3486 2667 3492 2668
rect 3486 2663 3487 2667
rect 3491 2663 3492 2667
rect 3486 2662 3492 2663
rect 327 2659 333 2660
rect 327 2658 328 2659
rect 110 2656 116 2657
rect 277 2656 328 2658
rect 110 2652 111 2656
rect 115 2652 116 2656
rect 327 2655 328 2656
rect 332 2655 333 2659
rect 455 2659 461 2660
rect 455 2658 456 2659
rect 397 2656 456 2658
rect 327 2654 333 2655
rect 455 2655 456 2656
rect 460 2655 461 2659
rect 575 2659 581 2660
rect 575 2658 576 2659
rect 525 2656 576 2658
rect 455 2654 461 2655
rect 575 2655 576 2656
rect 580 2655 581 2659
rect 814 2659 820 2660
rect 814 2658 815 2659
rect 765 2656 815 2658
rect 575 2654 581 2655
rect 814 2655 815 2656
rect 819 2655 820 2659
rect 927 2659 933 2660
rect 927 2658 928 2659
rect 885 2656 928 2658
rect 814 2654 820 2655
rect 927 2655 928 2656
rect 932 2655 933 2659
rect 1039 2659 1045 2660
rect 1039 2658 1040 2659
rect 997 2656 1040 2658
rect 927 2654 933 2655
rect 1039 2655 1040 2656
rect 1044 2655 1045 2659
rect 1138 2659 1144 2660
rect 1138 2658 1139 2659
rect 1109 2656 1139 2658
rect 1039 2654 1045 2655
rect 1138 2655 1139 2656
rect 1143 2655 1144 2659
rect 1263 2659 1269 2660
rect 1263 2658 1264 2659
rect 1221 2656 1264 2658
rect 1138 2654 1144 2655
rect 1263 2655 1264 2656
rect 1268 2655 1269 2659
rect 1263 2654 1269 2655
rect 1822 2656 1828 2657
rect 110 2651 116 2652
rect 1822 2652 1823 2656
rect 1827 2652 1828 2656
rect 1822 2651 1828 2652
rect 1903 2655 1909 2656
rect 1903 2651 1904 2655
rect 1908 2654 1909 2655
rect 1950 2655 1956 2656
rect 1950 2654 1951 2655
rect 1908 2652 1951 2654
rect 1908 2651 1909 2652
rect 1903 2650 1909 2651
rect 1950 2651 1951 2652
rect 1955 2651 1956 2655
rect 1950 2650 1956 2651
rect 1967 2655 1973 2656
rect 1967 2651 1968 2655
rect 1972 2654 1973 2655
rect 1991 2655 1997 2656
rect 1991 2654 1992 2655
rect 1972 2652 1992 2654
rect 1972 2651 1973 2652
rect 1967 2650 1973 2651
rect 1991 2651 1992 2652
rect 1996 2651 1997 2655
rect 1991 2650 1997 2651
rect 2042 2655 2048 2656
rect 2042 2651 2043 2655
rect 2047 2654 2048 2655
rect 2079 2655 2085 2656
rect 2079 2654 2080 2655
rect 2047 2652 2080 2654
rect 2047 2651 2048 2652
rect 2042 2650 2048 2651
rect 2079 2651 2080 2652
rect 2084 2651 2085 2655
rect 2079 2650 2085 2651
rect 2143 2655 2149 2656
rect 2143 2651 2144 2655
rect 2148 2654 2149 2655
rect 2167 2655 2173 2656
rect 2167 2654 2168 2655
rect 2148 2652 2168 2654
rect 2148 2651 2149 2652
rect 2143 2650 2149 2651
rect 2167 2651 2168 2652
rect 2172 2651 2173 2655
rect 2167 2650 2173 2651
rect 2231 2655 2237 2656
rect 2231 2651 2232 2655
rect 2236 2654 2237 2655
rect 2255 2655 2261 2656
rect 2255 2654 2256 2655
rect 2236 2652 2256 2654
rect 2236 2651 2237 2652
rect 2231 2650 2237 2651
rect 2255 2651 2256 2652
rect 2260 2651 2261 2655
rect 2255 2650 2261 2651
rect 2319 2655 2325 2656
rect 2319 2651 2320 2655
rect 2324 2654 2325 2655
rect 2343 2655 2349 2656
rect 2343 2654 2344 2655
rect 2324 2652 2344 2654
rect 2324 2651 2325 2652
rect 2319 2650 2325 2651
rect 2343 2651 2344 2652
rect 2348 2651 2349 2655
rect 2343 2650 2349 2651
rect 2407 2655 2413 2656
rect 2407 2651 2408 2655
rect 2412 2654 2413 2655
rect 2431 2655 2437 2656
rect 2431 2654 2432 2655
rect 2412 2652 2432 2654
rect 2412 2651 2413 2652
rect 2407 2650 2413 2651
rect 2431 2651 2432 2652
rect 2436 2651 2437 2655
rect 2431 2650 2437 2651
rect 2495 2655 2501 2656
rect 2495 2651 2496 2655
rect 2500 2654 2501 2655
rect 2519 2655 2525 2656
rect 2519 2654 2520 2655
rect 2500 2652 2520 2654
rect 2500 2651 2501 2652
rect 2495 2650 2501 2651
rect 2519 2651 2520 2652
rect 2524 2651 2525 2655
rect 2519 2650 2525 2651
rect 2583 2655 2589 2656
rect 2583 2651 2584 2655
rect 2588 2654 2589 2655
rect 2607 2655 2613 2656
rect 2607 2654 2608 2655
rect 2588 2652 2608 2654
rect 2588 2651 2589 2652
rect 2583 2650 2589 2651
rect 2607 2651 2608 2652
rect 2612 2651 2613 2655
rect 2607 2650 2613 2651
rect 2671 2655 2677 2656
rect 2671 2651 2672 2655
rect 2676 2654 2677 2655
rect 2695 2655 2701 2656
rect 2695 2654 2696 2655
rect 2676 2652 2696 2654
rect 2676 2651 2677 2652
rect 2671 2650 2677 2651
rect 2695 2651 2696 2652
rect 2700 2651 2701 2655
rect 2695 2650 2701 2651
rect 2759 2655 2765 2656
rect 2759 2651 2760 2655
rect 2764 2654 2765 2655
rect 2783 2655 2789 2656
rect 2783 2654 2784 2655
rect 2764 2652 2784 2654
rect 2764 2651 2765 2652
rect 2759 2650 2765 2651
rect 2783 2651 2784 2652
rect 2788 2651 2789 2655
rect 2783 2650 2789 2651
rect 2847 2655 2853 2656
rect 2847 2651 2848 2655
rect 2852 2654 2853 2655
rect 2871 2655 2877 2656
rect 2871 2654 2872 2655
rect 2852 2652 2872 2654
rect 2852 2651 2853 2652
rect 2847 2650 2853 2651
rect 2871 2651 2872 2652
rect 2876 2651 2877 2655
rect 2871 2650 2877 2651
rect 2935 2655 2941 2656
rect 2935 2651 2936 2655
rect 2940 2654 2941 2655
rect 2959 2655 2965 2656
rect 2959 2654 2960 2655
rect 2940 2652 2960 2654
rect 2940 2651 2941 2652
rect 2935 2650 2941 2651
rect 2959 2651 2960 2652
rect 2964 2651 2965 2655
rect 2959 2650 2965 2651
rect 3023 2655 3029 2656
rect 3023 2651 3024 2655
rect 3028 2654 3029 2655
rect 3047 2655 3053 2656
rect 3047 2654 3048 2655
rect 3028 2652 3048 2654
rect 3028 2651 3029 2652
rect 3023 2650 3029 2651
rect 3047 2651 3048 2652
rect 3052 2651 3053 2655
rect 3047 2650 3053 2651
rect 3111 2655 3117 2656
rect 3111 2651 3112 2655
rect 3116 2654 3117 2655
rect 3135 2655 3141 2656
rect 3135 2654 3136 2655
rect 3116 2652 3136 2654
rect 3116 2651 3117 2652
rect 3111 2650 3117 2651
rect 3135 2651 3136 2652
rect 3140 2651 3141 2655
rect 3135 2650 3141 2651
rect 3199 2655 3205 2656
rect 3199 2651 3200 2655
rect 3204 2654 3205 2655
rect 3223 2655 3229 2656
rect 3223 2654 3224 2655
rect 3204 2652 3224 2654
rect 3204 2651 3205 2652
rect 3199 2650 3205 2651
rect 3223 2651 3224 2652
rect 3228 2651 3229 2655
rect 3223 2650 3229 2651
rect 3287 2655 3293 2656
rect 3287 2651 3288 2655
rect 3292 2654 3293 2655
rect 3311 2655 3317 2656
rect 3311 2654 3312 2655
rect 3292 2652 3312 2654
rect 3292 2651 3293 2652
rect 3287 2650 3293 2651
rect 3311 2651 3312 2652
rect 3316 2651 3317 2655
rect 3311 2650 3317 2651
rect 3383 2655 3389 2656
rect 3383 2651 3384 2655
rect 3388 2654 3389 2655
rect 3407 2655 3413 2656
rect 3407 2654 3408 2655
rect 3388 2652 3408 2654
rect 3388 2651 3389 2652
rect 3383 2650 3389 2651
rect 3407 2651 3408 2652
rect 3412 2651 3413 2655
rect 3407 2650 3413 2651
rect 3495 2655 3504 2656
rect 3495 2651 3496 2655
rect 3503 2651 3504 2655
rect 3495 2650 3504 2651
rect 222 2643 228 2644
rect 222 2639 223 2643
rect 227 2639 228 2643
rect 222 2638 228 2639
rect 342 2643 348 2644
rect 342 2639 343 2643
rect 347 2639 348 2643
rect 342 2638 348 2639
rect 470 2643 476 2644
rect 470 2639 471 2643
rect 475 2639 476 2643
rect 470 2638 476 2639
rect 590 2643 596 2644
rect 590 2639 591 2643
rect 595 2639 596 2643
rect 590 2638 596 2639
rect 710 2643 716 2644
rect 710 2639 711 2643
rect 715 2639 716 2643
rect 710 2638 716 2639
rect 830 2643 836 2644
rect 830 2639 831 2643
rect 835 2639 836 2643
rect 830 2638 836 2639
rect 942 2643 948 2644
rect 942 2639 943 2643
rect 947 2639 948 2643
rect 942 2638 948 2639
rect 1054 2643 1060 2644
rect 1054 2639 1055 2643
rect 1059 2639 1060 2643
rect 1054 2638 1060 2639
rect 1166 2643 1172 2644
rect 1166 2639 1167 2643
rect 1171 2639 1172 2643
rect 1166 2638 1172 2639
rect 1278 2643 1284 2644
rect 1278 2639 1279 2643
rect 1283 2639 1284 2643
rect 1278 2638 1284 2639
rect 231 2631 240 2632
rect 231 2627 232 2631
rect 239 2627 240 2631
rect 231 2626 240 2627
rect 327 2631 333 2632
rect 327 2627 328 2631
rect 332 2630 333 2631
rect 351 2631 357 2632
rect 351 2630 352 2631
rect 332 2628 352 2630
rect 332 2627 333 2628
rect 327 2626 333 2627
rect 351 2627 352 2628
rect 356 2627 357 2631
rect 351 2626 357 2627
rect 455 2631 461 2632
rect 455 2627 456 2631
rect 460 2630 461 2631
rect 479 2631 485 2632
rect 479 2630 480 2631
rect 460 2628 480 2630
rect 460 2627 461 2628
rect 455 2626 461 2627
rect 479 2627 480 2628
rect 484 2627 485 2631
rect 479 2626 485 2627
rect 575 2631 581 2632
rect 575 2627 576 2631
rect 580 2630 581 2631
rect 599 2631 605 2632
rect 599 2630 600 2631
rect 580 2628 600 2630
rect 580 2627 581 2628
rect 575 2626 581 2627
rect 599 2627 600 2628
rect 604 2627 605 2631
rect 599 2626 605 2627
rect 711 2631 717 2632
rect 711 2627 712 2631
rect 716 2630 717 2631
rect 719 2631 725 2632
rect 719 2630 720 2631
rect 716 2628 720 2630
rect 716 2627 717 2628
rect 711 2626 717 2627
rect 719 2627 720 2628
rect 724 2627 725 2631
rect 719 2626 725 2627
rect 839 2631 848 2632
rect 839 2627 840 2631
rect 847 2627 848 2631
rect 839 2626 848 2627
rect 927 2631 933 2632
rect 927 2627 928 2631
rect 932 2630 933 2631
rect 951 2631 957 2632
rect 951 2630 952 2631
rect 932 2628 952 2630
rect 932 2627 933 2628
rect 927 2626 933 2627
rect 951 2627 952 2628
rect 956 2627 957 2631
rect 951 2626 957 2627
rect 1039 2631 1045 2632
rect 1039 2627 1040 2631
rect 1044 2630 1045 2631
rect 1063 2631 1069 2632
rect 1063 2630 1064 2631
rect 1044 2628 1064 2630
rect 1044 2627 1045 2628
rect 1039 2626 1045 2627
rect 1063 2627 1064 2628
rect 1068 2627 1069 2631
rect 1063 2626 1069 2627
rect 1175 2631 1184 2632
rect 1175 2627 1176 2631
rect 1183 2627 1184 2631
rect 1175 2626 1184 2627
rect 1263 2631 1269 2632
rect 1263 2627 1264 2631
rect 1268 2630 1269 2631
rect 1287 2631 1293 2632
rect 1287 2630 1288 2631
rect 1268 2628 1288 2630
rect 1268 2627 1269 2628
rect 1263 2626 1269 2627
rect 1287 2627 1288 2628
rect 1292 2627 1293 2631
rect 2498 2631 2504 2632
rect 2498 2630 2499 2631
rect 1287 2626 1293 2627
rect 2216 2628 2499 2630
rect 1247 2623 1253 2624
rect 1247 2622 1248 2623
rect 808 2620 1248 2622
rect 479 2615 488 2616
rect 479 2611 480 2615
rect 487 2611 488 2615
rect 479 2610 488 2611
rect 535 2615 541 2616
rect 535 2611 536 2615
rect 540 2614 541 2615
rect 567 2615 573 2616
rect 567 2614 568 2615
rect 540 2612 568 2614
rect 540 2611 541 2612
rect 535 2610 541 2611
rect 567 2611 568 2612
rect 572 2611 573 2615
rect 567 2610 573 2611
rect 623 2615 629 2616
rect 623 2611 624 2615
rect 628 2614 629 2615
rect 655 2615 661 2616
rect 655 2614 656 2615
rect 628 2612 656 2614
rect 628 2611 629 2612
rect 623 2610 629 2611
rect 655 2611 656 2612
rect 660 2611 661 2615
rect 655 2610 661 2611
rect 743 2615 749 2616
rect 743 2611 744 2615
rect 748 2614 749 2615
rect 808 2614 810 2620
rect 1247 2619 1248 2620
rect 1252 2619 1253 2623
rect 1247 2618 1253 2619
rect 2167 2623 2173 2624
rect 2167 2619 2168 2623
rect 2172 2622 2173 2623
rect 2216 2622 2218 2628
rect 2498 2627 2499 2628
rect 2503 2627 2504 2631
rect 3078 2631 3084 2632
rect 3078 2630 3079 2631
rect 2498 2626 2504 2627
rect 2920 2628 3079 2630
rect 2172 2620 2218 2622
rect 2223 2623 2229 2624
rect 2172 2619 2173 2620
rect 2167 2618 2173 2619
rect 2223 2619 2224 2623
rect 2228 2622 2229 2623
rect 2287 2623 2293 2624
rect 2287 2622 2288 2623
rect 2228 2620 2288 2622
rect 2228 2619 2229 2620
rect 2223 2618 2229 2619
rect 2287 2619 2288 2620
rect 2292 2619 2293 2623
rect 2287 2618 2293 2619
rect 2351 2623 2357 2624
rect 2351 2619 2352 2623
rect 2356 2622 2357 2623
rect 2423 2623 2429 2624
rect 2423 2622 2424 2623
rect 2356 2620 2424 2622
rect 2356 2619 2357 2620
rect 2351 2618 2357 2619
rect 2423 2619 2424 2620
rect 2428 2619 2429 2623
rect 2423 2618 2429 2619
rect 2487 2623 2493 2624
rect 2487 2619 2488 2623
rect 2492 2622 2493 2623
rect 2559 2623 2565 2624
rect 2559 2622 2560 2623
rect 2492 2620 2560 2622
rect 2492 2619 2493 2620
rect 2487 2618 2493 2619
rect 2559 2619 2560 2620
rect 2564 2619 2565 2623
rect 2559 2618 2565 2619
rect 2631 2623 2637 2624
rect 2631 2619 2632 2623
rect 2636 2622 2637 2623
rect 2703 2623 2709 2624
rect 2703 2622 2704 2623
rect 2636 2620 2704 2622
rect 2636 2619 2637 2620
rect 2631 2618 2637 2619
rect 2703 2619 2704 2620
rect 2708 2619 2709 2623
rect 2703 2618 2709 2619
rect 2855 2623 2861 2624
rect 2855 2619 2856 2623
rect 2860 2622 2861 2623
rect 2920 2622 2922 2628
rect 3078 2627 3079 2628
rect 3083 2627 3084 2631
rect 3078 2626 3084 2627
rect 2860 2620 2922 2622
rect 2927 2623 2933 2624
rect 2860 2619 2861 2620
rect 2855 2618 2861 2619
rect 2927 2619 2928 2623
rect 2932 2622 2933 2623
rect 3007 2623 3013 2624
rect 3007 2622 3008 2623
rect 2932 2620 3008 2622
rect 2932 2619 2933 2620
rect 2927 2618 2933 2619
rect 3007 2619 3008 2620
rect 3012 2619 3013 2623
rect 3007 2618 3013 2619
rect 3166 2623 3173 2624
rect 3166 2619 3167 2623
rect 3172 2619 3173 2623
rect 3166 2618 3173 2619
rect 748 2612 810 2614
rect 814 2615 820 2616
rect 748 2611 749 2612
rect 743 2610 749 2611
rect 814 2611 815 2615
rect 819 2614 820 2615
rect 831 2615 837 2616
rect 831 2614 832 2615
rect 819 2612 832 2614
rect 819 2611 820 2612
rect 814 2610 820 2611
rect 831 2611 832 2612
rect 836 2611 837 2615
rect 831 2610 837 2611
rect 887 2615 893 2616
rect 887 2611 888 2615
rect 892 2614 893 2615
rect 919 2615 925 2616
rect 919 2614 920 2615
rect 892 2612 920 2614
rect 892 2611 893 2612
rect 887 2610 893 2611
rect 919 2611 920 2612
rect 924 2611 925 2615
rect 919 2610 925 2611
rect 975 2615 981 2616
rect 975 2611 976 2615
rect 980 2614 981 2615
rect 1007 2615 1013 2616
rect 1007 2614 1008 2615
rect 980 2612 1008 2614
rect 980 2611 981 2612
rect 975 2610 981 2611
rect 1007 2611 1008 2612
rect 1012 2611 1013 2615
rect 1007 2610 1013 2611
rect 1063 2615 1069 2616
rect 1063 2611 1064 2615
rect 1068 2614 1069 2615
rect 1095 2615 1101 2616
rect 1095 2614 1096 2615
rect 1068 2612 1096 2614
rect 1068 2611 1069 2612
rect 1063 2610 1069 2611
rect 1095 2611 1096 2612
rect 1100 2611 1101 2615
rect 1095 2610 1101 2611
rect 1138 2615 1144 2616
rect 1138 2611 1139 2615
rect 1143 2614 1144 2615
rect 1183 2615 1189 2616
rect 1183 2614 1184 2615
rect 1143 2612 1184 2614
rect 1143 2611 1144 2612
rect 1138 2610 1144 2611
rect 1183 2611 1184 2612
rect 1188 2611 1189 2615
rect 1183 2610 1189 2611
rect 1239 2615 1245 2616
rect 1239 2611 1240 2615
rect 1244 2614 1245 2615
rect 1271 2615 1277 2616
rect 1271 2614 1272 2615
rect 1244 2612 1272 2614
rect 1244 2611 1245 2612
rect 1239 2610 1245 2611
rect 1271 2611 1272 2612
rect 1276 2611 1277 2615
rect 1271 2610 1277 2611
rect 2158 2613 2164 2614
rect 2158 2609 2159 2613
rect 2163 2609 2164 2613
rect 2158 2608 2164 2609
rect 2278 2613 2284 2614
rect 2278 2609 2279 2613
rect 2283 2609 2284 2613
rect 2278 2608 2284 2609
rect 2414 2613 2420 2614
rect 2414 2609 2415 2613
rect 2419 2609 2420 2613
rect 2414 2608 2420 2609
rect 2550 2613 2556 2614
rect 2550 2609 2551 2613
rect 2555 2609 2556 2613
rect 2550 2608 2556 2609
rect 2694 2613 2700 2614
rect 2694 2609 2695 2613
rect 2699 2609 2700 2613
rect 2694 2608 2700 2609
rect 2846 2613 2852 2614
rect 2846 2609 2847 2613
rect 2851 2609 2852 2613
rect 2846 2608 2852 2609
rect 2998 2613 3004 2614
rect 2998 2609 2999 2613
rect 3003 2609 3004 2613
rect 2998 2608 3004 2609
rect 3158 2613 3164 2614
rect 3158 2609 3159 2613
rect 3163 2609 3164 2613
rect 3158 2608 3164 2609
rect 470 2605 476 2606
rect 470 2601 471 2605
rect 475 2601 476 2605
rect 470 2600 476 2601
rect 558 2605 564 2606
rect 558 2601 559 2605
rect 563 2601 564 2605
rect 558 2600 564 2601
rect 646 2605 652 2606
rect 646 2601 647 2605
rect 651 2601 652 2605
rect 646 2600 652 2601
rect 734 2605 740 2606
rect 734 2601 735 2605
rect 739 2601 740 2605
rect 734 2600 740 2601
rect 822 2605 828 2606
rect 822 2601 823 2605
rect 827 2601 828 2605
rect 822 2600 828 2601
rect 910 2605 916 2606
rect 910 2601 911 2605
rect 915 2601 916 2605
rect 910 2600 916 2601
rect 998 2605 1004 2606
rect 998 2601 999 2605
rect 1003 2601 1004 2605
rect 998 2600 1004 2601
rect 1086 2605 1092 2606
rect 1086 2601 1087 2605
rect 1091 2601 1092 2605
rect 1086 2600 1092 2601
rect 1174 2605 1180 2606
rect 1174 2601 1175 2605
rect 1179 2601 1180 2605
rect 1174 2600 1180 2601
rect 1262 2605 1268 2606
rect 1262 2601 1263 2605
rect 1267 2601 1268 2605
rect 1262 2600 1268 2601
rect 1862 2600 1868 2601
rect 3574 2600 3580 2601
rect 1862 2596 1863 2600
rect 1867 2596 1868 2600
rect 2223 2599 2229 2600
rect 2223 2598 2224 2599
rect 2213 2596 2224 2598
rect 1862 2595 1868 2596
rect 2223 2595 2224 2596
rect 2228 2595 2229 2599
rect 2351 2599 2357 2600
rect 2351 2598 2352 2599
rect 2333 2596 2352 2598
rect 2223 2594 2229 2595
rect 2351 2595 2352 2596
rect 2356 2595 2357 2599
rect 2487 2599 2493 2600
rect 2487 2598 2488 2599
rect 2469 2596 2488 2598
rect 2351 2594 2357 2595
rect 2487 2595 2488 2596
rect 2492 2595 2493 2599
rect 2631 2599 2637 2600
rect 2631 2598 2632 2599
rect 2605 2596 2632 2598
rect 2487 2594 2493 2595
rect 2631 2595 2632 2596
rect 2636 2595 2637 2599
rect 2927 2599 2933 2600
rect 2927 2598 2928 2599
rect 2901 2596 2928 2598
rect 2631 2594 2637 2595
rect 2642 2595 2648 2596
rect 110 2592 116 2593
rect 1822 2592 1828 2593
rect 110 2588 111 2592
rect 115 2588 116 2592
rect 535 2591 541 2592
rect 535 2590 536 2591
rect 525 2588 536 2590
rect 110 2587 116 2588
rect 535 2587 536 2588
rect 540 2587 541 2591
rect 623 2591 629 2592
rect 623 2590 624 2591
rect 613 2588 624 2590
rect 535 2586 541 2587
rect 623 2587 624 2588
rect 628 2587 629 2591
rect 711 2591 717 2592
rect 711 2590 712 2591
rect 701 2588 712 2590
rect 623 2586 629 2587
rect 711 2587 712 2588
rect 716 2587 717 2591
rect 887 2591 893 2592
rect 887 2590 888 2591
rect 877 2588 888 2590
rect 711 2586 717 2587
rect 887 2587 888 2588
rect 892 2587 893 2591
rect 975 2591 981 2592
rect 975 2590 976 2591
rect 965 2588 976 2590
rect 887 2586 893 2587
rect 975 2587 976 2588
rect 980 2587 981 2591
rect 1063 2591 1069 2592
rect 1063 2590 1064 2591
rect 1053 2588 1064 2590
rect 975 2586 981 2587
rect 1063 2587 1064 2588
rect 1068 2587 1069 2591
rect 1239 2591 1245 2592
rect 1239 2590 1240 2591
rect 1229 2588 1240 2590
rect 1063 2586 1069 2587
rect 1239 2587 1240 2588
rect 1244 2587 1245 2591
rect 1822 2588 1823 2592
rect 1827 2588 1828 2592
rect 2642 2591 2643 2595
rect 2647 2594 2648 2595
rect 2927 2595 2928 2596
rect 2932 2595 2933 2599
rect 3574 2596 3575 2600
rect 3579 2596 3580 2600
rect 2927 2594 2933 2595
rect 3078 2595 3084 2596
rect 3574 2595 3580 2596
rect 2647 2592 2713 2594
rect 2647 2591 2648 2592
rect 2642 2590 2648 2591
rect 3078 2591 3079 2595
rect 3083 2594 3084 2595
rect 3083 2592 3177 2594
rect 3083 2591 3084 2592
rect 3078 2590 3084 2591
rect 1239 2586 1245 2587
rect 1247 2587 1253 2588
rect 1822 2587 1828 2588
rect 1247 2583 1248 2587
rect 1252 2586 1253 2587
rect 1252 2584 1281 2586
rect 1252 2583 1253 2584
rect 1247 2582 1253 2583
rect 1862 2583 1868 2584
rect 1862 2579 1863 2583
rect 1867 2579 1868 2583
rect 1862 2578 1868 2579
rect 3574 2583 3580 2584
rect 3574 2579 3575 2583
rect 3579 2579 3580 2583
rect 3574 2578 3580 2579
rect 110 2575 116 2576
rect 110 2571 111 2575
rect 115 2571 116 2575
rect 110 2570 116 2571
rect 714 2575 720 2576
rect 714 2571 715 2575
rect 719 2574 720 2575
rect 1822 2575 1828 2576
rect 719 2572 745 2574
rect 1060 2572 1097 2574
rect 719 2571 720 2572
rect 714 2570 720 2571
rect 462 2565 468 2566
rect 462 2561 463 2565
rect 467 2561 468 2565
rect 462 2560 468 2561
rect 550 2565 556 2566
rect 550 2561 551 2565
rect 555 2561 556 2565
rect 550 2560 556 2561
rect 638 2565 644 2566
rect 638 2561 639 2565
rect 643 2561 644 2565
rect 638 2560 644 2561
rect 726 2565 732 2566
rect 726 2561 727 2565
rect 731 2561 732 2565
rect 726 2560 732 2561
rect 814 2565 820 2566
rect 814 2561 815 2565
rect 819 2561 820 2565
rect 814 2560 820 2561
rect 902 2565 908 2566
rect 902 2561 903 2565
rect 907 2561 908 2565
rect 902 2560 908 2561
rect 990 2565 996 2566
rect 990 2561 991 2565
rect 995 2561 996 2565
rect 990 2560 996 2561
rect 954 2559 960 2560
rect 954 2555 955 2559
rect 959 2558 960 2559
rect 1060 2558 1062 2572
rect 1822 2571 1823 2575
rect 1827 2571 1828 2575
rect 1822 2570 1828 2571
rect 2150 2573 2156 2574
rect 2150 2569 2151 2573
rect 2155 2569 2156 2573
rect 2150 2568 2156 2569
rect 2270 2573 2276 2574
rect 2270 2569 2271 2573
rect 2275 2569 2276 2573
rect 2270 2568 2276 2569
rect 2406 2573 2412 2574
rect 2406 2569 2407 2573
rect 2411 2569 2412 2573
rect 2406 2568 2412 2569
rect 2542 2573 2548 2574
rect 2542 2569 2543 2573
rect 2547 2569 2548 2573
rect 2542 2568 2548 2569
rect 2686 2573 2692 2574
rect 2686 2569 2687 2573
rect 2691 2569 2692 2573
rect 2686 2568 2692 2569
rect 2838 2573 2844 2574
rect 2838 2569 2839 2573
rect 2843 2569 2844 2573
rect 2838 2568 2844 2569
rect 2990 2573 2996 2574
rect 2990 2569 2991 2573
rect 2995 2569 2996 2573
rect 2990 2568 2996 2569
rect 3150 2573 3156 2574
rect 3150 2569 3151 2573
rect 3155 2569 3156 2573
rect 3150 2568 3156 2569
rect 3018 2567 3024 2568
rect 1078 2565 1084 2566
rect 1078 2561 1079 2565
rect 1083 2561 1084 2565
rect 1078 2560 1084 2561
rect 1166 2565 1172 2566
rect 1166 2561 1167 2565
rect 1171 2561 1172 2565
rect 1166 2560 1172 2561
rect 1254 2565 1260 2566
rect 1254 2561 1255 2565
rect 1259 2561 1260 2565
rect 3018 2563 3019 2567
rect 3023 2566 3024 2567
rect 3039 2567 3045 2568
rect 3039 2566 3040 2567
rect 3023 2564 3040 2566
rect 3023 2563 3024 2564
rect 3018 2562 3024 2563
rect 3039 2563 3040 2564
rect 3044 2563 3045 2567
rect 3039 2562 3045 2563
rect 1254 2560 1260 2561
rect 959 2556 1062 2558
rect 959 2555 960 2556
rect 954 2554 960 2555
rect 2102 2551 2108 2552
rect 2102 2547 2103 2551
rect 2107 2547 2108 2551
rect 2102 2546 2108 2547
rect 2198 2551 2204 2552
rect 2198 2547 2199 2551
rect 2203 2547 2204 2551
rect 2198 2546 2204 2547
rect 2310 2551 2316 2552
rect 2310 2547 2311 2551
rect 2315 2547 2316 2551
rect 2310 2546 2316 2547
rect 2430 2551 2436 2552
rect 2430 2547 2431 2551
rect 2435 2547 2436 2551
rect 2430 2546 2436 2547
rect 2558 2551 2564 2552
rect 2558 2547 2559 2551
rect 2563 2547 2564 2551
rect 2558 2546 2564 2547
rect 2694 2551 2700 2552
rect 2694 2547 2695 2551
rect 2699 2547 2700 2551
rect 2694 2546 2700 2547
rect 2846 2551 2852 2552
rect 2846 2547 2847 2551
rect 2851 2547 2852 2551
rect 2846 2546 2852 2547
rect 2998 2551 3004 2552
rect 2998 2547 2999 2551
rect 3003 2547 3004 2551
rect 2998 2546 3004 2547
rect 3158 2551 3164 2552
rect 3158 2547 3159 2551
rect 3163 2547 3164 2551
rect 3158 2546 3164 2547
rect 3326 2551 3332 2552
rect 3326 2547 3327 2551
rect 3331 2547 3332 2551
rect 3326 2546 3332 2547
rect 3478 2551 3484 2552
rect 3478 2547 3479 2551
rect 3483 2547 3484 2551
rect 3478 2546 3484 2547
rect 2498 2543 2504 2544
rect 1862 2541 1868 2542
rect 1862 2537 1863 2541
rect 1867 2537 1868 2541
rect 2498 2539 2499 2543
rect 2503 2542 2504 2543
rect 2503 2540 2577 2542
rect 3168 2540 3177 2542
rect 3574 2541 3580 2542
rect 2503 2539 2504 2540
rect 2498 2538 2504 2539
rect 3166 2539 3172 2540
rect 1862 2536 1868 2537
rect 494 2535 500 2536
rect 494 2531 495 2535
rect 499 2531 500 2535
rect 494 2530 500 2531
rect 582 2535 588 2536
rect 582 2531 583 2535
rect 587 2531 588 2535
rect 582 2530 588 2531
rect 670 2535 676 2536
rect 670 2531 671 2535
rect 675 2531 676 2535
rect 670 2530 676 2531
rect 758 2535 764 2536
rect 758 2531 759 2535
rect 763 2531 764 2535
rect 758 2530 764 2531
rect 846 2535 852 2536
rect 846 2531 847 2535
rect 851 2531 852 2535
rect 846 2530 852 2531
rect 934 2535 940 2536
rect 934 2531 935 2535
rect 939 2531 940 2535
rect 934 2530 940 2531
rect 1022 2535 1028 2536
rect 1022 2531 1023 2535
rect 1027 2531 1028 2535
rect 1022 2530 1028 2531
rect 1110 2535 1116 2536
rect 1110 2531 1111 2535
rect 1115 2531 1116 2535
rect 1110 2530 1116 2531
rect 1198 2535 1204 2536
rect 1198 2531 1199 2535
rect 1203 2531 1204 2535
rect 1198 2530 1204 2531
rect 1286 2535 1292 2536
rect 1286 2531 1287 2535
rect 1291 2531 1292 2535
rect 3166 2535 3167 2539
rect 3171 2535 3172 2539
rect 3574 2537 3575 2541
rect 3579 2537 3580 2541
rect 3574 2536 3580 2537
rect 3166 2534 3172 2535
rect 1286 2530 1292 2531
rect 482 2527 488 2528
rect 110 2525 116 2526
rect 110 2521 111 2525
rect 115 2521 116 2525
rect 482 2523 483 2527
rect 487 2526 488 2527
rect 838 2527 844 2528
rect 487 2524 513 2526
rect 487 2523 488 2524
rect 482 2522 488 2523
rect 838 2523 839 2527
rect 843 2526 844 2527
rect 1266 2527 1272 2528
rect 843 2524 865 2526
rect 843 2523 844 2524
rect 838 2522 844 2523
rect 1266 2523 1267 2527
rect 1271 2526 1272 2527
rect 2191 2527 2197 2528
rect 2191 2526 2192 2527
rect 1271 2524 1305 2526
rect 1822 2525 1828 2526
rect 1271 2523 1272 2524
rect 1266 2522 1272 2523
rect 110 2520 116 2521
rect 1822 2521 1823 2525
rect 1827 2521 1828 2525
rect 1822 2520 1828 2521
rect 1862 2524 1868 2525
rect 2165 2524 2192 2526
rect 1862 2520 1863 2524
rect 1867 2520 1868 2524
rect 2191 2523 2192 2524
rect 2196 2523 2197 2527
rect 2303 2527 2309 2528
rect 2303 2526 2304 2527
rect 2261 2524 2304 2526
rect 2191 2522 2197 2523
rect 2303 2523 2304 2524
rect 2308 2523 2309 2527
rect 2423 2527 2429 2528
rect 2423 2526 2424 2527
rect 2373 2524 2424 2526
rect 2303 2522 2309 2523
rect 2423 2523 2424 2524
rect 2428 2523 2429 2527
rect 2551 2527 2557 2528
rect 2551 2526 2552 2527
rect 2493 2524 2552 2526
rect 2423 2522 2429 2523
rect 2551 2523 2552 2524
rect 2556 2523 2557 2527
rect 2551 2522 2557 2523
rect 2626 2527 2632 2528
rect 2626 2523 2627 2527
rect 2631 2526 2632 2527
rect 2762 2527 2768 2528
rect 2631 2524 2721 2526
rect 2631 2523 2632 2524
rect 2626 2522 2632 2523
rect 2762 2523 2763 2527
rect 2767 2526 2768 2527
rect 2914 2527 2920 2528
rect 2767 2524 2873 2526
rect 2767 2523 2768 2524
rect 2762 2522 2768 2523
rect 2914 2523 2915 2527
rect 2919 2526 2920 2527
rect 3226 2527 3232 2528
rect 2919 2524 3025 2526
rect 2919 2523 2920 2524
rect 2914 2522 2920 2523
rect 3226 2523 3227 2527
rect 3231 2526 3232 2527
rect 3471 2527 3477 2528
rect 3231 2524 3353 2526
rect 3231 2523 3232 2524
rect 3226 2522 3232 2523
rect 3471 2523 3472 2527
rect 3476 2526 3477 2527
rect 3476 2524 3505 2526
rect 3574 2524 3580 2525
rect 3476 2523 3477 2524
rect 3471 2522 3477 2523
rect 1862 2519 1868 2520
rect 3574 2520 3575 2524
rect 3579 2520 3580 2524
rect 3574 2519 3580 2520
rect 562 2511 568 2512
rect 110 2508 116 2509
rect 110 2504 111 2508
rect 115 2504 116 2508
rect 562 2507 563 2511
rect 567 2510 568 2511
rect 751 2511 757 2512
rect 751 2510 752 2511
rect 567 2508 609 2510
rect 733 2508 752 2510
rect 567 2507 568 2508
rect 562 2506 568 2507
rect 751 2507 752 2508
rect 756 2507 757 2511
rect 839 2511 845 2512
rect 839 2510 840 2511
rect 821 2508 840 2510
rect 751 2506 757 2507
rect 839 2507 840 2508
rect 844 2507 845 2511
rect 1015 2511 1021 2512
rect 1015 2510 1016 2511
rect 997 2508 1016 2510
rect 839 2506 845 2507
rect 1015 2507 1016 2508
rect 1020 2507 1021 2511
rect 1103 2511 1109 2512
rect 1103 2510 1104 2511
rect 1085 2508 1104 2510
rect 1015 2506 1021 2507
rect 1103 2507 1104 2508
rect 1108 2507 1109 2511
rect 1191 2511 1197 2512
rect 1191 2510 1192 2511
rect 1173 2508 1192 2510
rect 1103 2506 1109 2507
rect 1191 2507 1192 2508
rect 1196 2507 1197 2511
rect 1279 2511 1285 2512
rect 1279 2510 1280 2511
rect 1261 2508 1280 2510
rect 1191 2506 1197 2507
rect 1279 2507 1280 2508
rect 1284 2507 1285 2511
rect 2110 2511 2116 2512
rect 1279 2506 1285 2507
rect 1822 2508 1828 2509
rect 110 2503 116 2504
rect 1822 2504 1823 2508
rect 1827 2504 1828 2508
rect 2110 2507 2111 2511
rect 2115 2507 2116 2511
rect 2110 2506 2116 2507
rect 2206 2511 2212 2512
rect 2206 2507 2207 2511
rect 2211 2507 2212 2511
rect 2206 2506 2212 2507
rect 2318 2511 2324 2512
rect 2318 2507 2319 2511
rect 2323 2507 2324 2511
rect 2318 2506 2324 2507
rect 2438 2511 2444 2512
rect 2438 2507 2439 2511
rect 2443 2507 2444 2511
rect 2438 2506 2444 2507
rect 2566 2511 2572 2512
rect 2566 2507 2567 2511
rect 2571 2507 2572 2511
rect 2566 2506 2572 2507
rect 2702 2511 2708 2512
rect 2702 2507 2703 2511
rect 2707 2507 2708 2511
rect 2702 2506 2708 2507
rect 2854 2511 2860 2512
rect 2854 2507 2855 2511
rect 2859 2507 2860 2511
rect 2854 2506 2860 2507
rect 3006 2511 3012 2512
rect 3006 2507 3007 2511
rect 3011 2507 3012 2511
rect 3006 2506 3012 2507
rect 3166 2511 3172 2512
rect 3166 2507 3167 2511
rect 3171 2507 3172 2511
rect 3166 2506 3172 2507
rect 3334 2511 3340 2512
rect 3334 2507 3335 2511
rect 3339 2507 3340 2511
rect 3334 2506 3340 2507
rect 3486 2511 3492 2512
rect 3486 2507 3487 2511
rect 3491 2507 3492 2511
rect 3486 2506 3492 2507
rect 1822 2503 1828 2504
rect 2119 2499 2125 2500
rect 502 2495 508 2496
rect 502 2491 503 2495
rect 507 2491 508 2495
rect 502 2490 508 2491
rect 590 2495 596 2496
rect 590 2491 591 2495
rect 595 2491 596 2495
rect 590 2490 596 2491
rect 678 2495 684 2496
rect 678 2491 679 2495
rect 683 2491 684 2495
rect 678 2490 684 2491
rect 766 2495 772 2496
rect 766 2491 767 2495
rect 771 2491 772 2495
rect 766 2490 772 2491
rect 854 2495 860 2496
rect 854 2491 855 2495
rect 859 2491 860 2495
rect 854 2490 860 2491
rect 942 2495 948 2496
rect 942 2491 943 2495
rect 947 2491 948 2495
rect 942 2490 948 2491
rect 1030 2495 1036 2496
rect 1030 2491 1031 2495
rect 1035 2491 1036 2495
rect 1030 2490 1036 2491
rect 1118 2495 1124 2496
rect 1118 2491 1119 2495
rect 1123 2491 1124 2495
rect 1118 2490 1124 2491
rect 1206 2495 1212 2496
rect 1206 2491 1207 2495
rect 1211 2491 1212 2495
rect 1206 2490 1212 2491
rect 1294 2495 1300 2496
rect 1294 2491 1295 2495
rect 1299 2491 1300 2495
rect 2119 2495 2120 2499
rect 2124 2498 2125 2499
rect 2191 2499 2197 2500
rect 2124 2496 2186 2498
rect 2124 2495 2125 2496
rect 2119 2494 2125 2495
rect 1294 2490 1300 2491
rect 2184 2490 2186 2496
rect 2191 2495 2192 2499
rect 2196 2498 2197 2499
rect 2215 2499 2221 2500
rect 2215 2498 2216 2499
rect 2196 2496 2216 2498
rect 2196 2495 2197 2496
rect 2191 2494 2197 2495
rect 2215 2495 2216 2496
rect 2220 2495 2221 2499
rect 2215 2494 2221 2495
rect 2303 2499 2309 2500
rect 2303 2495 2304 2499
rect 2308 2498 2309 2499
rect 2327 2499 2333 2500
rect 2327 2498 2328 2499
rect 2308 2496 2328 2498
rect 2308 2495 2309 2496
rect 2303 2494 2309 2495
rect 2327 2495 2328 2496
rect 2332 2495 2333 2499
rect 2327 2494 2333 2495
rect 2423 2499 2429 2500
rect 2423 2495 2424 2499
rect 2428 2498 2429 2499
rect 2447 2499 2453 2500
rect 2447 2498 2448 2499
rect 2428 2496 2448 2498
rect 2428 2495 2429 2496
rect 2423 2494 2429 2495
rect 2447 2495 2448 2496
rect 2452 2495 2453 2499
rect 2447 2494 2453 2495
rect 2551 2499 2557 2500
rect 2551 2495 2552 2499
rect 2556 2498 2557 2499
rect 2575 2499 2581 2500
rect 2575 2498 2576 2499
rect 2556 2496 2576 2498
rect 2556 2495 2557 2496
rect 2551 2494 2557 2495
rect 2575 2495 2576 2496
rect 2580 2495 2581 2499
rect 2575 2494 2581 2495
rect 2711 2499 2717 2500
rect 2711 2495 2712 2499
rect 2716 2498 2717 2499
rect 2762 2499 2768 2500
rect 2762 2498 2763 2499
rect 2716 2496 2763 2498
rect 2716 2495 2717 2496
rect 2711 2494 2717 2495
rect 2762 2495 2763 2496
rect 2767 2495 2768 2499
rect 2762 2494 2768 2495
rect 2863 2499 2869 2500
rect 2863 2495 2864 2499
rect 2868 2498 2869 2499
rect 2914 2499 2920 2500
rect 2914 2498 2915 2499
rect 2868 2496 2915 2498
rect 2868 2495 2869 2496
rect 2863 2494 2869 2495
rect 2914 2495 2915 2496
rect 2919 2495 2920 2499
rect 2914 2494 2920 2495
rect 3015 2499 3024 2500
rect 3015 2495 3016 2499
rect 3023 2495 3024 2499
rect 3015 2494 3024 2495
rect 3175 2499 3181 2500
rect 3175 2495 3176 2499
rect 3180 2498 3181 2499
rect 3226 2499 3232 2500
rect 3226 2498 3227 2499
rect 3180 2496 3227 2498
rect 3180 2495 3181 2496
rect 3175 2494 3181 2495
rect 3226 2495 3227 2496
rect 3231 2495 3232 2499
rect 3226 2494 3232 2495
rect 3343 2499 3349 2500
rect 3343 2495 3344 2499
rect 3348 2498 3349 2499
rect 3354 2499 3360 2500
rect 3354 2498 3355 2499
rect 3348 2496 3355 2498
rect 3348 2495 3349 2496
rect 3343 2494 3349 2495
rect 3354 2495 3355 2496
rect 3359 2495 3360 2499
rect 3354 2494 3360 2495
rect 3470 2499 3476 2500
rect 3470 2495 3471 2499
rect 3475 2498 3476 2499
rect 3495 2499 3501 2500
rect 3495 2498 3496 2499
rect 3475 2496 3496 2498
rect 3475 2495 3476 2496
rect 3470 2494 3476 2495
rect 3495 2495 3496 2496
rect 3500 2495 3501 2499
rect 3495 2494 3501 2495
rect 2359 2491 2365 2492
rect 2359 2490 2360 2491
rect 2184 2488 2360 2490
rect 2359 2487 2360 2488
rect 2364 2487 2365 2491
rect 2359 2486 2365 2487
rect 511 2483 517 2484
rect 511 2479 512 2483
rect 516 2482 517 2483
rect 562 2483 568 2484
rect 562 2482 563 2483
rect 516 2480 563 2482
rect 516 2479 517 2480
rect 511 2478 517 2479
rect 562 2479 563 2480
rect 567 2479 568 2483
rect 562 2478 568 2479
rect 582 2483 588 2484
rect 582 2479 583 2483
rect 587 2482 588 2483
rect 599 2483 605 2484
rect 599 2482 600 2483
rect 587 2480 600 2482
rect 587 2479 588 2480
rect 582 2478 588 2479
rect 599 2479 600 2480
rect 604 2479 605 2483
rect 599 2478 605 2479
rect 687 2483 693 2484
rect 687 2479 688 2483
rect 692 2482 693 2483
rect 714 2483 720 2484
rect 714 2482 715 2483
rect 692 2480 715 2482
rect 692 2479 693 2480
rect 687 2478 693 2479
rect 714 2479 715 2480
rect 719 2479 720 2483
rect 714 2478 720 2479
rect 751 2483 757 2484
rect 751 2479 752 2483
rect 756 2482 757 2483
rect 775 2483 781 2484
rect 775 2482 776 2483
rect 756 2480 776 2482
rect 756 2479 757 2480
rect 751 2478 757 2479
rect 775 2479 776 2480
rect 780 2479 781 2483
rect 775 2478 781 2479
rect 839 2483 845 2484
rect 839 2479 840 2483
rect 844 2482 845 2483
rect 863 2483 869 2484
rect 863 2482 864 2483
rect 844 2480 864 2482
rect 844 2479 845 2480
rect 839 2478 845 2479
rect 863 2479 864 2480
rect 868 2479 869 2483
rect 863 2478 869 2479
rect 951 2483 960 2484
rect 951 2479 952 2483
rect 959 2479 960 2483
rect 951 2478 960 2479
rect 1015 2483 1021 2484
rect 1015 2479 1016 2483
rect 1020 2482 1021 2483
rect 1039 2483 1045 2484
rect 1039 2482 1040 2483
rect 1020 2480 1040 2482
rect 1020 2479 1021 2480
rect 1015 2478 1021 2479
rect 1039 2479 1040 2480
rect 1044 2479 1045 2483
rect 1039 2478 1045 2479
rect 1103 2483 1109 2484
rect 1103 2479 1104 2483
rect 1108 2482 1109 2483
rect 1127 2483 1133 2484
rect 1127 2482 1128 2483
rect 1108 2480 1128 2482
rect 1108 2479 1109 2480
rect 1103 2478 1109 2479
rect 1127 2479 1128 2480
rect 1132 2479 1133 2483
rect 1127 2478 1133 2479
rect 1191 2483 1197 2484
rect 1191 2479 1192 2483
rect 1196 2482 1197 2483
rect 1215 2483 1221 2484
rect 1215 2482 1216 2483
rect 1196 2480 1216 2482
rect 1196 2479 1197 2480
rect 1191 2478 1197 2479
rect 1215 2479 1216 2480
rect 1220 2479 1221 2483
rect 1215 2478 1221 2479
rect 1279 2483 1285 2484
rect 1279 2479 1280 2483
rect 1284 2482 1285 2483
rect 1303 2483 1309 2484
rect 1303 2482 1304 2483
rect 1284 2480 1304 2482
rect 1284 2479 1285 2480
rect 1279 2478 1285 2479
rect 1303 2479 1304 2480
rect 1308 2479 1309 2483
rect 1303 2478 1309 2479
rect 2095 2483 2104 2484
rect 2095 2479 2096 2483
rect 2103 2479 2104 2483
rect 2095 2478 2104 2479
rect 2151 2483 2157 2484
rect 2151 2479 2152 2483
rect 2156 2482 2157 2483
rect 2191 2483 2197 2484
rect 2191 2482 2192 2483
rect 2156 2480 2192 2482
rect 2156 2479 2157 2480
rect 2151 2478 2157 2479
rect 2191 2479 2192 2480
rect 2196 2479 2197 2483
rect 2191 2478 2197 2479
rect 2247 2483 2253 2484
rect 2247 2479 2248 2483
rect 2252 2482 2253 2483
rect 2295 2483 2301 2484
rect 2295 2482 2296 2483
rect 2252 2480 2296 2482
rect 2252 2479 2253 2480
rect 2247 2478 2253 2479
rect 2295 2479 2296 2480
rect 2300 2479 2301 2483
rect 2295 2478 2301 2479
rect 2351 2483 2357 2484
rect 2351 2479 2352 2483
rect 2356 2482 2357 2483
rect 2415 2483 2421 2484
rect 2415 2482 2416 2483
rect 2356 2480 2416 2482
rect 2356 2479 2357 2480
rect 2351 2478 2357 2479
rect 2415 2479 2416 2480
rect 2420 2479 2421 2483
rect 2415 2478 2421 2479
rect 2551 2483 2557 2484
rect 2551 2479 2552 2483
rect 2556 2482 2557 2483
rect 2622 2483 2628 2484
rect 2622 2482 2623 2483
rect 2556 2480 2623 2482
rect 2556 2479 2557 2480
rect 2551 2478 2557 2479
rect 2622 2479 2623 2480
rect 2627 2479 2628 2483
rect 2622 2478 2628 2479
rect 2631 2483 2637 2484
rect 2631 2479 2632 2483
rect 2636 2482 2637 2483
rect 2711 2483 2717 2484
rect 2711 2482 2712 2483
rect 2636 2480 2712 2482
rect 2636 2479 2637 2480
rect 2631 2478 2637 2479
rect 2711 2479 2712 2480
rect 2716 2479 2717 2483
rect 2711 2478 2717 2479
rect 2775 2483 2781 2484
rect 2775 2479 2776 2483
rect 2780 2482 2781 2483
rect 2895 2483 2901 2484
rect 2895 2482 2896 2483
rect 2780 2480 2896 2482
rect 2780 2479 2781 2480
rect 2775 2478 2781 2479
rect 2895 2479 2896 2480
rect 2900 2479 2901 2483
rect 2895 2478 2901 2479
rect 2991 2483 2997 2484
rect 2991 2479 2992 2483
rect 2996 2482 2997 2483
rect 3095 2483 3101 2484
rect 3095 2482 3096 2483
rect 2996 2480 3096 2482
rect 2996 2479 2997 2480
rect 2991 2478 2997 2479
rect 3095 2479 3096 2480
rect 3100 2479 3101 2483
rect 3095 2478 3101 2479
rect 3302 2483 3309 2484
rect 3302 2479 3303 2483
rect 3308 2479 3309 2483
rect 3302 2478 3309 2479
rect 3471 2483 3477 2484
rect 3471 2479 3472 2483
rect 3476 2482 3477 2483
rect 3495 2483 3501 2484
rect 3495 2482 3496 2483
rect 3476 2480 3496 2482
rect 3476 2479 3477 2480
rect 3471 2478 3477 2479
rect 3495 2479 3496 2480
rect 3500 2479 3501 2483
rect 3495 2478 3501 2479
rect 2086 2473 2092 2474
rect 2086 2469 2087 2473
rect 2091 2469 2092 2473
rect 2086 2468 2092 2469
rect 2182 2473 2188 2474
rect 2182 2469 2183 2473
rect 2187 2469 2188 2473
rect 2182 2468 2188 2469
rect 2286 2473 2292 2474
rect 2286 2469 2287 2473
rect 2291 2469 2292 2473
rect 2286 2468 2292 2469
rect 2406 2473 2412 2474
rect 2406 2469 2407 2473
rect 2411 2469 2412 2473
rect 2406 2468 2412 2469
rect 2542 2473 2548 2474
rect 2542 2469 2543 2473
rect 2547 2469 2548 2473
rect 2542 2468 2548 2469
rect 2702 2473 2708 2474
rect 2702 2469 2703 2473
rect 2707 2469 2708 2473
rect 2702 2468 2708 2469
rect 2886 2473 2892 2474
rect 2886 2469 2887 2473
rect 2891 2469 2892 2473
rect 2886 2468 2892 2469
rect 3086 2473 3092 2474
rect 3086 2469 3087 2473
rect 3091 2469 3092 2473
rect 3086 2468 3092 2469
rect 3294 2473 3300 2474
rect 3294 2469 3295 2473
rect 3299 2469 3300 2473
rect 3294 2468 3300 2469
rect 3486 2473 3492 2474
rect 3486 2469 3487 2473
rect 3491 2469 3492 2473
rect 3486 2468 3492 2469
rect 367 2467 373 2468
rect 367 2463 368 2467
rect 372 2466 373 2467
rect 423 2467 429 2468
rect 372 2464 418 2466
rect 372 2463 373 2464
rect 367 2462 373 2463
rect 414 2463 420 2464
rect 414 2459 415 2463
rect 419 2459 420 2463
rect 423 2463 424 2467
rect 428 2466 429 2467
rect 479 2467 485 2468
rect 479 2466 480 2467
rect 428 2464 480 2466
rect 428 2463 429 2464
rect 423 2462 429 2463
rect 479 2463 480 2464
rect 484 2463 485 2467
rect 479 2462 485 2463
rect 599 2467 605 2468
rect 599 2463 600 2467
rect 604 2466 605 2467
rect 663 2467 669 2468
rect 663 2466 664 2467
rect 604 2464 664 2466
rect 604 2463 605 2464
rect 599 2462 605 2463
rect 663 2463 664 2464
rect 668 2463 669 2467
rect 663 2462 669 2463
rect 727 2467 736 2468
rect 727 2463 728 2467
rect 735 2463 736 2467
rect 727 2462 736 2463
rect 838 2467 844 2468
rect 838 2463 839 2467
rect 843 2466 844 2467
rect 855 2467 861 2468
rect 855 2466 856 2467
rect 843 2464 856 2466
rect 843 2463 844 2464
rect 838 2462 844 2463
rect 855 2463 856 2464
rect 860 2463 861 2467
rect 855 2462 861 2463
rect 975 2467 984 2468
rect 975 2463 976 2467
rect 983 2463 984 2467
rect 975 2462 984 2463
rect 1031 2467 1037 2468
rect 1031 2463 1032 2467
rect 1036 2466 1037 2467
rect 1095 2467 1101 2468
rect 1095 2466 1096 2467
rect 1036 2464 1096 2466
rect 1036 2463 1037 2464
rect 1031 2462 1037 2463
rect 1095 2463 1096 2464
rect 1100 2463 1101 2467
rect 1095 2462 1101 2463
rect 1146 2467 1152 2468
rect 1146 2463 1147 2467
rect 1151 2466 1152 2467
rect 1215 2467 1221 2468
rect 1215 2466 1216 2467
rect 1151 2464 1216 2466
rect 1151 2463 1152 2464
rect 1146 2462 1152 2463
rect 1215 2463 1216 2464
rect 1220 2463 1221 2467
rect 1215 2462 1221 2463
rect 1279 2467 1285 2468
rect 1279 2463 1280 2467
rect 1284 2466 1285 2467
rect 1343 2467 1349 2468
rect 1343 2466 1344 2467
rect 1284 2464 1344 2466
rect 1284 2463 1285 2464
rect 1279 2462 1285 2463
rect 1343 2463 1344 2464
rect 1348 2463 1349 2467
rect 1343 2462 1349 2463
rect 1407 2467 1413 2468
rect 1407 2463 1408 2467
rect 1412 2466 1413 2467
rect 1471 2467 1477 2468
rect 1471 2466 1472 2467
rect 1412 2464 1472 2466
rect 1412 2463 1413 2464
rect 1407 2462 1413 2463
rect 1471 2463 1472 2464
rect 1476 2463 1477 2467
rect 1471 2462 1477 2463
rect 414 2458 420 2459
rect 1862 2460 1868 2461
rect 3574 2460 3580 2461
rect 358 2457 364 2458
rect 358 2453 359 2457
rect 363 2453 364 2457
rect 358 2452 364 2453
rect 470 2457 476 2458
rect 470 2453 471 2457
rect 475 2453 476 2457
rect 470 2452 476 2453
rect 590 2457 596 2458
rect 590 2453 591 2457
rect 595 2453 596 2457
rect 590 2452 596 2453
rect 718 2457 724 2458
rect 718 2453 719 2457
rect 723 2453 724 2457
rect 718 2452 724 2453
rect 846 2457 852 2458
rect 846 2453 847 2457
rect 851 2453 852 2457
rect 846 2452 852 2453
rect 966 2457 972 2458
rect 966 2453 967 2457
rect 971 2453 972 2457
rect 966 2452 972 2453
rect 1086 2457 1092 2458
rect 1086 2453 1087 2457
rect 1091 2453 1092 2457
rect 1086 2452 1092 2453
rect 1206 2457 1212 2458
rect 1206 2453 1207 2457
rect 1211 2453 1212 2457
rect 1206 2452 1212 2453
rect 1334 2457 1340 2458
rect 1334 2453 1335 2457
rect 1339 2453 1340 2457
rect 1334 2452 1340 2453
rect 1462 2457 1468 2458
rect 1462 2453 1463 2457
rect 1467 2453 1468 2457
rect 1862 2456 1863 2460
rect 1867 2456 1868 2460
rect 2151 2459 2157 2460
rect 2151 2458 2152 2459
rect 2141 2456 2152 2458
rect 1862 2455 1868 2456
rect 2151 2455 2152 2456
rect 2156 2455 2157 2459
rect 2247 2459 2253 2460
rect 2247 2458 2248 2459
rect 2237 2456 2248 2458
rect 2151 2454 2157 2455
rect 2247 2455 2248 2456
rect 2252 2455 2253 2459
rect 2351 2459 2357 2460
rect 2351 2458 2352 2459
rect 2341 2456 2352 2458
rect 2247 2454 2253 2455
rect 2351 2455 2352 2456
rect 2356 2455 2357 2459
rect 2631 2459 2637 2460
rect 2631 2458 2632 2459
rect 2597 2456 2632 2458
rect 2351 2454 2357 2455
rect 2359 2455 2365 2456
rect 1462 2452 1468 2453
rect 2359 2451 2360 2455
rect 2364 2454 2365 2455
rect 2631 2455 2632 2456
rect 2636 2455 2637 2459
rect 2775 2459 2781 2460
rect 2775 2458 2776 2459
rect 2757 2456 2776 2458
rect 2631 2454 2637 2455
rect 2775 2455 2776 2456
rect 2780 2455 2781 2459
rect 2991 2459 2997 2460
rect 2991 2458 2992 2459
rect 2941 2456 2992 2458
rect 2775 2454 2781 2455
rect 2991 2455 2992 2456
rect 2996 2455 2997 2459
rect 3354 2459 3360 2460
rect 3354 2458 3355 2459
rect 3349 2456 3355 2458
rect 2991 2454 2997 2455
rect 3354 2455 3355 2456
rect 3359 2455 3360 2459
rect 3574 2456 3575 2460
rect 3579 2456 3580 2460
rect 3574 2455 3580 2456
rect 3354 2454 3360 2455
rect 2364 2452 2425 2454
rect 2364 2451 2365 2452
rect 2359 2450 2365 2451
rect 110 2444 116 2445
rect 1822 2444 1828 2445
rect 110 2440 111 2444
rect 115 2440 116 2444
rect 423 2443 429 2444
rect 423 2442 424 2443
rect 413 2440 424 2442
rect 110 2439 116 2440
rect 423 2439 424 2440
rect 428 2439 429 2443
rect 1031 2443 1037 2444
rect 1031 2442 1032 2443
rect 1021 2440 1032 2442
rect 423 2438 429 2439
rect 582 2439 588 2440
rect 582 2435 583 2439
rect 587 2438 588 2439
rect 663 2439 669 2440
rect 587 2436 609 2438
rect 587 2435 588 2436
rect 582 2434 588 2435
rect 663 2435 664 2439
rect 668 2438 669 2439
rect 786 2439 792 2440
rect 668 2436 737 2438
rect 668 2435 669 2436
rect 663 2434 669 2435
rect 786 2435 787 2439
rect 791 2438 792 2439
rect 1031 2439 1032 2440
rect 1036 2439 1037 2443
rect 1146 2443 1152 2444
rect 1146 2442 1147 2443
rect 1141 2440 1147 2442
rect 1031 2438 1037 2439
rect 1146 2439 1147 2440
rect 1151 2439 1152 2443
rect 1279 2443 1285 2444
rect 1279 2442 1280 2443
rect 1261 2440 1280 2442
rect 1146 2438 1152 2439
rect 1279 2439 1280 2440
rect 1284 2439 1285 2443
rect 1407 2443 1413 2444
rect 1407 2442 1408 2443
rect 1389 2440 1408 2442
rect 1279 2438 1285 2439
rect 1407 2439 1408 2440
rect 1412 2439 1413 2443
rect 1822 2440 1823 2444
rect 1827 2440 1828 2444
rect 1822 2439 1828 2440
rect 1862 2443 1868 2444
rect 1862 2439 1863 2443
rect 1867 2439 1868 2443
rect 1407 2438 1413 2439
rect 1862 2438 1868 2439
rect 2954 2443 2960 2444
rect 2954 2439 2955 2443
rect 2959 2442 2960 2443
rect 3574 2443 3580 2444
rect 2959 2440 3097 2442
rect 2959 2439 2960 2440
rect 2954 2438 2960 2439
rect 3574 2439 3575 2443
rect 3579 2439 3580 2443
rect 3574 2438 3580 2439
rect 791 2436 865 2438
rect 791 2435 792 2436
rect 786 2434 792 2435
rect 2078 2433 2084 2434
rect 2078 2429 2079 2433
rect 2083 2429 2084 2433
rect 2078 2428 2084 2429
rect 2174 2433 2180 2434
rect 2174 2429 2175 2433
rect 2179 2429 2180 2433
rect 2174 2428 2180 2429
rect 2278 2433 2284 2434
rect 2278 2429 2279 2433
rect 2283 2429 2284 2433
rect 2278 2428 2284 2429
rect 2398 2433 2404 2434
rect 2398 2429 2399 2433
rect 2403 2429 2404 2433
rect 2398 2428 2404 2429
rect 2534 2433 2540 2434
rect 2534 2429 2535 2433
rect 2539 2429 2540 2433
rect 2534 2428 2540 2429
rect 2694 2433 2700 2434
rect 2694 2429 2695 2433
rect 2699 2429 2700 2433
rect 2694 2428 2700 2429
rect 2878 2433 2884 2434
rect 2878 2429 2879 2433
rect 2883 2429 2884 2433
rect 2878 2428 2884 2429
rect 3078 2433 3084 2434
rect 3078 2429 3079 2433
rect 3083 2429 3084 2433
rect 3078 2428 3084 2429
rect 3286 2433 3292 2434
rect 3286 2429 3287 2433
rect 3291 2429 3292 2433
rect 3286 2428 3292 2429
rect 3478 2433 3484 2434
rect 3478 2429 3479 2433
rect 3483 2429 3484 2433
rect 3478 2428 3484 2429
rect 110 2427 116 2428
rect 110 2423 111 2427
rect 115 2423 116 2427
rect 110 2422 116 2423
rect 1402 2427 1408 2428
rect 1402 2423 1403 2427
rect 1407 2426 1408 2427
rect 1822 2427 1828 2428
rect 1407 2424 1473 2426
rect 1407 2423 1408 2424
rect 1402 2422 1408 2423
rect 1822 2423 1823 2427
rect 1827 2423 1828 2427
rect 1822 2422 1828 2423
rect 3498 2427 3504 2428
rect 3498 2423 3499 2427
rect 3503 2426 3504 2427
rect 3527 2427 3533 2428
rect 3527 2426 3528 2427
rect 3503 2424 3528 2426
rect 3503 2423 3504 2424
rect 3498 2422 3504 2423
rect 3527 2423 3528 2424
rect 3532 2423 3533 2427
rect 3527 2422 3533 2423
rect 2610 2419 2616 2420
rect 350 2417 356 2418
rect 350 2413 351 2417
rect 355 2413 356 2417
rect 350 2412 356 2413
rect 462 2417 468 2418
rect 462 2413 463 2417
rect 467 2413 468 2417
rect 462 2412 468 2413
rect 582 2417 588 2418
rect 582 2413 583 2417
rect 587 2413 588 2417
rect 582 2412 588 2413
rect 710 2417 716 2418
rect 710 2413 711 2417
rect 715 2413 716 2417
rect 710 2412 716 2413
rect 838 2417 844 2418
rect 838 2413 839 2417
rect 843 2413 844 2417
rect 838 2412 844 2413
rect 958 2417 964 2418
rect 958 2413 959 2417
rect 963 2413 964 2417
rect 958 2412 964 2413
rect 1078 2417 1084 2418
rect 1078 2413 1079 2417
rect 1083 2413 1084 2417
rect 1078 2412 1084 2413
rect 1198 2417 1204 2418
rect 1198 2413 1199 2417
rect 1203 2413 1204 2417
rect 1198 2412 1204 2413
rect 1326 2417 1332 2418
rect 1326 2413 1327 2417
rect 1331 2413 1332 2417
rect 1326 2412 1332 2413
rect 1454 2417 1460 2418
rect 1454 2413 1455 2417
rect 1459 2413 1460 2417
rect 2610 2415 2611 2419
rect 2615 2418 2616 2419
rect 2954 2419 2960 2420
rect 2954 2418 2955 2419
rect 2615 2416 2955 2418
rect 2615 2415 2616 2416
rect 2610 2414 2616 2415
rect 2954 2415 2955 2416
rect 2959 2415 2960 2419
rect 2954 2414 2960 2415
rect 1454 2412 1460 2413
rect 490 2411 496 2412
rect 490 2407 491 2411
rect 495 2410 496 2411
rect 511 2411 517 2412
rect 511 2410 512 2411
rect 495 2408 512 2410
rect 495 2407 496 2408
rect 490 2406 496 2407
rect 511 2407 512 2408
rect 516 2407 517 2411
rect 511 2406 517 2407
rect 1950 2407 1956 2408
rect 1950 2403 1951 2407
rect 1955 2403 1956 2407
rect 1950 2402 1956 2403
rect 2062 2407 2068 2408
rect 2062 2403 2063 2407
rect 2067 2403 2068 2407
rect 2062 2402 2068 2403
rect 2182 2407 2188 2408
rect 2182 2403 2183 2407
rect 2187 2403 2188 2407
rect 2182 2402 2188 2403
rect 2310 2407 2316 2408
rect 2310 2403 2311 2407
rect 2315 2403 2316 2407
rect 2310 2402 2316 2403
rect 2446 2407 2452 2408
rect 2446 2403 2447 2407
rect 2451 2403 2452 2407
rect 2446 2402 2452 2403
rect 2590 2407 2596 2408
rect 2590 2403 2591 2407
rect 2595 2403 2596 2407
rect 2590 2402 2596 2403
rect 2750 2407 2756 2408
rect 2750 2403 2751 2407
rect 2755 2403 2756 2407
rect 2750 2402 2756 2403
rect 2926 2407 2932 2408
rect 2926 2403 2927 2407
rect 2931 2403 2932 2407
rect 2926 2402 2932 2403
rect 3110 2407 3116 2408
rect 3110 2403 3111 2407
rect 3115 2403 3116 2407
rect 3110 2402 3116 2403
rect 3302 2407 3308 2408
rect 3302 2403 3303 2407
rect 3307 2403 3308 2407
rect 3302 2402 3308 2403
rect 3478 2407 3484 2408
rect 3478 2403 3479 2407
rect 3483 2403 3484 2407
rect 3478 2402 3484 2403
rect 2378 2399 2384 2400
rect 1862 2397 1868 2398
rect 1862 2393 1863 2397
rect 1867 2393 1868 2397
rect 2378 2395 2379 2399
rect 2383 2398 2384 2399
rect 3018 2399 3024 2400
rect 2383 2396 2465 2398
rect 2383 2395 2384 2396
rect 2378 2394 2384 2395
rect 3018 2395 3019 2399
rect 3023 2398 3024 2399
rect 3294 2399 3300 2400
rect 3023 2396 3129 2398
rect 3023 2395 3024 2396
rect 3018 2394 3024 2395
rect 3294 2395 3295 2399
rect 3299 2398 3300 2399
rect 3299 2396 3321 2398
rect 3574 2397 3580 2398
rect 3299 2395 3300 2396
rect 3294 2394 3300 2395
rect 1862 2392 1868 2393
rect 3574 2393 3575 2397
rect 3579 2393 3580 2397
rect 3574 2392 3580 2393
rect 134 2391 140 2392
rect 134 2387 135 2391
rect 139 2387 140 2391
rect 134 2386 140 2387
rect 286 2391 292 2392
rect 286 2387 287 2391
rect 291 2387 292 2391
rect 286 2386 292 2387
rect 470 2391 476 2392
rect 470 2387 471 2391
rect 475 2387 476 2391
rect 470 2386 476 2387
rect 662 2391 668 2392
rect 662 2387 663 2391
rect 667 2387 668 2391
rect 662 2386 668 2387
rect 846 2391 852 2392
rect 846 2387 847 2391
rect 851 2387 852 2391
rect 846 2386 852 2387
rect 1030 2391 1036 2392
rect 1030 2387 1031 2391
rect 1035 2387 1036 2391
rect 1030 2386 1036 2387
rect 1206 2391 1212 2392
rect 1206 2387 1207 2391
rect 1211 2387 1212 2391
rect 1206 2386 1212 2387
rect 1374 2391 1380 2392
rect 1374 2387 1375 2391
rect 1379 2387 1380 2391
rect 1374 2386 1380 2387
rect 1542 2391 1548 2392
rect 1542 2387 1543 2391
rect 1547 2387 1548 2391
rect 1542 2386 1548 2387
rect 1710 2391 1716 2392
rect 1710 2387 1711 2391
rect 1715 2387 1716 2391
rect 1710 2386 1716 2387
rect 202 2383 208 2384
rect 110 2381 116 2382
rect 110 2377 111 2381
rect 115 2377 116 2381
rect 202 2379 203 2383
rect 207 2382 208 2383
rect 730 2383 736 2384
rect 730 2382 731 2383
rect 207 2380 305 2382
rect 721 2380 731 2382
rect 207 2379 208 2380
rect 202 2378 208 2379
rect 730 2379 731 2380
rect 735 2379 736 2383
rect 2055 2383 2061 2384
rect 2055 2382 2056 2383
rect 730 2378 736 2379
rect 1822 2381 1828 2382
rect 110 2376 116 2377
rect 1822 2377 1823 2381
rect 1827 2377 1828 2381
rect 1822 2376 1828 2377
rect 1862 2380 1868 2381
rect 2013 2380 2056 2382
rect 1862 2376 1863 2380
rect 1867 2376 1868 2380
rect 2055 2379 2056 2380
rect 2060 2379 2061 2383
rect 2175 2383 2181 2384
rect 2175 2382 2176 2383
rect 2125 2380 2176 2382
rect 2055 2378 2061 2379
rect 2175 2379 2176 2380
rect 2180 2379 2181 2383
rect 2303 2383 2309 2384
rect 2303 2382 2304 2383
rect 2245 2380 2304 2382
rect 2175 2378 2181 2379
rect 2303 2379 2304 2380
rect 2308 2379 2309 2383
rect 2439 2383 2445 2384
rect 2439 2382 2440 2383
rect 2373 2380 2440 2382
rect 2303 2378 2309 2379
rect 2439 2379 2440 2380
rect 2444 2379 2445 2383
rect 2743 2383 2749 2384
rect 2743 2382 2744 2383
rect 2653 2380 2744 2382
rect 2439 2378 2445 2379
rect 2743 2379 2744 2380
rect 2748 2379 2749 2383
rect 2919 2383 2925 2384
rect 2919 2382 2920 2383
rect 2813 2380 2920 2382
rect 2743 2378 2749 2379
rect 2919 2379 2920 2380
rect 2924 2379 2925 2383
rect 3103 2383 3109 2384
rect 3103 2382 3104 2383
rect 2989 2380 3104 2382
rect 2919 2378 2925 2379
rect 3103 2379 3104 2380
rect 3108 2379 3109 2383
rect 3103 2378 3109 2379
rect 3471 2383 3477 2384
rect 3471 2379 3472 2383
rect 3476 2382 3477 2383
rect 3476 2380 3505 2382
rect 3574 2380 3580 2381
rect 3476 2379 3477 2380
rect 3471 2378 3477 2379
rect 1862 2375 1868 2376
rect 3574 2376 3575 2380
rect 3579 2376 3580 2380
rect 3574 2375 3580 2376
rect 279 2367 285 2368
rect 279 2366 280 2367
rect 110 2364 116 2365
rect 197 2364 280 2366
rect 110 2360 111 2364
rect 115 2360 116 2364
rect 279 2363 280 2364
rect 284 2363 285 2367
rect 279 2362 285 2363
rect 362 2367 368 2368
rect 362 2363 363 2367
rect 367 2366 368 2367
rect 730 2367 736 2368
rect 367 2364 497 2366
rect 367 2363 368 2364
rect 362 2362 368 2363
rect 730 2363 731 2367
rect 735 2366 736 2367
rect 1199 2367 1205 2368
rect 1199 2366 1200 2367
rect 735 2364 873 2366
rect 1093 2364 1200 2366
rect 735 2363 736 2364
rect 730 2362 736 2363
rect 1199 2363 1200 2364
rect 1204 2363 1205 2367
rect 1367 2367 1373 2368
rect 1367 2366 1368 2367
rect 1269 2364 1368 2366
rect 1199 2362 1205 2363
rect 1367 2363 1368 2364
rect 1372 2363 1373 2367
rect 1535 2367 1541 2368
rect 1535 2366 1536 2367
rect 1437 2364 1536 2366
rect 1367 2362 1373 2363
rect 1535 2363 1536 2364
rect 1540 2363 1541 2367
rect 1703 2367 1709 2368
rect 1703 2366 1704 2367
rect 1605 2364 1704 2366
rect 1535 2362 1541 2363
rect 1703 2363 1704 2364
rect 1708 2363 1709 2367
rect 1778 2367 1784 2368
rect 1778 2366 1779 2367
rect 1773 2364 1779 2366
rect 1703 2362 1709 2363
rect 1778 2363 1779 2364
rect 1783 2363 1784 2367
rect 1958 2367 1964 2368
rect 1778 2362 1784 2363
rect 1822 2364 1828 2365
rect 110 2359 116 2360
rect 1822 2360 1823 2364
rect 1827 2360 1828 2364
rect 1958 2363 1959 2367
rect 1963 2363 1964 2367
rect 1958 2362 1964 2363
rect 2070 2367 2076 2368
rect 2070 2363 2071 2367
rect 2075 2363 2076 2367
rect 2070 2362 2076 2363
rect 2190 2367 2196 2368
rect 2190 2363 2191 2367
rect 2195 2363 2196 2367
rect 2190 2362 2196 2363
rect 2318 2367 2324 2368
rect 2318 2363 2319 2367
rect 2323 2363 2324 2367
rect 2318 2362 2324 2363
rect 2454 2367 2460 2368
rect 2454 2363 2455 2367
rect 2459 2363 2460 2367
rect 2454 2362 2460 2363
rect 2598 2367 2604 2368
rect 2598 2363 2599 2367
rect 2603 2363 2604 2367
rect 2598 2362 2604 2363
rect 2758 2367 2764 2368
rect 2758 2363 2759 2367
rect 2763 2363 2764 2367
rect 2758 2362 2764 2363
rect 2934 2367 2940 2368
rect 2934 2363 2935 2367
rect 2939 2363 2940 2367
rect 2934 2362 2940 2363
rect 3118 2367 3124 2368
rect 3118 2363 3119 2367
rect 3123 2363 3124 2367
rect 3118 2362 3124 2363
rect 3310 2367 3316 2368
rect 3310 2363 3311 2367
rect 3315 2363 3316 2367
rect 3310 2362 3316 2363
rect 3486 2367 3492 2368
rect 3486 2363 3487 2367
rect 3491 2363 3492 2367
rect 3486 2362 3492 2363
rect 1822 2359 1828 2360
rect 1967 2355 1973 2356
rect 142 2351 148 2352
rect 142 2347 143 2351
rect 147 2347 148 2351
rect 142 2346 148 2347
rect 294 2351 300 2352
rect 294 2347 295 2351
rect 299 2347 300 2351
rect 294 2346 300 2347
rect 478 2351 484 2352
rect 478 2347 479 2351
rect 483 2347 484 2351
rect 478 2346 484 2347
rect 670 2351 676 2352
rect 670 2347 671 2351
rect 675 2347 676 2351
rect 670 2346 676 2347
rect 854 2351 860 2352
rect 854 2347 855 2351
rect 859 2347 860 2351
rect 854 2346 860 2347
rect 1038 2351 1044 2352
rect 1038 2347 1039 2351
rect 1043 2347 1044 2351
rect 1038 2346 1044 2347
rect 1214 2351 1220 2352
rect 1214 2347 1215 2351
rect 1219 2347 1220 2351
rect 1214 2346 1220 2347
rect 1382 2351 1388 2352
rect 1382 2347 1383 2351
rect 1387 2347 1388 2351
rect 1382 2346 1388 2347
rect 1550 2351 1556 2352
rect 1550 2347 1551 2351
rect 1555 2347 1556 2351
rect 1550 2346 1556 2347
rect 1718 2351 1724 2352
rect 1718 2347 1719 2351
rect 1723 2347 1724 2351
rect 1967 2351 1968 2355
rect 1972 2354 1973 2355
rect 2046 2355 2052 2356
rect 2046 2354 2047 2355
rect 1972 2352 2047 2354
rect 1972 2351 1973 2352
rect 1967 2350 1973 2351
rect 2046 2351 2047 2352
rect 2051 2351 2052 2355
rect 2046 2350 2052 2351
rect 2055 2355 2061 2356
rect 2055 2351 2056 2355
rect 2060 2354 2061 2355
rect 2079 2355 2085 2356
rect 2079 2354 2080 2355
rect 2060 2352 2080 2354
rect 2060 2351 2061 2352
rect 2055 2350 2061 2351
rect 2079 2351 2080 2352
rect 2084 2351 2085 2355
rect 2079 2350 2085 2351
rect 2175 2355 2181 2356
rect 2175 2351 2176 2355
rect 2180 2354 2181 2355
rect 2199 2355 2205 2356
rect 2199 2354 2200 2355
rect 2180 2352 2200 2354
rect 2180 2351 2181 2352
rect 2175 2350 2181 2351
rect 2199 2351 2200 2352
rect 2204 2351 2205 2355
rect 2199 2350 2205 2351
rect 2303 2355 2309 2356
rect 2303 2351 2304 2355
rect 2308 2354 2309 2355
rect 2327 2355 2333 2356
rect 2327 2354 2328 2355
rect 2308 2352 2328 2354
rect 2308 2351 2309 2352
rect 2303 2350 2309 2351
rect 2327 2351 2328 2352
rect 2332 2351 2333 2355
rect 2327 2350 2333 2351
rect 2439 2355 2445 2356
rect 2439 2351 2440 2355
rect 2444 2354 2445 2355
rect 2463 2355 2469 2356
rect 2463 2354 2464 2355
rect 2444 2352 2464 2354
rect 2444 2351 2445 2352
rect 2439 2350 2445 2351
rect 2463 2351 2464 2352
rect 2468 2351 2469 2355
rect 2463 2350 2469 2351
rect 2607 2355 2616 2356
rect 2607 2351 2608 2355
rect 2615 2351 2616 2355
rect 2607 2350 2616 2351
rect 2743 2355 2749 2356
rect 2743 2351 2744 2355
rect 2748 2354 2749 2355
rect 2767 2355 2773 2356
rect 2767 2354 2768 2355
rect 2748 2352 2768 2354
rect 2748 2351 2749 2352
rect 2743 2350 2749 2351
rect 2767 2351 2768 2352
rect 2772 2351 2773 2355
rect 2767 2350 2773 2351
rect 2919 2355 2925 2356
rect 2919 2351 2920 2355
rect 2924 2354 2925 2355
rect 2943 2355 2949 2356
rect 2943 2354 2944 2355
rect 2924 2352 2944 2354
rect 2924 2351 2925 2352
rect 2919 2350 2925 2351
rect 2943 2351 2944 2352
rect 2948 2351 2949 2355
rect 2943 2350 2949 2351
rect 3103 2355 3109 2356
rect 3103 2351 3104 2355
rect 3108 2354 3109 2355
rect 3127 2355 3133 2356
rect 3127 2354 3128 2355
rect 3108 2352 3128 2354
rect 3108 2351 3109 2352
rect 3103 2350 3109 2351
rect 3127 2351 3128 2352
rect 3132 2351 3133 2355
rect 3127 2350 3133 2351
rect 3319 2355 3325 2356
rect 3319 2351 3320 2355
rect 3324 2354 3325 2355
rect 3359 2355 3365 2356
rect 3359 2354 3360 2355
rect 3324 2352 3360 2354
rect 3324 2351 3325 2352
rect 3319 2350 3325 2351
rect 3359 2351 3360 2352
rect 3364 2351 3365 2355
rect 3359 2350 3365 2351
rect 3495 2355 3504 2356
rect 3495 2351 3496 2355
rect 3503 2351 3504 2355
rect 3495 2350 3504 2351
rect 1718 2346 1724 2347
rect 3018 2343 3024 2344
rect 3018 2342 3019 2343
rect 2732 2340 3019 2342
rect 151 2339 157 2340
rect 151 2335 152 2339
rect 156 2338 157 2339
rect 202 2339 208 2340
rect 202 2338 203 2339
rect 156 2336 203 2338
rect 156 2335 157 2336
rect 151 2334 157 2335
rect 202 2335 203 2336
rect 207 2335 208 2339
rect 202 2334 208 2335
rect 303 2339 309 2340
rect 303 2335 304 2339
rect 308 2338 309 2339
rect 362 2339 368 2340
rect 362 2338 363 2339
rect 308 2336 363 2338
rect 308 2335 309 2336
rect 303 2334 309 2335
rect 362 2335 363 2336
rect 367 2335 368 2339
rect 362 2334 368 2335
rect 487 2339 496 2340
rect 487 2335 488 2339
rect 495 2335 496 2339
rect 487 2334 496 2335
rect 679 2339 685 2340
rect 679 2335 680 2339
rect 684 2338 685 2339
rect 730 2339 736 2340
rect 730 2338 731 2339
rect 684 2336 731 2338
rect 684 2335 685 2336
rect 679 2334 685 2335
rect 730 2335 731 2336
rect 735 2335 736 2339
rect 730 2334 736 2335
rect 846 2339 852 2340
rect 846 2335 847 2339
rect 851 2338 852 2339
rect 863 2339 869 2340
rect 863 2338 864 2339
rect 851 2336 864 2338
rect 851 2335 852 2336
rect 846 2334 852 2335
rect 863 2335 864 2336
rect 868 2335 869 2339
rect 863 2334 869 2335
rect 1047 2339 1053 2340
rect 1047 2335 1048 2339
rect 1052 2338 1053 2339
rect 1094 2339 1100 2340
rect 1094 2338 1095 2339
rect 1052 2336 1095 2338
rect 1052 2335 1053 2336
rect 1047 2334 1053 2335
rect 1094 2335 1095 2336
rect 1099 2335 1100 2339
rect 1094 2334 1100 2335
rect 1199 2339 1205 2340
rect 1199 2335 1200 2339
rect 1204 2338 1205 2339
rect 1223 2339 1229 2340
rect 1223 2338 1224 2339
rect 1204 2336 1224 2338
rect 1204 2335 1205 2336
rect 1199 2334 1205 2335
rect 1223 2335 1224 2336
rect 1228 2335 1229 2339
rect 1223 2334 1229 2335
rect 1367 2339 1373 2340
rect 1367 2335 1368 2339
rect 1372 2338 1373 2339
rect 1391 2339 1397 2340
rect 1391 2338 1392 2339
rect 1372 2336 1392 2338
rect 1372 2335 1373 2336
rect 1367 2334 1373 2335
rect 1391 2335 1392 2336
rect 1396 2335 1397 2339
rect 1391 2334 1397 2335
rect 1535 2339 1541 2340
rect 1535 2335 1536 2339
rect 1540 2338 1541 2339
rect 1559 2339 1565 2340
rect 1559 2338 1560 2339
rect 1540 2336 1560 2338
rect 1540 2335 1541 2336
rect 1535 2334 1541 2335
rect 1559 2335 1560 2336
rect 1564 2335 1565 2339
rect 1559 2334 1565 2335
rect 1703 2339 1709 2340
rect 1703 2335 1704 2339
rect 1708 2338 1709 2339
rect 1727 2339 1733 2340
rect 1727 2338 1728 2339
rect 1708 2336 1728 2338
rect 1708 2335 1709 2336
rect 1703 2334 1709 2335
rect 1727 2335 1728 2336
rect 1732 2335 1733 2339
rect 1727 2334 1733 2335
rect 1903 2335 1909 2336
rect 1903 2331 1904 2335
rect 1908 2334 1909 2335
rect 1950 2335 1956 2336
rect 1950 2334 1951 2335
rect 1908 2332 1951 2334
rect 1908 2331 1909 2332
rect 1903 2330 1909 2331
rect 1950 2331 1951 2332
rect 1955 2331 1956 2335
rect 1950 2330 1956 2331
rect 1959 2335 1965 2336
rect 1959 2331 1960 2335
rect 1964 2334 1965 2335
rect 2015 2335 2021 2336
rect 2015 2334 2016 2335
rect 1964 2332 2016 2334
rect 1964 2331 1965 2332
rect 1959 2330 1965 2331
rect 2015 2331 2016 2332
rect 2020 2331 2021 2335
rect 2015 2330 2021 2331
rect 2087 2335 2093 2336
rect 2087 2331 2088 2335
rect 2092 2334 2093 2335
rect 2167 2335 2173 2336
rect 2167 2334 2168 2335
rect 2092 2332 2168 2334
rect 2092 2331 2093 2332
rect 2087 2330 2093 2331
rect 2167 2331 2168 2332
rect 2172 2331 2173 2335
rect 2167 2330 2173 2331
rect 2239 2335 2245 2336
rect 2239 2331 2240 2335
rect 2244 2334 2245 2335
rect 2319 2335 2325 2336
rect 2319 2334 2320 2335
rect 2244 2332 2320 2334
rect 2244 2331 2245 2332
rect 2239 2330 2245 2331
rect 2319 2331 2320 2332
rect 2324 2331 2325 2335
rect 2319 2330 2325 2331
rect 2391 2335 2397 2336
rect 2391 2331 2392 2335
rect 2396 2334 2397 2335
rect 2471 2335 2477 2336
rect 2471 2334 2472 2335
rect 2396 2332 2472 2334
rect 2396 2331 2397 2332
rect 2391 2330 2397 2331
rect 2471 2331 2472 2332
rect 2476 2331 2477 2335
rect 2471 2330 2477 2331
rect 2623 2335 2629 2336
rect 2623 2331 2624 2335
rect 2628 2334 2629 2335
rect 2732 2334 2734 2340
rect 3018 2339 3019 2340
rect 3023 2339 3024 2343
rect 3018 2338 3024 2339
rect 2628 2332 2734 2334
rect 2743 2335 2749 2336
rect 2628 2331 2629 2332
rect 2623 2330 2629 2331
rect 2743 2331 2744 2335
rect 2748 2334 2749 2335
rect 2783 2335 2789 2336
rect 2783 2334 2784 2335
rect 2748 2332 2784 2334
rect 2748 2331 2749 2332
rect 2743 2330 2749 2331
rect 2783 2331 2784 2332
rect 2788 2331 2789 2335
rect 2783 2330 2789 2331
rect 2874 2335 2880 2336
rect 2874 2331 2875 2335
rect 2879 2334 2880 2335
rect 2951 2335 2957 2336
rect 2951 2334 2952 2335
rect 2879 2332 2952 2334
rect 2879 2331 2880 2332
rect 2874 2330 2880 2331
rect 2951 2331 2952 2332
rect 2956 2331 2957 2335
rect 2951 2330 2957 2331
rect 3031 2335 3037 2336
rect 3031 2331 3032 2335
rect 3036 2334 3037 2335
rect 3119 2335 3125 2336
rect 3119 2334 3120 2335
rect 3036 2332 3120 2334
rect 3036 2331 3037 2332
rect 3031 2330 3037 2331
rect 3119 2331 3120 2332
rect 3124 2331 3125 2335
rect 3119 2330 3125 2331
rect 3207 2335 3213 2336
rect 3207 2331 3208 2335
rect 3212 2334 3213 2335
rect 3295 2335 3301 2336
rect 3295 2334 3296 2335
rect 3212 2332 3296 2334
rect 3212 2331 3213 2332
rect 3207 2330 3213 2331
rect 3295 2331 3296 2332
rect 3300 2331 3301 2335
rect 3295 2330 3301 2331
rect 3471 2335 3477 2336
rect 3471 2331 3472 2335
rect 3476 2334 3477 2335
rect 3479 2335 3485 2336
rect 3479 2334 3480 2335
rect 3476 2332 3480 2334
rect 3476 2331 3477 2332
rect 3471 2330 3477 2331
rect 3479 2331 3480 2332
rect 3484 2331 3485 2335
rect 3479 2330 3485 2331
rect 1894 2325 1900 2326
rect 151 2323 157 2324
rect 151 2319 152 2323
rect 156 2322 157 2323
rect 226 2323 232 2324
rect 226 2322 227 2323
rect 156 2320 227 2322
rect 156 2319 157 2320
rect 151 2318 157 2319
rect 226 2319 227 2320
rect 231 2319 232 2323
rect 226 2318 232 2319
rect 279 2323 285 2324
rect 279 2319 280 2323
rect 284 2322 285 2323
rect 303 2323 309 2324
rect 303 2322 304 2323
rect 284 2320 304 2322
rect 284 2319 285 2320
rect 279 2318 285 2319
rect 303 2319 304 2320
rect 308 2319 309 2323
rect 303 2318 309 2319
rect 487 2323 496 2324
rect 487 2319 488 2323
rect 495 2319 496 2323
rect 487 2318 496 2319
rect 583 2323 589 2324
rect 583 2319 584 2323
rect 588 2322 589 2323
rect 679 2323 685 2324
rect 679 2322 680 2323
rect 588 2320 680 2322
rect 588 2319 589 2320
rect 583 2318 589 2319
rect 679 2319 680 2320
rect 684 2319 685 2323
rect 679 2318 685 2319
rect 775 2323 781 2324
rect 775 2319 776 2323
rect 780 2322 781 2323
rect 871 2323 877 2324
rect 871 2322 872 2323
rect 780 2320 872 2322
rect 780 2319 781 2320
rect 775 2318 781 2319
rect 871 2319 872 2320
rect 876 2319 877 2323
rect 871 2318 877 2319
rect 1063 2323 1069 2324
rect 1063 2319 1064 2323
rect 1068 2322 1069 2323
rect 1150 2323 1156 2324
rect 1150 2322 1151 2323
rect 1068 2320 1151 2322
rect 1068 2319 1069 2320
rect 1063 2318 1069 2319
rect 1150 2319 1151 2320
rect 1155 2319 1156 2323
rect 1239 2323 1245 2324
rect 1239 2322 1240 2323
rect 1150 2318 1156 2319
rect 1159 2320 1240 2322
rect 142 2313 148 2314
rect 142 2309 143 2313
rect 147 2309 148 2313
rect 142 2308 148 2309
rect 294 2313 300 2314
rect 294 2309 295 2313
rect 299 2309 300 2313
rect 294 2308 300 2309
rect 478 2313 484 2314
rect 478 2309 479 2313
rect 483 2309 484 2313
rect 478 2308 484 2309
rect 670 2313 676 2314
rect 670 2309 671 2313
rect 675 2309 676 2313
rect 670 2308 676 2309
rect 862 2313 868 2314
rect 862 2309 863 2313
rect 867 2309 868 2313
rect 862 2308 868 2309
rect 1054 2313 1060 2314
rect 1054 2309 1055 2313
rect 1059 2309 1060 2313
rect 1054 2308 1060 2309
rect 110 2300 116 2301
rect 110 2296 111 2300
rect 115 2296 116 2300
rect 583 2299 589 2300
rect 583 2298 584 2299
rect 533 2296 584 2298
rect 110 2295 116 2296
rect 226 2295 232 2296
rect 226 2291 227 2295
rect 231 2294 232 2295
rect 583 2295 584 2296
rect 588 2295 589 2299
rect 775 2299 781 2300
rect 775 2298 776 2299
rect 725 2296 776 2298
rect 583 2294 589 2295
rect 775 2295 776 2296
rect 780 2295 781 2299
rect 1159 2298 1161 2320
rect 1239 2319 1240 2320
rect 1244 2319 1245 2323
rect 1239 2318 1245 2319
rect 1415 2323 1421 2324
rect 1415 2319 1416 2323
rect 1420 2322 1421 2323
rect 1503 2323 1509 2324
rect 1503 2322 1504 2323
rect 1420 2320 1504 2322
rect 1420 2319 1421 2320
rect 1415 2318 1421 2319
rect 1503 2319 1504 2320
rect 1508 2319 1509 2323
rect 1503 2318 1509 2319
rect 1591 2323 1597 2324
rect 1591 2319 1592 2323
rect 1596 2322 1597 2323
rect 1650 2323 1656 2324
rect 1650 2322 1651 2323
rect 1596 2320 1651 2322
rect 1596 2319 1597 2320
rect 1591 2318 1597 2319
rect 1650 2319 1651 2320
rect 1655 2319 1656 2323
rect 1650 2318 1656 2319
rect 1743 2323 1749 2324
rect 1743 2319 1744 2323
rect 1748 2322 1749 2323
rect 1778 2323 1784 2324
rect 1778 2322 1779 2323
rect 1748 2320 1779 2322
rect 1748 2319 1749 2320
rect 1743 2318 1749 2319
rect 1778 2319 1779 2320
rect 1783 2319 1784 2323
rect 1894 2321 1895 2325
rect 1899 2321 1900 2325
rect 1894 2320 1900 2321
rect 2006 2325 2012 2326
rect 2006 2321 2007 2325
rect 2011 2321 2012 2325
rect 2006 2320 2012 2321
rect 2158 2325 2164 2326
rect 2158 2321 2159 2325
rect 2163 2321 2164 2325
rect 2158 2320 2164 2321
rect 2310 2325 2316 2326
rect 2310 2321 2311 2325
rect 2315 2321 2316 2325
rect 2310 2320 2316 2321
rect 2462 2325 2468 2326
rect 2462 2321 2463 2325
rect 2467 2321 2468 2325
rect 2462 2320 2468 2321
rect 2614 2325 2620 2326
rect 2614 2321 2615 2325
rect 2619 2321 2620 2325
rect 2614 2320 2620 2321
rect 2774 2325 2780 2326
rect 2774 2321 2775 2325
rect 2779 2321 2780 2325
rect 2774 2320 2780 2321
rect 2942 2325 2948 2326
rect 2942 2321 2943 2325
rect 2947 2321 2948 2325
rect 2942 2320 2948 2321
rect 3110 2325 3116 2326
rect 3110 2321 3111 2325
rect 3115 2321 3116 2325
rect 3110 2320 3116 2321
rect 3286 2325 3292 2326
rect 3286 2321 3287 2325
rect 3291 2321 3292 2325
rect 3286 2320 3292 2321
rect 3470 2325 3476 2326
rect 3470 2321 3471 2325
rect 3475 2321 3476 2325
rect 3470 2320 3476 2321
rect 1778 2318 1784 2319
rect 1230 2313 1236 2314
rect 1230 2309 1231 2313
rect 1235 2309 1236 2313
rect 1230 2308 1236 2309
rect 1406 2313 1412 2314
rect 1406 2309 1407 2313
rect 1411 2309 1412 2313
rect 1406 2308 1412 2309
rect 1582 2313 1588 2314
rect 1582 2309 1583 2313
rect 1587 2309 1588 2313
rect 1582 2308 1588 2309
rect 1734 2313 1740 2314
rect 1734 2309 1735 2313
rect 1739 2309 1740 2313
rect 1734 2308 1740 2309
rect 1862 2312 1868 2313
rect 3574 2312 3580 2313
rect 1862 2308 1863 2312
rect 1867 2308 1868 2312
rect 1959 2311 1965 2312
rect 1959 2310 1960 2311
rect 1949 2308 1960 2310
rect 1862 2307 1868 2308
rect 1959 2307 1960 2308
rect 1964 2307 1965 2311
rect 2087 2311 2093 2312
rect 2087 2310 2088 2311
rect 2061 2308 2088 2310
rect 1959 2306 1965 2307
rect 2087 2307 2088 2308
rect 2092 2307 2093 2311
rect 2239 2311 2245 2312
rect 2239 2310 2240 2311
rect 2213 2308 2240 2310
rect 2087 2306 2093 2307
rect 2239 2307 2240 2308
rect 2244 2307 2245 2311
rect 2391 2311 2397 2312
rect 2391 2310 2392 2311
rect 2365 2308 2392 2310
rect 2239 2306 2245 2307
rect 2391 2307 2392 2308
rect 2396 2307 2397 2311
rect 2743 2311 2749 2312
rect 2743 2310 2744 2311
rect 2669 2308 2744 2310
rect 2391 2306 2397 2307
rect 2402 2307 2408 2308
rect 2402 2303 2403 2307
rect 2407 2306 2408 2307
rect 2743 2307 2744 2308
rect 2748 2307 2749 2311
rect 2874 2311 2880 2312
rect 2874 2310 2875 2311
rect 2829 2308 2875 2310
rect 2743 2306 2749 2307
rect 2874 2307 2875 2308
rect 2879 2307 2880 2311
rect 3031 2311 3037 2312
rect 3031 2310 3032 2311
rect 2997 2308 3032 2310
rect 2874 2306 2880 2307
rect 3031 2307 3032 2308
rect 3036 2307 3037 2311
rect 3207 2311 3213 2312
rect 3207 2310 3208 2311
rect 3165 2308 3208 2310
rect 3031 2306 3037 2307
rect 3207 2307 3208 2308
rect 3212 2307 3213 2311
rect 3574 2308 3575 2312
rect 3579 2308 3580 2312
rect 3574 2307 3580 2308
rect 3207 2306 3213 2307
rect 2407 2304 2481 2306
rect 2407 2303 2408 2304
rect 2402 2302 2408 2303
rect 1109 2296 1161 2298
rect 1822 2300 1828 2301
rect 1822 2296 1823 2300
rect 1827 2296 1828 2300
rect 775 2294 781 2295
rect 846 2295 852 2296
rect 231 2292 313 2294
rect 231 2291 232 2292
rect 226 2290 232 2291
rect 846 2291 847 2295
rect 851 2294 852 2295
rect 1338 2295 1344 2296
rect 851 2292 881 2294
rect 851 2291 852 2292
rect 846 2290 852 2291
rect 1338 2291 1339 2295
rect 1343 2294 1344 2295
rect 1503 2295 1509 2296
rect 1343 2292 1425 2294
rect 1343 2291 1344 2292
rect 1338 2290 1344 2291
rect 1503 2291 1504 2295
rect 1508 2294 1509 2295
rect 1650 2295 1656 2296
rect 1822 2295 1828 2296
rect 1862 2295 1868 2296
rect 1508 2292 1601 2294
rect 1508 2291 1509 2292
rect 1503 2290 1509 2291
rect 1650 2291 1651 2295
rect 1655 2294 1656 2295
rect 1655 2292 1753 2294
rect 1655 2291 1656 2292
rect 1650 2290 1656 2291
rect 1862 2291 1863 2295
rect 1867 2291 1868 2295
rect 3574 2295 3580 2296
rect 1862 2290 1868 2291
rect 3204 2292 3297 2294
rect 1886 2285 1892 2286
rect 110 2283 116 2284
rect 110 2279 111 2283
rect 115 2279 116 2283
rect 1318 2283 1324 2284
rect 1318 2282 1319 2283
rect 1281 2280 1319 2282
rect 110 2278 116 2279
rect 1318 2279 1319 2280
rect 1323 2279 1324 2283
rect 1318 2278 1324 2279
rect 1822 2283 1828 2284
rect 1822 2279 1823 2283
rect 1827 2279 1828 2283
rect 1886 2281 1887 2285
rect 1891 2281 1892 2285
rect 1886 2280 1892 2281
rect 1998 2285 2004 2286
rect 1998 2281 1999 2285
rect 2003 2281 2004 2285
rect 1998 2280 2004 2281
rect 2150 2285 2156 2286
rect 2150 2281 2151 2285
rect 2155 2281 2156 2285
rect 2150 2280 2156 2281
rect 2302 2285 2308 2286
rect 2302 2281 2303 2285
rect 2307 2281 2308 2285
rect 2302 2280 2308 2281
rect 2454 2285 2460 2286
rect 2454 2281 2455 2285
rect 2459 2281 2460 2285
rect 2454 2280 2460 2281
rect 2606 2285 2612 2286
rect 2606 2281 2607 2285
rect 2611 2281 2612 2285
rect 2606 2280 2612 2281
rect 2766 2285 2772 2286
rect 2766 2281 2767 2285
rect 2771 2281 2772 2285
rect 2766 2280 2772 2281
rect 2934 2285 2940 2286
rect 2934 2281 2935 2285
rect 2939 2281 2940 2285
rect 2934 2280 2940 2281
rect 3102 2285 3108 2286
rect 3102 2281 3103 2285
rect 3107 2281 3108 2285
rect 3102 2280 3108 2281
rect 1822 2278 1828 2279
rect 2798 2279 2804 2280
rect 2798 2275 2799 2279
rect 2803 2278 2804 2279
rect 3204 2278 3206 2292
rect 3574 2291 3575 2295
rect 3579 2291 3580 2295
rect 3574 2290 3580 2291
rect 3278 2285 3284 2286
rect 3278 2281 3279 2285
rect 3283 2281 3284 2285
rect 3278 2280 3284 2281
rect 3462 2285 3468 2286
rect 3462 2281 3463 2285
rect 3467 2281 3468 2285
rect 3462 2280 3468 2281
rect 2803 2276 3206 2278
rect 3498 2279 3504 2280
rect 2803 2275 2804 2276
rect 2798 2274 2804 2275
rect 3498 2275 3499 2279
rect 3503 2278 3504 2279
rect 3511 2279 3517 2280
rect 3511 2278 3512 2279
rect 3503 2276 3512 2278
rect 3503 2275 3504 2276
rect 3498 2274 3504 2275
rect 3511 2275 3512 2276
rect 3516 2275 3517 2279
rect 3511 2274 3517 2275
rect 134 2273 140 2274
rect 134 2269 135 2273
rect 139 2269 140 2273
rect 134 2268 140 2269
rect 286 2273 292 2274
rect 286 2269 287 2273
rect 291 2269 292 2273
rect 286 2268 292 2269
rect 470 2273 476 2274
rect 470 2269 471 2273
rect 475 2269 476 2273
rect 470 2268 476 2269
rect 662 2273 668 2274
rect 662 2269 663 2273
rect 667 2269 668 2273
rect 662 2268 668 2269
rect 854 2273 860 2274
rect 854 2269 855 2273
rect 859 2269 860 2273
rect 854 2268 860 2269
rect 1046 2273 1052 2274
rect 1046 2269 1047 2273
rect 1051 2269 1052 2273
rect 1046 2268 1052 2269
rect 1222 2273 1228 2274
rect 1222 2269 1223 2273
rect 1227 2269 1228 2273
rect 1222 2268 1228 2269
rect 1398 2273 1404 2274
rect 1398 2269 1399 2273
rect 1403 2269 1404 2273
rect 1398 2268 1404 2269
rect 1574 2273 1580 2274
rect 1574 2269 1575 2273
rect 1579 2269 1580 2273
rect 1574 2268 1580 2269
rect 1726 2273 1732 2274
rect 1726 2269 1727 2273
rect 1731 2269 1732 2273
rect 1726 2268 1732 2269
rect 154 2267 160 2268
rect 154 2263 155 2267
rect 159 2266 160 2267
rect 183 2267 189 2268
rect 183 2266 184 2267
rect 159 2264 184 2266
rect 159 2263 160 2264
rect 154 2262 160 2263
rect 183 2263 184 2264
rect 188 2263 189 2267
rect 183 2262 189 2263
rect 1886 2259 1892 2260
rect 1886 2255 1887 2259
rect 1891 2255 1892 2259
rect 1886 2254 1892 2255
rect 2022 2259 2028 2260
rect 2022 2255 2023 2259
rect 2027 2255 2028 2259
rect 2022 2254 2028 2255
rect 2198 2259 2204 2260
rect 2198 2255 2199 2259
rect 2203 2255 2204 2259
rect 2198 2254 2204 2255
rect 2382 2259 2388 2260
rect 2382 2255 2383 2259
rect 2387 2255 2388 2259
rect 2382 2254 2388 2255
rect 2566 2259 2572 2260
rect 2566 2255 2567 2259
rect 2571 2255 2572 2259
rect 2566 2254 2572 2255
rect 2742 2259 2748 2260
rect 2742 2255 2743 2259
rect 2747 2255 2748 2259
rect 2742 2254 2748 2255
rect 2910 2259 2916 2260
rect 2910 2255 2911 2259
rect 2915 2255 2916 2259
rect 2910 2254 2916 2255
rect 3078 2259 3084 2260
rect 3078 2255 3079 2259
rect 3083 2255 3084 2259
rect 3078 2254 3084 2255
rect 3238 2259 3244 2260
rect 3238 2255 3239 2259
rect 3243 2255 3244 2259
rect 3238 2254 3244 2255
rect 3406 2259 3412 2260
rect 3406 2255 3407 2259
rect 3411 2255 3412 2259
rect 3406 2254 3412 2255
rect 2478 2251 2484 2252
rect 1862 2249 1868 2250
rect 1862 2245 1863 2249
rect 1867 2245 1868 2249
rect 2478 2247 2479 2251
rect 2483 2250 2484 2251
rect 3146 2251 3152 2252
rect 2483 2248 2585 2250
rect 2483 2247 2484 2248
rect 2478 2246 2484 2247
rect 3146 2247 3147 2251
rect 3151 2250 3152 2251
rect 3359 2251 3365 2252
rect 3151 2248 3257 2250
rect 3151 2247 3152 2248
rect 3146 2246 3152 2247
rect 3359 2247 3360 2251
rect 3364 2250 3365 2251
rect 3364 2248 3425 2250
rect 3574 2249 3580 2250
rect 3364 2247 3365 2248
rect 3359 2246 3365 2247
rect 1862 2244 1868 2245
rect 3574 2245 3575 2249
rect 3579 2245 3580 2249
rect 3574 2244 3580 2245
rect 134 2243 140 2244
rect 134 2239 135 2243
rect 139 2239 140 2243
rect 134 2238 140 2239
rect 254 2243 260 2244
rect 254 2239 255 2243
rect 259 2239 260 2243
rect 254 2238 260 2239
rect 406 2243 412 2244
rect 406 2239 407 2243
rect 411 2239 412 2243
rect 406 2238 412 2239
rect 558 2243 564 2244
rect 558 2239 559 2243
rect 563 2239 564 2243
rect 558 2238 564 2239
rect 718 2243 724 2244
rect 718 2239 719 2243
rect 723 2239 724 2243
rect 718 2238 724 2239
rect 870 2243 876 2244
rect 870 2239 871 2243
rect 875 2239 876 2243
rect 870 2238 876 2239
rect 1014 2243 1020 2244
rect 1014 2239 1015 2243
rect 1019 2239 1020 2243
rect 1014 2238 1020 2239
rect 1158 2243 1164 2244
rect 1158 2239 1159 2243
rect 1163 2239 1164 2243
rect 1158 2238 1164 2239
rect 1302 2243 1308 2244
rect 1302 2239 1303 2243
rect 1307 2239 1308 2243
rect 1302 2238 1308 2239
rect 1454 2243 1460 2244
rect 1454 2239 1455 2243
rect 1459 2239 1460 2243
rect 1454 2238 1460 2239
rect 374 2235 380 2236
rect 110 2233 116 2234
rect 110 2229 111 2233
rect 115 2229 116 2233
rect 374 2231 375 2235
rect 379 2234 380 2235
rect 490 2235 496 2236
rect 379 2232 425 2234
rect 379 2231 380 2232
rect 374 2230 380 2231
rect 490 2231 491 2235
rect 495 2234 496 2235
rect 1398 2235 1404 2236
rect 495 2232 577 2234
rect 495 2231 496 2232
rect 490 2230 496 2231
rect 1398 2231 1399 2235
rect 1403 2234 1404 2235
rect 2015 2235 2021 2236
rect 2015 2234 2016 2235
rect 1403 2232 1473 2234
rect 1822 2233 1828 2234
rect 1403 2231 1404 2232
rect 1398 2230 1404 2231
rect 110 2228 116 2229
rect 1822 2229 1823 2233
rect 1827 2229 1828 2233
rect 1822 2228 1828 2229
rect 1862 2232 1868 2233
rect 1949 2232 2016 2234
rect 1862 2228 1863 2232
rect 1867 2228 1868 2232
rect 2015 2231 2016 2232
rect 2020 2231 2021 2235
rect 2191 2235 2197 2236
rect 2191 2234 2192 2235
rect 2085 2232 2192 2234
rect 2015 2230 2021 2231
rect 2191 2231 2192 2232
rect 2196 2231 2197 2235
rect 2375 2235 2381 2236
rect 2375 2234 2376 2235
rect 2261 2232 2376 2234
rect 2191 2230 2197 2231
rect 2375 2231 2376 2232
rect 2380 2231 2381 2235
rect 2559 2235 2565 2236
rect 2559 2234 2560 2235
rect 2445 2232 2560 2234
rect 2375 2230 2381 2231
rect 2559 2231 2560 2232
rect 2564 2231 2565 2235
rect 2903 2235 2909 2236
rect 2903 2234 2904 2235
rect 2805 2232 2904 2234
rect 2559 2230 2565 2231
rect 2903 2231 2904 2232
rect 2908 2231 2909 2235
rect 3071 2235 3077 2236
rect 3071 2234 3072 2235
rect 2973 2232 3072 2234
rect 2903 2230 2909 2231
rect 3071 2231 3072 2232
rect 3076 2231 3077 2235
rect 3231 2235 3237 2236
rect 3231 2234 3232 2235
rect 3141 2232 3232 2234
rect 3071 2230 3077 2231
rect 3231 2231 3232 2232
rect 3236 2231 3237 2235
rect 3231 2230 3237 2231
rect 3574 2232 3580 2233
rect 1862 2227 1868 2228
rect 3574 2228 3575 2232
rect 3579 2228 3580 2232
rect 3574 2227 3580 2228
rect 247 2219 253 2220
rect 247 2218 248 2219
rect 110 2216 116 2217
rect 197 2216 248 2218
rect 110 2212 111 2216
rect 115 2212 116 2216
rect 247 2215 248 2216
rect 252 2215 253 2219
rect 399 2219 405 2220
rect 399 2218 400 2219
rect 317 2216 400 2218
rect 247 2214 253 2215
rect 399 2215 400 2216
rect 404 2215 405 2219
rect 399 2214 405 2215
rect 626 2219 632 2220
rect 626 2215 627 2219
rect 631 2218 632 2219
rect 1007 2219 1013 2220
rect 1007 2218 1008 2219
rect 631 2216 745 2218
rect 933 2216 1008 2218
rect 631 2215 632 2216
rect 626 2214 632 2215
rect 1007 2215 1008 2216
rect 1012 2215 1013 2219
rect 1082 2219 1088 2220
rect 1082 2218 1083 2219
rect 1077 2216 1083 2218
rect 1007 2214 1013 2215
rect 1082 2215 1083 2216
rect 1087 2215 1088 2219
rect 1082 2214 1088 2215
rect 1098 2219 1104 2220
rect 1098 2215 1099 2219
rect 1103 2218 1104 2219
rect 1447 2219 1453 2220
rect 1447 2218 1448 2219
rect 1103 2216 1185 2218
rect 1365 2216 1448 2218
rect 1103 2215 1104 2216
rect 1098 2214 1104 2215
rect 1447 2215 1448 2216
rect 1452 2215 1453 2219
rect 1894 2219 1900 2220
rect 1447 2214 1453 2215
rect 1822 2216 1828 2217
rect 110 2211 116 2212
rect 1822 2212 1823 2216
rect 1827 2212 1828 2216
rect 1894 2215 1895 2219
rect 1899 2215 1900 2219
rect 1894 2214 1900 2215
rect 2030 2219 2036 2220
rect 2030 2215 2031 2219
rect 2035 2215 2036 2219
rect 2030 2214 2036 2215
rect 2206 2219 2212 2220
rect 2206 2215 2207 2219
rect 2211 2215 2212 2219
rect 2206 2214 2212 2215
rect 2390 2219 2396 2220
rect 2390 2215 2391 2219
rect 2395 2215 2396 2219
rect 2390 2214 2396 2215
rect 2574 2219 2580 2220
rect 2574 2215 2575 2219
rect 2579 2215 2580 2219
rect 2574 2214 2580 2215
rect 2750 2219 2756 2220
rect 2750 2215 2751 2219
rect 2755 2215 2756 2219
rect 2750 2214 2756 2215
rect 2918 2219 2924 2220
rect 2918 2215 2919 2219
rect 2923 2215 2924 2219
rect 2918 2214 2924 2215
rect 3086 2219 3092 2220
rect 3086 2215 3087 2219
rect 3091 2215 3092 2219
rect 3086 2214 3092 2215
rect 3246 2219 3252 2220
rect 3246 2215 3247 2219
rect 3251 2215 3252 2219
rect 3246 2214 3252 2215
rect 3414 2219 3420 2220
rect 3414 2215 3415 2219
rect 3419 2215 3420 2219
rect 3414 2214 3420 2215
rect 1822 2211 1828 2212
rect 1903 2207 1909 2208
rect 142 2203 148 2204
rect 142 2199 143 2203
rect 147 2199 148 2203
rect 142 2198 148 2199
rect 262 2203 268 2204
rect 262 2199 263 2203
rect 267 2199 268 2203
rect 262 2198 268 2199
rect 414 2203 420 2204
rect 414 2199 415 2203
rect 419 2199 420 2203
rect 414 2198 420 2199
rect 566 2203 572 2204
rect 566 2199 567 2203
rect 571 2199 572 2203
rect 566 2198 572 2199
rect 726 2203 732 2204
rect 726 2199 727 2203
rect 731 2199 732 2203
rect 726 2198 732 2199
rect 878 2203 884 2204
rect 878 2199 879 2203
rect 883 2199 884 2203
rect 878 2198 884 2199
rect 1022 2203 1028 2204
rect 1022 2199 1023 2203
rect 1027 2199 1028 2203
rect 1022 2198 1028 2199
rect 1166 2203 1172 2204
rect 1166 2199 1167 2203
rect 1171 2199 1172 2203
rect 1166 2198 1172 2199
rect 1310 2203 1316 2204
rect 1310 2199 1311 2203
rect 1315 2199 1316 2203
rect 1310 2198 1316 2199
rect 1462 2203 1468 2204
rect 1462 2199 1463 2203
rect 1467 2199 1468 2203
rect 1903 2203 1904 2207
rect 1908 2206 1909 2207
rect 2006 2207 2012 2208
rect 2006 2206 2007 2207
rect 1908 2204 2007 2206
rect 1908 2203 1909 2204
rect 1903 2202 1909 2203
rect 2006 2203 2007 2204
rect 2011 2203 2012 2207
rect 2006 2202 2012 2203
rect 2015 2207 2021 2208
rect 2015 2203 2016 2207
rect 2020 2206 2021 2207
rect 2039 2207 2045 2208
rect 2039 2206 2040 2207
rect 2020 2204 2040 2206
rect 2020 2203 2021 2204
rect 2015 2202 2021 2203
rect 2039 2203 2040 2204
rect 2044 2203 2045 2207
rect 2039 2202 2045 2203
rect 2191 2207 2197 2208
rect 2191 2203 2192 2207
rect 2196 2206 2197 2207
rect 2215 2207 2221 2208
rect 2215 2206 2216 2207
rect 2196 2204 2216 2206
rect 2196 2203 2197 2204
rect 2191 2202 2197 2203
rect 2215 2203 2216 2204
rect 2220 2203 2221 2207
rect 2215 2202 2221 2203
rect 2375 2207 2381 2208
rect 2375 2203 2376 2207
rect 2380 2206 2381 2207
rect 2399 2207 2405 2208
rect 2399 2206 2400 2207
rect 2380 2204 2400 2206
rect 2380 2203 2381 2204
rect 2375 2202 2381 2203
rect 2399 2203 2400 2204
rect 2404 2203 2405 2207
rect 2399 2202 2405 2203
rect 2559 2207 2565 2208
rect 2559 2203 2560 2207
rect 2564 2206 2565 2207
rect 2583 2207 2589 2208
rect 2583 2206 2584 2207
rect 2564 2204 2584 2206
rect 2564 2203 2565 2204
rect 2559 2202 2565 2203
rect 2583 2203 2584 2204
rect 2588 2203 2589 2207
rect 2583 2202 2589 2203
rect 2759 2207 2765 2208
rect 2759 2203 2760 2207
rect 2764 2206 2765 2207
rect 2798 2207 2804 2208
rect 2798 2206 2799 2207
rect 2764 2204 2799 2206
rect 2764 2203 2765 2204
rect 2759 2202 2765 2203
rect 2798 2203 2799 2204
rect 2803 2203 2804 2207
rect 2798 2202 2804 2203
rect 2903 2207 2909 2208
rect 2903 2203 2904 2207
rect 2908 2206 2909 2207
rect 2927 2207 2933 2208
rect 2927 2206 2928 2207
rect 2908 2204 2928 2206
rect 2908 2203 2909 2204
rect 2903 2202 2909 2203
rect 2927 2203 2928 2204
rect 2932 2203 2933 2207
rect 2927 2202 2933 2203
rect 3071 2207 3077 2208
rect 3071 2203 3072 2207
rect 3076 2206 3077 2207
rect 3095 2207 3101 2208
rect 3095 2206 3096 2207
rect 3076 2204 3096 2206
rect 3076 2203 3077 2204
rect 3071 2202 3077 2203
rect 3095 2203 3096 2204
rect 3100 2203 3101 2207
rect 3095 2202 3101 2203
rect 3231 2207 3237 2208
rect 3231 2203 3232 2207
rect 3236 2206 3237 2207
rect 3255 2207 3261 2208
rect 3255 2206 3256 2207
rect 3236 2204 3256 2206
rect 3236 2203 3237 2204
rect 3231 2202 3237 2203
rect 3255 2203 3256 2204
rect 3260 2203 3261 2207
rect 3255 2202 3261 2203
rect 3423 2207 3432 2208
rect 3423 2203 3424 2207
rect 3431 2203 3432 2207
rect 3423 2202 3432 2203
rect 1462 2198 1468 2199
rect 151 2191 160 2192
rect 151 2187 152 2191
rect 159 2187 160 2191
rect 151 2186 160 2187
rect 247 2191 253 2192
rect 247 2187 248 2191
rect 252 2190 253 2191
rect 271 2191 277 2192
rect 271 2190 272 2191
rect 252 2188 272 2190
rect 252 2187 253 2188
rect 247 2186 253 2187
rect 271 2187 272 2188
rect 276 2187 277 2191
rect 271 2186 277 2187
rect 399 2191 405 2192
rect 399 2187 400 2191
rect 404 2190 405 2191
rect 423 2191 429 2192
rect 423 2190 424 2191
rect 404 2188 424 2190
rect 404 2187 405 2188
rect 399 2186 405 2187
rect 423 2187 424 2188
rect 428 2187 429 2191
rect 423 2186 429 2187
rect 575 2191 581 2192
rect 575 2187 576 2191
rect 580 2190 581 2191
rect 626 2191 632 2192
rect 626 2190 627 2191
rect 580 2188 627 2190
rect 580 2187 581 2188
rect 575 2186 581 2187
rect 626 2187 627 2188
rect 631 2187 632 2191
rect 626 2186 632 2187
rect 687 2191 693 2192
rect 687 2187 688 2191
rect 692 2190 693 2191
rect 735 2191 741 2192
rect 735 2190 736 2191
rect 692 2188 736 2190
rect 692 2187 693 2188
rect 687 2186 693 2187
rect 735 2187 736 2188
rect 740 2187 741 2191
rect 735 2186 741 2187
rect 887 2191 896 2192
rect 887 2187 888 2191
rect 895 2187 896 2191
rect 887 2186 896 2187
rect 1007 2191 1013 2192
rect 1007 2187 1008 2191
rect 1012 2190 1013 2191
rect 1031 2191 1037 2192
rect 1031 2190 1032 2191
rect 1012 2188 1032 2190
rect 1012 2187 1013 2188
rect 1007 2186 1013 2187
rect 1031 2187 1032 2188
rect 1036 2187 1037 2191
rect 1031 2186 1037 2187
rect 1175 2191 1181 2192
rect 1175 2187 1176 2191
rect 1180 2190 1181 2191
rect 1190 2191 1196 2192
rect 1190 2190 1191 2191
rect 1180 2188 1191 2190
rect 1180 2187 1181 2188
rect 1175 2186 1181 2187
rect 1190 2187 1191 2188
rect 1195 2187 1196 2191
rect 1190 2186 1196 2187
rect 1318 2191 1325 2192
rect 1318 2187 1319 2191
rect 1324 2187 1325 2191
rect 1318 2186 1325 2187
rect 1447 2191 1453 2192
rect 1447 2187 1448 2191
rect 1452 2190 1453 2191
rect 1471 2191 1477 2192
rect 1471 2190 1472 2191
rect 1452 2188 1472 2190
rect 1452 2187 1453 2188
rect 1447 2186 1453 2187
rect 1471 2187 1472 2188
rect 1476 2187 1477 2191
rect 1471 2186 1477 2187
rect 1879 2191 1885 2192
rect 1879 2187 1880 2191
rect 1884 2190 1885 2191
rect 1903 2191 1909 2192
rect 1903 2190 1904 2191
rect 1884 2188 1904 2190
rect 1884 2187 1885 2188
rect 1879 2186 1885 2187
rect 1903 2187 1904 2188
rect 1908 2187 1909 2191
rect 1903 2186 1909 2187
rect 1959 2191 1965 2192
rect 1959 2187 1960 2191
rect 1964 2190 1965 2191
rect 2047 2191 2053 2192
rect 2047 2190 2048 2191
rect 1964 2188 2048 2190
rect 1964 2187 1965 2188
rect 1959 2186 1965 2187
rect 2047 2187 2048 2188
rect 2052 2187 2053 2191
rect 2047 2186 2053 2187
rect 2135 2191 2141 2192
rect 2135 2187 2136 2191
rect 2140 2190 2141 2191
rect 2223 2191 2229 2192
rect 2223 2190 2224 2191
rect 2140 2188 2224 2190
rect 2140 2187 2141 2188
rect 2135 2186 2141 2187
rect 2223 2187 2224 2188
rect 2228 2187 2229 2191
rect 2223 2186 2229 2187
rect 2311 2191 2317 2192
rect 2311 2187 2312 2191
rect 2316 2190 2317 2191
rect 2407 2191 2413 2192
rect 2407 2190 2408 2191
rect 2316 2188 2408 2190
rect 2316 2187 2317 2188
rect 2311 2186 2317 2187
rect 2407 2187 2408 2188
rect 2412 2187 2413 2191
rect 2407 2186 2413 2187
rect 2495 2191 2501 2192
rect 2495 2187 2496 2191
rect 2500 2190 2501 2191
rect 2591 2191 2597 2192
rect 2591 2190 2592 2191
rect 2500 2188 2592 2190
rect 2500 2187 2501 2188
rect 2495 2186 2501 2187
rect 2591 2187 2592 2188
rect 2596 2187 2597 2191
rect 2591 2186 2597 2187
rect 2767 2191 2776 2192
rect 2767 2187 2768 2191
rect 2775 2187 2776 2191
rect 2767 2186 2776 2187
rect 2855 2191 2861 2192
rect 2855 2187 2856 2191
rect 2860 2190 2861 2191
rect 2927 2191 2933 2192
rect 2927 2190 2928 2191
rect 2860 2188 2928 2190
rect 2860 2187 2861 2188
rect 2855 2186 2861 2187
rect 2927 2187 2928 2188
rect 2932 2187 2933 2191
rect 2927 2186 2933 2187
rect 2999 2191 3005 2192
rect 2999 2187 3000 2191
rect 3004 2190 3005 2191
rect 3079 2191 3085 2192
rect 3079 2190 3080 2191
rect 3004 2188 3080 2190
rect 3004 2187 3005 2188
rect 2999 2186 3005 2187
rect 3079 2187 3080 2188
rect 3084 2187 3085 2191
rect 3079 2186 3085 2187
rect 3151 2191 3157 2192
rect 3151 2187 3152 2191
rect 3156 2190 3157 2191
rect 3223 2191 3229 2192
rect 3223 2190 3224 2191
rect 3156 2188 3224 2190
rect 3156 2187 3157 2188
rect 3151 2186 3157 2187
rect 3223 2187 3224 2188
rect 3228 2187 3229 2191
rect 3223 2186 3229 2187
rect 3295 2191 3301 2192
rect 3295 2187 3296 2191
rect 3300 2190 3301 2191
rect 3367 2191 3373 2192
rect 3367 2190 3368 2191
rect 3300 2188 3368 2190
rect 3300 2187 3301 2188
rect 3295 2186 3301 2187
rect 3367 2187 3368 2188
rect 3372 2187 3373 2191
rect 3367 2186 3373 2187
rect 3495 2191 3504 2192
rect 3495 2187 3496 2191
rect 3503 2187 3504 2191
rect 3495 2186 3504 2187
rect 374 2183 380 2184
rect 374 2182 375 2183
rect 272 2180 375 2182
rect 223 2175 229 2176
rect 223 2171 224 2175
rect 228 2174 229 2175
rect 272 2174 274 2180
rect 374 2179 375 2180
rect 379 2179 380 2183
rect 898 2183 904 2184
rect 898 2182 899 2183
rect 374 2178 380 2179
rect 784 2180 899 2182
rect 228 2172 274 2174
rect 279 2175 285 2176
rect 228 2171 229 2172
rect 223 2170 229 2171
rect 279 2171 280 2175
rect 284 2174 285 2175
rect 319 2175 325 2176
rect 319 2174 320 2175
rect 284 2172 320 2174
rect 284 2171 285 2172
rect 279 2170 285 2171
rect 319 2171 320 2172
rect 324 2171 325 2175
rect 319 2170 325 2171
rect 423 2175 429 2176
rect 423 2171 424 2175
rect 428 2174 429 2175
rect 479 2175 485 2176
rect 428 2172 474 2174
rect 428 2171 429 2172
rect 423 2170 429 2171
rect 472 2166 474 2172
rect 479 2171 480 2175
rect 484 2174 485 2175
rect 527 2175 533 2176
rect 527 2174 528 2175
rect 484 2172 528 2174
rect 484 2171 485 2172
rect 479 2170 485 2171
rect 527 2171 528 2172
rect 532 2171 533 2175
rect 527 2170 533 2171
rect 583 2175 589 2176
rect 583 2171 584 2175
rect 588 2174 589 2175
rect 631 2175 637 2176
rect 631 2174 632 2175
rect 588 2172 632 2174
rect 588 2171 589 2172
rect 583 2170 589 2171
rect 631 2171 632 2172
rect 636 2171 637 2175
rect 631 2170 637 2171
rect 735 2175 741 2176
rect 735 2171 736 2175
rect 740 2174 741 2175
rect 784 2174 786 2180
rect 898 2179 899 2180
rect 903 2179 904 2183
rect 1127 2183 1133 2184
rect 1127 2182 1128 2183
rect 898 2178 904 2179
rect 1056 2180 1128 2182
rect 740 2172 786 2174
rect 791 2175 797 2176
rect 740 2171 741 2172
rect 735 2170 741 2171
rect 791 2171 792 2175
rect 796 2174 797 2175
rect 839 2175 845 2176
rect 839 2174 840 2175
rect 796 2172 840 2174
rect 796 2171 797 2172
rect 791 2170 797 2171
rect 839 2171 840 2172
rect 844 2171 845 2175
rect 839 2170 845 2171
rect 951 2175 957 2176
rect 951 2171 952 2175
rect 956 2174 957 2175
rect 1056 2174 1058 2180
rect 1127 2179 1128 2180
rect 1132 2179 1133 2183
rect 1127 2178 1133 2179
rect 1894 2181 1900 2182
rect 1894 2177 1895 2181
rect 1899 2177 1900 2181
rect 1894 2176 1900 2177
rect 2038 2181 2044 2182
rect 2038 2177 2039 2181
rect 2043 2177 2044 2181
rect 2038 2176 2044 2177
rect 2214 2181 2220 2182
rect 2214 2177 2215 2181
rect 2219 2177 2220 2181
rect 2214 2176 2220 2177
rect 2398 2181 2404 2182
rect 2398 2177 2399 2181
rect 2403 2177 2404 2181
rect 2398 2176 2404 2177
rect 2582 2181 2588 2182
rect 2582 2177 2583 2181
rect 2587 2177 2588 2181
rect 2582 2176 2588 2177
rect 2758 2181 2764 2182
rect 2758 2177 2759 2181
rect 2763 2177 2764 2181
rect 2758 2176 2764 2177
rect 2918 2181 2924 2182
rect 2918 2177 2919 2181
rect 2923 2177 2924 2181
rect 2918 2176 2924 2177
rect 3070 2181 3076 2182
rect 3070 2177 3071 2181
rect 3075 2177 3076 2181
rect 3070 2176 3076 2177
rect 3214 2181 3220 2182
rect 3214 2177 3215 2181
rect 3219 2177 3220 2181
rect 3214 2176 3220 2177
rect 3358 2181 3364 2182
rect 3358 2177 3359 2181
rect 3363 2177 3364 2181
rect 3358 2176 3364 2177
rect 3486 2181 3492 2182
rect 3486 2177 3487 2181
rect 3491 2177 3492 2181
rect 3486 2176 3492 2177
rect 956 2172 1058 2174
rect 1063 2175 1069 2176
rect 956 2171 957 2172
rect 951 2170 957 2171
rect 1063 2171 1064 2175
rect 1068 2174 1069 2175
rect 1082 2175 1088 2176
rect 1082 2174 1083 2175
rect 1068 2172 1083 2174
rect 1068 2171 1069 2172
rect 1063 2170 1069 2171
rect 1082 2171 1083 2172
rect 1087 2171 1088 2175
rect 1082 2170 1088 2171
rect 1119 2175 1125 2176
rect 1119 2171 1120 2175
rect 1124 2174 1125 2175
rect 1175 2175 1181 2176
rect 1175 2174 1176 2175
rect 1124 2172 1176 2174
rect 1124 2171 1125 2172
rect 1119 2170 1125 2171
rect 1175 2171 1176 2172
rect 1180 2171 1181 2175
rect 1175 2170 1181 2171
rect 1862 2168 1868 2169
rect 3574 2168 3580 2169
rect 490 2167 496 2168
rect 490 2166 491 2167
rect 214 2165 220 2166
rect 214 2161 215 2165
rect 219 2161 220 2165
rect 214 2160 220 2161
rect 310 2165 316 2166
rect 310 2161 311 2165
rect 315 2161 316 2165
rect 310 2160 316 2161
rect 414 2165 420 2166
rect 414 2161 415 2165
rect 419 2161 420 2165
rect 472 2164 491 2166
rect 490 2163 491 2164
rect 495 2163 496 2167
rect 490 2162 496 2163
rect 518 2165 524 2166
rect 414 2160 420 2161
rect 518 2161 519 2165
rect 523 2161 524 2165
rect 518 2160 524 2161
rect 622 2165 628 2166
rect 622 2161 623 2165
rect 627 2161 628 2165
rect 622 2160 628 2161
rect 726 2165 732 2166
rect 726 2161 727 2165
rect 731 2161 732 2165
rect 726 2160 732 2161
rect 830 2165 836 2166
rect 830 2161 831 2165
rect 835 2161 836 2165
rect 830 2160 836 2161
rect 942 2165 948 2166
rect 942 2161 943 2165
rect 947 2161 948 2165
rect 942 2160 948 2161
rect 1054 2165 1060 2166
rect 1054 2161 1055 2165
rect 1059 2161 1060 2165
rect 1054 2160 1060 2161
rect 1166 2165 1172 2166
rect 1166 2161 1167 2165
rect 1171 2161 1172 2165
rect 1862 2164 1863 2168
rect 1867 2164 1868 2168
rect 1959 2167 1965 2168
rect 1959 2166 1960 2167
rect 1949 2164 1960 2166
rect 1862 2163 1868 2164
rect 1959 2163 1960 2164
rect 1964 2163 1965 2167
rect 2135 2167 2141 2168
rect 2135 2166 2136 2167
rect 2093 2164 2136 2166
rect 1959 2162 1965 2163
rect 2135 2163 2136 2164
rect 2140 2163 2141 2167
rect 2311 2167 2317 2168
rect 2311 2166 2312 2167
rect 2269 2164 2312 2166
rect 2135 2162 2141 2163
rect 2311 2163 2312 2164
rect 2316 2163 2317 2167
rect 2495 2167 2501 2168
rect 2495 2166 2496 2167
rect 2453 2164 2496 2166
rect 2311 2162 2317 2163
rect 2495 2163 2496 2164
rect 2500 2163 2501 2167
rect 2855 2167 2861 2168
rect 2855 2166 2856 2167
rect 2813 2164 2856 2166
rect 2495 2162 2501 2163
rect 2506 2163 2512 2164
rect 1166 2160 1172 2161
rect 2506 2159 2507 2163
rect 2511 2162 2512 2163
rect 2855 2163 2856 2164
rect 2860 2163 2861 2167
rect 2999 2167 3005 2168
rect 2999 2166 3000 2167
rect 2973 2164 3000 2166
rect 2855 2162 2861 2163
rect 2999 2163 3000 2164
rect 3004 2163 3005 2167
rect 3151 2167 3157 2168
rect 3151 2166 3152 2167
rect 3125 2164 3152 2166
rect 2999 2162 3005 2163
rect 3151 2163 3152 2164
rect 3156 2163 3157 2167
rect 3295 2167 3301 2168
rect 3295 2166 3296 2167
rect 3269 2164 3296 2166
rect 3151 2162 3157 2163
rect 3295 2163 3296 2164
rect 3300 2163 3301 2167
rect 3574 2164 3575 2168
rect 3579 2164 3580 2168
rect 3574 2163 3580 2164
rect 3295 2162 3301 2163
rect 2511 2160 2601 2162
rect 2511 2159 2512 2160
rect 2506 2158 2512 2159
rect 110 2152 116 2153
rect 1822 2152 1828 2153
rect 110 2148 111 2152
rect 115 2148 116 2152
rect 279 2151 285 2152
rect 279 2150 280 2151
rect 269 2148 280 2150
rect 110 2147 116 2148
rect 279 2147 280 2148
rect 284 2147 285 2151
rect 479 2151 485 2152
rect 479 2150 480 2151
rect 469 2148 480 2150
rect 279 2146 285 2147
rect 479 2147 480 2148
rect 484 2147 485 2151
rect 583 2151 589 2152
rect 583 2150 584 2151
rect 573 2148 584 2150
rect 479 2146 485 2147
rect 583 2147 584 2148
rect 588 2147 589 2151
rect 687 2151 693 2152
rect 687 2150 688 2151
rect 677 2148 688 2150
rect 583 2146 589 2147
rect 687 2147 688 2148
rect 692 2147 693 2151
rect 791 2151 797 2152
rect 791 2150 792 2151
rect 781 2148 792 2150
rect 687 2146 693 2147
rect 791 2147 792 2148
rect 796 2147 797 2151
rect 1119 2151 1125 2152
rect 1119 2150 1120 2151
rect 1109 2148 1120 2150
rect 791 2146 797 2147
rect 898 2147 904 2148
rect 898 2143 899 2147
rect 903 2146 904 2147
rect 1119 2147 1120 2148
rect 1124 2147 1125 2151
rect 1822 2148 1823 2152
rect 1827 2148 1828 2152
rect 1119 2146 1125 2147
rect 1127 2147 1133 2148
rect 1822 2147 1828 2148
rect 1862 2151 1868 2152
rect 1862 2147 1863 2151
rect 1867 2147 1868 2151
rect 903 2144 961 2146
rect 903 2143 904 2144
rect 898 2142 904 2143
rect 1127 2143 1128 2147
rect 1132 2146 1133 2147
rect 1862 2146 1868 2147
rect 3334 2151 3340 2152
rect 3334 2147 3335 2151
rect 3339 2150 3340 2151
rect 3574 2151 3580 2152
rect 3339 2148 3369 2150
rect 3339 2147 3340 2148
rect 3334 2146 3340 2147
rect 3574 2147 3575 2151
rect 3579 2147 3580 2151
rect 3574 2146 3580 2147
rect 1132 2144 1185 2146
rect 1132 2143 1133 2144
rect 1127 2142 1133 2143
rect 1886 2141 1892 2142
rect 1886 2137 1887 2141
rect 1891 2137 1892 2141
rect 1886 2136 1892 2137
rect 2030 2141 2036 2142
rect 2030 2137 2031 2141
rect 2035 2137 2036 2141
rect 2030 2136 2036 2137
rect 2206 2141 2212 2142
rect 2206 2137 2207 2141
rect 2211 2137 2212 2141
rect 2206 2136 2212 2137
rect 2390 2141 2396 2142
rect 2390 2137 2391 2141
rect 2395 2137 2396 2141
rect 2390 2136 2396 2137
rect 2574 2141 2580 2142
rect 2574 2137 2575 2141
rect 2579 2137 2580 2141
rect 2574 2136 2580 2137
rect 2750 2141 2756 2142
rect 2750 2137 2751 2141
rect 2755 2137 2756 2141
rect 2750 2136 2756 2137
rect 2910 2141 2916 2142
rect 2910 2137 2911 2141
rect 2915 2137 2916 2141
rect 2910 2136 2916 2137
rect 3062 2141 3068 2142
rect 3062 2137 3063 2141
rect 3067 2137 3068 2141
rect 3062 2136 3068 2137
rect 3206 2141 3212 2142
rect 3206 2137 3207 2141
rect 3211 2137 3212 2141
rect 3206 2136 3212 2137
rect 3350 2141 3356 2142
rect 3350 2137 3351 2141
rect 3355 2137 3356 2141
rect 3350 2136 3356 2137
rect 3478 2141 3484 2142
rect 3478 2137 3479 2141
rect 3483 2137 3484 2141
rect 3478 2136 3484 2137
rect 110 2135 116 2136
rect 110 2131 111 2135
rect 115 2131 116 2135
rect 110 2130 116 2131
rect 1822 2135 1828 2136
rect 1822 2131 1823 2135
rect 1827 2131 1828 2135
rect 1822 2130 1828 2131
rect 3498 2135 3504 2136
rect 3498 2131 3499 2135
rect 3503 2134 3504 2135
rect 3527 2135 3533 2136
rect 3527 2134 3528 2135
rect 3503 2132 3528 2134
rect 3503 2131 3504 2132
rect 3498 2130 3504 2131
rect 3527 2131 3528 2132
rect 3532 2131 3533 2135
rect 3527 2130 3533 2131
rect 206 2125 212 2126
rect 206 2121 207 2125
rect 211 2121 212 2125
rect 206 2120 212 2121
rect 302 2125 308 2126
rect 302 2121 303 2125
rect 307 2121 308 2125
rect 302 2120 308 2121
rect 406 2125 412 2126
rect 406 2121 407 2125
rect 411 2121 412 2125
rect 406 2120 412 2121
rect 510 2125 516 2126
rect 510 2121 511 2125
rect 515 2121 516 2125
rect 510 2120 516 2121
rect 614 2125 620 2126
rect 614 2121 615 2125
rect 619 2121 620 2125
rect 614 2120 620 2121
rect 718 2125 724 2126
rect 718 2121 719 2125
rect 723 2121 724 2125
rect 718 2120 724 2121
rect 822 2125 828 2126
rect 822 2121 823 2125
rect 827 2121 828 2125
rect 822 2120 828 2121
rect 934 2125 940 2126
rect 934 2121 935 2125
rect 939 2121 940 2125
rect 934 2120 940 2121
rect 1046 2125 1052 2126
rect 1046 2121 1047 2125
rect 1051 2121 1052 2125
rect 1046 2120 1052 2121
rect 1158 2125 1164 2126
rect 1158 2121 1159 2125
rect 1163 2121 1164 2125
rect 1158 2120 1164 2121
rect 338 2119 344 2120
rect 338 2115 339 2119
rect 343 2118 344 2119
rect 351 2119 357 2120
rect 351 2118 352 2119
rect 343 2116 352 2118
rect 343 2115 344 2116
rect 338 2114 344 2115
rect 351 2115 352 2116
rect 356 2115 357 2119
rect 351 2114 357 2115
rect 850 2119 856 2120
rect 850 2115 851 2119
rect 855 2118 856 2119
rect 871 2119 877 2120
rect 871 2118 872 2119
rect 855 2116 872 2118
rect 855 2115 856 2116
rect 850 2114 856 2115
rect 871 2115 872 2116
rect 876 2115 877 2119
rect 871 2114 877 2115
rect 1886 2115 1892 2116
rect 1886 2111 1887 2115
rect 1891 2111 1892 2115
rect 1886 2110 1892 2111
rect 2022 2115 2028 2116
rect 2022 2111 2023 2115
rect 2027 2111 2028 2115
rect 2022 2110 2028 2111
rect 2198 2115 2204 2116
rect 2198 2111 2199 2115
rect 2203 2111 2204 2115
rect 2198 2110 2204 2111
rect 2374 2115 2380 2116
rect 2374 2111 2375 2115
rect 2379 2111 2380 2115
rect 2374 2110 2380 2111
rect 2550 2115 2556 2116
rect 2550 2111 2551 2115
rect 2555 2111 2556 2115
rect 2550 2110 2556 2111
rect 2718 2115 2724 2116
rect 2718 2111 2719 2115
rect 2723 2111 2724 2115
rect 2718 2110 2724 2111
rect 2878 2115 2884 2116
rect 2878 2111 2879 2115
rect 2883 2111 2884 2115
rect 2878 2110 2884 2111
rect 3030 2115 3036 2116
rect 3030 2111 3031 2115
rect 3035 2111 3036 2115
rect 3030 2110 3036 2111
rect 3174 2115 3180 2116
rect 3174 2111 3175 2115
rect 3179 2111 3180 2115
rect 3174 2110 3180 2111
rect 3318 2115 3324 2116
rect 3318 2111 3319 2115
rect 3323 2111 3324 2115
rect 3318 2110 3324 2111
rect 3470 2115 3476 2116
rect 3470 2111 3471 2115
rect 3475 2111 3476 2115
rect 3470 2110 3476 2111
rect 1879 2107 1885 2108
rect 1862 2105 1868 2106
rect 1862 2101 1863 2105
rect 1867 2101 1868 2105
rect 1879 2103 1880 2107
rect 1884 2106 1885 2107
rect 2478 2107 2484 2108
rect 1884 2104 1905 2106
rect 1884 2103 1885 2104
rect 1879 2102 1885 2103
rect 2478 2103 2479 2107
rect 2483 2106 2484 2107
rect 3426 2107 3432 2108
rect 2483 2104 2569 2106
rect 2483 2103 2484 2104
rect 2478 2102 2484 2103
rect 3426 2103 3427 2107
rect 3431 2106 3432 2107
rect 3431 2104 3489 2106
rect 3574 2105 3580 2106
rect 3431 2103 3432 2104
rect 3426 2102 3432 2103
rect 1862 2100 1868 2101
rect 3574 2101 3575 2105
rect 3579 2101 3580 2105
rect 3574 2100 3580 2101
rect 318 2095 324 2096
rect 318 2091 319 2095
rect 323 2091 324 2095
rect 318 2090 324 2091
rect 422 2095 428 2096
rect 422 2091 423 2095
rect 427 2091 428 2095
rect 422 2090 428 2091
rect 526 2095 532 2096
rect 526 2091 527 2095
rect 531 2091 532 2095
rect 526 2090 532 2091
rect 630 2095 636 2096
rect 630 2091 631 2095
rect 635 2091 636 2095
rect 630 2090 636 2091
rect 734 2095 740 2096
rect 734 2091 735 2095
rect 739 2091 740 2095
rect 734 2090 740 2091
rect 830 2095 836 2096
rect 830 2091 831 2095
rect 835 2091 836 2095
rect 830 2090 836 2091
rect 926 2095 932 2096
rect 926 2091 927 2095
rect 931 2091 932 2095
rect 926 2090 932 2091
rect 1030 2095 1036 2096
rect 1030 2091 1031 2095
rect 1035 2091 1036 2095
rect 1030 2090 1036 2091
rect 1134 2095 1140 2096
rect 1134 2091 1135 2095
rect 1139 2091 1140 2095
rect 1134 2090 1140 2091
rect 1238 2095 1244 2096
rect 1238 2091 1239 2095
rect 1243 2091 1244 2095
rect 1238 2090 1244 2091
rect 1954 2091 1960 2092
rect 1862 2088 1868 2089
rect 407 2087 413 2088
rect 110 2085 116 2086
rect 110 2081 111 2085
rect 115 2081 116 2085
rect 407 2083 408 2087
rect 412 2086 413 2087
rect 490 2087 496 2088
rect 412 2084 441 2086
rect 412 2083 413 2084
rect 407 2082 413 2083
rect 490 2083 491 2087
rect 495 2086 496 2087
rect 495 2084 545 2086
rect 1822 2085 1828 2086
rect 495 2083 496 2084
rect 490 2082 496 2083
rect 110 2080 116 2081
rect 1822 2081 1823 2085
rect 1827 2081 1828 2085
rect 1862 2084 1863 2088
rect 1867 2084 1868 2088
rect 1954 2087 1955 2091
rect 1959 2090 1960 2091
rect 2367 2091 2373 2092
rect 2367 2090 2368 2091
rect 1959 2088 2049 2090
rect 2261 2088 2368 2090
rect 1959 2087 1960 2088
rect 1954 2086 1960 2087
rect 2367 2087 2368 2088
rect 2372 2087 2373 2091
rect 2543 2091 2549 2092
rect 2543 2090 2544 2091
rect 2437 2088 2544 2090
rect 2367 2086 2373 2087
rect 2543 2087 2544 2088
rect 2548 2087 2549 2091
rect 2543 2086 2549 2087
rect 2618 2091 2624 2092
rect 2618 2087 2619 2091
rect 2623 2090 2624 2091
rect 2790 2091 2796 2092
rect 2623 2088 2745 2090
rect 2623 2087 2624 2088
rect 2618 2086 2624 2087
rect 2790 2087 2791 2091
rect 2795 2090 2796 2091
rect 2946 2091 2952 2092
rect 2795 2088 2905 2090
rect 2795 2087 2796 2088
rect 2790 2086 2796 2087
rect 2946 2087 2947 2091
rect 2951 2090 2952 2091
rect 3098 2091 3104 2092
rect 2951 2088 3057 2090
rect 2951 2087 2952 2088
rect 2946 2086 2952 2087
rect 3098 2087 3099 2091
rect 3103 2090 3104 2091
rect 3242 2091 3248 2092
rect 3103 2088 3201 2090
rect 3103 2087 3104 2088
rect 3098 2086 3104 2087
rect 3242 2087 3243 2091
rect 3247 2090 3248 2091
rect 3247 2088 3345 2090
rect 3574 2088 3580 2089
rect 3247 2087 3248 2088
rect 3242 2086 3248 2087
rect 1862 2083 1868 2084
rect 3574 2084 3575 2088
rect 3579 2084 3580 2088
rect 3574 2083 3580 2084
rect 1822 2080 1828 2081
rect 1894 2075 1900 2076
rect 415 2071 421 2072
rect 415 2070 416 2071
rect 110 2068 116 2069
rect 381 2068 416 2070
rect 110 2064 111 2068
rect 115 2064 116 2068
rect 415 2067 416 2068
rect 420 2067 421 2071
rect 415 2066 421 2067
rect 599 2071 605 2072
rect 599 2067 600 2071
rect 604 2070 605 2071
rect 703 2071 709 2072
rect 604 2068 657 2070
rect 604 2067 605 2068
rect 599 2066 605 2067
rect 703 2067 704 2071
rect 708 2070 709 2071
rect 919 2071 925 2072
rect 919 2070 920 2071
rect 708 2068 761 2070
rect 893 2068 920 2070
rect 708 2067 709 2068
rect 703 2066 709 2067
rect 919 2067 920 2068
rect 924 2067 925 2071
rect 1023 2071 1029 2072
rect 1023 2070 1024 2071
rect 989 2068 1024 2070
rect 919 2066 925 2067
rect 1023 2067 1024 2068
rect 1028 2067 1029 2071
rect 1127 2071 1133 2072
rect 1127 2070 1128 2071
rect 1093 2068 1128 2070
rect 1023 2066 1029 2067
rect 1127 2067 1128 2068
rect 1132 2067 1133 2071
rect 1206 2071 1212 2072
rect 1206 2070 1207 2071
rect 1197 2068 1207 2070
rect 1127 2066 1133 2067
rect 1206 2067 1207 2068
rect 1211 2067 1212 2071
rect 1206 2066 1212 2067
rect 1214 2071 1220 2072
rect 1214 2067 1215 2071
rect 1219 2070 1220 2071
rect 1894 2071 1895 2075
rect 1899 2071 1900 2075
rect 1894 2070 1900 2071
rect 2030 2075 2036 2076
rect 2030 2071 2031 2075
rect 2035 2071 2036 2075
rect 2030 2070 2036 2071
rect 2206 2075 2212 2076
rect 2206 2071 2207 2075
rect 2211 2071 2212 2075
rect 2206 2070 2212 2071
rect 2382 2075 2388 2076
rect 2382 2071 2383 2075
rect 2387 2071 2388 2075
rect 2382 2070 2388 2071
rect 2558 2075 2564 2076
rect 2558 2071 2559 2075
rect 2563 2071 2564 2075
rect 2558 2070 2564 2071
rect 2726 2075 2732 2076
rect 2726 2071 2727 2075
rect 2731 2071 2732 2075
rect 2726 2070 2732 2071
rect 2886 2075 2892 2076
rect 2886 2071 2887 2075
rect 2891 2071 2892 2075
rect 2886 2070 2892 2071
rect 3038 2075 3044 2076
rect 3038 2071 3039 2075
rect 3043 2071 3044 2075
rect 3038 2070 3044 2071
rect 3182 2075 3188 2076
rect 3182 2071 3183 2075
rect 3187 2071 3188 2075
rect 3182 2070 3188 2071
rect 3326 2075 3332 2076
rect 3326 2071 3327 2075
rect 3331 2071 3332 2075
rect 3326 2070 3332 2071
rect 3478 2075 3484 2076
rect 3478 2071 3479 2075
rect 3483 2071 3484 2075
rect 3478 2070 3484 2071
rect 1219 2068 1265 2070
rect 1822 2068 1828 2069
rect 1219 2067 1220 2068
rect 1214 2066 1220 2067
rect 110 2063 116 2064
rect 1822 2064 1823 2068
rect 1827 2064 1828 2068
rect 1822 2063 1828 2064
rect 1903 2063 1909 2064
rect 1903 2059 1904 2063
rect 1908 2062 1909 2063
rect 1954 2063 1960 2064
rect 1954 2062 1955 2063
rect 1908 2060 1955 2062
rect 1908 2059 1909 2060
rect 1903 2058 1909 2059
rect 1954 2059 1955 2060
rect 1959 2059 1960 2063
rect 1954 2058 1960 2059
rect 2038 2063 2045 2064
rect 2038 2059 2039 2063
rect 2044 2059 2045 2063
rect 2038 2058 2045 2059
rect 2214 2063 2221 2064
rect 2214 2059 2215 2063
rect 2220 2059 2221 2063
rect 2214 2058 2221 2059
rect 2367 2063 2373 2064
rect 2367 2059 2368 2063
rect 2372 2062 2373 2063
rect 2391 2063 2397 2064
rect 2391 2062 2392 2063
rect 2372 2060 2392 2062
rect 2372 2059 2373 2060
rect 2367 2058 2373 2059
rect 2391 2059 2392 2060
rect 2396 2059 2397 2063
rect 2391 2058 2397 2059
rect 2543 2063 2549 2064
rect 2543 2059 2544 2063
rect 2548 2062 2549 2063
rect 2567 2063 2573 2064
rect 2567 2062 2568 2063
rect 2548 2060 2568 2062
rect 2548 2059 2549 2060
rect 2543 2058 2549 2059
rect 2567 2059 2568 2060
rect 2572 2059 2573 2063
rect 2567 2058 2573 2059
rect 2735 2063 2741 2064
rect 2735 2059 2736 2063
rect 2740 2062 2741 2063
rect 2790 2063 2796 2064
rect 2790 2062 2791 2063
rect 2740 2060 2791 2062
rect 2740 2059 2741 2060
rect 2735 2058 2741 2059
rect 2790 2059 2791 2060
rect 2795 2059 2796 2063
rect 2790 2058 2796 2059
rect 2895 2063 2901 2064
rect 2895 2059 2896 2063
rect 2900 2062 2901 2063
rect 2946 2063 2952 2064
rect 2946 2062 2947 2063
rect 2900 2060 2947 2062
rect 2900 2059 2901 2060
rect 2895 2058 2901 2059
rect 2946 2059 2947 2060
rect 2951 2059 2952 2063
rect 2946 2058 2952 2059
rect 3047 2063 3053 2064
rect 3047 2059 3048 2063
rect 3052 2062 3053 2063
rect 3098 2063 3104 2064
rect 3098 2062 3099 2063
rect 3052 2060 3099 2062
rect 3052 2059 3053 2060
rect 3047 2058 3053 2059
rect 3098 2059 3099 2060
rect 3103 2059 3104 2063
rect 3098 2058 3104 2059
rect 3191 2063 3197 2064
rect 3191 2059 3192 2063
rect 3196 2062 3197 2063
rect 3242 2063 3248 2064
rect 3242 2062 3243 2063
rect 3196 2060 3243 2062
rect 3196 2059 3197 2060
rect 3191 2058 3197 2059
rect 3242 2059 3243 2060
rect 3247 2059 3248 2063
rect 3242 2058 3248 2059
rect 3334 2063 3341 2064
rect 3334 2059 3335 2063
rect 3340 2059 3341 2063
rect 3334 2058 3341 2059
rect 3470 2063 3476 2064
rect 3470 2059 3471 2063
rect 3475 2062 3476 2063
rect 3487 2063 3493 2064
rect 3487 2062 3488 2063
rect 3475 2060 3488 2062
rect 3475 2059 3476 2060
rect 3470 2058 3476 2059
rect 3487 2059 3488 2060
rect 3492 2059 3493 2063
rect 3487 2058 3493 2059
rect 326 2055 332 2056
rect 326 2051 327 2055
rect 331 2051 332 2055
rect 326 2050 332 2051
rect 430 2055 436 2056
rect 430 2051 431 2055
rect 435 2051 436 2055
rect 430 2050 436 2051
rect 534 2055 540 2056
rect 534 2051 535 2055
rect 539 2051 540 2055
rect 534 2050 540 2051
rect 638 2055 644 2056
rect 638 2051 639 2055
rect 643 2051 644 2055
rect 638 2050 644 2051
rect 742 2055 748 2056
rect 742 2051 743 2055
rect 747 2051 748 2055
rect 742 2050 748 2051
rect 838 2055 844 2056
rect 838 2051 839 2055
rect 843 2051 844 2055
rect 838 2050 844 2051
rect 934 2055 940 2056
rect 934 2051 935 2055
rect 939 2051 940 2055
rect 934 2050 940 2051
rect 1038 2055 1044 2056
rect 1038 2051 1039 2055
rect 1043 2051 1044 2055
rect 1038 2050 1044 2051
rect 1142 2055 1148 2056
rect 1142 2051 1143 2055
rect 1147 2051 1148 2055
rect 1142 2050 1148 2051
rect 1246 2055 1252 2056
rect 1246 2051 1247 2055
rect 1251 2051 1252 2055
rect 1246 2050 1252 2051
rect 335 2043 344 2044
rect 335 2039 336 2043
rect 343 2039 344 2043
rect 335 2038 344 2039
rect 415 2043 421 2044
rect 415 2039 416 2043
rect 420 2042 421 2043
rect 439 2043 445 2044
rect 439 2042 440 2043
rect 420 2040 440 2042
rect 420 2039 421 2040
rect 415 2038 421 2039
rect 439 2039 440 2040
rect 444 2039 445 2043
rect 439 2038 445 2039
rect 543 2043 549 2044
rect 543 2039 544 2043
rect 548 2042 549 2043
rect 599 2043 605 2044
rect 599 2042 600 2043
rect 548 2040 600 2042
rect 548 2039 549 2040
rect 543 2038 549 2039
rect 599 2039 600 2040
rect 604 2039 605 2043
rect 599 2038 605 2039
rect 647 2043 653 2044
rect 647 2039 648 2043
rect 652 2042 653 2043
rect 703 2043 709 2044
rect 703 2042 704 2043
rect 652 2040 704 2042
rect 652 2039 653 2040
rect 647 2038 653 2039
rect 703 2039 704 2040
rect 708 2039 709 2043
rect 703 2038 709 2039
rect 751 2043 757 2044
rect 751 2039 752 2043
rect 756 2042 757 2043
rect 790 2043 796 2044
rect 790 2042 791 2043
rect 756 2040 791 2042
rect 756 2039 757 2040
rect 751 2038 757 2039
rect 790 2039 791 2040
rect 795 2039 796 2043
rect 790 2038 796 2039
rect 847 2043 856 2044
rect 847 2039 848 2043
rect 855 2039 856 2043
rect 847 2038 856 2039
rect 919 2043 925 2044
rect 919 2039 920 2043
rect 924 2042 925 2043
rect 943 2043 949 2044
rect 943 2042 944 2043
rect 924 2040 944 2042
rect 924 2039 925 2040
rect 919 2038 925 2039
rect 943 2039 944 2040
rect 948 2039 949 2043
rect 943 2038 949 2039
rect 1023 2043 1029 2044
rect 1023 2039 1024 2043
rect 1028 2042 1029 2043
rect 1047 2043 1053 2044
rect 1047 2042 1048 2043
rect 1028 2040 1048 2042
rect 1028 2039 1029 2040
rect 1023 2038 1029 2039
rect 1047 2039 1048 2040
rect 1052 2039 1053 2043
rect 1047 2038 1053 2039
rect 1127 2043 1133 2044
rect 1127 2039 1128 2043
rect 1132 2042 1133 2043
rect 1151 2043 1157 2044
rect 1151 2042 1152 2043
rect 1132 2040 1152 2042
rect 1132 2039 1133 2040
rect 1127 2038 1133 2039
rect 1151 2039 1152 2040
rect 1156 2039 1157 2043
rect 1151 2038 1157 2039
rect 1206 2043 1212 2044
rect 1206 2039 1207 2043
rect 1211 2042 1212 2043
rect 1255 2043 1261 2044
rect 1255 2042 1256 2043
rect 1211 2040 1256 2042
rect 1211 2039 1212 2040
rect 1206 2038 1212 2039
rect 1255 2039 1256 2040
rect 1260 2039 1261 2043
rect 1255 2038 1261 2039
rect 1903 2043 1909 2044
rect 1903 2039 1904 2043
rect 1908 2042 1909 2043
rect 1958 2043 1964 2044
rect 1908 2040 1954 2042
rect 1908 2039 1909 2040
rect 1903 2038 1909 2039
rect 1894 2033 1900 2034
rect 1214 2031 1220 2032
rect 1214 2030 1215 2031
rect 1068 2028 1215 2030
rect 223 2023 229 2024
rect 223 2019 224 2023
rect 228 2022 229 2023
rect 287 2023 293 2024
rect 287 2022 288 2023
rect 228 2020 288 2022
rect 228 2019 229 2020
rect 223 2018 229 2019
rect 287 2019 288 2020
rect 292 2019 293 2023
rect 287 2018 293 2019
rect 399 2023 405 2024
rect 399 2019 400 2023
rect 404 2022 405 2023
rect 407 2023 413 2024
rect 407 2022 408 2023
rect 404 2020 408 2022
rect 404 2019 405 2020
rect 399 2018 405 2019
rect 407 2019 408 2020
rect 412 2019 413 2023
rect 407 2018 413 2019
rect 567 2023 573 2024
rect 567 2019 568 2023
rect 572 2022 573 2023
rect 614 2023 620 2024
rect 614 2022 615 2023
rect 572 2020 615 2022
rect 572 2019 573 2020
rect 567 2018 573 2019
rect 614 2019 615 2020
rect 619 2019 620 2023
rect 614 2018 620 2019
rect 650 2023 656 2024
rect 650 2019 651 2023
rect 655 2022 656 2023
rect 727 2023 733 2024
rect 727 2022 728 2023
rect 655 2020 728 2022
rect 655 2019 656 2020
rect 650 2018 656 2019
rect 727 2019 728 2020
rect 732 2019 733 2023
rect 727 2018 733 2019
rect 782 2023 788 2024
rect 782 2019 783 2023
rect 787 2022 788 2023
rect 871 2023 877 2024
rect 871 2022 872 2023
rect 787 2020 872 2022
rect 787 2019 788 2020
rect 782 2018 788 2019
rect 871 2019 872 2020
rect 876 2019 877 2023
rect 871 2018 877 2019
rect 1007 2023 1013 2024
rect 1007 2019 1008 2023
rect 1012 2022 1013 2023
rect 1068 2022 1070 2028
rect 1214 2027 1215 2028
rect 1219 2027 1220 2031
rect 1894 2029 1895 2033
rect 1899 2029 1900 2033
rect 1894 2028 1900 2029
rect 1952 2030 1954 2040
rect 1958 2039 1959 2043
rect 1963 2042 1964 2043
rect 2023 2043 2029 2044
rect 2023 2042 2024 2043
rect 1963 2040 2024 2042
rect 1963 2039 1964 2040
rect 1958 2038 1964 2039
rect 2023 2039 2024 2040
rect 2028 2039 2029 2043
rect 2023 2038 2029 2039
rect 2090 2043 2096 2044
rect 2090 2039 2091 2043
rect 2095 2042 2096 2043
rect 2159 2043 2165 2044
rect 2159 2042 2160 2043
rect 2095 2040 2160 2042
rect 2095 2039 2096 2040
rect 2090 2038 2096 2039
rect 2159 2039 2160 2040
rect 2164 2039 2165 2043
rect 2159 2038 2165 2039
rect 2303 2043 2309 2044
rect 2303 2039 2304 2043
rect 2308 2042 2309 2043
rect 2362 2043 2368 2044
rect 2362 2042 2363 2043
rect 2308 2040 2363 2042
rect 2308 2039 2309 2040
rect 2303 2038 2309 2039
rect 2362 2039 2363 2040
rect 2367 2039 2368 2043
rect 2362 2038 2368 2039
rect 2447 2043 2456 2044
rect 2447 2039 2448 2043
rect 2455 2039 2456 2043
rect 2447 2038 2456 2039
rect 2599 2043 2605 2044
rect 2599 2039 2600 2043
rect 2604 2042 2605 2043
rect 2618 2043 2624 2044
rect 2618 2042 2619 2043
rect 2604 2040 2619 2042
rect 2604 2039 2605 2040
rect 2599 2038 2605 2039
rect 2618 2039 2619 2040
rect 2623 2039 2624 2043
rect 2618 2038 2624 2039
rect 2682 2043 2688 2044
rect 2682 2039 2683 2043
rect 2687 2042 2688 2043
rect 2767 2043 2773 2044
rect 2767 2042 2768 2043
rect 2687 2040 2768 2042
rect 2687 2039 2688 2040
rect 2682 2038 2688 2039
rect 2767 2039 2768 2040
rect 2772 2039 2773 2043
rect 2767 2038 2773 2039
rect 2870 2043 2876 2044
rect 2870 2039 2871 2043
rect 2875 2042 2876 2043
rect 2943 2043 2949 2044
rect 2943 2042 2944 2043
rect 2875 2040 2944 2042
rect 2875 2039 2876 2040
rect 2870 2038 2876 2039
rect 2943 2039 2944 2040
rect 2948 2039 2949 2043
rect 2943 2038 2949 2039
rect 3031 2043 3037 2044
rect 3031 2039 3032 2043
rect 3036 2042 3037 2043
rect 3127 2043 3133 2044
rect 3127 2042 3128 2043
rect 3036 2040 3128 2042
rect 3036 2039 3037 2040
rect 3031 2038 3037 2039
rect 3127 2039 3128 2040
rect 3132 2039 3133 2043
rect 3127 2038 3133 2039
rect 3222 2043 3228 2044
rect 3222 2039 3223 2043
rect 3227 2042 3228 2043
rect 3319 2043 3325 2044
rect 3319 2042 3320 2043
rect 3227 2040 3320 2042
rect 3227 2039 3228 2040
rect 3222 2038 3228 2039
rect 3319 2039 3320 2040
rect 3324 2039 3325 2043
rect 3319 2038 3325 2039
rect 3495 2043 3504 2044
rect 3495 2039 3496 2043
rect 3503 2039 3504 2043
rect 3495 2038 3504 2039
rect 2014 2033 2020 2034
rect 2006 2031 2012 2032
rect 2006 2030 2007 2031
rect 1952 2028 2007 2030
rect 1214 2026 1220 2027
rect 2006 2027 2007 2028
rect 2011 2027 2012 2031
rect 2014 2029 2015 2033
rect 2019 2029 2020 2033
rect 2014 2028 2020 2029
rect 2150 2033 2156 2034
rect 2150 2029 2151 2033
rect 2155 2029 2156 2033
rect 2150 2028 2156 2029
rect 2294 2033 2300 2034
rect 2294 2029 2295 2033
rect 2299 2029 2300 2033
rect 2294 2028 2300 2029
rect 2438 2033 2444 2034
rect 2438 2029 2439 2033
rect 2443 2029 2444 2033
rect 2438 2028 2444 2029
rect 2590 2033 2596 2034
rect 2590 2029 2591 2033
rect 2595 2029 2596 2033
rect 2590 2028 2596 2029
rect 2758 2033 2764 2034
rect 2758 2029 2759 2033
rect 2763 2029 2764 2033
rect 2758 2028 2764 2029
rect 2934 2033 2940 2034
rect 2934 2029 2935 2033
rect 2939 2029 2940 2033
rect 2934 2028 2940 2029
rect 3118 2033 3124 2034
rect 3118 2029 3119 2033
rect 3123 2029 3124 2033
rect 3118 2028 3124 2029
rect 3310 2033 3316 2034
rect 3310 2029 3311 2033
rect 3315 2029 3316 2033
rect 3310 2028 3316 2029
rect 3486 2033 3492 2034
rect 3486 2029 3487 2033
rect 3491 2029 3492 2033
rect 3486 2028 3492 2029
rect 2006 2026 2012 2027
rect 1012 2020 1070 2022
rect 1074 2023 1080 2024
rect 1012 2019 1013 2020
rect 1007 2018 1013 2019
rect 1074 2019 1075 2023
rect 1079 2022 1080 2023
rect 1135 2023 1141 2024
rect 1135 2022 1136 2023
rect 1079 2020 1136 2022
rect 1079 2019 1080 2020
rect 1074 2018 1080 2019
rect 1135 2019 1136 2020
rect 1140 2019 1141 2023
rect 1135 2018 1141 2019
rect 1215 2023 1221 2024
rect 1215 2019 1216 2023
rect 1220 2022 1221 2023
rect 1255 2023 1261 2024
rect 1255 2022 1256 2023
rect 1220 2020 1256 2022
rect 1220 2019 1221 2020
rect 1215 2018 1221 2019
rect 1255 2019 1256 2020
rect 1260 2019 1261 2023
rect 1255 2018 1261 2019
rect 1318 2023 1324 2024
rect 1318 2019 1319 2023
rect 1323 2022 1324 2023
rect 1375 2023 1381 2024
rect 1375 2022 1376 2023
rect 1323 2020 1376 2022
rect 1323 2019 1324 2020
rect 1318 2018 1324 2019
rect 1375 2019 1376 2020
rect 1380 2019 1381 2023
rect 1375 2018 1381 2019
rect 1442 2023 1448 2024
rect 1442 2019 1443 2023
rect 1447 2022 1448 2023
rect 1503 2023 1509 2024
rect 1503 2022 1504 2023
rect 1447 2020 1504 2022
rect 1447 2019 1448 2020
rect 1442 2018 1448 2019
rect 1503 2019 1504 2020
rect 1508 2019 1509 2023
rect 1503 2018 1509 2019
rect 1862 2020 1868 2021
rect 3574 2020 3580 2021
rect 1862 2016 1863 2020
rect 1867 2016 1868 2020
rect 1958 2019 1964 2020
rect 1958 2018 1959 2019
rect 1949 2016 1959 2018
rect 1862 2015 1868 2016
rect 1958 2015 1959 2016
rect 1963 2015 1964 2019
rect 2090 2019 2096 2020
rect 2090 2018 2091 2019
rect 2069 2016 2091 2018
rect 1958 2014 1964 2015
rect 2090 2015 2091 2016
rect 2095 2015 2096 2019
rect 2214 2019 2220 2020
rect 2214 2018 2215 2019
rect 2205 2016 2215 2018
rect 2090 2014 2096 2015
rect 2214 2015 2215 2016
rect 2219 2015 2220 2019
rect 2682 2019 2688 2020
rect 2682 2018 2683 2019
rect 2645 2016 2683 2018
rect 2214 2014 2220 2015
rect 2222 2015 2228 2016
rect 214 2013 220 2014
rect 214 2009 215 2013
rect 219 2009 220 2013
rect 214 2008 220 2009
rect 390 2013 396 2014
rect 390 2009 391 2013
rect 395 2009 396 2013
rect 390 2008 396 2009
rect 558 2013 564 2014
rect 558 2009 559 2013
rect 563 2009 564 2013
rect 558 2008 564 2009
rect 718 2013 724 2014
rect 718 2009 719 2013
rect 723 2009 724 2013
rect 718 2008 724 2009
rect 862 2013 868 2014
rect 862 2009 863 2013
rect 867 2009 868 2013
rect 862 2008 868 2009
rect 998 2013 1004 2014
rect 998 2009 999 2013
rect 1003 2009 1004 2013
rect 998 2008 1004 2009
rect 1126 2013 1132 2014
rect 1126 2009 1127 2013
rect 1131 2009 1132 2013
rect 1126 2008 1132 2009
rect 1246 2013 1252 2014
rect 1246 2009 1247 2013
rect 1251 2009 1252 2013
rect 1246 2008 1252 2009
rect 1366 2013 1372 2014
rect 1366 2009 1367 2013
rect 1371 2009 1372 2013
rect 1366 2008 1372 2009
rect 1494 2013 1500 2014
rect 1494 2009 1495 2013
rect 1499 2009 1500 2013
rect 2222 2011 2223 2015
rect 2227 2014 2228 2015
rect 2362 2015 2368 2016
rect 2227 2012 2313 2014
rect 2227 2011 2228 2012
rect 2222 2010 2228 2011
rect 2362 2011 2363 2015
rect 2367 2014 2368 2015
rect 2682 2015 2683 2016
rect 2687 2015 2688 2019
rect 2870 2019 2876 2020
rect 2870 2018 2871 2019
rect 2813 2016 2871 2018
rect 2682 2014 2688 2015
rect 2870 2015 2871 2016
rect 2875 2015 2876 2019
rect 3031 2019 3037 2020
rect 3031 2018 3032 2019
rect 2989 2016 3032 2018
rect 2870 2014 2876 2015
rect 3031 2015 3032 2016
rect 3036 2015 3037 2019
rect 3222 2019 3228 2020
rect 3222 2018 3223 2019
rect 3173 2016 3223 2018
rect 3031 2014 3037 2015
rect 3222 2015 3223 2016
rect 3227 2015 3228 2019
rect 3574 2016 3575 2020
rect 3579 2016 3580 2020
rect 3574 2015 3580 2016
rect 3222 2014 3228 2015
rect 2367 2012 2457 2014
rect 2367 2011 2368 2012
rect 2362 2010 2368 2011
rect 1494 2008 1500 2009
rect 1862 2003 1868 2004
rect 110 2000 116 2001
rect 1822 2000 1828 2001
rect 110 1996 111 2000
rect 115 1996 116 2000
rect 650 1999 656 2000
rect 650 1998 651 1999
rect 613 1996 651 1998
rect 110 1995 116 1996
rect 287 1995 293 1996
rect 287 1991 288 1995
rect 292 1994 293 1995
rect 650 1995 651 1996
rect 655 1995 656 1999
rect 782 1999 788 2000
rect 782 1998 783 1999
rect 773 1996 783 1998
rect 650 1994 656 1995
rect 782 1995 783 1996
rect 787 1995 788 1999
rect 1074 1999 1080 2000
rect 1074 1998 1075 1999
rect 1053 1996 1075 1998
rect 782 1994 788 1995
rect 790 1995 796 1996
rect 292 1992 409 1994
rect 292 1991 293 1992
rect 287 1990 293 1991
rect 790 1991 791 1995
rect 795 1994 796 1995
rect 1074 1995 1075 1996
rect 1079 1995 1080 1999
rect 1215 1999 1221 2000
rect 1215 1998 1216 1999
rect 1181 1996 1216 1998
rect 1074 1994 1080 1995
rect 1215 1995 1216 1996
rect 1220 1995 1221 1999
rect 1318 1999 1324 2000
rect 1318 1998 1319 1999
rect 1301 1996 1319 1998
rect 1215 1994 1221 1995
rect 1318 1995 1319 1996
rect 1323 1995 1324 1999
rect 1442 1999 1448 2000
rect 1442 1998 1443 1999
rect 1421 1996 1443 1998
rect 1318 1994 1324 1995
rect 1442 1995 1443 1996
rect 1447 1995 1448 1999
rect 1822 1996 1823 2000
rect 1827 1996 1828 2000
rect 1862 1999 1863 2003
rect 1867 1999 1868 2003
rect 1862 1998 1868 1999
rect 3310 2003 3316 2004
rect 3310 1999 3311 2003
rect 3315 2002 3316 2003
rect 3574 2003 3580 2004
rect 3315 2000 3321 2002
rect 3315 1999 3316 2000
rect 3310 1998 3316 1999
rect 3574 1999 3575 2003
rect 3579 1999 3580 2003
rect 3574 1998 3580 1999
rect 1822 1995 1828 1996
rect 1442 1994 1448 1995
rect 795 1992 881 1994
rect 1886 1993 1892 1994
rect 795 1991 796 1992
rect 790 1990 796 1991
rect 1886 1989 1887 1993
rect 1891 1989 1892 1993
rect 1886 1988 1892 1989
rect 2006 1993 2012 1994
rect 2006 1989 2007 1993
rect 2011 1989 2012 1993
rect 2006 1988 2012 1989
rect 2142 1993 2148 1994
rect 2142 1989 2143 1993
rect 2147 1989 2148 1993
rect 2142 1988 2148 1989
rect 2286 1993 2292 1994
rect 2286 1989 2287 1993
rect 2291 1989 2292 1993
rect 2286 1988 2292 1989
rect 2430 1993 2436 1994
rect 2430 1989 2431 1993
rect 2435 1989 2436 1993
rect 2430 1988 2436 1989
rect 2582 1993 2588 1994
rect 2582 1989 2583 1993
rect 2587 1989 2588 1993
rect 2582 1988 2588 1989
rect 2750 1993 2756 1994
rect 2750 1989 2751 1993
rect 2755 1989 2756 1993
rect 2750 1988 2756 1989
rect 2926 1993 2932 1994
rect 2926 1989 2927 1993
rect 2931 1989 2932 1993
rect 2926 1988 2932 1989
rect 3110 1993 3116 1994
rect 3110 1989 3111 1993
rect 3115 1989 3116 1993
rect 3110 1988 3116 1989
rect 3302 1993 3308 1994
rect 3302 1989 3303 1993
rect 3307 1989 3308 1993
rect 3302 1988 3308 1989
rect 3478 1993 3484 1994
rect 3478 1989 3479 1993
rect 3483 1989 3484 1993
rect 3478 1988 3484 1989
rect 3526 1987 3533 1988
rect 110 1983 116 1984
rect 110 1979 111 1983
rect 115 1979 116 1983
rect 110 1978 116 1979
rect 154 1983 160 1984
rect 154 1979 155 1983
rect 159 1982 160 1983
rect 1822 1983 1828 1984
rect 159 1980 225 1982
rect 1428 1980 1505 1982
rect 159 1979 160 1980
rect 154 1978 160 1979
rect 206 1973 212 1974
rect 206 1969 207 1973
rect 211 1969 212 1973
rect 206 1968 212 1969
rect 382 1973 388 1974
rect 382 1969 383 1973
rect 387 1969 388 1973
rect 382 1968 388 1969
rect 550 1973 556 1974
rect 550 1969 551 1973
rect 555 1969 556 1973
rect 550 1968 556 1969
rect 710 1973 716 1974
rect 710 1969 711 1973
rect 715 1969 716 1973
rect 710 1968 716 1969
rect 854 1973 860 1974
rect 854 1969 855 1973
rect 859 1969 860 1973
rect 854 1968 860 1969
rect 990 1973 996 1974
rect 990 1969 991 1973
rect 995 1969 996 1973
rect 990 1968 996 1969
rect 1118 1973 1124 1974
rect 1118 1969 1119 1973
rect 1123 1969 1124 1973
rect 1118 1968 1124 1969
rect 1238 1973 1244 1974
rect 1238 1969 1239 1973
rect 1243 1969 1244 1973
rect 1238 1968 1244 1969
rect 1358 1973 1364 1974
rect 1358 1969 1359 1973
rect 1363 1969 1364 1973
rect 1358 1968 1364 1969
rect 1134 1967 1140 1968
rect 1134 1963 1135 1967
rect 1139 1966 1140 1967
rect 1428 1966 1430 1980
rect 1822 1979 1823 1983
rect 1827 1979 1828 1983
rect 3526 1983 3527 1987
rect 3532 1983 3533 1987
rect 3526 1982 3533 1983
rect 1822 1978 1828 1979
rect 1486 1973 1492 1974
rect 1486 1969 1487 1973
rect 1491 1969 1492 1973
rect 1486 1968 1492 1969
rect 1139 1964 1430 1966
rect 2022 1967 2028 1968
rect 1139 1963 1140 1964
rect 1134 1962 1140 1963
rect 2022 1963 2023 1967
rect 2027 1963 2028 1967
rect 2022 1962 2028 1963
rect 2110 1967 2116 1968
rect 2110 1963 2111 1967
rect 2115 1963 2116 1967
rect 2110 1962 2116 1963
rect 2198 1967 2204 1968
rect 2198 1963 2199 1967
rect 2203 1963 2204 1967
rect 2198 1962 2204 1963
rect 2286 1967 2292 1968
rect 2286 1963 2287 1967
rect 2291 1963 2292 1967
rect 2286 1962 2292 1963
rect 2382 1967 2388 1968
rect 2382 1963 2383 1967
rect 2387 1963 2388 1967
rect 2382 1962 2388 1963
rect 2502 1967 2508 1968
rect 2502 1963 2503 1967
rect 2507 1963 2508 1967
rect 2502 1962 2508 1963
rect 2654 1967 2660 1968
rect 2654 1963 2655 1967
rect 2659 1963 2660 1967
rect 2654 1962 2660 1963
rect 2838 1967 2844 1968
rect 2838 1963 2839 1967
rect 2843 1963 2844 1967
rect 2838 1962 2844 1963
rect 3046 1967 3052 1968
rect 3046 1963 3047 1967
rect 3051 1963 3052 1967
rect 3046 1962 3052 1963
rect 3270 1967 3276 1968
rect 3270 1963 3271 1967
rect 3275 1963 3276 1967
rect 3270 1962 3276 1963
rect 3478 1967 3484 1968
rect 3478 1963 3479 1967
rect 3483 1963 3484 1967
rect 3478 1962 3484 1963
rect 2450 1959 2456 1960
rect 2450 1958 2451 1959
rect 1862 1957 1868 1958
rect 1862 1953 1863 1957
rect 1867 1953 1868 1957
rect 2441 1956 2451 1958
rect 2450 1955 2451 1956
rect 2455 1955 2456 1959
rect 2450 1954 2456 1955
rect 2570 1959 2576 1960
rect 2570 1955 2571 1959
rect 2575 1958 2576 1959
rect 2575 1956 2673 1958
rect 3574 1957 3580 1958
rect 2575 1955 2576 1956
rect 2570 1954 2576 1955
rect 1862 1952 1868 1953
rect 3574 1953 3575 1957
rect 3579 1953 3580 1957
rect 3574 1952 3580 1953
rect 134 1943 140 1944
rect 134 1939 135 1943
rect 139 1939 140 1943
rect 134 1938 140 1939
rect 310 1943 316 1944
rect 310 1939 311 1943
rect 315 1939 316 1943
rect 310 1938 316 1939
rect 518 1943 524 1944
rect 518 1939 519 1943
rect 523 1939 524 1943
rect 518 1938 524 1939
rect 718 1943 724 1944
rect 718 1939 719 1943
rect 723 1939 724 1943
rect 718 1938 724 1939
rect 910 1943 916 1944
rect 910 1939 911 1943
rect 915 1939 916 1943
rect 910 1938 916 1939
rect 1094 1943 1100 1944
rect 1094 1939 1095 1943
rect 1099 1939 1100 1943
rect 1094 1938 1100 1939
rect 1262 1943 1268 1944
rect 1262 1939 1263 1943
rect 1267 1939 1268 1943
rect 1262 1938 1268 1939
rect 1422 1943 1428 1944
rect 1422 1939 1423 1943
rect 1427 1939 1428 1943
rect 1422 1938 1428 1939
rect 1582 1943 1588 1944
rect 1582 1939 1583 1943
rect 1587 1939 1588 1943
rect 1582 1938 1588 1939
rect 1726 1943 1732 1944
rect 1726 1939 1727 1943
rect 1731 1939 1732 1943
rect 2103 1943 2109 1944
rect 2103 1942 2104 1943
rect 1726 1938 1732 1939
rect 1862 1940 1868 1941
rect 2085 1940 2104 1942
rect 1862 1936 1863 1940
rect 1867 1936 1868 1940
rect 2103 1939 2104 1940
rect 2108 1939 2109 1943
rect 2191 1943 2197 1944
rect 2191 1942 2192 1943
rect 2173 1940 2192 1942
rect 2103 1938 2109 1939
rect 2191 1939 2192 1940
rect 2196 1939 2197 1943
rect 2279 1943 2285 1944
rect 2279 1942 2280 1943
rect 2261 1940 2280 1942
rect 2191 1938 2197 1939
rect 2279 1939 2280 1940
rect 2284 1939 2285 1943
rect 2375 1943 2381 1944
rect 2375 1942 2376 1943
rect 2349 1940 2376 1942
rect 2279 1938 2285 1939
rect 2375 1939 2376 1940
rect 2380 1939 2381 1943
rect 2646 1943 2652 1944
rect 2646 1942 2647 1943
rect 2565 1940 2647 1942
rect 2375 1938 2381 1939
rect 2646 1939 2647 1940
rect 2651 1939 2652 1943
rect 2646 1938 2652 1939
rect 2722 1943 2728 1944
rect 2722 1939 2723 1943
rect 2727 1942 2728 1943
rect 2906 1943 2912 1944
rect 2727 1940 2865 1942
rect 2727 1939 2728 1940
rect 2722 1938 2728 1939
rect 2906 1939 2907 1943
rect 2911 1942 2912 1943
rect 3114 1943 3120 1944
rect 2911 1940 3073 1942
rect 2911 1939 2912 1940
rect 2906 1938 2912 1939
rect 3114 1939 3115 1943
rect 3119 1942 3120 1943
rect 3471 1943 3477 1944
rect 3119 1940 3297 1942
rect 3119 1939 3120 1940
rect 3114 1938 3120 1939
rect 3471 1939 3472 1943
rect 3476 1942 3477 1943
rect 3476 1940 3505 1942
rect 3574 1940 3580 1941
rect 3476 1939 3477 1940
rect 3471 1938 3477 1939
rect 378 1935 384 1936
rect 110 1933 116 1934
rect 110 1929 111 1933
rect 115 1929 116 1933
rect 378 1931 379 1935
rect 383 1934 384 1935
rect 614 1935 620 1936
rect 383 1932 537 1934
rect 383 1931 384 1932
rect 378 1930 384 1931
rect 614 1931 615 1935
rect 619 1934 620 1935
rect 1718 1935 1724 1936
rect 1862 1935 1868 1936
rect 3574 1936 3575 1940
rect 3579 1936 3580 1940
rect 3574 1935 3580 1936
rect 619 1932 737 1934
rect 619 1931 620 1932
rect 614 1930 620 1931
rect 1718 1931 1719 1935
rect 1723 1934 1724 1935
rect 1723 1932 1745 1934
rect 1822 1933 1828 1934
rect 1723 1931 1724 1932
rect 1718 1930 1724 1931
rect 110 1928 116 1929
rect 1822 1929 1823 1933
rect 1827 1929 1828 1933
rect 1822 1928 1828 1929
rect 2030 1927 2036 1928
rect 2030 1923 2031 1927
rect 2035 1923 2036 1927
rect 2030 1922 2036 1923
rect 2118 1927 2124 1928
rect 2118 1923 2119 1927
rect 2123 1923 2124 1927
rect 2118 1922 2124 1923
rect 2206 1927 2212 1928
rect 2206 1923 2207 1927
rect 2211 1923 2212 1927
rect 2206 1922 2212 1923
rect 2294 1927 2300 1928
rect 2294 1923 2295 1927
rect 2299 1923 2300 1927
rect 2294 1922 2300 1923
rect 2390 1927 2396 1928
rect 2390 1923 2391 1927
rect 2395 1923 2396 1927
rect 2390 1922 2396 1923
rect 2510 1927 2516 1928
rect 2510 1923 2511 1927
rect 2515 1923 2516 1927
rect 2510 1922 2516 1923
rect 2662 1927 2668 1928
rect 2662 1923 2663 1927
rect 2667 1923 2668 1927
rect 2662 1922 2668 1923
rect 2846 1927 2852 1928
rect 2846 1923 2847 1927
rect 2851 1923 2852 1927
rect 2846 1922 2852 1923
rect 3054 1927 3060 1928
rect 3054 1923 3055 1927
rect 3059 1923 3060 1927
rect 3054 1922 3060 1923
rect 3278 1927 3284 1928
rect 3278 1923 3279 1927
rect 3283 1923 3284 1927
rect 3278 1922 3284 1923
rect 3486 1927 3492 1928
rect 3486 1923 3487 1927
rect 3491 1923 3492 1927
rect 3486 1922 3492 1923
rect 242 1919 248 1920
rect 242 1918 243 1919
rect 110 1916 116 1917
rect 197 1916 243 1918
rect 110 1912 111 1916
rect 115 1912 116 1916
rect 242 1915 243 1916
rect 247 1915 248 1919
rect 511 1919 517 1920
rect 511 1918 512 1919
rect 373 1916 512 1918
rect 242 1914 248 1915
rect 511 1915 512 1916
rect 516 1915 517 1919
rect 511 1914 517 1915
rect 786 1919 792 1920
rect 786 1915 787 1919
rect 791 1918 792 1919
rect 1255 1919 1261 1920
rect 1255 1918 1256 1919
rect 791 1916 937 1918
rect 1157 1916 1256 1918
rect 791 1915 792 1916
rect 786 1914 792 1915
rect 1255 1915 1256 1916
rect 1260 1915 1261 1919
rect 1415 1919 1421 1920
rect 1415 1918 1416 1919
rect 1325 1916 1416 1918
rect 1255 1914 1261 1915
rect 1415 1915 1416 1916
rect 1420 1915 1421 1919
rect 1575 1919 1581 1920
rect 1575 1918 1576 1919
rect 1485 1916 1576 1918
rect 1415 1914 1421 1915
rect 1575 1915 1576 1916
rect 1580 1915 1581 1919
rect 1719 1919 1725 1920
rect 1719 1918 1720 1919
rect 1645 1916 1720 1918
rect 1575 1914 1581 1915
rect 1719 1915 1720 1916
rect 1724 1915 1725 1919
rect 1719 1914 1725 1915
rect 1822 1916 1828 1917
rect 110 1911 116 1912
rect 1822 1912 1823 1916
rect 1827 1912 1828 1916
rect 1822 1911 1828 1912
rect 2039 1915 2048 1916
rect 2039 1911 2040 1915
rect 2047 1911 2048 1915
rect 2039 1910 2048 1911
rect 2103 1915 2109 1916
rect 2103 1911 2104 1915
rect 2108 1914 2109 1915
rect 2127 1915 2133 1916
rect 2127 1914 2128 1915
rect 2108 1912 2128 1914
rect 2108 1911 2109 1912
rect 2103 1910 2109 1911
rect 2127 1911 2128 1912
rect 2132 1911 2133 1915
rect 2127 1910 2133 1911
rect 2191 1915 2197 1916
rect 2191 1911 2192 1915
rect 2196 1914 2197 1915
rect 2215 1915 2221 1916
rect 2215 1914 2216 1915
rect 2196 1912 2216 1914
rect 2196 1911 2197 1912
rect 2191 1910 2197 1911
rect 2215 1911 2216 1912
rect 2220 1911 2221 1915
rect 2215 1910 2221 1911
rect 2279 1915 2285 1916
rect 2279 1911 2280 1915
rect 2284 1914 2285 1915
rect 2303 1915 2309 1916
rect 2303 1914 2304 1915
rect 2284 1912 2304 1914
rect 2284 1911 2285 1912
rect 2279 1910 2285 1911
rect 2303 1911 2304 1912
rect 2308 1911 2309 1915
rect 2303 1910 2309 1911
rect 2375 1915 2381 1916
rect 2375 1911 2376 1915
rect 2380 1914 2381 1915
rect 2399 1915 2405 1916
rect 2399 1914 2400 1915
rect 2380 1912 2400 1914
rect 2380 1911 2381 1912
rect 2375 1910 2381 1911
rect 2399 1911 2400 1912
rect 2404 1911 2405 1915
rect 2399 1910 2405 1911
rect 2519 1915 2525 1916
rect 2519 1911 2520 1915
rect 2524 1914 2525 1915
rect 2570 1915 2576 1916
rect 2570 1914 2571 1915
rect 2524 1912 2571 1914
rect 2524 1911 2525 1912
rect 2519 1910 2525 1911
rect 2570 1911 2571 1912
rect 2575 1911 2576 1915
rect 2570 1910 2576 1911
rect 2671 1915 2677 1916
rect 2671 1911 2672 1915
rect 2676 1914 2677 1915
rect 2722 1915 2728 1916
rect 2722 1914 2723 1915
rect 2676 1912 2723 1914
rect 2676 1911 2677 1912
rect 2671 1910 2677 1911
rect 2722 1911 2723 1912
rect 2727 1911 2728 1915
rect 2722 1910 2728 1911
rect 2855 1915 2861 1916
rect 2855 1911 2856 1915
rect 2860 1914 2861 1915
rect 2906 1915 2912 1916
rect 2906 1914 2907 1915
rect 2860 1912 2907 1914
rect 2860 1911 2861 1912
rect 2855 1910 2861 1911
rect 2906 1911 2907 1912
rect 2911 1911 2912 1915
rect 2906 1910 2912 1911
rect 3063 1915 3069 1916
rect 3063 1911 3064 1915
rect 3068 1914 3069 1915
rect 3114 1915 3120 1916
rect 3114 1914 3115 1915
rect 3068 1912 3115 1914
rect 3068 1911 3069 1912
rect 3063 1910 3069 1911
rect 3114 1911 3115 1912
rect 3119 1911 3120 1915
rect 3114 1910 3120 1911
rect 3287 1915 3293 1916
rect 3287 1911 3288 1915
rect 3292 1914 3293 1915
rect 3310 1915 3316 1916
rect 3310 1914 3311 1915
rect 3292 1912 3311 1914
rect 3292 1911 3293 1912
rect 3287 1910 3293 1911
rect 3310 1911 3311 1912
rect 3315 1911 3316 1915
rect 3310 1910 3316 1911
rect 3495 1915 3501 1916
rect 3495 1911 3496 1915
rect 3500 1914 3501 1915
rect 3526 1915 3532 1916
rect 3526 1914 3527 1915
rect 3500 1912 3527 1914
rect 3500 1911 3501 1912
rect 3495 1910 3501 1911
rect 3526 1911 3527 1912
rect 3531 1911 3532 1915
rect 3526 1910 3532 1911
rect 142 1903 148 1904
rect 142 1899 143 1903
rect 147 1899 148 1903
rect 142 1898 148 1899
rect 318 1903 324 1904
rect 318 1899 319 1903
rect 323 1899 324 1903
rect 318 1898 324 1899
rect 526 1903 532 1904
rect 526 1899 527 1903
rect 531 1899 532 1903
rect 526 1898 532 1899
rect 726 1903 732 1904
rect 726 1899 727 1903
rect 731 1899 732 1903
rect 726 1898 732 1899
rect 918 1903 924 1904
rect 918 1899 919 1903
rect 923 1899 924 1903
rect 918 1898 924 1899
rect 1102 1903 1108 1904
rect 1102 1899 1103 1903
rect 1107 1899 1108 1903
rect 1102 1898 1108 1899
rect 1270 1903 1276 1904
rect 1270 1899 1271 1903
rect 1275 1899 1276 1903
rect 1270 1898 1276 1899
rect 1430 1903 1436 1904
rect 1430 1899 1431 1903
rect 1435 1899 1436 1903
rect 1430 1898 1436 1899
rect 1590 1903 1596 1904
rect 1590 1899 1591 1903
rect 1595 1899 1596 1903
rect 1590 1898 1596 1899
rect 1734 1903 1740 1904
rect 1734 1899 1735 1903
rect 1739 1899 1740 1903
rect 1734 1898 1740 1899
rect 2183 1895 2189 1896
rect 151 1891 160 1892
rect 151 1887 152 1891
rect 159 1887 160 1891
rect 151 1886 160 1887
rect 242 1891 248 1892
rect 242 1887 243 1891
rect 247 1890 248 1891
rect 327 1891 333 1892
rect 327 1890 328 1891
rect 247 1888 328 1890
rect 247 1887 248 1888
rect 242 1886 248 1887
rect 327 1887 328 1888
rect 332 1887 333 1891
rect 327 1886 333 1887
rect 511 1891 517 1892
rect 511 1887 512 1891
rect 516 1890 517 1891
rect 535 1891 541 1892
rect 535 1890 536 1891
rect 516 1888 536 1890
rect 516 1887 517 1888
rect 511 1886 517 1887
rect 535 1887 536 1888
rect 540 1887 541 1891
rect 535 1886 541 1887
rect 735 1891 741 1892
rect 735 1887 736 1891
rect 740 1890 741 1891
rect 786 1891 792 1892
rect 786 1890 787 1891
rect 740 1888 787 1890
rect 740 1887 741 1888
rect 735 1886 741 1887
rect 786 1887 787 1888
rect 791 1887 792 1891
rect 786 1886 792 1887
rect 927 1891 933 1892
rect 927 1887 928 1891
rect 932 1890 933 1891
rect 946 1891 952 1892
rect 946 1890 947 1891
rect 932 1888 947 1890
rect 932 1887 933 1888
rect 927 1886 933 1887
rect 946 1887 947 1888
rect 951 1887 952 1891
rect 946 1886 952 1887
rect 1111 1891 1117 1892
rect 1111 1887 1112 1891
rect 1116 1890 1117 1891
rect 1134 1891 1140 1892
rect 1134 1890 1135 1891
rect 1116 1888 1135 1890
rect 1116 1887 1117 1888
rect 1111 1886 1117 1887
rect 1134 1887 1135 1888
rect 1139 1887 1140 1891
rect 1134 1886 1140 1887
rect 1255 1891 1261 1892
rect 1255 1887 1256 1891
rect 1260 1890 1261 1891
rect 1279 1891 1285 1892
rect 1279 1890 1280 1891
rect 1260 1888 1280 1890
rect 1260 1887 1261 1888
rect 1255 1886 1261 1887
rect 1279 1887 1280 1888
rect 1284 1887 1285 1891
rect 1279 1886 1285 1887
rect 1415 1891 1421 1892
rect 1415 1887 1416 1891
rect 1420 1890 1421 1891
rect 1439 1891 1445 1892
rect 1439 1890 1440 1891
rect 1420 1888 1440 1890
rect 1420 1887 1421 1888
rect 1415 1886 1421 1887
rect 1439 1887 1440 1888
rect 1444 1887 1445 1891
rect 1439 1886 1445 1887
rect 1575 1891 1581 1892
rect 1575 1887 1576 1891
rect 1580 1890 1581 1891
rect 1599 1891 1605 1892
rect 1599 1890 1600 1891
rect 1580 1888 1600 1890
rect 1580 1887 1581 1888
rect 1575 1886 1581 1887
rect 1599 1887 1600 1888
rect 1604 1887 1605 1891
rect 1599 1886 1605 1887
rect 1719 1891 1725 1892
rect 1719 1887 1720 1891
rect 1724 1890 1725 1891
rect 1743 1891 1749 1892
rect 1743 1890 1744 1891
rect 1724 1888 1744 1890
rect 1724 1887 1725 1888
rect 1719 1886 1725 1887
rect 1743 1887 1744 1888
rect 1748 1887 1749 1891
rect 2183 1891 2184 1895
rect 2188 1894 2189 1895
rect 2242 1895 2248 1896
rect 2242 1894 2243 1895
rect 2188 1892 2243 1894
rect 2188 1891 2189 1892
rect 2183 1890 2189 1891
rect 2242 1891 2243 1892
rect 2247 1891 2248 1895
rect 2242 1890 2248 1891
rect 2271 1895 2277 1896
rect 2271 1891 2272 1895
rect 2276 1894 2277 1895
rect 2330 1895 2336 1896
rect 2330 1894 2331 1895
rect 2276 1892 2331 1894
rect 2276 1891 2277 1892
rect 2271 1890 2277 1891
rect 2330 1891 2331 1892
rect 2335 1891 2336 1895
rect 2330 1890 2336 1891
rect 2359 1895 2365 1896
rect 2359 1891 2360 1895
rect 2364 1894 2365 1895
rect 2418 1895 2424 1896
rect 2418 1894 2419 1895
rect 2364 1892 2419 1894
rect 2364 1891 2365 1892
rect 2359 1890 2365 1891
rect 2418 1891 2419 1892
rect 2423 1891 2424 1895
rect 2418 1890 2424 1891
rect 2447 1895 2453 1896
rect 2447 1891 2448 1895
rect 2452 1894 2453 1895
rect 2511 1895 2517 1896
rect 2511 1894 2512 1895
rect 2452 1892 2512 1894
rect 2452 1891 2453 1892
rect 2447 1890 2453 1891
rect 2511 1891 2512 1892
rect 2516 1891 2517 1895
rect 2511 1890 2517 1891
rect 2534 1895 2541 1896
rect 2534 1891 2535 1895
rect 2540 1891 2541 1895
rect 2534 1890 2541 1891
rect 2646 1895 2653 1896
rect 2646 1891 2647 1895
rect 2652 1891 2653 1895
rect 2646 1890 2653 1891
rect 2711 1895 2717 1896
rect 2711 1891 2712 1895
rect 2716 1894 2717 1895
rect 2783 1895 2789 1896
rect 2783 1894 2784 1895
rect 2716 1892 2784 1894
rect 2716 1891 2717 1892
rect 2711 1890 2717 1891
rect 2783 1891 2784 1892
rect 2788 1891 2789 1895
rect 2783 1890 2789 1891
rect 2890 1895 2896 1896
rect 2890 1891 2891 1895
rect 2895 1894 2896 1895
rect 2943 1895 2949 1896
rect 2943 1894 2944 1895
rect 2895 1892 2944 1894
rect 2895 1891 2896 1892
rect 2890 1890 2896 1891
rect 2943 1891 2944 1892
rect 2948 1891 2949 1895
rect 2943 1890 2949 1891
rect 3031 1895 3037 1896
rect 3031 1891 3032 1895
rect 3036 1894 3037 1895
rect 3127 1895 3133 1896
rect 3127 1894 3128 1895
rect 3036 1892 3128 1894
rect 3036 1891 3037 1892
rect 3031 1890 3037 1891
rect 3127 1891 3128 1892
rect 3132 1891 3133 1895
rect 3127 1890 3133 1891
rect 3223 1895 3229 1896
rect 3223 1891 3224 1895
rect 3228 1894 3229 1895
rect 3319 1895 3325 1896
rect 3319 1894 3320 1895
rect 3228 1892 3320 1894
rect 3228 1891 3229 1892
rect 3223 1890 3229 1891
rect 3319 1891 3320 1892
rect 3324 1891 3325 1895
rect 3319 1890 3325 1891
rect 3471 1895 3477 1896
rect 3471 1891 3472 1895
rect 3476 1894 3477 1895
rect 3495 1895 3501 1896
rect 3495 1894 3496 1895
rect 3476 1892 3496 1894
rect 3476 1891 3477 1892
rect 3471 1890 3477 1891
rect 3495 1891 3496 1892
rect 3500 1891 3501 1895
rect 3495 1890 3501 1891
rect 1743 1886 1749 1887
rect 2174 1885 2180 1886
rect 2174 1881 2175 1885
rect 2179 1881 2180 1885
rect 2174 1880 2180 1881
rect 2262 1885 2268 1886
rect 2262 1881 2263 1885
rect 2267 1881 2268 1885
rect 2262 1880 2268 1881
rect 2350 1885 2356 1886
rect 2350 1881 2351 1885
rect 2355 1881 2356 1885
rect 2350 1880 2356 1881
rect 2438 1885 2444 1886
rect 2438 1881 2439 1885
rect 2443 1881 2444 1885
rect 2438 1880 2444 1881
rect 2526 1885 2532 1886
rect 2526 1881 2527 1885
rect 2531 1881 2532 1885
rect 2526 1880 2532 1881
rect 2638 1885 2644 1886
rect 2638 1881 2639 1885
rect 2643 1881 2644 1885
rect 2638 1880 2644 1881
rect 2774 1885 2780 1886
rect 2774 1881 2775 1885
rect 2779 1881 2780 1885
rect 2774 1880 2780 1881
rect 2934 1885 2940 1886
rect 2934 1881 2935 1885
rect 2939 1881 2940 1885
rect 2934 1880 2940 1881
rect 3118 1885 3124 1886
rect 3118 1881 3119 1885
rect 3123 1881 3124 1885
rect 3118 1880 3124 1881
rect 3310 1885 3316 1886
rect 3310 1881 3311 1885
rect 3315 1881 3316 1885
rect 3310 1880 3316 1881
rect 3486 1885 3492 1886
rect 3486 1881 3487 1885
rect 3491 1881 3492 1885
rect 3486 1880 3492 1881
rect 1862 1872 1868 1873
rect 3574 1872 3580 1873
rect 151 1871 157 1872
rect 151 1867 152 1871
rect 156 1870 157 1871
rect 234 1871 240 1872
rect 234 1870 235 1871
rect 156 1868 235 1870
rect 156 1867 157 1868
rect 151 1866 157 1867
rect 234 1867 235 1868
rect 239 1867 240 1871
rect 234 1866 240 1867
rect 319 1871 325 1872
rect 319 1867 320 1871
rect 324 1870 325 1871
rect 378 1871 384 1872
rect 378 1870 379 1871
rect 324 1868 379 1870
rect 324 1867 325 1868
rect 319 1866 325 1867
rect 378 1867 379 1868
rect 383 1867 384 1871
rect 378 1866 384 1867
rect 519 1871 525 1872
rect 519 1867 520 1871
rect 524 1870 525 1871
rect 615 1871 621 1872
rect 524 1868 610 1870
rect 524 1867 525 1868
rect 519 1866 525 1867
rect 608 1862 610 1868
rect 615 1867 616 1871
rect 620 1870 621 1871
rect 711 1871 717 1872
rect 711 1870 712 1871
rect 620 1868 712 1870
rect 620 1867 621 1868
rect 615 1866 621 1867
rect 711 1867 712 1868
rect 716 1867 717 1871
rect 711 1866 717 1867
rect 799 1871 805 1872
rect 799 1867 800 1871
rect 804 1870 805 1871
rect 895 1871 901 1872
rect 895 1870 896 1871
rect 804 1868 896 1870
rect 804 1867 805 1868
rect 799 1866 805 1867
rect 895 1867 896 1868
rect 900 1867 901 1871
rect 895 1866 901 1867
rect 1071 1871 1077 1872
rect 1071 1867 1072 1871
rect 1076 1870 1077 1871
rect 1134 1871 1140 1872
rect 1134 1870 1135 1871
rect 1076 1868 1135 1870
rect 1076 1867 1077 1868
rect 1071 1866 1077 1867
rect 1134 1867 1135 1868
rect 1139 1867 1140 1871
rect 1134 1866 1140 1867
rect 1143 1871 1149 1872
rect 1143 1867 1144 1871
rect 1148 1870 1149 1871
rect 1239 1871 1245 1872
rect 1239 1870 1240 1871
rect 1148 1868 1240 1870
rect 1148 1867 1149 1868
rect 1143 1866 1149 1867
rect 1239 1867 1240 1868
rect 1244 1867 1245 1871
rect 1239 1866 1245 1867
rect 1399 1871 1405 1872
rect 1399 1867 1400 1871
rect 1404 1870 1405 1871
rect 1479 1871 1485 1872
rect 1479 1870 1480 1871
rect 1404 1868 1480 1870
rect 1404 1867 1405 1868
rect 1399 1866 1405 1867
rect 1479 1867 1480 1868
rect 1484 1867 1485 1871
rect 1479 1866 1485 1867
rect 1559 1871 1565 1872
rect 1559 1867 1560 1871
rect 1564 1870 1565 1871
rect 1639 1871 1645 1872
rect 1639 1870 1640 1871
rect 1564 1868 1640 1870
rect 1564 1867 1565 1868
rect 1559 1866 1565 1867
rect 1639 1867 1640 1868
rect 1644 1867 1645 1871
rect 1639 1866 1645 1867
rect 1718 1871 1725 1872
rect 1718 1867 1719 1871
rect 1724 1867 1725 1871
rect 1862 1868 1863 1872
rect 1867 1868 1868 1872
rect 2711 1871 2717 1872
rect 2711 1870 2712 1871
rect 2693 1868 2712 1870
rect 1862 1867 1868 1868
rect 2042 1867 2048 1868
rect 1718 1866 1725 1867
rect 634 1863 640 1864
rect 634 1862 635 1863
rect 142 1861 148 1862
rect 142 1857 143 1861
rect 147 1857 148 1861
rect 142 1856 148 1857
rect 310 1861 316 1862
rect 310 1857 311 1861
rect 315 1857 316 1861
rect 310 1856 316 1857
rect 510 1861 516 1862
rect 510 1857 511 1861
rect 515 1857 516 1861
rect 608 1860 635 1862
rect 634 1859 635 1860
rect 639 1859 640 1863
rect 2042 1863 2043 1867
rect 2047 1866 2048 1867
rect 2242 1867 2248 1868
rect 2047 1864 2193 1866
rect 2047 1863 2048 1864
rect 2042 1862 2048 1863
rect 2242 1863 2243 1867
rect 2247 1866 2248 1867
rect 2330 1867 2336 1868
rect 2247 1864 2281 1866
rect 2247 1863 2248 1864
rect 2242 1862 2248 1863
rect 2330 1863 2331 1867
rect 2335 1866 2336 1867
rect 2418 1867 2424 1868
rect 2335 1864 2369 1866
rect 2335 1863 2336 1864
rect 2330 1862 2336 1863
rect 2418 1863 2419 1867
rect 2423 1866 2424 1867
rect 2511 1867 2517 1868
rect 2423 1864 2457 1866
rect 2423 1863 2424 1864
rect 2418 1862 2424 1863
rect 2511 1863 2512 1867
rect 2516 1866 2517 1867
rect 2711 1867 2712 1868
rect 2716 1867 2717 1871
rect 2890 1871 2896 1872
rect 2890 1870 2891 1871
rect 2829 1868 2891 1870
rect 2711 1866 2717 1867
rect 2890 1867 2891 1868
rect 2895 1867 2896 1871
rect 3031 1871 3037 1872
rect 3031 1870 3032 1871
rect 2989 1868 3032 1870
rect 2890 1866 2896 1867
rect 3031 1867 3032 1868
rect 3036 1867 3037 1871
rect 3223 1871 3229 1872
rect 3223 1870 3224 1871
rect 3173 1868 3224 1870
rect 3031 1866 3037 1867
rect 3223 1867 3224 1868
rect 3228 1867 3229 1871
rect 3574 1868 3575 1872
rect 3579 1868 3580 1872
rect 3574 1867 3580 1868
rect 3223 1866 3229 1867
rect 2516 1864 2545 1866
rect 2516 1863 2517 1864
rect 2511 1862 2517 1863
rect 634 1858 640 1859
rect 702 1861 708 1862
rect 510 1856 516 1857
rect 702 1857 703 1861
rect 707 1857 708 1861
rect 702 1856 708 1857
rect 886 1861 892 1862
rect 886 1857 887 1861
rect 891 1857 892 1861
rect 886 1856 892 1857
rect 1062 1861 1068 1862
rect 1062 1857 1063 1861
rect 1067 1857 1068 1861
rect 1062 1856 1068 1857
rect 1230 1861 1236 1862
rect 1230 1857 1231 1861
rect 1235 1857 1236 1861
rect 1230 1856 1236 1857
rect 1390 1861 1396 1862
rect 1390 1857 1391 1861
rect 1395 1857 1396 1861
rect 1390 1856 1396 1857
rect 1550 1861 1556 1862
rect 1550 1857 1551 1861
rect 1555 1857 1556 1861
rect 1550 1856 1556 1857
rect 1710 1861 1716 1862
rect 1710 1857 1711 1861
rect 1715 1857 1716 1861
rect 1710 1856 1716 1857
rect 1862 1855 1868 1856
rect 1862 1851 1863 1855
rect 1867 1851 1868 1855
rect 1862 1850 1868 1851
rect 3198 1855 3204 1856
rect 3198 1851 3199 1855
rect 3203 1854 3204 1855
rect 3574 1855 3580 1856
rect 3203 1852 3321 1854
rect 3203 1851 3204 1852
rect 3198 1850 3204 1851
rect 3574 1851 3575 1855
rect 3579 1851 3580 1855
rect 3574 1850 3580 1851
rect 110 1848 116 1849
rect 1822 1848 1828 1849
rect 110 1844 111 1848
rect 115 1844 116 1848
rect 615 1847 621 1848
rect 615 1846 616 1847
rect 565 1844 616 1846
rect 110 1843 116 1844
rect 234 1843 240 1844
rect 234 1839 235 1843
rect 239 1842 240 1843
rect 615 1843 616 1844
rect 620 1843 621 1847
rect 799 1847 805 1848
rect 799 1846 800 1847
rect 757 1844 800 1846
rect 615 1842 621 1843
rect 799 1843 800 1844
rect 804 1843 805 1847
rect 946 1847 952 1848
rect 946 1846 947 1847
rect 941 1844 947 1846
rect 799 1842 805 1843
rect 946 1843 947 1844
rect 951 1843 952 1847
rect 1143 1847 1149 1848
rect 1143 1846 1144 1847
rect 1117 1844 1144 1846
rect 946 1842 952 1843
rect 1143 1843 1144 1844
rect 1148 1843 1149 1847
rect 1822 1844 1823 1848
rect 1827 1844 1828 1848
rect 1143 1842 1149 1843
rect 1298 1843 1304 1844
rect 239 1840 329 1842
rect 239 1839 240 1840
rect 234 1838 240 1839
rect 1298 1839 1299 1843
rect 1303 1842 1304 1843
rect 1479 1843 1485 1844
rect 1303 1840 1409 1842
rect 1303 1839 1304 1840
rect 1298 1838 1304 1839
rect 1479 1839 1480 1843
rect 1484 1842 1485 1843
rect 1639 1843 1645 1844
rect 1822 1843 1828 1844
rect 2166 1845 2172 1846
rect 1484 1840 1569 1842
rect 1484 1839 1485 1840
rect 1479 1838 1485 1839
rect 1639 1839 1640 1843
rect 1644 1842 1645 1843
rect 1644 1840 1729 1842
rect 2166 1841 2167 1845
rect 2171 1841 2172 1845
rect 2166 1840 2172 1841
rect 2254 1845 2260 1846
rect 2254 1841 2255 1845
rect 2259 1841 2260 1845
rect 2254 1840 2260 1841
rect 2342 1845 2348 1846
rect 2342 1841 2343 1845
rect 2347 1841 2348 1845
rect 2342 1840 2348 1841
rect 2430 1845 2436 1846
rect 2430 1841 2431 1845
rect 2435 1841 2436 1845
rect 2430 1840 2436 1841
rect 2518 1845 2524 1846
rect 2518 1841 2519 1845
rect 2523 1841 2524 1845
rect 2518 1840 2524 1841
rect 2630 1845 2636 1846
rect 2630 1841 2631 1845
rect 2635 1841 2636 1845
rect 2630 1840 2636 1841
rect 2766 1845 2772 1846
rect 2766 1841 2767 1845
rect 2771 1841 2772 1845
rect 2766 1840 2772 1841
rect 2926 1845 2932 1846
rect 2926 1841 2927 1845
rect 2931 1841 2932 1845
rect 2926 1840 2932 1841
rect 3110 1845 3116 1846
rect 3110 1841 3111 1845
rect 3115 1841 3116 1845
rect 3110 1840 3116 1841
rect 3302 1845 3308 1846
rect 3302 1841 3303 1845
rect 3307 1841 3308 1845
rect 3302 1840 3308 1841
rect 3478 1845 3484 1846
rect 3478 1841 3479 1845
rect 3483 1841 3484 1845
rect 3478 1840 3484 1841
rect 1644 1839 1645 1840
rect 1639 1838 1645 1839
rect 3498 1839 3504 1840
rect 3498 1835 3499 1839
rect 3503 1838 3504 1839
rect 3527 1839 3533 1840
rect 3527 1838 3528 1839
rect 3503 1836 3528 1838
rect 3503 1835 3504 1836
rect 3498 1834 3504 1835
rect 3527 1835 3528 1836
rect 3532 1835 3533 1839
rect 3527 1834 3533 1835
rect 110 1831 116 1832
rect 110 1827 111 1831
rect 115 1827 116 1831
rect 1298 1831 1304 1832
rect 1298 1830 1299 1831
rect 1281 1828 1299 1830
rect 110 1826 116 1827
rect 1298 1827 1299 1828
rect 1303 1827 1304 1831
rect 1298 1826 1304 1827
rect 1822 1831 1828 1832
rect 1822 1827 1823 1831
rect 1827 1827 1828 1831
rect 1822 1826 1828 1827
rect 134 1821 140 1822
rect 134 1817 135 1821
rect 139 1817 140 1821
rect 134 1816 140 1817
rect 302 1821 308 1822
rect 302 1817 303 1821
rect 307 1817 308 1821
rect 302 1816 308 1817
rect 502 1821 508 1822
rect 502 1817 503 1821
rect 507 1817 508 1821
rect 502 1816 508 1817
rect 694 1821 700 1822
rect 694 1817 695 1821
rect 699 1817 700 1821
rect 694 1816 700 1817
rect 878 1821 884 1822
rect 878 1817 879 1821
rect 883 1817 884 1821
rect 878 1816 884 1817
rect 1054 1821 1060 1822
rect 1054 1817 1055 1821
rect 1059 1817 1060 1821
rect 1054 1816 1060 1817
rect 1222 1821 1228 1822
rect 1222 1817 1223 1821
rect 1227 1817 1228 1821
rect 1222 1816 1228 1817
rect 1382 1821 1388 1822
rect 1382 1817 1383 1821
rect 1387 1817 1388 1821
rect 1382 1816 1388 1817
rect 1542 1821 1548 1822
rect 1542 1817 1543 1821
rect 1547 1817 1548 1821
rect 1542 1816 1548 1817
rect 1702 1821 1708 1822
rect 1702 1817 1703 1821
rect 1707 1817 1708 1821
rect 1702 1816 1708 1817
rect 2318 1819 2324 1820
rect 154 1815 160 1816
rect 154 1811 155 1815
rect 159 1814 160 1815
rect 183 1815 189 1816
rect 183 1814 184 1815
rect 159 1812 184 1814
rect 159 1811 160 1812
rect 154 1810 160 1811
rect 183 1811 184 1812
rect 188 1811 189 1815
rect 2318 1815 2319 1819
rect 2323 1815 2324 1819
rect 2318 1814 2324 1815
rect 2438 1819 2444 1820
rect 2438 1815 2439 1819
rect 2443 1815 2444 1819
rect 2438 1814 2444 1815
rect 2558 1819 2564 1820
rect 2558 1815 2559 1819
rect 2563 1815 2564 1819
rect 2558 1814 2564 1815
rect 2678 1819 2684 1820
rect 2678 1815 2679 1819
rect 2683 1815 2684 1819
rect 2678 1814 2684 1815
rect 2798 1819 2804 1820
rect 2798 1815 2799 1819
rect 2803 1815 2804 1819
rect 2798 1814 2804 1815
rect 2918 1819 2924 1820
rect 2918 1815 2919 1819
rect 2923 1815 2924 1819
rect 2918 1814 2924 1815
rect 3046 1819 3052 1820
rect 3046 1815 3047 1819
rect 3051 1815 3052 1819
rect 3046 1814 3052 1815
rect 3182 1819 3188 1820
rect 3182 1815 3183 1819
rect 3187 1815 3188 1819
rect 3182 1814 3188 1815
rect 3318 1819 3324 1820
rect 3318 1815 3319 1819
rect 3323 1815 3324 1819
rect 3318 1814 3324 1815
rect 3462 1819 3468 1820
rect 3462 1815 3463 1819
rect 3467 1815 3468 1819
rect 3462 1814 3468 1815
rect 183 1810 189 1811
rect 2534 1811 2540 1812
rect 2534 1810 2535 1811
rect 1862 1809 1868 1810
rect 1862 1805 1863 1809
rect 1867 1805 1868 1809
rect 2497 1808 2535 1810
rect 2534 1807 2535 1808
rect 2539 1807 2540 1811
rect 3472 1808 3481 1810
rect 3574 1809 3580 1810
rect 2534 1806 2540 1807
rect 3470 1807 3476 1808
rect 1862 1804 1868 1805
rect 3470 1803 3471 1807
rect 3475 1803 3476 1807
rect 3574 1805 3575 1809
rect 3579 1805 3580 1809
rect 3574 1804 3580 1805
rect 3470 1802 3476 1803
rect 2431 1795 2437 1796
rect 2431 1794 2432 1795
rect 1862 1792 1868 1793
rect 2381 1792 2432 1794
rect 134 1791 140 1792
rect 134 1787 135 1791
rect 139 1787 140 1791
rect 134 1786 140 1787
rect 262 1791 268 1792
rect 262 1787 263 1791
rect 267 1787 268 1791
rect 262 1786 268 1787
rect 414 1791 420 1792
rect 414 1787 415 1791
rect 419 1787 420 1791
rect 414 1786 420 1787
rect 566 1791 572 1792
rect 566 1787 567 1791
rect 571 1787 572 1791
rect 566 1786 572 1787
rect 718 1791 724 1792
rect 718 1787 719 1791
rect 723 1787 724 1791
rect 718 1786 724 1787
rect 862 1791 868 1792
rect 862 1787 863 1791
rect 867 1787 868 1791
rect 862 1786 868 1787
rect 1006 1791 1012 1792
rect 1006 1787 1007 1791
rect 1011 1787 1012 1791
rect 1006 1786 1012 1787
rect 1142 1791 1148 1792
rect 1142 1787 1143 1791
rect 1147 1787 1148 1791
rect 1142 1786 1148 1787
rect 1278 1791 1284 1792
rect 1278 1787 1279 1791
rect 1283 1787 1284 1791
rect 1278 1786 1284 1787
rect 1422 1791 1428 1792
rect 1422 1787 1423 1791
rect 1427 1787 1428 1791
rect 1862 1788 1863 1792
rect 1867 1788 1868 1792
rect 2431 1791 2432 1792
rect 2436 1791 2437 1795
rect 2431 1790 2437 1791
rect 2506 1795 2512 1796
rect 2506 1791 2507 1795
rect 2511 1794 2512 1795
rect 2626 1795 2632 1796
rect 2511 1792 2585 1794
rect 2511 1791 2512 1792
rect 2506 1790 2512 1791
rect 2626 1791 2627 1795
rect 2631 1794 2632 1795
rect 2911 1795 2917 1796
rect 2911 1794 2912 1795
rect 2631 1792 2705 1794
rect 2861 1792 2912 1794
rect 2631 1791 2632 1792
rect 2626 1790 2632 1791
rect 2911 1791 2912 1792
rect 2916 1791 2917 1795
rect 3039 1795 3045 1796
rect 3039 1794 3040 1795
rect 2981 1792 3040 1794
rect 2911 1790 2917 1791
rect 3039 1791 3040 1792
rect 3044 1791 3045 1795
rect 3175 1795 3181 1796
rect 3175 1794 3176 1795
rect 3109 1792 3176 1794
rect 3039 1790 3045 1791
rect 3175 1791 3176 1792
rect 3180 1791 3181 1795
rect 3311 1795 3317 1796
rect 3311 1794 3312 1795
rect 3245 1792 3312 1794
rect 3175 1790 3181 1791
rect 3311 1791 3312 1792
rect 3316 1791 3317 1795
rect 3390 1795 3396 1796
rect 3390 1794 3391 1795
rect 3381 1792 3391 1794
rect 3311 1790 3317 1791
rect 3390 1791 3391 1792
rect 3395 1791 3396 1795
rect 3390 1790 3396 1791
rect 3574 1792 3580 1793
rect 1862 1787 1868 1788
rect 3574 1788 3575 1792
rect 3579 1788 3580 1792
rect 3574 1787 3580 1788
rect 1422 1786 1428 1787
rect 634 1783 640 1784
rect 110 1781 116 1782
rect 110 1777 111 1781
rect 115 1777 116 1781
rect 634 1779 635 1783
rect 639 1782 640 1783
rect 1346 1783 1352 1784
rect 639 1780 737 1782
rect 639 1779 640 1780
rect 634 1778 640 1779
rect 1346 1779 1347 1783
rect 1351 1782 1352 1783
rect 1351 1780 1441 1782
rect 1822 1781 1828 1782
rect 1351 1779 1352 1780
rect 1346 1778 1352 1779
rect 110 1776 116 1777
rect 1822 1777 1823 1781
rect 1827 1777 1828 1781
rect 1822 1776 1828 1777
rect 2326 1779 2332 1780
rect 2326 1775 2327 1779
rect 2331 1775 2332 1779
rect 2326 1774 2332 1775
rect 2446 1779 2452 1780
rect 2446 1775 2447 1779
rect 2451 1775 2452 1779
rect 2446 1774 2452 1775
rect 2566 1779 2572 1780
rect 2566 1775 2567 1779
rect 2571 1775 2572 1779
rect 2566 1774 2572 1775
rect 2686 1779 2692 1780
rect 2686 1775 2687 1779
rect 2691 1775 2692 1779
rect 2686 1774 2692 1775
rect 2806 1779 2812 1780
rect 2806 1775 2807 1779
rect 2811 1775 2812 1779
rect 2806 1774 2812 1775
rect 2926 1779 2932 1780
rect 2926 1775 2927 1779
rect 2931 1775 2932 1779
rect 2926 1774 2932 1775
rect 3054 1779 3060 1780
rect 3054 1775 3055 1779
rect 3059 1775 3060 1779
rect 3054 1774 3060 1775
rect 3190 1779 3196 1780
rect 3190 1775 3191 1779
rect 3195 1775 3196 1779
rect 3190 1774 3196 1775
rect 3326 1779 3332 1780
rect 3326 1775 3327 1779
rect 3331 1775 3332 1779
rect 3326 1774 3332 1775
rect 3470 1779 3476 1780
rect 3470 1775 3471 1779
rect 3475 1775 3476 1779
rect 3470 1774 3476 1775
rect 255 1767 261 1768
rect 255 1766 256 1767
rect 110 1764 116 1765
rect 197 1764 256 1766
rect 110 1760 111 1764
rect 115 1760 116 1764
rect 255 1763 256 1764
rect 260 1763 261 1767
rect 330 1767 336 1768
rect 330 1766 331 1767
rect 325 1764 331 1766
rect 255 1762 261 1763
rect 330 1763 331 1764
rect 335 1763 336 1767
rect 559 1767 565 1768
rect 559 1766 560 1767
rect 477 1764 560 1766
rect 330 1762 336 1763
rect 559 1763 560 1764
rect 564 1763 565 1767
rect 711 1767 717 1768
rect 711 1766 712 1767
rect 629 1764 712 1766
rect 559 1762 565 1763
rect 711 1763 712 1764
rect 716 1763 717 1767
rect 711 1762 717 1763
rect 786 1767 792 1768
rect 786 1763 787 1767
rect 791 1766 792 1767
rect 930 1767 936 1768
rect 791 1764 889 1766
rect 791 1763 792 1764
rect 786 1762 792 1763
rect 930 1763 931 1767
rect 935 1766 936 1767
rect 1074 1767 1080 1768
rect 935 1764 1033 1766
rect 935 1763 936 1764
rect 930 1762 936 1763
rect 1074 1763 1075 1767
rect 1079 1766 1080 1767
rect 1415 1767 1421 1768
rect 1415 1766 1416 1767
rect 1079 1764 1169 1766
rect 1341 1764 1416 1766
rect 1079 1763 1080 1764
rect 1074 1762 1080 1763
rect 1415 1763 1416 1764
rect 1420 1763 1421 1767
rect 2335 1767 2341 1768
rect 1415 1762 1421 1763
rect 1822 1764 1828 1765
rect 110 1759 116 1760
rect 1822 1760 1823 1764
rect 1827 1760 1828 1764
rect 2335 1763 2336 1767
rect 2340 1766 2341 1767
rect 2431 1767 2437 1768
rect 2340 1764 2426 1766
rect 2340 1763 2341 1764
rect 2335 1762 2341 1763
rect 1822 1759 1828 1760
rect 2424 1758 2426 1764
rect 2431 1763 2432 1767
rect 2436 1766 2437 1767
rect 2455 1767 2461 1768
rect 2455 1766 2456 1767
rect 2436 1764 2456 1766
rect 2436 1763 2437 1764
rect 2431 1762 2437 1763
rect 2455 1763 2456 1764
rect 2460 1763 2461 1767
rect 2455 1762 2461 1763
rect 2575 1767 2581 1768
rect 2575 1763 2576 1767
rect 2580 1766 2581 1767
rect 2626 1767 2632 1768
rect 2626 1766 2627 1767
rect 2580 1764 2627 1766
rect 2580 1763 2581 1764
rect 2575 1762 2581 1763
rect 2626 1763 2627 1764
rect 2631 1763 2632 1767
rect 2626 1762 2632 1763
rect 2695 1767 2701 1768
rect 2695 1763 2696 1767
rect 2700 1766 2701 1767
rect 2722 1767 2728 1768
rect 2722 1766 2723 1767
rect 2700 1764 2723 1766
rect 2700 1763 2701 1764
rect 2695 1762 2701 1763
rect 2722 1763 2723 1764
rect 2727 1763 2728 1767
rect 2722 1762 2728 1763
rect 2815 1767 2824 1768
rect 2815 1763 2816 1767
rect 2823 1763 2824 1767
rect 2815 1762 2824 1763
rect 2911 1767 2917 1768
rect 2911 1763 2912 1767
rect 2916 1766 2917 1767
rect 2935 1767 2941 1768
rect 2935 1766 2936 1767
rect 2916 1764 2936 1766
rect 2916 1763 2917 1764
rect 2911 1762 2917 1763
rect 2935 1763 2936 1764
rect 2940 1763 2941 1767
rect 2935 1762 2941 1763
rect 3039 1767 3045 1768
rect 3039 1763 3040 1767
rect 3044 1766 3045 1767
rect 3063 1767 3069 1768
rect 3063 1766 3064 1767
rect 3044 1764 3064 1766
rect 3044 1763 3045 1764
rect 3039 1762 3045 1763
rect 3063 1763 3064 1764
rect 3068 1763 3069 1767
rect 3063 1762 3069 1763
rect 3175 1767 3181 1768
rect 3175 1763 3176 1767
rect 3180 1766 3181 1767
rect 3199 1767 3205 1768
rect 3199 1766 3200 1767
rect 3180 1764 3200 1766
rect 3180 1763 3181 1764
rect 3175 1762 3181 1763
rect 3199 1763 3200 1764
rect 3204 1763 3205 1767
rect 3199 1762 3205 1763
rect 3311 1767 3317 1768
rect 3311 1763 3312 1767
rect 3316 1766 3317 1767
rect 3335 1767 3341 1768
rect 3335 1766 3336 1767
rect 3316 1764 3336 1766
rect 3316 1763 3317 1764
rect 3311 1762 3317 1763
rect 3335 1763 3336 1764
rect 3340 1763 3341 1767
rect 3335 1762 3341 1763
rect 3462 1767 3468 1768
rect 3462 1763 3463 1767
rect 3467 1766 3468 1767
rect 3479 1767 3485 1768
rect 3479 1766 3480 1767
rect 3467 1764 3480 1766
rect 3467 1763 3468 1764
rect 3462 1762 3468 1763
rect 3479 1763 3480 1764
rect 3484 1763 3485 1767
rect 3479 1762 3485 1763
rect 2506 1759 2512 1760
rect 2506 1758 2507 1759
rect 2424 1756 2507 1758
rect 2506 1755 2507 1756
rect 2511 1755 2512 1759
rect 2506 1754 2512 1755
rect 3327 1755 3333 1756
rect 3327 1754 3328 1755
rect 3192 1752 3328 1754
rect 142 1751 148 1752
rect 142 1747 143 1751
rect 147 1747 148 1751
rect 142 1746 148 1747
rect 270 1751 276 1752
rect 270 1747 271 1751
rect 275 1747 276 1751
rect 270 1746 276 1747
rect 422 1751 428 1752
rect 422 1747 423 1751
rect 427 1747 428 1751
rect 422 1746 428 1747
rect 574 1751 580 1752
rect 574 1747 575 1751
rect 579 1747 580 1751
rect 574 1746 580 1747
rect 726 1751 732 1752
rect 726 1747 727 1751
rect 731 1747 732 1751
rect 726 1746 732 1747
rect 870 1751 876 1752
rect 870 1747 871 1751
rect 875 1747 876 1751
rect 870 1746 876 1747
rect 1014 1751 1020 1752
rect 1014 1747 1015 1751
rect 1019 1747 1020 1751
rect 1014 1746 1020 1747
rect 1150 1751 1156 1752
rect 1150 1747 1151 1751
rect 1155 1747 1156 1751
rect 1150 1746 1156 1747
rect 1286 1751 1292 1752
rect 1286 1747 1287 1751
rect 1291 1747 1292 1751
rect 1286 1746 1292 1747
rect 1430 1751 1436 1752
rect 1430 1747 1431 1751
rect 1435 1747 1436 1751
rect 1430 1746 1436 1747
rect 2303 1747 2312 1748
rect 2303 1743 2304 1747
rect 2311 1743 2312 1747
rect 2303 1742 2312 1743
rect 2359 1747 2365 1748
rect 2359 1743 2360 1747
rect 2364 1746 2365 1747
rect 2415 1747 2421 1748
rect 2415 1746 2416 1747
rect 2364 1744 2416 1746
rect 2364 1743 2365 1744
rect 2359 1742 2365 1743
rect 2415 1743 2416 1744
rect 2420 1743 2421 1747
rect 2415 1742 2421 1743
rect 2471 1747 2477 1748
rect 2471 1743 2472 1747
rect 2476 1746 2477 1747
rect 2535 1747 2541 1748
rect 2535 1746 2536 1747
rect 2476 1744 2536 1746
rect 2476 1743 2477 1744
rect 2471 1742 2477 1743
rect 2535 1743 2536 1744
rect 2540 1743 2541 1747
rect 2535 1742 2541 1743
rect 2599 1747 2605 1748
rect 2599 1743 2600 1747
rect 2604 1746 2605 1747
rect 2663 1747 2669 1748
rect 2663 1746 2664 1747
rect 2604 1744 2664 1746
rect 2604 1743 2605 1744
rect 2599 1742 2605 1743
rect 2663 1743 2664 1744
rect 2668 1743 2669 1747
rect 2663 1742 2669 1743
rect 2714 1747 2720 1748
rect 2714 1743 2715 1747
rect 2719 1746 2720 1747
rect 2783 1747 2789 1748
rect 2783 1746 2784 1747
rect 2719 1744 2784 1746
rect 2719 1743 2720 1744
rect 2714 1742 2720 1743
rect 2783 1743 2784 1744
rect 2788 1743 2789 1747
rect 2783 1742 2789 1743
rect 2903 1747 2909 1748
rect 2903 1743 2904 1747
rect 2908 1746 2909 1747
rect 2966 1747 2972 1748
rect 2966 1746 2967 1747
rect 2908 1744 2967 1746
rect 2908 1743 2909 1744
rect 2903 1742 2909 1743
rect 2966 1743 2967 1744
rect 2971 1743 2972 1747
rect 2966 1742 2972 1743
rect 3023 1747 3029 1748
rect 3023 1743 3024 1747
rect 3028 1746 3029 1747
rect 3042 1747 3048 1748
rect 3042 1746 3043 1747
rect 3028 1744 3043 1746
rect 3028 1743 3029 1744
rect 3023 1742 3029 1743
rect 3042 1743 3043 1744
rect 3047 1743 3048 1747
rect 3042 1742 3048 1743
rect 3143 1747 3149 1748
rect 3143 1743 3144 1747
rect 3148 1746 3149 1747
rect 3192 1746 3194 1752
rect 3327 1751 3328 1752
rect 3332 1751 3333 1755
rect 3327 1750 3333 1751
rect 3148 1744 3194 1746
rect 3199 1747 3205 1748
rect 3148 1743 3149 1744
rect 3143 1742 3149 1743
rect 3199 1743 3200 1747
rect 3204 1746 3205 1747
rect 3263 1747 3269 1748
rect 3263 1746 3264 1747
rect 3204 1744 3264 1746
rect 3204 1743 3205 1744
rect 3199 1742 3205 1743
rect 3263 1743 3264 1744
rect 3268 1743 3269 1747
rect 3263 1742 3269 1743
rect 3390 1747 3397 1748
rect 3390 1743 3391 1747
rect 3396 1743 3397 1747
rect 3390 1742 3397 1743
rect 3495 1747 3504 1748
rect 3495 1743 3496 1747
rect 3503 1743 3504 1747
rect 3495 1742 3504 1743
rect 151 1739 160 1740
rect 151 1735 152 1739
rect 159 1735 160 1739
rect 151 1734 160 1735
rect 255 1739 261 1740
rect 255 1735 256 1739
rect 260 1738 261 1739
rect 279 1739 285 1740
rect 279 1738 280 1739
rect 260 1736 280 1738
rect 260 1735 261 1736
rect 255 1734 261 1735
rect 279 1735 280 1736
rect 284 1735 285 1739
rect 279 1734 285 1735
rect 414 1739 420 1740
rect 414 1735 415 1739
rect 419 1738 420 1739
rect 431 1739 437 1740
rect 431 1738 432 1739
rect 419 1736 432 1738
rect 419 1735 420 1736
rect 414 1734 420 1735
rect 431 1735 432 1736
rect 436 1735 437 1739
rect 431 1734 437 1735
rect 559 1739 565 1740
rect 559 1735 560 1739
rect 564 1738 565 1739
rect 583 1739 589 1740
rect 583 1738 584 1739
rect 564 1736 584 1738
rect 564 1735 565 1736
rect 559 1734 565 1735
rect 583 1735 584 1736
rect 588 1735 589 1739
rect 583 1734 589 1735
rect 711 1739 717 1740
rect 711 1735 712 1739
rect 716 1738 717 1739
rect 735 1739 741 1740
rect 735 1738 736 1739
rect 716 1736 736 1738
rect 716 1735 717 1736
rect 711 1734 717 1735
rect 735 1735 736 1736
rect 740 1735 741 1739
rect 735 1734 741 1735
rect 879 1739 885 1740
rect 879 1735 880 1739
rect 884 1738 885 1739
rect 930 1739 936 1740
rect 930 1738 931 1739
rect 884 1736 931 1738
rect 884 1735 885 1736
rect 879 1734 885 1735
rect 930 1735 931 1736
rect 935 1735 936 1739
rect 930 1734 936 1735
rect 1023 1739 1029 1740
rect 1023 1735 1024 1739
rect 1028 1738 1029 1739
rect 1074 1739 1080 1740
rect 1074 1738 1075 1739
rect 1028 1736 1075 1738
rect 1028 1735 1029 1736
rect 1023 1734 1029 1735
rect 1074 1735 1075 1736
rect 1079 1735 1080 1739
rect 1074 1734 1080 1735
rect 1159 1739 1165 1740
rect 1159 1735 1160 1739
rect 1164 1738 1165 1739
rect 1295 1739 1304 1740
rect 1164 1736 1290 1738
rect 1164 1735 1165 1736
rect 1159 1734 1165 1735
rect 1288 1730 1290 1736
rect 1295 1735 1296 1739
rect 1303 1735 1304 1739
rect 1295 1734 1304 1735
rect 1415 1739 1421 1740
rect 1415 1735 1416 1739
rect 1420 1738 1421 1739
rect 1439 1739 1445 1740
rect 1439 1738 1440 1739
rect 1420 1736 1440 1738
rect 1420 1735 1421 1736
rect 1415 1734 1421 1735
rect 1439 1735 1440 1736
rect 1444 1735 1445 1739
rect 1439 1734 1445 1735
rect 2294 1737 2300 1738
rect 2294 1733 2295 1737
rect 2299 1733 2300 1737
rect 2294 1732 2300 1733
rect 2406 1737 2412 1738
rect 2406 1733 2407 1737
rect 2411 1733 2412 1737
rect 2406 1732 2412 1733
rect 2526 1737 2532 1738
rect 2526 1733 2527 1737
rect 2531 1733 2532 1737
rect 2526 1732 2532 1733
rect 2654 1737 2660 1738
rect 2654 1733 2655 1737
rect 2659 1733 2660 1737
rect 2654 1732 2660 1733
rect 2774 1737 2780 1738
rect 2774 1733 2775 1737
rect 2779 1733 2780 1737
rect 2774 1732 2780 1733
rect 2894 1737 2900 1738
rect 2894 1733 2895 1737
rect 2899 1733 2900 1737
rect 2894 1732 2900 1733
rect 3014 1737 3020 1738
rect 3014 1733 3015 1737
rect 3019 1733 3020 1737
rect 3014 1732 3020 1733
rect 3134 1737 3140 1738
rect 3134 1733 3135 1737
rect 3139 1733 3140 1737
rect 3134 1732 3140 1733
rect 3254 1737 3260 1738
rect 3254 1733 3255 1737
rect 3259 1733 3260 1737
rect 3254 1732 3260 1733
rect 3382 1737 3388 1738
rect 3382 1733 3383 1737
rect 3387 1733 3388 1737
rect 3382 1732 3388 1733
rect 3486 1737 3492 1738
rect 3486 1733 3487 1737
rect 3491 1733 3492 1737
rect 3486 1732 3492 1733
rect 1346 1731 1352 1732
rect 1346 1730 1347 1731
rect 1288 1728 1347 1730
rect 151 1727 157 1728
rect 151 1723 152 1727
rect 156 1726 157 1727
rect 218 1727 224 1728
rect 218 1726 219 1727
rect 156 1724 219 1726
rect 156 1723 157 1724
rect 151 1722 157 1723
rect 218 1723 219 1724
rect 223 1723 224 1727
rect 218 1722 224 1723
rect 287 1727 293 1728
rect 287 1723 288 1727
rect 292 1726 293 1727
rect 330 1727 336 1728
rect 330 1726 331 1727
rect 292 1724 331 1726
rect 292 1723 293 1724
rect 287 1722 293 1723
rect 330 1723 331 1724
rect 335 1723 336 1727
rect 330 1722 336 1723
rect 439 1727 445 1728
rect 439 1723 440 1727
rect 444 1726 445 1727
rect 498 1727 504 1728
rect 498 1726 499 1727
rect 444 1724 499 1726
rect 444 1723 445 1724
rect 439 1722 445 1723
rect 498 1723 499 1724
rect 503 1723 504 1727
rect 498 1722 504 1723
rect 567 1727 573 1728
rect 567 1723 568 1727
rect 572 1726 573 1727
rect 591 1727 597 1728
rect 591 1726 592 1727
rect 572 1724 592 1726
rect 572 1723 573 1724
rect 567 1722 573 1723
rect 591 1723 592 1724
rect 596 1723 597 1727
rect 591 1722 597 1723
rect 735 1727 741 1728
rect 735 1723 736 1727
rect 740 1726 741 1727
rect 786 1727 792 1728
rect 786 1726 787 1727
rect 740 1724 787 1726
rect 740 1723 741 1724
rect 735 1722 741 1723
rect 786 1723 787 1724
rect 791 1723 792 1727
rect 786 1722 792 1723
rect 799 1727 805 1728
rect 799 1723 800 1727
rect 804 1726 805 1727
rect 871 1727 877 1728
rect 871 1726 872 1727
rect 804 1724 872 1726
rect 804 1723 805 1724
rect 799 1722 805 1723
rect 871 1723 872 1724
rect 876 1723 877 1727
rect 871 1722 877 1723
rect 935 1727 941 1728
rect 935 1723 936 1727
rect 940 1726 941 1727
rect 999 1727 1005 1728
rect 999 1726 1000 1727
rect 940 1724 1000 1726
rect 940 1723 941 1724
rect 935 1722 941 1723
rect 999 1723 1000 1724
rect 1004 1723 1005 1727
rect 999 1722 1005 1723
rect 1063 1727 1069 1728
rect 1063 1723 1064 1727
rect 1068 1726 1069 1727
rect 1135 1727 1141 1728
rect 1135 1726 1136 1727
rect 1068 1724 1136 1726
rect 1068 1723 1069 1724
rect 1063 1722 1069 1723
rect 1135 1723 1136 1724
rect 1140 1723 1141 1727
rect 1135 1722 1141 1723
rect 1247 1727 1253 1728
rect 1247 1723 1248 1727
rect 1252 1726 1253 1727
rect 1271 1727 1277 1728
rect 1271 1726 1272 1727
rect 1252 1724 1272 1726
rect 1252 1723 1253 1724
rect 1247 1722 1253 1723
rect 1271 1723 1272 1724
rect 1276 1723 1277 1727
rect 1346 1727 1347 1728
rect 1351 1727 1352 1731
rect 1346 1726 1352 1727
rect 1271 1722 1277 1723
rect 1862 1724 1868 1725
rect 3574 1724 3580 1725
rect 1862 1720 1863 1724
rect 1867 1720 1868 1724
rect 2359 1723 2365 1724
rect 2359 1722 2360 1723
rect 2349 1720 2360 1722
rect 1862 1719 1868 1720
rect 2359 1719 2360 1720
rect 2364 1719 2365 1723
rect 2471 1723 2477 1724
rect 2471 1722 2472 1723
rect 2461 1720 2472 1722
rect 2359 1718 2365 1719
rect 2471 1719 2472 1720
rect 2476 1719 2477 1723
rect 2599 1723 2605 1724
rect 2599 1722 2600 1723
rect 2581 1720 2600 1722
rect 2471 1718 2477 1719
rect 2599 1719 2600 1720
rect 2604 1719 2605 1723
rect 2714 1723 2720 1724
rect 2714 1722 2715 1723
rect 2709 1720 2715 1722
rect 2599 1718 2605 1719
rect 2714 1719 2715 1720
rect 2719 1719 2720 1723
rect 3199 1723 3205 1724
rect 3199 1722 3200 1723
rect 3189 1720 3200 1722
rect 2714 1718 2720 1719
rect 2722 1719 2728 1720
rect 142 1717 148 1718
rect 142 1713 143 1717
rect 147 1713 148 1717
rect 142 1712 148 1713
rect 278 1717 284 1718
rect 278 1713 279 1717
rect 283 1713 284 1717
rect 278 1712 284 1713
rect 430 1717 436 1718
rect 430 1713 431 1717
rect 435 1713 436 1717
rect 430 1712 436 1713
rect 582 1717 588 1718
rect 582 1713 583 1717
rect 587 1713 588 1717
rect 582 1712 588 1713
rect 726 1717 732 1718
rect 726 1713 727 1717
rect 731 1713 732 1717
rect 726 1712 732 1713
rect 862 1717 868 1718
rect 862 1713 863 1717
rect 867 1713 868 1717
rect 862 1712 868 1713
rect 990 1717 996 1718
rect 990 1713 991 1717
rect 995 1713 996 1717
rect 990 1712 996 1713
rect 1126 1717 1132 1718
rect 1126 1713 1127 1717
rect 1131 1713 1132 1717
rect 1126 1712 1132 1713
rect 1262 1717 1268 1718
rect 1262 1713 1263 1717
rect 1267 1713 1268 1717
rect 2722 1715 2723 1719
rect 2727 1718 2728 1719
rect 2966 1719 2972 1720
rect 2727 1716 2793 1718
rect 2727 1715 2728 1716
rect 2722 1714 2728 1715
rect 2966 1715 2967 1719
rect 2971 1718 2972 1719
rect 3199 1719 3200 1720
rect 3204 1719 3205 1723
rect 3574 1720 3575 1724
rect 3579 1720 3580 1724
rect 3199 1718 3205 1719
rect 3327 1719 3333 1720
rect 3574 1719 3580 1720
rect 2971 1716 3033 1718
rect 2971 1715 2972 1716
rect 2966 1714 2972 1715
rect 3327 1715 3328 1719
rect 3332 1718 3333 1719
rect 3332 1716 3401 1718
rect 3332 1715 3333 1716
rect 3327 1714 3333 1715
rect 1262 1712 1268 1713
rect 1862 1707 1868 1708
rect 110 1704 116 1705
rect 1822 1704 1828 1705
rect 110 1700 111 1704
rect 115 1700 116 1704
rect 799 1703 805 1704
rect 799 1702 800 1703
rect 781 1700 800 1702
rect 110 1699 116 1700
rect 218 1699 224 1700
rect 218 1695 219 1699
rect 223 1698 224 1699
rect 414 1699 420 1700
rect 223 1696 297 1698
rect 223 1695 224 1696
rect 218 1694 224 1695
rect 414 1695 415 1699
rect 419 1698 420 1699
rect 498 1699 504 1700
rect 419 1696 449 1698
rect 419 1695 420 1696
rect 414 1694 420 1695
rect 498 1695 499 1699
rect 503 1698 504 1699
rect 799 1699 800 1700
rect 804 1699 805 1703
rect 935 1703 941 1704
rect 935 1702 936 1703
rect 917 1700 936 1702
rect 799 1698 805 1699
rect 935 1699 936 1700
rect 940 1699 941 1703
rect 1063 1703 1069 1704
rect 1063 1702 1064 1703
rect 1045 1700 1064 1702
rect 935 1698 941 1699
rect 1063 1699 1064 1700
rect 1068 1699 1069 1703
rect 1247 1703 1253 1704
rect 1247 1702 1248 1703
rect 1181 1700 1248 1702
rect 1063 1698 1069 1699
rect 1247 1699 1248 1700
rect 1252 1699 1253 1703
rect 1822 1700 1823 1704
rect 1827 1700 1828 1704
rect 1862 1703 1863 1707
rect 1867 1703 1868 1707
rect 1862 1702 1868 1703
rect 2854 1707 2860 1708
rect 2854 1703 2855 1707
rect 2859 1706 2860 1707
rect 3334 1707 3340 1708
rect 3334 1706 3335 1707
rect 2859 1704 2905 1706
rect 3305 1704 3335 1706
rect 2859 1703 2860 1704
rect 2854 1702 2860 1703
rect 3334 1703 3335 1704
rect 3339 1703 3340 1707
rect 3334 1702 3340 1703
rect 3574 1707 3580 1708
rect 3574 1703 3575 1707
rect 3579 1703 3580 1707
rect 3574 1702 3580 1703
rect 1822 1699 1828 1700
rect 1247 1698 1253 1699
rect 503 1696 601 1698
rect 2286 1697 2292 1698
rect 503 1695 504 1696
rect 498 1694 504 1695
rect 2286 1693 2287 1697
rect 2291 1693 2292 1697
rect 2286 1692 2292 1693
rect 2398 1697 2404 1698
rect 2398 1693 2399 1697
rect 2403 1693 2404 1697
rect 2398 1692 2404 1693
rect 2518 1697 2524 1698
rect 2518 1693 2519 1697
rect 2523 1693 2524 1697
rect 2518 1692 2524 1693
rect 2646 1697 2652 1698
rect 2646 1693 2647 1697
rect 2651 1693 2652 1697
rect 2646 1692 2652 1693
rect 2766 1697 2772 1698
rect 2766 1693 2767 1697
rect 2771 1693 2772 1697
rect 2766 1692 2772 1693
rect 2886 1697 2892 1698
rect 2886 1693 2887 1697
rect 2891 1693 2892 1697
rect 2886 1692 2892 1693
rect 3006 1697 3012 1698
rect 3006 1693 3007 1697
rect 3011 1693 3012 1697
rect 3006 1692 3012 1693
rect 3126 1697 3132 1698
rect 3126 1693 3127 1697
rect 3131 1693 3132 1697
rect 3126 1692 3132 1693
rect 3246 1697 3252 1698
rect 3246 1693 3247 1697
rect 3251 1693 3252 1697
rect 3246 1692 3252 1693
rect 3374 1697 3380 1698
rect 3374 1693 3375 1697
rect 3379 1693 3380 1697
rect 3374 1692 3380 1693
rect 3478 1697 3484 1698
rect 3478 1693 3479 1697
rect 3483 1693 3484 1697
rect 3478 1692 3484 1693
rect 3498 1691 3504 1692
rect 110 1687 116 1688
rect 110 1683 111 1687
rect 115 1683 116 1687
rect 110 1682 116 1683
rect 1210 1687 1216 1688
rect 1210 1683 1211 1687
rect 1215 1686 1216 1687
rect 1822 1687 1828 1688
rect 1215 1684 1273 1686
rect 1215 1683 1216 1684
rect 1210 1682 1216 1683
rect 1822 1683 1823 1687
rect 1827 1683 1828 1687
rect 3498 1687 3499 1691
rect 3503 1690 3504 1691
rect 3527 1691 3533 1692
rect 3527 1690 3528 1691
rect 3503 1688 3528 1690
rect 3503 1687 3504 1688
rect 3498 1686 3504 1687
rect 3527 1687 3528 1688
rect 3532 1687 3533 1691
rect 3527 1686 3533 1687
rect 1822 1682 1828 1683
rect 2306 1679 2312 1680
rect 134 1677 140 1678
rect 134 1673 135 1677
rect 139 1673 140 1677
rect 134 1672 140 1673
rect 270 1677 276 1678
rect 270 1673 271 1677
rect 275 1673 276 1677
rect 270 1672 276 1673
rect 422 1677 428 1678
rect 422 1673 423 1677
rect 427 1673 428 1677
rect 422 1672 428 1673
rect 574 1677 580 1678
rect 574 1673 575 1677
rect 579 1673 580 1677
rect 574 1672 580 1673
rect 718 1677 724 1678
rect 718 1673 719 1677
rect 723 1673 724 1677
rect 718 1672 724 1673
rect 854 1677 860 1678
rect 854 1673 855 1677
rect 859 1673 860 1677
rect 854 1672 860 1673
rect 982 1677 988 1678
rect 982 1673 983 1677
rect 987 1673 988 1677
rect 982 1672 988 1673
rect 1118 1677 1124 1678
rect 1118 1673 1119 1677
rect 1123 1673 1124 1677
rect 1118 1672 1124 1673
rect 1254 1677 1260 1678
rect 1254 1673 1255 1677
rect 1259 1673 1260 1677
rect 2306 1675 2307 1679
rect 2311 1678 2312 1679
rect 2311 1676 2574 1678
rect 2311 1675 2312 1676
rect 2306 1674 2312 1675
rect 1254 1672 1260 1673
rect 154 1671 160 1672
rect 154 1667 155 1671
rect 159 1670 160 1671
rect 183 1671 189 1672
rect 183 1670 184 1671
rect 159 1668 184 1670
rect 159 1667 160 1668
rect 154 1666 160 1667
rect 183 1667 184 1668
rect 188 1667 189 1671
rect 183 1666 189 1667
rect 2142 1671 2148 1672
rect 2142 1667 2143 1671
rect 2147 1667 2148 1671
rect 2142 1666 2148 1667
rect 2246 1671 2252 1672
rect 2246 1667 2247 1671
rect 2251 1667 2252 1671
rect 2246 1666 2252 1667
rect 2366 1671 2372 1672
rect 2366 1667 2367 1671
rect 2371 1667 2372 1671
rect 2366 1666 2372 1667
rect 2502 1671 2508 1672
rect 2502 1667 2503 1671
rect 2507 1667 2508 1671
rect 2502 1666 2508 1667
rect 2572 1662 2574 1676
rect 2646 1671 2652 1672
rect 2646 1667 2647 1671
rect 2651 1667 2652 1671
rect 2646 1666 2652 1667
rect 2806 1671 2812 1672
rect 2806 1667 2807 1671
rect 2811 1667 2812 1671
rect 2806 1666 2812 1667
rect 2974 1671 2980 1672
rect 2974 1667 2975 1671
rect 2979 1667 2980 1671
rect 2974 1666 2980 1667
rect 3142 1671 3148 1672
rect 3142 1667 3143 1671
rect 3147 1667 3148 1671
rect 3142 1666 3148 1667
rect 3318 1671 3324 1672
rect 3318 1667 3319 1671
rect 3323 1667 3324 1671
rect 3318 1666 3324 1667
rect 3478 1671 3484 1672
rect 3478 1667 3479 1671
rect 3483 1667 3484 1671
rect 3478 1666 3484 1667
rect 2954 1663 2960 1664
rect 1862 1661 1868 1662
rect 1862 1657 1863 1661
rect 1867 1657 1868 1661
rect 2572 1660 2665 1662
rect 2954 1659 2955 1663
rect 2959 1662 2960 1663
rect 3042 1663 3048 1664
rect 2959 1660 2993 1662
rect 2959 1659 2960 1660
rect 2954 1658 2960 1659
rect 3042 1659 3043 1663
rect 3047 1662 3048 1663
rect 3047 1660 3161 1662
rect 3574 1661 3580 1662
rect 3047 1659 3048 1660
rect 3042 1658 3048 1659
rect 1862 1656 1868 1657
rect 3574 1657 3575 1661
rect 3579 1657 3580 1661
rect 3574 1656 3580 1657
rect 134 1655 140 1656
rect 134 1651 135 1655
rect 139 1651 140 1655
rect 134 1650 140 1651
rect 262 1655 268 1656
rect 262 1651 263 1655
rect 267 1651 268 1655
rect 262 1650 268 1651
rect 422 1655 428 1656
rect 422 1651 423 1655
rect 427 1651 428 1655
rect 422 1650 428 1651
rect 574 1655 580 1656
rect 574 1651 575 1655
rect 579 1651 580 1655
rect 574 1650 580 1651
rect 726 1655 732 1656
rect 726 1651 727 1655
rect 731 1651 732 1655
rect 726 1650 732 1651
rect 870 1655 876 1656
rect 870 1651 871 1655
rect 875 1651 876 1655
rect 870 1650 876 1651
rect 1006 1655 1012 1656
rect 1006 1651 1007 1655
rect 1011 1651 1012 1655
rect 1006 1650 1012 1651
rect 1142 1655 1148 1656
rect 1142 1651 1143 1655
rect 1147 1651 1148 1655
rect 1142 1650 1148 1651
rect 1278 1655 1284 1656
rect 1278 1651 1279 1655
rect 1283 1651 1284 1655
rect 1278 1650 1284 1651
rect 1414 1655 1420 1656
rect 1414 1651 1415 1655
rect 1419 1651 1420 1655
rect 1414 1650 1420 1651
rect 202 1647 208 1648
rect 110 1645 116 1646
rect 110 1641 111 1645
rect 115 1641 116 1645
rect 202 1643 203 1647
rect 207 1646 208 1647
rect 567 1647 573 1648
rect 207 1644 281 1646
rect 207 1643 208 1644
rect 202 1642 208 1643
rect 567 1643 568 1647
rect 572 1646 573 1647
rect 1346 1647 1352 1648
rect 572 1644 593 1646
rect 572 1643 573 1644
rect 567 1642 573 1643
rect 1346 1643 1347 1647
rect 1351 1646 1352 1647
rect 2239 1647 2245 1648
rect 2239 1646 2240 1647
rect 1351 1644 1433 1646
rect 1822 1645 1828 1646
rect 1351 1643 1352 1644
rect 1346 1642 1352 1643
rect 110 1640 116 1641
rect 1822 1641 1823 1645
rect 1827 1641 1828 1645
rect 1822 1640 1828 1641
rect 1862 1644 1868 1645
rect 2205 1644 2240 1646
rect 1862 1640 1863 1644
rect 1867 1640 1868 1644
rect 2239 1643 2240 1644
rect 2244 1643 2245 1647
rect 2359 1647 2365 1648
rect 2359 1646 2360 1647
rect 2309 1644 2360 1646
rect 2239 1642 2245 1643
rect 2359 1643 2360 1644
rect 2364 1643 2365 1647
rect 2495 1647 2501 1648
rect 2495 1646 2496 1647
rect 2429 1644 2496 1646
rect 2359 1642 2365 1643
rect 2495 1643 2496 1644
rect 2500 1643 2501 1647
rect 2639 1647 2645 1648
rect 2639 1646 2640 1647
rect 2565 1644 2640 1646
rect 2495 1642 2501 1643
rect 2639 1643 2640 1644
rect 2644 1643 2645 1647
rect 2966 1647 2972 1648
rect 2966 1646 2967 1647
rect 2869 1644 2967 1646
rect 2639 1642 2645 1643
rect 2966 1643 2967 1644
rect 2971 1643 2972 1647
rect 3446 1647 3452 1648
rect 3446 1646 3447 1647
rect 3381 1644 3447 1646
rect 2966 1642 2972 1643
rect 3446 1643 3447 1644
rect 3451 1643 3452 1647
rect 3446 1642 3452 1643
rect 3471 1647 3477 1648
rect 3471 1643 3472 1647
rect 3476 1646 3477 1647
rect 3476 1644 3505 1646
rect 3574 1644 3580 1645
rect 3476 1643 3477 1644
rect 3471 1642 3477 1643
rect 1862 1639 1868 1640
rect 3574 1640 3575 1644
rect 3579 1640 3580 1644
rect 3574 1639 3580 1640
rect 255 1631 261 1632
rect 255 1630 256 1631
rect 110 1628 116 1629
rect 197 1628 256 1630
rect 110 1624 111 1628
rect 115 1624 116 1628
rect 255 1627 256 1628
rect 260 1627 261 1631
rect 567 1631 573 1632
rect 567 1630 568 1631
rect 485 1628 568 1630
rect 255 1626 261 1627
rect 567 1627 568 1628
rect 572 1627 573 1631
rect 567 1626 573 1627
rect 642 1631 648 1632
rect 642 1627 643 1631
rect 647 1630 648 1631
rect 999 1631 1005 1632
rect 999 1630 1000 1631
rect 647 1628 753 1630
rect 933 1628 1000 1630
rect 647 1627 648 1628
rect 642 1626 648 1627
rect 999 1627 1000 1628
rect 1004 1627 1005 1631
rect 1098 1631 1104 1632
rect 1098 1630 1099 1631
rect 1069 1628 1099 1630
rect 999 1626 1005 1627
rect 1098 1627 1099 1628
rect 1103 1627 1104 1631
rect 1271 1631 1277 1632
rect 1271 1630 1272 1631
rect 1205 1628 1272 1630
rect 1098 1626 1104 1627
rect 1271 1627 1272 1628
rect 1276 1627 1277 1631
rect 1407 1631 1413 1632
rect 1407 1630 1408 1631
rect 1341 1628 1408 1630
rect 1271 1626 1277 1627
rect 1407 1627 1408 1628
rect 1412 1627 1413 1631
rect 2150 1631 2156 1632
rect 1407 1626 1413 1627
rect 1822 1628 1828 1629
rect 110 1623 116 1624
rect 1822 1624 1823 1628
rect 1827 1624 1828 1628
rect 2150 1627 2151 1631
rect 2155 1627 2156 1631
rect 2150 1626 2156 1627
rect 2254 1631 2260 1632
rect 2254 1627 2255 1631
rect 2259 1627 2260 1631
rect 2254 1626 2260 1627
rect 2374 1631 2380 1632
rect 2374 1627 2375 1631
rect 2379 1627 2380 1631
rect 2374 1626 2380 1627
rect 2510 1631 2516 1632
rect 2510 1627 2511 1631
rect 2515 1627 2516 1631
rect 2510 1626 2516 1627
rect 2654 1631 2660 1632
rect 2654 1627 2655 1631
rect 2659 1627 2660 1631
rect 2654 1626 2660 1627
rect 2814 1631 2820 1632
rect 2814 1627 2815 1631
rect 2819 1627 2820 1631
rect 2814 1626 2820 1627
rect 2982 1631 2988 1632
rect 2982 1627 2983 1631
rect 2987 1627 2988 1631
rect 2982 1626 2988 1627
rect 3150 1631 3156 1632
rect 3150 1627 3151 1631
rect 3155 1627 3156 1631
rect 3150 1626 3156 1627
rect 3326 1631 3332 1632
rect 3326 1627 3327 1631
rect 3331 1627 3332 1631
rect 3326 1626 3332 1627
rect 3486 1631 3492 1632
rect 3486 1627 3487 1631
rect 3491 1627 3492 1631
rect 3486 1626 3492 1627
rect 1822 1623 1828 1624
rect 2159 1619 2165 1620
rect 142 1615 148 1616
rect 142 1611 143 1615
rect 147 1611 148 1615
rect 142 1610 148 1611
rect 270 1615 276 1616
rect 270 1611 271 1615
rect 275 1611 276 1615
rect 270 1610 276 1611
rect 430 1615 436 1616
rect 430 1611 431 1615
rect 435 1611 436 1615
rect 430 1610 436 1611
rect 582 1615 588 1616
rect 582 1611 583 1615
rect 587 1611 588 1615
rect 582 1610 588 1611
rect 734 1615 740 1616
rect 734 1611 735 1615
rect 739 1611 740 1615
rect 734 1610 740 1611
rect 878 1615 884 1616
rect 878 1611 879 1615
rect 883 1611 884 1615
rect 878 1610 884 1611
rect 1014 1615 1020 1616
rect 1014 1611 1015 1615
rect 1019 1611 1020 1615
rect 1014 1610 1020 1611
rect 1150 1615 1156 1616
rect 1150 1611 1151 1615
rect 1155 1611 1156 1615
rect 1150 1610 1156 1611
rect 1286 1615 1292 1616
rect 1286 1611 1287 1615
rect 1291 1611 1292 1615
rect 1286 1610 1292 1611
rect 1422 1615 1428 1616
rect 1422 1611 1423 1615
rect 1427 1611 1428 1615
rect 2159 1615 2160 1619
rect 2164 1618 2165 1619
rect 2226 1619 2232 1620
rect 2226 1618 2227 1619
rect 2164 1616 2227 1618
rect 2164 1615 2165 1616
rect 2159 1614 2165 1615
rect 2226 1615 2227 1616
rect 2231 1615 2232 1619
rect 2226 1614 2232 1615
rect 2239 1619 2245 1620
rect 2239 1615 2240 1619
rect 2244 1618 2245 1619
rect 2263 1619 2269 1620
rect 2263 1618 2264 1619
rect 2244 1616 2264 1618
rect 2244 1615 2245 1616
rect 2239 1614 2245 1615
rect 2263 1615 2264 1616
rect 2268 1615 2269 1619
rect 2263 1614 2269 1615
rect 2359 1619 2365 1620
rect 2359 1615 2360 1619
rect 2364 1618 2365 1619
rect 2383 1619 2389 1620
rect 2383 1618 2384 1619
rect 2364 1616 2384 1618
rect 2364 1615 2365 1616
rect 2359 1614 2365 1615
rect 2383 1615 2384 1616
rect 2388 1615 2389 1619
rect 2383 1614 2389 1615
rect 2495 1619 2501 1620
rect 2495 1615 2496 1619
rect 2500 1618 2501 1619
rect 2519 1619 2525 1620
rect 2519 1618 2520 1619
rect 2500 1616 2520 1618
rect 2500 1615 2501 1616
rect 2495 1614 2501 1615
rect 2519 1615 2520 1616
rect 2524 1615 2525 1619
rect 2519 1614 2525 1615
rect 2639 1619 2645 1620
rect 2639 1615 2640 1619
rect 2644 1618 2645 1619
rect 2663 1619 2669 1620
rect 2663 1618 2664 1619
rect 2644 1616 2664 1618
rect 2644 1615 2645 1616
rect 2639 1614 2645 1615
rect 2663 1615 2664 1616
rect 2668 1615 2669 1619
rect 2663 1614 2669 1615
rect 2823 1619 2829 1620
rect 2823 1615 2824 1619
rect 2828 1618 2829 1619
rect 2854 1619 2860 1620
rect 2854 1618 2855 1619
rect 2828 1616 2855 1618
rect 2828 1615 2829 1616
rect 2823 1614 2829 1615
rect 2854 1615 2855 1616
rect 2859 1615 2860 1619
rect 2854 1614 2860 1615
rect 2966 1619 2972 1620
rect 2966 1615 2967 1619
rect 2971 1618 2972 1619
rect 2991 1619 2997 1620
rect 2991 1618 2992 1619
rect 2971 1616 2992 1618
rect 2971 1615 2972 1616
rect 2966 1614 2972 1615
rect 2991 1615 2992 1616
rect 2996 1615 2997 1619
rect 2991 1614 2997 1615
rect 3159 1619 3165 1620
rect 3159 1615 3160 1619
rect 3164 1618 3165 1619
rect 3186 1619 3192 1620
rect 3186 1618 3187 1619
rect 3164 1616 3187 1618
rect 3164 1615 3165 1616
rect 3159 1614 3165 1615
rect 3186 1615 3187 1616
rect 3191 1615 3192 1619
rect 3186 1614 3192 1615
rect 3334 1619 3341 1620
rect 3334 1615 3335 1619
rect 3340 1615 3341 1619
rect 3334 1614 3341 1615
rect 3495 1619 3504 1620
rect 3495 1615 3496 1619
rect 3503 1615 3504 1619
rect 3495 1614 3504 1615
rect 1422 1610 1428 1611
rect 2015 1607 2024 1608
rect 151 1603 160 1604
rect 151 1599 152 1603
rect 159 1599 160 1603
rect 151 1598 160 1599
rect 255 1603 261 1604
rect 255 1599 256 1603
rect 260 1602 261 1603
rect 279 1603 285 1604
rect 279 1602 280 1603
rect 260 1600 280 1602
rect 260 1599 261 1600
rect 255 1598 261 1599
rect 279 1599 280 1600
rect 284 1599 285 1603
rect 279 1598 285 1599
rect 439 1603 448 1604
rect 439 1599 440 1603
rect 447 1599 448 1603
rect 439 1598 448 1599
rect 567 1603 573 1604
rect 567 1599 568 1603
rect 572 1602 573 1603
rect 591 1603 597 1604
rect 591 1602 592 1603
rect 572 1600 592 1602
rect 572 1599 573 1600
rect 567 1598 573 1599
rect 591 1599 592 1600
rect 596 1599 597 1603
rect 591 1598 597 1599
rect 742 1603 749 1604
rect 742 1599 743 1603
rect 748 1599 749 1603
rect 742 1598 749 1599
rect 887 1603 896 1604
rect 887 1599 888 1603
rect 895 1599 896 1603
rect 887 1598 896 1599
rect 999 1603 1005 1604
rect 999 1599 1000 1603
rect 1004 1602 1005 1603
rect 1023 1603 1029 1604
rect 1023 1602 1024 1603
rect 1004 1600 1024 1602
rect 1004 1599 1005 1600
rect 999 1598 1005 1599
rect 1023 1599 1024 1600
rect 1028 1599 1029 1603
rect 1023 1598 1029 1599
rect 1098 1603 1104 1604
rect 1098 1599 1099 1603
rect 1103 1602 1104 1603
rect 1159 1603 1165 1604
rect 1159 1602 1160 1603
rect 1103 1600 1160 1602
rect 1103 1599 1104 1600
rect 1098 1598 1104 1599
rect 1159 1599 1160 1600
rect 1164 1599 1165 1603
rect 1159 1598 1165 1599
rect 1271 1603 1277 1604
rect 1271 1599 1272 1603
rect 1276 1602 1277 1603
rect 1295 1603 1301 1604
rect 1295 1602 1296 1603
rect 1276 1600 1296 1602
rect 1276 1599 1277 1600
rect 1271 1598 1277 1599
rect 1295 1599 1296 1600
rect 1300 1599 1301 1603
rect 1295 1598 1301 1599
rect 1407 1603 1413 1604
rect 1407 1599 1408 1603
rect 1412 1602 1413 1603
rect 1431 1603 1437 1604
rect 1431 1602 1432 1603
rect 1412 1600 1432 1602
rect 1412 1599 1413 1600
rect 1407 1598 1413 1599
rect 1431 1599 1432 1600
rect 1436 1599 1437 1603
rect 2015 1603 2016 1607
rect 2023 1603 2024 1607
rect 2015 1602 2024 1603
rect 2071 1607 2077 1608
rect 2071 1603 2072 1607
rect 2076 1606 2077 1607
rect 2111 1607 2117 1608
rect 2111 1606 2112 1607
rect 2076 1604 2112 1606
rect 2076 1603 2077 1604
rect 2071 1602 2077 1603
rect 2111 1603 2112 1604
rect 2116 1603 2117 1607
rect 2111 1602 2117 1603
rect 2167 1607 2173 1608
rect 2167 1603 2168 1607
rect 2172 1606 2173 1607
rect 2215 1607 2221 1608
rect 2215 1606 2216 1607
rect 2172 1604 2216 1606
rect 2172 1603 2173 1604
rect 2167 1602 2173 1603
rect 2215 1603 2216 1604
rect 2220 1603 2221 1607
rect 2215 1602 2221 1603
rect 2271 1607 2277 1608
rect 2271 1603 2272 1607
rect 2276 1606 2277 1607
rect 2335 1607 2341 1608
rect 2335 1606 2336 1607
rect 2276 1604 2336 1606
rect 2276 1603 2277 1604
rect 2271 1602 2277 1603
rect 2335 1603 2336 1604
rect 2340 1603 2341 1607
rect 2335 1602 2341 1603
rect 2399 1607 2405 1608
rect 2399 1603 2400 1607
rect 2404 1606 2405 1607
rect 2471 1607 2477 1608
rect 2471 1606 2472 1607
rect 2404 1604 2472 1606
rect 2404 1603 2405 1604
rect 2399 1602 2405 1603
rect 2471 1603 2472 1604
rect 2476 1603 2477 1607
rect 2471 1602 2477 1603
rect 2615 1607 2621 1608
rect 2615 1603 2616 1607
rect 2620 1606 2621 1607
rect 2695 1607 2701 1608
rect 2695 1606 2696 1607
rect 2620 1604 2696 1606
rect 2620 1603 2621 1604
rect 2615 1602 2621 1603
rect 2695 1603 2696 1604
rect 2700 1603 2701 1607
rect 2695 1602 2701 1603
rect 2775 1607 2781 1608
rect 2775 1603 2776 1607
rect 2780 1606 2781 1607
rect 2847 1607 2853 1608
rect 2847 1606 2848 1607
rect 2780 1604 2848 1606
rect 2780 1603 2781 1604
rect 2775 1602 2781 1603
rect 2847 1603 2848 1604
rect 2852 1603 2853 1607
rect 2847 1602 2853 1603
rect 2951 1607 2960 1608
rect 2951 1603 2952 1607
rect 2959 1603 2960 1607
rect 2951 1602 2960 1603
rect 3135 1607 3141 1608
rect 3135 1603 3136 1607
rect 3140 1606 3141 1607
rect 3199 1607 3205 1608
rect 3199 1606 3200 1607
rect 3140 1604 3200 1606
rect 3140 1603 3141 1604
rect 3135 1602 3141 1603
rect 3199 1603 3200 1604
rect 3204 1603 3205 1607
rect 3327 1607 3333 1608
rect 3327 1604 3328 1607
rect 3199 1602 3205 1603
rect 3326 1603 3328 1604
rect 3332 1603 3333 1607
rect 1431 1598 1437 1599
rect 3326 1599 3327 1603
rect 3331 1602 3333 1603
rect 3471 1607 3477 1608
rect 3471 1603 3472 1607
rect 3476 1606 3477 1607
rect 3495 1607 3501 1608
rect 3495 1606 3496 1607
rect 3476 1604 3496 1606
rect 3476 1603 3477 1604
rect 3471 1602 3477 1603
rect 3495 1603 3496 1604
rect 3500 1603 3501 1607
rect 3495 1602 3501 1603
rect 3331 1599 3332 1602
rect 3326 1598 3332 1599
rect 2006 1597 2012 1598
rect 750 1595 756 1596
rect 750 1594 751 1595
rect 592 1592 751 1594
rect 175 1587 181 1588
rect 175 1583 176 1587
rect 180 1586 181 1587
rect 202 1587 208 1588
rect 202 1586 203 1587
rect 180 1584 203 1586
rect 180 1583 181 1584
rect 175 1582 181 1583
rect 202 1583 203 1584
rect 207 1583 208 1587
rect 202 1582 208 1583
rect 247 1587 253 1588
rect 247 1583 248 1587
rect 252 1586 253 1587
rect 343 1587 349 1588
rect 343 1586 344 1587
rect 252 1584 344 1586
rect 252 1583 253 1584
rect 247 1582 253 1583
rect 343 1583 344 1584
rect 348 1583 349 1587
rect 343 1582 349 1583
rect 519 1587 525 1588
rect 519 1583 520 1587
rect 524 1586 525 1587
rect 592 1586 594 1592
rect 750 1591 751 1592
rect 755 1591 756 1595
rect 2006 1593 2007 1597
rect 2011 1593 2012 1597
rect 2006 1592 2012 1593
rect 2102 1597 2108 1598
rect 2102 1593 2103 1597
rect 2107 1593 2108 1597
rect 2102 1592 2108 1593
rect 2206 1597 2212 1598
rect 2206 1593 2207 1597
rect 2211 1593 2212 1597
rect 2206 1592 2212 1593
rect 2326 1597 2332 1598
rect 2326 1593 2327 1597
rect 2331 1593 2332 1597
rect 2326 1592 2332 1593
rect 2462 1597 2468 1598
rect 2462 1593 2463 1597
rect 2467 1593 2468 1597
rect 2462 1592 2468 1593
rect 2606 1597 2612 1598
rect 2606 1593 2607 1597
rect 2611 1593 2612 1597
rect 2606 1592 2612 1593
rect 2766 1597 2772 1598
rect 2766 1593 2767 1597
rect 2771 1593 2772 1597
rect 2766 1592 2772 1593
rect 2942 1597 2948 1598
rect 2942 1593 2943 1597
rect 2947 1593 2948 1597
rect 2942 1592 2948 1593
rect 3126 1597 3132 1598
rect 3126 1593 3127 1597
rect 3131 1593 3132 1597
rect 3126 1592 3132 1593
rect 3318 1597 3324 1598
rect 3318 1593 3319 1597
rect 3323 1593 3324 1597
rect 3318 1592 3324 1593
rect 3486 1597 3492 1598
rect 3486 1593 3487 1597
rect 3491 1593 3492 1597
rect 3486 1592 3492 1593
rect 750 1590 756 1591
rect 524 1584 594 1586
rect 599 1587 605 1588
rect 524 1583 525 1584
rect 519 1582 525 1583
rect 599 1583 600 1587
rect 604 1586 605 1587
rect 687 1587 693 1588
rect 687 1586 688 1587
rect 604 1584 688 1586
rect 604 1583 605 1584
rect 599 1582 605 1583
rect 687 1583 688 1584
rect 692 1583 693 1587
rect 687 1582 693 1583
rect 855 1587 864 1588
rect 855 1583 856 1587
rect 863 1583 864 1587
rect 855 1582 864 1583
rect 1007 1587 1013 1588
rect 1007 1583 1008 1587
rect 1012 1586 1013 1587
rect 1022 1587 1028 1588
rect 1022 1586 1023 1587
rect 1012 1584 1023 1586
rect 1012 1583 1013 1584
rect 1007 1582 1013 1583
rect 1022 1583 1023 1584
rect 1027 1583 1028 1587
rect 1022 1582 1028 1583
rect 1079 1587 1085 1588
rect 1079 1583 1080 1587
rect 1084 1586 1085 1587
rect 1159 1587 1165 1588
rect 1159 1586 1160 1587
rect 1084 1584 1160 1586
rect 1084 1583 1085 1584
rect 1079 1582 1085 1583
rect 1159 1583 1160 1584
rect 1164 1583 1165 1587
rect 1159 1582 1165 1583
rect 1231 1587 1237 1588
rect 1231 1583 1232 1587
rect 1236 1586 1237 1587
rect 1303 1587 1309 1588
rect 1303 1586 1304 1587
rect 1236 1584 1304 1586
rect 1236 1583 1237 1584
rect 1231 1582 1237 1583
rect 1303 1583 1304 1584
rect 1308 1583 1309 1587
rect 1303 1582 1309 1583
rect 1375 1587 1381 1588
rect 1375 1583 1376 1587
rect 1380 1586 1381 1587
rect 1447 1587 1453 1588
rect 1447 1586 1448 1587
rect 1380 1584 1448 1586
rect 1380 1583 1381 1584
rect 1375 1582 1381 1583
rect 1447 1583 1448 1584
rect 1452 1583 1453 1587
rect 1447 1582 1453 1583
rect 1519 1587 1525 1588
rect 1519 1583 1520 1587
rect 1524 1586 1525 1587
rect 1591 1587 1597 1588
rect 1591 1586 1592 1587
rect 1524 1584 1592 1586
rect 1524 1583 1525 1584
rect 1519 1582 1525 1583
rect 1591 1583 1592 1584
rect 1596 1583 1597 1587
rect 1591 1582 1597 1583
rect 1862 1584 1868 1585
rect 3574 1584 3580 1585
rect 1862 1580 1863 1584
rect 1867 1580 1868 1584
rect 2071 1583 2077 1584
rect 2071 1582 2072 1583
rect 2061 1580 2072 1582
rect 1862 1579 1868 1580
rect 2071 1579 2072 1580
rect 2076 1579 2077 1583
rect 2167 1583 2173 1584
rect 2167 1582 2168 1583
rect 2157 1580 2168 1582
rect 2071 1578 2077 1579
rect 2167 1579 2168 1580
rect 2172 1579 2173 1583
rect 2271 1583 2277 1584
rect 2271 1582 2272 1583
rect 2261 1580 2272 1582
rect 2167 1578 2173 1579
rect 2271 1579 2272 1580
rect 2276 1579 2277 1583
rect 2399 1583 2405 1584
rect 2399 1582 2400 1583
rect 2381 1580 2400 1582
rect 2271 1578 2277 1579
rect 2399 1579 2400 1580
rect 2404 1579 2405 1583
rect 3186 1583 3192 1584
rect 3186 1582 3187 1583
rect 3181 1580 3187 1582
rect 2399 1578 2405 1579
rect 2695 1579 2701 1580
rect 166 1577 172 1578
rect 166 1573 167 1577
rect 171 1573 172 1577
rect 166 1572 172 1573
rect 334 1577 340 1578
rect 334 1573 335 1577
rect 339 1573 340 1577
rect 334 1572 340 1573
rect 510 1577 516 1578
rect 510 1573 511 1577
rect 515 1573 516 1577
rect 510 1572 516 1573
rect 678 1577 684 1578
rect 678 1573 679 1577
rect 683 1573 684 1577
rect 678 1572 684 1573
rect 846 1577 852 1578
rect 846 1573 847 1577
rect 851 1573 852 1577
rect 846 1572 852 1573
rect 998 1577 1004 1578
rect 998 1573 999 1577
rect 1003 1573 1004 1577
rect 998 1572 1004 1573
rect 1150 1577 1156 1578
rect 1150 1573 1151 1577
rect 1155 1573 1156 1577
rect 1150 1572 1156 1573
rect 1294 1577 1300 1578
rect 1294 1573 1295 1577
rect 1299 1573 1300 1577
rect 1294 1572 1300 1573
rect 1438 1577 1444 1578
rect 1438 1573 1439 1577
rect 1443 1573 1444 1577
rect 1438 1572 1444 1573
rect 1582 1577 1588 1578
rect 1582 1573 1583 1577
rect 1587 1573 1588 1577
rect 2695 1575 2696 1579
rect 2700 1578 2701 1579
rect 2847 1579 2853 1580
rect 2700 1576 2785 1578
rect 2700 1575 2701 1576
rect 2695 1574 2701 1575
rect 2847 1575 2848 1579
rect 2852 1578 2853 1579
rect 3186 1579 3187 1580
rect 3191 1579 3192 1583
rect 3574 1580 3575 1584
rect 3579 1580 3580 1584
rect 3186 1578 3192 1579
rect 3199 1579 3205 1580
rect 2852 1576 2961 1578
rect 2852 1575 2853 1576
rect 2847 1574 2853 1575
rect 3199 1575 3200 1579
rect 3204 1578 3205 1579
rect 3462 1579 3468 1580
rect 3574 1579 3580 1580
rect 3204 1576 3337 1578
rect 3204 1575 3205 1576
rect 3199 1574 3205 1575
rect 3462 1575 3463 1579
rect 3467 1578 3468 1579
rect 3467 1576 3505 1578
rect 3467 1575 3468 1576
rect 3462 1574 3468 1575
rect 1582 1572 1588 1573
rect 1862 1567 1868 1568
rect 110 1564 116 1565
rect 1822 1564 1828 1565
rect 110 1560 111 1564
rect 115 1560 116 1564
rect 247 1563 253 1564
rect 247 1562 248 1563
rect 221 1560 248 1562
rect 110 1559 116 1560
rect 247 1559 248 1560
rect 252 1559 253 1563
rect 599 1563 605 1564
rect 599 1562 600 1563
rect 565 1560 600 1562
rect 247 1558 253 1559
rect 599 1559 600 1560
rect 604 1559 605 1563
rect 742 1563 748 1564
rect 742 1562 743 1563
rect 733 1560 743 1562
rect 599 1558 605 1559
rect 742 1559 743 1560
rect 747 1559 748 1563
rect 1079 1563 1085 1564
rect 1079 1562 1080 1563
rect 1053 1560 1080 1562
rect 742 1558 748 1559
rect 750 1559 756 1560
rect 750 1555 751 1559
rect 755 1558 756 1559
rect 1079 1559 1080 1560
rect 1084 1559 1085 1563
rect 1231 1563 1237 1564
rect 1231 1562 1232 1563
rect 1205 1560 1232 1562
rect 1079 1558 1085 1559
rect 1231 1559 1232 1560
rect 1236 1559 1237 1563
rect 1375 1563 1381 1564
rect 1375 1562 1376 1563
rect 1349 1560 1376 1562
rect 1231 1558 1237 1559
rect 1375 1559 1376 1560
rect 1380 1559 1381 1563
rect 1519 1563 1525 1564
rect 1519 1562 1520 1563
rect 1493 1560 1520 1562
rect 1375 1558 1381 1559
rect 1519 1559 1520 1560
rect 1524 1559 1525 1563
rect 1822 1560 1823 1564
rect 1827 1560 1828 1564
rect 1862 1563 1863 1567
rect 1867 1563 1868 1567
rect 2726 1567 2732 1568
rect 2726 1566 2727 1567
rect 1862 1562 1868 1563
rect 2388 1564 2473 1566
rect 2657 1564 2727 1566
rect 1822 1559 1828 1560
rect 1519 1558 1525 1559
rect 755 1556 865 1558
rect 1998 1557 2004 1558
rect 755 1555 756 1556
rect 750 1554 756 1555
rect 1998 1553 1999 1557
rect 2003 1553 2004 1557
rect 1998 1552 2004 1553
rect 2094 1557 2100 1558
rect 2094 1553 2095 1557
rect 2099 1553 2100 1557
rect 2094 1552 2100 1553
rect 2198 1557 2204 1558
rect 2198 1553 2199 1557
rect 2203 1553 2204 1557
rect 2198 1552 2204 1553
rect 2318 1557 2324 1558
rect 2318 1553 2319 1557
rect 2323 1553 2324 1557
rect 2318 1552 2324 1553
rect 2226 1551 2232 1552
rect 110 1547 116 1548
rect 110 1543 111 1547
rect 115 1543 116 1547
rect 406 1547 412 1548
rect 406 1546 407 1547
rect 385 1544 407 1546
rect 110 1542 116 1543
rect 406 1543 407 1544
rect 411 1543 412 1547
rect 406 1542 412 1543
rect 1518 1547 1524 1548
rect 1518 1543 1519 1547
rect 1523 1546 1524 1547
rect 1822 1547 1828 1548
rect 1523 1544 1593 1546
rect 1523 1543 1524 1544
rect 1518 1542 1524 1543
rect 1822 1543 1823 1547
rect 1827 1543 1828 1547
rect 2226 1547 2227 1551
rect 2231 1550 2232 1551
rect 2388 1550 2390 1564
rect 2726 1563 2727 1564
rect 2731 1563 2732 1567
rect 2726 1562 2732 1563
rect 3574 1567 3580 1568
rect 3574 1563 3575 1567
rect 3579 1563 3580 1567
rect 3574 1562 3580 1563
rect 2454 1557 2460 1558
rect 2454 1553 2455 1557
rect 2459 1553 2460 1557
rect 2454 1552 2460 1553
rect 2598 1557 2604 1558
rect 2598 1553 2599 1557
rect 2603 1553 2604 1557
rect 2598 1552 2604 1553
rect 2758 1557 2764 1558
rect 2758 1553 2759 1557
rect 2763 1553 2764 1557
rect 2758 1552 2764 1553
rect 2934 1557 2940 1558
rect 2934 1553 2935 1557
rect 2939 1553 2940 1557
rect 2934 1552 2940 1553
rect 3118 1557 3124 1558
rect 3118 1553 3119 1557
rect 3123 1553 3124 1557
rect 3118 1552 3124 1553
rect 3310 1557 3316 1558
rect 3310 1553 3311 1557
rect 3315 1553 3316 1557
rect 3310 1552 3316 1553
rect 3478 1557 3484 1558
rect 3478 1553 3479 1557
rect 3483 1553 3484 1557
rect 3478 1552 3484 1553
rect 2231 1548 2390 1550
rect 2231 1547 2232 1548
rect 2226 1546 2232 1547
rect 1822 1542 1828 1543
rect 158 1537 164 1538
rect 158 1533 159 1537
rect 163 1533 164 1537
rect 158 1532 164 1533
rect 326 1537 332 1538
rect 326 1533 327 1537
rect 331 1533 332 1537
rect 326 1532 332 1533
rect 502 1537 508 1538
rect 502 1533 503 1537
rect 507 1533 508 1537
rect 502 1532 508 1533
rect 670 1537 676 1538
rect 670 1533 671 1537
rect 675 1533 676 1537
rect 670 1532 676 1533
rect 838 1537 844 1538
rect 838 1533 839 1537
rect 843 1533 844 1537
rect 838 1532 844 1533
rect 990 1537 996 1538
rect 990 1533 991 1537
rect 995 1533 996 1537
rect 990 1532 996 1533
rect 1142 1537 1148 1538
rect 1142 1533 1143 1537
rect 1147 1533 1148 1537
rect 1142 1532 1148 1533
rect 1286 1537 1292 1538
rect 1286 1533 1287 1537
rect 1291 1533 1292 1537
rect 1286 1532 1292 1533
rect 1430 1537 1436 1538
rect 1430 1533 1431 1537
rect 1435 1533 1436 1537
rect 1430 1532 1436 1533
rect 1574 1537 1580 1538
rect 1574 1533 1575 1537
rect 1579 1533 1580 1537
rect 1574 1532 1580 1533
rect 1886 1527 1892 1528
rect 1886 1523 1887 1527
rect 1891 1523 1892 1527
rect 1886 1522 1892 1523
rect 1974 1527 1980 1528
rect 1974 1523 1975 1527
rect 1979 1523 1980 1527
rect 1974 1522 1980 1523
rect 2102 1527 2108 1528
rect 2102 1523 2103 1527
rect 2107 1523 2108 1527
rect 2102 1522 2108 1523
rect 2238 1527 2244 1528
rect 2238 1523 2239 1527
rect 2243 1523 2244 1527
rect 2238 1522 2244 1523
rect 2382 1527 2388 1528
rect 2382 1523 2383 1527
rect 2387 1523 2388 1527
rect 2382 1522 2388 1523
rect 2542 1527 2548 1528
rect 2542 1523 2543 1527
rect 2547 1523 2548 1527
rect 2542 1522 2548 1523
rect 2710 1527 2716 1528
rect 2710 1523 2711 1527
rect 2715 1523 2716 1527
rect 2710 1522 2716 1523
rect 2878 1527 2884 1528
rect 2878 1523 2879 1527
rect 2883 1523 2884 1527
rect 2878 1522 2884 1523
rect 3054 1527 3060 1528
rect 3054 1523 3055 1527
rect 3059 1523 3060 1527
rect 3054 1522 3060 1523
rect 3238 1527 3244 1528
rect 3238 1523 3239 1527
rect 3243 1523 3244 1527
rect 3238 1522 3244 1523
rect 3430 1527 3436 1528
rect 3430 1523 3431 1527
rect 3435 1523 3436 1527
rect 3430 1522 3436 1523
rect 2306 1519 2312 1520
rect 1862 1517 1868 1518
rect 1862 1513 1863 1517
rect 1867 1513 1868 1517
rect 2306 1515 2307 1519
rect 2311 1518 2312 1519
rect 3326 1519 3332 1520
rect 3326 1518 3327 1519
rect 2311 1516 2401 1518
rect 3297 1516 3327 1518
rect 2311 1515 2312 1516
rect 2306 1514 2312 1515
rect 3326 1515 3327 1516
rect 3331 1515 3332 1519
rect 3326 1514 3332 1515
rect 3574 1517 3580 1518
rect 1862 1512 1868 1513
rect 3574 1513 3575 1517
rect 3579 1513 3580 1517
rect 3574 1512 3580 1513
rect 214 1511 220 1512
rect 214 1507 215 1511
rect 219 1507 220 1511
rect 214 1506 220 1507
rect 390 1511 396 1512
rect 390 1507 391 1511
rect 395 1507 396 1511
rect 390 1506 396 1507
rect 574 1511 580 1512
rect 574 1507 575 1511
rect 579 1507 580 1511
rect 574 1506 580 1507
rect 758 1511 764 1512
rect 758 1507 759 1511
rect 763 1507 764 1511
rect 758 1506 764 1507
rect 934 1511 940 1512
rect 934 1507 935 1511
rect 939 1507 940 1511
rect 934 1506 940 1507
rect 1094 1511 1100 1512
rect 1094 1507 1095 1511
rect 1099 1507 1100 1511
rect 1094 1506 1100 1507
rect 1254 1511 1260 1512
rect 1254 1507 1255 1511
rect 1259 1507 1260 1511
rect 1254 1506 1260 1507
rect 1406 1511 1412 1512
rect 1406 1507 1407 1511
rect 1411 1507 1412 1511
rect 1406 1506 1412 1507
rect 1558 1511 1564 1512
rect 1558 1507 1559 1511
rect 1563 1507 1564 1511
rect 1558 1506 1564 1507
rect 1710 1511 1716 1512
rect 1710 1507 1711 1511
rect 1715 1507 1716 1511
rect 1710 1506 1716 1507
rect 858 1503 864 1504
rect 110 1501 116 1502
rect 110 1497 111 1501
rect 115 1497 116 1501
rect 858 1499 859 1503
rect 863 1502 864 1503
rect 1626 1503 1632 1504
rect 863 1500 953 1502
rect 863 1499 864 1500
rect 858 1498 864 1499
rect 1626 1499 1627 1503
rect 1631 1502 1632 1503
rect 1967 1503 1973 1504
rect 1967 1502 1968 1503
rect 1631 1500 1729 1502
rect 1822 1501 1828 1502
rect 1631 1499 1632 1500
rect 1626 1498 1632 1499
rect 110 1496 116 1497
rect 1822 1497 1823 1501
rect 1827 1497 1828 1501
rect 1822 1496 1828 1497
rect 1862 1500 1868 1501
rect 1949 1500 1968 1502
rect 1862 1496 1863 1500
rect 1867 1496 1868 1500
rect 1967 1499 1968 1500
rect 1972 1499 1973 1503
rect 2042 1503 2048 1504
rect 2042 1502 2043 1503
rect 2037 1500 2043 1502
rect 1967 1498 1973 1499
rect 2042 1499 2043 1500
rect 2047 1499 2048 1503
rect 2231 1503 2237 1504
rect 2231 1502 2232 1503
rect 2165 1500 2232 1502
rect 2042 1498 2048 1499
rect 2231 1499 2232 1500
rect 2236 1499 2237 1503
rect 2375 1503 2381 1504
rect 2375 1502 2376 1503
rect 2301 1500 2376 1502
rect 2231 1498 2237 1499
rect 2375 1499 2376 1500
rect 2380 1499 2381 1503
rect 2375 1498 2381 1499
rect 2479 1503 2485 1504
rect 2479 1499 2480 1503
rect 2484 1502 2485 1503
rect 2610 1503 2616 1504
rect 2484 1500 2569 1502
rect 2484 1499 2485 1500
rect 2479 1498 2485 1499
rect 2610 1499 2611 1503
rect 2615 1502 2616 1503
rect 3047 1503 3053 1504
rect 3047 1502 3048 1503
rect 2615 1500 2737 1502
rect 2941 1500 3048 1502
rect 2615 1499 2616 1500
rect 2610 1498 2616 1499
rect 3047 1499 3048 1500
rect 3052 1499 3053 1503
rect 3122 1503 3128 1504
rect 3122 1502 3123 1503
rect 3117 1500 3123 1502
rect 3047 1498 3053 1499
rect 3122 1499 3123 1500
rect 3127 1499 3128 1503
rect 3498 1503 3504 1504
rect 3498 1502 3499 1503
rect 3493 1500 3499 1502
rect 3122 1498 3128 1499
rect 3498 1499 3499 1500
rect 3503 1499 3504 1503
rect 3498 1498 3504 1499
rect 3574 1500 3580 1501
rect 1862 1495 1868 1496
rect 3574 1496 3575 1500
rect 3579 1496 3580 1500
rect 3574 1495 3580 1496
rect 282 1487 288 1488
rect 282 1486 283 1487
rect 110 1484 116 1485
rect 277 1484 283 1486
rect 110 1480 111 1484
rect 115 1480 116 1484
rect 282 1483 283 1484
rect 287 1483 288 1487
rect 282 1482 288 1483
rect 290 1487 296 1488
rect 290 1483 291 1487
rect 295 1486 296 1487
rect 751 1487 757 1488
rect 751 1486 752 1487
rect 295 1484 417 1486
rect 637 1484 752 1486
rect 295 1483 296 1484
rect 290 1482 296 1483
rect 751 1483 752 1484
rect 756 1483 757 1487
rect 927 1487 933 1488
rect 927 1486 928 1487
rect 821 1484 928 1486
rect 751 1482 757 1483
rect 927 1483 928 1484
rect 932 1483 933 1487
rect 1247 1487 1253 1488
rect 1247 1486 1248 1487
rect 1157 1484 1248 1486
rect 927 1482 933 1483
rect 1247 1483 1248 1484
rect 1252 1483 1253 1487
rect 1399 1487 1405 1488
rect 1399 1486 1400 1487
rect 1317 1484 1400 1486
rect 1247 1482 1253 1483
rect 1399 1483 1400 1484
rect 1404 1483 1405 1487
rect 1551 1487 1557 1488
rect 1551 1486 1552 1487
rect 1469 1484 1552 1486
rect 1399 1482 1405 1483
rect 1551 1483 1552 1484
rect 1556 1483 1557 1487
rect 1703 1487 1709 1488
rect 1703 1486 1704 1487
rect 1621 1484 1704 1486
rect 1551 1482 1557 1483
rect 1703 1483 1704 1484
rect 1708 1483 1709 1487
rect 1894 1487 1900 1488
rect 1703 1482 1709 1483
rect 1822 1484 1828 1485
rect 110 1479 116 1480
rect 1822 1480 1823 1484
rect 1827 1480 1828 1484
rect 1894 1483 1895 1487
rect 1899 1483 1900 1487
rect 1894 1482 1900 1483
rect 1982 1487 1988 1488
rect 1982 1483 1983 1487
rect 1987 1483 1988 1487
rect 1982 1482 1988 1483
rect 2110 1487 2116 1488
rect 2110 1483 2111 1487
rect 2115 1483 2116 1487
rect 2110 1482 2116 1483
rect 2246 1487 2252 1488
rect 2246 1483 2247 1487
rect 2251 1483 2252 1487
rect 2246 1482 2252 1483
rect 2390 1487 2396 1488
rect 2390 1483 2391 1487
rect 2395 1483 2396 1487
rect 2390 1482 2396 1483
rect 2550 1487 2556 1488
rect 2550 1483 2551 1487
rect 2555 1483 2556 1487
rect 2550 1482 2556 1483
rect 2718 1487 2724 1488
rect 2718 1483 2719 1487
rect 2723 1483 2724 1487
rect 2718 1482 2724 1483
rect 2886 1487 2892 1488
rect 2886 1483 2887 1487
rect 2891 1483 2892 1487
rect 2886 1482 2892 1483
rect 3062 1487 3068 1488
rect 3062 1483 3063 1487
rect 3067 1483 3068 1487
rect 3062 1482 3068 1483
rect 3246 1487 3252 1488
rect 3246 1483 3247 1487
rect 3251 1483 3252 1487
rect 3246 1482 3252 1483
rect 3438 1487 3444 1488
rect 3438 1483 3439 1487
rect 3443 1483 3444 1487
rect 3438 1482 3444 1483
rect 1822 1479 1828 1480
rect 1903 1475 1909 1476
rect 222 1471 228 1472
rect 222 1467 223 1471
rect 227 1467 228 1471
rect 222 1466 228 1467
rect 398 1471 404 1472
rect 398 1467 399 1471
rect 403 1467 404 1471
rect 398 1466 404 1467
rect 582 1471 588 1472
rect 582 1467 583 1471
rect 587 1467 588 1471
rect 582 1466 588 1467
rect 766 1471 772 1472
rect 766 1467 767 1471
rect 771 1467 772 1471
rect 766 1466 772 1467
rect 942 1471 948 1472
rect 942 1467 943 1471
rect 947 1467 948 1471
rect 942 1466 948 1467
rect 1102 1471 1108 1472
rect 1102 1467 1103 1471
rect 1107 1467 1108 1471
rect 1102 1466 1108 1467
rect 1262 1471 1268 1472
rect 1262 1467 1263 1471
rect 1267 1467 1268 1471
rect 1262 1466 1268 1467
rect 1414 1471 1420 1472
rect 1414 1467 1415 1471
rect 1419 1467 1420 1471
rect 1414 1466 1420 1467
rect 1566 1471 1572 1472
rect 1566 1467 1567 1471
rect 1571 1467 1572 1471
rect 1566 1466 1572 1467
rect 1718 1471 1724 1472
rect 1718 1467 1719 1471
rect 1723 1467 1724 1471
rect 1903 1471 1904 1475
rect 1908 1474 1909 1475
rect 1950 1475 1956 1476
rect 1950 1474 1951 1475
rect 1908 1472 1951 1474
rect 1908 1471 1909 1472
rect 1903 1470 1909 1471
rect 1950 1471 1951 1472
rect 1955 1471 1956 1475
rect 1950 1470 1956 1471
rect 1967 1475 1973 1476
rect 1967 1471 1968 1475
rect 1972 1474 1973 1475
rect 1991 1475 1997 1476
rect 1991 1474 1992 1475
rect 1972 1472 1992 1474
rect 1972 1471 1973 1472
rect 1967 1470 1973 1471
rect 1991 1471 1992 1472
rect 1996 1471 1997 1475
rect 1991 1470 1997 1471
rect 2042 1475 2048 1476
rect 2042 1471 2043 1475
rect 2047 1474 2048 1475
rect 2119 1475 2125 1476
rect 2119 1474 2120 1475
rect 2047 1472 2120 1474
rect 2047 1471 2048 1472
rect 2042 1470 2048 1471
rect 2119 1471 2120 1472
rect 2124 1471 2125 1475
rect 2119 1470 2125 1471
rect 2231 1475 2237 1476
rect 2231 1471 2232 1475
rect 2236 1474 2237 1475
rect 2255 1475 2261 1476
rect 2255 1474 2256 1475
rect 2236 1472 2256 1474
rect 2236 1471 2237 1472
rect 2231 1470 2237 1471
rect 2255 1471 2256 1472
rect 2260 1471 2261 1475
rect 2255 1470 2261 1471
rect 2375 1475 2381 1476
rect 2375 1471 2376 1475
rect 2380 1474 2381 1475
rect 2399 1475 2405 1476
rect 2399 1474 2400 1475
rect 2380 1472 2400 1474
rect 2380 1471 2381 1472
rect 2375 1470 2381 1471
rect 2399 1471 2400 1472
rect 2404 1471 2405 1475
rect 2399 1470 2405 1471
rect 2559 1475 2565 1476
rect 2559 1471 2560 1475
rect 2564 1474 2565 1475
rect 2610 1475 2616 1476
rect 2610 1474 2611 1475
rect 2564 1472 2611 1474
rect 2564 1471 2565 1472
rect 2559 1470 2565 1471
rect 2610 1471 2611 1472
rect 2615 1471 2616 1475
rect 2610 1470 2616 1471
rect 2726 1475 2733 1476
rect 2726 1471 2727 1475
rect 2732 1471 2733 1475
rect 2726 1470 2733 1471
rect 2826 1475 2832 1476
rect 2826 1471 2827 1475
rect 2831 1474 2832 1475
rect 2895 1475 2901 1476
rect 2895 1474 2896 1475
rect 2831 1472 2896 1474
rect 2831 1471 2832 1472
rect 2826 1470 2832 1471
rect 2895 1471 2896 1472
rect 2900 1471 2901 1475
rect 2895 1470 2901 1471
rect 3047 1475 3053 1476
rect 3047 1471 3048 1475
rect 3052 1474 3053 1475
rect 3071 1475 3077 1476
rect 3071 1474 3072 1475
rect 3052 1472 3072 1474
rect 3052 1471 3053 1472
rect 3047 1470 3053 1471
rect 3071 1471 3072 1472
rect 3076 1471 3077 1475
rect 3071 1470 3077 1471
rect 3255 1475 3261 1476
rect 3255 1471 3256 1475
rect 3260 1474 3261 1475
rect 3263 1475 3269 1476
rect 3263 1474 3264 1475
rect 3260 1472 3264 1474
rect 3260 1471 3261 1472
rect 3255 1470 3261 1471
rect 3263 1471 3264 1472
rect 3268 1471 3269 1475
rect 3263 1470 3269 1471
rect 3446 1475 3453 1476
rect 3446 1471 3447 1475
rect 3452 1471 3453 1475
rect 3446 1470 3453 1471
rect 1718 1466 1724 1467
rect 3207 1467 3213 1468
rect 3207 1466 3208 1467
rect 3104 1464 3208 1466
rect 231 1459 237 1460
rect 231 1455 232 1459
rect 236 1458 237 1459
rect 290 1459 296 1460
rect 290 1458 291 1459
rect 236 1456 291 1458
rect 236 1455 237 1456
rect 231 1454 237 1455
rect 290 1455 291 1456
rect 295 1455 296 1459
rect 290 1454 296 1455
rect 406 1459 413 1460
rect 406 1455 407 1459
rect 412 1455 413 1459
rect 406 1454 413 1455
rect 591 1459 597 1460
rect 591 1455 592 1459
rect 596 1458 597 1459
rect 738 1459 744 1460
rect 738 1458 739 1459
rect 596 1456 739 1458
rect 596 1455 597 1456
rect 591 1454 597 1455
rect 738 1455 739 1456
rect 743 1455 744 1459
rect 738 1454 744 1455
rect 751 1459 757 1460
rect 751 1455 752 1459
rect 756 1458 757 1459
rect 775 1459 781 1460
rect 775 1458 776 1459
rect 756 1456 776 1458
rect 756 1455 757 1456
rect 751 1454 757 1455
rect 775 1455 776 1456
rect 780 1455 781 1459
rect 775 1454 781 1455
rect 927 1459 933 1460
rect 927 1455 928 1459
rect 932 1458 933 1459
rect 951 1459 957 1460
rect 951 1458 952 1459
rect 932 1456 952 1458
rect 932 1455 933 1456
rect 927 1454 933 1455
rect 951 1455 952 1456
rect 956 1455 957 1459
rect 951 1454 957 1455
rect 1111 1459 1120 1460
rect 1111 1455 1112 1459
rect 1119 1455 1120 1459
rect 1111 1454 1120 1455
rect 1247 1459 1253 1460
rect 1247 1455 1248 1459
rect 1252 1458 1253 1459
rect 1271 1459 1277 1460
rect 1271 1458 1272 1459
rect 1252 1456 1272 1458
rect 1252 1455 1253 1456
rect 1247 1454 1253 1455
rect 1271 1455 1272 1456
rect 1276 1455 1277 1459
rect 1271 1454 1277 1455
rect 1399 1459 1405 1460
rect 1399 1455 1400 1459
rect 1404 1458 1405 1459
rect 1423 1459 1429 1460
rect 1423 1458 1424 1459
rect 1404 1456 1424 1458
rect 1404 1455 1405 1456
rect 1399 1454 1405 1455
rect 1423 1455 1424 1456
rect 1428 1455 1429 1459
rect 1423 1454 1429 1455
rect 1551 1459 1557 1460
rect 1551 1455 1552 1459
rect 1556 1458 1557 1459
rect 1575 1459 1581 1460
rect 1575 1458 1576 1459
rect 1556 1456 1576 1458
rect 1556 1455 1557 1456
rect 1551 1454 1557 1455
rect 1575 1455 1576 1456
rect 1580 1455 1581 1459
rect 1575 1454 1581 1455
rect 1703 1459 1709 1460
rect 1703 1455 1704 1459
rect 1708 1458 1709 1459
rect 1727 1459 1733 1460
rect 1727 1458 1728 1459
rect 1708 1456 1728 1458
rect 1708 1455 1709 1456
rect 1703 1454 1709 1455
rect 1727 1455 1728 1456
rect 1732 1455 1733 1459
rect 1727 1454 1733 1455
rect 1807 1459 1813 1460
rect 1807 1455 1808 1459
rect 1812 1458 1813 1459
rect 1903 1459 1909 1460
rect 1903 1458 1904 1459
rect 1812 1456 1904 1458
rect 1812 1455 1813 1456
rect 1807 1454 1813 1455
rect 1903 1455 1904 1456
rect 1908 1455 1909 1459
rect 1903 1454 1909 1455
rect 1959 1459 1965 1460
rect 1959 1455 1960 1459
rect 1964 1458 1965 1459
rect 2031 1459 2037 1460
rect 2031 1458 2032 1459
rect 1964 1456 2032 1458
rect 1964 1455 1965 1456
rect 1959 1454 1965 1455
rect 2031 1455 2032 1456
rect 2036 1455 2037 1459
rect 2031 1454 2037 1455
rect 2103 1459 2109 1460
rect 2103 1455 2104 1459
rect 2108 1458 2109 1459
rect 2183 1459 2189 1460
rect 2183 1458 2184 1459
rect 2108 1456 2184 1458
rect 2108 1455 2109 1456
rect 2103 1454 2109 1455
rect 2183 1455 2184 1456
rect 2188 1455 2189 1459
rect 2183 1454 2189 1455
rect 2234 1459 2240 1460
rect 2234 1455 2235 1459
rect 2239 1458 2240 1459
rect 2327 1459 2333 1460
rect 2327 1458 2328 1459
rect 2239 1456 2328 1458
rect 2239 1455 2240 1456
rect 2234 1454 2240 1455
rect 2327 1455 2328 1456
rect 2332 1455 2333 1459
rect 2327 1454 2333 1455
rect 2471 1459 2477 1460
rect 2471 1455 2472 1459
rect 2476 1458 2477 1459
rect 2479 1459 2485 1460
rect 2479 1458 2480 1459
rect 2476 1456 2480 1458
rect 2476 1455 2477 1456
rect 2471 1454 2477 1455
rect 2479 1455 2480 1456
rect 2484 1455 2485 1459
rect 2479 1454 2485 1455
rect 2518 1459 2524 1460
rect 2518 1455 2519 1459
rect 2523 1458 2524 1459
rect 2623 1459 2629 1460
rect 2623 1458 2624 1459
rect 2523 1456 2624 1458
rect 2523 1455 2524 1456
rect 2518 1454 2524 1455
rect 2623 1455 2624 1456
rect 2628 1455 2629 1459
rect 2623 1454 2629 1455
rect 2695 1459 2701 1460
rect 2695 1455 2696 1459
rect 2700 1458 2701 1459
rect 2775 1459 2781 1460
rect 2775 1458 2776 1459
rect 2700 1456 2776 1458
rect 2700 1455 2701 1456
rect 2695 1454 2701 1455
rect 2775 1455 2776 1456
rect 2780 1455 2781 1459
rect 2775 1454 2781 1455
rect 2943 1459 2949 1460
rect 2943 1455 2944 1459
rect 2948 1458 2949 1459
rect 3104 1458 3106 1464
rect 3207 1463 3208 1464
rect 3212 1463 3213 1467
rect 3207 1462 3213 1463
rect 2948 1456 3106 1458
rect 3111 1459 3117 1460
rect 2948 1455 2949 1456
rect 2943 1454 2949 1455
rect 3111 1455 3112 1459
rect 3116 1458 3117 1459
rect 3122 1459 3128 1460
rect 3122 1458 3123 1459
rect 3116 1456 3123 1458
rect 3116 1455 3117 1456
rect 3111 1454 3117 1455
rect 3122 1455 3123 1456
rect 3127 1455 3128 1459
rect 3122 1454 3128 1455
rect 3199 1459 3205 1460
rect 3199 1455 3200 1459
rect 3204 1458 3205 1459
rect 3287 1459 3293 1460
rect 3287 1458 3288 1459
rect 3204 1456 3288 1458
rect 3204 1455 3205 1456
rect 3199 1454 3205 1455
rect 3287 1455 3288 1456
rect 3292 1455 3293 1459
rect 3287 1454 3293 1455
rect 3471 1459 3477 1460
rect 3471 1455 3472 1459
rect 3476 1458 3477 1459
rect 3498 1459 3504 1460
rect 3498 1458 3499 1459
rect 3476 1456 3499 1458
rect 3476 1455 3477 1456
rect 3471 1454 3477 1455
rect 3498 1455 3499 1456
rect 3503 1455 3504 1459
rect 3498 1454 3504 1455
rect 1626 1451 1632 1452
rect 1626 1450 1627 1451
rect 1369 1448 1627 1450
rect 263 1443 269 1444
rect 263 1439 264 1443
rect 268 1442 269 1443
rect 282 1443 288 1444
rect 282 1442 283 1443
rect 268 1440 283 1442
rect 268 1439 269 1440
rect 263 1438 269 1439
rect 282 1439 283 1440
rect 287 1439 288 1443
rect 282 1438 288 1439
rect 330 1443 336 1444
rect 330 1439 331 1443
rect 335 1442 336 1443
rect 391 1443 397 1444
rect 391 1442 392 1443
rect 335 1440 392 1442
rect 335 1439 336 1440
rect 330 1438 336 1439
rect 391 1439 392 1440
rect 396 1439 397 1443
rect 391 1438 397 1439
rect 455 1443 461 1444
rect 455 1439 456 1443
rect 460 1442 461 1443
rect 527 1443 533 1444
rect 527 1442 528 1443
rect 460 1440 528 1442
rect 460 1439 461 1440
rect 455 1438 461 1439
rect 527 1439 528 1440
rect 532 1439 533 1443
rect 527 1438 533 1439
rect 679 1443 685 1444
rect 679 1439 680 1443
rect 684 1442 685 1443
rect 690 1443 696 1444
rect 690 1442 691 1443
rect 684 1440 691 1442
rect 684 1439 685 1440
rect 679 1438 685 1439
rect 690 1439 691 1440
rect 695 1439 696 1443
rect 690 1438 696 1439
rect 759 1443 765 1444
rect 759 1439 760 1443
rect 764 1442 765 1443
rect 839 1443 845 1444
rect 839 1442 840 1443
rect 764 1440 840 1442
rect 764 1439 765 1440
rect 759 1438 765 1439
rect 839 1439 840 1440
rect 844 1439 845 1443
rect 839 1438 845 1439
rect 999 1443 1005 1444
rect 999 1439 1000 1443
rect 1004 1442 1005 1443
rect 1079 1443 1085 1444
rect 1079 1442 1080 1443
rect 1004 1440 1080 1442
rect 1004 1439 1005 1440
rect 999 1438 1005 1439
rect 1079 1439 1080 1440
rect 1084 1439 1085 1443
rect 1079 1438 1085 1439
rect 1151 1443 1157 1444
rect 1151 1439 1152 1443
rect 1156 1442 1157 1443
rect 1202 1443 1208 1444
rect 1202 1442 1203 1443
rect 1156 1440 1203 1442
rect 1156 1439 1157 1440
rect 1151 1438 1157 1439
rect 1202 1439 1203 1440
rect 1207 1439 1208 1443
rect 1202 1438 1208 1439
rect 1303 1443 1309 1444
rect 1303 1439 1304 1443
rect 1308 1442 1309 1443
rect 1369 1442 1371 1448
rect 1626 1447 1627 1448
rect 1631 1447 1632 1451
rect 1626 1446 1632 1447
rect 1894 1449 1900 1450
rect 1894 1445 1895 1449
rect 1899 1445 1900 1449
rect 1894 1444 1900 1445
rect 2022 1449 2028 1450
rect 2022 1445 2023 1449
rect 2027 1445 2028 1449
rect 2022 1444 2028 1445
rect 2174 1449 2180 1450
rect 2174 1445 2175 1449
rect 2179 1445 2180 1449
rect 2174 1444 2180 1445
rect 2318 1449 2324 1450
rect 2318 1445 2319 1449
rect 2323 1445 2324 1449
rect 2318 1444 2324 1445
rect 2462 1449 2468 1450
rect 2462 1445 2463 1449
rect 2467 1445 2468 1449
rect 2462 1444 2468 1445
rect 2614 1449 2620 1450
rect 2614 1445 2615 1449
rect 2619 1445 2620 1449
rect 2614 1444 2620 1445
rect 2766 1449 2772 1450
rect 2766 1445 2767 1449
rect 2771 1445 2772 1449
rect 2766 1444 2772 1445
rect 2934 1449 2940 1450
rect 2934 1445 2935 1449
rect 2939 1445 2940 1449
rect 2934 1444 2940 1445
rect 3102 1449 3108 1450
rect 3102 1445 3103 1449
rect 3107 1445 3108 1449
rect 3102 1444 3108 1445
rect 3278 1449 3284 1450
rect 3278 1445 3279 1449
rect 3283 1445 3284 1449
rect 3278 1444 3284 1445
rect 3462 1449 3468 1450
rect 3462 1445 3463 1449
rect 3467 1445 3468 1449
rect 3462 1444 3468 1445
rect 1308 1440 1371 1442
rect 1375 1443 1381 1444
rect 1308 1439 1309 1440
rect 1303 1438 1309 1439
rect 1375 1439 1376 1443
rect 1380 1442 1381 1443
rect 1455 1443 1461 1444
rect 1455 1442 1456 1443
rect 1380 1440 1456 1442
rect 1380 1439 1381 1440
rect 1375 1438 1381 1439
rect 1455 1439 1456 1440
rect 1460 1439 1461 1443
rect 1455 1438 1461 1439
rect 1527 1443 1533 1444
rect 1527 1439 1528 1443
rect 1532 1442 1533 1443
rect 1607 1443 1613 1444
rect 1607 1442 1608 1443
rect 1532 1440 1608 1442
rect 1532 1439 1533 1440
rect 1527 1438 1533 1439
rect 1607 1439 1608 1440
rect 1612 1439 1613 1443
rect 1607 1438 1613 1439
rect 1678 1443 1684 1444
rect 1678 1439 1679 1443
rect 1683 1442 1684 1443
rect 1743 1443 1749 1444
rect 1743 1442 1744 1443
rect 1683 1440 1744 1442
rect 1683 1439 1684 1440
rect 1678 1438 1684 1439
rect 1743 1439 1744 1440
rect 1748 1439 1749 1443
rect 1743 1438 1749 1439
rect 1862 1436 1868 1437
rect 3574 1436 3580 1437
rect 254 1433 260 1434
rect 254 1429 255 1433
rect 259 1429 260 1433
rect 254 1428 260 1429
rect 382 1433 388 1434
rect 382 1429 383 1433
rect 387 1429 388 1433
rect 382 1428 388 1429
rect 518 1433 524 1434
rect 518 1429 519 1433
rect 523 1429 524 1433
rect 518 1428 524 1429
rect 670 1433 676 1434
rect 670 1429 671 1433
rect 675 1429 676 1433
rect 670 1428 676 1429
rect 830 1433 836 1434
rect 830 1429 831 1433
rect 835 1429 836 1433
rect 830 1428 836 1429
rect 990 1433 996 1434
rect 990 1429 991 1433
rect 995 1429 996 1433
rect 990 1428 996 1429
rect 1142 1433 1148 1434
rect 1142 1429 1143 1433
rect 1147 1429 1148 1433
rect 1142 1428 1148 1429
rect 1294 1433 1300 1434
rect 1294 1429 1295 1433
rect 1299 1429 1300 1433
rect 1294 1428 1300 1429
rect 1446 1433 1452 1434
rect 1446 1429 1447 1433
rect 1451 1429 1452 1433
rect 1446 1428 1452 1429
rect 1598 1433 1604 1434
rect 1598 1429 1599 1433
rect 1603 1429 1604 1433
rect 1598 1428 1604 1429
rect 1734 1433 1740 1434
rect 1734 1429 1735 1433
rect 1739 1429 1740 1433
rect 1862 1432 1863 1436
rect 1867 1432 1868 1436
rect 1959 1435 1965 1436
rect 1959 1434 1960 1435
rect 1949 1432 1960 1434
rect 1862 1431 1868 1432
rect 1959 1431 1960 1432
rect 1964 1431 1965 1435
rect 2103 1435 2109 1436
rect 2103 1434 2104 1435
rect 2077 1432 2104 1434
rect 1959 1430 1965 1431
rect 2103 1431 2104 1432
rect 2108 1431 2109 1435
rect 2234 1435 2240 1436
rect 2234 1434 2235 1435
rect 2229 1432 2235 1434
rect 2103 1430 2109 1431
rect 2234 1431 2235 1432
rect 2239 1431 2240 1435
rect 2695 1435 2701 1436
rect 2695 1434 2696 1435
rect 2669 1432 2696 1434
rect 2234 1430 2240 1431
rect 2242 1431 2248 1432
rect 1734 1428 1740 1429
rect 2242 1427 2243 1431
rect 2247 1430 2248 1431
rect 2695 1431 2696 1432
rect 2700 1431 2701 1435
rect 2826 1435 2832 1436
rect 2826 1434 2827 1435
rect 2821 1432 2827 1434
rect 2695 1430 2701 1431
rect 2826 1431 2827 1432
rect 2831 1431 2832 1435
rect 3199 1435 3205 1436
rect 3199 1434 3200 1435
rect 3157 1432 3200 1434
rect 2826 1430 2832 1431
rect 3199 1431 3200 1432
rect 3204 1431 3205 1435
rect 3574 1432 3575 1436
rect 3579 1432 3580 1436
rect 3199 1430 3205 1431
rect 3207 1431 3213 1432
rect 3574 1431 3580 1432
rect 2247 1428 2337 1430
rect 2247 1427 2248 1428
rect 2242 1426 2248 1427
rect 3207 1427 3208 1431
rect 3212 1430 3213 1431
rect 3212 1428 3297 1430
rect 3212 1427 3213 1428
rect 3207 1426 3213 1427
rect 110 1420 116 1421
rect 1822 1420 1828 1421
rect 110 1416 111 1420
rect 115 1416 116 1420
rect 330 1419 336 1420
rect 330 1418 331 1419
rect 309 1416 331 1418
rect 110 1415 116 1416
rect 330 1415 331 1416
rect 335 1415 336 1419
rect 455 1419 461 1420
rect 455 1418 456 1419
rect 437 1416 456 1418
rect 330 1414 336 1415
rect 455 1415 456 1416
rect 460 1415 461 1419
rect 759 1419 765 1420
rect 759 1418 760 1419
rect 725 1416 760 1418
rect 455 1414 461 1415
rect 759 1415 760 1416
rect 764 1415 765 1419
rect 1375 1419 1381 1420
rect 1375 1418 1376 1419
rect 1349 1416 1376 1418
rect 759 1414 765 1415
rect 1079 1415 1085 1416
rect 1079 1411 1080 1415
rect 1084 1414 1085 1415
rect 1375 1415 1376 1416
rect 1380 1415 1381 1419
rect 1527 1419 1533 1420
rect 1527 1418 1528 1419
rect 1501 1416 1528 1418
rect 1375 1414 1381 1415
rect 1527 1415 1528 1416
rect 1532 1415 1533 1419
rect 1807 1419 1813 1420
rect 1807 1418 1808 1419
rect 1789 1416 1808 1418
rect 1527 1414 1533 1415
rect 1807 1415 1808 1416
rect 1812 1415 1813 1419
rect 1822 1416 1823 1420
rect 1827 1416 1828 1420
rect 1822 1415 1828 1416
rect 1862 1419 1868 1420
rect 1862 1415 1863 1419
rect 1867 1415 1868 1419
rect 2866 1419 2872 1420
rect 2380 1416 2473 1418
rect 1807 1414 1813 1415
rect 1862 1414 1868 1415
rect 2378 1415 2384 1416
rect 1084 1412 1161 1414
rect 1084 1411 1085 1412
rect 1079 1410 1085 1411
rect 2378 1411 2379 1415
rect 2383 1411 2384 1415
rect 2866 1415 2867 1419
rect 2871 1418 2872 1419
rect 3574 1419 3580 1420
rect 2871 1416 2945 1418
rect 2871 1415 2872 1416
rect 2866 1414 2872 1415
rect 3574 1415 3575 1419
rect 3579 1415 3580 1419
rect 3574 1414 3580 1415
rect 2378 1410 2384 1411
rect 1886 1409 1892 1410
rect 1886 1405 1887 1409
rect 1891 1405 1892 1409
rect 1886 1404 1892 1405
rect 2014 1409 2020 1410
rect 2014 1405 2015 1409
rect 2019 1405 2020 1409
rect 2014 1404 2020 1405
rect 2166 1409 2172 1410
rect 2166 1405 2167 1409
rect 2171 1405 2172 1409
rect 2166 1404 2172 1405
rect 2310 1409 2316 1410
rect 2310 1405 2311 1409
rect 2315 1405 2316 1409
rect 2310 1404 2316 1405
rect 2454 1409 2460 1410
rect 2454 1405 2455 1409
rect 2459 1405 2460 1409
rect 2454 1404 2460 1405
rect 2606 1409 2612 1410
rect 2606 1405 2607 1409
rect 2611 1405 2612 1409
rect 2606 1404 2612 1405
rect 2758 1409 2764 1410
rect 2758 1405 2759 1409
rect 2763 1405 2764 1409
rect 2758 1404 2764 1405
rect 2926 1409 2932 1410
rect 2926 1405 2927 1409
rect 2931 1405 2932 1409
rect 2926 1404 2932 1405
rect 3094 1409 3100 1410
rect 3094 1405 3095 1409
rect 3099 1405 3100 1409
rect 3094 1404 3100 1405
rect 3270 1409 3276 1410
rect 3270 1405 3271 1409
rect 3275 1405 3276 1409
rect 3270 1404 3276 1405
rect 3454 1409 3460 1410
rect 3454 1405 3455 1409
rect 3459 1405 3460 1409
rect 3454 1404 3460 1405
rect 110 1403 116 1404
rect 110 1399 111 1403
rect 115 1399 116 1403
rect 110 1398 116 1399
rect 738 1403 744 1404
rect 738 1399 739 1403
rect 743 1402 744 1403
rect 898 1403 904 1404
rect 743 1400 841 1402
rect 743 1399 744 1400
rect 738 1398 744 1399
rect 898 1399 899 1403
rect 903 1402 904 1403
rect 1718 1403 1724 1404
rect 1718 1402 1719 1403
rect 903 1400 1001 1402
rect 1649 1400 1719 1402
rect 903 1399 904 1400
rect 898 1398 904 1399
rect 1718 1399 1719 1400
rect 1723 1399 1724 1403
rect 1718 1398 1724 1399
rect 1822 1403 1828 1404
rect 1822 1399 1823 1403
rect 1827 1399 1828 1403
rect 1822 1398 1828 1399
rect 3498 1403 3509 1404
rect 3498 1399 3499 1403
rect 3503 1399 3504 1403
rect 3508 1399 3509 1403
rect 3498 1398 3509 1399
rect 246 1393 252 1394
rect 246 1389 247 1393
rect 251 1389 252 1393
rect 246 1388 252 1389
rect 374 1393 380 1394
rect 374 1389 375 1393
rect 379 1389 380 1393
rect 374 1388 380 1389
rect 510 1393 516 1394
rect 510 1389 511 1393
rect 515 1389 516 1393
rect 510 1388 516 1389
rect 662 1393 668 1394
rect 662 1389 663 1393
rect 667 1389 668 1393
rect 662 1388 668 1389
rect 822 1393 828 1394
rect 822 1389 823 1393
rect 827 1389 828 1393
rect 822 1388 828 1389
rect 982 1393 988 1394
rect 982 1389 983 1393
rect 987 1389 988 1393
rect 982 1388 988 1389
rect 1134 1393 1140 1394
rect 1134 1389 1135 1393
rect 1139 1389 1140 1393
rect 1134 1388 1140 1389
rect 1286 1393 1292 1394
rect 1286 1389 1287 1393
rect 1291 1389 1292 1393
rect 1286 1388 1292 1389
rect 1438 1393 1444 1394
rect 1438 1389 1439 1393
rect 1443 1389 1444 1393
rect 1438 1388 1444 1389
rect 1590 1393 1596 1394
rect 1590 1389 1591 1393
rect 1595 1389 1596 1393
rect 1590 1388 1596 1389
rect 1726 1393 1732 1394
rect 1726 1389 1727 1393
rect 1731 1389 1732 1393
rect 1726 1388 1732 1389
rect 542 1387 548 1388
rect 542 1383 543 1387
rect 547 1386 548 1387
rect 559 1387 565 1388
rect 559 1386 560 1387
rect 547 1384 560 1386
rect 547 1383 548 1384
rect 542 1382 548 1383
rect 559 1383 560 1384
rect 564 1383 565 1387
rect 559 1382 565 1383
rect 1886 1375 1892 1376
rect 350 1371 356 1372
rect 350 1367 351 1371
rect 355 1367 356 1371
rect 350 1366 356 1367
rect 438 1371 444 1372
rect 438 1367 439 1371
rect 443 1367 444 1371
rect 438 1366 444 1367
rect 526 1371 532 1372
rect 526 1367 527 1371
rect 531 1367 532 1371
rect 526 1366 532 1367
rect 622 1371 628 1372
rect 622 1367 623 1371
rect 627 1367 628 1371
rect 622 1366 628 1367
rect 726 1371 732 1372
rect 726 1367 727 1371
rect 731 1367 732 1371
rect 726 1366 732 1367
rect 846 1371 852 1372
rect 846 1367 847 1371
rect 851 1367 852 1371
rect 846 1366 852 1367
rect 982 1371 988 1372
rect 982 1367 983 1371
rect 987 1367 988 1371
rect 982 1366 988 1367
rect 1126 1371 1132 1372
rect 1126 1367 1127 1371
rect 1131 1367 1132 1371
rect 1126 1366 1132 1367
rect 1278 1371 1284 1372
rect 1278 1367 1279 1371
rect 1283 1367 1284 1371
rect 1278 1366 1284 1367
rect 1430 1371 1436 1372
rect 1430 1367 1431 1371
rect 1435 1367 1436 1371
rect 1430 1366 1436 1367
rect 1590 1371 1596 1372
rect 1590 1367 1591 1371
rect 1595 1367 1596 1371
rect 1590 1366 1596 1367
rect 1726 1371 1732 1372
rect 1726 1367 1727 1371
rect 1731 1367 1732 1371
rect 1886 1371 1887 1375
rect 1891 1371 1892 1375
rect 1886 1370 1892 1371
rect 2142 1375 2148 1376
rect 2142 1371 2143 1375
rect 2147 1371 2148 1375
rect 2142 1370 2148 1371
rect 2390 1375 2396 1376
rect 2390 1371 2391 1375
rect 2395 1371 2396 1375
rect 2390 1370 2396 1371
rect 2622 1375 2628 1376
rect 2622 1371 2623 1375
rect 2627 1371 2628 1375
rect 2622 1370 2628 1371
rect 2846 1375 2852 1376
rect 2846 1371 2847 1375
rect 2851 1371 2852 1375
rect 2846 1370 2852 1371
rect 3062 1375 3068 1376
rect 3062 1371 3063 1375
rect 3067 1371 3068 1375
rect 3062 1370 3068 1371
rect 3270 1375 3276 1376
rect 3270 1371 3271 1375
rect 3275 1371 3276 1375
rect 3270 1370 3276 1371
rect 3478 1375 3484 1376
rect 3478 1371 3479 1375
rect 3483 1371 3484 1375
rect 3478 1370 3484 1371
rect 1726 1366 1732 1367
rect 2518 1367 2524 1368
rect 2518 1366 2519 1367
rect 1862 1365 1868 1366
rect 690 1363 696 1364
rect 690 1362 691 1363
rect 110 1361 116 1362
rect 110 1357 111 1361
rect 115 1357 116 1361
rect 681 1360 691 1362
rect 690 1359 691 1360
rect 695 1359 696 1363
rect 690 1358 696 1359
rect 1202 1363 1208 1364
rect 1202 1359 1203 1363
rect 1207 1362 1208 1363
rect 1678 1363 1684 1364
rect 1678 1362 1679 1363
rect 1207 1360 1297 1362
rect 1649 1360 1679 1362
rect 1207 1359 1208 1360
rect 1202 1358 1208 1359
rect 1678 1359 1679 1360
rect 1683 1359 1684 1363
rect 1678 1358 1684 1359
rect 1822 1361 1828 1362
rect 110 1356 116 1357
rect 1822 1357 1823 1361
rect 1827 1357 1828 1361
rect 1862 1361 1863 1365
rect 1867 1361 1868 1365
rect 2449 1364 2519 1366
rect 2518 1363 2519 1364
rect 2523 1363 2524 1367
rect 2518 1362 2524 1363
rect 2970 1367 2976 1368
rect 2970 1363 2971 1367
rect 2975 1366 2976 1367
rect 3263 1367 3269 1368
rect 2975 1364 3081 1366
rect 2975 1363 2976 1364
rect 2970 1362 2976 1363
rect 3263 1363 3264 1367
rect 3268 1366 3269 1367
rect 3268 1364 3289 1366
rect 3574 1365 3580 1366
rect 3268 1363 3269 1364
rect 3263 1362 3269 1363
rect 1862 1360 1868 1361
rect 3574 1361 3575 1365
rect 3579 1361 3580 1365
rect 3574 1360 3580 1361
rect 1822 1356 1828 1357
rect 1870 1351 1876 1352
rect 1862 1348 1868 1349
rect 431 1347 437 1348
rect 431 1346 432 1347
rect 110 1344 116 1345
rect 413 1344 432 1346
rect 110 1340 111 1344
rect 115 1340 116 1344
rect 431 1343 432 1344
rect 436 1343 437 1347
rect 506 1347 512 1348
rect 506 1346 507 1347
rect 501 1344 507 1346
rect 431 1342 437 1343
rect 506 1343 507 1344
rect 511 1343 512 1347
rect 506 1342 512 1343
rect 514 1347 520 1348
rect 514 1343 515 1347
rect 519 1346 520 1347
rect 695 1347 701 1348
rect 519 1344 553 1346
rect 519 1343 520 1344
rect 514 1342 520 1343
rect 695 1343 696 1347
rect 700 1346 701 1347
rect 794 1347 800 1348
rect 700 1344 753 1346
rect 700 1343 701 1344
rect 695 1342 701 1343
rect 794 1343 795 1347
rect 799 1346 800 1347
rect 1119 1347 1125 1348
rect 1119 1346 1120 1347
rect 799 1344 873 1346
rect 1045 1344 1120 1346
rect 799 1343 800 1344
rect 794 1342 800 1343
rect 1119 1343 1120 1344
rect 1124 1343 1125 1347
rect 1271 1347 1277 1348
rect 1271 1346 1272 1347
rect 1189 1344 1272 1346
rect 1119 1342 1125 1343
rect 1271 1343 1272 1344
rect 1276 1343 1277 1347
rect 1583 1347 1589 1348
rect 1583 1346 1584 1347
rect 1493 1344 1584 1346
rect 1271 1342 1277 1343
rect 1583 1343 1584 1344
rect 1588 1343 1589 1347
rect 1583 1342 1589 1343
rect 1719 1347 1725 1348
rect 1719 1343 1720 1347
rect 1724 1346 1725 1347
rect 1724 1344 1753 1346
rect 1822 1344 1828 1345
rect 1724 1343 1725 1344
rect 1719 1342 1725 1343
rect 110 1339 116 1340
rect 1822 1340 1823 1344
rect 1827 1340 1828 1344
rect 1862 1344 1863 1348
rect 1867 1344 1868 1348
rect 1870 1347 1871 1351
rect 1875 1350 1876 1351
rect 2383 1351 2389 1352
rect 2383 1350 2384 1351
rect 1875 1348 1913 1350
rect 2205 1348 2384 1350
rect 1875 1347 1876 1348
rect 1870 1346 1876 1347
rect 2383 1347 2384 1348
rect 2388 1347 2389 1351
rect 2383 1346 2389 1347
rect 2462 1351 2468 1352
rect 2462 1347 2463 1351
rect 2467 1350 2468 1351
rect 3055 1351 3061 1352
rect 3055 1350 3056 1351
rect 2467 1348 2649 1350
rect 2909 1348 3056 1350
rect 2467 1347 2468 1348
rect 2462 1346 2468 1347
rect 3055 1347 3056 1348
rect 3060 1347 3061 1351
rect 3055 1346 3061 1347
rect 3471 1351 3477 1352
rect 3471 1347 3472 1351
rect 3476 1350 3477 1351
rect 3476 1348 3505 1350
rect 3574 1348 3580 1349
rect 3476 1347 3477 1348
rect 3471 1346 3477 1347
rect 1862 1343 1868 1344
rect 3574 1344 3575 1348
rect 3579 1344 3580 1348
rect 3574 1343 3580 1344
rect 1822 1339 1828 1340
rect 1894 1335 1900 1336
rect 358 1331 364 1332
rect 358 1327 359 1331
rect 363 1327 364 1331
rect 358 1326 364 1327
rect 446 1331 452 1332
rect 446 1327 447 1331
rect 451 1327 452 1331
rect 446 1326 452 1327
rect 534 1331 540 1332
rect 534 1327 535 1331
rect 539 1327 540 1331
rect 534 1326 540 1327
rect 630 1331 636 1332
rect 630 1327 631 1331
rect 635 1327 636 1331
rect 630 1326 636 1327
rect 734 1331 740 1332
rect 734 1327 735 1331
rect 739 1327 740 1331
rect 734 1326 740 1327
rect 854 1331 860 1332
rect 854 1327 855 1331
rect 859 1327 860 1331
rect 854 1326 860 1327
rect 990 1331 996 1332
rect 990 1327 991 1331
rect 995 1327 996 1331
rect 990 1326 996 1327
rect 1134 1331 1140 1332
rect 1134 1327 1135 1331
rect 1139 1327 1140 1331
rect 1134 1326 1140 1327
rect 1286 1331 1292 1332
rect 1286 1327 1287 1331
rect 1291 1327 1292 1331
rect 1286 1326 1292 1327
rect 1438 1331 1444 1332
rect 1438 1327 1439 1331
rect 1443 1327 1444 1331
rect 1438 1326 1444 1327
rect 1598 1331 1604 1332
rect 1598 1327 1599 1331
rect 1603 1327 1604 1331
rect 1598 1326 1604 1327
rect 1734 1331 1740 1332
rect 1734 1327 1735 1331
rect 1739 1327 1740 1331
rect 1894 1331 1895 1335
rect 1899 1331 1900 1335
rect 1894 1330 1900 1331
rect 2150 1335 2156 1336
rect 2150 1331 2151 1335
rect 2155 1331 2156 1335
rect 2150 1330 2156 1331
rect 2398 1335 2404 1336
rect 2398 1331 2399 1335
rect 2403 1331 2404 1335
rect 2398 1330 2404 1331
rect 2630 1335 2636 1336
rect 2630 1331 2631 1335
rect 2635 1331 2636 1335
rect 2630 1330 2636 1331
rect 2854 1335 2860 1336
rect 2854 1331 2855 1335
rect 2859 1331 2860 1335
rect 2854 1330 2860 1331
rect 3070 1335 3076 1336
rect 3070 1331 3071 1335
rect 3075 1331 3076 1335
rect 3070 1330 3076 1331
rect 3278 1335 3284 1336
rect 3278 1331 3279 1335
rect 3283 1331 3284 1335
rect 3278 1330 3284 1331
rect 3486 1335 3492 1336
rect 3486 1331 3487 1335
rect 3491 1331 3492 1335
rect 3486 1330 3492 1331
rect 1734 1326 1740 1327
rect 542 1323 548 1324
rect 366 1319 373 1320
rect 366 1315 367 1319
rect 372 1315 373 1319
rect 366 1314 373 1315
rect 431 1319 437 1320
rect 431 1315 432 1319
rect 436 1318 437 1319
rect 455 1319 461 1320
rect 455 1318 456 1319
rect 436 1316 456 1318
rect 436 1315 437 1316
rect 431 1314 437 1315
rect 455 1315 456 1316
rect 460 1315 461 1319
rect 542 1319 543 1323
rect 547 1322 548 1323
rect 1903 1323 1912 1324
rect 547 1321 549 1322
rect 542 1318 544 1319
rect 543 1317 544 1318
rect 548 1317 549 1321
rect 543 1316 549 1317
rect 639 1319 645 1320
rect 455 1314 461 1315
rect 639 1315 640 1319
rect 644 1318 645 1319
rect 695 1319 701 1320
rect 695 1318 696 1319
rect 644 1316 696 1318
rect 644 1315 645 1316
rect 639 1314 645 1315
rect 695 1315 696 1316
rect 700 1315 701 1319
rect 695 1314 701 1315
rect 743 1319 749 1320
rect 743 1315 744 1319
rect 748 1318 749 1319
rect 794 1319 800 1320
rect 794 1318 795 1319
rect 748 1316 795 1318
rect 748 1315 749 1316
rect 743 1314 749 1315
rect 794 1315 795 1316
rect 799 1315 800 1319
rect 794 1314 800 1315
rect 863 1319 869 1320
rect 863 1315 864 1319
rect 868 1318 869 1319
rect 898 1319 904 1320
rect 898 1318 899 1319
rect 868 1316 899 1318
rect 868 1315 869 1316
rect 863 1314 869 1315
rect 898 1315 899 1316
rect 903 1315 904 1319
rect 898 1314 904 1315
rect 999 1319 1005 1320
rect 999 1315 1000 1319
rect 1004 1318 1005 1319
rect 1026 1319 1032 1320
rect 1026 1318 1027 1319
rect 1004 1316 1027 1318
rect 1004 1315 1005 1316
rect 999 1314 1005 1315
rect 1026 1315 1027 1316
rect 1031 1315 1032 1319
rect 1026 1314 1032 1315
rect 1119 1319 1125 1320
rect 1119 1315 1120 1319
rect 1124 1318 1125 1319
rect 1143 1319 1149 1320
rect 1143 1318 1144 1319
rect 1124 1316 1144 1318
rect 1124 1315 1125 1316
rect 1119 1314 1125 1315
rect 1143 1315 1144 1316
rect 1148 1315 1149 1319
rect 1143 1314 1149 1315
rect 1271 1319 1277 1320
rect 1271 1315 1272 1319
rect 1276 1318 1277 1319
rect 1295 1319 1301 1320
rect 1295 1318 1296 1319
rect 1276 1316 1296 1318
rect 1276 1315 1277 1316
rect 1271 1314 1277 1315
rect 1295 1315 1296 1316
rect 1300 1315 1301 1319
rect 1295 1314 1301 1315
rect 1447 1319 1456 1320
rect 1447 1315 1448 1319
rect 1455 1315 1456 1319
rect 1447 1314 1456 1315
rect 1583 1319 1589 1320
rect 1583 1315 1584 1319
rect 1588 1318 1589 1319
rect 1607 1319 1613 1320
rect 1607 1318 1608 1319
rect 1588 1316 1608 1318
rect 1588 1315 1589 1316
rect 1583 1314 1589 1315
rect 1607 1315 1608 1316
rect 1612 1315 1613 1319
rect 1607 1314 1613 1315
rect 1718 1319 1724 1320
rect 1718 1315 1719 1319
rect 1723 1318 1724 1319
rect 1743 1319 1749 1320
rect 1743 1318 1744 1319
rect 1723 1316 1744 1318
rect 1723 1315 1724 1316
rect 1718 1314 1724 1315
rect 1743 1315 1744 1316
rect 1748 1315 1749 1319
rect 1903 1319 1904 1323
rect 1911 1319 1912 1323
rect 1903 1318 1912 1319
rect 2159 1323 2165 1324
rect 2159 1319 2160 1323
rect 2164 1322 2165 1323
rect 2378 1323 2384 1324
rect 2378 1322 2379 1323
rect 2164 1320 2379 1322
rect 2164 1319 2165 1320
rect 2159 1318 2165 1319
rect 2378 1319 2379 1320
rect 2383 1319 2384 1323
rect 2378 1318 2384 1319
rect 2407 1323 2413 1324
rect 2407 1319 2408 1323
rect 2412 1322 2413 1323
rect 2462 1323 2468 1324
rect 2462 1322 2463 1323
rect 2412 1320 2463 1322
rect 2412 1319 2413 1320
rect 2407 1318 2413 1319
rect 2462 1319 2463 1320
rect 2467 1319 2468 1323
rect 2462 1318 2468 1319
rect 2639 1323 2645 1324
rect 2639 1319 2640 1323
rect 2644 1322 2645 1323
rect 2682 1323 2688 1324
rect 2682 1322 2683 1323
rect 2644 1320 2683 1322
rect 2644 1319 2645 1320
rect 2639 1318 2645 1319
rect 2682 1319 2683 1320
rect 2687 1319 2688 1323
rect 2682 1318 2688 1319
rect 2863 1323 2872 1324
rect 2863 1319 2864 1323
rect 2871 1319 2872 1323
rect 2863 1318 2872 1319
rect 3055 1323 3061 1324
rect 3055 1319 3056 1323
rect 3060 1322 3061 1323
rect 3079 1323 3085 1324
rect 3079 1322 3080 1323
rect 3060 1320 3080 1322
rect 3060 1319 3061 1320
rect 3055 1318 3061 1319
rect 3079 1319 3080 1320
rect 3084 1319 3085 1323
rect 3079 1318 3085 1319
rect 3287 1323 3293 1324
rect 3287 1319 3288 1323
rect 3292 1322 3293 1323
rect 3418 1323 3424 1324
rect 3418 1322 3419 1323
rect 3292 1320 3419 1322
rect 3292 1319 3293 1320
rect 3287 1318 3293 1319
rect 3418 1319 3419 1320
rect 3423 1319 3424 1323
rect 3418 1318 3424 1319
rect 3495 1323 3504 1324
rect 3495 1319 3496 1323
rect 3503 1319 3504 1323
rect 3495 1318 3504 1319
rect 1743 1314 1749 1315
rect 1935 1311 1941 1312
rect 463 1307 469 1308
rect 463 1303 464 1307
rect 468 1306 469 1307
rect 506 1307 512 1308
rect 506 1306 507 1307
rect 468 1304 507 1306
rect 468 1303 469 1304
rect 463 1302 469 1303
rect 506 1303 507 1304
rect 511 1303 512 1307
rect 506 1302 512 1303
rect 519 1307 525 1308
rect 519 1303 520 1307
rect 524 1306 525 1307
rect 551 1307 557 1308
rect 551 1306 552 1307
rect 524 1304 552 1306
rect 524 1303 525 1304
rect 519 1302 525 1303
rect 551 1303 552 1304
rect 556 1303 557 1307
rect 551 1302 557 1303
rect 607 1307 613 1308
rect 607 1303 608 1307
rect 612 1306 613 1307
rect 639 1307 645 1308
rect 639 1306 640 1307
rect 612 1304 640 1306
rect 612 1303 613 1304
rect 607 1302 613 1303
rect 639 1303 640 1304
rect 644 1303 645 1307
rect 639 1302 645 1303
rect 695 1307 701 1308
rect 695 1303 696 1307
rect 700 1306 701 1307
rect 727 1307 733 1308
rect 727 1306 728 1307
rect 700 1304 728 1306
rect 700 1303 701 1304
rect 695 1302 701 1303
rect 727 1303 728 1304
rect 732 1303 733 1307
rect 727 1302 733 1303
rect 783 1307 789 1308
rect 783 1303 784 1307
rect 788 1306 789 1307
rect 839 1307 845 1308
rect 839 1306 840 1307
rect 788 1304 840 1306
rect 788 1303 789 1304
rect 783 1302 789 1303
rect 839 1303 840 1304
rect 844 1303 845 1307
rect 839 1302 845 1303
rect 975 1307 981 1308
rect 975 1303 976 1307
rect 980 1306 981 1307
rect 1058 1307 1064 1308
rect 1058 1306 1059 1307
rect 980 1304 1059 1306
rect 980 1303 981 1304
rect 975 1302 981 1303
rect 1058 1303 1059 1304
rect 1063 1303 1064 1307
rect 1058 1302 1064 1303
rect 1143 1307 1149 1308
rect 1143 1303 1144 1307
rect 1148 1306 1149 1307
rect 1230 1307 1236 1308
rect 1230 1306 1231 1307
rect 1148 1304 1231 1306
rect 1148 1303 1149 1304
rect 1143 1302 1149 1303
rect 1230 1303 1231 1304
rect 1235 1303 1236 1307
rect 1230 1302 1236 1303
rect 1335 1307 1341 1308
rect 1335 1303 1336 1307
rect 1340 1306 1341 1307
rect 1394 1307 1400 1308
rect 1394 1306 1395 1307
rect 1340 1304 1395 1306
rect 1340 1303 1341 1304
rect 1335 1302 1341 1303
rect 1394 1303 1395 1304
rect 1399 1303 1400 1307
rect 1394 1302 1400 1303
rect 1542 1307 1549 1308
rect 1542 1303 1543 1307
rect 1548 1303 1549 1307
rect 1542 1302 1549 1303
rect 1719 1307 1725 1308
rect 1719 1303 1720 1307
rect 1724 1306 1725 1307
rect 1743 1307 1749 1308
rect 1743 1306 1744 1307
rect 1724 1304 1744 1306
rect 1724 1303 1725 1304
rect 1719 1302 1725 1303
rect 1743 1303 1744 1304
rect 1748 1303 1749 1307
rect 1935 1307 1936 1311
rect 1940 1310 1941 1311
rect 2030 1311 2036 1312
rect 2030 1310 2031 1311
rect 1940 1308 2031 1310
rect 1940 1307 1941 1308
rect 1935 1306 1941 1307
rect 2030 1307 2031 1308
rect 2035 1307 2036 1311
rect 2030 1306 2036 1307
rect 2119 1311 2125 1312
rect 2119 1307 2120 1311
rect 2124 1310 2125 1311
rect 2207 1311 2213 1312
rect 2207 1310 2208 1311
rect 2124 1308 2208 1310
rect 2124 1307 2125 1308
rect 2119 1306 2125 1307
rect 2207 1307 2208 1308
rect 2212 1307 2213 1311
rect 2207 1306 2213 1307
rect 2230 1311 2236 1312
rect 2230 1307 2231 1311
rect 2235 1310 2236 1311
rect 2295 1311 2301 1312
rect 2295 1310 2296 1311
rect 2235 1308 2296 1310
rect 2235 1307 2236 1308
rect 2230 1306 2236 1307
rect 2295 1307 2296 1308
rect 2300 1307 2301 1311
rect 2295 1306 2301 1307
rect 2383 1311 2389 1312
rect 2383 1307 2384 1311
rect 2388 1310 2389 1311
rect 2463 1311 2469 1312
rect 2463 1310 2464 1311
rect 2388 1308 2464 1310
rect 2388 1307 2389 1308
rect 2383 1306 2389 1307
rect 2463 1307 2464 1308
rect 2468 1307 2469 1311
rect 2463 1306 2469 1307
rect 2631 1311 2637 1312
rect 2631 1307 2632 1311
rect 2636 1310 2637 1311
rect 2718 1311 2724 1312
rect 2718 1310 2719 1311
rect 2636 1308 2719 1310
rect 2636 1307 2637 1308
rect 2631 1306 2637 1307
rect 2718 1307 2719 1308
rect 2723 1307 2724 1311
rect 2718 1306 2724 1307
rect 2799 1311 2805 1312
rect 2799 1307 2800 1311
rect 2804 1310 2805 1311
rect 2814 1311 2820 1312
rect 2814 1310 2815 1311
rect 2804 1308 2815 1310
rect 2804 1307 2805 1308
rect 2799 1306 2805 1307
rect 2814 1307 2815 1308
rect 2819 1307 2820 1311
rect 2814 1306 2820 1307
rect 2967 1311 2976 1312
rect 2967 1307 2968 1311
rect 2975 1307 2976 1311
rect 2967 1306 2976 1307
rect 3055 1311 3061 1312
rect 3055 1307 3056 1311
rect 3060 1310 3061 1311
rect 3143 1311 3149 1312
rect 3143 1310 3144 1311
rect 3060 1308 3144 1310
rect 3060 1307 3061 1308
rect 3055 1306 3061 1307
rect 3143 1307 3144 1308
rect 3148 1307 3149 1311
rect 3143 1306 3149 1307
rect 3231 1311 3237 1312
rect 3231 1307 3232 1311
rect 3236 1310 3237 1311
rect 3327 1311 3333 1312
rect 3327 1310 3328 1311
rect 3236 1308 3328 1310
rect 3236 1307 3237 1308
rect 3231 1306 3237 1307
rect 3327 1307 3328 1308
rect 3332 1307 3333 1311
rect 3327 1306 3333 1307
rect 3471 1311 3477 1312
rect 3471 1307 3472 1311
rect 3476 1310 3477 1311
rect 3495 1311 3501 1312
rect 3495 1310 3496 1311
rect 3476 1308 3496 1310
rect 3476 1307 3477 1308
rect 3471 1306 3477 1307
rect 3495 1307 3496 1308
rect 3500 1307 3501 1311
rect 3495 1306 3501 1307
rect 1743 1302 1749 1303
rect 1926 1301 1932 1302
rect 454 1297 460 1298
rect 454 1293 455 1297
rect 459 1293 460 1297
rect 454 1292 460 1293
rect 542 1297 548 1298
rect 542 1293 543 1297
rect 547 1293 548 1297
rect 542 1292 548 1293
rect 630 1297 636 1298
rect 630 1293 631 1297
rect 635 1293 636 1297
rect 630 1292 636 1293
rect 718 1297 724 1298
rect 718 1293 719 1297
rect 723 1293 724 1297
rect 718 1292 724 1293
rect 830 1297 836 1298
rect 830 1293 831 1297
rect 835 1293 836 1297
rect 830 1292 836 1293
rect 966 1297 972 1298
rect 966 1293 967 1297
rect 971 1293 972 1297
rect 966 1292 972 1293
rect 1134 1297 1140 1298
rect 1134 1293 1135 1297
rect 1139 1293 1140 1297
rect 1134 1292 1140 1293
rect 1326 1297 1332 1298
rect 1326 1293 1327 1297
rect 1331 1293 1332 1297
rect 1326 1292 1332 1293
rect 1534 1297 1540 1298
rect 1534 1293 1535 1297
rect 1539 1293 1540 1297
rect 1534 1292 1540 1293
rect 1734 1297 1740 1298
rect 1734 1293 1735 1297
rect 1739 1293 1740 1297
rect 1926 1297 1927 1301
rect 1931 1297 1932 1301
rect 1926 1296 1932 1297
rect 2110 1301 2116 1302
rect 2110 1297 2111 1301
rect 2115 1297 2116 1301
rect 2110 1296 2116 1297
rect 2286 1301 2292 1302
rect 2286 1297 2287 1301
rect 2291 1297 2292 1301
rect 2286 1296 2292 1297
rect 2454 1301 2460 1302
rect 2454 1297 2455 1301
rect 2459 1297 2460 1301
rect 2454 1296 2460 1297
rect 2622 1301 2628 1302
rect 2622 1297 2623 1301
rect 2627 1297 2628 1301
rect 2622 1296 2628 1297
rect 2790 1301 2796 1302
rect 2790 1297 2791 1301
rect 2795 1297 2796 1301
rect 2790 1296 2796 1297
rect 2958 1301 2964 1302
rect 2958 1297 2959 1301
rect 2963 1297 2964 1301
rect 2958 1296 2964 1297
rect 3134 1301 3140 1302
rect 3134 1297 3135 1301
rect 3139 1297 3140 1301
rect 3134 1296 3140 1297
rect 3318 1301 3324 1302
rect 3318 1297 3319 1301
rect 3323 1297 3324 1301
rect 3318 1296 3324 1297
rect 3486 1301 3492 1302
rect 3486 1297 3487 1301
rect 3491 1297 3492 1301
rect 3486 1296 3492 1297
rect 1734 1292 1740 1293
rect 1862 1288 1868 1289
rect 3574 1288 3580 1289
rect 110 1284 116 1285
rect 1822 1284 1828 1285
rect 110 1280 111 1284
rect 115 1280 116 1284
rect 519 1283 525 1284
rect 519 1282 520 1283
rect 509 1280 520 1282
rect 110 1279 116 1280
rect 519 1279 520 1280
rect 524 1279 525 1283
rect 607 1283 613 1284
rect 607 1282 608 1283
rect 597 1280 608 1282
rect 519 1278 525 1279
rect 607 1279 608 1280
rect 612 1279 613 1283
rect 695 1283 701 1284
rect 695 1282 696 1283
rect 685 1280 696 1282
rect 607 1278 613 1279
rect 695 1279 696 1280
rect 700 1279 701 1283
rect 783 1283 789 1284
rect 783 1282 784 1283
rect 773 1280 784 1282
rect 695 1278 701 1279
rect 783 1279 784 1280
rect 788 1279 789 1283
rect 1026 1283 1032 1284
rect 1026 1282 1027 1283
rect 1021 1280 1027 1282
rect 783 1278 789 1279
rect 1026 1279 1027 1280
rect 1031 1279 1032 1283
rect 1822 1280 1823 1284
rect 1827 1280 1828 1284
rect 1862 1284 1863 1288
rect 1867 1284 1868 1288
rect 2682 1287 2688 1288
rect 2682 1286 2683 1287
rect 2677 1284 2683 1286
rect 1862 1283 1868 1284
rect 1906 1283 1912 1284
rect 1026 1278 1032 1279
rect 1058 1279 1064 1280
rect 1058 1275 1059 1279
rect 1063 1278 1064 1279
rect 1230 1279 1236 1280
rect 1063 1276 1153 1278
rect 1063 1275 1064 1276
rect 1058 1274 1064 1275
rect 1230 1275 1231 1279
rect 1235 1278 1236 1279
rect 1394 1279 1400 1280
rect 1822 1279 1828 1280
rect 1906 1279 1907 1283
rect 1911 1282 1912 1283
rect 2030 1283 2036 1284
rect 1911 1280 1945 1282
rect 1911 1279 1912 1280
rect 1235 1276 1345 1278
rect 1235 1275 1236 1276
rect 1230 1274 1236 1275
rect 1394 1275 1395 1279
rect 1399 1278 1400 1279
rect 1906 1278 1912 1279
rect 2030 1279 2031 1283
rect 2035 1282 2036 1283
rect 2207 1283 2213 1284
rect 2035 1280 2129 1282
rect 2035 1279 2036 1280
rect 2030 1278 2036 1279
rect 2207 1279 2208 1283
rect 2212 1282 2213 1283
rect 2682 1283 2683 1284
rect 2687 1283 2688 1287
rect 3055 1287 3061 1288
rect 3055 1286 3056 1287
rect 3013 1284 3056 1286
rect 2682 1282 2688 1283
rect 2718 1283 2724 1284
rect 2212 1280 2305 1282
rect 2212 1279 2213 1280
rect 2207 1278 2213 1279
rect 2718 1279 2719 1283
rect 2723 1282 2724 1283
rect 3055 1283 3056 1284
rect 3060 1283 3061 1287
rect 3231 1287 3237 1288
rect 3231 1286 3232 1287
rect 3189 1284 3232 1286
rect 3055 1282 3061 1283
rect 3231 1283 3232 1284
rect 3236 1283 3237 1287
rect 3574 1284 3575 1288
rect 3579 1284 3580 1288
rect 3574 1283 3580 1284
rect 3231 1282 3237 1283
rect 2723 1280 2809 1282
rect 2723 1279 2724 1280
rect 2718 1278 2724 1279
rect 1399 1276 1553 1278
rect 1399 1275 1400 1276
rect 1394 1274 1400 1275
rect 1862 1271 1868 1272
rect 110 1267 116 1268
rect 110 1263 111 1267
rect 115 1263 116 1267
rect 110 1262 116 1263
rect 830 1267 836 1268
rect 830 1263 831 1267
rect 835 1266 836 1267
rect 1626 1267 1632 1268
rect 835 1264 841 1266
rect 835 1263 836 1264
rect 830 1262 836 1263
rect 1626 1263 1627 1267
rect 1631 1266 1632 1267
rect 1822 1267 1828 1268
rect 1631 1264 1745 1266
rect 1631 1263 1632 1264
rect 1626 1262 1632 1263
rect 1822 1263 1823 1267
rect 1827 1263 1828 1267
rect 1862 1267 1863 1271
rect 1867 1267 1868 1271
rect 1862 1266 1868 1267
rect 3574 1271 3580 1272
rect 3574 1267 3575 1271
rect 3579 1267 3580 1271
rect 3574 1266 3580 1267
rect 1822 1262 1828 1263
rect 1918 1261 1924 1262
rect 446 1257 452 1258
rect 446 1253 447 1257
rect 451 1253 452 1257
rect 446 1252 452 1253
rect 534 1257 540 1258
rect 534 1253 535 1257
rect 539 1253 540 1257
rect 534 1252 540 1253
rect 622 1257 628 1258
rect 622 1253 623 1257
rect 627 1253 628 1257
rect 622 1252 628 1253
rect 710 1257 716 1258
rect 710 1253 711 1257
rect 715 1253 716 1257
rect 710 1252 716 1253
rect 822 1257 828 1258
rect 822 1253 823 1257
rect 827 1253 828 1257
rect 822 1252 828 1253
rect 958 1257 964 1258
rect 958 1253 959 1257
rect 963 1253 964 1257
rect 958 1252 964 1253
rect 1126 1257 1132 1258
rect 1126 1253 1127 1257
rect 1131 1253 1132 1257
rect 1126 1252 1132 1253
rect 1318 1257 1324 1258
rect 1318 1253 1319 1257
rect 1323 1253 1324 1257
rect 1318 1252 1324 1253
rect 1526 1257 1532 1258
rect 1526 1253 1527 1257
rect 1531 1253 1532 1257
rect 1526 1252 1532 1253
rect 1726 1257 1732 1258
rect 1726 1253 1727 1257
rect 1731 1253 1732 1257
rect 1918 1257 1919 1261
rect 1923 1257 1924 1261
rect 1918 1256 1924 1257
rect 2102 1261 2108 1262
rect 2102 1257 2103 1261
rect 2107 1257 2108 1261
rect 2102 1256 2108 1257
rect 2278 1261 2284 1262
rect 2278 1257 2279 1261
rect 2283 1257 2284 1261
rect 2278 1256 2284 1257
rect 2446 1261 2452 1262
rect 2446 1257 2447 1261
rect 2451 1257 2452 1261
rect 2446 1256 2452 1257
rect 2614 1261 2620 1262
rect 2614 1257 2615 1261
rect 2619 1257 2620 1261
rect 2614 1256 2620 1257
rect 2782 1261 2788 1262
rect 2782 1257 2783 1261
rect 2787 1257 2788 1261
rect 2782 1256 2788 1257
rect 2950 1261 2956 1262
rect 2950 1257 2951 1261
rect 2955 1257 2956 1261
rect 2950 1256 2956 1257
rect 3126 1261 3132 1262
rect 3126 1257 3127 1261
rect 3131 1257 3132 1261
rect 3126 1256 3132 1257
rect 3310 1261 3316 1262
rect 3310 1257 3311 1261
rect 3315 1257 3316 1261
rect 3310 1256 3316 1257
rect 3478 1261 3484 1262
rect 3478 1257 3479 1261
rect 3483 1257 3484 1261
rect 3478 1256 3484 1257
rect 1726 1252 1732 1253
rect 2495 1255 2501 1256
rect 2495 1251 2496 1255
rect 2500 1254 2501 1255
rect 2506 1255 2512 1256
rect 2506 1254 2507 1255
rect 2500 1252 2507 1254
rect 2500 1251 2501 1252
rect 2495 1250 2501 1251
rect 2506 1251 2507 1252
rect 2511 1251 2512 1255
rect 2506 1250 2512 1251
rect 3346 1255 3352 1256
rect 3346 1251 3347 1255
rect 3351 1254 3352 1255
rect 3359 1255 3365 1256
rect 3359 1254 3360 1255
rect 3351 1252 3360 1254
rect 3351 1251 3352 1252
rect 3346 1250 3352 1251
rect 3359 1251 3360 1252
rect 3364 1251 3365 1255
rect 3359 1250 3365 1251
rect 3498 1255 3504 1256
rect 3498 1251 3499 1255
rect 3503 1254 3504 1255
rect 3527 1255 3533 1256
rect 3527 1254 3528 1255
rect 3503 1252 3528 1254
rect 3503 1251 3504 1252
rect 3498 1250 3504 1251
rect 3527 1251 3528 1252
rect 3532 1251 3533 1255
rect 3527 1250 3533 1251
rect 542 1235 548 1236
rect 542 1231 543 1235
rect 547 1231 548 1235
rect 542 1230 548 1231
rect 630 1235 636 1236
rect 630 1231 631 1235
rect 635 1231 636 1235
rect 630 1230 636 1231
rect 718 1235 724 1236
rect 718 1231 719 1235
rect 723 1231 724 1235
rect 718 1230 724 1231
rect 806 1235 812 1236
rect 806 1231 807 1235
rect 811 1231 812 1235
rect 806 1230 812 1231
rect 894 1235 900 1236
rect 894 1231 895 1235
rect 899 1231 900 1235
rect 894 1230 900 1231
rect 990 1235 996 1236
rect 990 1231 991 1235
rect 995 1231 996 1235
rect 990 1230 996 1231
rect 1094 1235 1100 1236
rect 1094 1231 1095 1235
rect 1099 1231 1100 1235
rect 1094 1230 1100 1231
rect 1206 1235 1212 1236
rect 1206 1231 1207 1235
rect 1211 1231 1212 1235
rect 1206 1230 1212 1231
rect 1334 1235 1340 1236
rect 1334 1231 1335 1235
rect 1339 1231 1340 1235
rect 1334 1230 1340 1231
rect 1470 1235 1476 1236
rect 1470 1231 1471 1235
rect 1475 1231 1476 1235
rect 1470 1230 1476 1231
rect 1606 1235 1612 1236
rect 1606 1231 1607 1235
rect 1611 1231 1612 1235
rect 1606 1230 1612 1231
rect 1726 1235 1732 1236
rect 1726 1231 1727 1235
rect 1731 1231 1732 1235
rect 1726 1230 1732 1231
rect 2142 1231 2148 1232
rect 698 1227 704 1228
rect 110 1225 116 1226
rect 110 1221 111 1225
rect 115 1221 116 1225
rect 698 1223 699 1227
rect 703 1226 704 1227
rect 874 1227 880 1228
rect 703 1224 737 1226
rect 703 1223 704 1224
rect 698 1222 704 1223
rect 874 1223 875 1227
rect 879 1226 880 1227
rect 1542 1227 1548 1228
rect 1542 1226 1543 1227
rect 879 1224 913 1226
rect 1529 1224 1543 1226
rect 879 1223 880 1224
rect 874 1222 880 1223
rect 1542 1223 1543 1224
rect 1547 1223 1548 1227
rect 2142 1227 2143 1231
rect 2147 1227 2148 1231
rect 2142 1226 2148 1227
rect 2318 1231 2324 1232
rect 2318 1227 2319 1231
rect 2323 1227 2324 1231
rect 2318 1226 2324 1227
rect 2486 1231 2492 1232
rect 2486 1227 2487 1231
rect 2491 1227 2492 1231
rect 2486 1226 2492 1227
rect 2654 1231 2660 1232
rect 2654 1227 2655 1231
rect 2659 1227 2660 1231
rect 2654 1226 2660 1227
rect 2822 1231 2828 1232
rect 2822 1227 2823 1231
rect 2827 1227 2828 1231
rect 2822 1226 2828 1227
rect 2990 1231 2996 1232
rect 2990 1227 2991 1231
rect 2995 1227 2996 1231
rect 2990 1226 2996 1227
rect 3158 1231 3164 1232
rect 3158 1227 3159 1231
rect 3163 1227 3164 1231
rect 3158 1226 3164 1227
rect 3326 1231 3332 1232
rect 3326 1227 3327 1231
rect 3331 1227 3332 1231
rect 3326 1226 3332 1227
rect 3478 1231 3484 1232
rect 3478 1227 3479 1231
rect 3483 1227 3484 1231
rect 3478 1226 3484 1227
rect 1542 1222 1548 1223
rect 1822 1225 1828 1226
rect 110 1220 116 1221
rect 1822 1221 1823 1225
rect 1827 1221 1828 1225
rect 2230 1223 2236 1224
rect 2230 1222 2231 1223
rect 1822 1220 1828 1221
rect 1862 1221 1868 1222
rect 1862 1217 1863 1221
rect 1867 1217 1868 1221
rect 2201 1220 2231 1222
rect 2230 1219 2231 1220
rect 2235 1219 2236 1223
rect 2230 1218 2236 1219
rect 2814 1223 2820 1224
rect 2814 1219 2815 1223
rect 2819 1222 2820 1223
rect 3058 1223 3064 1224
rect 2819 1220 2841 1222
rect 2819 1219 2820 1220
rect 2814 1218 2820 1219
rect 3058 1219 3059 1223
rect 3063 1222 3064 1223
rect 3063 1220 3177 1222
rect 3574 1221 3580 1222
rect 3063 1219 3064 1220
rect 3058 1218 3064 1219
rect 1862 1216 1868 1217
rect 3574 1217 3575 1221
rect 3579 1217 3580 1221
rect 3574 1216 3580 1217
rect 623 1211 629 1212
rect 623 1210 624 1211
rect 110 1208 116 1209
rect 605 1208 624 1210
rect 110 1204 111 1208
rect 115 1204 116 1208
rect 623 1207 624 1208
rect 628 1207 629 1211
rect 711 1211 717 1212
rect 711 1210 712 1211
rect 693 1208 712 1210
rect 623 1206 629 1207
rect 711 1207 712 1208
rect 716 1207 717 1211
rect 887 1211 893 1212
rect 887 1210 888 1211
rect 869 1208 888 1210
rect 711 1206 717 1207
rect 887 1207 888 1208
rect 892 1207 893 1211
rect 1087 1211 1093 1212
rect 1087 1210 1088 1211
rect 1053 1208 1088 1210
rect 887 1206 893 1207
rect 1087 1207 1088 1208
rect 1092 1207 1093 1211
rect 1199 1211 1205 1212
rect 1199 1210 1200 1211
rect 1157 1208 1200 1210
rect 1087 1206 1093 1207
rect 1199 1207 1200 1208
rect 1204 1207 1205 1211
rect 1327 1211 1333 1212
rect 1327 1210 1328 1211
rect 1269 1208 1328 1210
rect 1199 1206 1205 1207
rect 1327 1207 1328 1208
rect 1332 1207 1333 1211
rect 1463 1211 1469 1212
rect 1463 1210 1464 1211
rect 1397 1208 1464 1210
rect 1327 1206 1333 1207
rect 1463 1207 1464 1208
rect 1468 1207 1469 1211
rect 1719 1211 1725 1212
rect 1719 1210 1720 1211
rect 1669 1208 1720 1210
rect 1463 1206 1469 1207
rect 1719 1207 1720 1208
rect 1724 1207 1725 1211
rect 1814 1211 1820 1212
rect 1814 1210 1815 1211
rect 1789 1208 1815 1210
rect 1719 1206 1725 1207
rect 1814 1207 1815 1208
rect 1819 1207 1820 1211
rect 1814 1206 1820 1207
rect 1822 1208 1828 1209
rect 110 1203 116 1204
rect 1822 1204 1823 1208
rect 1827 1204 1828 1208
rect 2210 1207 2216 1208
rect 1822 1203 1828 1204
rect 1862 1204 1868 1205
rect 1862 1200 1863 1204
rect 1867 1200 1868 1204
rect 2210 1203 2211 1207
rect 2215 1206 2216 1207
rect 2471 1207 2477 1208
rect 2215 1204 2345 1206
rect 2215 1203 2216 1204
rect 2210 1202 2216 1203
rect 2471 1203 2472 1207
rect 2476 1206 2477 1207
rect 2798 1207 2804 1208
rect 2798 1206 2799 1207
rect 2476 1204 2513 1206
rect 2717 1204 2799 1206
rect 2476 1203 2477 1204
rect 2471 1202 2477 1203
rect 2798 1203 2799 1204
rect 2803 1203 2804 1207
rect 3150 1207 3156 1208
rect 3150 1206 3151 1207
rect 3053 1204 3151 1206
rect 2798 1202 2804 1203
rect 3150 1203 3151 1204
rect 3155 1203 3156 1207
rect 3150 1202 3156 1203
rect 3226 1207 3232 1208
rect 3226 1203 3227 1207
rect 3231 1206 3232 1207
rect 3471 1207 3477 1208
rect 3231 1204 3353 1206
rect 3231 1203 3232 1204
rect 3226 1202 3232 1203
rect 3471 1203 3472 1207
rect 3476 1206 3477 1207
rect 3476 1204 3505 1206
rect 3574 1204 3580 1205
rect 3476 1203 3477 1204
rect 3471 1202 3477 1203
rect 1862 1199 1868 1200
rect 3574 1200 3575 1204
rect 3579 1200 3580 1204
rect 3574 1199 3580 1200
rect 550 1195 556 1196
rect 550 1191 551 1195
rect 555 1191 556 1195
rect 550 1190 556 1191
rect 638 1195 644 1196
rect 638 1191 639 1195
rect 643 1191 644 1195
rect 638 1190 644 1191
rect 726 1195 732 1196
rect 726 1191 727 1195
rect 731 1191 732 1195
rect 726 1190 732 1191
rect 814 1195 820 1196
rect 814 1191 815 1195
rect 819 1191 820 1195
rect 814 1190 820 1191
rect 902 1195 908 1196
rect 902 1191 903 1195
rect 907 1191 908 1195
rect 902 1190 908 1191
rect 998 1195 1004 1196
rect 998 1191 999 1195
rect 1003 1191 1004 1195
rect 998 1190 1004 1191
rect 1102 1195 1108 1196
rect 1102 1191 1103 1195
rect 1107 1191 1108 1195
rect 1102 1190 1108 1191
rect 1214 1195 1220 1196
rect 1214 1191 1215 1195
rect 1219 1191 1220 1195
rect 1214 1190 1220 1191
rect 1342 1195 1348 1196
rect 1342 1191 1343 1195
rect 1347 1191 1348 1195
rect 1342 1190 1348 1191
rect 1478 1195 1484 1196
rect 1478 1191 1479 1195
rect 1483 1191 1484 1195
rect 1478 1190 1484 1191
rect 1614 1195 1620 1196
rect 1614 1191 1615 1195
rect 1619 1191 1620 1195
rect 1614 1190 1620 1191
rect 1734 1195 1740 1196
rect 1734 1191 1735 1195
rect 1739 1191 1740 1195
rect 1734 1190 1740 1191
rect 2150 1191 2156 1192
rect 826 1187 832 1188
rect 826 1186 827 1187
rect 823 1185 827 1186
rect 559 1183 565 1184
rect 559 1179 560 1183
rect 564 1182 565 1183
rect 623 1183 629 1184
rect 564 1180 618 1182
rect 564 1179 565 1180
rect 559 1178 565 1179
rect 616 1174 618 1180
rect 623 1179 624 1183
rect 628 1182 629 1183
rect 647 1183 653 1184
rect 647 1182 648 1183
rect 628 1180 648 1182
rect 628 1179 629 1180
rect 623 1178 629 1179
rect 647 1179 648 1180
rect 652 1179 653 1183
rect 647 1178 653 1179
rect 735 1183 741 1184
rect 735 1179 736 1183
rect 740 1182 741 1183
rect 740 1180 818 1182
rect 823 1181 824 1185
rect 831 1183 832 1187
rect 2150 1187 2151 1191
rect 2155 1187 2156 1191
rect 2150 1186 2156 1187
rect 2326 1191 2332 1192
rect 2326 1187 2327 1191
rect 2331 1187 2332 1191
rect 2326 1186 2332 1187
rect 2494 1191 2500 1192
rect 2494 1187 2495 1191
rect 2499 1187 2500 1191
rect 2494 1186 2500 1187
rect 2662 1191 2668 1192
rect 2662 1187 2663 1191
rect 2667 1187 2668 1191
rect 2662 1186 2668 1187
rect 2830 1191 2836 1192
rect 2830 1187 2831 1191
rect 2835 1187 2836 1191
rect 2830 1186 2836 1187
rect 2998 1191 3004 1192
rect 2998 1187 2999 1191
rect 3003 1187 3004 1191
rect 2998 1186 3004 1187
rect 3166 1191 3172 1192
rect 3166 1187 3167 1191
rect 3171 1187 3172 1191
rect 3166 1186 3172 1187
rect 3334 1191 3340 1192
rect 3334 1187 3335 1191
rect 3339 1187 3340 1191
rect 3334 1186 3340 1187
rect 3486 1191 3492 1192
rect 3486 1187 3487 1191
rect 3491 1187 3492 1191
rect 3486 1186 3492 1187
rect 828 1182 832 1183
rect 887 1183 893 1184
rect 828 1181 829 1182
rect 823 1180 829 1181
rect 740 1179 741 1180
rect 735 1178 741 1179
rect 698 1175 704 1176
rect 698 1174 699 1175
rect 616 1172 699 1174
rect 698 1171 699 1172
rect 703 1171 704 1175
rect 816 1174 818 1180
rect 887 1179 888 1183
rect 892 1182 893 1183
rect 911 1183 917 1184
rect 911 1182 912 1183
rect 892 1180 912 1182
rect 892 1179 893 1180
rect 887 1178 893 1179
rect 911 1179 912 1180
rect 916 1179 917 1183
rect 911 1178 917 1179
rect 1007 1183 1016 1184
rect 1007 1179 1008 1183
rect 1015 1179 1016 1183
rect 1007 1178 1016 1179
rect 1087 1183 1093 1184
rect 1087 1179 1088 1183
rect 1092 1182 1093 1183
rect 1111 1183 1117 1184
rect 1111 1182 1112 1183
rect 1092 1180 1112 1182
rect 1092 1179 1093 1180
rect 1087 1178 1093 1179
rect 1111 1179 1112 1180
rect 1116 1179 1117 1183
rect 1111 1178 1117 1179
rect 1199 1183 1205 1184
rect 1199 1179 1200 1183
rect 1204 1182 1205 1183
rect 1223 1183 1229 1184
rect 1223 1182 1224 1183
rect 1204 1180 1224 1182
rect 1204 1179 1205 1180
rect 1199 1178 1205 1179
rect 1223 1179 1224 1180
rect 1228 1179 1229 1183
rect 1223 1178 1229 1179
rect 1327 1183 1333 1184
rect 1327 1179 1328 1183
rect 1332 1182 1333 1183
rect 1351 1183 1357 1184
rect 1351 1182 1352 1183
rect 1332 1180 1352 1182
rect 1332 1179 1333 1180
rect 1327 1178 1333 1179
rect 1351 1179 1352 1180
rect 1356 1179 1357 1183
rect 1351 1178 1357 1179
rect 1463 1183 1469 1184
rect 1463 1179 1464 1183
rect 1468 1182 1469 1183
rect 1487 1183 1493 1184
rect 1487 1182 1488 1183
rect 1468 1180 1488 1182
rect 1468 1179 1469 1180
rect 1463 1178 1469 1179
rect 1487 1179 1488 1180
rect 1492 1179 1493 1183
rect 1487 1178 1493 1179
rect 1623 1183 1632 1184
rect 1623 1179 1624 1183
rect 1631 1179 1632 1183
rect 1623 1178 1632 1179
rect 1719 1183 1725 1184
rect 1719 1179 1720 1183
rect 1724 1182 1725 1183
rect 1743 1183 1749 1184
rect 1743 1182 1744 1183
rect 1724 1180 1744 1182
rect 1724 1179 1725 1180
rect 1719 1178 1725 1179
rect 1743 1179 1744 1180
rect 1748 1179 1749 1183
rect 1743 1178 1749 1179
rect 2159 1179 2165 1180
rect 874 1175 880 1176
rect 874 1174 875 1175
rect 816 1172 875 1174
rect 698 1170 704 1171
rect 874 1171 875 1172
rect 879 1171 880 1175
rect 2159 1175 2160 1179
rect 2164 1178 2165 1179
rect 2210 1179 2216 1180
rect 2210 1178 2211 1179
rect 2164 1176 2211 1178
rect 2164 1175 2165 1176
rect 2159 1174 2165 1175
rect 2210 1175 2211 1176
rect 2215 1175 2216 1179
rect 2210 1174 2216 1175
rect 2335 1179 2341 1180
rect 2335 1175 2336 1179
rect 2340 1178 2341 1179
rect 2354 1179 2360 1180
rect 2354 1178 2355 1179
rect 2340 1176 2355 1178
rect 2340 1175 2341 1176
rect 2335 1174 2341 1175
rect 2354 1175 2355 1176
rect 2359 1175 2360 1179
rect 2354 1174 2360 1175
rect 2503 1179 2512 1180
rect 2503 1175 2504 1179
rect 2511 1175 2512 1179
rect 2503 1174 2512 1175
rect 2671 1179 2677 1180
rect 2671 1175 2672 1179
rect 2676 1178 2677 1179
rect 2682 1179 2688 1180
rect 2682 1178 2683 1179
rect 2676 1176 2683 1178
rect 2676 1175 2677 1176
rect 2671 1174 2677 1175
rect 2682 1175 2683 1176
rect 2687 1175 2688 1179
rect 2682 1174 2688 1175
rect 2798 1179 2804 1180
rect 2798 1175 2799 1179
rect 2803 1178 2804 1179
rect 2839 1179 2845 1180
rect 2839 1178 2840 1179
rect 2803 1176 2840 1178
rect 2803 1175 2804 1176
rect 2798 1174 2804 1175
rect 2839 1175 2840 1176
rect 2844 1175 2845 1179
rect 2839 1174 2845 1175
rect 3007 1179 3013 1180
rect 3007 1175 3008 1179
rect 3012 1178 3013 1179
rect 3058 1179 3064 1180
rect 3058 1178 3059 1179
rect 3012 1176 3059 1178
rect 3012 1175 3013 1176
rect 3007 1174 3013 1175
rect 3058 1175 3059 1176
rect 3063 1175 3064 1179
rect 3058 1174 3064 1175
rect 3175 1179 3181 1180
rect 3175 1175 3176 1179
rect 3180 1178 3181 1179
rect 3226 1179 3232 1180
rect 3226 1178 3227 1179
rect 3180 1176 3227 1178
rect 3180 1175 3181 1176
rect 3175 1174 3181 1175
rect 3226 1175 3227 1176
rect 3231 1175 3232 1179
rect 3226 1174 3232 1175
rect 3343 1179 3352 1180
rect 3343 1175 3344 1179
rect 3351 1175 3352 1179
rect 3343 1174 3352 1175
rect 3495 1179 3504 1180
rect 3495 1175 3496 1179
rect 3503 1175 3504 1179
rect 3495 1174 3504 1175
rect 874 1170 880 1171
rect 1375 1171 1381 1172
rect 1375 1170 1376 1171
rect 1193 1168 1376 1170
rect 1193 1164 1195 1168
rect 1375 1167 1376 1168
rect 1380 1167 1381 1171
rect 1375 1166 1381 1167
rect 1814 1167 1820 1168
rect 367 1163 373 1164
rect 367 1159 368 1163
rect 372 1162 373 1163
rect 414 1163 420 1164
rect 414 1162 415 1163
rect 372 1160 415 1162
rect 372 1159 373 1160
rect 367 1158 373 1159
rect 414 1159 415 1160
rect 419 1159 420 1163
rect 414 1158 420 1159
rect 423 1163 429 1164
rect 423 1159 424 1163
rect 428 1162 429 1163
rect 479 1163 485 1164
rect 479 1162 480 1163
rect 428 1160 480 1162
rect 428 1159 429 1160
rect 423 1158 429 1159
rect 479 1159 480 1160
rect 484 1159 485 1163
rect 479 1158 485 1159
rect 535 1163 541 1164
rect 535 1159 536 1163
rect 540 1162 541 1163
rect 599 1163 605 1164
rect 599 1162 600 1163
rect 540 1160 600 1162
rect 540 1159 541 1160
rect 535 1158 541 1159
rect 599 1159 600 1160
rect 604 1159 605 1163
rect 599 1158 605 1159
rect 711 1163 717 1164
rect 711 1159 712 1163
rect 716 1162 717 1163
rect 719 1163 725 1164
rect 719 1162 720 1163
rect 716 1160 720 1162
rect 716 1159 717 1160
rect 711 1158 717 1159
rect 719 1159 720 1160
rect 724 1159 725 1163
rect 719 1158 725 1159
rect 770 1163 776 1164
rect 770 1159 771 1163
rect 775 1162 776 1163
rect 839 1163 845 1164
rect 839 1162 840 1163
rect 775 1160 840 1162
rect 775 1159 776 1160
rect 770 1158 776 1159
rect 839 1159 840 1160
rect 844 1159 845 1163
rect 839 1158 845 1159
rect 959 1163 965 1164
rect 959 1159 960 1163
rect 964 1162 965 1163
rect 1018 1163 1024 1164
rect 1018 1162 1019 1163
rect 964 1160 1019 1162
rect 964 1159 965 1160
rect 959 1158 965 1159
rect 1018 1159 1019 1160
rect 1023 1159 1024 1163
rect 1018 1158 1024 1159
rect 1071 1163 1077 1164
rect 1071 1159 1072 1163
rect 1076 1162 1077 1163
rect 1134 1163 1140 1164
rect 1134 1162 1135 1163
rect 1076 1160 1135 1162
rect 1076 1159 1077 1160
rect 1071 1158 1077 1159
rect 1134 1159 1135 1160
rect 1139 1159 1140 1163
rect 1134 1158 1140 1159
rect 1191 1163 1197 1164
rect 1191 1159 1192 1163
rect 1196 1159 1197 1163
rect 1191 1158 1197 1159
rect 1311 1163 1317 1164
rect 1311 1159 1312 1163
rect 1316 1162 1317 1163
rect 1322 1163 1328 1164
rect 1322 1162 1323 1163
rect 1316 1160 1323 1162
rect 1316 1159 1317 1160
rect 1311 1158 1317 1159
rect 1322 1159 1323 1160
rect 1327 1159 1328 1163
rect 1322 1158 1328 1159
rect 1367 1163 1373 1164
rect 1367 1159 1368 1163
rect 1372 1162 1373 1163
rect 1431 1163 1437 1164
rect 1431 1162 1432 1163
rect 1372 1160 1432 1162
rect 1372 1159 1373 1160
rect 1367 1158 1373 1159
rect 1431 1159 1432 1160
rect 1436 1159 1437 1163
rect 1814 1163 1815 1167
rect 1819 1166 1820 1167
rect 1903 1167 1909 1168
rect 1903 1166 1904 1167
rect 1819 1164 1904 1166
rect 1819 1163 1820 1164
rect 1814 1162 1820 1163
rect 1903 1163 1904 1164
rect 1908 1163 1909 1167
rect 1903 1162 1909 1163
rect 1959 1167 1965 1168
rect 1959 1163 1960 1167
rect 1964 1166 1965 1167
rect 2015 1167 2021 1168
rect 2015 1166 2016 1167
rect 1964 1164 2016 1166
rect 1964 1163 1965 1164
rect 1959 1162 1965 1163
rect 2015 1163 2016 1164
rect 2020 1163 2021 1167
rect 2015 1162 2021 1163
rect 2079 1167 2085 1168
rect 2079 1163 2080 1167
rect 2084 1166 2085 1167
rect 2151 1167 2157 1168
rect 2151 1166 2152 1167
rect 2084 1164 2152 1166
rect 2084 1163 2085 1164
rect 2079 1162 2085 1163
rect 2151 1163 2152 1164
rect 2156 1163 2157 1167
rect 2151 1162 2157 1163
rect 2302 1167 2309 1168
rect 2302 1163 2303 1167
rect 2308 1163 2309 1167
rect 2302 1162 2309 1163
rect 2463 1167 2469 1168
rect 2463 1163 2464 1167
rect 2468 1166 2469 1167
rect 2471 1167 2477 1168
rect 2471 1166 2472 1167
rect 2468 1164 2472 1166
rect 2468 1163 2469 1164
rect 2463 1162 2469 1163
rect 2471 1163 2472 1164
rect 2476 1163 2477 1167
rect 2471 1162 2477 1163
rect 2631 1167 2640 1168
rect 2631 1163 2632 1167
rect 2639 1163 2640 1167
rect 2631 1162 2640 1163
rect 2799 1167 2808 1168
rect 2799 1163 2800 1167
rect 2807 1163 2808 1167
rect 2799 1162 2808 1163
rect 2887 1167 2893 1168
rect 2887 1163 2888 1167
rect 2892 1166 2893 1167
rect 2975 1167 2981 1168
rect 2975 1166 2976 1167
rect 2892 1164 2976 1166
rect 2892 1163 2893 1164
rect 2887 1162 2893 1163
rect 2975 1163 2976 1164
rect 2980 1163 2981 1167
rect 2975 1162 2981 1163
rect 3150 1167 3157 1168
rect 3150 1163 3151 1167
rect 3156 1163 3157 1167
rect 3150 1162 3157 1163
rect 3231 1167 3237 1168
rect 3231 1163 3232 1167
rect 3236 1166 3237 1167
rect 3335 1167 3341 1168
rect 3335 1166 3336 1167
rect 3236 1164 3336 1166
rect 3236 1163 3237 1164
rect 3231 1162 3237 1163
rect 3335 1163 3336 1164
rect 3340 1163 3341 1167
rect 3335 1162 3341 1163
rect 3471 1167 3477 1168
rect 3471 1163 3472 1167
rect 3476 1166 3477 1167
rect 3495 1167 3501 1168
rect 3495 1166 3496 1167
rect 3476 1164 3496 1166
rect 3476 1163 3477 1164
rect 3471 1162 3477 1163
rect 3495 1163 3496 1164
rect 3500 1163 3501 1167
rect 3495 1162 3501 1163
rect 1431 1158 1437 1159
rect 1894 1157 1900 1158
rect 358 1153 364 1154
rect 358 1149 359 1153
rect 363 1149 364 1153
rect 358 1148 364 1149
rect 470 1153 476 1154
rect 470 1149 471 1153
rect 475 1149 476 1153
rect 470 1148 476 1149
rect 590 1153 596 1154
rect 590 1149 591 1153
rect 595 1149 596 1153
rect 590 1148 596 1149
rect 710 1153 716 1154
rect 710 1149 711 1153
rect 715 1149 716 1153
rect 710 1148 716 1149
rect 830 1153 836 1154
rect 830 1149 831 1153
rect 835 1149 836 1153
rect 830 1148 836 1149
rect 950 1153 956 1154
rect 950 1149 951 1153
rect 955 1149 956 1153
rect 950 1148 956 1149
rect 1062 1153 1068 1154
rect 1062 1149 1063 1153
rect 1067 1149 1068 1153
rect 1062 1148 1068 1149
rect 1182 1153 1188 1154
rect 1182 1149 1183 1153
rect 1187 1149 1188 1153
rect 1182 1148 1188 1149
rect 1302 1153 1308 1154
rect 1302 1149 1303 1153
rect 1307 1149 1308 1153
rect 1302 1148 1308 1149
rect 1422 1153 1428 1154
rect 1422 1149 1423 1153
rect 1427 1149 1428 1153
rect 1894 1153 1895 1157
rect 1899 1153 1900 1157
rect 1894 1152 1900 1153
rect 2006 1157 2012 1158
rect 2006 1153 2007 1157
rect 2011 1153 2012 1157
rect 2006 1152 2012 1153
rect 2142 1157 2148 1158
rect 2142 1153 2143 1157
rect 2147 1153 2148 1157
rect 2142 1152 2148 1153
rect 2294 1157 2300 1158
rect 2294 1153 2295 1157
rect 2299 1153 2300 1157
rect 2294 1152 2300 1153
rect 2454 1157 2460 1158
rect 2454 1153 2455 1157
rect 2459 1153 2460 1157
rect 2454 1152 2460 1153
rect 2622 1157 2628 1158
rect 2622 1153 2623 1157
rect 2627 1153 2628 1157
rect 2622 1152 2628 1153
rect 2790 1157 2796 1158
rect 2790 1153 2791 1157
rect 2795 1153 2796 1157
rect 2790 1152 2796 1153
rect 2966 1157 2972 1158
rect 2966 1153 2967 1157
rect 2971 1153 2972 1157
rect 2966 1152 2972 1153
rect 3142 1157 3148 1158
rect 3142 1153 3143 1157
rect 3147 1153 3148 1157
rect 3142 1152 3148 1153
rect 3326 1157 3332 1158
rect 3326 1153 3327 1157
rect 3331 1153 3332 1157
rect 3326 1152 3332 1153
rect 3486 1157 3492 1158
rect 3486 1153 3487 1157
rect 3491 1153 3492 1157
rect 3486 1152 3492 1153
rect 1422 1148 1428 1149
rect 1862 1144 1868 1145
rect 3574 1144 3580 1145
rect 110 1140 116 1141
rect 1822 1140 1828 1141
rect 110 1136 111 1140
rect 115 1136 116 1140
rect 423 1139 429 1140
rect 423 1138 424 1139
rect 413 1136 424 1138
rect 110 1135 116 1136
rect 423 1135 424 1136
rect 428 1135 429 1139
rect 535 1139 541 1140
rect 535 1138 536 1139
rect 525 1136 536 1138
rect 423 1134 429 1135
rect 535 1135 536 1136
rect 540 1135 541 1139
rect 770 1139 776 1140
rect 770 1138 771 1139
rect 765 1136 771 1138
rect 535 1134 541 1135
rect 770 1135 771 1136
rect 775 1135 776 1139
rect 1010 1139 1016 1140
rect 1010 1138 1011 1139
rect 1005 1136 1011 1138
rect 770 1134 776 1135
rect 778 1135 784 1136
rect 778 1131 779 1135
rect 783 1134 784 1135
rect 1010 1135 1011 1136
rect 1015 1135 1016 1139
rect 1367 1139 1373 1140
rect 1367 1138 1368 1139
rect 1357 1136 1368 1138
rect 1010 1134 1016 1135
rect 1018 1135 1024 1136
rect 783 1132 849 1134
rect 783 1131 784 1132
rect 778 1130 784 1131
rect 1018 1131 1019 1135
rect 1023 1134 1024 1135
rect 1134 1135 1140 1136
rect 1023 1132 1081 1134
rect 1023 1131 1024 1132
rect 1018 1130 1024 1131
rect 1134 1131 1135 1135
rect 1139 1134 1140 1135
rect 1367 1135 1368 1136
rect 1372 1135 1373 1139
rect 1822 1136 1823 1140
rect 1827 1136 1828 1140
rect 1862 1140 1863 1144
rect 1867 1140 1868 1144
rect 1959 1143 1965 1144
rect 1959 1142 1960 1143
rect 1949 1140 1960 1142
rect 1862 1139 1868 1140
rect 1959 1139 1960 1140
rect 1964 1139 1965 1143
rect 2079 1143 2085 1144
rect 2079 1142 2080 1143
rect 2061 1140 2080 1142
rect 1959 1138 1965 1139
rect 2079 1139 2080 1140
rect 2084 1139 2085 1143
rect 2354 1143 2360 1144
rect 2354 1142 2355 1143
rect 2349 1140 2355 1142
rect 2079 1138 2085 1139
rect 2354 1139 2355 1140
rect 2359 1139 2360 1143
rect 2682 1143 2688 1144
rect 2682 1142 2683 1143
rect 2677 1140 2683 1142
rect 2354 1138 2360 1139
rect 2682 1139 2683 1140
rect 2687 1139 2688 1143
rect 2887 1143 2893 1144
rect 2887 1142 2888 1143
rect 2845 1140 2888 1142
rect 2682 1138 2688 1139
rect 2887 1139 2888 1140
rect 2892 1139 2893 1143
rect 3231 1143 3237 1144
rect 3231 1142 3232 1143
rect 3197 1140 3232 1142
rect 2887 1138 2893 1139
rect 3231 1139 3232 1140
rect 3236 1139 3237 1143
rect 3574 1140 3575 1144
rect 3579 1140 3580 1144
rect 3574 1139 3580 1140
rect 3231 1138 3237 1139
rect 1367 1134 1373 1135
rect 1375 1135 1381 1136
rect 1822 1135 1828 1136
rect 1139 1132 1201 1134
rect 1139 1131 1140 1132
rect 1134 1130 1140 1131
rect 1375 1131 1376 1135
rect 1380 1134 1381 1135
rect 1380 1132 1441 1134
rect 1380 1131 1381 1132
rect 1375 1130 1381 1131
rect 1862 1127 1868 1128
rect 110 1123 116 1124
rect 110 1119 111 1123
rect 115 1119 116 1123
rect 110 1118 116 1119
rect 1822 1123 1828 1124
rect 1822 1119 1823 1123
rect 1827 1119 1828 1123
rect 1862 1123 1863 1127
rect 1867 1123 1868 1127
rect 1862 1122 1868 1123
rect 2074 1127 2080 1128
rect 2074 1123 2075 1127
rect 2079 1126 2080 1127
rect 2582 1127 2588 1128
rect 2582 1126 2583 1127
rect 2079 1124 2153 1126
rect 2505 1124 2583 1126
rect 2079 1123 2080 1124
rect 2074 1122 2080 1123
rect 2582 1123 2583 1124
rect 2587 1123 2588 1127
rect 3574 1127 3580 1128
rect 2582 1122 2588 1123
rect 2908 1124 2977 1126
rect 1822 1118 1828 1119
rect 1886 1117 1892 1118
rect 350 1113 356 1114
rect 350 1109 351 1113
rect 355 1109 356 1113
rect 350 1108 356 1109
rect 462 1113 468 1114
rect 462 1109 463 1113
rect 467 1109 468 1113
rect 462 1108 468 1109
rect 582 1113 588 1114
rect 582 1109 583 1113
rect 587 1109 588 1113
rect 582 1108 588 1109
rect 702 1113 708 1114
rect 702 1109 703 1113
rect 707 1109 708 1113
rect 702 1108 708 1109
rect 822 1113 828 1114
rect 822 1109 823 1113
rect 827 1109 828 1113
rect 822 1108 828 1109
rect 942 1113 948 1114
rect 942 1109 943 1113
rect 947 1109 948 1113
rect 942 1108 948 1109
rect 1054 1113 1060 1114
rect 1054 1109 1055 1113
rect 1059 1109 1060 1113
rect 1054 1108 1060 1109
rect 1174 1113 1180 1114
rect 1174 1109 1175 1113
rect 1179 1109 1180 1113
rect 1174 1108 1180 1109
rect 1294 1113 1300 1114
rect 1294 1109 1295 1113
rect 1299 1109 1300 1113
rect 1294 1108 1300 1109
rect 1414 1113 1420 1114
rect 1414 1109 1415 1113
rect 1419 1109 1420 1113
rect 1886 1113 1887 1117
rect 1891 1113 1892 1117
rect 1886 1112 1892 1113
rect 1998 1117 2004 1118
rect 1998 1113 1999 1117
rect 2003 1113 2004 1117
rect 1998 1112 2004 1113
rect 2134 1117 2140 1118
rect 2134 1113 2135 1117
rect 2139 1113 2140 1117
rect 2134 1112 2140 1113
rect 2286 1117 2292 1118
rect 2286 1113 2287 1117
rect 2291 1113 2292 1117
rect 2286 1112 2292 1113
rect 2446 1117 2452 1118
rect 2446 1113 2447 1117
rect 2451 1113 2452 1117
rect 2446 1112 2452 1113
rect 2614 1117 2620 1118
rect 2614 1113 2615 1117
rect 2619 1113 2620 1117
rect 2614 1112 2620 1113
rect 2782 1117 2788 1118
rect 2782 1113 2783 1117
rect 2787 1113 2788 1117
rect 2782 1112 2788 1113
rect 1414 1108 1420 1109
rect 2634 1111 2640 1112
rect 630 1107 637 1108
rect 630 1103 631 1107
rect 636 1103 637 1107
rect 2634 1107 2635 1111
rect 2639 1110 2640 1111
rect 2908 1110 2910 1124
rect 3574 1123 3575 1127
rect 3579 1123 3580 1127
rect 3574 1122 3580 1123
rect 2958 1117 2964 1118
rect 2958 1113 2959 1117
rect 2963 1113 2964 1117
rect 2958 1112 2964 1113
rect 3134 1117 3140 1118
rect 3134 1113 3135 1117
rect 3139 1113 3140 1117
rect 3134 1112 3140 1113
rect 3318 1117 3324 1118
rect 3318 1113 3319 1117
rect 3323 1113 3324 1117
rect 3318 1112 3324 1113
rect 3478 1117 3484 1118
rect 3478 1113 3479 1117
rect 3483 1113 3484 1117
rect 3478 1112 3484 1113
rect 2639 1108 2910 1110
rect 3366 1111 3373 1112
rect 2639 1107 2640 1108
rect 2634 1106 2640 1107
rect 3366 1107 3367 1111
rect 3372 1107 3373 1111
rect 3366 1106 3373 1107
rect 3498 1111 3504 1112
rect 3498 1107 3499 1111
rect 3503 1110 3504 1111
rect 3527 1111 3533 1112
rect 3527 1110 3528 1111
rect 3503 1108 3528 1110
rect 3503 1107 3504 1108
rect 3498 1106 3504 1107
rect 3527 1107 3528 1108
rect 3532 1107 3533 1111
rect 3527 1106 3533 1107
rect 630 1102 637 1103
rect 142 1087 148 1088
rect 142 1083 143 1087
rect 147 1083 148 1087
rect 142 1082 148 1083
rect 286 1087 292 1088
rect 286 1083 287 1087
rect 291 1083 292 1087
rect 286 1082 292 1083
rect 446 1087 452 1088
rect 446 1083 447 1087
rect 451 1083 452 1087
rect 446 1082 452 1083
rect 614 1087 620 1088
rect 614 1083 615 1087
rect 619 1083 620 1087
rect 614 1082 620 1083
rect 782 1087 788 1088
rect 782 1083 783 1087
rect 787 1083 788 1087
rect 782 1082 788 1083
rect 942 1087 948 1088
rect 942 1083 943 1087
rect 947 1083 948 1087
rect 942 1082 948 1083
rect 1102 1087 1108 1088
rect 1102 1083 1103 1087
rect 1107 1083 1108 1087
rect 1102 1082 1108 1083
rect 1254 1087 1260 1088
rect 1254 1083 1255 1087
rect 1259 1083 1260 1087
rect 1254 1082 1260 1083
rect 1406 1087 1412 1088
rect 1406 1083 1407 1087
rect 1411 1083 1412 1087
rect 1406 1082 1412 1083
rect 1558 1087 1564 1088
rect 1558 1083 1559 1087
rect 1563 1083 1564 1087
rect 1558 1082 1564 1083
rect 1894 1087 1900 1088
rect 1894 1083 1895 1087
rect 1899 1083 1900 1087
rect 1894 1082 1900 1083
rect 2046 1087 2052 1088
rect 2046 1083 2047 1087
rect 2051 1083 2052 1087
rect 2046 1082 2052 1083
rect 2214 1087 2220 1088
rect 2214 1083 2215 1087
rect 2219 1083 2220 1087
rect 2214 1082 2220 1083
rect 2390 1087 2396 1088
rect 2390 1083 2391 1087
rect 2395 1083 2396 1087
rect 2390 1082 2396 1083
rect 2566 1087 2572 1088
rect 2566 1083 2567 1087
rect 2571 1083 2572 1087
rect 2566 1082 2572 1083
rect 2734 1087 2740 1088
rect 2734 1083 2735 1087
rect 2739 1083 2740 1087
rect 2734 1082 2740 1083
rect 2894 1087 2900 1088
rect 2894 1083 2895 1087
rect 2899 1083 2900 1087
rect 2894 1082 2900 1083
rect 3046 1087 3052 1088
rect 3046 1083 3047 1087
rect 3051 1083 3052 1087
rect 3046 1082 3052 1083
rect 3198 1087 3204 1088
rect 3198 1083 3199 1087
rect 3203 1083 3204 1087
rect 3198 1082 3204 1083
rect 3350 1087 3356 1088
rect 3350 1083 3351 1087
rect 3355 1083 3356 1087
rect 3350 1082 3356 1083
rect 3478 1087 3484 1088
rect 3478 1083 3479 1087
rect 3483 1083 3484 1087
rect 3478 1082 3484 1083
rect 682 1079 688 1080
rect 110 1077 116 1078
rect 110 1073 111 1077
rect 115 1073 116 1077
rect 682 1075 683 1079
rect 687 1078 688 1079
rect 1322 1079 1328 1080
rect 1322 1078 1323 1079
rect 687 1076 801 1078
rect 1313 1076 1323 1078
rect 687 1075 688 1076
rect 682 1074 688 1075
rect 1322 1075 1323 1076
rect 1327 1075 1328 1079
rect 1322 1074 1328 1075
rect 1474 1079 1480 1080
rect 1474 1075 1475 1079
rect 1479 1078 1480 1079
rect 2302 1079 2308 1080
rect 2302 1078 2303 1079
rect 1479 1076 1577 1078
rect 1822 1077 1828 1078
rect 1479 1075 1480 1076
rect 1474 1074 1480 1075
rect 110 1072 116 1073
rect 1822 1073 1823 1077
rect 1827 1073 1828 1077
rect 1822 1072 1828 1073
rect 1862 1077 1868 1078
rect 1862 1073 1863 1077
rect 1867 1073 1868 1077
rect 2273 1076 2303 1078
rect 2302 1075 2303 1076
rect 2307 1075 2308 1079
rect 2802 1079 2808 1080
rect 2802 1078 2803 1079
rect 2793 1076 2803 1078
rect 2302 1074 2308 1075
rect 2802 1075 2803 1076
rect 2807 1075 2808 1079
rect 2802 1074 2808 1075
rect 3418 1079 3424 1080
rect 3418 1075 3419 1079
rect 3423 1078 3424 1079
rect 3423 1076 3497 1078
rect 3574 1077 3580 1078
rect 3423 1075 3424 1076
rect 3418 1074 3424 1075
rect 1862 1072 1868 1073
rect 3574 1073 3575 1077
rect 3579 1073 3580 1077
rect 3574 1072 3580 1073
rect 279 1063 285 1064
rect 279 1062 280 1063
rect 110 1060 116 1061
rect 205 1060 280 1062
rect 110 1056 111 1060
rect 115 1056 116 1060
rect 279 1059 280 1060
rect 284 1059 285 1063
rect 439 1063 445 1064
rect 439 1062 440 1063
rect 349 1060 440 1062
rect 279 1058 285 1059
rect 439 1059 440 1060
rect 444 1059 445 1063
rect 514 1063 520 1064
rect 514 1062 515 1063
rect 509 1060 515 1062
rect 439 1058 445 1059
rect 514 1059 515 1060
rect 519 1059 520 1063
rect 775 1063 781 1064
rect 775 1062 776 1063
rect 677 1060 776 1062
rect 514 1058 520 1059
rect 775 1059 776 1060
rect 780 1059 781 1063
rect 1095 1063 1101 1064
rect 1095 1062 1096 1063
rect 1005 1060 1096 1062
rect 775 1058 781 1059
rect 1095 1059 1096 1060
rect 1100 1059 1101 1063
rect 1242 1063 1248 1064
rect 1242 1062 1243 1063
rect 1165 1060 1243 1062
rect 1095 1058 1101 1059
rect 1242 1059 1243 1060
rect 1247 1059 1248 1063
rect 1551 1063 1557 1064
rect 1551 1062 1552 1063
rect 1469 1060 1552 1062
rect 1242 1058 1248 1059
rect 1551 1059 1552 1060
rect 1556 1059 1557 1063
rect 1982 1063 1988 1064
rect 1982 1062 1983 1063
rect 1551 1058 1557 1059
rect 1822 1060 1828 1061
rect 110 1055 116 1056
rect 1822 1056 1823 1060
rect 1827 1056 1828 1060
rect 1822 1055 1828 1056
rect 1862 1060 1868 1061
rect 1957 1060 1983 1062
rect 1862 1056 1863 1060
rect 1867 1056 1868 1060
rect 1982 1059 1983 1060
rect 1987 1059 1988 1063
rect 1982 1058 1988 1059
rect 1990 1063 1996 1064
rect 1990 1059 1991 1063
rect 1995 1062 1996 1063
rect 2282 1063 2288 1064
rect 1995 1060 2073 1062
rect 1995 1059 1996 1060
rect 1990 1058 1996 1059
rect 2282 1059 2283 1063
rect 2287 1062 2288 1063
rect 2506 1063 2512 1064
rect 2287 1060 2417 1062
rect 2287 1059 2288 1060
rect 2282 1058 2288 1059
rect 2506 1059 2507 1063
rect 2511 1062 2512 1063
rect 2802 1063 2808 1064
rect 2511 1060 2593 1062
rect 2511 1059 2512 1060
rect 2506 1058 2512 1059
rect 2802 1059 2803 1063
rect 2807 1062 2808 1063
rect 2962 1063 2968 1064
rect 2807 1060 2921 1062
rect 2807 1059 2808 1060
rect 2802 1058 2808 1059
rect 2962 1059 2963 1063
rect 2967 1062 2968 1063
rect 3114 1063 3120 1064
rect 2967 1060 3073 1062
rect 2967 1059 2968 1060
rect 2962 1058 2968 1059
rect 3114 1059 3115 1063
rect 3119 1062 3120 1063
rect 3266 1063 3272 1064
rect 3119 1060 3225 1062
rect 3119 1059 3120 1060
rect 3114 1058 3120 1059
rect 3266 1059 3267 1063
rect 3271 1062 3272 1063
rect 3271 1060 3377 1062
rect 3574 1060 3580 1061
rect 3271 1059 3272 1060
rect 3266 1058 3272 1059
rect 1862 1055 1868 1056
rect 3574 1056 3575 1060
rect 3579 1056 3580 1060
rect 3574 1055 3580 1056
rect 150 1047 156 1048
rect 150 1043 151 1047
rect 155 1043 156 1047
rect 150 1042 156 1043
rect 294 1047 300 1048
rect 294 1043 295 1047
rect 299 1043 300 1047
rect 294 1042 300 1043
rect 454 1047 460 1048
rect 454 1043 455 1047
rect 459 1043 460 1047
rect 454 1042 460 1043
rect 622 1047 628 1048
rect 622 1043 623 1047
rect 627 1043 628 1047
rect 622 1042 628 1043
rect 790 1047 796 1048
rect 790 1043 791 1047
rect 795 1043 796 1047
rect 790 1042 796 1043
rect 950 1047 956 1048
rect 950 1043 951 1047
rect 955 1043 956 1047
rect 950 1042 956 1043
rect 1110 1047 1116 1048
rect 1110 1043 1111 1047
rect 1115 1043 1116 1047
rect 1110 1042 1116 1043
rect 1262 1047 1268 1048
rect 1262 1043 1263 1047
rect 1267 1043 1268 1047
rect 1262 1042 1268 1043
rect 1414 1047 1420 1048
rect 1414 1043 1415 1047
rect 1419 1043 1420 1047
rect 1414 1042 1420 1043
rect 1566 1047 1572 1048
rect 1566 1043 1567 1047
rect 1571 1043 1572 1047
rect 1566 1042 1572 1043
rect 1902 1047 1908 1048
rect 1902 1043 1903 1047
rect 1907 1043 1908 1047
rect 1902 1042 1908 1043
rect 2054 1047 2060 1048
rect 2054 1043 2055 1047
rect 2059 1043 2060 1047
rect 2054 1042 2060 1043
rect 2222 1047 2228 1048
rect 2222 1043 2223 1047
rect 2227 1043 2228 1047
rect 2222 1042 2228 1043
rect 2398 1047 2404 1048
rect 2398 1043 2399 1047
rect 2403 1043 2404 1047
rect 2398 1042 2404 1043
rect 2574 1047 2580 1048
rect 2574 1043 2575 1047
rect 2579 1043 2580 1047
rect 2574 1042 2580 1043
rect 2742 1047 2748 1048
rect 2742 1043 2743 1047
rect 2747 1043 2748 1047
rect 2742 1042 2748 1043
rect 2902 1047 2908 1048
rect 2902 1043 2903 1047
rect 2907 1043 2908 1047
rect 2902 1042 2908 1043
rect 3054 1047 3060 1048
rect 3054 1043 3055 1047
rect 3059 1043 3060 1047
rect 3054 1042 3060 1043
rect 3206 1047 3212 1048
rect 3206 1043 3207 1047
rect 3211 1043 3212 1047
rect 3206 1042 3212 1043
rect 3358 1047 3364 1048
rect 3358 1043 3359 1047
rect 3363 1043 3364 1047
rect 3358 1042 3364 1043
rect 3486 1047 3492 1048
rect 3486 1043 3487 1047
rect 3491 1043 3492 1047
rect 3486 1042 3492 1043
rect 159 1035 168 1036
rect 159 1031 160 1035
rect 167 1031 168 1035
rect 159 1030 168 1031
rect 279 1035 285 1036
rect 279 1031 280 1035
rect 284 1034 285 1035
rect 303 1035 309 1036
rect 303 1034 304 1035
rect 284 1032 304 1034
rect 284 1031 285 1032
rect 279 1030 285 1031
rect 303 1031 304 1032
rect 308 1031 309 1035
rect 303 1030 309 1031
rect 439 1035 445 1036
rect 439 1031 440 1035
rect 444 1034 445 1035
rect 463 1035 469 1036
rect 463 1034 464 1035
rect 444 1032 464 1034
rect 444 1031 445 1032
rect 439 1030 445 1031
rect 463 1031 464 1032
rect 468 1031 469 1035
rect 463 1030 469 1031
rect 630 1035 637 1036
rect 630 1031 631 1035
rect 636 1031 637 1035
rect 630 1030 637 1031
rect 775 1035 781 1036
rect 775 1031 776 1035
rect 780 1034 781 1035
rect 799 1035 805 1036
rect 799 1034 800 1035
rect 780 1032 800 1034
rect 780 1031 781 1032
rect 775 1030 781 1031
rect 799 1031 800 1032
rect 804 1031 805 1035
rect 799 1030 805 1031
rect 958 1035 965 1036
rect 958 1031 959 1035
rect 964 1031 965 1035
rect 958 1030 965 1031
rect 1095 1035 1101 1036
rect 1095 1031 1096 1035
rect 1100 1034 1101 1035
rect 1119 1035 1125 1036
rect 1119 1034 1120 1035
rect 1100 1032 1120 1034
rect 1100 1031 1101 1032
rect 1095 1030 1101 1031
rect 1119 1031 1120 1032
rect 1124 1031 1125 1035
rect 1119 1030 1125 1031
rect 1242 1035 1248 1036
rect 1242 1031 1243 1035
rect 1247 1034 1248 1035
rect 1271 1035 1277 1036
rect 1271 1034 1272 1035
rect 1247 1032 1272 1034
rect 1247 1031 1248 1032
rect 1242 1030 1248 1031
rect 1271 1031 1272 1032
rect 1276 1031 1277 1035
rect 1271 1030 1277 1031
rect 1423 1035 1429 1036
rect 1423 1031 1424 1035
rect 1428 1034 1429 1035
rect 1434 1035 1440 1036
rect 1434 1034 1435 1035
rect 1428 1032 1435 1034
rect 1428 1031 1429 1032
rect 1423 1030 1429 1031
rect 1434 1031 1435 1032
rect 1439 1031 1440 1035
rect 1434 1030 1440 1031
rect 1551 1035 1557 1036
rect 1551 1031 1552 1035
rect 1556 1034 1557 1035
rect 1575 1035 1581 1036
rect 1575 1034 1576 1035
rect 1556 1032 1576 1034
rect 1556 1031 1557 1032
rect 1551 1030 1557 1031
rect 1575 1031 1576 1032
rect 1580 1031 1581 1035
rect 1575 1030 1581 1031
rect 1911 1035 1917 1036
rect 1911 1031 1912 1035
rect 1916 1034 1917 1035
rect 1990 1035 1996 1036
rect 1990 1034 1991 1035
rect 1916 1032 1991 1034
rect 1916 1031 1917 1032
rect 1911 1030 1917 1031
rect 1990 1031 1991 1032
rect 1995 1031 1996 1035
rect 1990 1030 1996 1031
rect 2063 1035 2069 1036
rect 2063 1031 2064 1035
rect 2068 1034 2069 1035
rect 2074 1035 2080 1036
rect 2074 1034 2075 1035
rect 2068 1032 2075 1034
rect 2068 1031 2069 1032
rect 2063 1030 2069 1031
rect 2074 1031 2075 1032
rect 2079 1031 2080 1035
rect 2074 1030 2080 1031
rect 2231 1035 2237 1036
rect 2231 1031 2232 1035
rect 2236 1034 2237 1035
rect 2282 1035 2288 1036
rect 2282 1034 2283 1035
rect 2236 1032 2283 1034
rect 2236 1031 2237 1032
rect 2231 1030 2237 1031
rect 2282 1031 2283 1032
rect 2287 1031 2288 1035
rect 2282 1030 2288 1031
rect 2407 1035 2413 1036
rect 2407 1031 2408 1035
rect 2412 1034 2413 1035
rect 2418 1035 2424 1036
rect 2418 1034 2419 1035
rect 2412 1032 2419 1034
rect 2412 1031 2413 1032
rect 2407 1030 2413 1031
rect 2418 1031 2419 1032
rect 2423 1031 2424 1035
rect 2418 1030 2424 1031
rect 2582 1035 2589 1036
rect 2582 1031 2583 1035
rect 2588 1031 2589 1035
rect 2582 1030 2589 1031
rect 2703 1035 2709 1036
rect 2703 1031 2704 1035
rect 2708 1034 2709 1035
rect 2751 1035 2757 1036
rect 2751 1034 2752 1035
rect 2708 1032 2752 1034
rect 2708 1031 2709 1032
rect 2703 1030 2709 1031
rect 2751 1031 2752 1032
rect 2756 1031 2757 1035
rect 2751 1030 2757 1031
rect 2911 1035 2917 1036
rect 2911 1031 2912 1035
rect 2916 1034 2917 1035
rect 2962 1035 2968 1036
rect 2962 1034 2963 1035
rect 2916 1032 2963 1034
rect 2916 1031 2917 1032
rect 2911 1030 2917 1031
rect 2962 1031 2963 1032
rect 2967 1031 2968 1035
rect 2962 1030 2968 1031
rect 3063 1035 3069 1036
rect 3063 1031 3064 1035
rect 3068 1034 3069 1035
rect 3114 1035 3120 1036
rect 3114 1034 3115 1035
rect 3068 1032 3115 1034
rect 3068 1031 3069 1032
rect 3063 1030 3069 1031
rect 3114 1031 3115 1032
rect 3119 1031 3120 1035
rect 3114 1030 3120 1031
rect 3215 1035 3221 1036
rect 3215 1031 3216 1035
rect 3220 1034 3221 1035
rect 3266 1035 3272 1036
rect 3266 1034 3267 1035
rect 3220 1032 3267 1034
rect 3220 1031 3221 1032
rect 3215 1030 3221 1031
rect 3266 1031 3267 1032
rect 3271 1031 3272 1035
rect 3266 1030 3272 1031
rect 3366 1035 3373 1036
rect 3366 1031 3367 1035
rect 3372 1031 3373 1035
rect 3366 1030 3373 1031
rect 3495 1035 3501 1036
rect 3495 1031 3496 1035
rect 3500 1034 3501 1035
rect 3522 1035 3528 1036
rect 3522 1034 3523 1035
rect 3500 1032 3523 1034
rect 3500 1031 3501 1032
rect 3495 1030 3501 1031
rect 3522 1031 3523 1032
rect 3527 1031 3528 1035
rect 3522 1030 3528 1031
rect 151 1019 157 1020
rect 151 1015 152 1019
rect 156 1018 157 1019
rect 246 1019 252 1020
rect 246 1018 247 1019
rect 156 1016 247 1018
rect 156 1015 157 1016
rect 151 1014 157 1015
rect 246 1015 247 1016
rect 251 1015 252 1019
rect 246 1014 252 1015
rect 255 1019 261 1020
rect 255 1015 256 1019
rect 260 1018 261 1019
rect 295 1019 301 1020
rect 295 1018 296 1019
rect 260 1016 296 1018
rect 260 1015 261 1016
rect 255 1014 261 1015
rect 295 1015 296 1016
rect 300 1015 301 1019
rect 295 1014 301 1015
rect 479 1019 485 1020
rect 479 1015 480 1019
rect 484 1018 485 1019
rect 514 1019 520 1020
rect 514 1018 515 1019
rect 484 1016 515 1018
rect 484 1015 485 1016
rect 479 1014 485 1015
rect 514 1015 515 1016
rect 519 1015 520 1019
rect 514 1014 520 1015
rect 575 1019 581 1020
rect 575 1015 576 1019
rect 580 1018 581 1019
rect 671 1019 677 1020
rect 671 1018 672 1019
rect 580 1016 672 1018
rect 580 1015 581 1016
rect 575 1014 581 1015
rect 671 1015 672 1016
rect 676 1015 677 1019
rect 671 1014 677 1015
rect 759 1019 765 1020
rect 759 1015 760 1019
rect 764 1018 765 1019
rect 855 1019 861 1020
rect 855 1018 856 1019
rect 764 1016 856 1018
rect 764 1015 765 1016
rect 759 1014 765 1015
rect 855 1015 856 1016
rect 860 1015 861 1019
rect 855 1014 861 1015
rect 1039 1019 1045 1020
rect 1039 1015 1040 1019
rect 1044 1018 1045 1019
rect 1118 1019 1124 1020
rect 1118 1018 1119 1019
rect 1044 1016 1119 1018
rect 1044 1015 1045 1016
rect 1039 1014 1045 1015
rect 1118 1015 1119 1016
rect 1123 1015 1124 1019
rect 1118 1014 1124 1015
rect 1127 1019 1133 1020
rect 1127 1015 1128 1019
rect 1132 1018 1133 1019
rect 1215 1019 1221 1020
rect 1215 1018 1216 1019
rect 1132 1016 1216 1018
rect 1132 1015 1133 1016
rect 1127 1014 1133 1015
rect 1215 1015 1216 1016
rect 1220 1015 1221 1019
rect 1215 1014 1221 1015
rect 1295 1019 1301 1020
rect 1295 1015 1296 1019
rect 1300 1018 1301 1019
rect 1383 1019 1389 1020
rect 1383 1018 1384 1019
rect 1300 1016 1384 1018
rect 1300 1015 1301 1016
rect 1295 1014 1301 1015
rect 1383 1015 1384 1016
rect 1388 1015 1389 1019
rect 1383 1014 1389 1015
rect 1551 1019 1557 1020
rect 1551 1015 1552 1019
rect 1556 1018 1557 1019
rect 1610 1019 1616 1020
rect 1610 1018 1611 1019
rect 1556 1016 1611 1018
rect 1556 1015 1557 1016
rect 1551 1014 1557 1015
rect 1610 1015 1611 1016
rect 1615 1015 1616 1019
rect 1610 1014 1616 1015
rect 1718 1019 1725 1020
rect 1718 1015 1719 1019
rect 1724 1015 1725 1019
rect 1718 1014 1725 1015
rect 1982 1019 1989 1020
rect 1982 1015 1983 1019
rect 1988 1015 1989 1019
rect 1982 1014 1989 1015
rect 2066 1019 2072 1020
rect 2066 1015 2067 1019
rect 2071 1018 2072 1019
rect 2103 1019 2109 1020
rect 2103 1018 2104 1019
rect 2071 1016 2104 1018
rect 2071 1015 2072 1016
rect 2066 1014 2072 1015
rect 2103 1015 2104 1016
rect 2108 1015 2109 1019
rect 2103 1014 2109 1015
rect 2167 1019 2173 1020
rect 2167 1015 2168 1019
rect 2172 1018 2173 1019
rect 2231 1019 2237 1020
rect 2231 1018 2232 1019
rect 2172 1016 2232 1018
rect 2172 1015 2173 1016
rect 2167 1014 2173 1015
rect 2231 1015 2232 1016
rect 2236 1015 2237 1019
rect 2231 1014 2237 1015
rect 2295 1019 2301 1020
rect 2295 1015 2296 1019
rect 2300 1018 2301 1019
rect 2367 1019 2373 1020
rect 2367 1018 2368 1019
rect 2300 1016 2368 1018
rect 2300 1015 2301 1016
rect 2295 1014 2301 1015
rect 2367 1015 2368 1016
rect 2372 1015 2373 1019
rect 2367 1014 2373 1015
rect 2503 1019 2512 1020
rect 2503 1015 2504 1019
rect 2511 1015 2512 1019
rect 2503 1014 2512 1015
rect 2647 1019 2653 1020
rect 2647 1015 2648 1019
rect 2652 1018 2653 1019
rect 2682 1019 2688 1020
rect 2682 1018 2683 1019
rect 2652 1016 2683 1018
rect 2652 1015 2653 1016
rect 2647 1014 2653 1015
rect 2682 1015 2683 1016
rect 2687 1015 2688 1019
rect 2682 1014 2688 1015
rect 2799 1019 2808 1020
rect 2799 1015 2800 1019
rect 2807 1015 2808 1019
rect 2799 1014 2808 1015
rect 2903 1019 2909 1020
rect 2903 1015 2904 1019
rect 2908 1018 2909 1019
rect 2967 1019 2973 1020
rect 2967 1018 2968 1019
rect 2908 1016 2968 1018
rect 2908 1015 2909 1016
rect 2903 1014 2909 1015
rect 2967 1015 2968 1016
rect 2972 1015 2973 1019
rect 2967 1014 2973 1015
rect 3055 1019 3061 1020
rect 3055 1015 3056 1019
rect 3060 1018 3061 1019
rect 3143 1019 3149 1020
rect 3143 1018 3144 1019
rect 3060 1016 3144 1018
rect 3060 1015 3061 1016
rect 3055 1014 3061 1015
rect 3143 1015 3144 1016
rect 3148 1015 3149 1019
rect 3143 1014 3149 1015
rect 3231 1019 3237 1020
rect 3231 1015 3232 1019
rect 3236 1018 3237 1019
rect 3319 1019 3325 1020
rect 3319 1018 3320 1019
rect 3236 1016 3320 1018
rect 3236 1015 3237 1016
rect 3231 1014 3237 1015
rect 3319 1015 3320 1016
rect 3324 1015 3325 1019
rect 3319 1014 3325 1015
rect 3495 1019 3504 1020
rect 3495 1015 3496 1019
rect 3503 1015 3504 1019
rect 3495 1014 3504 1015
rect 142 1009 148 1010
rect 142 1005 143 1009
rect 147 1005 148 1009
rect 142 1004 148 1005
rect 286 1009 292 1010
rect 286 1005 287 1009
rect 291 1005 292 1009
rect 286 1004 292 1005
rect 470 1009 476 1010
rect 470 1005 471 1009
rect 475 1005 476 1009
rect 470 1004 476 1005
rect 662 1009 668 1010
rect 662 1005 663 1009
rect 667 1005 668 1009
rect 662 1004 668 1005
rect 846 1009 852 1010
rect 846 1005 847 1009
rect 851 1005 852 1009
rect 846 1004 852 1005
rect 1030 1009 1036 1010
rect 1030 1005 1031 1009
rect 1035 1005 1036 1009
rect 1030 1004 1036 1005
rect 1206 1009 1212 1010
rect 1206 1005 1207 1009
rect 1211 1005 1212 1009
rect 1206 1004 1212 1005
rect 1374 1009 1380 1010
rect 1374 1005 1375 1009
rect 1379 1005 1380 1009
rect 1374 1004 1380 1005
rect 1542 1009 1548 1010
rect 1542 1005 1543 1009
rect 1547 1005 1548 1009
rect 1542 1004 1548 1005
rect 1710 1009 1716 1010
rect 1710 1005 1711 1009
rect 1715 1005 1716 1009
rect 1710 1004 1716 1005
rect 1974 1009 1980 1010
rect 1974 1005 1975 1009
rect 1979 1005 1980 1009
rect 1974 1004 1980 1005
rect 2094 1009 2100 1010
rect 2094 1005 2095 1009
rect 2099 1005 2100 1009
rect 2094 1004 2100 1005
rect 2222 1009 2228 1010
rect 2222 1005 2223 1009
rect 2227 1005 2228 1009
rect 2222 1004 2228 1005
rect 2358 1009 2364 1010
rect 2358 1005 2359 1009
rect 2363 1005 2364 1009
rect 2358 1004 2364 1005
rect 2494 1009 2500 1010
rect 2494 1005 2495 1009
rect 2499 1005 2500 1009
rect 2494 1004 2500 1005
rect 2638 1009 2644 1010
rect 2638 1005 2639 1009
rect 2643 1005 2644 1009
rect 2638 1004 2644 1005
rect 2790 1009 2796 1010
rect 2790 1005 2791 1009
rect 2795 1005 2796 1009
rect 2790 1004 2796 1005
rect 2958 1009 2964 1010
rect 2958 1005 2959 1009
rect 2963 1005 2964 1009
rect 2958 1004 2964 1005
rect 3134 1009 3140 1010
rect 3134 1005 3135 1009
rect 3139 1005 3140 1009
rect 3134 1004 3140 1005
rect 3310 1009 3316 1010
rect 3310 1005 3311 1009
rect 3315 1005 3316 1009
rect 3310 1004 3316 1005
rect 3486 1009 3492 1010
rect 3486 1005 3487 1009
rect 3491 1005 3492 1009
rect 3486 1004 3492 1005
rect 110 996 116 997
rect 1822 996 1828 997
rect 110 992 111 996
rect 115 992 116 996
rect 255 995 261 996
rect 255 994 256 995
rect 197 992 256 994
rect 110 991 116 992
rect 255 991 256 992
rect 260 991 261 995
rect 575 995 581 996
rect 575 994 576 995
rect 525 992 576 994
rect 255 990 261 991
rect 575 991 576 992
rect 580 991 581 995
rect 759 995 765 996
rect 759 994 760 995
rect 717 992 760 994
rect 575 990 581 991
rect 759 991 760 992
rect 764 991 765 995
rect 1127 995 1133 996
rect 1127 994 1128 995
rect 1085 992 1128 994
rect 759 990 765 991
rect 770 991 776 992
rect 770 987 771 991
rect 775 990 776 991
rect 1127 991 1128 992
rect 1132 991 1133 995
rect 1295 995 1301 996
rect 1295 994 1296 995
rect 1261 992 1296 994
rect 1127 990 1133 991
rect 1295 991 1296 992
rect 1300 991 1301 995
rect 1434 995 1440 996
rect 1434 994 1435 995
rect 1429 992 1435 994
rect 1295 990 1301 991
rect 1434 991 1435 992
rect 1439 991 1440 995
rect 1822 992 1823 996
rect 1827 992 1828 996
rect 1434 990 1440 991
rect 1458 991 1464 992
rect 775 988 865 990
rect 775 987 776 988
rect 770 986 776 987
rect 1458 987 1459 991
rect 1463 990 1464 991
rect 1610 991 1616 992
rect 1822 991 1828 992
rect 1862 996 1868 997
rect 3574 996 3580 997
rect 1862 992 1863 996
rect 1867 992 1868 996
rect 2066 995 2072 996
rect 2066 994 2067 995
rect 2029 992 2067 994
rect 1862 991 1868 992
rect 2066 991 2067 992
rect 2071 991 2072 995
rect 2167 995 2173 996
rect 2167 994 2168 995
rect 2149 992 2168 994
rect 1463 988 1561 990
rect 1463 987 1464 988
rect 1458 986 1464 987
rect 1610 987 1611 991
rect 1615 990 1616 991
rect 2066 990 2072 991
rect 2167 991 2168 992
rect 2172 991 2173 995
rect 2295 995 2301 996
rect 2295 994 2296 995
rect 2277 992 2296 994
rect 2167 990 2173 991
rect 2295 991 2296 992
rect 2300 991 2301 995
rect 2418 995 2424 996
rect 2418 994 2419 995
rect 2413 992 2419 994
rect 2295 990 2301 991
rect 2418 991 2419 992
rect 2423 991 2424 995
rect 2703 995 2709 996
rect 2703 994 2704 995
rect 2693 992 2704 994
rect 2418 990 2424 991
rect 2703 991 2704 992
rect 2708 991 2709 995
rect 2903 995 2909 996
rect 2903 994 2904 995
rect 2845 992 2904 994
rect 2703 990 2709 991
rect 2903 991 2904 992
rect 2908 991 2909 995
rect 3055 995 3061 996
rect 3055 994 3056 995
rect 3013 992 3056 994
rect 2903 990 2909 991
rect 3055 991 3056 992
rect 3060 991 3061 995
rect 3231 995 3237 996
rect 3231 994 3232 995
rect 3189 992 3232 994
rect 3055 990 3061 991
rect 3231 991 3232 992
rect 3236 991 3237 995
rect 3574 992 3575 996
rect 3579 992 3580 996
rect 3574 991 3580 992
rect 3231 990 3237 991
rect 1615 988 1729 990
rect 1615 987 1616 988
rect 1610 986 1616 987
rect 110 979 116 980
rect 110 975 111 979
rect 115 975 116 979
rect 455 979 461 980
rect 455 978 456 979
rect 337 976 456 978
rect 110 974 116 975
rect 455 975 456 976
rect 460 975 461 979
rect 455 974 461 975
rect 1822 979 1828 980
rect 1822 975 1823 979
rect 1827 975 1828 979
rect 1822 974 1828 975
rect 1862 979 1868 980
rect 1862 975 1863 979
rect 1867 975 1868 979
rect 1862 974 1868 975
rect 3282 979 3288 980
rect 3282 975 3283 979
rect 3287 978 3288 979
rect 3486 979 3492 980
rect 3287 976 3321 978
rect 3287 975 3288 976
rect 3282 974 3288 975
rect 3486 975 3487 979
rect 3491 978 3492 979
rect 3574 979 3580 980
rect 3491 976 3497 978
rect 3491 975 3492 976
rect 3486 974 3492 975
rect 3574 975 3575 979
rect 3579 975 3580 979
rect 3574 974 3580 975
rect 134 969 140 970
rect 134 965 135 969
rect 139 965 140 969
rect 134 964 140 965
rect 278 969 284 970
rect 278 965 279 969
rect 283 965 284 969
rect 278 964 284 965
rect 462 969 468 970
rect 462 965 463 969
rect 467 965 468 969
rect 462 964 468 965
rect 654 969 660 970
rect 654 965 655 969
rect 659 965 660 969
rect 654 964 660 965
rect 838 969 844 970
rect 838 965 839 969
rect 843 965 844 969
rect 838 964 844 965
rect 1022 969 1028 970
rect 1022 965 1023 969
rect 1027 965 1028 969
rect 1022 964 1028 965
rect 1198 969 1204 970
rect 1198 965 1199 969
rect 1203 965 1204 969
rect 1198 964 1204 965
rect 1366 969 1372 970
rect 1366 965 1367 969
rect 1371 965 1372 969
rect 1366 964 1372 965
rect 1534 969 1540 970
rect 1534 965 1535 969
rect 1539 965 1540 969
rect 1534 964 1540 965
rect 1702 969 1708 970
rect 1702 965 1703 969
rect 1707 965 1708 969
rect 1702 964 1708 965
rect 1966 969 1972 970
rect 1966 965 1967 969
rect 1971 965 1972 969
rect 1966 964 1972 965
rect 2086 969 2092 970
rect 2086 965 2087 969
rect 2091 965 2092 969
rect 2086 964 2092 965
rect 2214 969 2220 970
rect 2214 965 2215 969
rect 2219 965 2220 969
rect 2214 964 2220 965
rect 2350 969 2356 970
rect 2350 965 2351 969
rect 2355 965 2356 969
rect 2350 964 2356 965
rect 2486 969 2492 970
rect 2486 965 2487 969
rect 2491 965 2492 969
rect 2486 964 2492 965
rect 2630 969 2636 970
rect 2630 965 2631 969
rect 2635 965 2636 969
rect 2630 964 2636 965
rect 2782 969 2788 970
rect 2782 965 2783 969
rect 2787 965 2788 969
rect 2782 964 2788 965
rect 2950 969 2956 970
rect 2950 965 2951 969
rect 2955 965 2956 969
rect 2950 964 2956 965
rect 3126 969 3132 970
rect 3126 965 3127 969
rect 3131 965 3132 969
rect 3126 964 3132 965
rect 3302 969 3308 970
rect 3302 965 3303 969
rect 3307 965 3308 969
rect 3302 964 3308 965
rect 3478 969 3484 970
rect 3478 965 3479 969
rect 3483 965 3484 969
rect 3478 964 3484 965
rect 2522 963 2528 964
rect 2522 959 2523 963
rect 2527 962 2528 963
rect 2535 963 2541 964
rect 2535 962 2536 963
rect 2527 960 2536 962
rect 2527 959 2528 960
rect 2522 958 2528 959
rect 2535 959 2536 960
rect 2540 959 2541 963
rect 2535 958 2541 959
rect 134 943 140 944
rect 134 939 135 943
rect 139 939 140 943
rect 134 938 140 939
rect 286 943 292 944
rect 286 939 287 943
rect 291 939 292 943
rect 286 938 292 939
rect 470 943 476 944
rect 470 939 471 943
rect 475 939 476 943
rect 470 938 476 939
rect 662 943 668 944
rect 662 939 663 943
rect 667 939 668 943
rect 662 938 668 939
rect 854 943 860 944
rect 854 939 855 943
rect 859 939 860 943
rect 854 938 860 939
rect 1046 943 1052 944
rect 1046 939 1047 943
rect 1051 939 1052 943
rect 1046 938 1052 939
rect 1222 943 1228 944
rect 1222 939 1223 943
rect 1227 939 1228 943
rect 1222 938 1228 939
rect 1398 943 1404 944
rect 1398 939 1399 943
rect 1403 939 1404 943
rect 1398 938 1404 939
rect 1574 943 1580 944
rect 1574 939 1575 943
rect 1579 939 1580 943
rect 1574 938 1580 939
rect 1726 943 1732 944
rect 1726 939 1727 943
rect 1731 939 1732 943
rect 1726 938 1732 939
rect 2142 943 2148 944
rect 2142 939 2143 943
rect 2147 939 2148 943
rect 2142 938 2148 939
rect 2230 943 2236 944
rect 2230 939 2231 943
rect 2235 939 2236 943
rect 2230 938 2236 939
rect 2318 943 2324 944
rect 2318 939 2319 943
rect 2323 939 2324 943
rect 2318 938 2324 939
rect 2406 943 2412 944
rect 2406 939 2407 943
rect 2411 939 2412 943
rect 2406 938 2412 939
rect 2502 943 2508 944
rect 2502 939 2503 943
rect 2507 939 2508 943
rect 2502 938 2508 939
rect 2614 943 2620 944
rect 2614 939 2615 943
rect 2619 939 2620 943
rect 2614 938 2620 939
rect 2750 943 2756 944
rect 2750 939 2751 943
rect 2755 939 2756 943
rect 2750 938 2756 939
rect 2902 943 2908 944
rect 2902 939 2903 943
rect 2907 939 2908 943
rect 2902 938 2908 939
rect 3078 943 3084 944
rect 3078 939 3079 943
rect 3083 939 3084 943
rect 3078 938 3084 939
rect 3262 943 3268 944
rect 3262 939 3263 943
rect 3267 939 3268 943
rect 3262 938 3268 939
rect 3454 943 3460 944
rect 3454 939 3455 943
rect 3459 939 3460 943
rect 3454 938 3460 939
rect 798 935 804 936
rect 110 933 116 934
rect 110 929 111 933
rect 115 929 116 933
rect 798 931 799 935
rect 803 934 804 935
rect 1718 935 1724 936
rect 803 932 873 934
rect 803 931 804 932
rect 798 930 804 931
rect 1718 931 1719 935
rect 1723 934 1724 935
rect 2682 935 2688 936
rect 2682 934 2683 935
rect 1723 932 1745 934
rect 1822 933 1828 934
rect 1723 931 1724 932
rect 1718 930 1724 931
rect 110 928 116 929
rect 1822 929 1823 933
rect 1827 929 1828 933
rect 1822 928 1828 929
rect 1862 933 1868 934
rect 1862 929 1863 933
rect 1867 929 1868 933
rect 2673 932 2683 934
rect 2682 931 2683 932
rect 2687 931 2688 935
rect 3522 935 3528 936
rect 3522 934 3523 935
rect 3513 932 3523 934
rect 2682 930 2688 931
rect 3522 931 3523 932
rect 3527 931 3528 935
rect 3522 930 3528 931
rect 3574 933 3580 934
rect 1862 928 1868 929
rect 3574 929 3575 933
rect 3579 929 3580 933
rect 3574 928 3580 929
rect 127 919 133 920
rect 110 916 116 917
rect 110 912 111 916
rect 115 912 116 916
rect 127 915 128 919
rect 132 918 133 919
rect 202 919 208 920
rect 132 916 161 918
rect 132 915 133 916
rect 127 914 133 915
rect 202 915 203 919
rect 207 918 208 919
rect 655 919 661 920
rect 655 918 656 919
rect 207 916 313 918
rect 533 916 656 918
rect 207 915 208 916
rect 202 914 208 915
rect 655 915 656 916
rect 660 915 661 919
rect 847 919 853 920
rect 847 918 848 919
rect 725 916 848 918
rect 655 914 661 915
rect 847 915 848 916
rect 852 915 853 919
rect 1215 919 1221 920
rect 1215 918 1216 919
rect 1109 916 1216 918
rect 847 914 853 915
rect 1215 915 1216 916
rect 1220 915 1221 919
rect 1391 919 1397 920
rect 1391 918 1392 919
rect 1285 916 1392 918
rect 1215 914 1221 915
rect 1391 915 1392 916
rect 1396 915 1397 919
rect 1567 919 1573 920
rect 1567 918 1568 919
rect 1461 916 1568 918
rect 1391 914 1397 915
rect 1567 915 1568 916
rect 1572 915 1573 919
rect 1719 919 1725 920
rect 1719 918 1720 919
rect 1637 916 1720 918
rect 1567 914 1573 915
rect 1719 915 1720 916
rect 1724 915 1725 919
rect 2119 919 2125 920
rect 1719 914 1725 915
rect 1822 916 1828 917
rect 110 911 116 912
rect 1822 912 1823 916
rect 1827 912 1828 916
rect 1822 911 1828 912
rect 1862 916 1868 917
rect 1862 912 1863 916
rect 1867 912 1868 916
rect 2119 915 2120 919
rect 2124 918 2125 919
rect 2210 919 2216 920
rect 2124 916 2169 918
rect 2124 915 2125 916
rect 2119 914 2125 915
rect 2210 915 2211 919
rect 2215 918 2216 919
rect 2298 919 2304 920
rect 2215 916 2257 918
rect 2215 915 2216 916
rect 2210 914 2216 915
rect 2298 915 2299 919
rect 2303 918 2304 919
rect 2386 919 2392 920
rect 2303 916 2345 918
rect 2303 915 2304 916
rect 2298 914 2304 915
rect 2386 915 2387 919
rect 2391 918 2392 919
rect 2474 919 2480 920
rect 2391 916 2433 918
rect 2391 915 2392 916
rect 2386 914 2392 915
rect 2474 915 2475 919
rect 2479 918 2480 919
rect 2682 919 2688 920
rect 2479 916 2529 918
rect 2479 915 2480 916
rect 2474 914 2480 915
rect 2682 915 2683 919
rect 2687 918 2688 919
rect 2818 919 2824 920
rect 2687 916 2777 918
rect 2687 915 2688 916
rect 2682 914 2688 915
rect 2818 915 2819 919
rect 2823 918 2824 919
rect 2970 919 2976 920
rect 2823 916 2929 918
rect 2823 915 2824 916
rect 2818 914 2824 915
rect 2970 915 2971 919
rect 2975 918 2976 919
rect 3146 919 3152 920
rect 2975 916 3105 918
rect 2975 915 2976 916
rect 2970 914 2976 915
rect 3146 915 3147 919
rect 3151 918 3152 919
rect 3151 916 3289 918
rect 3574 916 3580 917
rect 3151 915 3152 916
rect 3146 914 3152 915
rect 1862 911 1868 912
rect 3574 912 3575 916
rect 3579 912 3580 916
rect 3574 911 3580 912
rect 142 903 148 904
rect 142 899 143 903
rect 147 899 148 903
rect 142 898 148 899
rect 294 903 300 904
rect 294 899 295 903
rect 299 899 300 903
rect 294 898 300 899
rect 478 903 484 904
rect 478 899 479 903
rect 483 899 484 903
rect 478 898 484 899
rect 670 903 676 904
rect 670 899 671 903
rect 675 899 676 903
rect 670 898 676 899
rect 862 903 868 904
rect 862 899 863 903
rect 867 899 868 903
rect 862 898 868 899
rect 1054 903 1060 904
rect 1054 899 1055 903
rect 1059 899 1060 903
rect 1054 898 1060 899
rect 1230 903 1236 904
rect 1230 899 1231 903
rect 1235 899 1236 903
rect 1230 898 1236 899
rect 1406 903 1412 904
rect 1406 899 1407 903
rect 1411 899 1412 903
rect 1406 898 1412 899
rect 1582 903 1588 904
rect 1582 899 1583 903
rect 1587 899 1588 903
rect 1582 898 1588 899
rect 1734 903 1740 904
rect 1734 899 1735 903
rect 1739 899 1740 903
rect 1734 898 1740 899
rect 2150 903 2156 904
rect 2150 899 2151 903
rect 2155 899 2156 903
rect 2150 898 2156 899
rect 2238 903 2244 904
rect 2238 899 2239 903
rect 2243 899 2244 903
rect 2238 898 2244 899
rect 2326 903 2332 904
rect 2326 899 2327 903
rect 2331 899 2332 903
rect 2326 898 2332 899
rect 2414 903 2420 904
rect 2414 899 2415 903
rect 2419 899 2420 903
rect 2414 898 2420 899
rect 2510 903 2516 904
rect 2510 899 2511 903
rect 2515 899 2516 903
rect 2510 898 2516 899
rect 2622 903 2628 904
rect 2622 899 2623 903
rect 2627 899 2628 903
rect 2622 898 2628 899
rect 2758 903 2764 904
rect 2758 899 2759 903
rect 2763 899 2764 903
rect 2758 898 2764 899
rect 2910 903 2916 904
rect 2910 899 2911 903
rect 2915 899 2916 903
rect 2910 898 2916 899
rect 3086 903 3092 904
rect 3086 899 3087 903
rect 3091 899 3092 903
rect 3086 898 3092 899
rect 3270 903 3276 904
rect 3270 899 3271 903
rect 3275 899 3276 903
rect 3270 898 3276 899
rect 3462 903 3468 904
rect 3462 899 3463 903
rect 3467 899 3468 903
rect 3462 898 3468 899
rect 151 891 157 892
rect 151 887 152 891
rect 156 890 157 891
rect 202 891 208 892
rect 202 890 203 891
rect 156 888 203 890
rect 156 887 157 888
rect 151 886 157 887
rect 202 887 203 888
rect 207 887 208 891
rect 202 886 208 887
rect 302 891 309 892
rect 302 887 303 891
rect 308 887 309 891
rect 302 886 309 887
rect 455 891 461 892
rect 455 887 456 891
rect 460 890 461 891
rect 487 891 493 892
rect 487 890 488 891
rect 460 888 488 890
rect 460 887 461 888
rect 455 886 461 887
rect 487 887 488 888
rect 492 887 493 891
rect 487 886 493 887
rect 655 891 661 892
rect 655 887 656 891
rect 660 890 661 891
rect 679 891 685 892
rect 679 890 680 891
rect 660 888 680 890
rect 660 887 661 888
rect 655 886 661 887
rect 679 887 680 888
rect 684 887 685 891
rect 679 886 685 887
rect 847 891 853 892
rect 847 887 848 891
rect 852 890 853 891
rect 871 891 877 892
rect 871 890 872 891
rect 852 888 872 890
rect 852 887 853 888
rect 847 886 853 887
rect 871 887 872 888
rect 876 887 877 891
rect 871 886 877 887
rect 1063 891 1069 892
rect 1063 887 1064 891
rect 1068 890 1069 891
rect 1206 891 1212 892
rect 1206 890 1207 891
rect 1068 888 1207 890
rect 1068 887 1069 888
rect 1063 886 1069 887
rect 1206 887 1207 888
rect 1211 887 1212 891
rect 1206 886 1212 887
rect 1215 891 1221 892
rect 1215 887 1216 891
rect 1220 890 1221 891
rect 1239 891 1245 892
rect 1239 890 1240 891
rect 1220 888 1240 890
rect 1220 887 1221 888
rect 1215 886 1221 887
rect 1239 887 1240 888
rect 1244 887 1245 891
rect 1239 886 1245 887
rect 1391 891 1397 892
rect 1391 887 1392 891
rect 1396 890 1397 891
rect 1415 891 1421 892
rect 1415 890 1416 891
rect 1396 888 1416 890
rect 1396 887 1397 888
rect 1391 886 1397 887
rect 1415 887 1416 888
rect 1420 887 1421 891
rect 1415 886 1421 887
rect 1567 891 1573 892
rect 1567 887 1568 891
rect 1572 890 1573 891
rect 1591 891 1597 892
rect 1591 890 1592 891
rect 1572 888 1592 890
rect 1572 887 1573 888
rect 1567 886 1573 887
rect 1591 887 1592 888
rect 1596 887 1597 891
rect 1591 886 1597 887
rect 1719 891 1725 892
rect 1719 887 1720 891
rect 1724 890 1725 891
rect 1743 891 1749 892
rect 1743 890 1744 891
rect 1724 888 1744 890
rect 1724 887 1725 888
rect 1719 886 1725 887
rect 1743 887 1744 888
rect 1748 887 1749 891
rect 1743 886 1749 887
rect 2159 891 2165 892
rect 2159 887 2160 891
rect 2164 890 2165 891
rect 2210 891 2216 892
rect 2210 890 2211 891
rect 2164 888 2211 890
rect 2164 887 2165 888
rect 2159 886 2165 887
rect 2210 887 2211 888
rect 2215 887 2216 891
rect 2210 886 2216 887
rect 2247 891 2253 892
rect 2247 887 2248 891
rect 2252 890 2253 891
rect 2298 891 2304 892
rect 2298 890 2299 891
rect 2252 888 2299 890
rect 2252 887 2253 888
rect 2247 886 2253 887
rect 2298 887 2299 888
rect 2303 887 2304 891
rect 2298 886 2304 887
rect 2335 891 2341 892
rect 2335 887 2336 891
rect 2340 890 2341 891
rect 2386 891 2392 892
rect 2386 890 2387 891
rect 2340 888 2387 890
rect 2340 887 2341 888
rect 2335 886 2341 887
rect 2386 887 2387 888
rect 2391 887 2392 891
rect 2386 886 2392 887
rect 2423 891 2429 892
rect 2423 887 2424 891
rect 2428 890 2429 891
rect 2474 891 2480 892
rect 2474 890 2475 891
rect 2428 888 2475 890
rect 2428 887 2429 888
rect 2423 886 2429 887
rect 2474 887 2475 888
rect 2479 887 2480 891
rect 2474 886 2480 887
rect 2519 891 2528 892
rect 2519 887 2520 891
rect 2527 887 2528 891
rect 2519 886 2528 887
rect 2551 891 2557 892
rect 2551 887 2552 891
rect 2556 890 2557 891
rect 2631 891 2637 892
rect 2631 890 2632 891
rect 2556 888 2632 890
rect 2556 887 2557 888
rect 2551 886 2557 887
rect 2631 887 2632 888
rect 2636 887 2637 891
rect 2631 886 2637 887
rect 2767 891 2773 892
rect 2767 887 2768 891
rect 2772 890 2773 891
rect 2818 891 2824 892
rect 2818 890 2819 891
rect 2772 888 2819 890
rect 2772 887 2773 888
rect 2767 886 2773 887
rect 2818 887 2819 888
rect 2823 887 2824 891
rect 2818 886 2824 887
rect 2919 891 2925 892
rect 2919 887 2920 891
rect 2924 890 2925 891
rect 2970 891 2976 892
rect 2970 890 2971 891
rect 2924 888 2971 890
rect 2924 887 2925 888
rect 2919 886 2925 887
rect 2970 887 2971 888
rect 2975 887 2976 891
rect 2970 886 2976 887
rect 3095 891 3101 892
rect 3095 887 3096 891
rect 3100 890 3101 891
rect 3146 891 3152 892
rect 3146 890 3147 891
rect 3100 888 3147 890
rect 3100 887 3101 888
rect 3095 886 3101 887
rect 3146 887 3147 888
rect 3151 887 3152 891
rect 3146 886 3152 887
rect 3279 891 3288 892
rect 3279 887 3280 891
rect 3287 887 3288 891
rect 3279 886 3288 887
rect 3471 891 3477 892
rect 3471 887 3472 891
rect 3476 890 3477 891
rect 3486 891 3492 892
rect 3486 890 3487 891
rect 3476 888 3487 890
rect 3476 887 3477 888
rect 3471 886 3477 887
rect 3486 887 3487 888
rect 3491 887 3492 891
rect 3486 886 3492 887
rect 2682 883 2688 884
rect 2682 882 2683 883
rect 2633 880 2683 882
rect 127 875 133 876
rect 127 871 128 875
rect 132 874 133 875
rect 151 875 157 876
rect 151 874 152 875
rect 132 872 152 874
rect 132 871 133 872
rect 127 870 133 871
rect 151 871 152 872
rect 156 871 157 875
rect 151 870 157 871
rect 223 875 229 876
rect 223 871 224 875
rect 228 874 229 875
rect 295 875 301 876
rect 295 874 296 875
rect 228 872 296 874
rect 228 871 229 872
rect 223 870 229 871
rect 295 871 296 872
rect 300 871 301 875
rect 295 870 301 871
rect 455 875 461 876
rect 455 871 456 875
rect 460 874 461 875
rect 479 875 485 876
rect 479 874 480 875
rect 460 872 480 874
rect 460 871 461 872
rect 455 870 461 871
rect 479 871 480 872
rect 484 871 485 875
rect 479 870 485 871
rect 567 875 573 876
rect 567 871 568 875
rect 572 874 573 875
rect 663 875 669 876
rect 663 874 664 875
rect 572 872 664 874
rect 572 871 573 872
rect 567 870 573 871
rect 663 871 664 872
rect 668 871 669 875
rect 663 870 669 871
rect 751 875 757 876
rect 751 871 752 875
rect 756 874 757 875
rect 847 875 853 876
rect 847 874 848 875
rect 756 872 848 874
rect 756 871 757 872
rect 751 870 757 871
rect 847 871 848 872
rect 852 871 853 875
rect 847 870 853 871
rect 1031 875 1037 876
rect 1031 871 1032 875
rect 1036 874 1037 875
rect 1086 875 1092 876
rect 1086 874 1087 875
rect 1036 872 1087 874
rect 1036 871 1037 872
rect 1031 870 1037 871
rect 1086 871 1087 872
rect 1091 871 1092 875
rect 1086 870 1092 871
rect 1095 875 1101 876
rect 1095 871 1096 875
rect 1100 874 1101 875
rect 1199 875 1205 876
rect 1199 874 1200 875
rect 1100 872 1200 874
rect 1100 871 1101 872
rect 1095 870 1101 871
rect 1199 871 1200 872
rect 1204 871 1205 875
rect 1199 870 1205 871
rect 1279 875 1285 876
rect 1279 871 1280 875
rect 1284 874 1285 875
rect 1367 875 1373 876
rect 1367 874 1368 875
rect 1284 872 1368 874
rect 1284 871 1285 872
rect 1279 870 1285 871
rect 1367 871 1368 872
rect 1372 871 1373 875
rect 1367 870 1373 871
rect 1447 875 1453 876
rect 1447 871 1448 875
rect 1452 874 1453 875
rect 1535 875 1541 876
rect 1535 874 1536 875
rect 1452 872 1536 874
rect 1452 871 1453 872
rect 1447 870 1453 871
rect 1535 871 1536 872
rect 1540 871 1541 875
rect 1535 870 1541 871
rect 1615 875 1621 876
rect 1615 871 1616 875
rect 1620 874 1621 875
rect 1703 875 1709 876
rect 1703 874 1704 875
rect 1620 872 1704 874
rect 1620 871 1621 872
rect 1615 870 1621 871
rect 1703 871 1704 872
rect 1708 871 1709 875
rect 1703 870 1709 871
rect 2111 875 2117 876
rect 2111 871 2112 875
rect 2116 874 2117 875
rect 2119 875 2125 876
rect 2119 874 2120 875
rect 2116 872 2120 874
rect 2116 871 2117 872
rect 2111 870 2117 871
rect 2119 871 2120 872
rect 2124 871 2125 875
rect 2119 870 2125 871
rect 2167 875 2173 876
rect 2167 871 2168 875
rect 2172 874 2173 875
rect 2199 875 2205 876
rect 2199 874 2200 875
rect 2172 872 2200 874
rect 2172 871 2173 872
rect 2167 870 2173 871
rect 2199 871 2200 872
rect 2204 871 2205 875
rect 2199 870 2205 871
rect 2255 875 2261 876
rect 2255 871 2256 875
rect 2260 874 2261 875
rect 2287 875 2293 876
rect 2287 874 2288 875
rect 2260 872 2288 874
rect 2260 871 2261 872
rect 2255 870 2261 871
rect 2287 871 2288 872
rect 2292 871 2293 875
rect 2287 870 2293 871
rect 2375 875 2381 876
rect 2375 871 2376 875
rect 2380 874 2381 875
rect 2431 875 2437 876
rect 2380 872 2426 874
rect 2380 871 2381 872
rect 2375 870 2381 871
rect 2424 866 2426 872
rect 2431 871 2432 875
rect 2436 874 2437 875
rect 2463 875 2469 876
rect 2463 874 2464 875
rect 2436 872 2464 874
rect 2436 871 2437 872
rect 2431 870 2437 871
rect 2463 871 2464 872
rect 2468 871 2469 875
rect 2463 870 2469 871
rect 2575 875 2581 876
rect 2575 871 2576 875
rect 2580 874 2581 875
rect 2633 874 2635 880
rect 2682 879 2683 880
rect 2687 879 2688 883
rect 2682 878 2688 879
rect 2580 872 2635 874
rect 2639 875 2645 876
rect 2580 871 2581 872
rect 2575 870 2581 871
rect 2639 871 2640 875
rect 2644 874 2645 875
rect 2711 875 2717 876
rect 2711 874 2712 875
rect 2644 872 2712 874
rect 2644 871 2645 872
rect 2639 870 2645 871
rect 2711 871 2712 872
rect 2716 871 2717 875
rect 2711 870 2717 871
rect 2775 875 2781 876
rect 2775 871 2776 875
rect 2780 874 2781 875
rect 2879 875 2885 876
rect 2879 874 2880 875
rect 2780 872 2880 874
rect 2780 871 2781 872
rect 2775 870 2781 871
rect 2879 871 2880 872
rect 2884 871 2885 875
rect 2879 870 2885 871
rect 2967 875 2973 876
rect 2967 871 2968 875
rect 2972 874 2973 875
rect 3063 875 3069 876
rect 3063 874 3064 875
rect 2972 872 3064 874
rect 2972 871 2973 872
rect 2967 870 2973 871
rect 3063 871 3064 872
rect 3068 871 3069 875
rect 3063 870 3069 871
rect 3159 875 3165 876
rect 3159 871 3160 875
rect 3164 874 3165 875
rect 3263 875 3269 876
rect 3263 874 3264 875
rect 3164 872 3264 874
rect 3164 871 3165 872
rect 3159 870 3165 871
rect 3263 871 3264 872
rect 3268 871 3269 875
rect 3263 870 3269 871
rect 3471 875 3477 876
rect 3471 871 3472 875
rect 3476 874 3477 875
rect 3506 875 3512 876
rect 3506 874 3507 875
rect 3476 872 3507 874
rect 3476 871 3477 872
rect 3471 870 3477 871
rect 3506 871 3507 872
rect 3511 871 3512 875
rect 3506 870 3512 871
rect 2438 867 2444 868
rect 2438 866 2439 867
rect 142 865 148 866
rect 142 861 143 865
rect 147 861 148 865
rect 142 860 148 861
rect 286 865 292 866
rect 286 861 287 865
rect 291 861 292 865
rect 286 860 292 861
rect 470 865 476 866
rect 470 861 471 865
rect 475 861 476 865
rect 470 860 476 861
rect 654 865 660 866
rect 654 861 655 865
rect 659 861 660 865
rect 654 860 660 861
rect 838 865 844 866
rect 838 861 839 865
rect 843 861 844 865
rect 838 860 844 861
rect 1022 865 1028 866
rect 1022 861 1023 865
rect 1027 861 1028 865
rect 1022 860 1028 861
rect 1190 865 1196 866
rect 1190 861 1191 865
rect 1195 861 1196 865
rect 1190 860 1196 861
rect 1358 865 1364 866
rect 1358 861 1359 865
rect 1363 861 1364 865
rect 1358 860 1364 861
rect 1526 865 1532 866
rect 1526 861 1527 865
rect 1531 861 1532 865
rect 1526 860 1532 861
rect 1694 865 1700 866
rect 1694 861 1695 865
rect 1699 861 1700 865
rect 1694 860 1700 861
rect 2102 865 2108 866
rect 2102 861 2103 865
rect 2107 861 2108 865
rect 2102 860 2108 861
rect 2190 865 2196 866
rect 2190 861 2191 865
rect 2195 861 2196 865
rect 2190 860 2196 861
rect 2278 865 2284 866
rect 2278 861 2279 865
rect 2283 861 2284 865
rect 2278 860 2284 861
rect 2366 865 2372 866
rect 2366 861 2367 865
rect 2371 861 2372 865
rect 2424 864 2439 866
rect 2438 863 2439 864
rect 2443 863 2444 867
rect 2438 862 2444 863
rect 2454 865 2460 866
rect 2366 860 2372 861
rect 2454 861 2455 865
rect 2459 861 2460 865
rect 2454 860 2460 861
rect 2566 865 2572 866
rect 2566 861 2567 865
rect 2571 861 2572 865
rect 2566 860 2572 861
rect 2702 865 2708 866
rect 2702 861 2703 865
rect 2707 861 2708 865
rect 2702 860 2708 861
rect 2870 865 2876 866
rect 2870 861 2871 865
rect 2875 861 2876 865
rect 2870 860 2876 861
rect 3054 865 3060 866
rect 3054 861 3055 865
rect 3059 861 3060 865
rect 3054 860 3060 861
rect 3254 865 3260 866
rect 3254 861 3255 865
rect 3259 861 3260 865
rect 3254 860 3260 861
rect 3462 865 3468 866
rect 3462 861 3463 865
rect 3467 861 3468 865
rect 3462 860 3468 861
rect 110 852 116 853
rect 1822 852 1828 853
rect 110 848 111 852
rect 115 848 116 852
rect 223 851 229 852
rect 223 850 224 851
rect 197 848 224 850
rect 110 847 116 848
rect 223 847 224 848
rect 228 847 229 851
rect 455 851 461 852
rect 455 850 456 851
rect 341 848 456 850
rect 223 846 229 847
rect 455 847 456 848
rect 460 847 461 851
rect 567 851 573 852
rect 567 850 568 851
rect 525 848 568 850
rect 455 846 461 847
rect 567 847 568 848
rect 572 847 573 851
rect 751 851 757 852
rect 751 850 752 851
rect 709 848 752 850
rect 567 846 573 847
rect 751 847 752 848
rect 756 847 757 851
rect 1095 851 1101 852
rect 1095 850 1096 851
rect 1077 848 1096 850
rect 751 846 757 847
rect 1095 847 1096 848
rect 1100 847 1101 851
rect 1279 851 1285 852
rect 1279 850 1280 851
rect 1245 848 1280 850
rect 1095 846 1101 847
rect 1279 847 1280 848
rect 1284 847 1285 851
rect 1447 851 1453 852
rect 1447 850 1448 851
rect 1413 848 1448 850
rect 1279 846 1285 847
rect 1447 847 1448 848
rect 1452 847 1453 851
rect 1615 851 1621 852
rect 1615 850 1616 851
rect 1581 848 1616 850
rect 1447 846 1453 847
rect 1615 847 1616 848
rect 1620 847 1621 851
rect 1822 848 1823 852
rect 1827 848 1828 852
rect 1615 846 1621 847
rect 1626 847 1632 848
rect 1822 847 1828 848
rect 1862 852 1868 853
rect 3574 852 3580 853
rect 1862 848 1863 852
rect 1867 848 1868 852
rect 2167 851 2173 852
rect 2167 850 2168 851
rect 2157 848 2168 850
rect 1862 847 1868 848
rect 2167 847 2168 848
rect 2172 847 2173 851
rect 2255 851 2261 852
rect 2255 850 2256 851
rect 2245 848 2256 850
rect 1626 843 1627 847
rect 1631 846 1632 847
rect 2167 846 2173 847
rect 2255 847 2256 848
rect 2260 847 2261 851
rect 2431 851 2437 852
rect 2431 850 2432 851
rect 2421 848 2432 850
rect 2255 846 2261 847
rect 2431 847 2432 848
rect 2436 847 2437 851
rect 2551 851 2557 852
rect 2551 850 2552 851
rect 2509 848 2552 850
rect 2431 846 2437 847
rect 2551 847 2552 848
rect 2556 847 2557 851
rect 2639 851 2645 852
rect 2639 850 2640 851
rect 2621 848 2640 850
rect 2551 846 2557 847
rect 2639 847 2640 848
rect 2644 847 2645 851
rect 2775 851 2781 852
rect 2775 850 2776 851
rect 2757 848 2776 850
rect 2639 846 2645 847
rect 2775 847 2776 848
rect 2780 847 2781 851
rect 2967 851 2973 852
rect 2967 850 2968 851
rect 2925 848 2968 850
rect 2775 846 2781 847
rect 2967 847 2968 848
rect 2972 847 2973 851
rect 3159 851 3165 852
rect 3159 850 3160 851
rect 3109 848 3160 850
rect 2967 846 2973 847
rect 3159 847 3160 848
rect 3164 847 3165 851
rect 3574 848 3575 852
rect 3579 848 3580 852
rect 3574 847 3580 848
rect 3159 846 3165 847
rect 1631 844 1713 846
rect 1631 843 1632 844
rect 1626 842 1632 843
rect 110 835 116 836
rect 110 831 111 835
rect 115 831 116 835
rect 110 830 116 831
rect 750 835 756 836
rect 750 831 751 835
rect 755 834 756 835
rect 1822 835 1828 836
rect 755 832 849 834
rect 755 831 756 832
rect 750 830 756 831
rect 1822 831 1823 835
rect 1827 831 1828 835
rect 1822 830 1828 831
rect 1862 835 1868 836
rect 1862 831 1863 835
rect 1867 831 1868 835
rect 1862 830 1868 831
rect 3138 835 3144 836
rect 3138 831 3139 835
rect 3143 834 3144 835
rect 3574 835 3580 836
rect 3143 832 3265 834
rect 3143 831 3144 832
rect 3138 830 3144 831
rect 3574 831 3575 835
rect 3579 831 3580 835
rect 3574 830 3580 831
rect 134 825 140 826
rect 134 821 135 825
rect 139 821 140 825
rect 134 820 140 821
rect 278 825 284 826
rect 278 821 279 825
rect 283 821 284 825
rect 278 820 284 821
rect 462 825 468 826
rect 462 821 463 825
rect 467 821 468 825
rect 462 820 468 821
rect 646 825 652 826
rect 646 821 647 825
rect 651 821 652 825
rect 646 820 652 821
rect 830 825 836 826
rect 830 821 831 825
rect 835 821 836 825
rect 830 820 836 821
rect 1014 825 1020 826
rect 1014 821 1015 825
rect 1019 821 1020 825
rect 1014 820 1020 821
rect 1182 825 1188 826
rect 1182 821 1183 825
rect 1187 821 1188 825
rect 1182 820 1188 821
rect 1350 825 1356 826
rect 1350 821 1351 825
rect 1355 821 1356 825
rect 1350 820 1356 821
rect 1518 825 1524 826
rect 1518 821 1519 825
rect 1523 821 1524 825
rect 1518 820 1524 821
rect 1686 825 1692 826
rect 1686 821 1687 825
rect 1691 821 1692 825
rect 1686 820 1692 821
rect 2094 825 2100 826
rect 2094 821 2095 825
rect 2099 821 2100 825
rect 2094 820 2100 821
rect 2182 825 2188 826
rect 2182 821 2183 825
rect 2187 821 2188 825
rect 2182 820 2188 821
rect 2270 825 2276 826
rect 2270 821 2271 825
rect 2275 821 2276 825
rect 2270 820 2276 821
rect 2358 825 2364 826
rect 2358 821 2359 825
rect 2363 821 2364 825
rect 2358 820 2364 821
rect 2446 825 2452 826
rect 2446 821 2447 825
rect 2451 821 2452 825
rect 2446 820 2452 821
rect 2558 825 2564 826
rect 2558 821 2559 825
rect 2563 821 2564 825
rect 2558 820 2564 821
rect 2694 825 2700 826
rect 2694 821 2695 825
rect 2699 821 2700 825
rect 2694 820 2700 821
rect 2862 825 2868 826
rect 2862 821 2863 825
rect 2867 821 2868 825
rect 2862 820 2868 821
rect 3046 825 3052 826
rect 3046 821 3047 825
rect 3051 821 3052 825
rect 3046 820 3052 821
rect 3246 825 3252 826
rect 3246 821 3247 825
rect 3251 821 3252 825
rect 3246 820 3252 821
rect 3454 825 3460 826
rect 3454 821 3455 825
rect 3459 821 3460 825
rect 3454 820 3460 821
rect 2306 819 2312 820
rect 2306 815 2307 819
rect 2311 818 2312 819
rect 2319 819 2325 820
rect 2319 818 2320 819
rect 2311 816 2320 818
rect 2311 815 2312 816
rect 2306 814 2312 815
rect 2319 815 2320 816
rect 2324 815 2325 819
rect 2319 814 2325 815
rect 3498 819 3509 820
rect 3498 815 3499 819
rect 3503 815 3504 819
rect 3508 815 3509 819
rect 3498 814 3509 815
rect 134 803 140 804
rect 134 799 135 803
rect 139 799 140 803
rect 134 798 140 799
rect 270 803 276 804
rect 270 799 271 803
rect 275 799 276 803
rect 270 798 276 799
rect 422 803 428 804
rect 422 799 423 803
rect 427 799 428 803
rect 422 798 428 799
rect 582 803 588 804
rect 582 799 583 803
rect 587 799 588 803
rect 582 798 588 799
rect 742 803 748 804
rect 742 799 743 803
rect 747 799 748 803
rect 742 798 748 799
rect 894 803 900 804
rect 894 799 895 803
rect 899 799 900 803
rect 894 798 900 799
rect 1038 803 1044 804
rect 1038 799 1039 803
rect 1043 799 1044 803
rect 1038 798 1044 799
rect 1182 803 1188 804
rect 1182 799 1183 803
rect 1187 799 1188 803
rect 1182 798 1188 799
rect 1326 803 1332 804
rect 1326 799 1327 803
rect 1331 799 1332 803
rect 1326 798 1332 799
rect 1478 803 1484 804
rect 1478 799 1479 803
rect 1483 799 1484 803
rect 1478 798 1484 799
rect 2198 803 2204 804
rect 2198 799 2199 803
rect 2203 799 2204 803
rect 2198 798 2204 799
rect 2286 803 2292 804
rect 2286 799 2287 803
rect 2291 799 2292 803
rect 2286 798 2292 799
rect 2374 803 2380 804
rect 2374 799 2375 803
rect 2379 799 2380 803
rect 2374 798 2380 799
rect 2462 803 2468 804
rect 2462 799 2463 803
rect 2467 799 2468 803
rect 2462 798 2468 799
rect 2550 803 2556 804
rect 2550 799 2551 803
rect 2555 799 2556 803
rect 2550 798 2556 799
rect 2654 803 2660 804
rect 2654 799 2655 803
rect 2659 799 2660 803
rect 2654 798 2660 799
rect 2782 803 2788 804
rect 2782 799 2783 803
rect 2787 799 2788 803
rect 2782 798 2788 799
rect 2934 803 2940 804
rect 2934 799 2935 803
rect 2939 799 2940 803
rect 2934 798 2940 799
rect 3110 803 3116 804
rect 3110 799 3111 803
rect 3115 799 3116 803
rect 3110 798 3116 799
rect 3294 803 3300 804
rect 3294 799 3295 803
rect 3299 799 3300 803
rect 3294 798 3300 799
rect 3478 803 3484 804
rect 3478 799 3479 803
rect 3483 799 3484 803
rect 3478 798 3484 799
rect 678 795 684 796
rect 110 793 116 794
rect 110 789 111 793
rect 115 789 116 793
rect 678 791 679 795
rect 683 794 684 795
rect 1398 795 1404 796
rect 683 792 761 794
rect 683 791 684 792
rect 678 790 684 791
rect 1398 791 1399 795
rect 1403 794 1404 795
rect 2354 795 2360 796
rect 1403 792 1497 794
rect 1822 793 1828 794
rect 1403 791 1404 792
rect 1398 790 1404 791
rect 110 788 116 789
rect 1822 789 1823 793
rect 1827 789 1828 793
rect 1822 788 1828 789
rect 1862 793 1868 794
rect 1862 789 1863 793
rect 1867 789 1868 793
rect 2354 791 2355 795
rect 2359 794 2360 795
rect 2442 795 2448 796
rect 2359 792 2393 794
rect 2359 791 2360 792
rect 2354 790 2360 791
rect 2442 791 2443 795
rect 2447 794 2448 795
rect 3198 795 3204 796
rect 2447 792 2481 794
rect 2447 791 2448 792
rect 2442 790 2448 791
rect 3198 791 3199 795
rect 3203 794 3204 795
rect 3203 792 3313 794
rect 3574 793 3580 794
rect 3203 791 3204 792
rect 3198 790 3204 791
rect 1862 788 1868 789
rect 3574 789 3575 793
rect 3579 789 3580 793
rect 3574 788 3580 789
rect 263 779 269 780
rect 263 778 264 779
rect 110 776 116 777
rect 197 776 264 778
rect 110 772 111 776
rect 115 772 116 776
rect 263 775 264 776
rect 268 775 269 779
rect 415 779 421 780
rect 415 778 416 779
rect 333 776 416 778
rect 263 774 269 775
rect 415 775 416 776
rect 420 775 421 779
rect 575 779 581 780
rect 575 778 576 779
rect 485 776 576 778
rect 415 774 421 775
rect 575 775 576 776
rect 580 775 581 779
rect 735 779 741 780
rect 735 778 736 779
rect 645 776 736 778
rect 575 774 581 775
rect 735 775 736 776
rect 740 775 741 779
rect 1031 779 1037 780
rect 1031 778 1032 779
rect 957 776 1032 778
rect 735 774 741 775
rect 1031 775 1032 776
rect 1036 775 1037 779
rect 1175 779 1181 780
rect 1175 778 1176 779
rect 1101 776 1176 778
rect 1031 774 1037 775
rect 1175 775 1176 776
rect 1180 775 1181 779
rect 1319 779 1325 780
rect 1319 778 1320 779
rect 1245 776 1320 778
rect 1175 774 1181 775
rect 1319 775 1320 776
rect 1324 775 1325 779
rect 1471 779 1477 780
rect 1471 778 1472 779
rect 1389 776 1472 778
rect 1319 774 1325 775
rect 1471 775 1472 776
rect 1476 775 1477 779
rect 2266 779 2272 780
rect 2266 778 2267 779
rect 1471 774 1477 775
rect 1822 776 1828 777
rect 110 771 116 772
rect 1822 772 1823 776
rect 1827 772 1828 776
rect 1822 771 1828 772
rect 1862 776 1868 777
rect 2261 776 2267 778
rect 1862 772 1863 776
rect 1867 772 1868 776
rect 2266 775 2267 776
rect 2271 775 2272 779
rect 2367 779 2373 780
rect 2367 778 2368 779
rect 2349 776 2368 778
rect 2266 774 2272 775
rect 2367 775 2368 776
rect 2372 775 2373 779
rect 2367 774 2373 775
rect 2530 779 2536 780
rect 2530 775 2531 779
rect 2535 778 2536 779
rect 2775 779 2781 780
rect 2775 778 2776 779
rect 2535 776 2577 778
rect 2717 776 2776 778
rect 2535 775 2536 776
rect 2530 774 2536 775
rect 2775 775 2776 776
rect 2780 775 2781 779
rect 2927 779 2933 780
rect 2927 778 2928 779
rect 2845 776 2928 778
rect 2775 774 2781 775
rect 2927 775 2928 776
rect 2932 775 2933 779
rect 3103 779 3109 780
rect 3103 778 3104 779
rect 2997 776 3104 778
rect 2927 774 2933 775
rect 3103 775 3104 776
rect 3108 775 3109 779
rect 3287 779 3293 780
rect 3287 778 3288 779
rect 3173 776 3288 778
rect 3103 774 3109 775
rect 3287 775 3288 776
rect 3292 775 3293 779
rect 3287 774 3293 775
rect 3470 779 3476 780
rect 3470 775 3471 779
rect 3475 778 3476 779
rect 3475 776 3505 778
rect 3574 776 3580 777
rect 3475 775 3476 776
rect 3470 774 3476 775
rect 1862 771 1868 772
rect 3574 772 3575 776
rect 3579 772 3580 776
rect 3574 771 3580 772
rect 142 763 148 764
rect 142 759 143 763
rect 147 759 148 763
rect 142 758 148 759
rect 278 763 284 764
rect 278 759 279 763
rect 283 759 284 763
rect 278 758 284 759
rect 430 763 436 764
rect 430 759 431 763
rect 435 759 436 763
rect 430 758 436 759
rect 590 763 596 764
rect 590 759 591 763
rect 595 759 596 763
rect 590 758 596 759
rect 750 763 756 764
rect 750 759 751 763
rect 755 759 756 763
rect 750 758 756 759
rect 902 763 908 764
rect 902 759 903 763
rect 907 759 908 763
rect 902 758 908 759
rect 1046 763 1052 764
rect 1046 759 1047 763
rect 1051 759 1052 763
rect 1046 758 1052 759
rect 1190 763 1196 764
rect 1190 759 1191 763
rect 1195 759 1196 763
rect 1190 758 1196 759
rect 1334 763 1340 764
rect 1334 759 1335 763
rect 1339 759 1340 763
rect 1334 758 1340 759
rect 1486 763 1492 764
rect 1486 759 1487 763
rect 1491 759 1492 763
rect 1486 758 1492 759
rect 2206 763 2212 764
rect 2206 759 2207 763
rect 2211 759 2212 763
rect 2206 758 2212 759
rect 2294 763 2300 764
rect 2294 759 2295 763
rect 2299 759 2300 763
rect 2294 758 2300 759
rect 2382 763 2388 764
rect 2382 759 2383 763
rect 2387 759 2388 763
rect 2382 758 2388 759
rect 2470 763 2476 764
rect 2470 759 2471 763
rect 2475 759 2476 763
rect 2470 758 2476 759
rect 2558 763 2564 764
rect 2558 759 2559 763
rect 2563 759 2564 763
rect 2558 758 2564 759
rect 2662 763 2668 764
rect 2662 759 2663 763
rect 2667 759 2668 763
rect 2662 758 2668 759
rect 2790 763 2796 764
rect 2790 759 2791 763
rect 2795 759 2796 763
rect 2790 758 2796 759
rect 2942 763 2948 764
rect 2942 759 2943 763
rect 2947 759 2948 763
rect 2942 758 2948 759
rect 3118 763 3124 764
rect 3118 759 3119 763
rect 3123 759 3124 763
rect 3118 758 3124 759
rect 3302 763 3308 764
rect 3302 759 3303 763
rect 3307 759 3308 763
rect 3302 758 3308 759
rect 3486 763 3492 764
rect 3486 759 3487 763
rect 3491 759 3492 763
rect 3486 758 3492 759
rect 151 751 160 752
rect 151 747 152 751
rect 159 747 160 751
rect 151 746 160 747
rect 263 751 269 752
rect 263 747 264 751
rect 268 750 269 751
rect 287 751 293 752
rect 287 750 288 751
rect 268 748 288 750
rect 268 747 269 748
rect 263 746 269 747
rect 287 747 288 748
rect 292 747 293 751
rect 287 746 293 747
rect 415 751 421 752
rect 415 747 416 751
rect 420 750 421 751
rect 439 751 445 752
rect 439 750 440 751
rect 420 748 440 750
rect 420 747 421 748
rect 415 746 421 747
rect 439 747 440 748
rect 444 747 445 751
rect 439 746 445 747
rect 575 751 581 752
rect 575 747 576 751
rect 580 750 581 751
rect 599 751 605 752
rect 599 750 600 751
rect 580 748 600 750
rect 580 747 581 748
rect 575 746 581 747
rect 599 747 600 748
rect 604 747 605 751
rect 599 746 605 747
rect 735 751 741 752
rect 735 747 736 751
rect 740 750 741 751
rect 759 751 765 752
rect 759 750 760 751
rect 740 748 760 750
rect 740 747 741 748
rect 735 746 741 747
rect 759 747 760 748
rect 764 747 765 751
rect 759 746 765 747
rect 911 751 917 752
rect 911 747 912 751
rect 916 750 917 751
rect 1022 751 1028 752
rect 1022 750 1023 751
rect 916 748 1023 750
rect 916 747 917 748
rect 911 746 917 747
rect 1022 747 1023 748
rect 1027 747 1028 751
rect 1022 746 1028 747
rect 1031 751 1037 752
rect 1031 747 1032 751
rect 1036 750 1037 751
rect 1055 751 1061 752
rect 1055 750 1056 751
rect 1036 748 1056 750
rect 1036 747 1037 748
rect 1031 746 1037 747
rect 1055 747 1056 748
rect 1060 747 1061 751
rect 1055 746 1061 747
rect 1175 751 1181 752
rect 1175 747 1176 751
rect 1180 750 1181 751
rect 1199 751 1205 752
rect 1199 750 1200 751
rect 1180 748 1200 750
rect 1180 747 1181 748
rect 1175 746 1181 747
rect 1199 747 1200 748
rect 1204 747 1205 751
rect 1199 746 1205 747
rect 1319 751 1325 752
rect 1319 747 1320 751
rect 1324 750 1325 751
rect 1343 751 1349 752
rect 1343 750 1344 751
rect 1324 748 1344 750
rect 1324 747 1325 748
rect 1319 746 1325 747
rect 1343 747 1344 748
rect 1348 747 1349 751
rect 1343 746 1349 747
rect 1471 751 1477 752
rect 1471 747 1472 751
rect 1476 750 1477 751
rect 1495 751 1501 752
rect 1495 750 1496 751
rect 1476 748 1496 750
rect 1476 747 1477 748
rect 1471 746 1477 747
rect 1495 747 1496 748
rect 1500 747 1501 751
rect 1495 746 1501 747
rect 2215 751 2221 752
rect 2215 747 2216 751
rect 2220 750 2221 751
rect 2303 751 2312 752
rect 2220 748 2298 750
rect 2220 747 2221 748
rect 2215 746 2221 747
rect 2296 742 2298 748
rect 2303 747 2304 751
rect 2311 747 2312 751
rect 2303 746 2312 747
rect 2367 751 2373 752
rect 2367 747 2368 751
rect 2372 750 2373 751
rect 2391 751 2397 752
rect 2391 750 2392 751
rect 2372 748 2392 750
rect 2372 747 2373 748
rect 2367 746 2373 747
rect 2391 747 2392 748
rect 2396 747 2397 751
rect 2391 746 2397 747
rect 2479 751 2485 752
rect 2479 747 2480 751
rect 2484 750 2485 751
rect 2530 751 2536 752
rect 2530 750 2531 751
rect 2484 748 2531 750
rect 2484 747 2485 748
rect 2479 746 2485 747
rect 2530 747 2531 748
rect 2535 747 2536 751
rect 2530 746 2536 747
rect 2567 751 2573 752
rect 2567 747 2568 751
rect 2572 750 2573 751
rect 2610 751 2616 752
rect 2610 750 2611 751
rect 2572 748 2611 750
rect 2572 747 2573 748
rect 2567 746 2573 747
rect 2610 747 2611 748
rect 2615 747 2616 751
rect 2610 746 2616 747
rect 2671 751 2680 752
rect 2671 747 2672 751
rect 2679 747 2680 751
rect 2671 746 2680 747
rect 2775 751 2781 752
rect 2775 747 2776 751
rect 2780 750 2781 751
rect 2799 751 2805 752
rect 2799 750 2800 751
rect 2780 748 2800 750
rect 2780 747 2781 748
rect 2775 746 2781 747
rect 2799 747 2800 748
rect 2804 747 2805 751
rect 2799 746 2805 747
rect 2927 751 2933 752
rect 2927 747 2928 751
rect 2932 750 2933 751
rect 2951 751 2957 752
rect 2951 750 2952 751
rect 2932 748 2952 750
rect 2932 747 2933 748
rect 2927 746 2933 747
rect 2951 747 2952 748
rect 2956 747 2957 751
rect 2951 746 2957 747
rect 3103 751 3109 752
rect 3103 747 3104 751
rect 3108 750 3109 751
rect 3127 751 3133 752
rect 3127 750 3128 751
rect 3108 748 3128 750
rect 3108 747 3109 748
rect 3103 746 3109 747
rect 3127 747 3128 748
rect 3132 747 3133 751
rect 3127 746 3133 747
rect 3287 751 3293 752
rect 3287 747 3288 751
rect 3292 750 3293 751
rect 3311 751 3317 752
rect 3311 750 3312 751
rect 3292 748 3312 750
rect 3292 747 3293 748
rect 3287 746 3293 747
rect 3311 747 3312 748
rect 3316 747 3317 751
rect 3311 746 3317 747
rect 3495 751 3504 752
rect 3495 747 3496 751
rect 3503 747 3504 751
rect 3495 746 3504 747
rect 2354 743 2360 744
rect 2354 742 2355 743
rect 2296 740 2355 742
rect 2354 739 2355 740
rect 2359 739 2360 743
rect 2354 738 2360 739
rect 367 735 376 736
rect 367 731 368 735
rect 375 731 376 735
rect 367 730 376 731
rect 423 735 429 736
rect 423 731 424 735
rect 428 734 429 735
rect 455 735 461 736
rect 455 734 456 735
rect 428 732 456 734
rect 428 731 429 732
rect 423 730 429 731
rect 455 731 456 732
rect 460 731 461 735
rect 455 730 461 731
rect 511 735 517 736
rect 511 731 512 735
rect 516 734 517 735
rect 551 735 557 736
rect 551 734 552 735
rect 516 732 552 734
rect 516 731 517 732
rect 511 730 517 731
rect 551 731 552 732
rect 556 731 557 735
rect 551 730 557 731
rect 607 735 613 736
rect 607 731 608 735
rect 612 734 613 735
rect 647 735 653 736
rect 647 734 648 735
rect 612 732 648 734
rect 612 731 613 732
rect 607 730 613 731
rect 647 731 648 732
rect 652 731 653 735
rect 647 730 653 731
rect 703 735 709 736
rect 703 731 704 735
rect 708 734 709 735
rect 743 735 749 736
rect 743 734 744 735
rect 708 732 744 734
rect 708 731 709 732
rect 703 730 709 731
rect 743 731 744 732
rect 748 731 749 735
rect 743 730 749 731
rect 839 735 845 736
rect 839 731 840 735
rect 844 734 845 735
rect 895 735 901 736
rect 844 732 890 734
rect 844 731 845 732
rect 839 730 845 731
rect 888 726 890 732
rect 895 731 896 735
rect 900 734 901 735
rect 935 735 941 736
rect 935 734 936 735
rect 900 732 936 734
rect 900 731 901 732
rect 895 730 901 731
rect 935 731 936 732
rect 940 731 941 735
rect 935 730 941 731
rect 991 735 997 736
rect 991 731 992 735
rect 996 734 997 735
rect 1039 735 1045 736
rect 1039 734 1040 735
rect 996 732 1040 734
rect 996 731 997 732
rect 991 730 997 731
rect 1039 731 1040 732
rect 1044 731 1045 735
rect 1039 730 1045 731
rect 1095 735 1101 736
rect 1095 731 1096 735
rect 1100 734 1101 735
rect 1143 735 1149 736
rect 1143 734 1144 735
rect 1100 732 1144 734
rect 1100 731 1101 732
rect 1095 730 1101 731
rect 1143 731 1144 732
rect 1148 731 1149 735
rect 1143 730 1149 731
rect 1223 735 1229 736
rect 1223 731 1224 735
rect 1228 734 1229 735
rect 1247 735 1253 736
rect 1247 734 1248 735
rect 1228 732 1248 734
rect 1228 731 1229 732
rect 1223 730 1229 731
rect 1247 731 1248 732
rect 1252 731 1253 735
rect 1247 730 1253 731
rect 1951 735 1957 736
rect 1951 731 1952 735
rect 1956 734 1957 735
rect 2046 735 2052 736
rect 2046 734 2047 735
rect 1956 732 2047 734
rect 1956 731 1957 732
rect 1951 730 1957 731
rect 2046 731 2047 732
rect 2051 731 2052 735
rect 2046 730 2052 731
rect 2111 735 2120 736
rect 2111 731 2112 735
rect 2119 731 2120 735
rect 2111 730 2120 731
rect 2263 735 2272 736
rect 2263 731 2264 735
rect 2271 731 2272 735
rect 2263 730 2272 731
rect 2335 735 2341 736
rect 2335 731 2336 735
rect 2340 734 2341 735
rect 2415 735 2421 736
rect 2415 734 2416 735
rect 2340 732 2416 734
rect 2340 731 2341 732
rect 2335 730 2341 731
rect 2415 731 2416 732
rect 2420 731 2421 735
rect 2415 730 2421 731
rect 2487 735 2493 736
rect 2487 731 2488 735
rect 2492 734 2493 735
rect 2559 735 2565 736
rect 2559 734 2560 735
rect 2492 732 2560 734
rect 2492 731 2493 732
rect 2487 730 2493 731
rect 2559 731 2560 732
rect 2564 731 2565 735
rect 2559 730 2565 731
rect 2703 735 2712 736
rect 2703 731 2704 735
rect 2711 731 2712 735
rect 2703 730 2712 731
rect 2767 735 2773 736
rect 2767 731 2768 735
rect 2772 734 2773 735
rect 2847 735 2853 736
rect 2847 734 2848 735
rect 2772 732 2848 734
rect 2772 731 2773 732
rect 2767 730 2773 731
rect 2847 731 2848 732
rect 2852 731 2853 735
rect 2847 730 2853 731
rect 2919 735 2925 736
rect 2919 731 2920 735
rect 2924 734 2925 735
rect 2991 735 2997 736
rect 2991 734 2992 735
rect 2924 732 2992 734
rect 2924 731 2925 732
rect 2919 730 2925 731
rect 2991 731 2992 732
rect 2996 731 2997 735
rect 2991 730 2997 731
rect 3063 735 3069 736
rect 3063 731 3064 735
rect 3068 734 3069 735
rect 3143 735 3149 736
rect 3143 734 3144 735
rect 3068 732 3144 734
rect 3068 731 3069 732
rect 3063 730 3069 731
rect 3143 731 3144 732
rect 3148 731 3149 735
rect 3143 730 3149 731
rect 3190 735 3196 736
rect 3190 731 3191 735
rect 3195 734 3196 735
rect 3295 735 3301 736
rect 3295 734 3296 735
rect 3195 732 3296 734
rect 3195 731 3196 732
rect 3190 730 3196 731
rect 3295 731 3296 732
rect 3300 731 3301 735
rect 3295 730 3301 731
rect 3447 735 3456 736
rect 3447 731 3448 735
rect 3455 731 3456 735
rect 3447 730 3456 731
rect 898 727 904 728
rect 898 726 899 727
rect 358 725 364 726
rect 358 721 359 725
rect 363 721 364 725
rect 358 720 364 721
rect 446 725 452 726
rect 446 721 447 725
rect 451 721 452 725
rect 446 720 452 721
rect 542 725 548 726
rect 542 721 543 725
rect 547 721 548 725
rect 542 720 548 721
rect 638 725 644 726
rect 638 721 639 725
rect 643 721 644 725
rect 638 720 644 721
rect 734 725 740 726
rect 734 721 735 725
rect 739 721 740 725
rect 734 720 740 721
rect 830 725 836 726
rect 830 721 831 725
rect 835 721 836 725
rect 888 724 899 726
rect 898 723 899 724
rect 903 723 904 727
rect 898 722 904 723
rect 926 725 932 726
rect 830 720 836 721
rect 926 721 927 725
rect 931 721 932 725
rect 926 720 932 721
rect 1030 725 1036 726
rect 1030 721 1031 725
rect 1035 721 1036 725
rect 1030 720 1036 721
rect 1134 725 1140 726
rect 1134 721 1135 725
rect 1139 721 1140 725
rect 1134 720 1140 721
rect 1238 725 1244 726
rect 1238 721 1239 725
rect 1243 721 1244 725
rect 1238 720 1244 721
rect 1942 725 1948 726
rect 1942 721 1943 725
rect 1947 721 1948 725
rect 1942 720 1948 721
rect 2102 725 2108 726
rect 2102 721 2103 725
rect 2107 721 2108 725
rect 2102 720 2108 721
rect 2254 725 2260 726
rect 2254 721 2255 725
rect 2259 721 2260 725
rect 2254 720 2260 721
rect 2406 725 2412 726
rect 2406 721 2407 725
rect 2411 721 2412 725
rect 2406 720 2412 721
rect 2550 725 2556 726
rect 2550 721 2551 725
rect 2555 721 2556 725
rect 2550 720 2556 721
rect 2694 725 2700 726
rect 2694 721 2695 725
rect 2699 721 2700 725
rect 2694 720 2700 721
rect 2838 725 2844 726
rect 2838 721 2839 725
rect 2843 721 2844 725
rect 2838 720 2844 721
rect 2982 725 2988 726
rect 2982 721 2983 725
rect 2987 721 2988 725
rect 2982 720 2988 721
rect 3134 725 3140 726
rect 3134 721 3135 725
rect 3139 721 3140 725
rect 3134 720 3140 721
rect 3286 725 3292 726
rect 3286 721 3287 725
rect 3291 721 3292 725
rect 3286 720 3292 721
rect 3438 725 3444 726
rect 3438 721 3439 725
rect 3443 721 3444 725
rect 3438 720 3444 721
rect 110 712 116 713
rect 1822 712 1828 713
rect 110 708 111 712
rect 115 708 116 712
rect 423 711 429 712
rect 423 710 424 711
rect 413 708 424 710
rect 110 707 116 708
rect 423 707 424 708
rect 428 707 429 711
rect 511 711 517 712
rect 511 710 512 711
rect 501 708 512 710
rect 423 706 429 707
rect 511 707 512 708
rect 516 707 517 711
rect 607 711 613 712
rect 607 710 608 711
rect 597 708 608 710
rect 511 706 517 707
rect 607 707 608 708
rect 612 707 613 711
rect 703 711 709 712
rect 703 710 704 711
rect 693 708 704 710
rect 607 706 613 707
rect 703 707 704 708
rect 708 707 709 711
rect 895 711 901 712
rect 895 710 896 711
rect 885 708 896 710
rect 703 706 709 707
rect 895 707 896 708
rect 900 707 901 711
rect 991 711 997 712
rect 991 710 992 711
rect 981 708 992 710
rect 895 706 901 707
rect 991 707 992 708
rect 996 707 997 711
rect 1095 711 1101 712
rect 1095 710 1096 711
rect 1085 708 1096 710
rect 991 706 997 707
rect 1095 707 1096 708
rect 1100 707 1101 711
rect 1223 711 1229 712
rect 1223 710 1224 711
rect 1189 708 1224 710
rect 1095 706 1101 707
rect 1223 707 1224 708
rect 1228 707 1229 711
rect 1822 708 1823 712
rect 1827 708 1828 712
rect 1822 707 1828 708
rect 1862 712 1868 713
rect 3574 712 3580 713
rect 1862 708 1863 712
rect 1867 708 1868 712
rect 2335 711 2341 712
rect 2335 710 2336 711
rect 2309 708 2336 710
rect 1862 707 1868 708
rect 2046 707 2052 708
rect 1223 706 1229 707
rect 2046 703 2047 707
rect 2051 706 2052 707
rect 2335 707 2336 708
rect 2340 707 2341 711
rect 2487 711 2493 712
rect 2487 710 2488 711
rect 2461 708 2488 710
rect 2335 706 2341 707
rect 2487 707 2488 708
rect 2492 707 2493 711
rect 2610 711 2616 712
rect 2610 710 2611 711
rect 2605 708 2611 710
rect 2487 706 2493 707
rect 2610 707 2611 708
rect 2615 707 2616 711
rect 2767 711 2773 712
rect 2767 710 2768 711
rect 2749 708 2768 710
rect 2610 706 2616 707
rect 2767 707 2768 708
rect 2772 707 2773 711
rect 2919 711 2925 712
rect 2919 710 2920 711
rect 2893 708 2920 710
rect 2767 706 2773 707
rect 2919 707 2920 708
rect 2924 707 2925 711
rect 3063 711 3069 712
rect 3063 710 3064 711
rect 3037 708 3064 710
rect 2919 706 2925 707
rect 3063 707 3064 708
rect 3068 707 3069 711
rect 3506 711 3512 712
rect 3506 710 3507 711
rect 3493 708 3507 710
rect 3063 706 3069 707
rect 3506 707 3507 708
rect 3511 707 3512 711
rect 3574 708 3575 712
rect 3579 708 3580 712
rect 3574 707 3580 708
rect 3506 706 3512 707
rect 2051 704 2121 706
rect 2051 703 2052 704
rect 2046 702 2052 703
rect 110 695 116 696
rect 110 691 111 695
rect 115 691 116 695
rect 1202 695 1208 696
rect 110 690 116 691
rect 700 692 745 694
rect 350 685 356 686
rect 350 681 351 685
rect 355 681 356 685
rect 350 680 356 681
rect 438 685 444 686
rect 438 681 439 685
rect 443 681 444 685
rect 438 680 444 681
rect 534 685 540 686
rect 534 681 535 685
rect 539 681 540 685
rect 534 680 540 681
rect 630 685 636 686
rect 630 681 631 685
rect 635 681 636 685
rect 630 680 636 681
rect 510 679 516 680
rect 510 675 511 679
rect 515 678 516 679
rect 700 678 702 692
rect 1202 691 1203 695
rect 1207 694 1208 695
rect 1822 695 1828 696
rect 1207 692 1249 694
rect 1207 691 1208 692
rect 1202 690 1208 691
rect 1822 691 1823 695
rect 1827 691 1828 695
rect 1822 690 1828 691
rect 1862 695 1868 696
rect 1862 691 1863 695
rect 1867 691 1868 695
rect 1862 690 1868 691
rect 1906 695 1912 696
rect 1906 691 1907 695
rect 1911 694 1912 695
rect 3078 695 3084 696
rect 1911 692 1953 694
rect 1911 691 1912 692
rect 1906 690 1912 691
rect 3078 691 3079 695
rect 3083 694 3084 695
rect 3226 695 3232 696
rect 3083 692 3145 694
rect 3083 691 3084 692
rect 3078 690 3084 691
rect 3226 691 3227 695
rect 3231 694 3232 695
rect 3574 695 3580 696
rect 3231 692 3297 694
rect 3231 691 3232 692
rect 3226 690 3232 691
rect 3574 691 3575 695
rect 3579 691 3580 695
rect 3574 690 3580 691
rect 726 685 732 686
rect 726 681 727 685
rect 731 681 732 685
rect 726 680 732 681
rect 822 685 828 686
rect 822 681 823 685
rect 827 681 828 685
rect 822 680 828 681
rect 918 685 924 686
rect 918 681 919 685
rect 923 681 924 685
rect 918 680 924 681
rect 1022 685 1028 686
rect 1022 681 1023 685
rect 1027 681 1028 685
rect 1022 680 1028 681
rect 1126 685 1132 686
rect 1126 681 1127 685
rect 1131 681 1132 685
rect 1126 680 1132 681
rect 1230 685 1236 686
rect 1230 681 1231 685
rect 1235 681 1236 685
rect 1230 680 1236 681
rect 1934 685 1940 686
rect 1934 681 1935 685
rect 1939 681 1940 685
rect 1934 680 1940 681
rect 2094 685 2100 686
rect 2094 681 2095 685
rect 2099 681 2100 685
rect 2094 680 2100 681
rect 2246 685 2252 686
rect 2246 681 2247 685
rect 2251 681 2252 685
rect 2246 680 2252 681
rect 2398 685 2404 686
rect 2398 681 2399 685
rect 2403 681 2404 685
rect 2398 680 2404 681
rect 2542 685 2548 686
rect 2542 681 2543 685
rect 2547 681 2548 685
rect 2542 680 2548 681
rect 2686 685 2692 686
rect 2686 681 2687 685
rect 2691 681 2692 685
rect 2686 680 2692 681
rect 2830 685 2836 686
rect 2830 681 2831 685
rect 2835 681 2836 685
rect 2830 680 2836 681
rect 2974 685 2980 686
rect 2974 681 2975 685
rect 2979 681 2980 685
rect 2974 680 2980 681
rect 3126 685 3132 686
rect 3126 681 3127 685
rect 3131 681 3132 685
rect 3126 680 3132 681
rect 3278 685 3284 686
rect 3278 681 3279 685
rect 3283 681 3284 685
rect 3278 680 3284 681
rect 3430 685 3436 686
rect 3430 681 3431 685
rect 3435 681 3436 685
rect 3430 680 3436 681
rect 515 676 702 678
rect 515 675 516 676
rect 510 674 516 675
rect 2114 667 2120 668
rect 2114 663 2115 667
rect 2119 666 2120 667
rect 2119 664 2270 666
rect 2119 663 2120 664
rect 2114 662 2120 663
rect 478 659 484 660
rect 478 655 479 659
rect 483 655 484 659
rect 478 654 484 655
rect 566 659 572 660
rect 566 655 567 659
rect 571 655 572 659
rect 566 654 572 655
rect 654 659 660 660
rect 654 655 655 659
rect 659 655 660 659
rect 654 654 660 655
rect 742 659 748 660
rect 742 655 743 659
rect 747 655 748 659
rect 742 654 748 655
rect 830 659 836 660
rect 830 655 831 659
rect 835 655 836 659
rect 830 654 836 655
rect 918 659 924 660
rect 918 655 919 659
rect 923 655 924 659
rect 918 654 924 655
rect 1006 659 1012 660
rect 1006 655 1007 659
rect 1011 655 1012 659
rect 1006 654 1012 655
rect 1094 659 1100 660
rect 1094 655 1095 659
rect 1099 655 1100 659
rect 1094 654 1100 655
rect 1182 659 1188 660
rect 1182 655 1183 659
rect 1187 655 1188 659
rect 1182 654 1188 655
rect 1270 659 1276 660
rect 1270 655 1271 659
rect 1275 655 1276 659
rect 1270 654 1276 655
rect 1886 659 1892 660
rect 1886 655 1887 659
rect 1891 655 1892 659
rect 1886 654 1892 655
rect 2022 659 2028 660
rect 2022 655 2023 659
rect 2027 655 2028 659
rect 2022 654 2028 655
rect 2198 659 2204 660
rect 2198 655 2199 659
rect 2203 655 2204 659
rect 2198 654 2204 655
rect 898 651 904 652
rect 110 649 116 650
rect 110 645 111 649
rect 115 645 116 649
rect 898 647 899 651
rect 903 650 904 651
rect 2098 651 2104 652
rect 903 648 937 650
rect 1822 649 1828 650
rect 903 647 904 648
rect 898 646 904 647
rect 110 644 116 645
rect 1822 645 1823 649
rect 1827 645 1828 649
rect 1822 644 1828 645
rect 1862 649 1868 650
rect 1862 645 1863 649
rect 1867 645 1868 649
rect 2098 647 2099 651
rect 2103 650 2104 651
rect 2268 650 2270 664
rect 2382 659 2388 660
rect 2382 655 2383 659
rect 2387 655 2388 659
rect 2382 654 2388 655
rect 2566 659 2572 660
rect 2566 655 2567 659
rect 2571 655 2572 659
rect 2566 654 2572 655
rect 2742 659 2748 660
rect 2742 655 2743 659
rect 2747 655 2748 659
rect 2742 654 2748 655
rect 2910 659 2916 660
rect 2910 655 2911 659
rect 2915 655 2916 659
rect 2910 654 2916 655
rect 3062 659 3068 660
rect 3062 655 3063 659
rect 3067 655 3068 659
rect 3062 654 3068 655
rect 3206 659 3212 660
rect 3206 655 3207 659
rect 3211 655 3212 659
rect 3206 654 3212 655
rect 3350 659 3356 660
rect 3350 655 3351 659
rect 3355 655 3356 659
rect 3350 654 3356 655
rect 3478 659 3484 660
rect 3478 655 3479 659
rect 3483 655 3484 659
rect 3478 654 3484 655
rect 3190 651 3196 652
rect 3190 650 3191 651
rect 2103 648 2217 650
rect 2268 648 2401 650
rect 3121 648 3191 650
rect 2103 647 2104 648
rect 2098 646 2104 647
rect 3190 647 3191 648
rect 3195 647 3196 651
rect 3190 646 3196 647
rect 3342 651 3348 652
rect 3342 647 3343 651
rect 3347 650 3348 651
rect 3347 648 3369 650
rect 3574 649 3580 650
rect 3347 647 3348 648
rect 3342 646 3348 647
rect 1862 644 1868 645
rect 3574 645 3575 649
rect 3579 645 3580 649
rect 3574 644 3580 645
rect 559 635 565 636
rect 559 634 560 635
rect 110 632 116 633
rect 541 632 560 634
rect 110 628 111 632
rect 115 628 116 632
rect 559 631 560 632
rect 564 631 565 635
rect 647 635 653 636
rect 647 634 648 635
rect 629 632 648 634
rect 559 630 565 631
rect 647 631 648 632
rect 652 631 653 635
rect 735 635 741 636
rect 735 634 736 635
rect 717 632 736 634
rect 647 630 653 631
rect 735 631 736 632
rect 740 631 741 635
rect 823 635 829 636
rect 823 634 824 635
rect 805 632 824 634
rect 735 630 741 631
rect 823 631 824 632
rect 828 631 829 635
rect 911 635 917 636
rect 911 634 912 635
rect 893 632 912 634
rect 823 630 829 631
rect 911 631 912 632
rect 916 631 917 635
rect 911 630 917 631
rect 986 635 992 636
rect 986 631 987 635
rect 991 634 992 635
rect 1074 635 1080 636
rect 991 632 1033 634
rect 991 631 992 632
rect 986 630 992 631
rect 1074 631 1075 635
rect 1079 634 1080 635
rect 1175 635 1181 636
rect 1079 632 1121 634
rect 1079 631 1080 632
rect 1074 630 1080 631
rect 1175 631 1176 635
rect 1180 634 1181 635
rect 1250 635 1256 636
rect 1180 632 1209 634
rect 1180 631 1181 632
rect 1175 630 1181 631
rect 1250 631 1251 635
rect 1255 634 1256 635
rect 2015 635 2021 636
rect 2015 634 2016 635
rect 1255 632 1297 634
rect 1822 632 1828 633
rect 1255 631 1256 632
rect 1250 630 1256 631
rect 110 627 116 628
rect 1822 628 1823 632
rect 1827 628 1828 632
rect 1822 627 1828 628
rect 1862 632 1868 633
rect 1949 632 2016 634
rect 1862 628 1863 632
rect 1867 628 1868 632
rect 2015 631 2016 632
rect 2020 631 2021 635
rect 2191 635 2197 636
rect 2191 634 2192 635
rect 2085 632 2192 634
rect 2015 630 2021 631
rect 2191 631 2192 632
rect 2196 631 2197 635
rect 2191 630 2197 631
rect 2450 635 2456 636
rect 2450 631 2451 635
rect 2455 634 2456 635
rect 2714 635 2720 636
rect 2455 632 2593 634
rect 2455 631 2456 632
rect 2450 630 2456 631
rect 2714 631 2715 635
rect 2719 634 2720 635
rect 3055 635 3061 636
rect 3055 634 3056 635
rect 2719 632 2769 634
rect 2973 632 3056 634
rect 2719 631 2720 632
rect 2714 630 2720 631
rect 3055 631 3056 632
rect 3060 631 3061 635
rect 3343 635 3349 636
rect 3343 634 3344 635
rect 3269 632 3344 634
rect 3055 630 3061 631
rect 3343 631 3344 632
rect 3348 631 3349 635
rect 3343 630 3349 631
rect 3471 635 3477 636
rect 3471 631 3472 635
rect 3476 634 3477 635
rect 3476 632 3505 634
rect 3574 632 3580 633
rect 3476 631 3477 632
rect 3471 630 3477 631
rect 1862 627 1868 628
rect 3574 628 3575 632
rect 3579 628 3580 632
rect 3574 627 3580 628
rect 486 619 492 620
rect 486 615 487 619
rect 491 615 492 619
rect 486 614 492 615
rect 574 619 580 620
rect 574 615 575 619
rect 579 615 580 619
rect 574 614 580 615
rect 662 619 668 620
rect 662 615 663 619
rect 667 615 668 619
rect 662 614 668 615
rect 750 619 756 620
rect 750 615 751 619
rect 755 615 756 619
rect 750 614 756 615
rect 838 619 844 620
rect 838 615 839 619
rect 843 615 844 619
rect 838 614 844 615
rect 926 619 932 620
rect 926 615 927 619
rect 931 615 932 619
rect 926 614 932 615
rect 1014 619 1020 620
rect 1014 615 1015 619
rect 1019 615 1020 619
rect 1014 614 1020 615
rect 1102 619 1108 620
rect 1102 615 1103 619
rect 1107 615 1108 619
rect 1102 614 1108 615
rect 1190 619 1196 620
rect 1190 615 1191 619
rect 1195 615 1196 619
rect 1190 614 1196 615
rect 1278 619 1284 620
rect 1278 615 1279 619
rect 1283 615 1284 619
rect 1278 614 1284 615
rect 1894 619 1900 620
rect 1894 615 1895 619
rect 1899 615 1900 619
rect 1894 614 1900 615
rect 2030 619 2036 620
rect 2030 615 2031 619
rect 2035 615 2036 619
rect 2030 614 2036 615
rect 2206 619 2212 620
rect 2206 615 2207 619
rect 2211 615 2212 619
rect 2206 614 2212 615
rect 2390 619 2396 620
rect 2390 615 2391 619
rect 2395 615 2396 619
rect 2390 614 2396 615
rect 2574 619 2580 620
rect 2574 615 2575 619
rect 2579 615 2580 619
rect 2574 614 2580 615
rect 2750 619 2756 620
rect 2750 615 2751 619
rect 2755 615 2756 619
rect 2750 614 2756 615
rect 2918 619 2924 620
rect 2918 615 2919 619
rect 2923 615 2924 619
rect 2918 614 2924 615
rect 3070 619 3076 620
rect 3070 615 3071 619
rect 3075 615 3076 619
rect 3070 614 3076 615
rect 3214 619 3220 620
rect 3214 615 3215 619
rect 3219 615 3220 619
rect 3214 614 3220 615
rect 3358 619 3364 620
rect 3358 615 3359 619
rect 3363 615 3364 619
rect 3358 614 3364 615
rect 3486 619 3492 620
rect 3486 615 3487 619
rect 3491 615 3492 619
rect 3486 614 3492 615
rect 495 607 501 608
rect 495 603 496 607
rect 500 606 501 607
rect 510 607 516 608
rect 510 606 511 607
rect 500 604 511 606
rect 500 603 501 604
rect 495 602 501 603
rect 510 603 511 604
rect 515 603 516 607
rect 510 602 516 603
rect 559 607 565 608
rect 559 603 560 607
rect 564 606 565 607
rect 583 607 589 608
rect 583 606 584 607
rect 564 604 584 606
rect 564 603 565 604
rect 559 602 565 603
rect 583 603 584 604
rect 588 603 589 607
rect 583 602 589 603
rect 647 607 653 608
rect 647 603 648 607
rect 652 606 653 607
rect 671 607 677 608
rect 671 606 672 607
rect 652 604 672 606
rect 652 603 653 604
rect 647 602 653 603
rect 671 603 672 604
rect 676 603 677 607
rect 671 602 677 603
rect 735 607 741 608
rect 735 603 736 607
rect 740 606 741 607
rect 759 607 765 608
rect 759 606 760 607
rect 740 604 760 606
rect 740 603 741 604
rect 735 602 741 603
rect 759 603 760 604
rect 764 603 765 607
rect 759 602 765 603
rect 823 607 829 608
rect 823 603 824 607
rect 828 606 829 607
rect 847 607 853 608
rect 847 606 848 607
rect 828 604 848 606
rect 828 603 829 604
rect 823 602 829 603
rect 847 603 848 604
rect 852 603 853 607
rect 847 602 853 603
rect 935 607 941 608
rect 935 603 936 607
rect 940 606 941 607
rect 986 607 992 608
rect 986 606 987 607
rect 940 604 987 606
rect 940 603 941 604
rect 935 602 941 603
rect 986 603 987 604
rect 991 603 992 607
rect 986 602 992 603
rect 1023 607 1029 608
rect 1023 603 1024 607
rect 1028 606 1029 607
rect 1074 607 1080 608
rect 1074 606 1075 607
rect 1028 604 1075 606
rect 1028 603 1029 604
rect 1023 602 1029 603
rect 1074 603 1075 604
rect 1079 603 1080 607
rect 1074 602 1080 603
rect 1111 607 1117 608
rect 1111 603 1112 607
rect 1116 606 1117 607
rect 1175 607 1181 608
rect 1175 606 1176 607
rect 1116 604 1176 606
rect 1116 603 1117 604
rect 1111 602 1117 603
rect 1175 603 1176 604
rect 1180 603 1181 607
rect 1175 602 1181 603
rect 1199 607 1205 608
rect 1199 603 1200 607
rect 1204 606 1205 607
rect 1250 607 1256 608
rect 1250 606 1251 607
rect 1204 604 1251 606
rect 1204 603 1205 604
rect 1199 602 1205 603
rect 1250 603 1251 604
rect 1255 603 1256 607
rect 1250 602 1256 603
rect 1287 607 1293 608
rect 1287 603 1288 607
rect 1292 606 1293 607
rect 1415 607 1421 608
rect 1415 606 1416 607
rect 1292 604 1416 606
rect 1292 603 1293 604
rect 1287 602 1293 603
rect 1415 603 1416 604
rect 1420 603 1421 607
rect 1415 602 1421 603
rect 1903 607 1912 608
rect 1903 603 1904 607
rect 1911 603 1912 607
rect 1903 602 1912 603
rect 2015 607 2021 608
rect 2015 603 2016 607
rect 2020 606 2021 607
rect 2039 607 2045 608
rect 2039 606 2040 607
rect 2020 604 2040 606
rect 2020 603 2021 604
rect 2015 602 2021 603
rect 2039 603 2040 604
rect 2044 603 2045 607
rect 2039 602 2045 603
rect 2191 607 2197 608
rect 2191 603 2192 607
rect 2196 606 2197 607
rect 2215 607 2221 608
rect 2215 606 2216 607
rect 2196 604 2216 606
rect 2196 603 2197 604
rect 2191 602 2197 603
rect 2215 603 2216 604
rect 2220 603 2221 607
rect 2215 602 2221 603
rect 2399 607 2405 608
rect 2399 603 2400 607
rect 2404 606 2405 607
rect 2450 607 2456 608
rect 2450 606 2451 607
rect 2404 604 2451 606
rect 2404 603 2405 604
rect 2399 602 2405 603
rect 2450 603 2451 604
rect 2455 603 2456 607
rect 2450 602 2456 603
rect 2575 607 2581 608
rect 2575 603 2576 607
rect 2580 606 2581 607
rect 2583 607 2589 608
rect 2583 606 2584 607
rect 2580 604 2584 606
rect 2580 603 2581 604
rect 2575 602 2581 603
rect 2583 603 2584 604
rect 2588 603 2589 607
rect 2583 602 2589 603
rect 2759 607 2768 608
rect 2759 603 2760 607
rect 2767 603 2768 607
rect 2759 602 2768 603
rect 2927 607 2933 608
rect 2927 603 2928 607
rect 2932 606 2933 607
rect 2938 607 2944 608
rect 2938 606 2939 607
rect 2932 604 2939 606
rect 2932 603 2933 604
rect 2927 602 2933 603
rect 2938 603 2939 604
rect 2943 603 2944 607
rect 2938 602 2944 603
rect 3055 607 3061 608
rect 3055 603 3056 607
rect 3060 606 3061 607
rect 3079 607 3085 608
rect 3079 606 3080 607
rect 3060 604 3080 606
rect 3060 603 3061 604
rect 3055 602 3061 603
rect 3079 603 3080 604
rect 3084 603 3085 607
rect 3079 602 3085 603
rect 3223 607 3232 608
rect 3223 603 3224 607
rect 3231 603 3232 607
rect 3223 602 3232 603
rect 3343 607 3349 608
rect 3343 603 3344 607
rect 3348 606 3349 607
rect 3367 607 3373 608
rect 3367 606 3368 607
rect 3348 604 3368 606
rect 3348 603 3349 604
rect 3343 602 3349 603
rect 3367 603 3368 604
rect 3372 603 3373 607
rect 3367 602 3373 603
rect 3470 607 3476 608
rect 3470 603 3471 607
rect 3475 606 3476 607
rect 3495 607 3501 608
rect 3495 606 3496 607
rect 3475 604 3496 606
rect 3475 603 3476 604
rect 3470 602 3476 603
rect 3495 603 3496 604
rect 3500 603 3501 607
rect 3495 602 3501 603
rect 3120 600 3218 602
rect 511 595 517 596
rect 511 591 512 595
rect 516 594 517 595
rect 558 595 564 596
rect 558 594 559 595
rect 516 592 559 594
rect 516 591 517 592
rect 511 590 517 591
rect 558 591 559 592
rect 563 591 564 595
rect 558 590 564 591
rect 567 595 573 596
rect 567 591 568 595
rect 572 594 573 595
rect 607 595 613 596
rect 607 594 608 595
rect 572 592 608 594
rect 572 591 573 592
rect 567 590 573 591
rect 607 591 608 592
rect 612 591 613 595
rect 607 590 613 591
rect 663 595 669 596
rect 663 591 664 595
rect 668 594 669 595
rect 711 595 717 596
rect 711 594 712 595
rect 668 592 712 594
rect 668 591 669 592
rect 663 590 669 591
rect 711 591 712 592
rect 716 591 717 595
rect 711 590 717 591
rect 823 595 829 596
rect 823 591 824 595
rect 828 594 829 595
rect 886 595 892 596
rect 886 594 887 595
rect 828 592 887 594
rect 828 591 829 592
rect 823 590 829 591
rect 886 591 887 592
rect 891 591 892 595
rect 886 590 892 591
rect 911 595 917 596
rect 911 591 912 595
rect 916 594 917 595
rect 943 595 949 596
rect 943 594 944 595
rect 916 592 944 594
rect 916 591 917 592
rect 911 590 917 591
rect 943 591 944 592
rect 948 591 949 595
rect 943 590 949 591
rect 1026 595 1032 596
rect 1026 591 1027 595
rect 1031 594 1032 595
rect 1071 595 1077 596
rect 1071 594 1072 595
rect 1031 592 1072 594
rect 1031 591 1032 592
rect 1026 590 1032 591
rect 1071 591 1072 592
rect 1076 591 1077 595
rect 1071 590 1077 591
rect 1127 595 1133 596
rect 1127 591 1128 595
rect 1132 594 1133 595
rect 1199 595 1205 596
rect 1199 594 1200 595
rect 1132 592 1200 594
rect 1132 591 1133 592
rect 1127 590 1133 591
rect 1199 591 1200 592
rect 1204 591 1205 595
rect 1199 590 1205 591
rect 1263 595 1269 596
rect 1263 591 1264 595
rect 1268 594 1269 595
rect 1335 595 1341 596
rect 1335 594 1336 595
rect 1268 592 1336 594
rect 1268 591 1269 592
rect 1263 590 1269 591
rect 1335 591 1336 592
rect 1340 591 1341 595
rect 1335 590 1341 591
rect 1407 595 1413 596
rect 1407 591 1408 595
rect 1412 594 1413 595
rect 1479 595 1485 596
rect 1479 594 1480 595
rect 1412 592 1480 594
rect 1412 591 1413 592
rect 1407 590 1413 591
rect 1479 591 1480 592
rect 1484 591 1485 595
rect 1479 590 1485 591
rect 1623 595 1629 596
rect 1623 591 1624 595
rect 1628 594 1629 595
rect 1686 595 1692 596
rect 1686 594 1687 595
rect 1628 592 1687 594
rect 1628 591 1629 592
rect 1623 590 1629 591
rect 1686 591 1687 592
rect 1691 591 1692 595
rect 1686 590 1692 591
rect 1694 595 1700 596
rect 1694 591 1695 595
rect 1699 594 1700 595
rect 1743 595 1749 596
rect 1743 594 1744 595
rect 1699 592 1744 594
rect 1699 591 1700 592
rect 1694 590 1700 591
rect 1743 591 1744 592
rect 1748 591 1749 595
rect 1743 590 1749 591
rect 1903 595 1909 596
rect 1903 591 1904 595
rect 1908 594 1909 595
rect 1970 595 1976 596
rect 1970 594 1971 595
rect 1908 592 1971 594
rect 1908 591 1909 592
rect 1903 590 1909 591
rect 1970 591 1971 592
rect 1975 591 1976 595
rect 1970 590 1976 591
rect 2095 595 2104 596
rect 2095 591 2096 595
rect 2103 591 2104 595
rect 2095 590 2104 591
rect 2279 595 2285 596
rect 2279 591 2280 595
rect 2284 594 2285 595
rect 2311 595 2317 596
rect 2311 594 2312 595
rect 2284 592 2312 594
rect 2284 591 2285 592
rect 2279 590 2285 591
rect 2311 591 2312 592
rect 2316 591 2317 595
rect 2311 590 2317 591
rect 2415 595 2421 596
rect 2415 591 2416 595
rect 2420 594 2421 595
rect 2519 595 2525 596
rect 2519 594 2520 595
rect 2420 592 2520 594
rect 2420 591 2421 592
rect 2415 590 2421 591
rect 2519 591 2520 592
rect 2524 591 2525 595
rect 2519 590 2525 591
rect 2711 595 2720 596
rect 2711 591 2712 595
rect 2719 591 2720 595
rect 2711 590 2720 591
rect 2775 595 2781 596
rect 2775 591 2776 595
rect 2780 594 2781 595
rect 2887 595 2893 596
rect 2887 594 2888 595
rect 2780 592 2888 594
rect 2780 591 2781 592
rect 2775 590 2781 591
rect 2887 591 2888 592
rect 2892 591 2893 595
rect 2887 590 2893 591
rect 3047 595 3053 596
rect 3047 591 3048 595
rect 3052 594 3053 595
rect 3120 594 3122 600
rect 3216 598 3218 600
rect 3266 599 3272 600
rect 3266 598 3267 599
rect 3216 596 3267 598
rect 3052 592 3122 594
rect 3127 595 3133 596
rect 3052 591 3053 592
rect 3047 590 3053 591
rect 3127 591 3128 595
rect 3132 594 3133 595
rect 3207 595 3213 596
rect 3207 594 3208 595
rect 3132 592 3208 594
rect 3132 591 3133 592
rect 3127 590 3133 591
rect 3207 591 3208 592
rect 3212 591 3213 595
rect 3266 595 3267 596
rect 3271 595 3272 599
rect 3266 594 3272 595
rect 3342 595 3348 596
rect 3207 590 3213 591
rect 3342 591 3343 595
rect 3347 594 3348 595
rect 3359 595 3365 596
rect 3359 594 3360 595
rect 3347 592 3360 594
rect 3347 591 3348 592
rect 3342 590 3348 591
rect 3359 591 3360 592
rect 3364 591 3365 595
rect 3359 590 3365 591
rect 3471 595 3477 596
rect 3471 591 3472 595
rect 3476 594 3477 595
rect 3495 595 3501 596
rect 3495 594 3496 595
rect 3476 592 3496 594
rect 3476 591 3477 592
rect 3471 590 3477 591
rect 3495 591 3496 592
rect 3500 591 3501 595
rect 3495 590 3501 591
rect 502 585 508 586
rect 502 581 503 585
rect 507 581 508 585
rect 502 580 508 581
rect 598 585 604 586
rect 598 581 599 585
rect 603 581 604 585
rect 598 580 604 581
rect 702 585 708 586
rect 702 581 703 585
rect 707 581 708 585
rect 702 580 708 581
rect 814 585 820 586
rect 814 581 815 585
rect 819 581 820 585
rect 814 580 820 581
rect 934 585 940 586
rect 934 581 935 585
rect 939 581 940 585
rect 934 580 940 581
rect 1062 585 1068 586
rect 1062 581 1063 585
rect 1067 581 1068 585
rect 1062 580 1068 581
rect 1190 585 1196 586
rect 1190 581 1191 585
rect 1195 581 1196 585
rect 1190 580 1196 581
rect 1326 585 1332 586
rect 1326 581 1327 585
rect 1331 581 1332 585
rect 1326 580 1332 581
rect 1470 585 1476 586
rect 1470 581 1471 585
rect 1475 581 1476 585
rect 1470 580 1476 581
rect 1614 585 1620 586
rect 1614 581 1615 585
rect 1619 581 1620 585
rect 1614 580 1620 581
rect 1734 585 1740 586
rect 1734 581 1735 585
rect 1739 581 1740 585
rect 1734 580 1740 581
rect 1894 585 1900 586
rect 1894 581 1895 585
rect 1899 581 1900 585
rect 1894 580 1900 581
rect 2086 585 2092 586
rect 2086 581 2087 585
rect 2091 581 2092 585
rect 2086 580 2092 581
rect 2302 585 2308 586
rect 2302 581 2303 585
rect 2307 581 2308 585
rect 2302 580 2308 581
rect 2510 585 2516 586
rect 2510 581 2511 585
rect 2515 581 2516 585
rect 2510 580 2516 581
rect 2702 585 2708 586
rect 2702 581 2703 585
rect 2707 581 2708 585
rect 2702 580 2708 581
rect 2878 585 2884 586
rect 2878 581 2879 585
rect 2883 581 2884 585
rect 2878 580 2884 581
rect 3038 585 3044 586
rect 3038 581 3039 585
rect 3043 581 3044 585
rect 3038 580 3044 581
rect 3198 585 3204 586
rect 3198 581 3199 585
rect 3203 581 3204 585
rect 3198 580 3204 581
rect 3350 585 3356 586
rect 3350 581 3351 585
rect 3355 581 3356 585
rect 3350 580 3356 581
rect 3486 585 3492 586
rect 3486 581 3487 585
rect 3491 581 3492 585
rect 3486 580 3492 581
rect 110 572 116 573
rect 1822 572 1828 573
rect 110 568 111 572
rect 115 568 116 572
rect 567 571 573 572
rect 567 570 568 571
rect 557 568 568 570
rect 110 567 116 568
rect 567 567 568 568
rect 572 567 573 571
rect 663 571 669 572
rect 663 570 664 571
rect 653 568 664 570
rect 567 566 573 567
rect 663 567 664 568
rect 668 567 669 571
rect 1127 571 1133 572
rect 1127 570 1128 571
rect 1117 568 1128 570
rect 663 566 669 567
rect 770 567 776 568
rect 770 563 771 567
rect 775 566 776 567
rect 886 567 892 568
rect 775 564 833 566
rect 775 563 776 564
rect 770 562 776 563
rect 886 563 887 567
rect 891 566 892 567
rect 1127 567 1128 568
rect 1132 567 1133 571
rect 1263 571 1269 572
rect 1263 570 1264 571
rect 1245 568 1264 570
rect 1127 566 1133 567
rect 1263 567 1264 568
rect 1268 567 1269 571
rect 1407 571 1413 572
rect 1407 570 1408 571
rect 1381 568 1408 570
rect 1263 566 1269 567
rect 1407 567 1408 568
rect 1412 567 1413 571
rect 1822 568 1823 572
rect 1827 568 1828 572
rect 1407 566 1413 567
rect 1415 567 1421 568
rect 891 564 953 566
rect 891 563 892 564
rect 886 562 892 563
rect 1415 563 1416 567
rect 1420 566 1421 567
rect 1686 567 1692 568
rect 1822 567 1828 568
rect 1862 572 1868 573
rect 3574 572 3580 573
rect 1862 568 1863 572
rect 1867 568 1868 572
rect 2415 571 2421 572
rect 2415 570 2416 571
rect 2357 568 2416 570
rect 1862 567 1868 568
rect 1970 567 1976 568
rect 1420 564 1489 566
rect 1420 563 1421 564
rect 1415 562 1421 563
rect 1686 563 1687 567
rect 1691 566 1692 567
rect 1691 564 1753 566
rect 1691 563 1692 564
rect 1686 562 1692 563
rect 1970 563 1971 567
rect 1975 566 1976 567
rect 2415 567 2416 568
rect 2420 567 2421 571
rect 2575 571 2581 572
rect 2575 570 2576 571
rect 2565 568 2576 570
rect 2415 566 2421 567
rect 2575 567 2576 568
rect 2580 567 2581 571
rect 2775 571 2781 572
rect 2775 570 2776 571
rect 2757 568 2776 570
rect 2575 566 2581 567
rect 2775 567 2776 568
rect 2780 567 2781 571
rect 2938 571 2944 572
rect 2938 570 2939 571
rect 2933 568 2939 570
rect 2775 566 2781 567
rect 2938 567 2939 568
rect 2943 567 2944 571
rect 3127 571 3133 572
rect 3127 570 3128 571
rect 3093 568 3128 570
rect 2938 566 2944 567
rect 3127 567 3128 568
rect 3132 567 3133 571
rect 3574 568 3575 572
rect 3579 568 3580 572
rect 3127 566 3133 567
rect 3266 567 3272 568
rect 3574 567 3580 568
rect 1975 564 2105 566
rect 1975 563 1976 564
rect 1970 562 1976 563
rect 3266 563 3267 567
rect 3271 566 3272 567
rect 3271 564 3369 566
rect 3271 563 3272 564
rect 3266 562 3272 563
rect 110 555 116 556
rect 110 551 111 555
rect 115 551 116 555
rect 814 555 820 556
rect 814 554 815 555
rect 753 552 815 554
rect 110 550 116 551
rect 814 551 815 552
rect 819 551 820 555
rect 814 550 820 551
rect 1538 555 1544 556
rect 1538 551 1539 555
rect 1543 554 1544 555
rect 1822 555 1828 556
rect 1543 552 1625 554
rect 1543 551 1544 552
rect 1538 550 1544 551
rect 1822 551 1823 555
rect 1827 551 1828 555
rect 1822 550 1828 551
rect 1862 555 1868 556
rect 1862 551 1863 555
rect 1867 551 1868 555
rect 1862 550 1868 551
rect 1870 555 1876 556
rect 1870 551 1871 555
rect 1875 554 1876 555
rect 3350 555 3356 556
rect 3350 554 3351 555
rect 1875 552 1905 554
rect 3249 552 3351 554
rect 1875 551 1876 552
rect 1870 550 1876 551
rect 3350 551 3351 552
rect 3355 551 3356 555
rect 3350 550 3356 551
rect 3574 555 3580 556
rect 3574 551 3575 555
rect 3579 551 3580 555
rect 3574 550 3580 551
rect 494 545 500 546
rect 494 541 495 545
rect 499 541 500 545
rect 494 540 500 541
rect 590 545 596 546
rect 590 541 591 545
rect 595 541 596 545
rect 590 540 596 541
rect 694 545 700 546
rect 694 541 695 545
rect 699 541 700 545
rect 694 540 700 541
rect 806 545 812 546
rect 806 541 807 545
rect 811 541 812 545
rect 806 540 812 541
rect 926 545 932 546
rect 926 541 927 545
rect 931 541 932 545
rect 926 540 932 541
rect 1054 545 1060 546
rect 1054 541 1055 545
rect 1059 541 1060 545
rect 1054 540 1060 541
rect 1182 545 1188 546
rect 1182 541 1183 545
rect 1187 541 1188 545
rect 1182 540 1188 541
rect 1318 545 1324 546
rect 1318 541 1319 545
rect 1323 541 1324 545
rect 1318 540 1324 541
rect 1462 545 1468 546
rect 1462 541 1463 545
rect 1467 541 1468 545
rect 1462 540 1468 541
rect 1606 545 1612 546
rect 1606 541 1607 545
rect 1611 541 1612 545
rect 1606 540 1612 541
rect 1726 545 1732 546
rect 1726 541 1727 545
rect 1731 541 1732 545
rect 1726 540 1732 541
rect 1886 545 1892 546
rect 1886 541 1887 545
rect 1891 541 1892 545
rect 1886 540 1892 541
rect 2078 545 2084 546
rect 2078 541 2079 545
rect 2083 541 2084 545
rect 2078 540 2084 541
rect 2294 545 2300 546
rect 2294 541 2295 545
rect 2299 541 2300 545
rect 2294 540 2300 541
rect 2502 545 2508 546
rect 2502 541 2503 545
rect 2507 541 2508 545
rect 2502 540 2508 541
rect 2694 545 2700 546
rect 2694 541 2695 545
rect 2699 541 2700 545
rect 2694 540 2700 541
rect 2870 545 2876 546
rect 2870 541 2871 545
rect 2875 541 2876 545
rect 2870 540 2876 541
rect 3030 545 3036 546
rect 3030 541 3031 545
rect 3035 541 3036 545
rect 3030 540 3036 541
rect 3190 545 3196 546
rect 3190 541 3191 545
rect 3195 541 3196 545
rect 3190 540 3196 541
rect 3342 545 3348 546
rect 3342 541 3343 545
rect 3347 541 3348 545
rect 3342 540 3348 541
rect 3478 545 3484 546
rect 3478 541 3479 545
rect 3483 541 3484 545
rect 3478 540 3484 541
rect 158 523 164 524
rect 158 519 159 523
rect 163 519 164 523
rect 158 518 164 519
rect 302 523 308 524
rect 302 519 303 523
rect 307 519 308 523
rect 302 518 308 519
rect 462 523 468 524
rect 462 519 463 523
rect 467 519 468 523
rect 462 518 468 519
rect 630 523 636 524
rect 630 519 631 523
rect 635 519 636 523
rect 630 518 636 519
rect 798 523 804 524
rect 798 519 799 523
rect 803 519 804 523
rect 798 518 804 519
rect 958 523 964 524
rect 958 519 959 523
rect 963 519 964 523
rect 958 518 964 519
rect 1102 523 1108 524
rect 1102 519 1103 523
rect 1107 519 1108 523
rect 1102 518 1108 519
rect 1238 523 1244 524
rect 1238 519 1239 523
rect 1243 519 1244 523
rect 1238 518 1244 519
rect 1366 523 1372 524
rect 1366 519 1367 523
rect 1371 519 1372 523
rect 1366 518 1372 519
rect 1494 523 1500 524
rect 1494 519 1495 523
rect 1499 519 1500 523
rect 1494 518 1500 519
rect 1622 523 1628 524
rect 1622 519 1623 523
rect 1627 519 1628 523
rect 1622 518 1628 519
rect 1726 523 1732 524
rect 1726 519 1727 523
rect 1731 519 1732 523
rect 1726 518 1732 519
rect 1026 515 1032 516
rect 1026 514 1027 515
rect 110 513 116 514
rect 110 509 111 513
rect 115 509 116 513
rect 1017 512 1027 514
rect 1026 511 1027 512
rect 1031 511 1032 515
rect 1694 515 1700 516
rect 1694 514 1695 515
rect 1681 512 1695 514
rect 1026 510 1032 511
rect 1694 511 1695 512
rect 1699 511 1700 515
rect 2078 515 2084 516
rect 1694 510 1700 511
rect 1822 513 1828 514
rect 110 508 116 509
rect 1822 509 1823 513
rect 1827 509 1828 513
rect 2078 511 2079 515
rect 2083 511 2084 515
rect 2078 510 2084 511
rect 2286 515 2292 516
rect 2286 511 2287 515
rect 2291 511 2292 515
rect 2286 510 2292 511
rect 2486 515 2492 516
rect 2486 511 2487 515
rect 2491 511 2492 515
rect 2486 510 2492 511
rect 2670 515 2676 516
rect 2670 511 2671 515
rect 2675 511 2676 515
rect 2670 510 2676 511
rect 2846 515 2852 516
rect 2846 511 2847 515
rect 2851 511 2852 515
rect 2846 510 2852 511
rect 3014 515 3020 516
rect 3014 511 3015 515
rect 3019 511 3020 515
rect 3014 510 3020 511
rect 3174 515 3180 516
rect 3174 511 3175 515
rect 3179 511 3180 515
rect 3174 510 3180 511
rect 3334 515 3340 516
rect 3334 511 3335 515
rect 3339 511 3340 515
rect 3334 510 3340 511
rect 3478 515 3484 516
rect 3478 511 3479 515
rect 3483 511 3484 515
rect 3478 510 3484 511
rect 1822 508 1828 509
rect 2279 507 2285 508
rect 1862 505 1868 506
rect 1862 501 1863 505
rect 1867 501 1868 505
rect 2279 503 2280 507
rect 2284 506 2285 507
rect 3082 507 3088 508
rect 2284 504 2305 506
rect 2284 503 2285 504
rect 2279 502 2285 503
rect 3082 503 3083 507
rect 3087 506 3088 507
rect 3450 507 3456 508
rect 3087 504 3193 506
rect 3087 503 3088 504
rect 3082 502 3088 503
rect 3450 503 3451 507
rect 3455 506 3456 507
rect 3455 504 3497 506
rect 3574 505 3580 506
rect 3455 503 3456 504
rect 3450 502 3456 503
rect 1862 500 1868 501
rect 3574 501 3575 505
rect 3579 501 3580 505
rect 3574 500 3580 501
rect 150 499 156 500
rect 110 496 116 497
rect 110 492 111 496
rect 115 492 116 496
rect 150 495 151 499
rect 155 498 156 499
rect 226 499 232 500
rect 155 496 185 498
rect 155 495 156 496
rect 150 494 156 495
rect 226 495 227 499
rect 231 498 232 499
rect 370 499 376 500
rect 231 496 329 498
rect 231 495 232 496
rect 226 494 232 495
rect 370 495 371 499
rect 375 498 376 499
rect 530 499 536 500
rect 375 496 489 498
rect 375 495 376 496
rect 370 494 376 495
rect 530 495 531 499
rect 535 498 536 499
rect 698 499 704 500
rect 535 496 657 498
rect 535 495 536 496
rect 530 494 536 495
rect 698 495 699 499
rect 703 498 704 499
rect 1026 499 1032 500
rect 703 496 825 498
rect 703 495 704 496
rect 698 494 704 495
rect 1026 495 1027 499
rect 1031 498 1032 499
rect 1359 499 1365 500
rect 1359 498 1360 499
rect 1031 496 1129 498
rect 1301 496 1360 498
rect 1031 495 1032 496
rect 1026 494 1032 495
rect 1359 495 1360 496
rect 1364 495 1365 499
rect 1454 499 1460 500
rect 1454 498 1455 499
rect 1429 496 1455 498
rect 1359 494 1365 495
rect 1454 495 1455 496
rect 1459 495 1460 499
rect 1454 494 1460 495
rect 1462 499 1468 500
rect 1462 495 1463 499
rect 1467 498 1468 499
rect 1695 499 1701 500
rect 1467 496 1521 498
rect 1467 495 1468 496
rect 1462 494 1468 495
rect 1695 495 1696 499
rect 1700 498 1701 499
rect 1700 496 1753 498
rect 1822 496 1828 497
rect 1700 495 1701 496
rect 1695 494 1701 495
rect 110 491 116 492
rect 1822 492 1823 496
rect 1827 492 1828 496
rect 1822 491 1828 492
rect 2279 491 2285 492
rect 2279 490 2280 491
rect 1862 488 1868 489
rect 2141 488 2280 490
rect 1862 484 1863 488
rect 1867 484 1868 488
rect 2279 487 2280 488
rect 2284 487 2285 491
rect 2279 486 2285 487
rect 2418 491 2424 492
rect 2418 487 2419 491
rect 2423 490 2424 491
rect 2839 491 2845 492
rect 2839 490 2840 491
rect 2423 488 2513 490
rect 2733 488 2840 490
rect 2423 487 2424 488
rect 2418 486 2424 487
rect 2839 487 2840 488
rect 2844 487 2845 491
rect 3007 491 3013 492
rect 3007 490 3008 491
rect 2909 488 3008 490
rect 2839 486 2845 487
rect 3007 487 3008 488
rect 3012 487 3013 491
rect 3167 491 3173 492
rect 3167 490 3168 491
rect 3077 488 3168 490
rect 3007 486 3013 487
rect 3167 487 3168 488
rect 3172 487 3173 491
rect 3167 486 3173 487
rect 3242 491 3248 492
rect 3242 487 3243 491
rect 3247 490 3248 491
rect 3247 488 3361 490
rect 3574 488 3580 489
rect 3247 487 3248 488
rect 3242 486 3248 487
rect 166 483 172 484
rect 166 479 167 483
rect 171 479 172 483
rect 166 478 172 479
rect 310 483 316 484
rect 310 479 311 483
rect 315 479 316 483
rect 310 478 316 479
rect 470 483 476 484
rect 470 479 471 483
rect 475 479 476 483
rect 470 478 476 479
rect 638 483 644 484
rect 638 479 639 483
rect 643 479 644 483
rect 638 478 644 479
rect 806 483 812 484
rect 806 479 807 483
rect 811 479 812 483
rect 806 478 812 479
rect 966 483 972 484
rect 966 479 967 483
rect 971 479 972 483
rect 966 478 972 479
rect 1110 483 1116 484
rect 1110 479 1111 483
rect 1115 479 1116 483
rect 1110 478 1116 479
rect 1246 483 1252 484
rect 1246 479 1247 483
rect 1251 479 1252 483
rect 1246 478 1252 479
rect 1374 483 1380 484
rect 1374 479 1375 483
rect 1379 479 1380 483
rect 1374 478 1380 479
rect 1502 483 1508 484
rect 1502 479 1503 483
rect 1507 479 1508 483
rect 1502 478 1508 479
rect 1630 483 1636 484
rect 1630 479 1631 483
rect 1635 479 1636 483
rect 1630 478 1636 479
rect 1734 483 1740 484
rect 1862 483 1868 484
rect 3574 484 3575 488
rect 3579 484 3580 488
rect 3574 483 3580 484
rect 1734 479 1735 483
rect 1739 479 1740 483
rect 1734 478 1740 479
rect 2086 475 2092 476
rect 175 471 181 472
rect 175 467 176 471
rect 180 470 181 471
rect 226 471 232 472
rect 226 470 227 471
rect 180 468 227 470
rect 180 467 181 468
rect 175 466 181 467
rect 226 467 227 468
rect 231 467 232 471
rect 226 466 232 467
rect 319 471 325 472
rect 319 467 320 471
rect 324 470 325 471
rect 370 471 376 472
rect 370 470 371 471
rect 324 468 371 470
rect 324 467 325 468
rect 319 466 325 467
rect 370 467 371 468
rect 375 467 376 471
rect 370 466 376 467
rect 479 471 485 472
rect 479 467 480 471
rect 484 470 485 471
rect 530 471 536 472
rect 530 470 531 471
rect 484 468 531 470
rect 484 467 485 468
rect 479 466 485 467
rect 530 467 531 468
rect 535 467 536 471
rect 530 466 536 467
rect 647 471 653 472
rect 647 467 648 471
rect 652 470 653 471
rect 698 471 704 472
rect 698 470 699 471
rect 652 468 699 470
rect 652 467 653 468
rect 647 466 653 467
rect 698 467 699 468
rect 703 467 704 471
rect 698 466 704 467
rect 814 471 821 472
rect 814 467 815 471
rect 820 467 821 471
rect 814 466 821 467
rect 975 471 981 472
rect 975 467 976 471
rect 980 470 981 471
rect 1026 471 1032 472
rect 1026 470 1027 471
rect 980 468 1027 470
rect 980 467 981 468
rect 975 466 981 467
rect 1026 467 1027 468
rect 1031 467 1032 471
rect 1026 466 1032 467
rect 1119 471 1125 472
rect 1119 467 1120 471
rect 1124 470 1125 471
rect 1238 471 1244 472
rect 1238 470 1239 471
rect 1124 468 1239 470
rect 1124 467 1125 468
rect 1119 466 1125 467
rect 1238 467 1239 468
rect 1243 467 1244 471
rect 1238 466 1244 467
rect 1255 471 1261 472
rect 1255 467 1256 471
rect 1260 470 1261 471
rect 1359 471 1365 472
rect 1260 468 1355 470
rect 1260 467 1261 468
rect 1255 466 1261 467
rect 1353 462 1355 468
rect 1359 467 1360 471
rect 1364 470 1365 471
rect 1383 471 1389 472
rect 1383 470 1384 471
rect 1364 468 1384 470
rect 1364 467 1365 468
rect 1359 466 1365 467
rect 1383 467 1384 468
rect 1388 467 1389 471
rect 1383 466 1389 467
rect 1511 471 1517 472
rect 1511 467 1512 471
rect 1516 470 1517 471
rect 1538 471 1544 472
rect 1538 470 1539 471
rect 1516 468 1539 470
rect 1516 467 1517 468
rect 1511 466 1517 467
rect 1538 467 1539 468
rect 1543 467 1544 471
rect 1538 466 1544 467
rect 1639 471 1645 472
rect 1639 467 1640 471
rect 1644 470 1645 471
rect 1695 471 1701 472
rect 1695 470 1696 471
rect 1644 468 1696 470
rect 1644 467 1645 468
rect 1639 466 1645 467
rect 1695 467 1696 468
rect 1700 467 1701 471
rect 1695 466 1701 467
rect 1743 471 1749 472
rect 1743 467 1744 471
rect 1748 470 1749 471
rect 1870 471 1876 472
rect 1870 470 1871 471
rect 1748 468 1871 470
rect 1748 467 1749 468
rect 1743 466 1749 467
rect 1870 467 1871 468
rect 1875 467 1876 471
rect 2086 471 2087 475
rect 2091 471 2092 475
rect 2086 470 2092 471
rect 2294 475 2300 476
rect 2294 471 2295 475
rect 2299 471 2300 475
rect 2294 470 2300 471
rect 2494 475 2500 476
rect 2494 471 2495 475
rect 2499 471 2500 475
rect 2494 470 2500 471
rect 2678 475 2684 476
rect 2678 471 2679 475
rect 2683 471 2684 475
rect 2678 470 2684 471
rect 2854 475 2860 476
rect 2854 471 2855 475
rect 2859 471 2860 475
rect 2854 470 2860 471
rect 3022 475 3028 476
rect 3022 471 3023 475
rect 3027 471 3028 475
rect 3022 470 3028 471
rect 3182 475 3188 476
rect 3182 471 3183 475
rect 3187 471 3188 475
rect 3182 470 3188 471
rect 3342 475 3348 476
rect 3342 471 3343 475
rect 3347 471 3348 475
rect 3342 470 3348 471
rect 3486 475 3492 476
rect 3486 471 3487 475
rect 3491 471 3492 475
rect 3486 470 3492 471
rect 1870 466 1876 467
rect 1462 463 1468 464
rect 1462 462 1463 463
rect 1353 460 1463 462
rect 1462 459 1463 460
rect 1467 459 1468 463
rect 1462 458 1468 459
rect 2094 463 2101 464
rect 2094 459 2095 463
rect 2100 459 2101 463
rect 2094 458 2101 459
rect 2279 463 2285 464
rect 2279 459 2280 463
rect 2284 462 2285 463
rect 2303 463 2309 464
rect 2303 462 2304 463
rect 2284 460 2304 462
rect 2284 459 2285 460
rect 2279 458 2285 459
rect 2303 459 2304 460
rect 2308 459 2309 463
rect 2303 458 2309 459
rect 2503 463 2512 464
rect 2503 459 2504 463
rect 2511 459 2512 463
rect 2503 458 2512 459
rect 2686 463 2693 464
rect 2686 459 2687 463
rect 2692 459 2693 463
rect 2686 458 2693 459
rect 2839 463 2845 464
rect 2839 459 2840 463
rect 2844 462 2845 463
rect 2863 463 2869 464
rect 2863 462 2864 463
rect 2844 460 2864 462
rect 2844 459 2845 460
rect 2839 458 2845 459
rect 2863 459 2864 460
rect 2868 459 2869 463
rect 2863 458 2869 459
rect 3007 463 3013 464
rect 3007 459 3008 463
rect 3012 462 3013 463
rect 3031 463 3037 464
rect 3031 462 3032 463
rect 3012 460 3032 462
rect 3012 459 3013 460
rect 3007 458 3013 459
rect 3031 459 3032 460
rect 3036 459 3037 463
rect 3031 458 3037 459
rect 3191 463 3197 464
rect 3191 459 3192 463
rect 3196 462 3197 463
rect 3242 463 3248 464
rect 3242 462 3243 463
rect 3196 460 3243 462
rect 3196 459 3197 460
rect 3191 458 3197 459
rect 3242 459 3243 460
rect 3247 459 3248 463
rect 3242 458 3248 459
rect 3350 463 3357 464
rect 3350 459 3351 463
rect 3356 459 3357 463
rect 3350 458 3357 459
rect 3478 463 3484 464
rect 3478 459 3479 463
rect 3483 462 3484 463
rect 3495 463 3501 464
rect 3495 462 3496 463
rect 3483 460 3496 462
rect 3483 459 3484 460
rect 3478 458 3484 459
rect 3495 459 3496 460
rect 3500 459 3501 463
rect 3495 458 3501 459
rect 3160 456 3186 458
rect 150 451 157 452
rect 150 447 151 451
rect 156 447 157 451
rect 150 446 157 447
rect 215 451 221 452
rect 215 447 216 451
rect 220 450 221 451
rect 279 451 285 452
rect 279 450 280 451
rect 220 448 280 450
rect 220 447 221 448
rect 215 446 221 447
rect 279 447 280 448
rect 284 447 285 451
rect 279 446 285 447
rect 382 451 388 452
rect 382 447 383 451
rect 387 450 388 451
rect 447 451 453 452
rect 447 450 448 451
rect 387 448 448 450
rect 387 447 388 448
rect 382 446 388 447
rect 447 447 448 448
rect 452 447 453 451
rect 447 446 453 447
rect 535 451 541 452
rect 535 447 536 451
rect 540 450 541 451
rect 623 451 629 452
rect 623 450 624 451
rect 540 448 624 450
rect 540 447 541 448
rect 535 446 541 447
rect 623 447 624 448
rect 628 447 629 451
rect 623 446 629 447
rect 711 451 717 452
rect 711 447 712 451
rect 716 450 717 451
rect 799 451 805 452
rect 799 450 800 451
rect 716 448 800 450
rect 716 447 717 448
rect 711 446 717 447
rect 799 447 800 448
rect 804 447 805 451
rect 799 446 805 447
rect 943 451 949 452
rect 943 447 944 451
rect 948 450 949 451
rect 975 451 981 452
rect 975 450 976 451
rect 948 448 976 450
rect 948 447 949 448
rect 943 446 949 447
rect 975 447 976 448
rect 980 447 981 451
rect 975 446 981 447
rect 1055 451 1061 452
rect 1055 447 1056 451
rect 1060 450 1061 451
rect 1135 451 1141 452
rect 1135 450 1136 451
rect 1060 448 1136 450
rect 1060 447 1061 448
rect 1055 446 1061 447
rect 1135 447 1136 448
rect 1140 447 1141 451
rect 1135 446 1141 447
rect 1271 451 1277 452
rect 1271 447 1272 451
rect 1276 450 1277 451
rect 1295 451 1301 452
rect 1295 450 1296 451
rect 1276 448 1296 450
rect 1276 447 1277 448
rect 1271 446 1277 447
rect 1295 447 1296 448
rect 1300 447 1301 451
rect 1295 446 1301 447
rect 1454 451 1461 452
rect 1454 447 1455 451
rect 1460 447 1461 451
rect 1454 446 1461 447
rect 1535 451 1541 452
rect 1535 447 1536 451
rect 1540 450 1541 451
rect 1615 451 1621 452
rect 1615 450 1616 451
rect 1540 448 1616 450
rect 1540 447 1541 448
rect 1535 446 1541 447
rect 1615 447 1616 448
rect 1620 447 1621 451
rect 1615 446 1621 447
rect 2255 451 2261 452
rect 2255 447 2256 451
rect 2260 450 2261 451
rect 2311 451 2317 452
rect 2260 448 2306 450
rect 2260 447 2261 448
rect 2255 446 2261 447
rect 2302 447 2308 448
rect 2302 443 2303 447
rect 2307 443 2308 447
rect 2311 447 2312 451
rect 2316 450 2317 451
rect 2343 451 2349 452
rect 2343 450 2344 451
rect 2316 448 2344 450
rect 2316 447 2317 448
rect 2311 446 2317 447
rect 2343 447 2344 448
rect 2348 447 2349 451
rect 2343 446 2349 447
rect 2399 451 2405 452
rect 2399 447 2400 451
rect 2404 450 2405 451
rect 2439 451 2445 452
rect 2439 450 2440 451
rect 2404 448 2440 450
rect 2404 447 2405 448
rect 2399 446 2405 447
rect 2439 447 2440 448
rect 2444 447 2445 451
rect 2439 446 2445 447
rect 2495 451 2501 452
rect 2495 447 2496 451
rect 2500 450 2501 451
rect 2535 451 2541 452
rect 2535 450 2536 451
rect 2500 448 2536 450
rect 2500 447 2501 448
rect 2495 446 2501 447
rect 2535 447 2536 448
rect 2540 447 2541 451
rect 2535 446 2541 447
rect 2578 451 2584 452
rect 2578 447 2579 451
rect 2583 450 2584 451
rect 2631 451 2637 452
rect 2631 450 2632 451
rect 2583 448 2632 450
rect 2583 447 2584 448
rect 2578 446 2584 447
rect 2631 447 2632 448
rect 2636 447 2637 451
rect 2631 446 2637 447
rect 2743 451 2749 452
rect 2743 447 2744 451
rect 2748 450 2749 451
rect 2790 451 2796 452
rect 2790 450 2791 451
rect 2748 448 2791 450
rect 2748 447 2749 448
rect 2743 446 2749 447
rect 2790 447 2791 448
rect 2795 447 2796 451
rect 2790 446 2796 447
rect 2799 451 2805 452
rect 2799 447 2800 451
rect 2804 450 2805 451
rect 2871 451 2877 452
rect 2871 450 2872 451
rect 2804 448 2872 450
rect 2804 447 2805 448
rect 2799 446 2805 447
rect 2871 447 2872 448
rect 2876 447 2877 451
rect 2871 446 2877 447
rect 3015 451 3021 452
rect 3015 447 3016 451
rect 3020 450 3021 451
rect 3160 450 3162 456
rect 3184 454 3186 456
rect 3184 452 3222 454
rect 3020 448 3162 450
rect 3167 451 3173 452
rect 3020 447 3021 448
rect 3015 446 3021 447
rect 3167 447 3168 451
rect 3172 450 3173 451
rect 3175 451 3181 452
rect 3175 450 3176 451
rect 3172 448 3176 450
rect 3172 447 3173 448
rect 3167 446 3173 447
rect 3175 447 3176 448
rect 3180 447 3181 451
rect 3175 446 3181 447
rect 2302 442 2308 443
rect 3220 442 3222 452
rect 3255 451 3261 452
rect 3255 447 3256 451
rect 3260 450 3261 451
rect 3343 451 3349 452
rect 3343 450 3344 451
rect 3260 448 3344 450
rect 3260 447 3261 448
rect 3255 446 3261 447
rect 3343 447 3344 448
rect 3348 447 3349 451
rect 3343 446 3349 447
rect 3471 451 3477 452
rect 3471 447 3472 451
rect 3476 450 3477 451
rect 3495 451 3501 452
rect 3495 450 3496 451
rect 3476 448 3496 450
rect 3476 447 3477 448
rect 3471 446 3477 447
rect 3495 447 3496 448
rect 3500 447 3501 451
rect 3495 446 3501 447
rect 3263 443 3269 444
rect 3263 442 3264 443
rect 142 441 148 442
rect 142 437 143 441
rect 147 437 148 441
rect 142 436 148 437
rect 270 441 276 442
rect 270 437 271 441
rect 275 437 276 441
rect 270 436 276 437
rect 438 441 444 442
rect 438 437 439 441
rect 443 437 444 441
rect 438 436 444 437
rect 614 441 620 442
rect 614 437 615 441
rect 619 437 620 441
rect 614 436 620 437
rect 790 441 796 442
rect 790 437 791 441
rect 795 437 796 441
rect 790 436 796 437
rect 966 441 972 442
rect 966 437 967 441
rect 971 437 972 441
rect 966 436 972 437
rect 1126 441 1132 442
rect 1126 437 1127 441
rect 1131 437 1132 441
rect 1126 436 1132 437
rect 1286 441 1292 442
rect 1286 437 1287 441
rect 1291 437 1292 441
rect 1286 436 1292 437
rect 1446 441 1452 442
rect 1446 437 1447 441
rect 1451 437 1452 441
rect 1446 436 1452 437
rect 1606 441 1612 442
rect 1606 437 1607 441
rect 1611 437 1612 441
rect 1606 436 1612 437
rect 2246 441 2252 442
rect 2246 437 2247 441
rect 2251 437 2252 441
rect 2246 436 2252 437
rect 2334 441 2340 442
rect 2334 437 2335 441
rect 2339 437 2340 441
rect 2334 436 2340 437
rect 2430 441 2436 442
rect 2430 437 2431 441
rect 2435 437 2436 441
rect 2430 436 2436 437
rect 2526 441 2532 442
rect 2526 437 2527 441
rect 2531 437 2532 441
rect 2526 436 2532 437
rect 2622 441 2628 442
rect 2622 437 2623 441
rect 2627 437 2628 441
rect 2622 436 2628 437
rect 2734 441 2740 442
rect 2734 437 2735 441
rect 2739 437 2740 441
rect 2734 436 2740 437
rect 2862 441 2868 442
rect 2862 437 2863 441
rect 2867 437 2868 441
rect 2862 436 2868 437
rect 3006 441 3012 442
rect 3006 437 3007 441
rect 3011 437 3012 441
rect 3006 436 3012 437
rect 3166 441 3172 442
rect 3166 437 3167 441
rect 3171 437 3172 441
rect 3220 440 3264 442
rect 3263 439 3264 440
rect 3268 439 3269 443
rect 3263 438 3269 439
rect 3334 441 3340 442
rect 3166 436 3172 437
rect 3334 437 3335 441
rect 3339 437 3340 441
rect 3334 436 3340 437
rect 3486 441 3492 442
rect 3486 437 3487 441
rect 3491 437 3492 441
rect 3486 436 3492 437
rect 110 428 116 429
rect 1822 428 1828 429
rect 110 424 111 428
rect 115 424 116 428
rect 215 427 221 428
rect 215 426 216 427
rect 197 424 216 426
rect 110 423 116 424
rect 215 423 216 424
rect 220 423 221 427
rect 382 427 388 428
rect 382 426 383 427
rect 325 424 383 426
rect 215 422 221 423
rect 382 423 383 424
rect 387 423 388 427
rect 535 427 541 428
rect 535 426 536 427
rect 493 424 536 426
rect 382 422 388 423
rect 535 423 536 424
rect 540 423 541 427
rect 711 427 717 428
rect 711 426 712 427
rect 669 424 712 426
rect 535 422 541 423
rect 711 423 712 424
rect 716 423 717 427
rect 1055 427 1061 428
rect 1055 426 1056 427
rect 1021 424 1056 426
rect 711 422 717 423
rect 1055 423 1056 424
rect 1060 423 1061 427
rect 1271 427 1277 428
rect 1271 426 1272 427
rect 1181 424 1272 426
rect 1055 422 1061 423
rect 1271 423 1272 424
rect 1276 423 1277 427
rect 1535 427 1541 428
rect 1535 426 1536 427
rect 1501 424 1536 426
rect 1271 422 1277 423
rect 1535 423 1536 424
rect 1540 423 1541 427
rect 1822 424 1823 428
rect 1827 424 1828 428
rect 1535 422 1541 423
rect 1546 423 1552 424
rect 1822 423 1828 424
rect 1862 428 1868 429
rect 3574 428 3580 429
rect 1862 424 1863 428
rect 1867 424 1868 428
rect 2311 427 2317 428
rect 2311 426 2312 427
rect 2301 424 2312 426
rect 1862 423 1868 424
rect 2311 423 2312 424
rect 2316 423 2317 427
rect 2399 427 2405 428
rect 2399 426 2400 427
rect 2389 424 2400 426
rect 1546 419 1547 423
rect 1551 422 1552 423
rect 2311 422 2317 423
rect 2399 423 2400 424
rect 2404 423 2405 427
rect 2495 427 2501 428
rect 2495 426 2496 427
rect 2485 424 2496 426
rect 2399 422 2405 423
rect 2495 423 2496 424
rect 2500 423 2501 427
rect 2799 427 2805 428
rect 2799 426 2800 427
rect 2789 424 2800 426
rect 2495 422 2501 423
rect 2506 423 2512 424
rect 1551 420 1625 422
rect 1551 419 1552 420
rect 1546 418 1552 419
rect 2506 419 2507 423
rect 2511 422 2512 423
rect 2594 423 2600 424
rect 2511 420 2545 422
rect 2511 419 2512 420
rect 2506 418 2512 419
rect 2594 419 2595 423
rect 2599 422 2600 423
rect 2799 423 2800 424
rect 2804 423 2805 427
rect 3255 427 3261 428
rect 3255 426 3256 427
rect 3221 424 3256 426
rect 2799 422 2805 423
rect 3255 423 3256 424
rect 3260 423 3261 427
rect 3574 424 3575 428
rect 3579 424 3580 428
rect 3255 422 3261 423
rect 3263 423 3269 424
rect 2599 420 2641 422
rect 2599 419 2600 420
rect 2594 418 2600 419
rect 3263 419 3264 423
rect 3268 422 3269 423
rect 3478 423 3484 424
rect 3574 423 3580 424
rect 3268 420 3353 422
rect 3268 419 3269 420
rect 3263 418 3269 419
rect 3478 419 3479 423
rect 3483 422 3484 423
rect 3483 420 3505 422
rect 3483 419 3484 420
rect 3478 418 3484 419
rect 110 411 116 412
rect 110 407 111 411
rect 115 407 116 411
rect 110 406 116 407
rect 682 411 688 412
rect 682 407 683 411
rect 687 410 688 411
rect 1286 411 1292 412
rect 687 408 801 410
rect 687 407 688 408
rect 682 406 688 407
rect 1286 407 1287 411
rect 1291 410 1292 411
rect 1822 411 1828 412
rect 1291 408 1297 410
rect 1291 407 1292 408
rect 1286 406 1292 407
rect 1822 407 1823 411
rect 1827 407 1828 411
rect 1822 406 1828 407
rect 1862 411 1868 412
rect 1862 407 1863 411
rect 1867 407 1868 411
rect 2934 411 2940 412
rect 2934 410 2935 411
rect 2913 408 2935 410
rect 1862 406 1868 407
rect 2934 407 2935 408
rect 2939 407 2940 411
rect 3574 411 3580 412
rect 2934 406 2940 407
rect 2944 408 3017 410
rect 134 401 140 402
rect 134 397 135 401
rect 139 397 140 401
rect 134 396 140 397
rect 262 401 268 402
rect 262 397 263 401
rect 267 397 268 401
rect 262 396 268 397
rect 430 401 436 402
rect 430 397 431 401
rect 435 397 436 401
rect 430 396 436 397
rect 606 401 612 402
rect 606 397 607 401
rect 611 397 612 401
rect 606 396 612 397
rect 782 401 788 402
rect 782 397 783 401
rect 787 397 788 401
rect 782 396 788 397
rect 958 401 964 402
rect 958 397 959 401
rect 963 397 964 401
rect 958 396 964 397
rect 1118 401 1124 402
rect 1118 397 1119 401
rect 1123 397 1124 401
rect 1118 396 1124 397
rect 1278 401 1284 402
rect 1278 397 1279 401
rect 1283 397 1284 401
rect 1278 396 1284 397
rect 1438 401 1444 402
rect 1438 397 1439 401
rect 1443 397 1444 401
rect 1438 396 1444 397
rect 1598 401 1604 402
rect 1598 397 1599 401
rect 1603 397 1604 401
rect 1598 396 1604 397
rect 2238 401 2244 402
rect 2238 397 2239 401
rect 2243 397 2244 401
rect 2238 396 2244 397
rect 2326 401 2332 402
rect 2326 397 2327 401
rect 2331 397 2332 401
rect 2326 396 2332 397
rect 2422 401 2428 402
rect 2422 397 2423 401
rect 2427 397 2428 401
rect 2422 396 2428 397
rect 2518 401 2524 402
rect 2518 397 2519 401
rect 2523 397 2524 401
rect 2518 396 2524 397
rect 2614 401 2620 402
rect 2614 397 2615 401
rect 2619 397 2620 401
rect 2614 396 2620 397
rect 2726 401 2732 402
rect 2726 397 2727 401
rect 2731 397 2732 401
rect 2726 396 2732 397
rect 2854 401 2860 402
rect 2854 397 2855 401
rect 2859 397 2860 401
rect 2854 396 2860 397
rect 2790 395 2796 396
rect 2790 391 2791 395
rect 2795 394 2796 395
rect 2944 394 2946 408
rect 3574 407 3575 411
rect 3579 407 3580 411
rect 3574 406 3580 407
rect 2998 401 3004 402
rect 2998 397 2999 401
rect 3003 397 3004 401
rect 2998 396 3004 397
rect 3158 401 3164 402
rect 3158 397 3159 401
rect 3163 397 3164 401
rect 3158 396 3164 397
rect 3326 401 3332 402
rect 3326 397 3327 401
rect 3331 397 3332 401
rect 3326 396 3332 397
rect 3478 401 3484 402
rect 3478 397 3479 401
rect 3483 397 3484 401
rect 3478 396 3484 397
rect 2795 392 2946 394
rect 2795 391 2796 392
rect 2790 390 2796 391
rect 134 379 140 380
rect 134 375 135 379
rect 139 375 140 379
rect 134 374 140 375
rect 262 379 268 380
rect 262 375 263 379
rect 267 375 268 379
rect 262 374 268 375
rect 430 379 436 380
rect 430 375 431 379
rect 435 375 436 379
rect 430 374 436 375
rect 606 379 612 380
rect 606 375 607 379
rect 611 375 612 379
rect 606 374 612 375
rect 782 379 788 380
rect 782 375 783 379
rect 787 375 788 379
rect 782 374 788 375
rect 950 379 956 380
rect 950 375 951 379
rect 955 375 956 379
rect 950 374 956 375
rect 1110 379 1116 380
rect 1110 375 1111 379
rect 1115 375 1116 379
rect 1110 374 1116 375
rect 1270 379 1276 380
rect 1270 375 1271 379
rect 1275 375 1276 379
rect 1270 374 1276 375
rect 1430 379 1436 380
rect 1430 375 1431 379
rect 1435 375 1436 379
rect 1430 374 1436 375
rect 1590 379 1596 380
rect 1590 375 1591 379
rect 1595 375 1596 379
rect 1590 374 1596 375
rect 2150 379 2156 380
rect 2150 375 2151 379
rect 2155 375 2156 379
rect 2150 374 2156 375
rect 2238 379 2244 380
rect 2238 375 2239 379
rect 2243 375 2244 379
rect 2238 374 2244 375
rect 2326 379 2332 380
rect 2326 375 2327 379
rect 2331 375 2332 379
rect 2326 374 2332 375
rect 2414 379 2420 380
rect 2414 375 2415 379
rect 2419 375 2420 379
rect 2414 374 2420 375
rect 2502 379 2508 380
rect 2502 375 2503 379
rect 2507 375 2508 379
rect 2502 374 2508 375
rect 2614 379 2620 380
rect 2614 375 2615 379
rect 2619 375 2620 379
rect 2614 374 2620 375
rect 2750 379 2756 380
rect 2750 375 2751 379
rect 2755 375 2756 379
rect 2750 374 2756 375
rect 2918 379 2924 380
rect 2918 375 2919 379
rect 2923 375 2924 379
rect 2918 374 2924 375
rect 3102 379 3108 380
rect 3102 375 3103 379
rect 3107 375 3108 379
rect 3102 374 3108 375
rect 3302 379 3308 380
rect 3302 375 3303 379
rect 3307 375 3308 379
rect 3302 374 3308 375
rect 3478 379 3484 380
rect 3478 375 3479 379
rect 3483 375 3484 379
rect 3478 374 3484 375
rect 690 371 696 372
rect 110 369 116 370
rect 110 365 111 369
rect 115 365 116 369
rect 690 367 691 371
rect 695 370 696 371
rect 943 371 949 372
rect 695 368 801 370
rect 695 367 696 368
rect 690 366 696 367
rect 943 367 944 371
rect 948 370 949 371
rect 2578 371 2584 372
rect 2578 370 2579 371
rect 948 368 969 370
rect 1822 369 1828 370
rect 948 367 949 368
rect 943 366 949 367
rect 110 364 116 365
rect 1822 365 1823 369
rect 1827 365 1828 369
rect 1822 364 1828 365
rect 1862 369 1868 370
rect 1862 365 1863 369
rect 1867 365 1868 369
rect 2561 368 2579 370
rect 2578 367 2579 368
rect 2583 367 2584 371
rect 2578 366 2584 367
rect 3198 371 3204 372
rect 3198 367 3199 371
rect 3203 370 3204 371
rect 3471 371 3477 372
rect 3203 368 3321 370
rect 3203 367 3204 368
rect 3198 366 3204 367
rect 3471 367 3472 371
rect 3476 370 3477 371
rect 3476 368 3497 370
rect 3574 369 3580 370
rect 3476 367 3477 368
rect 3471 366 3477 367
rect 1862 364 1868 365
rect 3574 365 3575 369
rect 3579 365 3580 369
rect 3574 364 3580 365
rect 255 355 261 356
rect 255 354 256 355
rect 110 352 116 353
rect 197 352 256 354
rect 110 348 111 352
rect 115 348 116 352
rect 255 351 256 352
rect 260 351 261 355
rect 423 355 429 356
rect 423 354 424 355
rect 325 352 424 354
rect 255 350 261 351
rect 423 351 424 352
rect 428 351 429 355
rect 599 355 605 356
rect 599 354 600 355
rect 493 352 600 354
rect 423 350 429 351
rect 599 351 600 352
rect 604 351 605 355
rect 775 355 781 356
rect 775 354 776 355
rect 669 352 776 354
rect 599 350 605 351
rect 775 351 776 352
rect 780 351 781 355
rect 775 350 781 351
rect 1018 355 1024 356
rect 1018 351 1019 355
rect 1023 354 1024 355
rect 1423 355 1429 356
rect 1423 354 1424 355
rect 1023 352 1137 354
rect 1333 352 1424 354
rect 1023 351 1024 352
rect 1018 350 1024 351
rect 1423 351 1424 352
rect 1428 351 1429 355
rect 1583 355 1589 356
rect 1583 354 1584 355
rect 1493 352 1584 354
rect 1423 350 1429 351
rect 1583 351 1584 352
rect 1588 351 1589 355
rect 1694 355 1700 356
rect 1694 354 1695 355
rect 1653 352 1695 354
rect 1583 350 1589 351
rect 1694 351 1695 352
rect 1699 351 1700 355
rect 2231 355 2237 356
rect 2231 354 2232 355
rect 1694 350 1700 351
rect 1822 352 1828 353
rect 110 347 116 348
rect 1822 348 1823 352
rect 1827 348 1828 352
rect 1822 347 1828 348
rect 1862 352 1868 353
rect 2213 352 2232 354
rect 1862 348 1863 352
rect 1867 348 1868 352
rect 2231 351 2232 352
rect 2236 351 2237 355
rect 2319 355 2325 356
rect 2319 354 2320 355
rect 2301 352 2320 354
rect 2231 350 2237 351
rect 2319 351 2320 352
rect 2324 351 2325 355
rect 2407 355 2413 356
rect 2407 354 2408 355
rect 2389 352 2408 354
rect 2319 350 2325 351
rect 2407 351 2408 352
rect 2412 351 2413 355
rect 2495 355 2501 356
rect 2495 354 2496 355
rect 2477 352 2496 354
rect 2407 350 2413 351
rect 2495 351 2496 352
rect 2500 351 2501 355
rect 2495 350 2501 351
rect 2570 355 2576 356
rect 2570 351 2571 355
rect 2575 354 2576 355
rect 2682 355 2688 356
rect 2575 352 2641 354
rect 2575 351 2576 352
rect 2570 350 2576 351
rect 2682 351 2683 355
rect 2687 354 2688 355
rect 3095 355 3101 356
rect 3095 354 3096 355
rect 2687 352 2777 354
rect 2981 352 3096 354
rect 2687 351 2688 352
rect 2682 350 2688 351
rect 3095 351 3096 352
rect 3100 351 3101 355
rect 3295 355 3301 356
rect 3295 354 3296 355
rect 3165 352 3296 354
rect 3095 350 3101 351
rect 3295 351 3296 352
rect 3300 351 3301 355
rect 3295 350 3301 351
rect 3574 352 3580 353
rect 1862 347 1868 348
rect 3574 348 3575 352
rect 3579 348 3580 352
rect 3574 347 3580 348
rect 142 339 148 340
rect 142 335 143 339
rect 147 335 148 339
rect 142 334 148 335
rect 270 339 276 340
rect 270 335 271 339
rect 275 335 276 339
rect 270 334 276 335
rect 438 339 444 340
rect 438 335 439 339
rect 443 335 444 339
rect 438 334 444 335
rect 614 339 620 340
rect 614 335 615 339
rect 619 335 620 339
rect 614 334 620 335
rect 790 339 796 340
rect 790 335 791 339
rect 795 335 796 339
rect 790 334 796 335
rect 958 339 964 340
rect 958 335 959 339
rect 963 335 964 339
rect 958 334 964 335
rect 1118 339 1124 340
rect 1118 335 1119 339
rect 1123 335 1124 339
rect 1118 334 1124 335
rect 1278 339 1284 340
rect 1278 335 1279 339
rect 1283 335 1284 339
rect 1278 334 1284 335
rect 1438 339 1444 340
rect 1438 335 1439 339
rect 1443 335 1444 339
rect 1438 334 1444 335
rect 1598 339 1604 340
rect 1598 335 1599 339
rect 1603 335 1604 339
rect 1598 334 1604 335
rect 2158 339 2164 340
rect 2158 335 2159 339
rect 2163 335 2164 339
rect 2158 334 2164 335
rect 2246 339 2252 340
rect 2246 335 2247 339
rect 2251 335 2252 339
rect 2246 334 2252 335
rect 2334 339 2340 340
rect 2334 335 2335 339
rect 2339 335 2340 339
rect 2334 334 2340 335
rect 2422 339 2428 340
rect 2422 335 2423 339
rect 2427 335 2428 339
rect 2422 334 2428 335
rect 2510 339 2516 340
rect 2510 335 2511 339
rect 2515 335 2516 339
rect 2510 334 2516 335
rect 2622 339 2628 340
rect 2622 335 2623 339
rect 2627 335 2628 339
rect 2622 334 2628 335
rect 2758 339 2764 340
rect 2758 335 2759 339
rect 2763 335 2764 339
rect 2758 334 2764 335
rect 2926 339 2932 340
rect 2926 335 2927 339
rect 2931 335 2932 339
rect 2926 334 2932 335
rect 3110 339 3116 340
rect 3110 335 3111 339
rect 3115 335 3116 339
rect 3110 334 3116 335
rect 3310 339 3316 340
rect 3310 335 3311 339
rect 3315 335 3316 339
rect 3310 334 3316 335
rect 3486 339 3492 340
rect 3486 335 3487 339
rect 3491 335 3492 339
rect 3486 334 3492 335
rect 151 327 160 328
rect 151 323 152 327
rect 159 323 160 327
rect 151 322 160 323
rect 255 327 261 328
rect 255 323 256 327
rect 260 326 261 327
rect 279 327 285 328
rect 279 326 280 327
rect 260 324 280 326
rect 260 323 261 324
rect 255 322 261 323
rect 279 323 280 324
rect 284 323 285 327
rect 279 322 285 323
rect 423 327 429 328
rect 423 323 424 327
rect 428 326 429 327
rect 447 327 453 328
rect 447 326 448 327
rect 428 324 448 326
rect 428 323 429 324
rect 423 322 429 323
rect 447 323 448 324
rect 452 323 453 327
rect 447 322 453 323
rect 599 327 605 328
rect 599 323 600 327
rect 604 326 605 327
rect 623 327 629 328
rect 623 326 624 327
rect 604 324 624 326
rect 604 323 605 324
rect 599 322 605 323
rect 623 323 624 324
rect 628 323 629 327
rect 623 322 629 323
rect 775 327 781 328
rect 775 323 776 327
rect 780 326 781 327
rect 799 327 805 328
rect 799 326 800 327
rect 780 324 800 326
rect 780 323 781 324
rect 775 322 781 323
rect 799 323 800 324
rect 804 323 805 327
rect 799 322 805 323
rect 967 327 973 328
rect 967 323 968 327
rect 972 326 973 327
rect 1018 327 1024 328
rect 1018 326 1019 327
rect 972 324 1019 326
rect 972 323 973 324
rect 967 322 973 323
rect 1018 323 1019 324
rect 1023 323 1024 327
rect 1018 322 1024 323
rect 1127 327 1133 328
rect 1127 323 1128 327
rect 1132 326 1133 327
rect 1242 327 1248 328
rect 1242 326 1243 327
rect 1132 324 1243 326
rect 1132 323 1133 324
rect 1127 322 1133 323
rect 1242 323 1243 324
rect 1247 323 1248 327
rect 1242 322 1248 323
rect 1286 327 1293 328
rect 1286 323 1287 327
rect 1292 323 1293 327
rect 1286 322 1293 323
rect 1423 327 1429 328
rect 1423 323 1424 327
rect 1428 326 1429 327
rect 1447 327 1453 328
rect 1447 326 1448 327
rect 1428 324 1448 326
rect 1428 323 1429 324
rect 1423 322 1429 323
rect 1447 323 1448 324
rect 1452 323 1453 327
rect 1447 322 1453 323
rect 1583 327 1589 328
rect 1583 323 1584 327
rect 1588 326 1589 327
rect 1607 327 1613 328
rect 1607 326 1608 327
rect 1588 324 1608 326
rect 1588 323 1589 324
rect 1583 322 1589 323
rect 1607 323 1608 324
rect 1612 323 1613 327
rect 1607 322 1613 323
rect 2167 327 2173 328
rect 2167 323 2168 327
rect 2172 326 2173 327
rect 2214 327 2220 328
rect 2214 326 2215 327
rect 2172 324 2215 326
rect 2172 323 2173 324
rect 2167 322 2173 323
rect 2214 323 2215 324
rect 2219 323 2220 327
rect 2214 322 2220 323
rect 2231 327 2237 328
rect 2231 323 2232 327
rect 2236 326 2237 327
rect 2255 327 2261 328
rect 2255 326 2256 327
rect 2236 324 2256 326
rect 2236 323 2237 324
rect 2231 322 2237 323
rect 2255 323 2256 324
rect 2260 323 2261 327
rect 2255 322 2261 323
rect 2319 327 2325 328
rect 2319 323 2320 327
rect 2324 326 2325 327
rect 2343 327 2349 328
rect 2343 326 2344 327
rect 2324 324 2344 326
rect 2324 323 2325 324
rect 2319 322 2325 323
rect 2343 323 2344 324
rect 2348 323 2349 327
rect 2343 322 2349 323
rect 2407 327 2413 328
rect 2407 323 2408 327
rect 2412 326 2413 327
rect 2431 327 2437 328
rect 2431 326 2432 327
rect 2412 324 2432 326
rect 2412 323 2413 324
rect 2407 322 2413 323
rect 2431 323 2432 324
rect 2436 323 2437 327
rect 2431 322 2437 323
rect 2495 327 2501 328
rect 2495 323 2496 327
rect 2500 326 2501 327
rect 2519 327 2525 328
rect 2519 326 2520 327
rect 2500 324 2520 326
rect 2500 323 2501 324
rect 2495 322 2501 323
rect 2519 323 2520 324
rect 2524 323 2525 327
rect 2519 322 2525 323
rect 2631 327 2637 328
rect 2631 323 2632 327
rect 2636 326 2637 327
rect 2682 327 2688 328
rect 2682 326 2683 327
rect 2636 324 2683 326
rect 2636 323 2637 324
rect 2631 322 2637 323
rect 2682 323 2683 324
rect 2687 323 2688 327
rect 2682 322 2688 323
rect 2767 327 2776 328
rect 2767 323 2768 327
rect 2775 323 2776 327
rect 2767 322 2776 323
rect 2934 327 2941 328
rect 2934 323 2935 327
rect 2940 323 2941 327
rect 2934 322 2941 323
rect 3095 327 3101 328
rect 3095 323 3096 327
rect 3100 326 3101 327
rect 3119 327 3125 328
rect 3119 326 3120 327
rect 3100 324 3120 326
rect 3100 323 3101 324
rect 3095 322 3101 323
rect 3119 323 3120 324
rect 3124 323 3125 327
rect 3119 322 3125 323
rect 3295 327 3301 328
rect 3295 323 3296 327
rect 3300 326 3301 327
rect 3319 327 3325 328
rect 3319 326 3320 327
rect 3300 324 3320 326
rect 3300 323 3301 324
rect 3295 322 3301 323
rect 3319 323 3320 324
rect 3324 323 3325 327
rect 3319 322 3325 323
rect 3471 327 3477 328
rect 3471 323 3472 327
rect 3476 326 3477 327
rect 3495 327 3501 328
rect 3495 326 3496 327
rect 3476 324 3496 326
rect 3476 323 3477 324
rect 3471 322 3477 323
rect 3495 323 3496 324
rect 3500 323 3501 327
rect 3495 322 3501 323
rect 350 315 356 316
rect 350 314 351 315
rect 272 312 351 314
rect 271 311 277 312
rect 271 307 272 311
rect 276 307 277 311
rect 350 311 351 312
rect 355 311 356 315
rect 2030 315 2037 316
rect 350 310 356 311
rect 358 311 364 312
rect 271 306 277 307
rect 358 307 359 311
rect 363 310 364 311
rect 399 311 405 312
rect 399 310 400 311
rect 363 308 400 310
rect 363 307 364 308
rect 358 306 364 307
rect 399 307 400 308
rect 404 307 405 311
rect 399 306 405 307
rect 463 311 469 312
rect 463 307 464 311
rect 468 310 469 311
rect 535 311 541 312
rect 535 310 536 311
rect 468 308 536 310
rect 468 307 469 308
rect 463 306 469 307
rect 535 307 536 308
rect 540 307 541 311
rect 535 306 541 307
rect 607 311 613 312
rect 607 307 608 311
rect 612 310 613 311
rect 687 311 693 312
rect 687 310 688 311
rect 612 308 688 310
rect 612 307 613 308
rect 607 306 613 307
rect 687 307 688 308
rect 692 307 693 311
rect 687 306 693 307
rect 767 311 773 312
rect 767 307 768 311
rect 772 310 773 311
rect 847 311 853 312
rect 847 310 848 311
rect 772 308 848 310
rect 772 307 773 308
rect 767 306 773 307
rect 847 307 848 308
rect 852 307 853 311
rect 847 306 853 307
rect 983 311 989 312
rect 983 307 984 311
rect 988 310 989 311
rect 1015 311 1021 312
rect 1015 310 1016 311
rect 988 308 1016 310
rect 988 307 989 308
rect 983 306 989 307
rect 1015 307 1016 308
rect 1020 307 1021 311
rect 1015 306 1021 307
rect 1087 311 1093 312
rect 1087 307 1088 311
rect 1092 310 1093 311
rect 1183 311 1189 312
rect 1183 310 1184 311
rect 1092 308 1184 310
rect 1092 307 1093 308
rect 1087 306 1093 307
rect 1183 307 1184 308
rect 1188 307 1189 311
rect 1183 306 1189 307
rect 1234 311 1240 312
rect 1234 307 1235 311
rect 1239 310 1240 311
rect 1351 311 1357 312
rect 1351 310 1352 311
rect 1239 308 1352 310
rect 1239 307 1240 308
rect 1234 306 1240 307
rect 1351 307 1352 308
rect 1356 307 1357 311
rect 1351 306 1357 307
rect 1519 311 1525 312
rect 1519 307 1520 311
rect 1524 310 1525 311
rect 1607 311 1613 312
rect 1607 310 1608 311
rect 1524 308 1608 310
rect 1524 307 1525 308
rect 1519 306 1525 307
rect 1607 307 1608 308
rect 1612 307 1613 311
rect 1607 306 1613 307
rect 1694 311 1701 312
rect 1694 307 1695 311
rect 1700 307 1701 311
rect 2030 311 2031 315
rect 2036 311 2037 315
rect 2030 310 2037 311
rect 2087 315 2093 316
rect 2087 311 2088 315
rect 2092 314 2093 315
rect 2127 315 2133 316
rect 2127 314 2128 315
rect 2092 312 2128 314
rect 2092 311 2093 312
rect 2087 310 2093 311
rect 2127 311 2128 312
rect 2132 311 2133 315
rect 2127 310 2133 311
rect 2183 315 2189 316
rect 2183 311 2184 315
rect 2188 314 2189 315
rect 2231 315 2237 316
rect 2231 314 2232 315
rect 2188 312 2232 314
rect 2188 311 2189 312
rect 2183 310 2189 311
rect 2231 311 2232 312
rect 2236 311 2237 315
rect 2231 310 2237 311
rect 2287 315 2293 316
rect 2287 311 2288 315
rect 2292 314 2293 315
rect 2335 315 2341 316
rect 2335 314 2336 315
rect 2292 312 2336 314
rect 2292 311 2293 312
rect 2287 310 2293 311
rect 2335 311 2336 312
rect 2340 311 2341 315
rect 2335 310 2341 311
rect 2390 315 2396 316
rect 2390 311 2391 315
rect 2395 314 2396 315
rect 2439 315 2445 316
rect 2439 314 2440 315
rect 2395 312 2440 314
rect 2395 311 2396 312
rect 2390 310 2396 311
rect 2439 311 2440 312
rect 2444 311 2445 315
rect 2439 310 2445 311
rect 2543 315 2549 316
rect 2543 311 2544 315
rect 2548 314 2549 315
rect 2570 315 2576 316
rect 2570 314 2571 315
rect 2548 312 2571 314
rect 2548 311 2549 312
rect 2543 310 2549 311
rect 2570 311 2571 312
rect 2575 311 2576 315
rect 2570 310 2576 311
rect 2599 315 2605 316
rect 2599 311 2600 315
rect 2604 314 2605 315
rect 2647 315 2653 316
rect 2647 314 2648 315
rect 2604 312 2648 314
rect 2604 311 2605 312
rect 2599 310 2605 311
rect 2647 311 2648 312
rect 2652 311 2653 315
rect 2647 310 2653 311
rect 2703 315 2709 316
rect 2703 311 2704 315
rect 2708 314 2709 315
rect 2751 315 2757 316
rect 2751 314 2752 315
rect 2708 312 2752 314
rect 2708 311 2709 312
rect 2703 310 2709 311
rect 2751 311 2752 312
rect 2756 311 2757 315
rect 2751 310 2757 311
rect 2807 315 2813 316
rect 2807 311 2808 315
rect 2812 314 2813 315
rect 2863 315 2869 316
rect 2863 314 2864 315
rect 2812 312 2864 314
rect 2812 311 2813 312
rect 2807 310 2813 311
rect 2863 311 2864 312
rect 2868 311 2869 315
rect 2863 310 2869 311
rect 2919 315 2925 316
rect 2919 311 2920 315
rect 2924 314 2925 315
rect 2975 315 2981 316
rect 2975 314 2976 315
rect 2924 312 2976 314
rect 2924 311 2925 312
rect 2919 310 2925 311
rect 2975 311 2976 312
rect 2980 311 2981 315
rect 2975 310 2981 311
rect 1694 306 1701 307
rect 2022 305 2028 306
rect 262 301 268 302
rect 262 297 263 301
rect 267 297 268 301
rect 262 296 268 297
rect 390 301 396 302
rect 390 297 391 301
rect 395 297 396 301
rect 390 296 396 297
rect 526 301 532 302
rect 526 297 527 301
rect 531 297 532 301
rect 526 296 532 297
rect 678 301 684 302
rect 678 297 679 301
rect 683 297 684 301
rect 678 296 684 297
rect 838 301 844 302
rect 838 297 839 301
rect 843 297 844 301
rect 838 296 844 297
rect 1006 301 1012 302
rect 1006 297 1007 301
rect 1011 297 1012 301
rect 1006 296 1012 297
rect 1174 301 1180 302
rect 1174 297 1175 301
rect 1179 297 1180 301
rect 1174 296 1180 297
rect 1342 301 1348 302
rect 1342 297 1343 301
rect 1347 297 1348 301
rect 1342 296 1348 297
rect 1510 301 1516 302
rect 1510 297 1511 301
rect 1515 297 1516 301
rect 1510 296 1516 297
rect 1686 301 1692 302
rect 1686 297 1687 301
rect 1691 297 1692 301
rect 2022 301 2023 305
rect 2027 301 2028 305
rect 2022 300 2028 301
rect 2118 305 2124 306
rect 2118 301 2119 305
rect 2123 301 2124 305
rect 2118 300 2124 301
rect 2222 305 2228 306
rect 2222 301 2223 305
rect 2227 301 2228 305
rect 2222 300 2228 301
rect 2326 305 2332 306
rect 2326 301 2327 305
rect 2331 301 2332 305
rect 2326 300 2332 301
rect 2430 305 2436 306
rect 2430 301 2431 305
rect 2435 301 2436 305
rect 2430 300 2436 301
rect 2534 305 2540 306
rect 2534 301 2535 305
rect 2539 301 2540 305
rect 2534 300 2540 301
rect 2638 305 2644 306
rect 2638 301 2639 305
rect 2643 301 2644 305
rect 2638 300 2644 301
rect 2742 305 2748 306
rect 2742 301 2743 305
rect 2747 301 2748 305
rect 2742 300 2748 301
rect 2854 305 2860 306
rect 2854 301 2855 305
rect 2859 301 2860 305
rect 2854 300 2860 301
rect 2966 305 2972 306
rect 2966 301 2967 305
rect 2971 301 2972 305
rect 2966 300 2972 301
rect 1686 296 1692 297
rect 1862 292 1868 293
rect 3574 292 3580 293
rect 110 288 116 289
rect 1822 288 1828 289
rect 110 284 111 288
rect 115 284 116 288
rect 358 287 364 288
rect 358 286 359 287
rect 317 284 359 286
rect 110 283 116 284
rect 358 283 359 284
rect 363 283 364 287
rect 463 287 469 288
rect 463 286 464 287
rect 445 284 464 286
rect 358 282 364 283
rect 463 283 464 284
rect 468 283 469 287
rect 607 287 613 288
rect 607 286 608 287
rect 581 284 608 286
rect 463 282 469 283
rect 607 283 608 284
rect 612 283 613 287
rect 767 287 773 288
rect 767 286 768 287
rect 733 284 768 286
rect 607 282 613 283
rect 767 283 768 284
rect 772 283 773 287
rect 1087 287 1093 288
rect 1087 286 1088 287
rect 1061 284 1088 286
rect 767 282 773 283
rect 1087 283 1088 284
rect 1092 283 1093 287
rect 1234 287 1240 288
rect 1234 286 1235 287
rect 1229 284 1235 286
rect 1087 282 1093 283
rect 1234 283 1235 284
rect 1239 283 1240 287
rect 1822 284 1823 288
rect 1827 284 1828 288
rect 1862 288 1863 292
rect 1867 288 1868 292
rect 2087 291 2093 292
rect 2087 290 2088 291
rect 2077 288 2088 290
rect 1862 287 1868 288
rect 2087 287 2088 288
rect 2092 287 2093 291
rect 2183 291 2189 292
rect 2183 290 2184 291
rect 2173 288 2184 290
rect 2087 286 2093 287
rect 2183 287 2184 288
rect 2188 287 2189 291
rect 2287 291 2293 292
rect 2287 290 2288 291
rect 2277 288 2288 290
rect 2183 286 2189 287
rect 2287 287 2288 288
rect 2292 287 2293 291
rect 2390 291 2396 292
rect 2390 290 2391 291
rect 2381 288 2391 290
rect 2287 286 2293 287
rect 2390 287 2391 288
rect 2395 287 2396 291
rect 2599 291 2605 292
rect 2599 290 2600 291
rect 2589 288 2600 290
rect 2390 286 2396 287
rect 2398 287 2404 288
rect 1234 282 1240 283
rect 1242 283 1248 284
rect 1242 279 1243 283
rect 1247 282 1248 283
rect 1607 283 1613 284
rect 1822 283 1828 284
rect 2398 283 2399 287
rect 2403 286 2404 287
rect 2599 287 2600 288
rect 2604 287 2605 291
rect 2703 291 2709 292
rect 2703 290 2704 291
rect 2693 288 2704 290
rect 2599 286 2605 287
rect 2703 287 2704 288
rect 2708 287 2709 291
rect 2807 291 2813 292
rect 2807 290 2808 291
rect 2797 288 2808 290
rect 2703 286 2709 287
rect 2807 287 2808 288
rect 2812 287 2813 291
rect 2919 291 2925 292
rect 2919 290 2920 291
rect 2909 288 2920 290
rect 2807 286 2813 287
rect 2919 287 2920 288
rect 2924 287 2925 291
rect 3574 288 3575 292
rect 3579 288 3580 292
rect 3574 287 3580 288
rect 2919 286 2925 287
rect 2403 284 2449 286
rect 2403 283 2404 284
rect 1247 280 1361 282
rect 1247 279 1248 280
rect 1242 278 1248 279
rect 1607 279 1608 283
rect 1612 282 1613 283
rect 2398 282 2404 283
rect 1612 280 1705 282
rect 1612 279 1613 280
rect 1607 278 1613 279
rect 1862 275 1868 276
rect 110 271 116 272
rect 110 267 111 271
rect 115 267 116 271
rect 110 266 116 267
rect 810 271 816 272
rect 810 267 811 271
rect 815 270 816 271
rect 1410 271 1416 272
rect 815 268 849 270
rect 815 267 816 268
rect 810 266 816 267
rect 1410 267 1411 271
rect 1415 270 1416 271
rect 1822 271 1828 272
rect 1415 268 1521 270
rect 1415 267 1416 268
rect 1410 266 1416 267
rect 1822 267 1823 271
rect 1827 267 1828 271
rect 1862 271 1863 275
rect 1867 271 1868 275
rect 1862 270 1868 271
rect 2922 275 2928 276
rect 2922 271 2923 275
rect 2927 274 2928 275
rect 3574 275 3580 276
rect 2927 272 2977 274
rect 2927 271 2928 272
rect 2922 270 2928 271
rect 3574 271 3575 275
rect 3579 271 3580 275
rect 3574 270 3580 271
rect 1822 266 1828 267
rect 2014 265 2020 266
rect 254 261 260 262
rect 254 257 255 261
rect 259 257 260 261
rect 254 256 260 257
rect 382 261 388 262
rect 382 257 383 261
rect 387 257 388 261
rect 382 256 388 257
rect 518 261 524 262
rect 518 257 519 261
rect 523 257 524 261
rect 518 256 524 257
rect 670 261 676 262
rect 670 257 671 261
rect 675 257 676 261
rect 670 256 676 257
rect 830 261 836 262
rect 830 257 831 261
rect 835 257 836 261
rect 830 256 836 257
rect 998 261 1004 262
rect 998 257 999 261
rect 1003 257 1004 261
rect 998 256 1004 257
rect 1166 261 1172 262
rect 1166 257 1167 261
rect 1171 257 1172 261
rect 1166 256 1172 257
rect 1334 261 1340 262
rect 1334 257 1335 261
rect 1339 257 1340 261
rect 1334 256 1340 257
rect 1502 261 1508 262
rect 1502 257 1503 261
rect 1507 257 1508 261
rect 1502 256 1508 257
rect 1678 261 1684 262
rect 1678 257 1679 261
rect 1683 257 1684 261
rect 2014 261 2015 265
rect 2019 261 2020 265
rect 2014 260 2020 261
rect 2110 265 2116 266
rect 2110 261 2111 265
rect 2115 261 2116 265
rect 2110 260 2116 261
rect 2214 265 2220 266
rect 2214 261 2215 265
rect 2219 261 2220 265
rect 2214 260 2220 261
rect 2318 265 2324 266
rect 2318 261 2319 265
rect 2323 261 2324 265
rect 2318 260 2324 261
rect 2422 265 2428 266
rect 2422 261 2423 265
rect 2427 261 2428 265
rect 2422 260 2428 261
rect 2526 265 2532 266
rect 2526 261 2527 265
rect 2531 261 2532 265
rect 2526 260 2532 261
rect 2630 265 2636 266
rect 2630 261 2631 265
rect 2635 261 2636 265
rect 2630 260 2636 261
rect 2734 265 2740 266
rect 2734 261 2735 265
rect 2739 261 2740 265
rect 2734 260 2740 261
rect 2846 265 2852 266
rect 2846 261 2847 265
rect 2851 261 2852 265
rect 2846 260 2852 261
rect 2958 265 2964 266
rect 2958 261 2959 265
rect 2963 261 2964 265
rect 2958 260 2964 261
rect 1678 256 1684 257
rect 1958 243 1964 244
rect 1958 239 1959 243
rect 1963 239 1964 243
rect 1958 238 1964 239
rect 2174 243 2180 244
rect 2174 239 2175 243
rect 2179 239 2180 243
rect 2174 238 2180 239
rect 2382 243 2388 244
rect 2382 239 2383 243
rect 2387 239 2388 243
rect 2382 238 2388 239
rect 2582 243 2588 244
rect 2582 239 2583 243
rect 2587 239 2588 243
rect 2582 238 2588 239
rect 2766 243 2772 244
rect 2766 239 2767 243
rect 2771 239 2772 243
rect 2766 238 2772 239
rect 2950 243 2956 244
rect 2950 239 2951 243
rect 2955 239 2956 243
rect 2950 238 2956 239
rect 3126 243 3132 244
rect 3126 239 3127 243
rect 3131 239 3132 243
rect 3126 238 3132 239
rect 3310 243 3316 244
rect 3310 239 3311 243
rect 3315 239 3316 243
rect 3310 238 3316 239
rect 3478 243 3484 244
rect 3478 239 3479 243
rect 3483 239 3484 243
rect 3478 238 3484 239
rect 398 235 404 236
rect 398 231 399 235
rect 403 231 404 235
rect 398 230 404 231
rect 502 235 508 236
rect 502 231 503 235
rect 507 231 508 235
rect 502 230 508 231
rect 614 235 620 236
rect 614 231 615 235
rect 619 231 620 235
rect 614 230 620 231
rect 734 235 740 236
rect 734 231 735 235
rect 739 231 740 235
rect 734 230 740 231
rect 862 235 868 236
rect 862 231 863 235
rect 867 231 868 235
rect 862 230 868 231
rect 990 235 996 236
rect 990 231 991 235
rect 995 231 996 235
rect 990 230 996 231
rect 1118 235 1124 236
rect 1118 231 1119 235
rect 1123 231 1124 235
rect 1118 230 1124 231
rect 1246 235 1252 236
rect 1246 231 1247 235
rect 1251 231 1252 235
rect 1246 230 1252 231
rect 1374 235 1380 236
rect 1374 231 1375 235
rect 1379 231 1380 235
rect 1374 230 1380 231
rect 1494 235 1500 236
rect 1494 231 1495 235
rect 1499 231 1500 235
rect 1494 230 1500 231
rect 1622 235 1628 236
rect 1622 231 1623 235
rect 1627 231 1628 235
rect 1622 230 1628 231
rect 1726 235 1732 236
rect 1726 231 1727 235
rect 1731 231 1732 235
rect 2030 235 2036 236
rect 2030 234 2031 235
rect 1726 230 1732 231
rect 1862 233 1868 234
rect 1862 229 1863 233
rect 1867 229 1868 233
rect 2017 232 2031 234
rect 2030 231 2031 232
rect 2035 231 2036 235
rect 2030 230 2036 231
rect 3198 235 3204 236
rect 3198 231 3199 235
rect 3203 234 3204 235
rect 3471 235 3477 236
rect 3203 232 3329 234
rect 3203 231 3204 232
rect 3198 230 3204 231
rect 3471 231 3472 235
rect 3476 234 3477 235
rect 3476 232 3497 234
rect 3574 233 3580 234
rect 3476 231 3477 232
rect 3471 230 3477 231
rect 1862 228 1868 229
rect 3574 229 3575 233
rect 3579 229 3580 233
rect 3574 228 3580 229
rect 802 227 808 228
rect 110 225 116 226
rect 110 221 111 225
rect 115 221 116 225
rect 802 223 803 227
rect 807 226 808 227
rect 983 227 989 228
rect 807 224 881 226
rect 807 223 808 224
rect 802 222 808 223
rect 983 223 984 227
rect 988 226 989 227
rect 988 224 1009 226
rect 1728 224 1745 226
rect 1822 225 1828 226
rect 988 223 989 224
rect 983 222 989 223
rect 1726 223 1732 224
rect 110 220 116 221
rect 1726 219 1727 223
rect 1731 219 1732 223
rect 1822 221 1823 225
rect 1827 221 1828 225
rect 1822 220 1828 221
rect 1726 218 1732 219
rect 2094 219 2100 220
rect 1862 216 1868 217
rect 1862 212 1863 216
rect 1867 212 1868 216
rect 2094 215 2095 219
rect 2099 218 2100 219
rect 2242 219 2248 220
rect 2099 216 2201 218
rect 2099 215 2100 216
rect 2094 214 2100 215
rect 2242 215 2243 219
rect 2247 218 2248 219
rect 2759 219 2765 220
rect 2759 218 2760 219
rect 2247 216 2409 218
rect 2645 216 2760 218
rect 2247 215 2248 216
rect 2242 214 2248 215
rect 2759 215 2760 216
rect 2764 215 2765 219
rect 2943 219 2949 220
rect 2943 218 2944 219
rect 2829 216 2944 218
rect 2759 214 2765 215
rect 2943 215 2944 216
rect 2948 215 2949 219
rect 3119 219 3125 220
rect 3119 218 3120 219
rect 3013 216 3120 218
rect 2943 214 2949 215
rect 3119 215 3120 216
rect 3124 215 3125 219
rect 3303 219 3309 220
rect 3303 218 3304 219
rect 3189 216 3304 218
rect 3119 214 3125 215
rect 3303 215 3304 216
rect 3308 215 3309 219
rect 3303 214 3309 215
rect 3574 216 3580 217
rect 495 211 501 212
rect 495 210 496 211
rect 110 208 116 209
rect 461 208 496 210
rect 110 204 111 208
rect 115 204 116 208
rect 495 207 496 208
rect 500 207 501 211
rect 607 211 613 212
rect 607 210 608 211
rect 565 208 608 210
rect 495 206 501 207
rect 607 207 608 208
rect 612 207 613 211
rect 727 211 733 212
rect 727 210 728 211
rect 677 208 728 210
rect 607 206 613 207
rect 727 207 728 208
rect 732 207 733 211
rect 855 211 861 212
rect 855 210 856 211
rect 797 208 856 210
rect 727 206 733 207
rect 855 207 856 208
rect 860 207 861 211
rect 855 206 861 207
rect 1058 211 1064 212
rect 1058 207 1059 211
rect 1063 210 1064 211
rect 1214 211 1220 212
rect 1063 208 1145 210
rect 1063 207 1064 208
rect 1058 206 1064 207
rect 1214 207 1215 211
rect 1219 210 1220 211
rect 1487 211 1493 212
rect 1487 210 1488 211
rect 1219 208 1273 210
rect 1437 208 1488 210
rect 1219 207 1220 208
rect 1214 206 1220 207
rect 1487 207 1488 208
rect 1492 207 1493 211
rect 1615 211 1621 212
rect 1615 210 1616 211
rect 1557 208 1616 210
rect 1487 206 1493 207
rect 1615 207 1616 208
rect 1620 207 1621 211
rect 1719 211 1725 212
rect 1862 211 1868 212
rect 3574 212 3575 216
rect 3579 212 3580 216
rect 3574 211 3580 212
rect 1719 210 1720 211
rect 1685 208 1720 210
rect 1615 206 1621 207
rect 1719 207 1720 208
rect 1724 207 1725 211
rect 1719 206 1725 207
rect 1822 208 1828 209
rect 110 203 116 204
rect 1822 204 1823 208
rect 1827 204 1828 208
rect 1822 203 1828 204
rect 1966 203 1972 204
rect 1966 199 1967 203
rect 1971 199 1972 203
rect 1966 198 1972 199
rect 2182 203 2188 204
rect 2182 199 2183 203
rect 2187 199 2188 203
rect 2182 198 2188 199
rect 2390 203 2396 204
rect 2390 199 2391 203
rect 2395 199 2396 203
rect 2390 198 2396 199
rect 2590 203 2596 204
rect 2590 199 2591 203
rect 2595 199 2596 203
rect 2590 198 2596 199
rect 2774 203 2780 204
rect 2774 199 2775 203
rect 2779 199 2780 203
rect 2774 198 2780 199
rect 2958 203 2964 204
rect 2958 199 2959 203
rect 2963 199 2964 203
rect 2958 198 2964 199
rect 3134 203 3140 204
rect 3134 199 3135 203
rect 3139 199 3140 203
rect 3134 198 3140 199
rect 3318 203 3324 204
rect 3318 199 3319 203
rect 3323 199 3324 203
rect 3318 198 3324 199
rect 3486 203 3492 204
rect 3486 199 3487 203
rect 3491 199 3492 203
rect 3486 198 3492 199
rect 406 195 412 196
rect 406 191 407 195
rect 411 191 412 195
rect 406 190 412 191
rect 510 195 516 196
rect 510 191 511 195
rect 515 191 516 195
rect 510 190 516 191
rect 622 195 628 196
rect 622 191 623 195
rect 627 191 628 195
rect 622 190 628 191
rect 742 195 748 196
rect 742 191 743 195
rect 747 191 748 195
rect 742 190 748 191
rect 870 195 876 196
rect 870 191 871 195
rect 875 191 876 195
rect 870 190 876 191
rect 998 195 1004 196
rect 998 191 999 195
rect 1003 191 1004 195
rect 998 190 1004 191
rect 1126 195 1132 196
rect 1126 191 1127 195
rect 1131 191 1132 195
rect 1126 190 1132 191
rect 1254 195 1260 196
rect 1254 191 1255 195
rect 1259 191 1260 195
rect 1254 190 1260 191
rect 1382 195 1388 196
rect 1382 191 1383 195
rect 1387 191 1388 195
rect 1382 190 1388 191
rect 1502 195 1508 196
rect 1502 191 1503 195
rect 1507 191 1508 195
rect 1502 190 1508 191
rect 1630 195 1636 196
rect 1630 191 1631 195
rect 1635 191 1636 195
rect 1630 190 1636 191
rect 1734 195 1740 196
rect 1734 191 1735 195
rect 1739 191 1740 195
rect 1734 190 1740 191
rect 1975 191 1981 192
rect 1975 187 1976 191
rect 1980 190 1981 191
rect 2094 191 2100 192
rect 2094 190 2095 191
rect 1980 188 2095 190
rect 1980 187 1981 188
rect 1975 186 1981 187
rect 2094 187 2095 188
rect 2099 187 2100 191
rect 2094 186 2100 187
rect 2191 191 2197 192
rect 2191 187 2192 191
rect 2196 190 2197 191
rect 2242 191 2248 192
rect 2242 190 2243 191
rect 2196 188 2243 190
rect 2196 187 2197 188
rect 2191 186 2197 187
rect 2242 187 2243 188
rect 2247 187 2248 191
rect 2242 186 2248 187
rect 2399 191 2405 192
rect 2399 187 2400 191
rect 2404 190 2405 191
rect 2450 191 2456 192
rect 2450 190 2451 191
rect 2404 188 2451 190
rect 2404 187 2405 188
rect 2399 186 2405 187
rect 2450 187 2451 188
rect 2455 187 2456 191
rect 2450 186 2456 187
rect 2599 191 2608 192
rect 2599 187 2600 191
rect 2607 187 2608 191
rect 2599 186 2608 187
rect 2759 191 2765 192
rect 2759 187 2760 191
rect 2764 190 2765 191
rect 2783 191 2789 192
rect 2783 190 2784 191
rect 2764 188 2784 190
rect 2764 187 2765 188
rect 2759 186 2765 187
rect 2783 187 2784 188
rect 2788 187 2789 191
rect 2783 186 2789 187
rect 2943 191 2949 192
rect 2943 187 2944 191
rect 2948 190 2949 191
rect 2967 191 2973 192
rect 2967 190 2968 191
rect 2948 188 2968 190
rect 2948 187 2949 188
rect 2943 186 2949 187
rect 2967 187 2968 188
rect 2972 187 2973 191
rect 2967 186 2973 187
rect 3119 191 3125 192
rect 3119 187 3120 191
rect 3124 190 3125 191
rect 3143 191 3149 192
rect 3143 190 3144 191
rect 3124 188 3144 190
rect 3124 187 3125 188
rect 3119 186 3125 187
rect 3143 187 3144 188
rect 3148 187 3149 191
rect 3143 186 3149 187
rect 3303 191 3309 192
rect 3303 187 3304 191
rect 3308 190 3309 191
rect 3327 191 3333 192
rect 3327 190 3328 191
rect 3308 188 3328 190
rect 3308 187 3309 188
rect 3303 186 3309 187
rect 3327 187 3328 188
rect 3332 187 3333 191
rect 3327 186 3333 187
rect 3478 191 3484 192
rect 3478 187 3479 191
rect 3483 190 3484 191
rect 3495 191 3501 192
rect 3495 190 3496 191
rect 3483 188 3496 190
rect 3483 187 3484 188
rect 3478 186 3484 187
rect 3495 187 3496 188
rect 3500 187 3501 191
rect 3495 186 3501 187
rect 415 183 424 184
rect 415 179 416 183
rect 423 179 424 183
rect 415 178 424 179
rect 495 183 501 184
rect 495 179 496 183
rect 500 182 501 183
rect 519 183 525 184
rect 519 182 520 183
rect 500 180 520 182
rect 500 179 501 180
rect 495 178 501 179
rect 519 179 520 180
rect 524 179 525 183
rect 519 178 525 179
rect 607 183 613 184
rect 607 179 608 183
rect 612 182 613 183
rect 631 183 637 184
rect 631 182 632 183
rect 612 180 632 182
rect 612 179 613 180
rect 607 178 613 179
rect 631 179 632 180
rect 636 179 637 183
rect 631 178 637 179
rect 727 183 733 184
rect 727 179 728 183
rect 732 182 733 183
rect 751 183 757 184
rect 751 182 752 183
rect 732 180 752 182
rect 732 179 733 180
rect 727 178 733 179
rect 751 179 752 180
rect 756 179 757 183
rect 751 178 757 179
rect 855 183 861 184
rect 855 179 856 183
rect 860 182 861 183
rect 879 183 885 184
rect 879 182 880 183
rect 860 180 880 182
rect 860 179 861 180
rect 855 178 861 179
rect 879 179 880 180
rect 884 179 885 183
rect 879 178 885 179
rect 1007 183 1013 184
rect 1007 179 1008 183
rect 1012 182 1013 183
rect 1058 183 1064 184
rect 1058 182 1059 183
rect 1012 180 1059 182
rect 1012 179 1013 180
rect 1007 178 1013 179
rect 1058 179 1059 180
rect 1063 179 1064 183
rect 1058 178 1064 179
rect 1135 183 1141 184
rect 1135 179 1136 183
rect 1140 182 1141 183
rect 1214 183 1220 184
rect 1214 182 1215 183
rect 1140 180 1215 182
rect 1140 179 1141 180
rect 1135 178 1141 179
rect 1214 179 1215 180
rect 1219 179 1220 183
rect 1214 178 1220 179
rect 1263 183 1269 184
rect 1263 179 1264 183
rect 1268 182 1269 183
rect 1391 183 1397 184
rect 1268 180 1386 182
rect 1268 179 1269 180
rect 1263 178 1269 179
rect 1384 174 1386 180
rect 1391 179 1392 183
rect 1396 182 1397 183
rect 1410 183 1416 184
rect 1410 182 1411 183
rect 1396 180 1411 182
rect 1396 179 1397 180
rect 1391 178 1397 179
rect 1410 179 1411 180
rect 1415 179 1416 183
rect 1410 178 1416 179
rect 1487 183 1493 184
rect 1487 179 1488 183
rect 1492 182 1493 183
rect 1511 183 1517 184
rect 1511 182 1512 183
rect 1492 180 1512 182
rect 1492 179 1493 180
rect 1487 178 1493 179
rect 1511 179 1512 180
rect 1516 179 1517 183
rect 1511 178 1517 179
rect 1615 183 1621 184
rect 1615 179 1616 183
rect 1620 182 1621 183
rect 1639 183 1645 184
rect 1639 182 1640 183
rect 1620 180 1640 182
rect 1620 179 1621 180
rect 1615 178 1621 179
rect 1639 179 1640 180
rect 1644 179 1645 183
rect 1639 178 1645 179
rect 1719 183 1725 184
rect 1719 179 1720 183
rect 1724 182 1725 183
rect 1743 183 1749 184
rect 1743 182 1744 183
rect 1724 180 1744 182
rect 1724 179 1725 180
rect 1719 178 1725 179
rect 1743 179 1744 180
rect 1748 179 1749 183
rect 1743 178 1749 179
rect 1583 175 1589 176
rect 1583 174 1584 175
rect 1384 172 1584 174
rect 1583 171 1584 172
rect 1588 171 1589 175
rect 1583 170 1589 171
rect 802 159 808 160
rect 802 158 803 159
rect 276 156 803 158
rect 231 151 237 152
rect 231 147 232 151
rect 236 150 237 151
rect 276 150 278 156
rect 802 155 803 156
rect 807 155 808 159
rect 802 154 808 155
rect 236 148 278 150
rect 287 151 293 152
rect 236 147 237 148
rect 231 146 237 147
rect 287 147 288 151
rect 292 150 293 151
rect 319 151 325 152
rect 319 150 320 151
rect 292 148 320 150
rect 292 147 293 148
rect 287 146 293 147
rect 319 147 320 148
rect 324 147 325 151
rect 319 146 325 147
rect 375 151 381 152
rect 375 147 376 151
rect 380 150 381 151
rect 407 151 413 152
rect 407 150 408 151
rect 380 148 408 150
rect 380 147 381 148
rect 375 146 381 147
rect 407 147 408 148
rect 412 147 413 151
rect 407 146 413 147
rect 463 151 469 152
rect 463 147 464 151
rect 468 150 469 151
rect 495 151 501 152
rect 495 150 496 151
rect 468 148 496 150
rect 468 147 469 148
rect 463 146 469 147
rect 495 147 496 148
rect 500 147 501 151
rect 495 146 501 147
rect 551 151 557 152
rect 551 147 552 151
rect 556 150 557 151
rect 583 151 589 152
rect 583 150 584 151
rect 556 148 584 150
rect 556 147 557 148
rect 551 146 557 147
rect 583 147 584 148
rect 588 147 589 151
rect 583 146 589 147
rect 639 151 645 152
rect 639 147 640 151
rect 644 150 645 151
rect 671 151 677 152
rect 671 150 672 151
rect 644 148 672 150
rect 644 147 645 148
rect 639 146 645 147
rect 671 147 672 148
rect 676 147 677 151
rect 671 146 677 147
rect 727 151 733 152
rect 727 147 728 151
rect 732 150 733 151
rect 759 151 765 152
rect 759 150 760 151
rect 732 148 760 150
rect 732 147 733 148
rect 727 146 733 147
rect 759 147 760 148
rect 764 147 765 151
rect 759 146 765 147
rect 815 151 821 152
rect 815 147 816 151
rect 820 150 821 151
rect 847 151 853 152
rect 847 150 848 151
rect 820 148 848 150
rect 820 147 821 148
rect 815 146 821 147
rect 847 147 848 148
rect 852 147 853 151
rect 847 146 853 147
rect 903 151 909 152
rect 903 147 904 151
rect 908 150 909 151
rect 935 151 941 152
rect 935 150 936 151
rect 908 148 936 150
rect 908 147 909 148
rect 903 146 909 147
rect 935 147 936 148
rect 940 147 941 151
rect 935 146 941 147
rect 991 151 997 152
rect 991 147 992 151
rect 996 150 997 151
rect 1023 151 1029 152
rect 1023 150 1024 151
rect 996 148 1024 150
rect 996 147 997 148
rect 991 146 997 147
rect 1023 147 1024 148
rect 1028 147 1029 151
rect 1023 146 1029 147
rect 1079 151 1085 152
rect 1079 147 1080 151
rect 1084 150 1085 151
rect 1111 151 1117 152
rect 1111 150 1112 151
rect 1084 148 1112 150
rect 1084 147 1085 148
rect 1079 146 1085 147
rect 1111 147 1112 148
rect 1116 147 1117 151
rect 1111 146 1117 147
rect 1162 151 1168 152
rect 1162 147 1163 151
rect 1167 150 1168 151
rect 1199 151 1205 152
rect 1199 150 1200 151
rect 1167 148 1200 150
rect 1167 147 1168 148
rect 1162 146 1168 147
rect 1199 147 1200 148
rect 1204 147 1205 151
rect 1199 146 1205 147
rect 1255 151 1261 152
rect 1255 147 1256 151
rect 1260 150 1261 151
rect 1303 151 1309 152
rect 1303 150 1304 151
rect 1260 148 1304 150
rect 1260 147 1261 148
rect 1255 146 1261 147
rect 1303 147 1304 148
rect 1308 147 1309 151
rect 1303 146 1309 147
rect 1359 151 1365 152
rect 1359 147 1360 151
rect 1364 150 1365 151
rect 1407 151 1413 152
rect 1407 150 1408 151
rect 1364 148 1408 150
rect 1364 147 1365 148
rect 1359 146 1365 147
rect 1407 147 1408 148
rect 1412 147 1413 151
rect 1407 146 1413 147
rect 1463 151 1469 152
rect 1463 147 1464 151
rect 1468 150 1469 151
rect 1519 151 1525 152
rect 1519 150 1520 151
rect 1468 148 1520 150
rect 1468 147 1469 148
rect 1463 146 1469 147
rect 1519 147 1520 148
rect 1524 147 1525 151
rect 1519 146 1525 147
rect 1575 151 1581 152
rect 1575 147 1576 151
rect 1580 150 1581 151
rect 1639 151 1645 152
rect 1639 150 1640 151
rect 1580 148 1640 150
rect 1580 147 1581 148
rect 1575 146 1581 147
rect 1639 147 1640 148
rect 1644 147 1645 151
rect 1639 146 1645 147
rect 1726 151 1732 152
rect 1726 147 1727 151
rect 1731 150 1732 151
rect 1743 151 1749 152
rect 1743 150 1744 151
rect 1731 148 1744 150
rect 1731 147 1732 148
rect 1726 146 1732 147
rect 1743 147 1744 148
rect 1748 147 1749 151
rect 1743 146 1749 147
rect 1807 147 1813 148
rect 1807 143 1808 147
rect 1812 146 1813 147
rect 1903 147 1909 148
rect 1903 146 1904 147
rect 1812 144 1904 146
rect 1812 143 1813 144
rect 1807 142 1813 143
rect 1903 143 1904 144
rect 1908 143 1909 147
rect 1903 142 1909 143
rect 1959 147 1965 148
rect 1959 143 1960 147
rect 1964 146 1965 147
rect 1991 147 1997 148
rect 1991 146 1992 147
rect 1964 144 1992 146
rect 1964 143 1965 144
rect 1959 142 1965 143
rect 1991 143 1992 144
rect 1996 143 1997 147
rect 1991 142 1997 143
rect 2055 147 2061 148
rect 2055 143 2056 147
rect 2060 146 2061 147
rect 2079 147 2085 148
rect 2079 146 2080 147
rect 2060 144 2080 146
rect 2060 143 2061 144
rect 2055 142 2061 143
rect 2079 143 2080 144
rect 2084 143 2085 147
rect 2079 142 2085 143
rect 2135 147 2141 148
rect 2135 143 2136 147
rect 2140 146 2141 147
rect 2167 147 2173 148
rect 2167 146 2168 147
rect 2140 144 2168 146
rect 2140 143 2141 144
rect 2135 142 2141 143
rect 2167 143 2168 144
rect 2172 143 2173 147
rect 2167 142 2173 143
rect 2223 147 2229 148
rect 2223 143 2224 147
rect 2228 146 2229 147
rect 2279 147 2285 148
rect 2279 146 2280 147
rect 2228 144 2280 146
rect 2228 143 2229 144
rect 2223 142 2229 143
rect 2279 143 2280 144
rect 2284 143 2285 147
rect 2279 142 2285 143
rect 2335 147 2341 148
rect 2335 143 2336 147
rect 2340 146 2341 147
rect 2391 147 2397 148
rect 2391 146 2392 147
rect 2340 144 2392 146
rect 2340 143 2341 144
rect 2335 142 2341 143
rect 2391 143 2392 144
rect 2396 143 2397 147
rect 2391 142 2397 143
rect 2442 147 2448 148
rect 2442 143 2443 147
rect 2447 146 2448 147
rect 2503 147 2509 148
rect 2503 146 2504 147
rect 2447 144 2504 146
rect 2447 143 2448 144
rect 2442 142 2448 143
rect 2503 143 2504 144
rect 2508 143 2509 147
rect 2503 142 2509 143
rect 2615 147 2624 148
rect 2615 143 2616 147
rect 2623 143 2624 147
rect 2615 142 2624 143
rect 2671 147 2677 148
rect 2671 143 2672 147
rect 2676 146 2677 147
rect 2727 147 2733 148
rect 2727 146 2728 147
rect 2676 144 2728 146
rect 2676 143 2677 144
rect 2671 142 2677 143
rect 2727 143 2728 144
rect 2732 143 2733 147
rect 2727 142 2733 143
rect 2783 147 2789 148
rect 2783 143 2784 147
rect 2788 146 2789 147
rect 2831 147 2837 148
rect 2831 146 2832 147
rect 2788 144 2832 146
rect 2788 143 2789 144
rect 2783 142 2789 143
rect 2831 143 2832 144
rect 2836 143 2837 147
rect 2831 142 2837 143
rect 2911 147 2917 148
rect 2911 143 2912 147
rect 2916 146 2917 147
rect 2935 147 2941 148
rect 2935 146 2936 147
rect 2916 144 2936 146
rect 2916 143 2917 144
rect 2911 142 2917 143
rect 2935 143 2936 144
rect 2940 143 2941 147
rect 2935 142 2941 143
rect 2991 147 2997 148
rect 2991 143 2992 147
rect 2996 146 2997 147
rect 3031 147 3037 148
rect 3031 146 3032 147
rect 2996 144 3032 146
rect 2996 143 2997 144
rect 2991 142 2997 143
rect 3031 143 3032 144
rect 3036 143 3037 147
rect 3031 142 3037 143
rect 3087 147 3093 148
rect 3087 143 3088 147
rect 3092 146 3093 147
rect 3127 147 3133 148
rect 3127 146 3128 147
rect 3092 144 3128 146
rect 3092 143 3093 144
rect 3087 142 3093 143
rect 3127 143 3128 144
rect 3132 143 3133 147
rect 3127 142 3133 143
rect 3183 147 3189 148
rect 3183 143 3184 147
rect 3188 146 3189 147
rect 3223 147 3229 148
rect 3223 146 3224 147
rect 3188 144 3224 146
rect 3188 143 3189 144
rect 3183 142 3189 143
rect 3223 143 3224 144
rect 3228 143 3229 147
rect 3223 142 3229 143
rect 3279 147 3285 148
rect 3279 143 3280 147
rect 3284 146 3285 147
rect 3319 147 3325 148
rect 3319 146 3320 147
rect 3284 144 3320 146
rect 3284 143 3285 144
rect 3279 142 3285 143
rect 3319 143 3320 144
rect 3324 143 3325 147
rect 3319 142 3325 143
rect 3375 147 3381 148
rect 3375 143 3376 147
rect 3380 146 3381 147
rect 3407 147 3413 148
rect 3407 146 3408 147
rect 3380 144 3408 146
rect 3380 143 3381 144
rect 3375 142 3381 143
rect 3407 143 3408 144
rect 3412 143 3413 147
rect 3407 142 3413 143
rect 3463 147 3469 148
rect 3463 143 3464 147
rect 3468 146 3469 147
rect 3495 147 3501 148
rect 3495 146 3496 147
rect 3468 144 3496 146
rect 3468 143 3469 144
rect 3463 142 3469 143
rect 3495 143 3496 144
rect 3500 143 3501 147
rect 3495 142 3501 143
rect 222 141 228 142
rect 222 137 223 141
rect 227 137 228 141
rect 222 136 228 137
rect 310 141 316 142
rect 310 137 311 141
rect 315 137 316 141
rect 310 136 316 137
rect 398 141 404 142
rect 398 137 399 141
rect 403 137 404 141
rect 398 136 404 137
rect 486 141 492 142
rect 486 137 487 141
rect 491 137 492 141
rect 486 136 492 137
rect 574 141 580 142
rect 574 137 575 141
rect 579 137 580 141
rect 574 136 580 137
rect 662 141 668 142
rect 662 137 663 141
rect 667 137 668 141
rect 662 136 668 137
rect 750 141 756 142
rect 750 137 751 141
rect 755 137 756 141
rect 750 136 756 137
rect 838 141 844 142
rect 838 137 839 141
rect 843 137 844 141
rect 838 136 844 137
rect 926 141 932 142
rect 926 137 927 141
rect 931 137 932 141
rect 926 136 932 137
rect 1014 141 1020 142
rect 1014 137 1015 141
rect 1019 137 1020 141
rect 1014 136 1020 137
rect 1102 141 1108 142
rect 1102 137 1103 141
rect 1107 137 1108 141
rect 1102 136 1108 137
rect 1190 141 1196 142
rect 1190 137 1191 141
rect 1195 137 1196 141
rect 1190 136 1196 137
rect 1294 141 1300 142
rect 1294 137 1295 141
rect 1299 137 1300 141
rect 1294 136 1300 137
rect 1398 141 1404 142
rect 1398 137 1399 141
rect 1403 137 1404 141
rect 1398 136 1404 137
rect 1510 141 1516 142
rect 1510 137 1511 141
rect 1515 137 1516 141
rect 1510 136 1516 137
rect 1630 141 1636 142
rect 1630 137 1631 141
rect 1635 137 1636 141
rect 1630 136 1636 137
rect 1734 141 1740 142
rect 1734 137 1735 141
rect 1739 137 1740 141
rect 1734 136 1740 137
rect 1894 137 1900 138
rect 1894 133 1895 137
rect 1899 133 1900 137
rect 1894 132 1900 133
rect 1982 137 1988 138
rect 1982 133 1983 137
rect 1987 133 1988 137
rect 1982 132 1988 133
rect 2070 137 2076 138
rect 2070 133 2071 137
rect 2075 133 2076 137
rect 2070 132 2076 133
rect 2158 137 2164 138
rect 2158 133 2159 137
rect 2163 133 2164 137
rect 2158 132 2164 133
rect 2270 137 2276 138
rect 2270 133 2271 137
rect 2275 133 2276 137
rect 2270 132 2276 133
rect 2382 137 2388 138
rect 2382 133 2383 137
rect 2387 133 2388 137
rect 2382 132 2388 133
rect 2494 137 2500 138
rect 2494 133 2495 137
rect 2499 133 2500 137
rect 2494 132 2500 133
rect 2606 137 2612 138
rect 2606 133 2607 137
rect 2611 133 2612 137
rect 2606 132 2612 133
rect 2718 137 2724 138
rect 2718 133 2719 137
rect 2723 133 2724 137
rect 2718 132 2724 133
rect 2822 137 2828 138
rect 2822 133 2823 137
rect 2827 133 2828 137
rect 2822 132 2828 133
rect 2926 137 2932 138
rect 2926 133 2927 137
rect 2931 133 2932 137
rect 2926 132 2932 133
rect 3022 137 3028 138
rect 3022 133 3023 137
rect 3027 133 3028 137
rect 3022 132 3028 133
rect 3118 137 3124 138
rect 3118 133 3119 137
rect 3123 133 3124 137
rect 3118 132 3124 133
rect 3214 137 3220 138
rect 3214 133 3215 137
rect 3219 133 3220 137
rect 3214 132 3220 133
rect 3310 137 3316 138
rect 3310 133 3311 137
rect 3315 133 3316 137
rect 3310 132 3316 133
rect 3398 137 3404 138
rect 3398 133 3399 137
rect 3403 133 3404 137
rect 3398 132 3404 133
rect 3486 137 3492 138
rect 3486 133 3487 137
rect 3491 133 3492 137
rect 3486 132 3492 133
rect 110 128 116 129
rect 1822 128 1828 129
rect 110 124 111 128
rect 115 124 116 128
rect 287 127 293 128
rect 287 126 288 127
rect 277 124 288 126
rect 110 123 116 124
rect 287 123 288 124
rect 292 123 293 127
rect 375 127 381 128
rect 375 126 376 127
rect 365 124 376 126
rect 287 122 293 123
rect 375 123 376 124
rect 380 123 381 127
rect 463 127 469 128
rect 463 126 464 127
rect 453 124 464 126
rect 375 122 381 123
rect 463 123 464 124
rect 468 123 469 127
rect 551 127 557 128
rect 551 126 552 127
rect 541 124 552 126
rect 463 122 469 123
rect 551 123 552 124
rect 556 123 557 127
rect 639 127 645 128
rect 639 126 640 127
rect 629 124 640 126
rect 551 122 557 123
rect 639 123 640 124
rect 644 123 645 127
rect 727 127 733 128
rect 727 126 728 127
rect 717 124 728 126
rect 639 122 645 123
rect 727 123 728 124
rect 732 123 733 127
rect 815 127 821 128
rect 815 126 816 127
rect 805 124 816 126
rect 727 122 733 123
rect 815 123 816 124
rect 820 123 821 127
rect 903 127 909 128
rect 903 126 904 127
rect 893 124 904 126
rect 815 122 821 123
rect 903 123 904 124
rect 908 123 909 127
rect 991 127 997 128
rect 991 126 992 127
rect 981 124 992 126
rect 903 122 909 123
rect 991 123 992 124
rect 996 123 997 127
rect 1079 127 1085 128
rect 1079 126 1080 127
rect 1069 124 1080 126
rect 991 122 997 123
rect 1079 123 1080 124
rect 1084 123 1085 127
rect 1162 127 1168 128
rect 1162 126 1163 127
rect 1157 124 1163 126
rect 1079 122 1085 123
rect 1162 123 1163 124
rect 1167 123 1168 127
rect 1255 127 1261 128
rect 1255 126 1256 127
rect 1245 124 1256 126
rect 1162 122 1168 123
rect 1255 123 1256 124
rect 1260 123 1261 127
rect 1359 127 1365 128
rect 1359 126 1360 127
rect 1349 124 1360 126
rect 1255 122 1261 123
rect 1359 123 1360 124
rect 1364 123 1365 127
rect 1463 127 1469 128
rect 1463 126 1464 127
rect 1453 124 1464 126
rect 1359 122 1365 123
rect 1463 123 1464 124
rect 1468 123 1469 127
rect 1575 127 1581 128
rect 1575 126 1576 127
rect 1565 124 1576 126
rect 1463 122 1469 123
rect 1575 123 1576 124
rect 1580 123 1581 127
rect 1807 127 1813 128
rect 1807 126 1808 127
rect 1789 124 1808 126
rect 1575 122 1581 123
rect 1583 123 1589 124
rect 1583 119 1584 123
rect 1588 122 1589 123
rect 1807 123 1808 124
rect 1812 123 1813 127
rect 1822 124 1823 128
rect 1827 124 1828 128
rect 1822 123 1828 124
rect 1862 124 1868 125
rect 3574 124 3580 125
rect 1807 122 1813 123
rect 1588 120 1649 122
rect 1862 120 1863 124
rect 1867 120 1868 124
rect 1959 123 1965 124
rect 1959 122 1960 123
rect 1949 120 1960 122
rect 1588 119 1589 120
rect 1862 119 1868 120
rect 1959 119 1960 120
rect 1964 119 1965 123
rect 2055 123 2061 124
rect 2055 122 2056 123
rect 2037 120 2056 122
rect 1583 118 1589 119
rect 1959 118 1965 119
rect 2055 119 2056 120
rect 2060 119 2061 123
rect 2135 123 2141 124
rect 2135 122 2136 123
rect 2125 120 2136 122
rect 2055 118 2061 119
rect 2135 119 2136 120
rect 2140 119 2141 123
rect 2223 123 2229 124
rect 2223 122 2224 123
rect 2213 120 2224 122
rect 2135 118 2141 119
rect 2223 119 2224 120
rect 2228 119 2229 123
rect 2335 123 2341 124
rect 2335 122 2336 123
rect 2325 120 2336 122
rect 2223 118 2229 119
rect 2335 119 2336 120
rect 2340 119 2341 123
rect 2442 123 2448 124
rect 2442 122 2443 123
rect 2437 120 2443 122
rect 2335 118 2341 119
rect 2442 119 2443 120
rect 2447 119 2448 123
rect 2671 123 2677 124
rect 2671 122 2672 123
rect 2661 120 2672 122
rect 2442 118 2448 119
rect 2450 119 2456 120
rect 2450 115 2451 119
rect 2455 118 2456 119
rect 2671 119 2672 120
rect 2676 119 2677 123
rect 2783 123 2789 124
rect 2783 122 2784 123
rect 2773 120 2784 122
rect 2671 118 2677 119
rect 2783 119 2784 120
rect 2788 119 2789 123
rect 2911 123 2917 124
rect 2911 122 2912 123
rect 2877 120 2912 122
rect 2783 118 2789 119
rect 2911 119 2912 120
rect 2916 119 2917 123
rect 2991 123 2997 124
rect 2991 122 2992 123
rect 2981 120 2992 122
rect 2911 118 2917 119
rect 2991 119 2992 120
rect 2996 119 2997 123
rect 3087 123 3093 124
rect 3087 122 3088 123
rect 3077 120 3088 122
rect 2991 118 2997 119
rect 3087 119 3088 120
rect 3092 119 3093 123
rect 3183 123 3189 124
rect 3183 122 3184 123
rect 3173 120 3184 122
rect 3087 118 3093 119
rect 3183 119 3184 120
rect 3188 119 3189 123
rect 3279 123 3285 124
rect 3279 122 3280 123
rect 3269 120 3280 122
rect 3183 118 3189 119
rect 3279 119 3280 120
rect 3284 119 3285 123
rect 3375 123 3381 124
rect 3375 122 3376 123
rect 3365 120 3376 122
rect 3279 118 3285 119
rect 3375 119 3376 120
rect 3380 119 3381 123
rect 3463 123 3469 124
rect 3463 122 3464 123
rect 3453 120 3464 122
rect 3375 118 3381 119
rect 3463 119 3464 120
rect 3468 119 3469 123
rect 3574 120 3575 124
rect 3579 120 3580 124
rect 3463 118 3469 119
rect 3478 119 3484 120
rect 3574 119 3580 120
rect 2455 116 2513 118
rect 2455 115 2456 116
rect 2450 114 2456 115
rect 3478 115 3479 119
rect 3483 118 3484 119
rect 3483 116 3505 118
rect 3483 115 3484 116
rect 3478 114 3484 115
rect 110 111 116 112
rect 110 107 111 111
rect 115 107 116 111
rect 110 106 116 107
rect 1822 111 1828 112
rect 1822 107 1823 111
rect 1827 107 1828 111
rect 1822 106 1828 107
rect 1862 107 1868 108
rect 1862 103 1863 107
rect 1867 103 1868 107
rect 1862 102 1868 103
rect 3574 107 3580 108
rect 3574 103 3575 107
rect 3579 103 3580 107
rect 3574 102 3580 103
rect 214 101 220 102
rect 214 97 215 101
rect 219 97 220 101
rect 214 96 220 97
rect 302 101 308 102
rect 302 97 303 101
rect 307 97 308 101
rect 302 96 308 97
rect 390 101 396 102
rect 390 97 391 101
rect 395 97 396 101
rect 390 96 396 97
rect 478 101 484 102
rect 478 97 479 101
rect 483 97 484 101
rect 478 96 484 97
rect 566 101 572 102
rect 566 97 567 101
rect 571 97 572 101
rect 566 96 572 97
rect 654 101 660 102
rect 654 97 655 101
rect 659 97 660 101
rect 654 96 660 97
rect 742 101 748 102
rect 742 97 743 101
rect 747 97 748 101
rect 742 96 748 97
rect 830 101 836 102
rect 830 97 831 101
rect 835 97 836 101
rect 830 96 836 97
rect 918 101 924 102
rect 918 97 919 101
rect 923 97 924 101
rect 918 96 924 97
rect 1006 101 1012 102
rect 1006 97 1007 101
rect 1011 97 1012 101
rect 1006 96 1012 97
rect 1094 101 1100 102
rect 1094 97 1095 101
rect 1099 97 1100 101
rect 1094 96 1100 97
rect 1182 101 1188 102
rect 1182 97 1183 101
rect 1187 97 1188 101
rect 1182 96 1188 97
rect 1286 101 1292 102
rect 1286 97 1287 101
rect 1291 97 1292 101
rect 1286 96 1292 97
rect 1390 101 1396 102
rect 1390 97 1391 101
rect 1395 97 1396 101
rect 1390 96 1396 97
rect 1502 101 1508 102
rect 1502 97 1503 101
rect 1507 97 1508 101
rect 1502 96 1508 97
rect 1622 101 1628 102
rect 1622 97 1623 101
rect 1627 97 1628 101
rect 1622 96 1628 97
rect 1726 101 1732 102
rect 1726 97 1727 101
rect 1731 97 1732 101
rect 1726 96 1732 97
rect 1886 97 1892 98
rect 1886 93 1887 97
rect 1891 93 1892 97
rect 1886 92 1892 93
rect 1974 97 1980 98
rect 1974 93 1975 97
rect 1979 93 1980 97
rect 1974 92 1980 93
rect 2062 97 2068 98
rect 2062 93 2063 97
rect 2067 93 2068 97
rect 2062 92 2068 93
rect 2150 97 2156 98
rect 2150 93 2151 97
rect 2155 93 2156 97
rect 2150 92 2156 93
rect 2262 97 2268 98
rect 2262 93 2263 97
rect 2267 93 2268 97
rect 2262 92 2268 93
rect 2374 97 2380 98
rect 2374 93 2375 97
rect 2379 93 2380 97
rect 2374 92 2380 93
rect 2486 97 2492 98
rect 2486 93 2487 97
rect 2491 93 2492 97
rect 2486 92 2492 93
rect 2598 97 2604 98
rect 2598 93 2599 97
rect 2603 93 2604 97
rect 2598 92 2604 93
rect 2710 97 2716 98
rect 2710 93 2711 97
rect 2715 93 2716 97
rect 2710 92 2716 93
rect 2814 97 2820 98
rect 2814 93 2815 97
rect 2819 93 2820 97
rect 2814 92 2820 93
rect 2918 97 2924 98
rect 2918 93 2919 97
rect 2923 93 2924 97
rect 2918 92 2924 93
rect 3014 97 3020 98
rect 3014 93 3015 97
rect 3019 93 3020 97
rect 3014 92 3020 93
rect 3110 97 3116 98
rect 3110 93 3111 97
rect 3115 93 3116 97
rect 3110 92 3116 93
rect 3206 97 3212 98
rect 3206 93 3207 97
rect 3211 93 3212 97
rect 3206 92 3212 93
rect 3302 97 3308 98
rect 3302 93 3303 97
rect 3307 93 3308 97
rect 3302 92 3308 93
rect 3390 97 3396 98
rect 3390 93 3391 97
rect 3395 93 3396 97
rect 3390 92 3396 93
rect 3478 97 3484 98
rect 3478 93 3479 97
rect 3483 93 3484 97
rect 3478 92 3484 93
<< m3c >>
rect 143 3629 147 3633
rect 231 3629 235 3633
rect 319 3629 323 3633
rect 407 3629 411 3633
rect 495 3629 499 3633
rect 583 3629 587 3633
rect 671 3629 675 3633
rect 111 3616 115 3620
rect 1823 3616 1827 3620
rect 111 3599 115 3603
rect 651 3599 655 3603
rect 1823 3599 1827 3603
rect 135 3589 139 3593
rect 223 3589 227 3593
rect 311 3589 315 3593
rect 399 3589 403 3593
rect 487 3589 491 3593
rect 575 3589 579 3593
rect 663 3589 667 3593
rect 1547 3567 1551 3571
rect 135 3559 139 3563
rect 287 3559 291 3563
rect 463 3559 467 3563
rect 631 3559 635 3563
rect 791 3559 795 3563
rect 935 3559 939 3563
rect 1071 3559 1075 3563
rect 1191 3559 1195 3563
rect 1311 3559 1315 3563
rect 1423 3559 1427 3563
rect 1527 3559 1531 3563
rect 1639 3559 1643 3563
rect 111 3549 115 3553
rect 559 3551 563 3555
rect 1727 3559 1731 3563
rect 1823 3549 1827 3553
rect 111 3532 115 3536
rect 1823 3532 1827 3536
rect 143 3519 147 3523
rect 295 3519 299 3523
rect 471 3519 475 3523
rect 639 3519 643 3523
rect 799 3519 803 3523
rect 943 3519 947 3523
rect 1079 3519 1083 3523
rect 1199 3519 1203 3523
rect 1319 3519 1323 3523
rect 1431 3519 1435 3523
rect 1535 3519 1539 3523
rect 1647 3519 1651 3523
rect 1735 3519 1739 3523
rect 167 3507 171 3511
rect 807 3513 811 3515
rect 807 3511 808 3513
rect 808 3511 811 3513
rect 159 3495 160 3499
rect 160 3495 163 3499
rect 879 3495 883 3499
rect 1147 3495 1151 3499
rect 1547 3495 1548 3499
rect 1548 3495 1551 3499
rect 151 3485 155 3489
rect 327 3485 331 3489
rect 495 3485 499 3489
rect 655 3485 659 3489
rect 807 3485 811 3489
rect 951 3485 955 3489
rect 1087 3485 1091 3489
rect 1207 3485 1211 3489
rect 1319 3485 1323 3489
rect 1431 3485 1435 3489
rect 1535 3485 1539 3489
rect 1647 3485 1651 3489
rect 1735 3485 1739 3489
rect 1895 3481 1899 3485
rect 1983 3481 1987 3485
rect 2071 3481 2075 3485
rect 2159 3481 2163 3485
rect 111 3472 115 3476
rect 1147 3471 1151 3475
rect 1395 3467 1399 3471
rect 1823 3472 1827 3476
rect 1863 3468 1867 3472
rect 3575 3468 3579 3472
rect 111 3455 115 3459
rect 563 3455 567 3459
rect 1823 3455 1827 3459
rect 1863 3451 1867 3455
rect 2139 3451 2143 3455
rect 3575 3451 3579 3455
rect 143 3445 147 3449
rect 319 3445 323 3449
rect 487 3445 491 3449
rect 647 3445 651 3449
rect 799 3445 803 3449
rect 943 3445 947 3449
rect 1079 3445 1083 3449
rect 1199 3445 1203 3449
rect 1311 3445 1315 3449
rect 1423 3445 1427 3449
rect 1527 3445 1531 3449
rect 1639 3445 1643 3449
rect 1727 3445 1731 3449
rect 1887 3441 1891 3445
rect 1975 3441 1979 3445
rect 2063 3441 2067 3445
rect 2151 3441 2155 3445
rect 1915 3435 1919 3439
rect 215 3423 219 3427
rect 431 3423 435 3427
rect 639 3423 643 3427
rect 847 3423 851 3427
rect 1039 3423 1043 3427
rect 1223 3423 1227 3427
rect 1399 3423 1403 3427
rect 1567 3423 1571 3427
rect 1727 3423 1731 3427
rect 2139 3427 2143 3431
rect 111 3413 115 3417
rect 739 3415 743 3419
rect 1647 3415 1651 3419
rect 1887 3419 1891 3423
rect 1991 3419 1995 3423
rect 2119 3419 2123 3423
rect 2255 3419 2259 3423
rect 2391 3419 2395 3423
rect 2527 3419 2531 3423
rect 2655 3419 2659 3423
rect 2783 3419 2787 3423
rect 2919 3419 2923 3423
rect 3055 3419 3059 3423
rect 1823 3413 1827 3417
rect 1863 3409 1867 3413
rect 2323 3411 2327 3415
rect 3575 3409 3579 3413
rect 111 3396 115 3400
rect 1823 3396 1827 3400
rect 1863 3392 1867 3396
rect 1955 3395 1959 3399
rect 3123 3395 3127 3399
rect 3575 3392 3579 3396
rect 223 3383 227 3387
rect 439 3383 443 3387
rect 647 3383 651 3387
rect 855 3383 859 3387
rect 1047 3383 1051 3387
rect 1231 3383 1235 3387
rect 1407 3383 1411 3387
rect 1575 3383 1579 3387
rect 1735 3383 1739 3387
rect 1895 3379 1899 3383
rect 1999 3379 2003 3383
rect 2127 3379 2131 3383
rect 2263 3379 2267 3383
rect 2399 3379 2403 3383
rect 2535 3379 2539 3383
rect 2663 3379 2667 3383
rect 2791 3379 2795 3383
rect 2927 3379 2931 3383
rect 3063 3379 3067 3383
rect 235 3371 236 3375
rect 236 3371 239 3375
rect 1207 3371 1211 3375
rect 1915 3367 1919 3371
rect 1955 3367 1959 3371
rect 2547 3367 2548 3371
rect 2548 3367 2551 3371
rect 739 3359 743 3363
rect 1087 3351 1091 3355
rect 1907 3355 1908 3359
rect 1908 3355 1911 3359
rect 2627 3355 2631 3359
rect 2707 3355 2708 3359
rect 2708 3355 2711 3359
rect 2899 3355 2903 3359
rect 3035 3355 3039 3359
rect 3123 3355 3127 3359
rect 239 3341 243 3345
rect 383 3341 387 3345
rect 543 3341 547 3345
rect 711 3341 715 3345
rect 871 3341 875 3345
rect 1031 3341 1035 3345
rect 1183 3341 1187 3345
rect 1335 3341 1339 3345
rect 1487 3341 1491 3345
rect 1639 3341 1643 3345
rect 1895 3345 1899 3349
rect 1999 3345 2003 3349
rect 2135 3345 2139 3349
rect 2279 3345 2283 3349
rect 2423 3345 2427 3349
rect 2559 3345 2563 3349
rect 2695 3345 2699 3349
rect 2831 3345 2835 3349
rect 2967 3345 2971 3349
rect 3103 3345 3107 3349
rect 111 3328 115 3332
rect 1823 3328 1827 3332
rect 1863 3332 1867 3336
rect 3575 3332 3579 3336
rect 2547 3327 2551 3331
rect 1583 3323 1587 3327
rect 2627 3327 2631 3331
rect 2899 3327 2903 3331
rect 3035 3327 3039 3331
rect 111 3311 115 3315
rect 779 3311 783 3315
rect 1823 3311 1827 3315
rect 1863 3315 1867 3319
rect 2359 3315 2363 3319
rect 2903 3315 2907 3319
rect 3575 3315 3579 3319
rect 231 3301 235 3305
rect 375 3301 379 3305
rect 535 3301 539 3305
rect 703 3301 707 3305
rect 863 3301 867 3305
rect 1023 3301 1027 3305
rect 1175 3301 1179 3305
rect 1327 3301 1331 3305
rect 1479 3301 1483 3305
rect 1631 3301 1635 3305
rect 1887 3305 1891 3309
rect 1991 3305 1995 3309
rect 2127 3305 2131 3309
rect 2271 3305 2275 3309
rect 2415 3305 2419 3309
rect 2551 3305 2555 3309
rect 2687 3305 2691 3309
rect 2823 3305 2827 3309
rect 2959 3305 2963 3309
rect 3095 3305 3099 3309
rect 1087 3283 1091 3287
rect 239 3275 243 3279
rect 407 3275 411 3279
rect 575 3275 579 3279
rect 743 3275 747 3279
rect 895 3275 899 3279
rect 1047 3275 1051 3279
rect 1191 3275 1195 3279
rect 1335 3275 1339 3279
rect 111 3265 115 3269
rect 499 3267 503 3271
rect 1927 3283 1931 3287
rect 2047 3283 2051 3287
rect 2175 3283 2179 3287
rect 2311 3283 2315 3287
rect 2455 3283 2459 3287
rect 2599 3283 2603 3287
rect 2743 3283 2747 3287
rect 2887 3283 2891 3287
rect 3031 3283 3035 3287
rect 3183 3283 3187 3287
rect 1487 3275 1491 3279
rect 1863 3273 1867 3277
rect 2383 3275 2387 3279
rect 2707 3275 2711 3279
rect 3575 3273 3579 3277
rect 1823 3265 1827 3269
rect 1863 3256 1867 3260
rect 3287 3259 3291 3263
rect 111 3248 115 3252
rect 567 3251 571 3255
rect 643 3251 647 3255
rect 3575 3256 3579 3260
rect 1823 3248 1827 3252
rect 1935 3243 1939 3247
rect 2055 3243 2059 3247
rect 2183 3243 2187 3247
rect 2319 3243 2323 3247
rect 2463 3243 2467 3247
rect 2607 3243 2611 3247
rect 2751 3243 2755 3247
rect 2895 3243 2899 3247
rect 3039 3243 3043 3247
rect 3191 3243 3195 3247
rect 247 3235 251 3239
rect 415 3235 419 3239
rect 583 3235 587 3239
rect 751 3235 755 3239
rect 903 3235 907 3239
rect 1055 3235 1059 3239
rect 1199 3235 1203 3239
rect 1343 3235 1347 3239
rect 1495 3235 1499 3239
rect 1947 3231 1948 3235
rect 1948 3231 1951 3235
rect 2619 3231 2620 3235
rect 2620 3231 2623 3235
rect 2903 3231 2904 3235
rect 2904 3231 2907 3235
rect 259 3223 260 3227
rect 260 3223 263 3227
rect 643 3223 647 3227
rect 779 3223 783 3227
rect 1031 3223 1035 3227
rect 2383 3219 2387 3223
rect 3047 3211 3051 3215
rect 3287 3211 3288 3215
rect 3288 3211 3291 3215
rect 259 3199 263 3203
rect 479 3199 483 3203
rect 567 3199 568 3203
rect 568 3199 571 3203
rect 807 3199 811 3203
rect 2007 3201 2011 3205
rect 2119 3201 2123 3205
rect 2239 3201 2243 3205
rect 2375 3201 2379 3205
rect 2519 3201 2523 3205
rect 2663 3201 2667 3205
rect 2815 3201 2819 3205
rect 2967 3201 2971 3205
rect 3119 3201 3123 3205
rect 3279 3201 3283 3205
rect 175 3189 179 3193
rect 375 3189 379 3193
rect 559 3189 563 3193
rect 727 3189 731 3193
rect 887 3189 891 3193
rect 1039 3189 1043 3193
rect 1191 3189 1195 3193
rect 1351 3189 1355 3193
rect 1863 3188 1867 3192
rect 3575 3188 3579 3192
rect 2619 3183 2623 3187
rect 3047 3183 3051 3187
rect 111 3176 115 3180
rect 259 3171 263 3175
rect 479 3171 483 3175
rect 1823 3176 1827 3180
rect 1279 3171 1283 3175
rect 1863 3171 1867 3175
rect 3575 3171 3579 3175
rect 111 3159 115 3163
rect 155 3159 159 3163
rect 1823 3159 1827 3163
rect 1999 3161 2003 3165
rect 2111 3161 2115 3165
rect 2231 3161 2235 3165
rect 2367 3161 2371 3165
rect 2511 3161 2515 3165
rect 2655 3161 2659 3165
rect 2807 3161 2811 3165
rect 2959 3161 2963 3165
rect 3111 3161 3115 3165
rect 3271 3161 3275 3165
rect 2531 3155 2535 3159
rect 167 3149 171 3153
rect 367 3149 371 3153
rect 551 3149 555 3153
rect 719 3149 723 3153
rect 879 3149 883 3153
rect 1031 3149 1035 3153
rect 1183 3149 1187 3153
rect 1343 3149 1347 3153
rect 2055 3135 2059 3139
rect 2207 3135 2211 3139
rect 2359 3135 2363 3139
rect 2511 3135 2515 3139
rect 2655 3135 2659 3139
rect 2791 3135 2795 3139
rect 2919 3135 2923 3139
rect 3039 3135 3043 3139
rect 3159 3135 3163 3139
rect 3271 3135 3275 3139
rect 3383 3135 3387 3139
rect 3479 3135 3483 3139
rect 611 3123 615 3127
rect 1863 3125 1867 3129
rect 3451 3127 3455 3131
rect 3575 3125 3579 3129
rect 135 3115 139 3119
rect 263 3115 267 3119
rect 399 3115 403 3119
rect 527 3115 531 3119
rect 647 3115 651 3119
rect 111 3105 115 3109
rect 255 3107 259 3111
rect 759 3115 763 3119
rect 863 3115 867 3119
rect 967 3115 971 3119
rect 1071 3115 1075 3119
rect 1175 3115 1179 3119
rect 1279 3115 1283 3119
rect 1243 3107 1247 3111
rect 1823 3105 1827 3109
rect 1863 3108 1867 3112
rect 1963 3111 1967 3115
rect 2123 3111 2127 3115
rect 2275 3111 2279 3115
rect 2427 3111 2431 3115
rect 3119 3111 3123 3115
rect 3575 3108 3579 3112
rect 111 3088 115 3092
rect 2063 3095 2067 3099
rect 2215 3095 2219 3099
rect 2367 3095 2371 3099
rect 2519 3095 2523 3099
rect 2663 3095 2667 3099
rect 2799 3095 2803 3099
rect 2927 3095 2931 3099
rect 3047 3095 3051 3099
rect 3167 3095 3171 3099
rect 3279 3095 3283 3099
rect 3391 3095 3395 3099
rect 3487 3095 3491 3099
rect 1823 3088 1827 3092
rect 2123 3083 2127 3087
rect 2275 3083 2279 3087
rect 2427 3083 2431 3087
rect 2531 3083 2532 3087
rect 2532 3083 2535 3087
rect 2671 3083 2672 3087
rect 2672 3083 2675 3087
rect 3179 3083 3180 3087
rect 3180 3083 3183 3087
rect 143 3075 147 3079
rect 271 3075 275 3079
rect 407 3075 411 3079
rect 535 3075 539 3079
rect 655 3075 659 3079
rect 767 3075 771 3079
rect 871 3075 875 3079
rect 975 3075 979 3079
rect 1079 3075 1083 3079
rect 1183 3075 1187 3079
rect 1287 3075 1291 3079
rect 155 3063 156 3067
rect 156 3063 159 3067
rect 427 3063 431 3067
rect 951 3063 955 3067
rect 1963 3067 1964 3071
rect 1964 3067 1967 3071
rect 2043 3067 2047 3071
rect 2767 3067 2771 3071
rect 2867 3067 2871 3071
rect 3119 3067 3120 3071
rect 3120 3067 3123 3071
rect 3359 3067 3363 3071
rect 3451 3075 3455 3079
rect 1951 3057 1955 3061
rect 2079 3057 2083 3061
rect 2215 3057 2219 3061
rect 2367 3057 2371 3061
rect 2527 3057 2531 3061
rect 2679 3057 2683 3061
rect 2831 3057 2835 3061
rect 2975 3057 2979 3061
rect 3111 3057 3115 3061
rect 3239 3057 3243 3061
rect 3375 3057 3379 3061
rect 3487 3057 3491 3061
rect 211 3051 215 3055
rect 255 3051 256 3055
rect 256 3051 259 3055
rect 439 3051 443 3055
rect 523 3051 527 3055
rect 611 3051 612 3055
rect 612 3051 615 3055
rect 999 3051 1000 3055
rect 1000 3051 1003 3055
rect 1147 3051 1151 3055
rect 1243 3051 1247 3055
rect 143 3041 147 3045
rect 247 3041 251 3045
rect 367 3041 371 3045
rect 487 3041 491 3045
rect 599 3041 603 3045
rect 703 3041 707 3045
rect 799 3041 803 3045
rect 895 3041 899 3045
rect 991 3041 995 3045
rect 1087 3041 1091 3045
rect 1183 3041 1187 3045
rect 1287 3041 1291 3045
rect 1863 3044 1867 3048
rect 2043 3043 2047 3047
rect 2671 3039 2675 3043
rect 2767 3039 2771 3043
rect 3179 3039 3183 3043
rect 3575 3044 3579 3048
rect 111 3028 115 3032
rect 211 3023 215 3027
rect 427 3027 431 3031
rect 439 3023 443 3027
rect 1147 3027 1151 3031
rect 1243 3027 1247 3031
rect 1823 3028 1827 3032
rect 1863 3027 1867 3031
rect 1251 3023 1255 3027
rect 2595 3027 2599 3031
rect 1943 3017 1947 3021
rect 2071 3017 2075 3021
rect 2207 3017 2211 3021
rect 2359 3017 2363 3021
rect 2519 3017 2523 3021
rect 2671 3017 2675 3021
rect 2823 3017 2827 3021
rect 111 3011 115 3015
rect 1823 3011 1827 3015
rect 2707 3011 2711 3015
rect 3575 3027 3579 3031
rect 2967 3017 2971 3021
rect 3103 3017 3107 3021
rect 3231 3017 3235 3021
rect 3367 3017 3371 3021
rect 3479 3017 3483 3021
rect 3499 3011 3503 3015
rect 135 3001 139 3005
rect 239 3001 243 3005
rect 359 3001 363 3005
rect 479 3001 483 3005
rect 591 3001 595 3005
rect 695 3001 699 3005
rect 791 3001 795 3005
rect 887 3001 891 3005
rect 983 3001 987 3005
rect 1079 3001 1083 3005
rect 1175 3001 1179 3005
rect 1279 3001 1283 3005
rect 155 2995 159 2999
rect 947 2995 951 2999
rect 1887 2983 1891 2987
rect 1975 2983 1979 2987
rect 2063 2983 2067 2987
rect 2151 2983 2155 2987
rect 2239 2983 2243 2987
rect 2351 2983 2355 2987
rect 2463 2983 2467 2987
rect 2575 2983 2579 2987
rect 2687 2983 2691 2987
rect 2799 2983 2803 2987
rect 2903 2983 2907 2987
rect 3007 2983 3011 2987
rect 3103 2983 3107 2987
rect 3199 2983 3203 2987
rect 3295 2983 3299 2987
rect 3391 2983 3395 2987
rect 3479 2983 3483 2987
rect 1863 2973 1867 2977
rect 2867 2975 2871 2979
rect 3363 2975 3367 2979
rect 3575 2973 3579 2977
rect 135 2967 139 2971
rect 287 2967 291 2971
rect 455 2967 459 2971
rect 623 2967 627 2971
rect 783 2967 787 2971
rect 927 2967 931 2971
rect 1063 2967 1067 2971
rect 1191 2967 1195 2971
rect 1311 2967 1315 2971
rect 1423 2967 1427 2971
rect 1527 2967 1531 2971
rect 1639 2967 1643 2971
rect 1727 2967 1731 2971
rect 111 2957 115 2961
rect 523 2959 527 2963
rect 691 2959 695 2963
rect 999 2959 1003 2963
rect 1823 2957 1827 2961
rect 1863 2956 1867 2960
rect 1871 2959 1875 2963
rect 1955 2959 1959 2963
rect 2043 2959 2047 2963
rect 2131 2959 2135 2963
rect 2219 2959 2223 2963
rect 2307 2959 2311 2963
rect 2419 2959 2423 2963
rect 2531 2959 2535 2963
rect 3575 2956 3579 2960
rect 111 2940 115 2944
rect 355 2943 359 2947
rect 1407 2943 1411 2947
rect 1415 2943 1419 2947
rect 1491 2943 1495 2947
rect 1595 2943 1599 2947
rect 1823 2940 1827 2944
rect 1895 2943 1899 2947
rect 1983 2943 1987 2947
rect 2071 2943 2075 2947
rect 2159 2943 2163 2947
rect 2247 2943 2251 2947
rect 2359 2943 2363 2947
rect 2471 2943 2475 2947
rect 2583 2943 2587 2947
rect 2695 2943 2699 2947
rect 2807 2943 2811 2947
rect 2911 2943 2915 2947
rect 3015 2943 3019 2947
rect 3111 2943 3115 2947
rect 3207 2943 3211 2947
rect 3303 2943 3307 2947
rect 3399 2943 3403 2947
rect 3487 2943 3491 2947
rect 143 2927 147 2931
rect 295 2927 299 2931
rect 463 2927 467 2931
rect 631 2927 635 2931
rect 791 2927 795 2931
rect 935 2927 939 2931
rect 1071 2927 1075 2931
rect 1199 2927 1203 2931
rect 1319 2927 1323 2931
rect 1431 2927 1435 2931
rect 1535 2927 1539 2931
rect 1647 2927 1651 2931
rect 1735 2927 1739 2931
rect 1955 2931 1959 2935
rect 2043 2931 2047 2935
rect 2131 2931 2135 2935
rect 2219 2931 2223 2935
rect 2307 2931 2311 2935
rect 2419 2931 2423 2935
rect 2531 2931 2535 2935
rect 2595 2931 2596 2935
rect 2596 2931 2599 2935
rect 2707 2931 2708 2935
rect 2708 2931 2711 2935
rect 2955 2931 2959 2935
rect 3499 2931 3500 2935
rect 3500 2931 3503 2935
rect 155 2915 156 2919
rect 156 2915 159 2919
rect 475 2915 476 2919
rect 476 2915 479 2919
rect 947 2915 948 2919
rect 948 2915 951 2919
rect 1119 2915 1123 2919
rect 1491 2915 1495 2919
rect 1595 2915 1599 2919
rect 1871 2915 1875 2919
rect 3163 2911 3167 2915
rect 235 2903 239 2907
rect 355 2903 359 2907
rect 779 2903 783 2907
rect 903 2903 904 2907
rect 904 2903 907 2907
rect 1119 2903 1123 2907
rect 1163 2903 1167 2907
rect 1407 2903 1408 2907
rect 1408 2903 1411 2907
rect 2895 2901 2899 2905
rect 3199 2901 3203 2905
rect 3487 2901 3491 2905
rect 143 2893 147 2897
rect 319 2893 323 2897
rect 519 2893 523 2897
rect 711 2893 715 2897
rect 895 2893 899 2897
rect 1071 2893 1075 2897
rect 1239 2893 1243 2897
rect 1399 2893 1403 2897
rect 1551 2893 1555 2897
rect 1711 2893 1715 2897
rect 1863 2888 1867 2892
rect 2955 2887 2959 2891
rect 3575 2888 3579 2892
rect 111 2880 115 2884
rect 235 2875 239 2879
rect 779 2875 783 2879
rect 1163 2879 1167 2883
rect 1823 2880 1827 2884
rect 1651 2875 1655 2879
rect 1863 2871 1867 2875
rect 3575 2871 3579 2875
rect 111 2863 115 2867
rect 1823 2863 1827 2867
rect 2887 2861 2891 2865
rect 3191 2861 3195 2865
rect 3479 2861 3483 2865
rect 135 2853 139 2857
rect 311 2853 315 2857
rect 511 2853 515 2857
rect 703 2853 707 2857
rect 887 2853 891 2857
rect 1063 2853 1067 2857
rect 1231 2853 1235 2857
rect 1391 2853 1395 2857
rect 1543 2853 1547 2857
rect 1703 2853 1707 2857
rect 3499 2855 3503 2859
rect 179 2847 183 2851
rect 1291 2847 1295 2851
rect 2831 2839 2835 2843
rect 2919 2839 2923 2843
rect 3007 2839 3011 2843
rect 3095 2839 3099 2843
rect 159 2827 163 2831
rect 319 2827 323 2831
rect 487 2827 491 2831
rect 655 2827 659 2831
rect 823 2827 827 2831
rect 975 2827 979 2831
rect 1127 2827 1131 2831
rect 1271 2827 1275 2831
rect 1415 2827 1419 2831
rect 1559 2827 1563 2831
rect 1863 2829 1867 2833
rect 3163 2831 3167 2835
rect 3575 2829 3579 2833
rect 111 2817 115 2821
rect 903 2819 907 2823
rect 1483 2819 1487 2823
rect 1823 2817 1827 2821
rect 1863 2812 1867 2816
rect 2899 2815 2903 2819
rect 2987 2815 2991 2819
rect 3075 2815 3079 2819
rect 3575 2812 3579 2816
rect 111 2800 115 2804
rect 251 2803 255 2807
rect 387 2803 391 2807
rect 1823 2800 1827 2804
rect 2839 2799 2843 2803
rect 2927 2799 2931 2803
rect 3015 2799 3019 2803
rect 3103 2799 3107 2803
rect 167 2787 171 2791
rect 327 2787 331 2791
rect 495 2787 499 2791
rect 663 2787 667 2791
rect 831 2787 835 2791
rect 983 2787 987 2791
rect 1135 2787 1139 2791
rect 1279 2787 1283 2791
rect 1423 2787 1427 2791
rect 1567 2787 1571 2791
rect 2851 2787 2852 2791
rect 2852 2787 2855 2791
rect 2899 2787 2903 2791
rect 2987 2787 2991 2791
rect 3075 2787 3079 2791
rect 179 2775 180 2779
rect 180 2775 183 2779
rect 251 2775 255 2779
rect 531 2775 535 2779
rect 995 2775 996 2779
rect 996 2775 999 2779
rect 1291 2775 1292 2779
rect 1292 2775 1295 2779
rect 2735 2775 2739 2779
rect 3499 2775 3500 2779
rect 3500 2775 3503 2779
rect 303 2755 307 2759
rect 387 2755 391 2759
rect 651 2755 655 2759
rect 2671 2765 2675 2769
rect 2807 2765 2811 2769
rect 2967 2765 2971 2769
rect 3143 2765 3147 2769
rect 3327 2765 3331 2769
rect 3487 2765 3491 2769
rect 1863 2752 1867 2756
rect 207 2745 211 2749
rect 335 2745 339 2749
rect 471 2745 475 2749
rect 607 2745 611 2749
rect 751 2745 755 2749
rect 887 2745 891 2749
rect 111 2732 115 2736
rect 303 2727 307 2731
rect 531 2731 535 2735
rect 3575 2752 3579 2756
rect 1023 2745 1027 2749
rect 1151 2745 1155 2749
rect 1287 2745 1291 2749
rect 1423 2745 1427 2749
rect 3259 2747 3263 2751
rect 1823 2732 1827 2736
rect 1863 2735 1867 2739
rect 3575 2735 3579 2739
rect 2663 2725 2667 2729
rect 2799 2725 2803 2729
rect 2959 2725 2963 2729
rect 3135 2725 3139 2729
rect 3319 2725 3323 2729
rect 3479 2725 3483 2729
rect 111 2715 115 2719
rect 1823 2715 1827 2719
rect 3499 2719 3503 2723
rect 199 2705 203 2709
rect 327 2705 331 2709
rect 463 2705 467 2709
rect 599 2705 603 2709
rect 743 2705 747 2709
rect 879 2705 883 2709
rect 1015 2705 1019 2709
rect 1143 2705 1147 2709
rect 1279 2705 1283 2709
rect 1415 2705 1419 2709
rect 235 2699 239 2703
rect 1179 2699 1183 2703
rect 1887 2703 1891 2707
rect 1975 2703 1979 2707
rect 2063 2703 2067 2707
rect 2151 2703 2155 2707
rect 2239 2703 2243 2707
rect 2327 2703 2331 2707
rect 2415 2703 2419 2707
rect 2503 2703 2507 2707
rect 2591 2703 2595 2707
rect 2679 2703 2683 2707
rect 2767 2703 2771 2707
rect 2855 2703 2859 2707
rect 2943 2703 2947 2707
rect 3031 2703 3035 2707
rect 3119 2703 3123 2707
rect 3207 2703 3211 2707
rect 3295 2703 3299 2707
rect 3391 2703 3395 2707
rect 3479 2703 3483 2707
rect 1863 2693 1867 2697
rect 3363 2695 3367 2699
rect 3575 2693 3579 2697
rect 215 2679 219 2683
rect 335 2679 339 2683
rect 463 2679 467 2683
rect 583 2679 587 2683
rect 703 2679 707 2683
rect 823 2679 827 2683
rect 935 2679 939 2683
rect 1047 2679 1051 2683
rect 1159 2679 1163 2683
rect 1271 2679 1275 2683
rect 1863 2676 1867 2680
rect 2043 2679 2047 2683
rect 3471 2679 3475 2683
rect 111 2669 115 2673
rect 651 2671 655 2675
rect 3575 2676 3579 2680
rect 1227 2671 1231 2675
rect 1823 2669 1827 2673
rect 1895 2663 1899 2667
rect 1983 2663 1987 2667
rect 2071 2663 2075 2667
rect 2159 2663 2163 2667
rect 2247 2663 2251 2667
rect 2335 2663 2339 2667
rect 2423 2663 2427 2667
rect 2511 2663 2515 2667
rect 2599 2663 2603 2667
rect 2687 2663 2691 2667
rect 2775 2663 2779 2667
rect 2863 2663 2867 2667
rect 2951 2663 2955 2667
rect 3039 2663 3043 2667
rect 3127 2663 3131 2667
rect 3215 2663 3219 2667
rect 3303 2663 3307 2667
rect 3399 2663 3403 2667
rect 3487 2663 3491 2667
rect 111 2652 115 2656
rect 815 2655 819 2659
rect 1139 2655 1143 2659
rect 1823 2652 1827 2656
rect 1951 2651 1955 2655
rect 2043 2651 2047 2655
rect 3499 2651 3500 2655
rect 3500 2651 3503 2655
rect 223 2639 227 2643
rect 343 2639 347 2643
rect 471 2639 475 2643
rect 591 2639 595 2643
rect 711 2639 715 2643
rect 831 2639 835 2643
rect 943 2639 947 2643
rect 1055 2639 1059 2643
rect 1167 2639 1171 2643
rect 1279 2639 1283 2643
rect 235 2627 236 2631
rect 236 2627 239 2631
rect 843 2627 844 2631
rect 844 2627 847 2631
rect 1179 2627 1180 2631
rect 1180 2627 1183 2631
rect 483 2611 484 2615
rect 484 2611 487 2615
rect 2499 2627 2503 2631
rect 3079 2627 3083 2631
rect 3167 2619 3168 2623
rect 3168 2619 3171 2623
rect 815 2611 819 2615
rect 1139 2611 1143 2615
rect 2159 2609 2163 2613
rect 2279 2609 2283 2613
rect 2415 2609 2419 2613
rect 2551 2609 2555 2613
rect 2695 2609 2699 2613
rect 2847 2609 2851 2613
rect 2999 2609 3003 2613
rect 3159 2609 3163 2613
rect 471 2601 475 2605
rect 559 2601 563 2605
rect 647 2601 651 2605
rect 735 2601 739 2605
rect 823 2601 827 2605
rect 911 2601 915 2605
rect 999 2601 1003 2605
rect 1087 2601 1091 2605
rect 1175 2601 1179 2605
rect 1263 2601 1267 2605
rect 1863 2596 1867 2600
rect 111 2588 115 2592
rect 1823 2588 1827 2592
rect 2643 2591 2647 2595
rect 3575 2596 3579 2600
rect 3079 2591 3083 2595
rect 1863 2579 1867 2583
rect 3575 2579 3579 2583
rect 111 2571 115 2575
rect 715 2571 719 2575
rect 463 2561 467 2565
rect 551 2561 555 2565
rect 639 2561 643 2565
rect 727 2561 731 2565
rect 815 2561 819 2565
rect 903 2561 907 2565
rect 991 2561 995 2565
rect 955 2555 959 2559
rect 1823 2571 1827 2575
rect 2151 2569 2155 2573
rect 2271 2569 2275 2573
rect 2407 2569 2411 2573
rect 2543 2569 2547 2573
rect 2687 2569 2691 2573
rect 2839 2569 2843 2573
rect 2991 2569 2995 2573
rect 3151 2569 3155 2573
rect 1079 2561 1083 2565
rect 1167 2561 1171 2565
rect 1255 2561 1259 2565
rect 3019 2563 3023 2567
rect 2103 2547 2107 2551
rect 2199 2547 2203 2551
rect 2311 2547 2315 2551
rect 2431 2547 2435 2551
rect 2559 2547 2563 2551
rect 2695 2547 2699 2551
rect 2847 2547 2851 2551
rect 2999 2547 3003 2551
rect 3159 2547 3163 2551
rect 3327 2547 3331 2551
rect 3479 2547 3483 2551
rect 1863 2537 1867 2541
rect 2499 2539 2503 2543
rect 495 2531 499 2535
rect 583 2531 587 2535
rect 671 2531 675 2535
rect 759 2531 763 2535
rect 847 2531 851 2535
rect 935 2531 939 2535
rect 1023 2531 1027 2535
rect 1111 2531 1115 2535
rect 1199 2531 1203 2535
rect 1287 2531 1291 2535
rect 3167 2535 3171 2539
rect 3575 2537 3579 2541
rect 111 2521 115 2525
rect 483 2523 487 2527
rect 839 2523 843 2527
rect 1267 2523 1271 2527
rect 1823 2521 1827 2525
rect 1863 2520 1867 2524
rect 2627 2523 2631 2527
rect 2763 2523 2767 2527
rect 2915 2523 2919 2527
rect 3227 2523 3231 2527
rect 3575 2520 3579 2524
rect 111 2504 115 2508
rect 563 2507 567 2511
rect 1823 2504 1827 2508
rect 2111 2507 2115 2511
rect 2207 2507 2211 2511
rect 2319 2507 2323 2511
rect 2439 2507 2443 2511
rect 2567 2507 2571 2511
rect 2703 2507 2707 2511
rect 2855 2507 2859 2511
rect 3007 2507 3011 2511
rect 3167 2507 3171 2511
rect 3335 2507 3339 2511
rect 3487 2507 3491 2511
rect 503 2491 507 2495
rect 591 2491 595 2495
rect 679 2491 683 2495
rect 767 2491 771 2495
rect 855 2491 859 2495
rect 943 2491 947 2495
rect 1031 2491 1035 2495
rect 1119 2491 1123 2495
rect 1207 2491 1211 2495
rect 1295 2491 1299 2495
rect 2763 2495 2767 2499
rect 2915 2495 2919 2499
rect 3019 2495 3020 2499
rect 3020 2495 3023 2499
rect 3227 2495 3231 2499
rect 3355 2495 3359 2499
rect 3471 2495 3475 2499
rect 563 2479 567 2483
rect 583 2479 587 2483
rect 715 2479 719 2483
rect 955 2479 956 2483
rect 956 2479 959 2483
rect 2099 2479 2100 2483
rect 2100 2479 2103 2483
rect 2623 2479 2627 2483
rect 3303 2479 3304 2483
rect 3304 2479 3307 2483
rect 2087 2469 2091 2473
rect 2183 2469 2187 2473
rect 2287 2469 2291 2473
rect 2407 2469 2411 2473
rect 2543 2469 2547 2473
rect 2703 2469 2707 2473
rect 2887 2469 2891 2473
rect 3087 2469 3091 2473
rect 3295 2469 3299 2473
rect 3487 2469 3491 2473
rect 415 2459 419 2463
rect 731 2463 732 2467
rect 732 2463 735 2467
rect 839 2463 843 2467
rect 979 2463 980 2467
rect 980 2463 983 2467
rect 1147 2463 1151 2467
rect 359 2453 363 2457
rect 471 2453 475 2457
rect 591 2453 595 2457
rect 719 2453 723 2457
rect 847 2453 851 2457
rect 967 2453 971 2457
rect 1087 2453 1091 2457
rect 1207 2453 1211 2457
rect 1335 2453 1339 2457
rect 1463 2453 1467 2457
rect 1863 2456 1867 2460
rect 3355 2455 3359 2459
rect 3575 2456 3579 2460
rect 111 2440 115 2444
rect 583 2435 587 2439
rect 787 2435 791 2439
rect 1147 2439 1151 2443
rect 1823 2440 1827 2444
rect 1863 2439 1867 2443
rect 2955 2439 2959 2443
rect 3575 2439 3579 2443
rect 2079 2429 2083 2433
rect 2175 2429 2179 2433
rect 2279 2429 2283 2433
rect 2399 2429 2403 2433
rect 2535 2429 2539 2433
rect 2695 2429 2699 2433
rect 2879 2429 2883 2433
rect 3079 2429 3083 2433
rect 3287 2429 3291 2433
rect 3479 2429 3483 2433
rect 111 2423 115 2427
rect 1403 2423 1407 2427
rect 1823 2423 1827 2427
rect 3499 2423 3503 2427
rect 351 2413 355 2417
rect 463 2413 467 2417
rect 583 2413 587 2417
rect 711 2413 715 2417
rect 839 2413 843 2417
rect 959 2413 963 2417
rect 1079 2413 1083 2417
rect 1199 2413 1203 2417
rect 1327 2413 1331 2417
rect 1455 2413 1459 2417
rect 2611 2415 2615 2419
rect 2955 2415 2959 2419
rect 491 2407 495 2411
rect 1951 2403 1955 2407
rect 2063 2403 2067 2407
rect 2183 2403 2187 2407
rect 2311 2403 2315 2407
rect 2447 2403 2451 2407
rect 2591 2403 2595 2407
rect 2751 2403 2755 2407
rect 2927 2403 2931 2407
rect 3111 2403 3115 2407
rect 3303 2403 3307 2407
rect 3479 2403 3483 2407
rect 1863 2393 1867 2397
rect 2379 2395 2383 2399
rect 3019 2395 3023 2399
rect 3295 2395 3299 2399
rect 3575 2393 3579 2397
rect 135 2387 139 2391
rect 287 2387 291 2391
rect 471 2387 475 2391
rect 663 2387 667 2391
rect 847 2387 851 2391
rect 1031 2387 1035 2391
rect 1207 2387 1211 2391
rect 1375 2387 1379 2391
rect 1543 2387 1547 2391
rect 1711 2387 1715 2391
rect 111 2377 115 2381
rect 203 2379 207 2383
rect 731 2379 735 2383
rect 1823 2377 1827 2381
rect 1863 2376 1867 2380
rect 3575 2376 3579 2380
rect 111 2360 115 2364
rect 363 2363 367 2367
rect 731 2363 735 2367
rect 1779 2363 1783 2367
rect 1823 2360 1827 2364
rect 1959 2363 1963 2367
rect 2071 2363 2075 2367
rect 2191 2363 2195 2367
rect 2319 2363 2323 2367
rect 2455 2363 2459 2367
rect 2599 2363 2603 2367
rect 2759 2363 2763 2367
rect 2935 2363 2939 2367
rect 3119 2363 3123 2367
rect 3311 2363 3315 2367
rect 3487 2363 3491 2367
rect 143 2347 147 2351
rect 295 2347 299 2351
rect 479 2347 483 2351
rect 671 2347 675 2351
rect 855 2347 859 2351
rect 1039 2347 1043 2351
rect 1215 2347 1219 2351
rect 1383 2347 1387 2351
rect 1551 2347 1555 2351
rect 1719 2347 1723 2351
rect 2047 2351 2051 2355
rect 2611 2351 2612 2355
rect 2612 2351 2615 2355
rect 3499 2351 3500 2355
rect 3500 2351 3503 2355
rect 203 2335 207 2339
rect 363 2335 367 2339
rect 491 2335 492 2339
rect 492 2335 495 2339
rect 731 2335 735 2339
rect 847 2335 851 2339
rect 1095 2335 1099 2339
rect 1951 2331 1955 2335
rect 3019 2339 3023 2343
rect 2875 2331 2879 2335
rect 227 2319 231 2323
rect 491 2319 492 2323
rect 492 2319 495 2323
rect 1151 2319 1155 2323
rect 143 2309 147 2313
rect 295 2309 299 2313
rect 479 2309 483 2313
rect 671 2309 675 2313
rect 863 2309 867 2313
rect 1055 2309 1059 2313
rect 111 2296 115 2300
rect 227 2291 231 2295
rect 1651 2319 1655 2323
rect 1779 2319 1783 2323
rect 1895 2321 1899 2325
rect 2007 2321 2011 2325
rect 2159 2321 2163 2325
rect 2311 2321 2315 2325
rect 2463 2321 2467 2325
rect 2615 2321 2619 2325
rect 2775 2321 2779 2325
rect 2943 2321 2947 2325
rect 3111 2321 3115 2325
rect 3287 2321 3291 2325
rect 3471 2321 3475 2325
rect 1231 2309 1235 2313
rect 1407 2309 1411 2313
rect 1583 2309 1587 2313
rect 1735 2309 1739 2313
rect 1863 2308 1867 2312
rect 2403 2303 2407 2307
rect 2875 2307 2879 2311
rect 3575 2308 3579 2312
rect 1823 2296 1827 2300
rect 847 2291 851 2295
rect 1339 2291 1343 2295
rect 1651 2291 1655 2295
rect 1863 2291 1867 2295
rect 111 2279 115 2283
rect 1319 2279 1323 2283
rect 1823 2279 1827 2283
rect 1887 2281 1891 2285
rect 1999 2281 2003 2285
rect 2151 2281 2155 2285
rect 2303 2281 2307 2285
rect 2455 2281 2459 2285
rect 2607 2281 2611 2285
rect 2767 2281 2771 2285
rect 2935 2281 2939 2285
rect 3103 2281 3107 2285
rect 2799 2275 2803 2279
rect 3575 2291 3579 2295
rect 3279 2281 3283 2285
rect 3463 2281 3467 2285
rect 3499 2275 3503 2279
rect 135 2269 139 2273
rect 287 2269 291 2273
rect 471 2269 475 2273
rect 663 2269 667 2273
rect 855 2269 859 2273
rect 1047 2269 1051 2273
rect 1223 2269 1227 2273
rect 1399 2269 1403 2273
rect 1575 2269 1579 2273
rect 1727 2269 1731 2273
rect 155 2263 159 2267
rect 1887 2255 1891 2259
rect 2023 2255 2027 2259
rect 2199 2255 2203 2259
rect 2383 2255 2387 2259
rect 2567 2255 2571 2259
rect 2743 2255 2747 2259
rect 2911 2255 2915 2259
rect 3079 2255 3083 2259
rect 3239 2255 3243 2259
rect 3407 2255 3411 2259
rect 1863 2245 1867 2249
rect 2479 2247 2483 2251
rect 3147 2247 3151 2251
rect 3575 2245 3579 2249
rect 135 2239 139 2243
rect 255 2239 259 2243
rect 407 2239 411 2243
rect 559 2239 563 2243
rect 719 2239 723 2243
rect 871 2239 875 2243
rect 1015 2239 1019 2243
rect 1159 2239 1163 2243
rect 1303 2239 1307 2243
rect 1455 2239 1459 2243
rect 111 2229 115 2233
rect 375 2231 379 2235
rect 491 2231 495 2235
rect 1399 2231 1403 2235
rect 1823 2229 1827 2233
rect 1863 2228 1867 2232
rect 3575 2228 3579 2232
rect 111 2212 115 2216
rect 627 2215 631 2219
rect 1083 2215 1087 2219
rect 1099 2215 1103 2219
rect 1823 2212 1827 2216
rect 1895 2215 1899 2219
rect 2031 2215 2035 2219
rect 2207 2215 2211 2219
rect 2391 2215 2395 2219
rect 2575 2215 2579 2219
rect 2751 2215 2755 2219
rect 2919 2215 2923 2219
rect 3087 2215 3091 2219
rect 3247 2215 3251 2219
rect 3415 2215 3419 2219
rect 143 2199 147 2203
rect 263 2199 267 2203
rect 415 2199 419 2203
rect 567 2199 571 2203
rect 727 2199 731 2203
rect 879 2199 883 2203
rect 1023 2199 1027 2203
rect 1167 2199 1171 2203
rect 1311 2199 1315 2203
rect 1463 2199 1467 2203
rect 2007 2203 2011 2207
rect 2799 2203 2803 2207
rect 3427 2203 3428 2207
rect 3428 2203 3431 2207
rect 155 2187 156 2191
rect 156 2187 159 2191
rect 627 2187 631 2191
rect 891 2187 892 2191
rect 892 2187 895 2191
rect 1191 2187 1195 2191
rect 1319 2187 1320 2191
rect 1320 2187 1323 2191
rect 2771 2187 2772 2191
rect 2772 2187 2775 2191
rect 3499 2187 3500 2191
rect 3500 2187 3503 2191
rect 375 2179 379 2183
rect 899 2179 903 2183
rect 1895 2177 1899 2181
rect 2039 2177 2043 2181
rect 2215 2177 2219 2181
rect 2399 2177 2403 2181
rect 2583 2177 2587 2181
rect 2759 2177 2763 2181
rect 2919 2177 2923 2181
rect 3071 2177 3075 2181
rect 3215 2177 3219 2181
rect 3359 2177 3363 2181
rect 3487 2177 3491 2181
rect 1083 2171 1087 2175
rect 215 2161 219 2165
rect 311 2161 315 2165
rect 415 2161 419 2165
rect 491 2163 495 2167
rect 519 2161 523 2165
rect 623 2161 627 2165
rect 727 2161 731 2165
rect 831 2161 835 2165
rect 943 2161 947 2165
rect 1055 2161 1059 2165
rect 1167 2161 1171 2165
rect 1863 2164 1867 2168
rect 2507 2159 2511 2163
rect 3575 2164 3579 2168
rect 111 2148 115 2152
rect 899 2143 903 2147
rect 1823 2148 1827 2152
rect 1863 2147 1867 2151
rect 3335 2147 3339 2151
rect 3575 2147 3579 2151
rect 1887 2137 1891 2141
rect 2031 2137 2035 2141
rect 2207 2137 2211 2141
rect 2391 2137 2395 2141
rect 2575 2137 2579 2141
rect 2751 2137 2755 2141
rect 2911 2137 2915 2141
rect 3063 2137 3067 2141
rect 3207 2137 3211 2141
rect 3351 2137 3355 2141
rect 3479 2137 3483 2141
rect 111 2131 115 2135
rect 1823 2131 1827 2135
rect 3499 2131 3503 2135
rect 207 2121 211 2125
rect 303 2121 307 2125
rect 407 2121 411 2125
rect 511 2121 515 2125
rect 615 2121 619 2125
rect 719 2121 723 2125
rect 823 2121 827 2125
rect 935 2121 939 2125
rect 1047 2121 1051 2125
rect 1159 2121 1163 2125
rect 339 2115 343 2119
rect 851 2115 855 2119
rect 1887 2111 1891 2115
rect 2023 2111 2027 2115
rect 2199 2111 2203 2115
rect 2375 2111 2379 2115
rect 2551 2111 2555 2115
rect 2719 2111 2723 2115
rect 2879 2111 2883 2115
rect 3031 2111 3035 2115
rect 3175 2111 3179 2115
rect 3319 2111 3323 2115
rect 3471 2111 3475 2115
rect 1863 2101 1867 2105
rect 2479 2103 2483 2107
rect 3427 2103 3431 2107
rect 3575 2101 3579 2105
rect 319 2091 323 2095
rect 423 2091 427 2095
rect 527 2091 531 2095
rect 631 2091 635 2095
rect 735 2091 739 2095
rect 831 2091 835 2095
rect 927 2091 931 2095
rect 1031 2091 1035 2095
rect 1135 2091 1139 2095
rect 1239 2091 1243 2095
rect 111 2081 115 2085
rect 491 2083 495 2087
rect 1823 2081 1827 2085
rect 1863 2084 1867 2088
rect 1955 2087 1959 2091
rect 2619 2087 2623 2091
rect 2791 2087 2795 2091
rect 2947 2087 2951 2091
rect 3099 2087 3103 2091
rect 3243 2087 3247 2091
rect 3575 2084 3579 2088
rect 111 2064 115 2068
rect 1207 2067 1211 2071
rect 1215 2067 1219 2071
rect 1895 2071 1899 2075
rect 2031 2071 2035 2075
rect 2207 2071 2211 2075
rect 2383 2071 2387 2075
rect 2559 2071 2563 2075
rect 2727 2071 2731 2075
rect 2887 2071 2891 2075
rect 3039 2071 3043 2075
rect 3183 2071 3187 2075
rect 3327 2071 3331 2075
rect 3479 2071 3483 2075
rect 1823 2064 1827 2068
rect 1955 2059 1959 2063
rect 2039 2059 2040 2063
rect 2040 2059 2043 2063
rect 2215 2059 2216 2063
rect 2216 2059 2219 2063
rect 2791 2059 2795 2063
rect 2947 2059 2951 2063
rect 3099 2059 3103 2063
rect 3243 2059 3247 2063
rect 3335 2059 3336 2063
rect 3336 2059 3339 2063
rect 3471 2059 3475 2063
rect 327 2051 331 2055
rect 431 2051 435 2055
rect 535 2051 539 2055
rect 639 2051 643 2055
rect 743 2051 747 2055
rect 839 2051 843 2055
rect 935 2051 939 2055
rect 1039 2051 1043 2055
rect 1143 2051 1147 2055
rect 1247 2051 1251 2055
rect 339 2039 340 2043
rect 340 2039 343 2043
rect 791 2039 795 2043
rect 851 2039 852 2043
rect 852 2039 855 2043
rect 1207 2039 1211 2043
rect 615 2019 619 2023
rect 651 2019 655 2023
rect 783 2019 787 2023
rect 1215 2027 1219 2031
rect 1895 2029 1899 2033
rect 1959 2039 1963 2043
rect 2091 2039 2095 2043
rect 2363 2039 2367 2043
rect 2451 2039 2452 2043
rect 2452 2039 2455 2043
rect 2619 2039 2623 2043
rect 2683 2039 2687 2043
rect 2871 2039 2875 2043
rect 3223 2039 3227 2043
rect 3499 2039 3500 2043
rect 3500 2039 3503 2043
rect 2007 2027 2011 2031
rect 2015 2029 2019 2033
rect 2151 2029 2155 2033
rect 2295 2029 2299 2033
rect 2439 2029 2443 2033
rect 2591 2029 2595 2033
rect 2759 2029 2763 2033
rect 2935 2029 2939 2033
rect 3119 2029 3123 2033
rect 3311 2029 3315 2033
rect 3487 2029 3491 2033
rect 1075 2019 1079 2023
rect 1319 2019 1323 2023
rect 1443 2019 1447 2023
rect 1863 2016 1867 2020
rect 1959 2015 1963 2019
rect 2091 2015 2095 2019
rect 2215 2015 2219 2019
rect 215 2009 219 2013
rect 391 2009 395 2013
rect 559 2009 563 2013
rect 719 2009 723 2013
rect 863 2009 867 2013
rect 999 2009 1003 2013
rect 1127 2009 1131 2013
rect 1247 2009 1251 2013
rect 1367 2009 1371 2013
rect 1495 2009 1499 2013
rect 2223 2011 2227 2015
rect 2363 2011 2367 2015
rect 2683 2015 2687 2019
rect 2871 2015 2875 2019
rect 3223 2015 3227 2019
rect 3575 2016 3579 2020
rect 111 1996 115 2000
rect 651 1995 655 1999
rect 783 1995 787 1999
rect 791 1991 795 1995
rect 1075 1995 1079 1999
rect 1319 1995 1323 1999
rect 1443 1995 1447 1999
rect 1823 1996 1827 2000
rect 1863 1999 1867 2003
rect 3311 1999 3315 2003
rect 3575 1999 3579 2003
rect 1887 1989 1891 1993
rect 2007 1989 2011 1993
rect 2143 1989 2147 1993
rect 2287 1989 2291 1993
rect 2431 1989 2435 1993
rect 2583 1989 2587 1993
rect 2751 1989 2755 1993
rect 2927 1989 2931 1993
rect 3111 1989 3115 1993
rect 3303 1989 3307 1993
rect 3479 1989 3483 1993
rect 111 1979 115 1983
rect 155 1979 159 1983
rect 207 1969 211 1973
rect 383 1969 387 1973
rect 551 1969 555 1973
rect 711 1969 715 1973
rect 855 1969 859 1973
rect 991 1969 995 1973
rect 1119 1969 1123 1973
rect 1239 1969 1243 1973
rect 1359 1969 1363 1973
rect 1135 1963 1139 1967
rect 1823 1979 1827 1983
rect 3527 1983 3528 1987
rect 3528 1983 3531 1987
rect 1487 1969 1491 1973
rect 2023 1963 2027 1967
rect 2111 1963 2115 1967
rect 2199 1963 2203 1967
rect 2287 1963 2291 1967
rect 2383 1963 2387 1967
rect 2503 1963 2507 1967
rect 2655 1963 2659 1967
rect 2839 1963 2843 1967
rect 3047 1963 3051 1967
rect 3271 1963 3275 1967
rect 3479 1963 3483 1967
rect 1863 1953 1867 1957
rect 2451 1955 2455 1959
rect 2571 1955 2575 1959
rect 3575 1953 3579 1957
rect 135 1939 139 1943
rect 311 1939 315 1943
rect 519 1939 523 1943
rect 719 1939 723 1943
rect 911 1939 915 1943
rect 1095 1939 1099 1943
rect 1263 1939 1267 1943
rect 1423 1939 1427 1943
rect 1583 1939 1587 1943
rect 1727 1939 1731 1943
rect 1863 1936 1867 1940
rect 2647 1939 2651 1943
rect 2723 1939 2727 1943
rect 2907 1939 2911 1943
rect 3115 1939 3119 1943
rect 111 1929 115 1933
rect 379 1931 383 1935
rect 615 1931 619 1935
rect 3575 1936 3579 1940
rect 1719 1931 1723 1935
rect 1823 1929 1827 1933
rect 2031 1923 2035 1927
rect 2119 1923 2123 1927
rect 2207 1923 2211 1927
rect 2295 1923 2299 1927
rect 2391 1923 2395 1927
rect 2511 1923 2515 1927
rect 2663 1923 2667 1927
rect 2847 1923 2851 1927
rect 3055 1923 3059 1927
rect 3279 1923 3283 1927
rect 3487 1923 3491 1927
rect 111 1912 115 1916
rect 243 1915 247 1919
rect 787 1915 791 1919
rect 1823 1912 1827 1916
rect 2043 1911 2044 1915
rect 2044 1911 2047 1915
rect 2571 1911 2575 1915
rect 2723 1911 2727 1915
rect 2907 1911 2911 1915
rect 3115 1911 3119 1915
rect 3311 1911 3315 1915
rect 3527 1911 3531 1915
rect 143 1899 147 1903
rect 319 1899 323 1903
rect 527 1899 531 1903
rect 727 1899 731 1903
rect 919 1899 923 1903
rect 1103 1899 1107 1903
rect 1271 1899 1275 1903
rect 1431 1899 1435 1903
rect 1591 1899 1595 1903
rect 1735 1899 1739 1903
rect 155 1887 156 1891
rect 156 1887 159 1891
rect 243 1887 247 1891
rect 787 1887 791 1891
rect 947 1887 951 1891
rect 1135 1887 1139 1891
rect 2243 1891 2247 1895
rect 2331 1891 2335 1895
rect 2419 1891 2423 1895
rect 2535 1891 2536 1895
rect 2536 1891 2539 1895
rect 2647 1891 2648 1895
rect 2648 1891 2651 1895
rect 2891 1891 2895 1895
rect 2175 1881 2179 1885
rect 2263 1881 2267 1885
rect 2351 1881 2355 1885
rect 2439 1881 2443 1885
rect 2527 1881 2531 1885
rect 2639 1881 2643 1885
rect 2775 1881 2779 1885
rect 2935 1881 2939 1885
rect 3119 1881 3123 1885
rect 3311 1881 3315 1885
rect 3487 1881 3491 1885
rect 235 1867 239 1871
rect 379 1867 383 1871
rect 1135 1867 1139 1871
rect 1719 1867 1720 1871
rect 1720 1867 1723 1871
rect 1863 1868 1867 1872
rect 143 1857 147 1861
rect 311 1857 315 1861
rect 511 1857 515 1861
rect 635 1859 639 1863
rect 2043 1863 2047 1867
rect 2243 1863 2247 1867
rect 2331 1863 2335 1867
rect 2419 1863 2423 1867
rect 2891 1867 2895 1871
rect 3575 1868 3579 1872
rect 703 1857 707 1861
rect 887 1857 891 1861
rect 1063 1857 1067 1861
rect 1231 1857 1235 1861
rect 1391 1857 1395 1861
rect 1551 1857 1555 1861
rect 1711 1857 1715 1861
rect 1863 1851 1867 1855
rect 3199 1851 3203 1855
rect 3575 1851 3579 1855
rect 111 1844 115 1848
rect 235 1839 239 1843
rect 947 1843 951 1847
rect 1823 1844 1827 1848
rect 1299 1839 1303 1843
rect 2167 1841 2171 1845
rect 2255 1841 2259 1845
rect 2343 1841 2347 1845
rect 2431 1841 2435 1845
rect 2519 1841 2523 1845
rect 2631 1841 2635 1845
rect 2767 1841 2771 1845
rect 2927 1841 2931 1845
rect 3111 1841 3115 1845
rect 3303 1841 3307 1845
rect 3479 1841 3483 1845
rect 3499 1835 3503 1839
rect 111 1827 115 1831
rect 1299 1827 1303 1831
rect 1823 1827 1827 1831
rect 135 1817 139 1821
rect 303 1817 307 1821
rect 503 1817 507 1821
rect 695 1817 699 1821
rect 879 1817 883 1821
rect 1055 1817 1059 1821
rect 1223 1817 1227 1821
rect 1383 1817 1387 1821
rect 1543 1817 1547 1821
rect 1703 1817 1707 1821
rect 155 1811 159 1815
rect 2319 1815 2323 1819
rect 2439 1815 2443 1819
rect 2559 1815 2563 1819
rect 2679 1815 2683 1819
rect 2799 1815 2803 1819
rect 2919 1815 2923 1819
rect 3047 1815 3051 1819
rect 3183 1815 3187 1819
rect 3319 1815 3323 1819
rect 3463 1815 3467 1819
rect 1863 1805 1867 1809
rect 2535 1807 2539 1811
rect 3471 1803 3475 1807
rect 3575 1805 3579 1809
rect 135 1787 139 1791
rect 263 1787 267 1791
rect 415 1787 419 1791
rect 567 1787 571 1791
rect 719 1787 723 1791
rect 863 1787 867 1791
rect 1007 1787 1011 1791
rect 1143 1787 1147 1791
rect 1279 1787 1283 1791
rect 1423 1787 1427 1791
rect 1863 1788 1867 1792
rect 2507 1791 2511 1795
rect 2627 1791 2631 1795
rect 3391 1791 3395 1795
rect 3575 1788 3579 1792
rect 111 1777 115 1781
rect 635 1779 639 1783
rect 1347 1779 1351 1783
rect 1823 1777 1827 1781
rect 2327 1775 2331 1779
rect 2447 1775 2451 1779
rect 2567 1775 2571 1779
rect 2687 1775 2691 1779
rect 2807 1775 2811 1779
rect 2927 1775 2931 1779
rect 3055 1775 3059 1779
rect 3191 1775 3195 1779
rect 3327 1775 3331 1779
rect 3471 1775 3475 1779
rect 111 1760 115 1764
rect 331 1763 335 1767
rect 787 1763 791 1767
rect 931 1763 935 1767
rect 1075 1763 1079 1767
rect 1823 1760 1827 1764
rect 2627 1763 2631 1767
rect 2723 1763 2727 1767
rect 2819 1763 2820 1767
rect 2820 1763 2823 1767
rect 3463 1763 3467 1767
rect 2507 1755 2511 1759
rect 143 1747 147 1751
rect 271 1747 275 1751
rect 423 1747 427 1751
rect 575 1747 579 1751
rect 727 1747 731 1751
rect 871 1747 875 1751
rect 1015 1747 1019 1751
rect 1151 1747 1155 1751
rect 1287 1747 1291 1751
rect 1431 1747 1435 1751
rect 2307 1743 2308 1747
rect 2308 1743 2311 1747
rect 2715 1743 2719 1747
rect 2967 1743 2971 1747
rect 3043 1743 3047 1747
rect 3391 1743 3392 1747
rect 3392 1743 3395 1747
rect 3499 1743 3500 1747
rect 3500 1743 3503 1747
rect 155 1735 156 1739
rect 156 1735 159 1739
rect 415 1735 419 1739
rect 931 1735 935 1739
rect 1075 1735 1079 1739
rect 1299 1735 1300 1739
rect 1300 1735 1303 1739
rect 2295 1733 2299 1737
rect 2407 1733 2411 1737
rect 2527 1733 2531 1737
rect 2655 1733 2659 1737
rect 2775 1733 2779 1737
rect 2895 1733 2899 1737
rect 3015 1733 3019 1737
rect 3135 1733 3139 1737
rect 3255 1733 3259 1737
rect 3383 1733 3387 1737
rect 3487 1733 3491 1737
rect 219 1723 223 1727
rect 331 1723 335 1727
rect 499 1723 503 1727
rect 787 1723 791 1727
rect 1347 1727 1351 1731
rect 1863 1720 1867 1724
rect 2715 1719 2719 1723
rect 143 1713 147 1717
rect 279 1713 283 1717
rect 431 1713 435 1717
rect 583 1713 587 1717
rect 727 1713 731 1717
rect 863 1713 867 1717
rect 991 1713 995 1717
rect 1127 1713 1131 1717
rect 1263 1713 1267 1717
rect 2723 1715 2727 1719
rect 2967 1715 2971 1719
rect 3575 1720 3579 1724
rect 111 1700 115 1704
rect 219 1695 223 1699
rect 415 1695 419 1699
rect 499 1695 503 1699
rect 1823 1700 1827 1704
rect 1863 1703 1867 1707
rect 2855 1703 2859 1707
rect 3335 1703 3339 1707
rect 3575 1703 3579 1707
rect 2287 1693 2291 1697
rect 2399 1693 2403 1697
rect 2519 1693 2523 1697
rect 2647 1693 2651 1697
rect 2767 1693 2771 1697
rect 2887 1693 2891 1697
rect 3007 1693 3011 1697
rect 3127 1693 3131 1697
rect 3247 1693 3251 1697
rect 3375 1693 3379 1697
rect 3479 1693 3483 1697
rect 111 1683 115 1687
rect 1211 1683 1215 1687
rect 1823 1683 1827 1687
rect 3499 1687 3503 1691
rect 135 1673 139 1677
rect 271 1673 275 1677
rect 423 1673 427 1677
rect 575 1673 579 1677
rect 719 1673 723 1677
rect 855 1673 859 1677
rect 983 1673 987 1677
rect 1119 1673 1123 1677
rect 1255 1673 1259 1677
rect 2307 1675 2311 1679
rect 155 1667 159 1671
rect 2143 1667 2147 1671
rect 2247 1667 2251 1671
rect 2367 1667 2371 1671
rect 2503 1667 2507 1671
rect 2647 1667 2651 1671
rect 2807 1667 2811 1671
rect 2975 1667 2979 1671
rect 3143 1667 3147 1671
rect 3319 1667 3323 1671
rect 3479 1667 3483 1671
rect 1863 1657 1867 1661
rect 2955 1659 2959 1663
rect 3043 1659 3047 1663
rect 3575 1657 3579 1661
rect 135 1651 139 1655
rect 263 1651 267 1655
rect 423 1651 427 1655
rect 575 1651 579 1655
rect 727 1651 731 1655
rect 871 1651 875 1655
rect 1007 1651 1011 1655
rect 1143 1651 1147 1655
rect 1279 1651 1283 1655
rect 1415 1651 1419 1655
rect 111 1641 115 1645
rect 203 1643 207 1647
rect 1347 1643 1351 1647
rect 1823 1641 1827 1645
rect 1863 1640 1867 1644
rect 2967 1643 2971 1647
rect 3447 1643 3451 1647
rect 3575 1640 3579 1644
rect 111 1624 115 1628
rect 643 1627 647 1631
rect 1099 1627 1103 1631
rect 1823 1624 1827 1628
rect 2151 1627 2155 1631
rect 2255 1627 2259 1631
rect 2375 1627 2379 1631
rect 2511 1627 2515 1631
rect 2655 1627 2659 1631
rect 2815 1627 2819 1631
rect 2983 1627 2987 1631
rect 3151 1627 3155 1631
rect 3327 1627 3331 1631
rect 3487 1627 3491 1631
rect 143 1611 147 1615
rect 271 1611 275 1615
rect 431 1611 435 1615
rect 583 1611 587 1615
rect 735 1611 739 1615
rect 879 1611 883 1615
rect 1015 1611 1019 1615
rect 1151 1611 1155 1615
rect 1287 1611 1291 1615
rect 1423 1611 1427 1615
rect 2227 1615 2231 1619
rect 2855 1615 2859 1619
rect 2967 1615 2971 1619
rect 3187 1615 3191 1619
rect 3335 1615 3336 1619
rect 3336 1615 3339 1619
rect 3499 1615 3500 1619
rect 3500 1615 3503 1619
rect 155 1599 156 1603
rect 156 1599 159 1603
rect 443 1599 444 1603
rect 444 1599 447 1603
rect 743 1599 744 1603
rect 744 1599 747 1603
rect 891 1599 892 1603
rect 892 1599 895 1603
rect 1099 1599 1103 1603
rect 2019 1603 2020 1607
rect 2020 1603 2023 1607
rect 2955 1603 2956 1607
rect 2956 1603 2959 1607
rect 3327 1599 3331 1603
rect 203 1583 207 1587
rect 751 1591 755 1595
rect 2007 1593 2011 1597
rect 2103 1593 2107 1597
rect 2207 1593 2211 1597
rect 2327 1593 2331 1597
rect 2463 1593 2467 1597
rect 2607 1593 2611 1597
rect 2767 1593 2771 1597
rect 2943 1593 2947 1597
rect 3127 1593 3131 1597
rect 3319 1593 3323 1597
rect 3487 1593 3491 1597
rect 859 1583 860 1587
rect 860 1583 863 1587
rect 1023 1583 1027 1587
rect 1863 1580 1867 1584
rect 167 1573 171 1577
rect 335 1573 339 1577
rect 511 1573 515 1577
rect 679 1573 683 1577
rect 847 1573 851 1577
rect 999 1573 1003 1577
rect 1151 1573 1155 1577
rect 1295 1573 1299 1577
rect 1439 1573 1443 1577
rect 1583 1573 1587 1577
rect 3187 1579 3191 1583
rect 3575 1580 3579 1584
rect 3463 1575 3467 1579
rect 111 1560 115 1564
rect 743 1559 747 1563
rect 751 1555 755 1559
rect 1823 1560 1827 1564
rect 1863 1563 1867 1567
rect 1999 1553 2003 1557
rect 2095 1553 2099 1557
rect 2199 1553 2203 1557
rect 2319 1553 2323 1557
rect 111 1543 115 1547
rect 407 1543 411 1547
rect 1519 1543 1523 1547
rect 1823 1543 1827 1547
rect 2227 1547 2231 1551
rect 2727 1563 2731 1567
rect 3575 1563 3579 1567
rect 2455 1553 2459 1557
rect 2599 1553 2603 1557
rect 2759 1553 2763 1557
rect 2935 1553 2939 1557
rect 3119 1553 3123 1557
rect 3311 1553 3315 1557
rect 3479 1553 3483 1557
rect 159 1533 163 1537
rect 327 1533 331 1537
rect 503 1533 507 1537
rect 671 1533 675 1537
rect 839 1533 843 1537
rect 991 1533 995 1537
rect 1143 1533 1147 1537
rect 1287 1533 1291 1537
rect 1431 1533 1435 1537
rect 1575 1533 1579 1537
rect 1887 1523 1891 1527
rect 1975 1523 1979 1527
rect 2103 1523 2107 1527
rect 2239 1523 2243 1527
rect 2383 1523 2387 1527
rect 2543 1523 2547 1527
rect 2711 1523 2715 1527
rect 2879 1523 2883 1527
rect 3055 1523 3059 1527
rect 3239 1523 3243 1527
rect 3431 1523 3435 1527
rect 1863 1513 1867 1517
rect 2307 1515 2311 1519
rect 3327 1515 3331 1519
rect 3575 1513 3579 1517
rect 215 1507 219 1511
rect 391 1507 395 1511
rect 575 1507 579 1511
rect 759 1507 763 1511
rect 935 1507 939 1511
rect 1095 1507 1099 1511
rect 1255 1507 1259 1511
rect 1407 1507 1411 1511
rect 1559 1507 1563 1511
rect 1711 1507 1715 1511
rect 111 1497 115 1501
rect 859 1499 863 1503
rect 1627 1499 1631 1503
rect 1823 1497 1827 1501
rect 1863 1496 1867 1500
rect 2043 1499 2047 1503
rect 2611 1499 2615 1503
rect 3123 1499 3127 1503
rect 3499 1499 3503 1503
rect 3575 1496 3579 1500
rect 111 1480 115 1484
rect 283 1483 287 1487
rect 291 1483 295 1487
rect 1823 1480 1827 1484
rect 1895 1483 1899 1487
rect 1983 1483 1987 1487
rect 2111 1483 2115 1487
rect 2247 1483 2251 1487
rect 2391 1483 2395 1487
rect 2551 1483 2555 1487
rect 2719 1483 2723 1487
rect 2887 1483 2891 1487
rect 3063 1483 3067 1487
rect 3247 1483 3251 1487
rect 3439 1483 3443 1487
rect 223 1467 227 1471
rect 399 1467 403 1471
rect 583 1467 587 1471
rect 767 1467 771 1471
rect 943 1467 947 1471
rect 1103 1467 1107 1471
rect 1263 1467 1267 1471
rect 1415 1467 1419 1471
rect 1567 1467 1571 1471
rect 1719 1467 1723 1471
rect 1951 1471 1955 1475
rect 2043 1471 2047 1475
rect 2611 1471 2615 1475
rect 2727 1471 2728 1475
rect 2728 1471 2731 1475
rect 2827 1471 2831 1475
rect 3447 1471 3448 1475
rect 3448 1471 3451 1475
rect 291 1455 295 1459
rect 407 1455 408 1459
rect 408 1455 411 1459
rect 739 1455 743 1459
rect 1115 1455 1116 1459
rect 1116 1455 1119 1459
rect 2235 1455 2239 1459
rect 2519 1455 2523 1459
rect 3123 1455 3127 1459
rect 3499 1455 3503 1459
rect 283 1439 287 1443
rect 331 1439 335 1443
rect 691 1439 695 1443
rect 1203 1439 1207 1443
rect 1627 1447 1631 1451
rect 1895 1445 1899 1449
rect 2023 1445 2027 1449
rect 2175 1445 2179 1449
rect 2319 1445 2323 1449
rect 2463 1445 2467 1449
rect 2615 1445 2619 1449
rect 2767 1445 2771 1449
rect 2935 1445 2939 1449
rect 3103 1445 3107 1449
rect 3279 1445 3283 1449
rect 3463 1445 3467 1449
rect 1679 1439 1683 1443
rect 255 1429 259 1433
rect 383 1429 387 1433
rect 519 1429 523 1433
rect 671 1429 675 1433
rect 831 1429 835 1433
rect 991 1429 995 1433
rect 1143 1429 1147 1433
rect 1295 1429 1299 1433
rect 1447 1429 1451 1433
rect 1599 1429 1603 1433
rect 1735 1429 1739 1433
rect 1863 1432 1867 1436
rect 2235 1431 2239 1435
rect 2243 1427 2247 1431
rect 2827 1431 2831 1435
rect 3575 1432 3579 1436
rect 111 1416 115 1420
rect 331 1415 335 1419
rect 1823 1416 1827 1420
rect 1863 1415 1867 1419
rect 2379 1411 2383 1415
rect 2867 1415 2871 1419
rect 3575 1415 3579 1419
rect 1887 1405 1891 1409
rect 2015 1405 2019 1409
rect 2167 1405 2171 1409
rect 2311 1405 2315 1409
rect 2455 1405 2459 1409
rect 2607 1405 2611 1409
rect 2759 1405 2763 1409
rect 2927 1405 2931 1409
rect 3095 1405 3099 1409
rect 3271 1405 3275 1409
rect 3455 1405 3459 1409
rect 111 1399 115 1403
rect 739 1399 743 1403
rect 899 1399 903 1403
rect 1719 1399 1723 1403
rect 1823 1399 1827 1403
rect 3499 1399 3503 1403
rect 247 1389 251 1393
rect 375 1389 379 1393
rect 511 1389 515 1393
rect 663 1389 667 1393
rect 823 1389 827 1393
rect 983 1389 987 1393
rect 1135 1389 1139 1393
rect 1287 1389 1291 1393
rect 1439 1389 1443 1393
rect 1591 1389 1595 1393
rect 1727 1389 1731 1393
rect 543 1383 547 1387
rect 351 1367 355 1371
rect 439 1367 443 1371
rect 527 1367 531 1371
rect 623 1367 627 1371
rect 727 1367 731 1371
rect 847 1367 851 1371
rect 983 1367 987 1371
rect 1127 1367 1131 1371
rect 1279 1367 1283 1371
rect 1431 1367 1435 1371
rect 1591 1367 1595 1371
rect 1727 1367 1731 1371
rect 1887 1371 1891 1375
rect 2143 1371 2147 1375
rect 2391 1371 2395 1375
rect 2623 1371 2627 1375
rect 2847 1371 2851 1375
rect 3063 1371 3067 1375
rect 3271 1371 3275 1375
rect 3479 1371 3483 1375
rect 111 1357 115 1361
rect 691 1359 695 1363
rect 1203 1359 1207 1363
rect 1679 1359 1683 1363
rect 1823 1357 1827 1361
rect 1863 1361 1867 1365
rect 2519 1363 2523 1367
rect 2971 1363 2975 1367
rect 3575 1361 3579 1365
rect 111 1340 115 1344
rect 507 1343 511 1347
rect 515 1343 519 1347
rect 795 1343 799 1347
rect 1823 1340 1827 1344
rect 1863 1344 1867 1348
rect 1871 1347 1875 1351
rect 2463 1347 2467 1351
rect 3575 1344 3579 1348
rect 359 1327 363 1331
rect 447 1327 451 1331
rect 535 1327 539 1331
rect 631 1327 635 1331
rect 735 1327 739 1331
rect 855 1327 859 1331
rect 991 1327 995 1331
rect 1135 1327 1139 1331
rect 1287 1327 1291 1331
rect 1439 1327 1443 1331
rect 1599 1327 1603 1331
rect 1735 1327 1739 1331
rect 1895 1331 1899 1335
rect 2151 1331 2155 1335
rect 2399 1331 2403 1335
rect 2631 1331 2635 1335
rect 2855 1331 2859 1335
rect 3071 1331 3075 1335
rect 3279 1331 3283 1335
rect 3487 1331 3491 1335
rect 367 1315 368 1319
rect 368 1315 371 1319
rect 543 1321 547 1323
rect 543 1319 544 1321
rect 544 1319 547 1321
rect 795 1315 799 1319
rect 899 1315 903 1319
rect 1027 1315 1031 1319
rect 1451 1315 1452 1319
rect 1452 1315 1455 1319
rect 1719 1315 1723 1319
rect 1907 1319 1908 1323
rect 1908 1319 1911 1323
rect 2379 1319 2383 1323
rect 2463 1319 2467 1323
rect 2683 1319 2687 1323
rect 2867 1319 2868 1323
rect 2868 1319 2871 1323
rect 3419 1319 3423 1323
rect 3499 1319 3500 1323
rect 3500 1319 3503 1323
rect 507 1303 511 1307
rect 1059 1303 1063 1307
rect 1231 1303 1235 1307
rect 1395 1303 1399 1307
rect 1543 1303 1544 1307
rect 1544 1303 1547 1307
rect 2031 1307 2035 1311
rect 2231 1307 2235 1311
rect 2719 1307 2723 1311
rect 2815 1307 2819 1311
rect 2971 1307 2972 1311
rect 2972 1307 2975 1311
rect 455 1293 459 1297
rect 543 1293 547 1297
rect 631 1293 635 1297
rect 719 1293 723 1297
rect 831 1293 835 1297
rect 967 1293 971 1297
rect 1135 1293 1139 1297
rect 1327 1293 1331 1297
rect 1535 1293 1539 1297
rect 1735 1293 1739 1297
rect 1927 1297 1931 1301
rect 2111 1297 2115 1301
rect 2287 1297 2291 1301
rect 2455 1297 2459 1301
rect 2623 1297 2627 1301
rect 2791 1297 2795 1301
rect 2959 1297 2963 1301
rect 3135 1297 3139 1301
rect 3319 1297 3323 1301
rect 3487 1297 3491 1301
rect 111 1280 115 1284
rect 1027 1279 1031 1283
rect 1823 1280 1827 1284
rect 1863 1284 1867 1288
rect 1059 1275 1063 1279
rect 1231 1275 1235 1279
rect 1907 1279 1911 1283
rect 1395 1275 1399 1279
rect 2031 1279 2035 1283
rect 2683 1283 2687 1287
rect 2719 1279 2723 1283
rect 3575 1284 3579 1288
rect 111 1263 115 1267
rect 831 1263 835 1267
rect 1627 1263 1631 1267
rect 1823 1263 1827 1267
rect 1863 1267 1867 1271
rect 3575 1267 3579 1271
rect 447 1253 451 1257
rect 535 1253 539 1257
rect 623 1253 627 1257
rect 711 1253 715 1257
rect 823 1253 827 1257
rect 959 1253 963 1257
rect 1127 1253 1131 1257
rect 1319 1253 1323 1257
rect 1527 1253 1531 1257
rect 1727 1253 1731 1257
rect 1919 1257 1923 1261
rect 2103 1257 2107 1261
rect 2279 1257 2283 1261
rect 2447 1257 2451 1261
rect 2615 1257 2619 1261
rect 2783 1257 2787 1261
rect 2951 1257 2955 1261
rect 3127 1257 3131 1261
rect 3311 1257 3315 1261
rect 3479 1257 3483 1261
rect 2507 1251 2511 1255
rect 3347 1251 3351 1255
rect 3499 1251 3503 1255
rect 543 1231 547 1235
rect 631 1231 635 1235
rect 719 1231 723 1235
rect 807 1231 811 1235
rect 895 1231 899 1235
rect 991 1231 995 1235
rect 1095 1231 1099 1235
rect 1207 1231 1211 1235
rect 1335 1231 1339 1235
rect 1471 1231 1475 1235
rect 1607 1231 1611 1235
rect 1727 1231 1731 1235
rect 111 1221 115 1225
rect 699 1223 703 1227
rect 875 1223 879 1227
rect 1543 1223 1547 1227
rect 2143 1227 2147 1231
rect 2319 1227 2323 1231
rect 2487 1227 2491 1231
rect 2655 1227 2659 1231
rect 2823 1227 2827 1231
rect 2991 1227 2995 1231
rect 3159 1227 3163 1231
rect 3327 1227 3331 1231
rect 3479 1227 3483 1231
rect 1823 1221 1827 1225
rect 1863 1217 1867 1221
rect 2231 1219 2235 1223
rect 2815 1219 2819 1223
rect 3059 1219 3063 1223
rect 3575 1217 3579 1221
rect 111 1204 115 1208
rect 1815 1207 1819 1211
rect 1823 1204 1827 1208
rect 1863 1200 1867 1204
rect 2211 1203 2215 1207
rect 2799 1203 2803 1207
rect 3151 1203 3155 1207
rect 3227 1203 3231 1207
rect 3575 1200 3579 1204
rect 551 1191 555 1195
rect 639 1191 643 1195
rect 727 1191 731 1195
rect 815 1191 819 1195
rect 903 1191 907 1195
rect 999 1191 1003 1195
rect 1103 1191 1107 1195
rect 1215 1191 1219 1195
rect 1343 1191 1347 1195
rect 1479 1191 1483 1195
rect 1615 1191 1619 1195
rect 1735 1191 1739 1195
rect 827 1185 831 1187
rect 827 1183 828 1185
rect 828 1183 831 1185
rect 2151 1187 2155 1191
rect 2327 1187 2331 1191
rect 2495 1187 2499 1191
rect 2663 1187 2667 1191
rect 2831 1187 2835 1191
rect 2999 1187 3003 1191
rect 3167 1187 3171 1191
rect 3335 1187 3339 1191
rect 3487 1187 3491 1191
rect 699 1171 703 1175
rect 1011 1179 1012 1183
rect 1012 1179 1015 1183
rect 1627 1179 1628 1183
rect 1628 1179 1631 1183
rect 875 1171 879 1175
rect 2211 1175 2215 1179
rect 2355 1175 2359 1179
rect 2507 1175 2508 1179
rect 2508 1175 2511 1179
rect 2683 1175 2687 1179
rect 2799 1175 2803 1179
rect 3059 1175 3063 1179
rect 3227 1175 3231 1179
rect 3347 1175 3348 1179
rect 3348 1175 3351 1179
rect 3499 1175 3500 1179
rect 3500 1175 3503 1179
rect 415 1159 419 1163
rect 771 1159 775 1163
rect 1019 1159 1023 1163
rect 1135 1159 1139 1163
rect 1323 1159 1327 1163
rect 1815 1163 1819 1167
rect 2303 1163 2304 1167
rect 2304 1163 2307 1167
rect 2635 1163 2636 1167
rect 2636 1163 2639 1167
rect 2803 1163 2804 1167
rect 2804 1163 2807 1167
rect 3151 1163 3152 1167
rect 3152 1163 3155 1167
rect 359 1149 363 1153
rect 471 1149 475 1153
rect 591 1149 595 1153
rect 711 1149 715 1153
rect 831 1149 835 1153
rect 951 1149 955 1153
rect 1063 1149 1067 1153
rect 1183 1149 1187 1153
rect 1303 1149 1307 1153
rect 1423 1149 1427 1153
rect 1895 1153 1899 1157
rect 2007 1153 2011 1157
rect 2143 1153 2147 1157
rect 2295 1153 2299 1157
rect 2455 1153 2459 1157
rect 2623 1153 2627 1157
rect 2791 1153 2795 1157
rect 2967 1153 2971 1157
rect 3143 1153 3147 1157
rect 3327 1153 3331 1157
rect 3487 1153 3491 1157
rect 111 1136 115 1140
rect 771 1135 775 1139
rect 779 1131 783 1135
rect 1011 1135 1015 1139
rect 1019 1131 1023 1135
rect 1135 1131 1139 1135
rect 1823 1136 1827 1140
rect 1863 1140 1867 1144
rect 2355 1139 2359 1143
rect 2683 1139 2687 1143
rect 3575 1140 3579 1144
rect 111 1119 115 1123
rect 1823 1119 1827 1123
rect 1863 1123 1867 1127
rect 2075 1123 2079 1127
rect 2583 1123 2587 1127
rect 351 1109 355 1113
rect 463 1109 467 1113
rect 583 1109 587 1113
rect 703 1109 707 1113
rect 823 1109 827 1113
rect 943 1109 947 1113
rect 1055 1109 1059 1113
rect 1175 1109 1179 1113
rect 1295 1109 1299 1113
rect 1415 1109 1419 1113
rect 1887 1113 1891 1117
rect 1999 1113 2003 1117
rect 2135 1113 2139 1117
rect 2287 1113 2291 1117
rect 2447 1113 2451 1117
rect 2615 1113 2619 1117
rect 2783 1113 2787 1117
rect 631 1103 632 1107
rect 632 1103 635 1107
rect 2635 1107 2639 1111
rect 3575 1123 3579 1127
rect 2959 1113 2963 1117
rect 3135 1113 3139 1117
rect 3319 1113 3323 1117
rect 3479 1113 3483 1117
rect 3367 1107 3368 1111
rect 3368 1107 3371 1111
rect 3499 1107 3503 1111
rect 143 1083 147 1087
rect 287 1083 291 1087
rect 447 1083 451 1087
rect 615 1083 619 1087
rect 783 1083 787 1087
rect 943 1083 947 1087
rect 1103 1083 1107 1087
rect 1255 1083 1259 1087
rect 1407 1083 1411 1087
rect 1559 1083 1563 1087
rect 1895 1083 1899 1087
rect 2047 1083 2051 1087
rect 2215 1083 2219 1087
rect 2391 1083 2395 1087
rect 2567 1083 2571 1087
rect 2735 1083 2739 1087
rect 2895 1083 2899 1087
rect 3047 1083 3051 1087
rect 3199 1083 3203 1087
rect 3351 1083 3355 1087
rect 3479 1083 3483 1087
rect 111 1073 115 1077
rect 683 1075 687 1079
rect 1323 1075 1327 1079
rect 1475 1075 1479 1079
rect 1823 1073 1827 1077
rect 1863 1073 1867 1077
rect 2303 1075 2307 1079
rect 2803 1075 2807 1079
rect 3419 1075 3423 1079
rect 3575 1073 3579 1077
rect 111 1056 115 1060
rect 515 1059 519 1063
rect 1243 1059 1247 1063
rect 1823 1056 1827 1060
rect 1863 1056 1867 1060
rect 1983 1059 1987 1063
rect 1991 1059 1995 1063
rect 2283 1059 2287 1063
rect 2507 1059 2511 1063
rect 2803 1059 2807 1063
rect 2963 1059 2967 1063
rect 3115 1059 3119 1063
rect 3267 1059 3271 1063
rect 3575 1056 3579 1060
rect 151 1043 155 1047
rect 295 1043 299 1047
rect 455 1043 459 1047
rect 623 1043 627 1047
rect 791 1043 795 1047
rect 951 1043 955 1047
rect 1111 1043 1115 1047
rect 1263 1043 1267 1047
rect 1415 1043 1419 1047
rect 1567 1043 1571 1047
rect 1903 1043 1907 1047
rect 2055 1043 2059 1047
rect 2223 1043 2227 1047
rect 2399 1043 2403 1047
rect 2575 1043 2579 1047
rect 2743 1043 2747 1047
rect 2903 1043 2907 1047
rect 3055 1043 3059 1047
rect 3207 1043 3211 1047
rect 3359 1043 3363 1047
rect 3487 1043 3491 1047
rect 163 1031 164 1035
rect 164 1031 167 1035
rect 631 1031 632 1035
rect 632 1031 635 1035
rect 959 1031 960 1035
rect 960 1031 963 1035
rect 1243 1031 1247 1035
rect 1435 1031 1439 1035
rect 1991 1031 1995 1035
rect 2075 1031 2079 1035
rect 2283 1031 2287 1035
rect 2419 1031 2423 1035
rect 2583 1031 2584 1035
rect 2584 1031 2587 1035
rect 2963 1031 2967 1035
rect 3115 1031 3119 1035
rect 3267 1031 3271 1035
rect 3367 1031 3368 1035
rect 3368 1031 3371 1035
rect 3523 1031 3527 1035
rect 247 1015 251 1019
rect 515 1015 519 1019
rect 1119 1015 1123 1019
rect 1611 1015 1615 1019
rect 1719 1015 1720 1019
rect 1720 1015 1723 1019
rect 1983 1015 1984 1019
rect 1984 1015 1987 1019
rect 2067 1015 2071 1019
rect 2507 1015 2508 1019
rect 2508 1015 2511 1019
rect 2683 1015 2687 1019
rect 2803 1015 2804 1019
rect 2804 1015 2807 1019
rect 3499 1015 3500 1019
rect 3500 1015 3503 1019
rect 143 1005 147 1009
rect 287 1005 291 1009
rect 471 1005 475 1009
rect 663 1005 667 1009
rect 847 1005 851 1009
rect 1031 1005 1035 1009
rect 1207 1005 1211 1009
rect 1375 1005 1379 1009
rect 1543 1005 1547 1009
rect 1711 1005 1715 1009
rect 1975 1005 1979 1009
rect 2095 1005 2099 1009
rect 2223 1005 2227 1009
rect 2359 1005 2363 1009
rect 2495 1005 2499 1009
rect 2639 1005 2643 1009
rect 2791 1005 2795 1009
rect 2959 1005 2963 1009
rect 3135 1005 3139 1009
rect 3311 1005 3315 1009
rect 3487 1005 3491 1009
rect 111 992 115 996
rect 771 987 775 991
rect 1435 991 1439 995
rect 1823 992 1827 996
rect 1459 987 1463 991
rect 1863 992 1867 996
rect 2067 991 2071 995
rect 1611 987 1615 991
rect 2419 991 2423 995
rect 3575 992 3579 996
rect 111 975 115 979
rect 1823 975 1827 979
rect 1863 975 1867 979
rect 3283 975 3287 979
rect 3487 975 3491 979
rect 3575 975 3579 979
rect 135 965 139 969
rect 279 965 283 969
rect 463 965 467 969
rect 655 965 659 969
rect 839 965 843 969
rect 1023 965 1027 969
rect 1199 965 1203 969
rect 1367 965 1371 969
rect 1535 965 1539 969
rect 1703 965 1707 969
rect 1967 965 1971 969
rect 2087 965 2091 969
rect 2215 965 2219 969
rect 2351 965 2355 969
rect 2487 965 2491 969
rect 2631 965 2635 969
rect 2783 965 2787 969
rect 2951 965 2955 969
rect 3127 965 3131 969
rect 3303 965 3307 969
rect 3479 965 3483 969
rect 2523 959 2527 963
rect 135 939 139 943
rect 287 939 291 943
rect 471 939 475 943
rect 663 939 667 943
rect 855 939 859 943
rect 1047 939 1051 943
rect 1223 939 1227 943
rect 1399 939 1403 943
rect 1575 939 1579 943
rect 1727 939 1731 943
rect 2143 939 2147 943
rect 2231 939 2235 943
rect 2319 939 2323 943
rect 2407 939 2411 943
rect 2503 939 2507 943
rect 2615 939 2619 943
rect 2751 939 2755 943
rect 2903 939 2907 943
rect 3079 939 3083 943
rect 3263 939 3267 943
rect 3455 939 3459 943
rect 111 929 115 933
rect 799 931 803 935
rect 1719 931 1723 935
rect 1823 929 1827 933
rect 1863 929 1867 933
rect 2683 931 2687 935
rect 3523 931 3527 935
rect 3575 929 3579 933
rect 111 912 115 916
rect 203 915 207 919
rect 1823 912 1827 916
rect 1863 912 1867 916
rect 2211 915 2215 919
rect 2299 915 2303 919
rect 2387 915 2391 919
rect 2475 915 2479 919
rect 2683 915 2687 919
rect 2819 915 2823 919
rect 2971 915 2975 919
rect 3147 915 3151 919
rect 3575 912 3579 916
rect 143 899 147 903
rect 295 899 299 903
rect 479 899 483 903
rect 671 899 675 903
rect 863 899 867 903
rect 1055 899 1059 903
rect 1231 899 1235 903
rect 1407 899 1411 903
rect 1583 899 1587 903
rect 1735 899 1739 903
rect 2151 899 2155 903
rect 2239 899 2243 903
rect 2327 899 2331 903
rect 2415 899 2419 903
rect 2511 899 2515 903
rect 2623 899 2627 903
rect 2759 899 2763 903
rect 2911 899 2915 903
rect 3087 899 3091 903
rect 3271 899 3275 903
rect 3463 899 3467 903
rect 203 887 207 891
rect 303 887 304 891
rect 304 887 307 891
rect 1207 887 1211 891
rect 2211 887 2215 891
rect 2299 887 2303 891
rect 2387 887 2391 891
rect 2475 887 2479 891
rect 2523 887 2524 891
rect 2524 887 2527 891
rect 2819 887 2823 891
rect 2971 887 2975 891
rect 3147 887 3151 891
rect 3283 887 3284 891
rect 3284 887 3287 891
rect 3487 887 3491 891
rect 1087 871 1091 875
rect 2683 879 2687 883
rect 3507 871 3511 875
rect 143 861 147 865
rect 287 861 291 865
rect 471 861 475 865
rect 655 861 659 865
rect 839 861 843 865
rect 1023 861 1027 865
rect 1191 861 1195 865
rect 1359 861 1363 865
rect 1527 861 1531 865
rect 1695 861 1699 865
rect 2103 861 2107 865
rect 2191 861 2195 865
rect 2279 861 2283 865
rect 2367 861 2371 865
rect 2439 863 2443 867
rect 2455 861 2459 865
rect 2567 861 2571 865
rect 2703 861 2707 865
rect 2871 861 2875 865
rect 3055 861 3059 865
rect 3255 861 3259 865
rect 3463 861 3467 865
rect 111 848 115 852
rect 1823 848 1827 852
rect 1863 848 1867 852
rect 1627 843 1631 847
rect 3575 848 3579 852
rect 111 831 115 835
rect 751 831 755 835
rect 1823 831 1827 835
rect 1863 831 1867 835
rect 3139 831 3143 835
rect 3575 831 3579 835
rect 135 821 139 825
rect 279 821 283 825
rect 463 821 467 825
rect 647 821 651 825
rect 831 821 835 825
rect 1015 821 1019 825
rect 1183 821 1187 825
rect 1351 821 1355 825
rect 1519 821 1523 825
rect 1687 821 1691 825
rect 2095 821 2099 825
rect 2183 821 2187 825
rect 2271 821 2275 825
rect 2359 821 2363 825
rect 2447 821 2451 825
rect 2559 821 2563 825
rect 2695 821 2699 825
rect 2863 821 2867 825
rect 3047 821 3051 825
rect 3247 821 3251 825
rect 3455 821 3459 825
rect 2307 815 2311 819
rect 3499 815 3503 819
rect 135 799 139 803
rect 271 799 275 803
rect 423 799 427 803
rect 583 799 587 803
rect 743 799 747 803
rect 895 799 899 803
rect 1039 799 1043 803
rect 1183 799 1187 803
rect 1327 799 1331 803
rect 1479 799 1483 803
rect 2199 799 2203 803
rect 2287 799 2291 803
rect 2375 799 2379 803
rect 2463 799 2467 803
rect 2551 799 2555 803
rect 2655 799 2659 803
rect 2783 799 2787 803
rect 2935 799 2939 803
rect 3111 799 3115 803
rect 3295 799 3299 803
rect 3479 799 3483 803
rect 111 789 115 793
rect 679 791 683 795
rect 1399 791 1403 795
rect 1823 789 1827 793
rect 1863 789 1867 793
rect 2355 791 2359 795
rect 2443 791 2447 795
rect 3199 791 3203 795
rect 3575 789 3579 793
rect 111 772 115 776
rect 1823 772 1827 776
rect 1863 772 1867 776
rect 2267 775 2271 779
rect 2531 775 2535 779
rect 3471 775 3475 779
rect 3575 772 3579 776
rect 143 759 147 763
rect 279 759 283 763
rect 431 759 435 763
rect 591 759 595 763
rect 751 759 755 763
rect 903 759 907 763
rect 1047 759 1051 763
rect 1191 759 1195 763
rect 1335 759 1339 763
rect 1487 759 1491 763
rect 2207 759 2211 763
rect 2295 759 2299 763
rect 2383 759 2387 763
rect 2471 759 2475 763
rect 2559 759 2563 763
rect 2663 759 2667 763
rect 2791 759 2795 763
rect 2943 759 2947 763
rect 3119 759 3123 763
rect 3303 759 3307 763
rect 3487 759 3491 763
rect 155 747 156 751
rect 156 747 159 751
rect 1023 747 1027 751
rect 2307 747 2308 751
rect 2308 747 2311 751
rect 2531 747 2535 751
rect 2611 747 2615 751
rect 2675 747 2676 751
rect 2676 747 2679 751
rect 3499 747 3500 751
rect 3500 747 3503 751
rect 2355 739 2359 743
rect 371 731 372 735
rect 372 731 375 735
rect 2047 731 2051 735
rect 2115 731 2116 735
rect 2116 731 2119 735
rect 2267 731 2268 735
rect 2268 731 2271 735
rect 2707 731 2708 735
rect 2708 731 2711 735
rect 3191 731 3195 735
rect 3451 731 3452 735
rect 3452 731 3455 735
rect 359 721 363 725
rect 447 721 451 725
rect 543 721 547 725
rect 639 721 643 725
rect 735 721 739 725
rect 831 721 835 725
rect 899 723 903 727
rect 927 721 931 725
rect 1031 721 1035 725
rect 1135 721 1139 725
rect 1239 721 1243 725
rect 1943 721 1947 725
rect 2103 721 2107 725
rect 2255 721 2259 725
rect 2407 721 2411 725
rect 2551 721 2555 725
rect 2695 721 2699 725
rect 2839 721 2843 725
rect 2983 721 2987 725
rect 3135 721 3139 725
rect 3287 721 3291 725
rect 3439 721 3443 725
rect 111 708 115 712
rect 1823 708 1827 712
rect 1863 708 1867 712
rect 2047 703 2051 707
rect 2611 707 2615 711
rect 3507 707 3511 711
rect 3575 708 3579 712
rect 111 691 115 695
rect 351 681 355 685
rect 439 681 443 685
rect 535 681 539 685
rect 631 681 635 685
rect 511 675 515 679
rect 1203 691 1207 695
rect 1823 691 1827 695
rect 1863 691 1867 695
rect 1907 691 1911 695
rect 3079 691 3083 695
rect 3227 691 3231 695
rect 3575 691 3579 695
rect 727 681 731 685
rect 823 681 827 685
rect 919 681 923 685
rect 1023 681 1027 685
rect 1127 681 1131 685
rect 1231 681 1235 685
rect 1935 681 1939 685
rect 2095 681 2099 685
rect 2247 681 2251 685
rect 2399 681 2403 685
rect 2543 681 2547 685
rect 2687 681 2691 685
rect 2831 681 2835 685
rect 2975 681 2979 685
rect 3127 681 3131 685
rect 3279 681 3283 685
rect 3431 681 3435 685
rect 2115 663 2119 667
rect 479 655 483 659
rect 567 655 571 659
rect 655 655 659 659
rect 743 655 747 659
rect 831 655 835 659
rect 919 655 923 659
rect 1007 655 1011 659
rect 1095 655 1099 659
rect 1183 655 1187 659
rect 1271 655 1275 659
rect 1887 655 1891 659
rect 2023 655 2027 659
rect 2199 655 2203 659
rect 111 645 115 649
rect 899 647 903 651
rect 1823 645 1827 649
rect 1863 645 1867 649
rect 2099 647 2103 651
rect 2383 655 2387 659
rect 2567 655 2571 659
rect 2743 655 2747 659
rect 2911 655 2915 659
rect 3063 655 3067 659
rect 3207 655 3211 659
rect 3351 655 3355 659
rect 3479 655 3483 659
rect 3191 647 3195 651
rect 3343 647 3347 651
rect 3575 645 3579 649
rect 111 628 115 632
rect 987 631 991 635
rect 1075 631 1079 635
rect 1251 631 1255 635
rect 1823 628 1827 632
rect 1863 628 1867 632
rect 2451 631 2455 635
rect 2715 631 2719 635
rect 3575 628 3579 632
rect 487 615 491 619
rect 575 615 579 619
rect 663 615 667 619
rect 751 615 755 619
rect 839 615 843 619
rect 927 615 931 619
rect 1015 615 1019 619
rect 1103 615 1107 619
rect 1191 615 1195 619
rect 1279 615 1283 619
rect 1895 615 1899 619
rect 2031 615 2035 619
rect 2207 615 2211 619
rect 2391 615 2395 619
rect 2575 615 2579 619
rect 2751 615 2755 619
rect 2919 615 2923 619
rect 3071 615 3075 619
rect 3215 615 3219 619
rect 3359 615 3363 619
rect 3487 615 3491 619
rect 511 603 515 607
rect 987 603 991 607
rect 1075 603 1079 607
rect 1251 603 1255 607
rect 1907 603 1908 607
rect 1908 603 1911 607
rect 2451 603 2455 607
rect 2763 603 2764 607
rect 2764 603 2767 607
rect 2939 603 2943 607
rect 3227 603 3228 607
rect 3228 603 3231 607
rect 3471 603 3475 607
rect 559 591 563 595
rect 887 591 891 595
rect 1027 591 1031 595
rect 1687 591 1691 595
rect 1695 591 1699 595
rect 1971 591 1975 595
rect 2099 591 2100 595
rect 2100 591 2103 595
rect 2715 591 2716 595
rect 2716 591 2719 595
rect 3267 595 3271 599
rect 3343 591 3347 595
rect 503 581 507 585
rect 599 581 603 585
rect 703 581 707 585
rect 815 581 819 585
rect 935 581 939 585
rect 1063 581 1067 585
rect 1191 581 1195 585
rect 1327 581 1331 585
rect 1471 581 1475 585
rect 1615 581 1619 585
rect 1735 581 1739 585
rect 1895 581 1899 585
rect 2087 581 2091 585
rect 2303 581 2307 585
rect 2511 581 2515 585
rect 2703 581 2707 585
rect 2879 581 2883 585
rect 3039 581 3043 585
rect 3199 581 3203 585
rect 3351 581 3355 585
rect 3487 581 3491 585
rect 111 568 115 572
rect 771 563 775 567
rect 887 563 891 567
rect 1823 568 1827 572
rect 1863 568 1867 572
rect 1687 563 1691 567
rect 1971 563 1975 567
rect 2939 567 2943 571
rect 3575 568 3579 572
rect 3267 563 3271 567
rect 111 551 115 555
rect 815 551 819 555
rect 1539 551 1543 555
rect 1823 551 1827 555
rect 1863 551 1867 555
rect 1871 551 1875 555
rect 3351 551 3355 555
rect 3575 551 3579 555
rect 495 541 499 545
rect 591 541 595 545
rect 695 541 699 545
rect 807 541 811 545
rect 927 541 931 545
rect 1055 541 1059 545
rect 1183 541 1187 545
rect 1319 541 1323 545
rect 1463 541 1467 545
rect 1607 541 1611 545
rect 1727 541 1731 545
rect 1887 541 1891 545
rect 2079 541 2083 545
rect 2295 541 2299 545
rect 2503 541 2507 545
rect 2695 541 2699 545
rect 2871 541 2875 545
rect 3031 541 3035 545
rect 3191 541 3195 545
rect 3343 541 3347 545
rect 3479 541 3483 545
rect 159 519 163 523
rect 303 519 307 523
rect 463 519 467 523
rect 631 519 635 523
rect 799 519 803 523
rect 959 519 963 523
rect 1103 519 1107 523
rect 1239 519 1243 523
rect 1367 519 1371 523
rect 1495 519 1499 523
rect 1623 519 1627 523
rect 1727 519 1731 523
rect 111 509 115 513
rect 1027 511 1031 515
rect 1695 511 1699 515
rect 1823 509 1827 513
rect 2079 511 2083 515
rect 2287 511 2291 515
rect 2487 511 2491 515
rect 2671 511 2675 515
rect 2847 511 2851 515
rect 3015 511 3019 515
rect 3175 511 3179 515
rect 3335 511 3339 515
rect 3479 511 3483 515
rect 1863 501 1867 505
rect 3083 503 3087 507
rect 3451 503 3455 507
rect 3575 501 3579 505
rect 111 492 115 496
rect 151 495 155 499
rect 227 495 231 499
rect 371 495 375 499
rect 531 495 535 499
rect 699 495 703 499
rect 1027 495 1031 499
rect 1455 495 1459 499
rect 1463 495 1467 499
rect 1823 492 1827 496
rect 1863 484 1867 488
rect 2419 487 2423 491
rect 3243 487 3247 491
rect 167 479 171 483
rect 311 479 315 483
rect 471 479 475 483
rect 639 479 643 483
rect 807 479 811 483
rect 967 479 971 483
rect 1111 479 1115 483
rect 1247 479 1251 483
rect 1375 479 1379 483
rect 1503 479 1507 483
rect 1631 479 1635 483
rect 3575 484 3579 488
rect 1735 479 1739 483
rect 227 467 231 471
rect 371 467 375 471
rect 531 467 535 471
rect 699 467 703 471
rect 815 467 816 471
rect 816 467 819 471
rect 1027 467 1031 471
rect 1239 467 1243 471
rect 1539 467 1543 471
rect 1871 467 1875 471
rect 2087 471 2091 475
rect 2295 471 2299 475
rect 2495 471 2499 475
rect 2679 471 2683 475
rect 2855 471 2859 475
rect 3023 471 3027 475
rect 3183 471 3187 475
rect 3343 471 3347 475
rect 3487 471 3491 475
rect 1463 459 1467 463
rect 2095 459 2096 463
rect 2096 459 2099 463
rect 2507 459 2508 463
rect 2508 459 2511 463
rect 2687 459 2688 463
rect 2688 459 2691 463
rect 3243 459 3247 463
rect 3351 459 3352 463
rect 3352 459 3355 463
rect 3479 459 3483 463
rect 151 447 152 451
rect 152 447 155 451
rect 383 447 387 451
rect 1455 447 1456 451
rect 1456 447 1459 451
rect 2303 443 2307 447
rect 2579 447 2583 451
rect 2791 447 2795 451
rect 143 437 147 441
rect 271 437 275 441
rect 439 437 443 441
rect 615 437 619 441
rect 791 437 795 441
rect 967 437 971 441
rect 1127 437 1131 441
rect 1287 437 1291 441
rect 1447 437 1451 441
rect 1607 437 1611 441
rect 2247 437 2251 441
rect 2335 437 2339 441
rect 2431 437 2435 441
rect 2527 437 2531 441
rect 2623 437 2627 441
rect 2735 437 2739 441
rect 2863 437 2867 441
rect 3007 437 3011 441
rect 3167 437 3171 441
rect 3335 437 3339 441
rect 3487 437 3491 441
rect 111 424 115 428
rect 383 423 387 427
rect 1823 424 1827 428
rect 1863 424 1867 428
rect 1547 419 1551 423
rect 2507 419 2511 423
rect 2595 419 2599 423
rect 3575 424 3579 428
rect 3479 419 3483 423
rect 111 407 115 411
rect 683 407 687 411
rect 1287 407 1291 411
rect 1823 407 1827 411
rect 1863 407 1867 411
rect 2935 407 2939 411
rect 135 397 139 401
rect 263 397 267 401
rect 431 397 435 401
rect 607 397 611 401
rect 783 397 787 401
rect 959 397 963 401
rect 1119 397 1123 401
rect 1279 397 1283 401
rect 1439 397 1443 401
rect 1599 397 1603 401
rect 2239 397 2243 401
rect 2327 397 2331 401
rect 2423 397 2427 401
rect 2519 397 2523 401
rect 2615 397 2619 401
rect 2727 397 2731 401
rect 2855 397 2859 401
rect 2791 391 2795 395
rect 3575 407 3579 411
rect 2999 397 3003 401
rect 3159 397 3163 401
rect 3327 397 3331 401
rect 3479 397 3483 401
rect 135 375 139 379
rect 263 375 267 379
rect 431 375 435 379
rect 607 375 611 379
rect 783 375 787 379
rect 951 375 955 379
rect 1111 375 1115 379
rect 1271 375 1275 379
rect 1431 375 1435 379
rect 1591 375 1595 379
rect 2151 375 2155 379
rect 2239 375 2243 379
rect 2327 375 2331 379
rect 2415 375 2419 379
rect 2503 375 2507 379
rect 2615 375 2619 379
rect 2751 375 2755 379
rect 2919 375 2923 379
rect 3103 375 3107 379
rect 3303 375 3307 379
rect 3479 375 3483 379
rect 111 365 115 369
rect 691 367 695 371
rect 1823 365 1827 369
rect 1863 365 1867 369
rect 2579 367 2583 371
rect 3199 367 3203 371
rect 3575 365 3579 369
rect 111 348 115 352
rect 1019 351 1023 355
rect 1695 351 1699 355
rect 1823 348 1827 352
rect 1863 348 1867 352
rect 2571 351 2575 355
rect 2683 351 2687 355
rect 3575 348 3579 352
rect 143 335 147 339
rect 271 335 275 339
rect 439 335 443 339
rect 615 335 619 339
rect 791 335 795 339
rect 959 335 963 339
rect 1119 335 1123 339
rect 1279 335 1283 339
rect 1439 335 1443 339
rect 1599 335 1603 339
rect 2159 335 2163 339
rect 2247 335 2251 339
rect 2335 335 2339 339
rect 2423 335 2427 339
rect 2511 335 2515 339
rect 2623 335 2627 339
rect 2759 335 2763 339
rect 2927 335 2931 339
rect 3111 335 3115 339
rect 3311 335 3315 339
rect 3487 335 3491 339
rect 155 323 156 327
rect 156 323 159 327
rect 1019 323 1023 327
rect 1243 323 1247 327
rect 1287 323 1288 327
rect 1288 323 1291 327
rect 2215 323 2219 327
rect 2683 323 2687 327
rect 2771 323 2772 327
rect 2772 323 2775 327
rect 2935 323 2936 327
rect 2936 323 2939 327
rect 351 311 355 315
rect 359 307 363 311
rect 1235 307 1239 311
rect 1695 307 1696 311
rect 1696 307 1699 311
rect 2031 311 2032 315
rect 2032 311 2035 315
rect 2391 311 2395 315
rect 2571 311 2575 315
rect 263 297 267 301
rect 391 297 395 301
rect 527 297 531 301
rect 679 297 683 301
rect 839 297 843 301
rect 1007 297 1011 301
rect 1175 297 1179 301
rect 1343 297 1347 301
rect 1511 297 1515 301
rect 1687 297 1691 301
rect 2023 301 2027 305
rect 2119 301 2123 305
rect 2223 301 2227 305
rect 2327 301 2331 305
rect 2431 301 2435 305
rect 2535 301 2539 305
rect 2639 301 2643 305
rect 2743 301 2747 305
rect 2855 301 2859 305
rect 2967 301 2971 305
rect 111 284 115 288
rect 359 283 363 287
rect 1235 283 1239 287
rect 1823 284 1827 288
rect 1863 288 1867 292
rect 2391 287 2395 291
rect 1243 279 1247 283
rect 2399 283 2403 287
rect 3575 288 3579 292
rect 111 267 115 271
rect 811 267 815 271
rect 1411 267 1415 271
rect 1823 267 1827 271
rect 1863 271 1867 275
rect 2923 271 2927 275
rect 3575 271 3579 275
rect 255 257 259 261
rect 383 257 387 261
rect 519 257 523 261
rect 671 257 675 261
rect 831 257 835 261
rect 999 257 1003 261
rect 1167 257 1171 261
rect 1335 257 1339 261
rect 1503 257 1507 261
rect 1679 257 1683 261
rect 2015 261 2019 265
rect 2111 261 2115 265
rect 2215 261 2219 265
rect 2319 261 2323 265
rect 2423 261 2427 265
rect 2527 261 2531 265
rect 2631 261 2635 265
rect 2735 261 2739 265
rect 2847 261 2851 265
rect 2959 261 2963 265
rect 1959 239 1963 243
rect 2175 239 2179 243
rect 2383 239 2387 243
rect 2583 239 2587 243
rect 2767 239 2771 243
rect 2951 239 2955 243
rect 3127 239 3131 243
rect 3311 239 3315 243
rect 3479 239 3483 243
rect 399 231 403 235
rect 503 231 507 235
rect 615 231 619 235
rect 735 231 739 235
rect 863 231 867 235
rect 991 231 995 235
rect 1119 231 1123 235
rect 1247 231 1251 235
rect 1375 231 1379 235
rect 1495 231 1499 235
rect 1623 231 1627 235
rect 1727 231 1731 235
rect 1863 229 1867 233
rect 2031 231 2035 235
rect 3199 231 3203 235
rect 3575 229 3579 233
rect 111 221 115 225
rect 803 223 807 227
rect 1727 219 1731 223
rect 1823 221 1827 225
rect 1863 212 1867 216
rect 2095 215 2099 219
rect 2243 215 2247 219
rect 111 204 115 208
rect 1059 207 1063 211
rect 1215 207 1219 211
rect 3575 212 3579 216
rect 1823 204 1827 208
rect 1967 199 1971 203
rect 2183 199 2187 203
rect 2391 199 2395 203
rect 2591 199 2595 203
rect 2775 199 2779 203
rect 2959 199 2963 203
rect 3135 199 3139 203
rect 3319 199 3323 203
rect 3487 199 3491 203
rect 407 191 411 195
rect 511 191 515 195
rect 623 191 627 195
rect 743 191 747 195
rect 871 191 875 195
rect 999 191 1003 195
rect 1127 191 1131 195
rect 1255 191 1259 195
rect 1383 191 1387 195
rect 1503 191 1507 195
rect 1631 191 1635 195
rect 1735 191 1739 195
rect 2095 187 2099 191
rect 2243 187 2247 191
rect 2451 187 2455 191
rect 2603 187 2604 191
rect 2604 187 2607 191
rect 3479 187 3483 191
rect 419 179 420 183
rect 420 179 423 183
rect 1059 179 1063 183
rect 1215 179 1219 183
rect 1411 179 1415 183
rect 803 155 807 159
rect 1163 147 1167 151
rect 1727 147 1731 151
rect 2443 143 2447 147
rect 2619 143 2620 147
rect 2620 143 2623 147
rect 223 137 227 141
rect 311 137 315 141
rect 399 137 403 141
rect 487 137 491 141
rect 575 137 579 141
rect 663 137 667 141
rect 751 137 755 141
rect 839 137 843 141
rect 927 137 931 141
rect 1015 137 1019 141
rect 1103 137 1107 141
rect 1191 137 1195 141
rect 1295 137 1299 141
rect 1399 137 1403 141
rect 1511 137 1515 141
rect 1631 137 1635 141
rect 1735 137 1739 141
rect 1895 133 1899 137
rect 1983 133 1987 137
rect 2071 133 2075 137
rect 2159 133 2163 137
rect 2271 133 2275 137
rect 2383 133 2387 137
rect 2495 133 2499 137
rect 2607 133 2611 137
rect 2719 133 2723 137
rect 2823 133 2827 137
rect 2927 133 2931 137
rect 3023 133 3027 137
rect 3119 133 3123 137
rect 3215 133 3219 137
rect 3311 133 3315 137
rect 3399 133 3403 137
rect 3487 133 3491 137
rect 111 124 115 128
rect 1163 123 1167 127
rect 1823 124 1827 128
rect 1863 120 1867 124
rect 2443 119 2447 123
rect 2451 115 2455 119
rect 3575 120 3579 124
rect 3479 115 3483 119
rect 111 107 115 111
rect 1823 107 1827 111
rect 1863 103 1867 107
rect 3575 103 3579 107
rect 215 97 219 101
rect 303 97 307 101
rect 391 97 395 101
rect 479 97 483 101
rect 567 97 571 101
rect 655 97 659 101
rect 743 97 747 101
rect 831 97 835 101
rect 919 97 923 101
rect 1007 97 1011 101
rect 1095 97 1099 101
rect 1183 97 1187 101
rect 1287 97 1291 101
rect 1391 97 1395 101
rect 1503 97 1507 101
rect 1623 97 1627 101
rect 1727 97 1731 101
rect 1887 93 1891 97
rect 1975 93 1979 97
rect 2063 93 2067 97
rect 2151 93 2155 97
rect 2263 93 2267 97
rect 2375 93 2379 97
rect 2487 93 2491 97
rect 2599 93 2603 97
rect 2711 93 2715 97
rect 2815 93 2819 97
rect 2919 93 2923 97
rect 3015 93 3019 97
rect 3111 93 3115 97
rect 3207 93 3211 97
rect 3303 93 3307 97
rect 3391 93 3395 97
rect 3479 93 3483 97
<< m3 >>
rect 111 3650 115 3651
rect 111 3645 115 3646
rect 143 3650 147 3651
rect 143 3645 147 3646
rect 231 3650 235 3651
rect 231 3645 235 3646
rect 319 3650 323 3651
rect 319 3645 323 3646
rect 407 3650 411 3651
rect 407 3645 411 3646
rect 495 3650 499 3651
rect 495 3645 499 3646
rect 583 3650 587 3651
rect 583 3645 587 3646
rect 671 3650 675 3651
rect 671 3645 675 3646
rect 1823 3650 1827 3651
rect 1823 3645 1827 3646
rect 112 3621 114 3645
rect 144 3634 146 3645
rect 232 3634 234 3645
rect 320 3634 322 3645
rect 408 3634 410 3645
rect 496 3634 498 3645
rect 584 3634 586 3645
rect 672 3634 674 3645
rect 142 3633 148 3634
rect 142 3629 143 3633
rect 147 3629 148 3633
rect 142 3628 148 3629
rect 230 3633 236 3634
rect 230 3629 231 3633
rect 235 3629 236 3633
rect 230 3628 236 3629
rect 318 3633 324 3634
rect 318 3629 319 3633
rect 323 3629 324 3633
rect 318 3628 324 3629
rect 406 3633 412 3634
rect 406 3629 407 3633
rect 411 3629 412 3633
rect 406 3628 412 3629
rect 494 3633 500 3634
rect 494 3629 495 3633
rect 499 3629 500 3633
rect 494 3628 500 3629
rect 582 3633 588 3634
rect 582 3629 583 3633
rect 587 3629 588 3633
rect 582 3628 588 3629
rect 670 3633 676 3634
rect 670 3629 671 3633
rect 675 3629 676 3633
rect 670 3628 676 3629
rect 1824 3621 1826 3645
rect 110 3620 116 3621
rect 110 3616 111 3620
rect 115 3616 116 3620
rect 110 3615 116 3616
rect 1822 3620 1828 3621
rect 1822 3616 1823 3620
rect 1827 3616 1828 3620
rect 1822 3615 1828 3616
rect 110 3603 116 3604
rect 110 3599 111 3603
rect 115 3599 116 3603
rect 110 3598 116 3599
rect 650 3603 656 3604
rect 650 3599 651 3603
rect 655 3599 656 3603
rect 650 3598 656 3599
rect 1822 3603 1828 3604
rect 1822 3599 1823 3603
rect 1827 3599 1828 3603
rect 1822 3598 1828 3599
rect 112 3575 114 3598
rect 134 3593 140 3594
rect 134 3589 135 3593
rect 139 3589 140 3593
rect 134 3588 140 3589
rect 222 3593 228 3594
rect 222 3589 223 3593
rect 227 3589 228 3593
rect 222 3588 228 3589
rect 310 3593 316 3594
rect 310 3589 311 3593
rect 315 3589 316 3593
rect 310 3588 316 3589
rect 398 3593 404 3594
rect 398 3589 399 3593
rect 403 3589 404 3593
rect 398 3588 404 3589
rect 486 3593 492 3594
rect 486 3589 487 3593
rect 491 3589 492 3593
rect 486 3588 492 3589
rect 574 3593 580 3594
rect 574 3589 575 3593
rect 579 3589 580 3593
rect 574 3588 580 3589
rect 136 3575 138 3588
rect 224 3575 226 3588
rect 312 3575 314 3588
rect 400 3575 402 3588
rect 488 3575 490 3588
rect 576 3575 578 3588
rect 111 3574 115 3575
rect 111 3569 115 3570
rect 135 3574 139 3575
rect 135 3569 139 3570
rect 223 3574 227 3575
rect 223 3569 227 3570
rect 287 3574 291 3575
rect 287 3569 291 3570
rect 311 3574 315 3575
rect 311 3569 315 3570
rect 399 3574 403 3575
rect 399 3569 403 3570
rect 463 3574 467 3575
rect 463 3569 467 3570
rect 487 3574 491 3575
rect 487 3569 491 3570
rect 575 3574 579 3575
rect 575 3569 579 3570
rect 631 3574 635 3575
rect 631 3569 635 3570
rect 112 3554 114 3569
rect 136 3564 138 3569
rect 288 3564 290 3569
rect 464 3564 466 3569
rect 632 3564 634 3569
rect 134 3563 140 3564
rect 134 3559 135 3563
rect 139 3559 140 3563
rect 134 3558 140 3559
rect 286 3563 292 3564
rect 286 3559 287 3563
rect 291 3559 292 3563
rect 286 3558 292 3559
rect 462 3563 468 3564
rect 462 3559 463 3563
rect 467 3559 468 3563
rect 462 3558 468 3559
rect 630 3563 636 3564
rect 630 3559 631 3563
rect 635 3559 636 3563
rect 630 3558 636 3559
rect 652 3557 654 3598
rect 662 3593 668 3594
rect 662 3589 663 3593
rect 667 3589 668 3593
rect 662 3588 668 3589
rect 664 3575 666 3588
rect 1824 3575 1826 3598
rect 663 3574 667 3575
rect 663 3569 667 3570
rect 791 3574 795 3575
rect 791 3569 795 3570
rect 935 3574 939 3575
rect 935 3569 939 3570
rect 1071 3574 1075 3575
rect 1071 3569 1075 3570
rect 1191 3574 1195 3575
rect 1191 3569 1195 3570
rect 1311 3574 1315 3575
rect 1311 3569 1315 3570
rect 1423 3574 1427 3575
rect 1423 3569 1427 3570
rect 1527 3574 1531 3575
rect 1639 3574 1643 3575
rect 1527 3569 1531 3570
rect 1546 3571 1552 3572
rect 792 3564 794 3569
rect 936 3564 938 3569
rect 1072 3564 1074 3569
rect 1192 3564 1194 3569
rect 1312 3564 1314 3569
rect 1424 3564 1426 3569
rect 1528 3564 1530 3569
rect 1546 3567 1547 3571
rect 1551 3567 1552 3571
rect 1639 3569 1643 3570
rect 1727 3574 1731 3575
rect 1727 3569 1731 3570
rect 1823 3574 1827 3575
rect 1823 3569 1827 3570
rect 1546 3566 1552 3567
rect 790 3563 796 3564
rect 790 3559 791 3563
rect 795 3559 796 3563
rect 790 3558 796 3559
rect 934 3563 940 3564
rect 934 3559 935 3563
rect 939 3559 940 3563
rect 934 3558 940 3559
rect 1070 3563 1076 3564
rect 1070 3559 1071 3563
rect 1075 3559 1076 3563
rect 1070 3558 1076 3559
rect 1190 3563 1196 3564
rect 1190 3559 1191 3563
rect 1195 3559 1196 3563
rect 1190 3558 1196 3559
rect 1310 3563 1316 3564
rect 1310 3559 1311 3563
rect 1315 3559 1316 3563
rect 1310 3558 1316 3559
rect 1422 3563 1428 3564
rect 1422 3559 1423 3563
rect 1427 3559 1428 3563
rect 1422 3558 1428 3559
rect 1526 3563 1532 3564
rect 1526 3559 1527 3563
rect 1531 3559 1532 3563
rect 1526 3558 1532 3559
rect 167 3556 171 3557
rect 651 3556 655 3557
rect 110 3553 116 3554
rect 110 3549 111 3553
rect 115 3549 116 3553
rect 167 3551 171 3552
rect 558 3555 564 3556
rect 558 3551 559 3555
rect 563 3551 564 3555
rect 651 3551 655 3552
rect 110 3548 116 3549
rect 110 3536 116 3537
rect 110 3532 111 3536
rect 115 3532 116 3536
rect 110 3531 116 3532
rect 112 3507 114 3531
rect 142 3523 148 3524
rect 142 3519 143 3523
rect 147 3519 148 3523
rect 142 3518 148 3519
rect 144 3507 146 3518
rect 159 3516 163 3517
rect 168 3512 170 3551
rect 558 3550 564 3551
rect 294 3523 300 3524
rect 294 3519 295 3523
rect 299 3519 300 3523
rect 294 3518 300 3519
rect 470 3523 476 3524
rect 470 3519 471 3523
rect 475 3519 476 3523
rect 470 3518 476 3519
rect 159 3511 163 3512
rect 166 3511 172 3512
rect 111 3506 115 3507
rect 111 3501 115 3502
rect 143 3506 147 3507
rect 143 3501 147 3502
rect 151 3506 155 3507
rect 151 3501 155 3502
rect 112 3477 114 3501
rect 152 3490 154 3501
rect 160 3500 162 3511
rect 166 3507 167 3511
rect 171 3507 172 3511
rect 296 3507 298 3518
rect 472 3507 474 3518
rect 560 3517 562 3550
rect 638 3523 644 3524
rect 638 3519 639 3523
rect 643 3519 644 3523
rect 638 3518 644 3519
rect 798 3523 804 3524
rect 798 3519 799 3523
rect 803 3519 804 3523
rect 798 3518 804 3519
rect 942 3523 948 3524
rect 942 3519 943 3523
rect 947 3519 948 3523
rect 942 3518 948 3519
rect 1078 3523 1084 3524
rect 1078 3519 1079 3523
rect 1083 3519 1084 3523
rect 1078 3518 1084 3519
rect 1198 3523 1204 3524
rect 1198 3519 1199 3523
rect 1203 3519 1204 3523
rect 1198 3518 1204 3519
rect 1318 3523 1324 3524
rect 1318 3519 1319 3523
rect 1323 3519 1324 3523
rect 1318 3518 1324 3519
rect 1430 3523 1436 3524
rect 1430 3519 1431 3523
rect 1435 3519 1436 3523
rect 1430 3518 1436 3519
rect 1534 3523 1540 3524
rect 1534 3519 1535 3523
rect 1539 3519 1540 3523
rect 1534 3518 1540 3519
rect 559 3516 563 3517
rect 559 3511 563 3512
rect 640 3507 642 3518
rect 800 3507 802 3518
rect 807 3516 811 3517
rect 806 3511 807 3516
rect 811 3511 812 3516
rect 806 3510 812 3511
rect 944 3507 946 3518
rect 1080 3507 1082 3518
rect 1200 3507 1202 3518
rect 1320 3507 1322 3518
rect 1395 3516 1399 3517
rect 1395 3511 1399 3512
rect 166 3506 172 3507
rect 295 3506 299 3507
rect 295 3501 299 3502
rect 327 3506 331 3507
rect 327 3501 331 3502
rect 471 3506 475 3507
rect 471 3501 475 3502
rect 495 3506 499 3507
rect 495 3501 499 3502
rect 639 3506 643 3507
rect 639 3501 643 3502
rect 655 3506 659 3507
rect 655 3501 659 3502
rect 799 3506 803 3507
rect 799 3501 803 3502
rect 807 3506 811 3507
rect 807 3501 811 3502
rect 943 3506 947 3507
rect 943 3501 947 3502
rect 951 3506 955 3507
rect 951 3501 955 3502
rect 1079 3506 1083 3507
rect 1079 3501 1083 3502
rect 1087 3506 1091 3507
rect 1087 3501 1091 3502
rect 1199 3506 1203 3507
rect 1199 3501 1203 3502
rect 1207 3506 1211 3507
rect 1207 3501 1211 3502
rect 1319 3506 1323 3507
rect 1319 3501 1323 3502
rect 158 3499 164 3500
rect 158 3495 159 3499
rect 163 3495 164 3499
rect 158 3494 164 3495
rect 328 3490 330 3501
rect 496 3490 498 3501
rect 656 3490 658 3501
rect 808 3490 810 3501
rect 878 3499 884 3500
rect 878 3495 879 3499
rect 883 3495 884 3499
rect 878 3494 884 3495
rect 150 3489 156 3490
rect 150 3485 151 3489
rect 155 3485 156 3489
rect 150 3484 156 3485
rect 326 3489 332 3490
rect 326 3485 327 3489
rect 331 3485 332 3489
rect 326 3484 332 3485
rect 494 3489 500 3490
rect 494 3485 495 3489
rect 499 3485 500 3489
rect 494 3484 500 3485
rect 654 3489 660 3490
rect 654 3485 655 3489
rect 659 3485 660 3489
rect 654 3484 660 3485
rect 806 3489 812 3490
rect 806 3485 807 3489
rect 811 3485 812 3489
rect 806 3484 812 3485
rect 110 3476 116 3477
rect 110 3472 111 3476
rect 115 3472 116 3476
rect 110 3471 116 3472
rect 880 3461 882 3494
rect 952 3490 954 3501
rect 1088 3490 1090 3501
rect 1146 3499 1152 3500
rect 1146 3495 1147 3499
rect 1151 3495 1152 3499
rect 1146 3494 1152 3495
rect 950 3489 956 3490
rect 950 3485 951 3489
rect 955 3485 956 3489
rect 950 3484 956 3485
rect 1086 3489 1092 3490
rect 1086 3485 1087 3489
rect 1091 3485 1092 3489
rect 1086 3484 1092 3485
rect 1148 3476 1150 3494
rect 1208 3490 1210 3501
rect 1320 3490 1322 3501
rect 1206 3489 1212 3490
rect 1206 3485 1207 3489
rect 1211 3485 1212 3489
rect 1206 3484 1212 3485
rect 1318 3489 1324 3490
rect 1318 3485 1319 3489
rect 1323 3485 1324 3489
rect 1318 3484 1324 3485
rect 1146 3475 1152 3476
rect 1146 3471 1147 3475
rect 1151 3471 1152 3475
rect 1396 3472 1398 3511
rect 1432 3507 1434 3518
rect 1536 3507 1538 3518
rect 1431 3506 1435 3507
rect 1431 3501 1435 3502
rect 1535 3506 1539 3507
rect 1535 3501 1539 3502
rect 1432 3490 1434 3501
rect 1536 3490 1538 3501
rect 1548 3500 1550 3566
rect 1640 3564 1642 3569
rect 1728 3564 1730 3569
rect 1638 3563 1644 3564
rect 1638 3559 1639 3563
rect 1643 3559 1644 3563
rect 1638 3558 1644 3559
rect 1726 3563 1732 3564
rect 1726 3559 1727 3563
rect 1731 3559 1732 3563
rect 1726 3558 1732 3559
rect 1824 3554 1826 3569
rect 1822 3553 1828 3554
rect 1822 3549 1823 3553
rect 1827 3549 1828 3553
rect 1822 3548 1828 3549
rect 1822 3536 1828 3537
rect 1822 3532 1823 3536
rect 1827 3532 1828 3536
rect 1822 3531 1828 3532
rect 1646 3523 1652 3524
rect 1646 3519 1647 3523
rect 1651 3519 1652 3523
rect 1646 3518 1652 3519
rect 1734 3523 1740 3524
rect 1734 3519 1735 3523
rect 1739 3519 1740 3523
rect 1734 3518 1740 3519
rect 1648 3507 1650 3518
rect 1736 3507 1738 3518
rect 1824 3507 1826 3531
rect 1647 3506 1651 3507
rect 1647 3501 1651 3502
rect 1735 3506 1739 3507
rect 1735 3501 1739 3502
rect 1823 3506 1827 3507
rect 1823 3501 1827 3502
rect 1863 3502 1867 3503
rect 1546 3499 1552 3500
rect 1546 3495 1547 3499
rect 1551 3495 1552 3499
rect 1546 3494 1552 3495
rect 1648 3490 1650 3501
rect 1736 3490 1738 3501
rect 1430 3489 1436 3490
rect 1430 3485 1431 3489
rect 1435 3485 1436 3489
rect 1430 3484 1436 3485
rect 1534 3489 1540 3490
rect 1534 3485 1535 3489
rect 1539 3485 1540 3489
rect 1534 3484 1540 3485
rect 1646 3489 1652 3490
rect 1646 3485 1647 3489
rect 1651 3485 1652 3489
rect 1646 3484 1652 3485
rect 1734 3489 1740 3490
rect 1734 3485 1735 3489
rect 1739 3485 1740 3489
rect 1734 3484 1740 3485
rect 1824 3477 1826 3501
rect 1863 3497 1867 3498
rect 1895 3502 1899 3503
rect 1895 3497 1899 3498
rect 1983 3502 1987 3503
rect 1983 3497 1987 3498
rect 2071 3502 2075 3503
rect 2071 3497 2075 3498
rect 2159 3502 2163 3503
rect 2159 3497 2163 3498
rect 3575 3502 3579 3503
rect 3575 3497 3579 3498
rect 1822 3476 1828 3477
rect 1822 3472 1823 3476
rect 1827 3472 1828 3476
rect 1864 3473 1866 3497
rect 1896 3486 1898 3497
rect 1984 3486 1986 3497
rect 2072 3486 2074 3497
rect 2160 3486 2162 3497
rect 1894 3485 1900 3486
rect 1894 3481 1895 3485
rect 1899 3481 1900 3485
rect 1894 3480 1900 3481
rect 1982 3485 1988 3486
rect 1982 3481 1983 3485
rect 1987 3481 1988 3485
rect 1982 3480 1988 3481
rect 2070 3485 2076 3486
rect 2070 3481 2071 3485
rect 2075 3481 2076 3485
rect 2070 3480 2076 3481
rect 2158 3485 2164 3486
rect 2158 3481 2159 3485
rect 2163 3481 2164 3485
rect 2158 3480 2164 3481
rect 3576 3473 3578 3497
rect 1146 3470 1152 3471
rect 1394 3471 1400 3472
rect 1822 3471 1828 3472
rect 1862 3472 1868 3473
rect 1394 3467 1395 3471
rect 1399 3467 1400 3471
rect 1862 3468 1863 3472
rect 1867 3468 1868 3472
rect 1862 3467 1868 3468
rect 3574 3472 3580 3473
rect 3574 3468 3575 3472
rect 3579 3468 3580 3472
rect 3574 3467 3580 3468
rect 1394 3466 1400 3467
rect 879 3460 883 3461
rect 110 3459 116 3460
rect 110 3455 111 3459
rect 115 3455 116 3459
rect 110 3454 116 3455
rect 562 3459 568 3460
rect 562 3455 563 3459
rect 567 3455 568 3459
rect 879 3455 883 3456
rect 1647 3460 1651 3461
rect 1647 3455 1651 3456
rect 1822 3459 1828 3460
rect 1822 3455 1823 3459
rect 1827 3455 1828 3459
rect 562 3454 568 3455
rect 112 3439 114 3454
rect 142 3449 148 3450
rect 142 3445 143 3449
rect 147 3445 148 3449
rect 142 3444 148 3445
rect 318 3449 324 3450
rect 318 3445 319 3449
rect 323 3445 324 3449
rect 318 3444 324 3445
rect 486 3449 492 3450
rect 486 3445 487 3449
rect 491 3445 492 3449
rect 486 3444 492 3445
rect 144 3439 146 3444
rect 320 3439 322 3444
rect 488 3439 490 3444
rect 111 3438 115 3439
rect 111 3433 115 3434
rect 143 3438 147 3439
rect 143 3433 147 3434
rect 215 3438 219 3439
rect 215 3433 219 3434
rect 319 3438 323 3439
rect 319 3433 323 3434
rect 431 3438 435 3439
rect 431 3433 435 3434
rect 487 3438 491 3439
rect 487 3433 491 3434
rect 112 3418 114 3433
rect 216 3428 218 3433
rect 432 3428 434 3433
rect 214 3427 220 3428
rect 214 3423 215 3427
rect 219 3423 220 3427
rect 214 3422 220 3423
rect 430 3427 436 3428
rect 430 3423 431 3427
rect 435 3423 436 3427
rect 430 3422 436 3423
rect 110 3417 116 3418
rect 110 3413 111 3417
rect 115 3413 116 3417
rect 110 3412 116 3413
rect 110 3400 116 3401
rect 110 3396 111 3400
rect 115 3396 116 3400
rect 110 3395 116 3396
rect 112 3363 114 3395
rect 222 3387 228 3388
rect 222 3383 223 3387
rect 227 3383 228 3387
rect 222 3382 228 3383
rect 438 3387 444 3388
rect 438 3383 439 3387
rect 443 3383 444 3387
rect 438 3382 444 3383
rect 224 3363 226 3382
rect 235 3380 239 3381
rect 234 3375 240 3376
rect 234 3371 235 3375
rect 239 3371 240 3375
rect 234 3370 240 3371
rect 440 3363 442 3382
rect 564 3381 566 3454
rect 646 3449 652 3450
rect 646 3445 647 3449
rect 651 3445 652 3449
rect 646 3444 652 3445
rect 798 3449 804 3450
rect 798 3445 799 3449
rect 803 3445 804 3449
rect 798 3444 804 3445
rect 942 3449 948 3450
rect 942 3445 943 3449
rect 947 3445 948 3449
rect 942 3444 948 3445
rect 1078 3449 1084 3450
rect 1078 3445 1079 3449
rect 1083 3445 1084 3449
rect 1078 3444 1084 3445
rect 1198 3449 1204 3450
rect 1198 3445 1199 3449
rect 1203 3445 1204 3449
rect 1198 3444 1204 3445
rect 1310 3449 1316 3450
rect 1310 3445 1311 3449
rect 1315 3445 1316 3449
rect 1310 3444 1316 3445
rect 1422 3449 1428 3450
rect 1422 3445 1423 3449
rect 1427 3445 1428 3449
rect 1422 3444 1428 3445
rect 1526 3449 1532 3450
rect 1526 3445 1527 3449
rect 1531 3445 1532 3449
rect 1526 3444 1532 3445
rect 1638 3449 1644 3450
rect 1638 3445 1639 3449
rect 1643 3445 1644 3449
rect 1638 3444 1644 3445
rect 648 3439 650 3444
rect 800 3439 802 3444
rect 944 3439 946 3444
rect 1080 3439 1082 3444
rect 1200 3439 1202 3444
rect 1312 3439 1314 3444
rect 1424 3439 1426 3444
rect 1528 3439 1530 3444
rect 1640 3439 1642 3444
rect 639 3438 643 3439
rect 639 3433 643 3434
rect 647 3438 651 3439
rect 647 3433 651 3434
rect 799 3438 803 3439
rect 799 3433 803 3434
rect 847 3438 851 3439
rect 847 3433 851 3434
rect 943 3438 947 3439
rect 943 3433 947 3434
rect 1039 3438 1043 3439
rect 1039 3433 1043 3434
rect 1079 3438 1083 3439
rect 1079 3433 1083 3434
rect 1199 3438 1203 3439
rect 1199 3433 1203 3434
rect 1223 3438 1227 3439
rect 1223 3433 1227 3434
rect 1311 3438 1315 3439
rect 1311 3433 1315 3434
rect 1399 3438 1403 3439
rect 1399 3433 1403 3434
rect 1423 3438 1427 3439
rect 1423 3433 1427 3434
rect 1527 3438 1531 3439
rect 1527 3433 1531 3434
rect 1567 3438 1571 3439
rect 1567 3433 1571 3434
rect 1639 3438 1643 3439
rect 1639 3433 1643 3434
rect 640 3428 642 3433
rect 848 3428 850 3433
rect 1040 3428 1042 3433
rect 1224 3428 1226 3433
rect 1400 3428 1402 3433
rect 1568 3428 1570 3433
rect 638 3427 644 3428
rect 638 3423 639 3427
rect 643 3423 644 3427
rect 638 3422 644 3423
rect 846 3427 852 3428
rect 846 3423 847 3427
rect 851 3423 852 3427
rect 846 3422 852 3423
rect 1038 3427 1044 3428
rect 1038 3423 1039 3427
rect 1043 3423 1044 3427
rect 1038 3422 1044 3423
rect 1222 3427 1228 3428
rect 1222 3423 1223 3427
rect 1227 3423 1228 3427
rect 1222 3422 1228 3423
rect 1398 3427 1404 3428
rect 1398 3423 1399 3427
rect 1403 3423 1404 3427
rect 1398 3422 1404 3423
rect 1566 3427 1572 3428
rect 1566 3423 1567 3427
rect 1571 3423 1572 3427
rect 1566 3422 1572 3423
rect 1648 3420 1650 3455
rect 1822 3454 1828 3455
rect 1862 3455 1868 3456
rect 1726 3449 1732 3450
rect 1726 3445 1727 3449
rect 1731 3445 1732 3449
rect 1726 3444 1732 3445
rect 1728 3439 1730 3444
rect 1824 3439 1826 3454
rect 1862 3451 1863 3455
rect 1867 3451 1868 3455
rect 1862 3450 1868 3451
rect 2138 3455 2144 3456
rect 2138 3451 2139 3455
rect 2143 3451 2144 3455
rect 2138 3450 2144 3451
rect 3574 3455 3580 3456
rect 3574 3451 3575 3455
rect 3579 3451 3580 3455
rect 3574 3450 3580 3451
rect 1727 3438 1731 3439
rect 1727 3433 1731 3434
rect 1823 3438 1827 3439
rect 1864 3435 1866 3450
rect 1886 3445 1892 3446
rect 1886 3441 1887 3445
rect 1891 3441 1892 3445
rect 1886 3440 1892 3441
rect 1974 3445 1980 3446
rect 1974 3441 1975 3445
rect 1979 3441 1980 3445
rect 1974 3440 1980 3441
rect 2062 3445 2068 3446
rect 2062 3441 2063 3445
rect 2067 3441 2068 3445
rect 2062 3440 2068 3441
rect 1888 3435 1890 3440
rect 1914 3439 1920 3440
rect 1914 3435 1915 3439
rect 1919 3435 1920 3439
rect 1976 3435 1978 3440
rect 2064 3435 2066 3440
rect 1823 3433 1827 3434
rect 1863 3434 1867 3435
rect 1728 3428 1730 3433
rect 1726 3427 1732 3428
rect 1726 3423 1727 3427
rect 1731 3423 1732 3427
rect 1726 3422 1732 3423
rect 738 3419 744 3420
rect 738 3415 739 3419
rect 743 3415 744 3419
rect 738 3414 744 3415
rect 1646 3419 1652 3420
rect 1646 3415 1647 3419
rect 1651 3415 1652 3419
rect 1824 3418 1826 3433
rect 1863 3429 1867 3430
rect 1887 3434 1891 3435
rect 1914 3434 1920 3435
rect 1975 3434 1979 3435
rect 1887 3429 1891 3430
rect 1646 3414 1652 3415
rect 1822 3417 1828 3418
rect 646 3387 652 3388
rect 646 3383 647 3387
rect 651 3383 652 3387
rect 646 3382 652 3383
rect 563 3380 567 3381
rect 563 3375 567 3376
rect 648 3363 650 3382
rect 740 3364 742 3414
rect 1822 3413 1823 3417
rect 1827 3413 1828 3417
rect 1864 3414 1866 3429
rect 1888 3424 1890 3429
rect 1886 3423 1892 3424
rect 1886 3419 1887 3423
rect 1891 3419 1892 3423
rect 1886 3418 1892 3419
rect 1822 3412 1828 3413
rect 1862 3413 1868 3414
rect 1862 3409 1863 3413
rect 1867 3409 1868 3413
rect 1862 3408 1868 3409
rect 1822 3400 1828 3401
rect 1822 3396 1823 3400
rect 1827 3396 1828 3400
rect 1822 3395 1828 3396
rect 1862 3396 1868 3397
rect 854 3387 860 3388
rect 854 3383 855 3387
rect 859 3383 860 3387
rect 854 3382 860 3383
rect 1046 3387 1052 3388
rect 1046 3383 1047 3387
rect 1051 3383 1052 3387
rect 1046 3382 1052 3383
rect 1230 3387 1236 3388
rect 1230 3383 1231 3387
rect 1235 3383 1236 3387
rect 1230 3382 1236 3383
rect 1406 3387 1412 3388
rect 1406 3383 1407 3387
rect 1411 3383 1412 3387
rect 1406 3382 1412 3383
rect 1574 3387 1580 3388
rect 1574 3383 1575 3387
rect 1579 3383 1580 3387
rect 1574 3382 1580 3383
rect 1734 3387 1740 3388
rect 1734 3383 1735 3387
rect 1739 3383 1740 3387
rect 1734 3382 1740 3383
rect 738 3363 744 3364
rect 856 3363 858 3382
rect 1048 3363 1050 3382
rect 1206 3375 1212 3376
rect 1206 3370 1207 3375
rect 1211 3370 1212 3375
rect 1207 3367 1211 3368
rect 1232 3363 1234 3382
rect 1408 3363 1410 3382
rect 1576 3363 1578 3382
rect 1583 3372 1587 3373
rect 1583 3367 1587 3368
rect 111 3362 115 3363
rect 111 3357 115 3358
rect 223 3362 227 3363
rect 223 3357 227 3358
rect 239 3362 243 3363
rect 239 3357 243 3358
rect 383 3362 387 3363
rect 383 3357 387 3358
rect 439 3362 443 3363
rect 439 3357 443 3358
rect 543 3362 547 3363
rect 543 3357 547 3358
rect 647 3362 651 3363
rect 647 3357 651 3358
rect 711 3362 715 3363
rect 738 3359 739 3363
rect 743 3359 744 3363
rect 738 3358 744 3359
rect 855 3362 859 3363
rect 711 3357 715 3358
rect 855 3357 859 3358
rect 871 3362 875 3363
rect 871 3357 875 3358
rect 1031 3362 1035 3363
rect 1031 3357 1035 3358
rect 1047 3362 1051 3363
rect 1047 3357 1051 3358
rect 1183 3362 1187 3363
rect 1183 3357 1187 3358
rect 1231 3362 1235 3363
rect 1231 3357 1235 3358
rect 1335 3362 1339 3363
rect 1335 3357 1339 3358
rect 1407 3362 1411 3363
rect 1407 3357 1411 3358
rect 1487 3362 1491 3363
rect 1487 3357 1491 3358
rect 1575 3362 1579 3363
rect 1575 3357 1579 3358
rect 112 3333 114 3357
rect 240 3346 242 3357
rect 384 3346 386 3357
rect 544 3346 546 3357
rect 712 3346 714 3357
rect 872 3346 874 3357
rect 1032 3346 1034 3357
rect 1086 3355 1092 3356
rect 1086 3351 1087 3355
rect 1091 3351 1092 3355
rect 1086 3350 1092 3351
rect 238 3345 244 3346
rect 238 3341 239 3345
rect 243 3341 244 3345
rect 238 3340 244 3341
rect 382 3345 388 3346
rect 382 3341 383 3345
rect 387 3341 388 3345
rect 382 3340 388 3341
rect 542 3345 548 3346
rect 542 3341 543 3345
rect 547 3341 548 3345
rect 542 3340 548 3341
rect 710 3345 716 3346
rect 710 3341 711 3345
rect 715 3341 716 3345
rect 710 3340 716 3341
rect 870 3345 876 3346
rect 870 3341 871 3345
rect 875 3341 876 3345
rect 870 3340 876 3341
rect 1030 3345 1036 3346
rect 1030 3341 1031 3345
rect 1035 3341 1036 3345
rect 1030 3340 1036 3341
rect 110 3332 116 3333
rect 110 3328 111 3332
rect 115 3328 116 3332
rect 110 3327 116 3328
rect 110 3315 116 3316
rect 110 3311 111 3315
rect 115 3311 116 3315
rect 110 3310 116 3311
rect 778 3315 784 3316
rect 778 3311 779 3315
rect 783 3311 784 3315
rect 778 3310 784 3311
rect 112 3291 114 3310
rect 230 3305 236 3306
rect 230 3301 231 3305
rect 235 3301 236 3305
rect 230 3300 236 3301
rect 374 3305 380 3306
rect 374 3301 375 3305
rect 379 3301 380 3305
rect 374 3300 380 3301
rect 534 3305 540 3306
rect 534 3301 535 3305
rect 539 3301 540 3305
rect 534 3300 540 3301
rect 702 3305 708 3306
rect 702 3301 703 3305
rect 707 3301 708 3305
rect 702 3300 708 3301
rect 232 3291 234 3300
rect 376 3291 378 3300
rect 536 3291 538 3300
rect 704 3291 706 3300
rect 111 3290 115 3291
rect 111 3285 115 3286
rect 231 3290 235 3291
rect 231 3285 235 3286
rect 239 3290 243 3291
rect 239 3285 243 3286
rect 375 3290 379 3291
rect 375 3285 379 3286
rect 407 3290 411 3291
rect 407 3285 411 3286
rect 535 3290 539 3291
rect 535 3285 539 3286
rect 575 3290 579 3291
rect 575 3285 579 3286
rect 703 3290 707 3291
rect 703 3285 707 3286
rect 743 3290 747 3291
rect 743 3285 747 3286
rect 112 3270 114 3285
rect 240 3280 242 3285
rect 408 3280 410 3285
rect 576 3280 578 3285
rect 744 3280 746 3285
rect 238 3279 244 3280
rect 238 3275 239 3279
rect 243 3275 244 3279
rect 238 3274 244 3275
rect 406 3279 412 3280
rect 406 3275 407 3279
rect 411 3275 412 3279
rect 406 3274 412 3275
rect 574 3279 580 3280
rect 574 3275 575 3279
rect 579 3275 580 3279
rect 574 3274 580 3275
rect 742 3279 748 3280
rect 742 3275 743 3279
rect 747 3275 748 3279
rect 742 3274 748 3275
rect 498 3271 504 3272
rect 110 3269 116 3270
rect 110 3265 111 3269
rect 115 3265 116 3269
rect 498 3267 499 3271
rect 503 3267 504 3271
rect 498 3266 504 3267
rect 110 3264 116 3265
rect 110 3252 116 3253
rect 110 3248 111 3252
rect 115 3248 116 3252
rect 110 3247 116 3248
rect 112 3211 114 3247
rect 246 3239 252 3240
rect 246 3235 247 3239
rect 251 3235 252 3239
rect 414 3239 420 3240
rect 246 3234 252 3235
rect 259 3236 263 3237
rect 248 3211 250 3234
rect 414 3235 415 3239
rect 419 3235 420 3239
rect 500 3237 502 3266
rect 566 3255 572 3256
rect 566 3251 567 3255
rect 571 3251 572 3255
rect 566 3250 572 3251
rect 642 3255 648 3256
rect 642 3251 643 3255
rect 647 3251 648 3255
rect 642 3250 648 3251
rect 414 3234 420 3235
rect 499 3236 503 3237
rect 259 3231 263 3232
rect 260 3228 262 3231
rect 258 3227 264 3228
rect 258 3223 259 3227
rect 263 3223 264 3227
rect 258 3222 264 3223
rect 416 3211 418 3234
rect 499 3231 503 3232
rect 111 3210 115 3211
rect 111 3205 115 3206
rect 175 3210 179 3211
rect 175 3205 179 3206
rect 247 3210 251 3211
rect 247 3205 251 3206
rect 375 3210 379 3211
rect 375 3205 379 3206
rect 415 3210 419 3211
rect 415 3205 419 3206
rect 559 3210 563 3211
rect 559 3205 563 3206
rect 112 3181 114 3205
rect 176 3194 178 3205
rect 258 3203 264 3204
rect 258 3199 259 3203
rect 263 3199 264 3203
rect 258 3198 264 3199
rect 174 3193 180 3194
rect 174 3189 175 3193
rect 179 3189 180 3193
rect 174 3188 180 3189
rect 110 3180 116 3181
rect 110 3176 111 3180
rect 115 3176 116 3180
rect 260 3176 262 3198
rect 376 3194 378 3205
rect 478 3203 484 3204
rect 478 3199 479 3203
rect 483 3199 484 3203
rect 478 3198 484 3199
rect 374 3193 380 3194
rect 374 3189 375 3193
rect 379 3189 380 3193
rect 374 3188 380 3189
rect 480 3176 482 3198
rect 560 3194 562 3205
rect 568 3204 570 3250
rect 582 3239 588 3240
rect 582 3235 583 3239
rect 587 3235 588 3239
rect 582 3234 588 3235
rect 584 3211 586 3234
rect 644 3228 646 3250
rect 750 3239 756 3240
rect 750 3235 751 3239
rect 755 3235 756 3239
rect 750 3234 756 3235
rect 642 3227 648 3228
rect 642 3223 643 3227
rect 647 3223 648 3227
rect 642 3222 648 3223
rect 752 3211 754 3234
rect 780 3228 782 3310
rect 862 3305 868 3306
rect 862 3301 863 3305
rect 867 3301 868 3305
rect 862 3300 868 3301
rect 1022 3305 1028 3306
rect 1022 3301 1023 3305
rect 1027 3301 1028 3305
rect 1022 3300 1028 3301
rect 864 3291 866 3300
rect 1024 3291 1026 3300
rect 863 3290 867 3291
rect 863 3285 867 3286
rect 895 3290 899 3291
rect 895 3285 899 3286
rect 1023 3290 1027 3291
rect 1023 3285 1027 3286
rect 1047 3290 1051 3291
rect 1088 3288 1090 3350
rect 1184 3346 1186 3357
rect 1336 3346 1338 3357
rect 1488 3346 1490 3357
rect 1182 3345 1188 3346
rect 1182 3341 1183 3345
rect 1187 3341 1188 3345
rect 1182 3340 1188 3341
rect 1334 3345 1340 3346
rect 1334 3341 1335 3345
rect 1339 3341 1340 3345
rect 1334 3340 1340 3341
rect 1486 3345 1492 3346
rect 1486 3341 1487 3345
rect 1491 3341 1492 3345
rect 1486 3340 1492 3341
rect 1584 3328 1586 3367
rect 1736 3363 1738 3382
rect 1824 3363 1826 3395
rect 1862 3392 1863 3396
rect 1867 3392 1868 3396
rect 1862 3391 1868 3392
rect 1864 3367 1866 3391
rect 1894 3383 1900 3384
rect 1894 3379 1895 3383
rect 1899 3379 1900 3383
rect 1894 3378 1900 3379
rect 1907 3380 1911 3381
rect 1896 3367 1898 3378
rect 1907 3375 1911 3376
rect 1863 3366 1867 3367
rect 1639 3362 1643 3363
rect 1639 3357 1643 3358
rect 1735 3362 1739 3363
rect 1735 3357 1739 3358
rect 1823 3362 1827 3363
rect 1863 3361 1867 3362
rect 1895 3366 1899 3367
rect 1895 3361 1899 3362
rect 1823 3357 1827 3358
rect 1640 3346 1642 3357
rect 1638 3345 1644 3346
rect 1638 3341 1639 3345
rect 1643 3341 1644 3345
rect 1638 3340 1644 3341
rect 1824 3333 1826 3357
rect 1864 3337 1866 3361
rect 1896 3350 1898 3361
rect 1908 3360 1910 3375
rect 1916 3372 1918 3434
rect 1975 3429 1979 3430
rect 1991 3434 1995 3435
rect 1991 3429 1995 3430
rect 2063 3434 2067 3435
rect 2063 3429 2067 3430
rect 2119 3434 2123 3435
rect 2140 3432 2142 3450
rect 2150 3445 2156 3446
rect 2150 3441 2151 3445
rect 2155 3441 2156 3445
rect 2150 3440 2156 3441
rect 2152 3435 2154 3440
rect 3576 3435 3578 3450
rect 2151 3434 2155 3435
rect 2119 3429 2123 3430
rect 2138 3431 2144 3432
rect 1992 3424 1994 3429
rect 2120 3424 2122 3429
rect 2138 3427 2139 3431
rect 2143 3427 2144 3431
rect 2151 3429 2155 3430
rect 2255 3434 2259 3435
rect 2255 3429 2259 3430
rect 2391 3434 2395 3435
rect 2391 3429 2395 3430
rect 2527 3434 2531 3435
rect 2527 3429 2531 3430
rect 2655 3434 2659 3435
rect 2655 3429 2659 3430
rect 2783 3434 2787 3435
rect 2783 3429 2787 3430
rect 2919 3434 2923 3435
rect 2919 3429 2923 3430
rect 3055 3434 3059 3435
rect 3055 3429 3059 3430
rect 3575 3434 3579 3435
rect 3575 3429 3579 3430
rect 2138 3426 2144 3427
rect 2256 3424 2258 3429
rect 2392 3424 2394 3429
rect 2528 3424 2530 3429
rect 2656 3424 2658 3429
rect 2784 3424 2786 3429
rect 2920 3424 2922 3429
rect 3056 3424 3058 3429
rect 1990 3423 1996 3424
rect 1990 3419 1991 3423
rect 1995 3419 1996 3423
rect 1990 3418 1996 3419
rect 2118 3423 2124 3424
rect 2118 3419 2119 3423
rect 2123 3419 2124 3423
rect 2118 3418 2124 3419
rect 2254 3423 2260 3424
rect 2254 3419 2255 3423
rect 2259 3419 2260 3423
rect 2254 3418 2260 3419
rect 2390 3423 2396 3424
rect 2390 3419 2391 3423
rect 2395 3419 2396 3423
rect 2390 3418 2396 3419
rect 2526 3423 2532 3424
rect 2526 3419 2527 3423
rect 2531 3419 2532 3423
rect 2526 3418 2532 3419
rect 2654 3423 2660 3424
rect 2654 3419 2655 3423
rect 2659 3419 2660 3423
rect 2654 3418 2660 3419
rect 2782 3423 2788 3424
rect 2782 3419 2783 3423
rect 2787 3419 2788 3423
rect 2782 3418 2788 3419
rect 2918 3423 2924 3424
rect 2918 3419 2919 3423
rect 2923 3419 2924 3423
rect 2918 3418 2924 3419
rect 3054 3423 3060 3424
rect 3054 3419 3055 3423
rect 3059 3419 3060 3423
rect 3054 3418 3060 3419
rect 2322 3415 2328 3416
rect 2322 3411 2323 3415
rect 2327 3411 2328 3415
rect 3576 3414 3578 3429
rect 2322 3410 2328 3411
rect 3574 3413 3580 3414
rect 1954 3399 1960 3400
rect 1954 3395 1955 3399
rect 1959 3395 1960 3399
rect 1954 3394 1960 3395
rect 1956 3372 1958 3394
rect 1998 3383 2004 3384
rect 1998 3379 1999 3383
rect 2003 3379 2004 3383
rect 1998 3378 2004 3379
rect 2126 3383 2132 3384
rect 2126 3379 2127 3383
rect 2131 3379 2132 3383
rect 2126 3378 2132 3379
rect 2262 3383 2268 3384
rect 2262 3379 2263 3383
rect 2267 3379 2268 3383
rect 2324 3381 2326 3410
rect 3574 3409 3575 3413
rect 3579 3409 3580 3413
rect 3574 3408 3580 3409
rect 3122 3399 3128 3400
rect 3122 3395 3123 3399
rect 3127 3395 3128 3399
rect 3122 3394 3128 3395
rect 3574 3396 3580 3397
rect 2398 3383 2404 3384
rect 2262 3378 2268 3379
rect 2323 3380 2327 3381
rect 1914 3371 1920 3372
rect 1914 3367 1915 3371
rect 1919 3367 1920 3371
rect 1914 3366 1920 3367
rect 1954 3371 1960 3372
rect 1954 3367 1955 3371
rect 1959 3367 1960 3371
rect 2000 3367 2002 3378
rect 2128 3367 2130 3378
rect 2264 3367 2266 3378
rect 2398 3379 2399 3383
rect 2403 3379 2404 3383
rect 2398 3378 2404 3379
rect 2534 3383 2540 3384
rect 2534 3379 2535 3383
rect 2539 3379 2540 3383
rect 2534 3378 2540 3379
rect 2662 3383 2668 3384
rect 2662 3379 2663 3383
rect 2667 3379 2668 3383
rect 2662 3378 2668 3379
rect 2790 3383 2796 3384
rect 2790 3379 2791 3383
rect 2795 3379 2796 3383
rect 2790 3378 2796 3379
rect 2926 3383 2932 3384
rect 2926 3379 2927 3383
rect 2931 3379 2932 3383
rect 2926 3378 2932 3379
rect 3062 3383 3068 3384
rect 3062 3379 3063 3383
rect 3067 3379 3068 3383
rect 3062 3378 3068 3379
rect 2323 3375 2327 3376
rect 2400 3367 2402 3378
rect 2536 3367 2538 3378
rect 2546 3371 2552 3372
rect 2546 3367 2547 3371
rect 2551 3367 2552 3371
rect 2664 3367 2666 3378
rect 2792 3367 2794 3378
rect 2928 3367 2930 3378
rect 3064 3367 3066 3378
rect 1954 3366 1960 3367
rect 1999 3366 2003 3367
rect 1999 3361 2003 3362
rect 2127 3366 2131 3367
rect 2127 3361 2131 3362
rect 2135 3366 2139 3367
rect 2135 3361 2139 3362
rect 2263 3366 2267 3367
rect 2263 3361 2267 3362
rect 2279 3366 2283 3367
rect 2279 3361 2283 3362
rect 2399 3366 2403 3367
rect 2399 3361 2403 3362
rect 2423 3366 2427 3367
rect 2423 3361 2427 3362
rect 2535 3366 2539 3367
rect 2546 3366 2552 3367
rect 2559 3366 2563 3367
rect 2535 3361 2539 3362
rect 1906 3359 1912 3360
rect 1906 3355 1907 3359
rect 1911 3355 1912 3359
rect 1906 3354 1912 3355
rect 2000 3350 2002 3361
rect 2136 3350 2138 3361
rect 2280 3350 2282 3361
rect 2424 3350 2426 3361
rect 1894 3349 1900 3350
rect 1894 3345 1895 3349
rect 1899 3345 1900 3349
rect 1894 3344 1900 3345
rect 1998 3349 2004 3350
rect 1998 3345 1999 3349
rect 2003 3345 2004 3349
rect 1998 3344 2004 3345
rect 2134 3349 2140 3350
rect 2134 3345 2135 3349
rect 2139 3345 2140 3349
rect 2134 3344 2140 3345
rect 2278 3349 2284 3350
rect 2278 3345 2279 3349
rect 2283 3345 2284 3349
rect 2278 3344 2284 3345
rect 2422 3349 2428 3350
rect 2422 3345 2423 3349
rect 2427 3345 2428 3349
rect 2422 3344 2428 3345
rect 1862 3336 1868 3337
rect 1822 3332 1828 3333
rect 1822 3328 1823 3332
rect 1827 3328 1828 3332
rect 1862 3332 1863 3336
rect 1867 3332 1868 3336
rect 2548 3332 2550 3366
rect 2559 3361 2563 3362
rect 2663 3366 2667 3367
rect 2663 3361 2667 3362
rect 2695 3366 2699 3367
rect 2695 3361 2699 3362
rect 2791 3366 2795 3367
rect 2791 3361 2795 3362
rect 2831 3366 2835 3367
rect 2831 3361 2835 3362
rect 2927 3366 2931 3367
rect 2927 3361 2931 3362
rect 2967 3366 2971 3367
rect 2967 3361 2971 3362
rect 3063 3366 3067 3367
rect 3063 3361 3067 3362
rect 3103 3366 3107 3367
rect 3103 3361 3107 3362
rect 2560 3350 2562 3361
rect 2626 3359 2632 3360
rect 2626 3355 2627 3359
rect 2631 3355 2632 3359
rect 2626 3354 2632 3355
rect 2558 3349 2564 3350
rect 2558 3345 2559 3349
rect 2563 3345 2564 3349
rect 2558 3344 2564 3345
rect 2628 3332 2630 3354
rect 2696 3350 2698 3361
rect 2706 3359 2712 3360
rect 2706 3355 2707 3359
rect 2711 3355 2712 3359
rect 2706 3354 2712 3355
rect 2694 3349 2700 3350
rect 2694 3345 2695 3349
rect 2699 3345 2700 3349
rect 2694 3344 2700 3345
rect 1862 3331 1868 3332
rect 2546 3331 2552 3332
rect 1582 3327 1588 3328
rect 1822 3327 1828 3328
rect 2546 3327 2547 3331
rect 2551 3327 2552 3331
rect 1582 3323 1583 3327
rect 1587 3323 1588 3327
rect 2546 3326 2552 3327
rect 2626 3331 2632 3332
rect 2626 3327 2627 3331
rect 2631 3327 2632 3331
rect 2626 3326 2632 3327
rect 1582 3322 1588 3323
rect 1862 3319 1868 3320
rect 1822 3315 1828 3316
rect 1822 3311 1823 3315
rect 1827 3311 1828 3315
rect 1862 3315 1863 3319
rect 1867 3315 1868 3319
rect 1862 3314 1868 3315
rect 2358 3319 2364 3320
rect 2358 3315 2359 3319
rect 2363 3315 2364 3319
rect 2358 3314 2364 3315
rect 1822 3310 1828 3311
rect 1174 3305 1180 3306
rect 1174 3301 1175 3305
rect 1179 3301 1180 3305
rect 1174 3300 1180 3301
rect 1326 3305 1332 3306
rect 1326 3301 1327 3305
rect 1331 3301 1332 3305
rect 1326 3300 1332 3301
rect 1478 3305 1484 3306
rect 1478 3301 1479 3305
rect 1483 3301 1484 3305
rect 1478 3300 1484 3301
rect 1630 3305 1636 3306
rect 1630 3301 1631 3305
rect 1635 3301 1636 3305
rect 1630 3300 1636 3301
rect 1176 3291 1178 3300
rect 1328 3291 1330 3300
rect 1480 3291 1482 3300
rect 1632 3291 1634 3300
rect 1824 3291 1826 3310
rect 1864 3299 1866 3314
rect 1886 3309 1892 3310
rect 1886 3305 1887 3309
rect 1891 3305 1892 3309
rect 1886 3304 1892 3305
rect 1990 3309 1996 3310
rect 1990 3305 1991 3309
rect 1995 3305 1996 3309
rect 1990 3304 1996 3305
rect 2126 3309 2132 3310
rect 2126 3305 2127 3309
rect 2131 3305 2132 3309
rect 2126 3304 2132 3305
rect 2270 3309 2276 3310
rect 2270 3305 2271 3309
rect 2275 3305 2276 3309
rect 2270 3304 2276 3305
rect 1888 3299 1890 3304
rect 1992 3299 1994 3304
rect 2128 3299 2130 3304
rect 2272 3299 2274 3304
rect 1863 3298 1867 3299
rect 1863 3293 1867 3294
rect 1887 3298 1891 3299
rect 1887 3293 1891 3294
rect 1927 3298 1931 3299
rect 1927 3293 1931 3294
rect 1991 3298 1995 3299
rect 1991 3293 1995 3294
rect 2047 3298 2051 3299
rect 2047 3293 2051 3294
rect 2127 3298 2131 3299
rect 2127 3293 2131 3294
rect 2175 3298 2179 3299
rect 2175 3293 2179 3294
rect 2271 3298 2275 3299
rect 2271 3293 2275 3294
rect 2311 3298 2315 3299
rect 2311 3293 2315 3294
rect 1175 3290 1179 3291
rect 1047 3285 1051 3286
rect 1086 3287 1092 3288
rect 896 3280 898 3285
rect 1048 3280 1050 3285
rect 1086 3283 1087 3287
rect 1091 3283 1092 3287
rect 1175 3285 1179 3286
rect 1191 3290 1195 3291
rect 1191 3285 1195 3286
rect 1327 3290 1331 3291
rect 1327 3285 1331 3286
rect 1335 3290 1339 3291
rect 1335 3285 1339 3286
rect 1479 3290 1483 3291
rect 1479 3285 1483 3286
rect 1487 3290 1491 3291
rect 1487 3285 1491 3286
rect 1631 3290 1635 3291
rect 1631 3285 1635 3286
rect 1823 3290 1827 3291
rect 1823 3285 1827 3286
rect 1086 3282 1092 3283
rect 1192 3280 1194 3285
rect 1336 3280 1338 3285
rect 1488 3280 1490 3285
rect 894 3279 900 3280
rect 894 3275 895 3279
rect 899 3275 900 3279
rect 894 3274 900 3275
rect 1046 3279 1052 3280
rect 1046 3275 1047 3279
rect 1051 3275 1052 3279
rect 1046 3274 1052 3275
rect 1190 3279 1196 3280
rect 1190 3275 1191 3279
rect 1195 3275 1196 3279
rect 1190 3274 1196 3275
rect 1334 3279 1340 3280
rect 1334 3275 1335 3279
rect 1339 3275 1340 3279
rect 1334 3274 1340 3275
rect 1486 3279 1492 3280
rect 1486 3275 1487 3279
rect 1491 3275 1492 3279
rect 1486 3274 1492 3275
rect 1824 3270 1826 3285
rect 1864 3278 1866 3293
rect 1928 3288 1930 3293
rect 2048 3288 2050 3293
rect 2176 3288 2178 3293
rect 2312 3288 2314 3293
rect 1926 3287 1932 3288
rect 1926 3283 1927 3287
rect 1931 3283 1932 3287
rect 1926 3282 1932 3283
rect 2046 3287 2052 3288
rect 2046 3283 2047 3287
rect 2051 3283 2052 3287
rect 2046 3282 2052 3283
rect 2174 3287 2180 3288
rect 2174 3283 2175 3287
rect 2179 3283 2180 3287
rect 2174 3282 2180 3283
rect 2310 3287 2316 3288
rect 2310 3283 2311 3287
rect 2315 3283 2316 3287
rect 2310 3282 2316 3283
rect 1862 3277 1868 3278
rect 1862 3273 1863 3277
rect 1867 3273 1868 3277
rect 1862 3272 1868 3273
rect 1822 3269 1828 3270
rect 1822 3265 1823 3269
rect 1827 3265 1828 3269
rect 1822 3264 1828 3265
rect 1862 3260 1868 3261
rect 1862 3256 1863 3260
rect 1867 3256 1868 3260
rect 1862 3255 1868 3256
rect 1822 3252 1828 3253
rect 1822 3248 1823 3252
rect 1827 3248 1828 3252
rect 1822 3247 1828 3248
rect 902 3239 908 3240
rect 902 3235 903 3239
rect 907 3235 908 3239
rect 902 3234 908 3235
rect 1054 3239 1060 3240
rect 1054 3235 1055 3239
rect 1059 3235 1060 3239
rect 1054 3234 1060 3235
rect 1198 3239 1204 3240
rect 1198 3235 1199 3239
rect 1203 3235 1204 3239
rect 1198 3234 1204 3235
rect 1342 3239 1348 3240
rect 1342 3235 1343 3239
rect 1347 3235 1348 3239
rect 1342 3234 1348 3235
rect 1494 3239 1500 3240
rect 1494 3235 1495 3239
rect 1499 3235 1500 3239
rect 1494 3234 1500 3235
rect 778 3227 784 3228
rect 778 3223 779 3227
rect 783 3223 784 3227
rect 778 3222 784 3223
rect 904 3211 906 3234
rect 1030 3227 1036 3228
rect 1030 3223 1031 3227
rect 1035 3223 1036 3227
rect 1030 3222 1036 3223
rect 583 3210 587 3211
rect 583 3205 587 3206
rect 727 3210 731 3211
rect 727 3205 731 3206
rect 751 3210 755 3211
rect 751 3205 755 3206
rect 887 3210 891 3211
rect 887 3205 891 3206
rect 903 3210 907 3211
rect 903 3205 907 3206
rect 566 3203 572 3204
rect 566 3199 567 3203
rect 571 3199 572 3203
rect 566 3198 572 3199
rect 728 3194 730 3205
rect 806 3203 812 3204
rect 806 3199 807 3203
rect 811 3199 812 3203
rect 806 3198 812 3199
rect 558 3193 564 3194
rect 558 3189 559 3193
rect 563 3189 564 3193
rect 558 3188 564 3189
rect 726 3193 732 3194
rect 726 3189 727 3193
rect 731 3189 732 3193
rect 726 3188 732 3189
rect 110 3175 116 3176
rect 258 3175 264 3176
rect 258 3171 259 3175
rect 263 3171 264 3175
rect 258 3170 264 3171
rect 478 3175 484 3176
rect 478 3171 479 3175
rect 483 3171 484 3175
rect 478 3170 484 3171
rect 110 3163 116 3164
rect 110 3159 111 3163
rect 115 3159 116 3163
rect 110 3158 116 3159
rect 154 3163 160 3164
rect 154 3159 155 3163
rect 159 3159 160 3163
rect 154 3158 160 3159
rect 112 3131 114 3158
rect 111 3130 115 3131
rect 111 3125 115 3126
rect 135 3130 139 3131
rect 135 3125 139 3126
rect 112 3110 114 3125
rect 136 3120 138 3125
rect 134 3119 140 3120
rect 134 3115 135 3119
rect 139 3115 140 3119
rect 134 3114 140 3115
rect 110 3109 116 3110
rect 110 3105 111 3109
rect 115 3105 116 3109
rect 110 3104 116 3105
rect 110 3092 116 3093
rect 110 3088 111 3092
rect 115 3088 116 3092
rect 110 3087 116 3088
rect 112 3063 114 3087
rect 142 3079 148 3080
rect 142 3075 143 3079
rect 147 3075 148 3079
rect 142 3074 148 3075
rect 144 3063 146 3074
rect 156 3068 158 3158
rect 166 3153 172 3154
rect 166 3149 167 3153
rect 171 3149 172 3153
rect 166 3148 172 3149
rect 366 3153 372 3154
rect 366 3149 367 3153
rect 371 3149 372 3153
rect 366 3148 372 3149
rect 550 3153 556 3154
rect 550 3149 551 3153
rect 555 3149 556 3153
rect 550 3148 556 3149
rect 718 3153 724 3154
rect 718 3149 719 3153
rect 723 3149 724 3153
rect 808 3149 810 3198
rect 888 3194 890 3205
rect 1032 3197 1034 3222
rect 1056 3211 1058 3234
rect 1200 3211 1202 3234
rect 1344 3211 1346 3234
rect 1496 3211 1498 3234
rect 1824 3211 1826 3247
rect 1864 3223 1866 3255
rect 1934 3247 1940 3248
rect 1934 3243 1935 3247
rect 1939 3243 1940 3247
rect 2054 3247 2060 3248
rect 1934 3242 1940 3243
rect 1947 3244 1951 3245
rect 1936 3223 1938 3242
rect 2054 3243 2055 3247
rect 2059 3243 2060 3247
rect 2054 3242 2060 3243
rect 2182 3247 2188 3248
rect 2182 3243 2183 3247
rect 2187 3243 2188 3247
rect 2182 3242 2188 3243
rect 2318 3247 2324 3248
rect 2318 3243 2319 3247
rect 2323 3243 2324 3247
rect 2360 3245 2362 3314
rect 2414 3309 2420 3310
rect 2414 3305 2415 3309
rect 2419 3305 2420 3309
rect 2414 3304 2420 3305
rect 2550 3309 2556 3310
rect 2550 3305 2551 3309
rect 2555 3305 2556 3309
rect 2550 3304 2556 3305
rect 2686 3309 2692 3310
rect 2686 3305 2687 3309
rect 2691 3305 2692 3309
rect 2686 3304 2692 3305
rect 2416 3299 2418 3304
rect 2552 3299 2554 3304
rect 2688 3299 2690 3304
rect 2415 3298 2419 3299
rect 2415 3293 2419 3294
rect 2455 3298 2459 3299
rect 2455 3293 2459 3294
rect 2551 3298 2555 3299
rect 2551 3293 2555 3294
rect 2599 3298 2603 3299
rect 2599 3293 2603 3294
rect 2687 3298 2691 3299
rect 2687 3293 2691 3294
rect 2456 3288 2458 3293
rect 2600 3288 2602 3293
rect 2454 3287 2460 3288
rect 2454 3283 2455 3287
rect 2459 3283 2460 3287
rect 2454 3282 2460 3283
rect 2598 3287 2604 3288
rect 2598 3283 2599 3287
rect 2603 3283 2604 3287
rect 2598 3282 2604 3283
rect 2708 3280 2710 3354
rect 2832 3350 2834 3361
rect 2898 3359 2904 3360
rect 2898 3355 2899 3359
rect 2903 3355 2904 3359
rect 2898 3354 2904 3355
rect 2830 3349 2836 3350
rect 2830 3345 2831 3349
rect 2835 3345 2836 3349
rect 2830 3344 2836 3345
rect 2900 3332 2902 3354
rect 2968 3350 2970 3361
rect 3034 3359 3040 3360
rect 3034 3355 3035 3359
rect 3039 3355 3040 3359
rect 3034 3354 3040 3355
rect 2966 3349 2972 3350
rect 2966 3345 2967 3349
rect 2971 3345 2972 3349
rect 2966 3344 2972 3345
rect 3036 3332 3038 3354
rect 3104 3350 3106 3361
rect 3124 3360 3126 3394
rect 3574 3392 3575 3396
rect 3579 3392 3580 3396
rect 3574 3391 3580 3392
rect 3576 3367 3578 3391
rect 3575 3366 3579 3367
rect 3575 3361 3579 3362
rect 3122 3359 3128 3360
rect 3122 3355 3123 3359
rect 3127 3355 3128 3359
rect 3122 3354 3128 3355
rect 3102 3349 3108 3350
rect 3102 3345 3103 3349
rect 3107 3345 3108 3349
rect 3102 3344 3108 3345
rect 3576 3337 3578 3361
rect 3574 3336 3580 3337
rect 3574 3332 3575 3336
rect 3579 3332 3580 3336
rect 2898 3331 2904 3332
rect 2898 3327 2899 3331
rect 2903 3327 2904 3331
rect 2898 3326 2904 3327
rect 3034 3331 3040 3332
rect 3574 3331 3580 3332
rect 3034 3327 3035 3331
rect 3039 3327 3040 3331
rect 3034 3326 3040 3327
rect 2902 3319 2908 3320
rect 2902 3315 2903 3319
rect 2907 3315 2908 3319
rect 2902 3314 2908 3315
rect 3574 3319 3580 3320
rect 3574 3315 3575 3319
rect 3579 3315 3580 3319
rect 3574 3314 3580 3315
rect 2822 3309 2828 3310
rect 2822 3305 2823 3309
rect 2827 3305 2828 3309
rect 2822 3304 2828 3305
rect 2824 3299 2826 3304
rect 2743 3298 2747 3299
rect 2743 3293 2747 3294
rect 2823 3298 2827 3299
rect 2823 3293 2827 3294
rect 2887 3298 2891 3299
rect 2887 3293 2891 3294
rect 2744 3288 2746 3293
rect 2888 3288 2890 3293
rect 2742 3287 2748 3288
rect 2742 3283 2743 3287
rect 2747 3283 2748 3287
rect 2742 3282 2748 3283
rect 2886 3287 2892 3288
rect 2886 3283 2887 3287
rect 2891 3283 2892 3287
rect 2886 3282 2892 3283
rect 2382 3279 2388 3280
rect 2382 3275 2383 3279
rect 2387 3275 2388 3279
rect 2382 3274 2388 3275
rect 2706 3279 2712 3280
rect 2706 3275 2707 3279
rect 2711 3275 2712 3279
rect 2706 3274 2712 3275
rect 2318 3242 2324 3243
rect 2359 3244 2363 3245
rect 1947 3239 1951 3240
rect 1948 3236 1950 3239
rect 1946 3235 1952 3236
rect 1946 3231 1947 3235
rect 1951 3231 1952 3235
rect 1946 3230 1952 3231
rect 2056 3223 2058 3242
rect 2184 3223 2186 3242
rect 2320 3223 2322 3242
rect 2359 3239 2363 3240
rect 2384 3224 2386 3274
rect 2462 3247 2468 3248
rect 2462 3243 2463 3247
rect 2467 3243 2468 3247
rect 2462 3242 2468 3243
rect 2606 3247 2612 3248
rect 2606 3243 2607 3247
rect 2611 3243 2612 3247
rect 2606 3242 2612 3243
rect 2750 3247 2756 3248
rect 2750 3243 2751 3247
rect 2755 3243 2756 3247
rect 2750 3242 2756 3243
rect 2894 3247 2900 3248
rect 2894 3243 2895 3247
rect 2899 3243 2900 3247
rect 2894 3242 2900 3243
rect 2382 3223 2388 3224
rect 2464 3223 2466 3242
rect 2608 3223 2610 3242
rect 2618 3235 2624 3236
rect 2618 3231 2619 3235
rect 2623 3231 2624 3235
rect 2618 3230 2624 3231
rect 1863 3222 1867 3223
rect 1863 3217 1867 3218
rect 1935 3222 1939 3223
rect 1935 3217 1939 3218
rect 2007 3222 2011 3223
rect 2007 3217 2011 3218
rect 2055 3222 2059 3223
rect 2055 3217 2059 3218
rect 2119 3222 2123 3223
rect 2119 3217 2123 3218
rect 2183 3222 2187 3223
rect 2183 3217 2187 3218
rect 2239 3222 2243 3223
rect 2239 3217 2243 3218
rect 2319 3222 2323 3223
rect 2319 3217 2323 3218
rect 2375 3222 2379 3223
rect 2382 3219 2383 3223
rect 2387 3219 2388 3223
rect 2382 3218 2388 3219
rect 2463 3222 2467 3223
rect 2375 3217 2379 3218
rect 2463 3217 2467 3218
rect 2519 3222 2523 3223
rect 2519 3217 2523 3218
rect 2607 3222 2611 3223
rect 2607 3217 2611 3218
rect 1039 3210 1043 3211
rect 1039 3205 1043 3206
rect 1055 3210 1059 3211
rect 1055 3205 1059 3206
rect 1191 3210 1195 3211
rect 1191 3205 1195 3206
rect 1199 3210 1203 3211
rect 1199 3205 1203 3206
rect 1343 3210 1347 3211
rect 1343 3205 1347 3206
rect 1351 3210 1355 3211
rect 1351 3205 1355 3206
rect 1495 3210 1499 3211
rect 1495 3205 1499 3206
rect 1823 3210 1827 3211
rect 1823 3205 1827 3206
rect 1031 3196 1035 3197
rect 886 3193 892 3194
rect 886 3189 887 3193
rect 891 3189 892 3193
rect 1040 3194 1042 3205
rect 1192 3194 1194 3205
rect 1279 3196 1283 3197
rect 1031 3191 1035 3192
rect 1038 3193 1044 3194
rect 886 3188 892 3189
rect 1038 3189 1039 3193
rect 1043 3189 1044 3193
rect 1038 3188 1044 3189
rect 1190 3193 1196 3194
rect 1190 3189 1191 3193
rect 1195 3189 1196 3193
rect 1352 3194 1354 3205
rect 1279 3191 1283 3192
rect 1350 3193 1356 3194
rect 1190 3188 1196 3189
rect 1280 3176 1282 3191
rect 1350 3189 1351 3193
rect 1355 3189 1356 3193
rect 1350 3188 1356 3189
rect 1824 3181 1826 3205
rect 1864 3193 1866 3217
rect 2008 3206 2010 3217
rect 2120 3206 2122 3217
rect 2240 3206 2242 3217
rect 2376 3206 2378 3217
rect 2520 3206 2522 3217
rect 2006 3205 2012 3206
rect 2006 3201 2007 3205
rect 2011 3201 2012 3205
rect 2006 3200 2012 3201
rect 2118 3205 2124 3206
rect 2118 3201 2119 3205
rect 2123 3201 2124 3205
rect 2118 3200 2124 3201
rect 2238 3205 2244 3206
rect 2238 3201 2239 3205
rect 2243 3201 2244 3205
rect 2238 3200 2244 3201
rect 2374 3205 2380 3206
rect 2374 3201 2375 3205
rect 2379 3201 2380 3205
rect 2374 3200 2380 3201
rect 2518 3205 2524 3206
rect 2518 3201 2519 3205
rect 2523 3201 2524 3205
rect 2518 3200 2524 3201
rect 1862 3192 1868 3193
rect 1862 3188 1863 3192
rect 1867 3188 1868 3192
rect 2620 3188 2622 3230
rect 2752 3223 2754 3242
rect 2896 3223 2898 3242
rect 2904 3236 2906 3314
rect 2958 3309 2964 3310
rect 2958 3305 2959 3309
rect 2963 3305 2964 3309
rect 2958 3304 2964 3305
rect 3094 3309 3100 3310
rect 3094 3305 3095 3309
rect 3099 3305 3100 3309
rect 3094 3304 3100 3305
rect 2960 3299 2962 3304
rect 3096 3299 3098 3304
rect 3576 3299 3578 3314
rect 2959 3298 2963 3299
rect 2959 3293 2963 3294
rect 3031 3298 3035 3299
rect 3031 3293 3035 3294
rect 3095 3298 3099 3299
rect 3095 3293 3099 3294
rect 3183 3298 3187 3299
rect 3183 3293 3187 3294
rect 3575 3298 3579 3299
rect 3575 3293 3579 3294
rect 3032 3288 3034 3293
rect 3184 3288 3186 3293
rect 3030 3287 3036 3288
rect 3030 3283 3031 3287
rect 3035 3283 3036 3287
rect 3030 3282 3036 3283
rect 3182 3287 3188 3288
rect 3182 3283 3183 3287
rect 3187 3283 3188 3287
rect 3182 3282 3188 3283
rect 3576 3278 3578 3293
rect 3574 3277 3580 3278
rect 3574 3273 3575 3277
rect 3579 3273 3580 3277
rect 3574 3272 3580 3273
rect 3286 3263 3292 3264
rect 3286 3259 3287 3263
rect 3291 3259 3292 3263
rect 3286 3258 3292 3259
rect 3574 3260 3580 3261
rect 3038 3247 3044 3248
rect 3038 3243 3039 3247
rect 3043 3243 3044 3247
rect 3038 3242 3044 3243
rect 3190 3247 3196 3248
rect 3190 3243 3191 3247
rect 3195 3243 3196 3247
rect 3190 3242 3196 3243
rect 2902 3235 2908 3236
rect 2902 3231 2903 3235
rect 2907 3231 2908 3235
rect 2902 3230 2908 3231
rect 3040 3223 3042 3242
rect 3192 3223 3194 3242
rect 2663 3222 2667 3223
rect 2663 3217 2667 3218
rect 2751 3222 2755 3223
rect 2751 3217 2755 3218
rect 2815 3222 2819 3223
rect 2815 3217 2819 3218
rect 2895 3222 2899 3223
rect 2895 3217 2899 3218
rect 2967 3222 2971 3223
rect 2967 3217 2971 3218
rect 3039 3222 3043 3223
rect 3039 3217 3043 3218
rect 3119 3222 3123 3223
rect 3119 3217 3123 3218
rect 3191 3222 3195 3223
rect 3191 3217 3195 3218
rect 3279 3222 3283 3223
rect 3279 3217 3283 3218
rect 2664 3206 2666 3217
rect 2816 3206 2818 3217
rect 2968 3206 2970 3217
rect 3046 3215 3052 3216
rect 3046 3211 3047 3215
rect 3051 3211 3052 3215
rect 3046 3210 3052 3211
rect 2662 3205 2668 3206
rect 2662 3201 2663 3205
rect 2667 3201 2668 3205
rect 2662 3200 2668 3201
rect 2814 3205 2820 3206
rect 2814 3201 2815 3205
rect 2819 3201 2820 3205
rect 2814 3200 2820 3201
rect 2966 3205 2972 3206
rect 2966 3201 2967 3205
rect 2971 3201 2972 3205
rect 2966 3200 2972 3201
rect 3048 3188 3050 3210
rect 3120 3206 3122 3217
rect 3280 3206 3282 3217
rect 3288 3216 3290 3258
rect 3574 3256 3575 3260
rect 3579 3256 3580 3260
rect 3574 3255 3580 3256
rect 3576 3223 3578 3255
rect 3575 3222 3579 3223
rect 3575 3217 3579 3218
rect 3286 3215 3292 3216
rect 3286 3211 3287 3215
rect 3291 3211 3292 3215
rect 3286 3210 3292 3211
rect 3118 3205 3124 3206
rect 3118 3201 3119 3205
rect 3123 3201 3124 3205
rect 3118 3200 3124 3201
rect 3278 3205 3284 3206
rect 3278 3201 3279 3205
rect 3283 3201 3284 3205
rect 3278 3200 3284 3201
rect 3576 3193 3578 3217
rect 3574 3192 3580 3193
rect 3574 3188 3575 3192
rect 3579 3188 3580 3192
rect 1862 3187 1868 3188
rect 2618 3187 2624 3188
rect 2618 3183 2619 3187
rect 2623 3183 2624 3187
rect 2618 3182 2624 3183
rect 3046 3187 3052 3188
rect 3574 3187 3580 3188
rect 3046 3183 3047 3187
rect 3051 3183 3052 3187
rect 3046 3182 3052 3183
rect 1822 3180 1828 3181
rect 1822 3176 1823 3180
rect 1827 3176 1828 3180
rect 1278 3175 1284 3176
rect 1822 3175 1828 3176
rect 1862 3175 1868 3176
rect 1278 3171 1279 3175
rect 1283 3171 1284 3175
rect 1278 3170 1284 3171
rect 1862 3171 1863 3175
rect 1867 3171 1868 3175
rect 1862 3170 1868 3171
rect 3574 3175 3580 3176
rect 3574 3171 3575 3175
rect 3579 3171 3580 3175
rect 3574 3170 3580 3171
rect 1822 3163 1828 3164
rect 1822 3159 1823 3163
rect 1827 3159 1828 3163
rect 1822 3158 1828 3159
rect 878 3153 884 3154
rect 878 3149 879 3153
rect 883 3149 884 3153
rect 718 3148 724 3149
rect 807 3148 811 3149
rect 878 3148 884 3149
rect 1030 3153 1036 3154
rect 1030 3149 1031 3153
rect 1035 3149 1036 3153
rect 1030 3148 1036 3149
rect 1182 3153 1188 3154
rect 1182 3149 1183 3153
rect 1187 3149 1188 3153
rect 1342 3153 1348 3154
rect 1342 3149 1343 3153
rect 1347 3149 1348 3153
rect 1182 3148 1188 3149
rect 1243 3148 1247 3149
rect 1342 3148 1348 3149
rect 168 3131 170 3148
rect 368 3131 370 3148
rect 552 3131 554 3148
rect 720 3131 722 3148
rect 807 3143 811 3144
rect 880 3131 882 3148
rect 1032 3131 1034 3148
rect 1184 3131 1186 3148
rect 1243 3143 1247 3144
rect 167 3130 171 3131
rect 167 3125 171 3126
rect 263 3130 267 3131
rect 263 3125 267 3126
rect 367 3130 371 3131
rect 367 3125 371 3126
rect 399 3130 403 3131
rect 399 3125 403 3126
rect 527 3130 531 3131
rect 527 3125 531 3126
rect 551 3130 555 3131
rect 647 3130 651 3131
rect 551 3125 555 3126
rect 610 3127 616 3128
rect 264 3120 266 3125
rect 400 3120 402 3125
rect 528 3120 530 3125
rect 610 3123 611 3127
rect 615 3123 616 3127
rect 647 3125 651 3126
rect 719 3130 723 3131
rect 719 3125 723 3126
rect 759 3130 763 3131
rect 759 3125 763 3126
rect 863 3130 867 3131
rect 863 3125 867 3126
rect 879 3130 883 3131
rect 879 3125 883 3126
rect 967 3130 971 3131
rect 967 3125 971 3126
rect 1031 3130 1035 3131
rect 1031 3125 1035 3126
rect 1071 3130 1075 3131
rect 1071 3125 1075 3126
rect 1175 3130 1179 3131
rect 1175 3125 1179 3126
rect 1183 3130 1187 3131
rect 1183 3125 1187 3126
rect 610 3122 616 3123
rect 262 3119 268 3120
rect 262 3115 263 3119
rect 267 3115 268 3119
rect 262 3114 268 3115
rect 398 3119 404 3120
rect 398 3115 399 3119
rect 403 3115 404 3119
rect 398 3114 404 3115
rect 526 3119 532 3120
rect 526 3115 527 3119
rect 531 3115 532 3119
rect 526 3114 532 3115
rect 254 3111 260 3112
rect 254 3107 255 3111
rect 259 3107 260 3111
rect 254 3106 260 3107
rect 154 3067 160 3068
rect 154 3063 155 3067
rect 159 3063 160 3067
rect 111 3062 115 3063
rect 111 3057 115 3058
rect 143 3062 147 3063
rect 154 3062 160 3063
rect 247 3062 251 3063
rect 143 3057 147 3058
rect 247 3057 251 3058
rect 112 3033 114 3057
rect 144 3046 146 3057
rect 210 3055 216 3056
rect 210 3051 211 3055
rect 215 3051 216 3055
rect 210 3050 216 3051
rect 142 3045 148 3046
rect 142 3041 143 3045
rect 147 3041 148 3045
rect 142 3040 148 3041
rect 110 3032 116 3033
rect 110 3028 111 3032
rect 115 3028 116 3032
rect 212 3028 214 3050
rect 248 3046 250 3057
rect 256 3056 258 3106
rect 270 3079 276 3080
rect 270 3075 271 3079
rect 275 3075 276 3079
rect 270 3074 276 3075
rect 406 3079 412 3080
rect 406 3075 407 3079
rect 411 3075 412 3079
rect 406 3074 412 3075
rect 534 3079 540 3080
rect 534 3075 535 3079
rect 539 3075 540 3079
rect 534 3074 540 3075
rect 272 3063 274 3074
rect 408 3063 410 3074
rect 426 3067 432 3068
rect 426 3063 427 3067
rect 431 3063 432 3067
rect 536 3063 538 3074
rect 271 3062 275 3063
rect 271 3057 275 3058
rect 367 3062 371 3063
rect 367 3057 371 3058
rect 407 3062 411 3063
rect 426 3062 432 3063
rect 487 3062 491 3063
rect 407 3057 411 3058
rect 254 3055 260 3056
rect 254 3051 255 3055
rect 259 3051 260 3055
rect 254 3050 260 3051
rect 368 3046 370 3057
rect 246 3045 252 3046
rect 246 3041 247 3045
rect 251 3041 252 3045
rect 246 3040 252 3041
rect 366 3045 372 3046
rect 366 3041 367 3045
rect 371 3041 372 3045
rect 366 3040 372 3041
rect 428 3032 430 3062
rect 487 3057 491 3058
rect 535 3062 539 3063
rect 535 3057 539 3058
rect 599 3062 603 3063
rect 599 3057 603 3058
rect 438 3055 444 3056
rect 438 3051 439 3055
rect 443 3051 444 3055
rect 438 3050 444 3051
rect 426 3031 432 3032
rect 110 3027 116 3028
rect 210 3027 216 3028
rect 210 3023 211 3027
rect 215 3023 216 3027
rect 426 3027 427 3031
rect 431 3027 432 3031
rect 440 3028 442 3050
rect 488 3046 490 3057
rect 522 3055 528 3056
rect 522 3051 523 3055
rect 527 3051 528 3055
rect 522 3050 528 3051
rect 486 3045 492 3046
rect 486 3041 487 3045
rect 491 3041 492 3045
rect 486 3040 492 3041
rect 426 3026 432 3027
rect 438 3027 444 3028
rect 210 3022 216 3023
rect 438 3023 439 3027
rect 443 3023 444 3027
rect 438 3022 444 3023
rect 110 3015 116 3016
rect 110 3011 111 3015
rect 115 3011 116 3015
rect 110 3010 116 3011
rect 112 2983 114 3010
rect 134 3005 140 3006
rect 134 3001 135 3005
rect 139 3001 140 3005
rect 134 3000 140 3001
rect 238 3005 244 3006
rect 238 3001 239 3005
rect 243 3001 244 3005
rect 238 3000 244 3001
rect 358 3005 364 3006
rect 358 3001 359 3005
rect 363 3001 364 3005
rect 358 3000 364 3001
rect 478 3005 484 3006
rect 478 3001 479 3005
rect 483 3001 484 3005
rect 478 3000 484 3001
rect 136 2983 138 3000
rect 154 2999 160 3000
rect 154 2995 155 2999
rect 159 2995 160 2999
rect 154 2994 160 2995
rect 111 2982 115 2983
rect 111 2977 115 2978
rect 135 2982 139 2983
rect 135 2977 139 2978
rect 112 2962 114 2977
rect 136 2972 138 2977
rect 134 2971 140 2972
rect 134 2967 135 2971
rect 139 2967 140 2971
rect 134 2966 140 2967
rect 110 2961 116 2962
rect 110 2957 111 2961
rect 115 2957 116 2961
rect 110 2956 116 2957
rect 110 2944 116 2945
rect 110 2940 111 2944
rect 115 2940 116 2944
rect 110 2939 116 2940
rect 112 2915 114 2939
rect 142 2931 148 2932
rect 142 2927 143 2931
rect 147 2927 148 2931
rect 142 2926 148 2927
rect 144 2915 146 2926
rect 156 2920 158 2994
rect 240 2983 242 3000
rect 360 2983 362 3000
rect 480 2983 482 3000
rect 239 2982 243 2983
rect 239 2977 243 2978
rect 287 2982 291 2983
rect 287 2977 291 2978
rect 359 2982 363 2983
rect 359 2977 363 2978
rect 455 2982 459 2983
rect 455 2977 459 2978
rect 479 2982 483 2983
rect 479 2977 483 2978
rect 288 2972 290 2977
rect 456 2972 458 2977
rect 286 2971 292 2972
rect 286 2967 287 2971
rect 291 2967 292 2971
rect 286 2966 292 2967
rect 454 2971 460 2972
rect 454 2967 455 2971
rect 459 2967 460 2971
rect 454 2966 460 2967
rect 524 2964 526 3050
rect 600 3046 602 3057
rect 612 3056 614 3122
rect 648 3120 650 3125
rect 760 3120 762 3125
rect 864 3120 866 3125
rect 968 3120 970 3125
rect 1072 3120 1074 3125
rect 1176 3120 1178 3125
rect 646 3119 652 3120
rect 646 3115 647 3119
rect 651 3115 652 3119
rect 646 3114 652 3115
rect 758 3119 764 3120
rect 758 3115 759 3119
rect 763 3115 764 3119
rect 758 3114 764 3115
rect 862 3119 868 3120
rect 862 3115 863 3119
rect 867 3115 868 3119
rect 862 3114 868 3115
rect 966 3119 972 3120
rect 966 3115 967 3119
rect 971 3115 972 3119
rect 966 3114 972 3115
rect 1070 3119 1076 3120
rect 1070 3115 1071 3119
rect 1075 3115 1076 3119
rect 1070 3114 1076 3115
rect 1174 3119 1180 3120
rect 1174 3115 1175 3119
rect 1179 3115 1180 3119
rect 1174 3114 1180 3115
rect 1244 3112 1246 3143
rect 1344 3131 1346 3148
rect 1824 3131 1826 3158
rect 1864 3151 1866 3170
rect 1998 3165 2004 3166
rect 1998 3161 1999 3165
rect 2003 3161 2004 3165
rect 1998 3160 2004 3161
rect 2110 3165 2116 3166
rect 2110 3161 2111 3165
rect 2115 3161 2116 3165
rect 2110 3160 2116 3161
rect 2230 3165 2236 3166
rect 2230 3161 2231 3165
rect 2235 3161 2236 3165
rect 2230 3160 2236 3161
rect 2366 3165 2372 3166
rect 2366 3161 2367 3165
rect 2371 3161 2372 3165
rect 2366 3160 2372 3161
rect 2510 3165 2516 3166
rect 2510 3161 2511 3165
rect 2515 3161 2516 3165
rect 2510 3160 2516 3161
rect 2654 3165 2660 3166
rect 2654 3161 2655 3165
rect 2659 3161 2660 3165
rect 2654 3160 2660 3161
rect 2806 3165 2812 3166
rect 2806 3161 2807 3165
rect 2811 3161 2812 3165
rect 2806 3160 2812 3161
rect 2958 3165 2964 3166
rect 2958 3161 2959 3165
rect 2963 3161 2964 3165
rect 2958 3160 2964 3161
rect 3110 3165 3116 3166
rect 3110 3161 3111 3165
rect 3115 3161 3116 3165
rect 3110 3160 3116 3161
rect 3270 3165 3276 3166
rect 3270 3161 3271 3165
rect 3275 3161 3276 3165
rect 3270 3160 3276 3161
rect 2000 3151 2002 3160
rect 2112 3151 2114 3160
rect 2232 3151 2234 3160
rect 2368 3151 2370 3160
rect 2512 3151 2514 3160
rect 2530 3159 2536 3160
rect 2530 3155 2531 3159
rect 2535 3155 2536 3159
rect 2530 3154 2536 3155
rect 1863 3150 1867 3151
rect 1863 3145 1867 3146
rect 1999 3150 2003 3151
rect 1999 3145 2003 3146
rect 2055 3150 2059 3151
rect 2055 3145 2059 3146
rect 2111 3150 2115 3151
rect 2111 3145 2115 3146
rect 2207 3150 2211 3151
rect 2207 3145 2211 3146
rect 2231 3150 2235 3151
rect 2231 3145 2235 3146
rect 2359 3150 2363 3151
rect 2359 3145 2363 3146
rect 2367 3150 2371 3151
rect 2367 3145 2371 3146
rect 2511 3150 2515 3151
rect 2511 3145 2515 3146
rect 1279 3130 1283 3131
rect 1279 3125 1283 3126
rect 1343 3130 1347 3131
rect 1343 3125 1347 3126
rect 1823 3130 1827 3131
rect 1864 3130 1866 3145
rect 2056 3140 2058 3145
rect 2208 3140 2210 3145
rect 2360 3140 2362 3145
rect 2512 3140 2514 3145
rect 2054 3139 2060 3140
rect 2054 3135 2055 3139
rect 2059 3135 2060 3139
rect 2054 3134 2060 3135
rect 2206 3139 2212 3140
rect 2206 3135 2207 3139
rect 2211 3135 2212 3139
rect 2206 3134 2212 3135
rect 2358 3139 2364 3140
rect 2358 3135 2359 3139
rect 2363 3135 2364 3139
rect 2358 3134 2364 3135
rect 2510 3139 2516 3140
rect 2510 3135 2511 3139
rect 2515 3135 2516 3139
rect 2510 3134 2516 3135
rect 1823 3125 1827 3126
rect 1862 3129 1868 3130
rect 1862 3125 1863 3129
rect 1867 3125 1868 3129
rect 1280 3120 1282 3125
rect 1278 3119 1284 3120
rect 1278 3115 1279 3119
rect 1283 3115 1284 3119
rect 1278 3114 1284 3115
rect 1242 3111 1248 3112
rect 1242 3107 1243 3111
rect 1247 3107 1248 3111
rect 1824 3110 1826 3125
rect 1862 3124 1868 3125
rect 1962 3115 1968 3116
rect 1862 3112 1868 3113
rect 1242 3106 1248 3107
rect 1822 3109 1828 3110
rect 1822 3105 1823 3109
rect 1827 3105 1828 3109
rect 1862 3108 1863 3112
rect 1867 3108 1868 3112
rect 1962 3111 1963 3115
rect 1967 3111 1968 3115
rect 1962 3110 1968 3111
rect 2122 3115 2128 3116
rect 2122 3111 2123 3115
rect 2127 3111 2128 3115
rect 2122 3110 2128 3111
rect 2274 3115 2280 3116
rect 2274 3111 2275 3115
rect 2279 3111 2280 3115
rect 2274 3110 2280 3111
rect 2426 3115 2432 3116
rect 2426 3111 2427 3115
rect 2431 3111 2432 3115
rect 2426 3110 2432 3111
rect 1862 3107 1868 3108
rect 1822 3104 1828 3105
rect 1822 3092 1828 3093
rect 1822 3088 1823 3092
rect 1827 3088 1828 3092
rect 1822 3087 1828 3088
rect 654 3079 660 3080
rect 654 3075 655 3079
rect 659 3075 660 3079
rect 654 3074 660 3075
rect 766 3079 772 3080
rect 766 3075 767 3079
rect 771 3075 772 3079
rect 766 3074 772 3075
rect 870 3079 876 3080
rect 870 3075 871 3079
rect 875 3075 876 3079
rect 870 3074 876 3075
rect 974 3079 980 3080
rect 974 3075 975 3079
rect 979 3075 980 3079
rect 974 3074 980 3075
rect 1078 3079 1084 3080
rect 1078 3075 1079 3079
rect 1083 3075 1084 3079
rect 1078 3074 1084 3075
rect 1182 3079 1188 3080
rect 1182 3075 1183 3079
rect 1187 3075 1188 3079
rect 1182 3074 1188 3075
rect 1286 3079 1292 3080
rect 1286 3075 1287 3079
rect 1291 3075 1292 3079
rect 1286 3074 1292 3075
rect 656 3063 658 3074
rect 768 3063 770 3074
rect 872 3063 874 3074
rect 950 3067 956 3068
rect 950 3063 951 3067
rect 955 3063 956 3067
rect 976 3063 978 3074
rect 1080 3063 1082 3074
rect 1184 3063 1186 3074
rect 1288 3063 1290 3074
rect 1824 3063 1826 3087
rect 1864 3079 1866 3107
rect 1863 3078 1867 3079
rect 1863 3073 1867 3074
rect 1951 3078 1955 3079
rect 1951 3073 1955 3074
rect 655 3062 659 3063
rect 655 3057 659 3058
rect 703 3062 707 3063
rect 703 3057 707 3058
rect 767 3062 771 3063
rect 767 3057 771 3058
rect 799 3062 803 3063
rect 799 3057 803 3058
rect 871 3062 875 3063
rect 871 3057 875 3058
rect 895 3062 899 3063
rect 950 3062 956 3063
rect 975 3062 979 3063
rect 895 3057 899 3058
rect 610 3055 616 3056
rect 610 3051 611 3055
rect 615 3051 616 3055
rect 610 3050 616 3051
rect 704 3046 706 3057
rect 800 3046 802 3057
rect 896 3046 898 3057
rect 952 3053 954 3062
rect 975 3057 979 3058
rect 991 3062 995 3063
rect 991 3057 995 3058
rect 1079 3062 1083 3063
rect 1079 3057 1083 3058
rect 1087 3062 1091 3063
rect 1087 3057 1091 3058
rect 1183 3062 1187 3063
rect 1183 3057 1187 3058
rect 1287 3062 1291 3063
rect 1287 3057 1291 3058
rect 1823 3062 1827 3063
rect 1823 3057 1827 3058
rect 951 3052 955 3053
rect 951 3047 955 3048
rect 992 3046 994 3057
rect 998 3055 1004 3056
rect 998 3051 999 3055
rect 1003 3051 1004 3055
rect 998 3050 1004 3051
rect 598 3045 604 3046
rect 598 3041 599 3045
rect 603 3041 604 3045
rect 598 3040 604 3041
rect 702 3045 708 3046
rect 702 3041 703 3045
rect 707 3041 708 3045
rect 702 3040 708 3041
rect 798 3045 804 3046
rect 798 3041 799 3045
rect 803 3041 804 3045
rect 798 3040 804 3041
rect 894 3045 900 3046
rect 894 3041 895 3045
rect 899 3041 900 3045
rect 894 3040 900 3041
rect 990 3045 996 3046
rect 990 3041 991 3045
rect 995 3041 996 3045
rect 990 3040 996 3041
rect 590 3005 596 3006
rect 590 3001 591 3005
rect 595 3001 596 3005
rect 590 3000 596 3001
rect 694 3005 700 3006
rect 694 3001 695 3005
rect 699 3001 700 3005
rect 694 3000 700 3001
rect 790 3005 796 3006
rect 790 3001 791 3005
rect 795 3001 796 3005
rect 790 3000 796 3001
rect 886 3005 892 3006
rect 886 3001 887 3005
rect 891 3001 892 3005
rect 886 3000 892 3001
rect 982 3005 988 3006
rect 982 3001 983 3005
rect 987 3001 988 3005
rect 982 3000 988 3001
rect 592 2983 594 3000
rect 696 2983 698 3000
rect 792 2983 794 3000
rect 888 2983 890 3000
rect 946 2999 952 3000
rect 946 2995 947 2999
rect 951 2995 952 2999
rect 946 2994 952 2995
rect 591 2982 595 2983
rect 591 2977 595 2978
rect 623 2982 627 2983
rect 623 2977 627 2978
rect 695 2982 699 2983
rect 695 2977 699 2978
rect 783 2982 787 2983
rect 783 2977 787 2978
rect 791 2982 795 2983
rect 791 2977 795 2978
rect 887 2982 891 2983
rect 887 2977 891 2978
rect 927 2982 931 2983
rect 927 2977 931 2978
rect 624 2972 626 2977
rect 784 2972 786 2977
rect 928 2972 930 2977
rect 622 2971 628 2972
rect 622 2967 623 2971
rect 627 2967 628 2971
rect 622 2966 628 2967
rect 782 2971 788 2972
rect 782 2967 783 2971
rect 787 2967 788 2971
rect 782 2966 788 2967
rect 926 2971 932 2972
rect 926 2967 927 2971
rect 931 2967 932 2971
rect 926 2966 932 2967
rect 522 2963 528 2964
rect 522 2959 523 2963
rect 527 2959 528 2963
rect 522 2958 528 2959
rect 690 2963 696 2964
rect 690 2959 691 2963
rect 695 2959 696 2963
rect 690 2958 696 2959
rect 354 2947 360 2948
rect 354 2943 355 2947
rect 359 2943 360 2947
rect 354 2942 360 2943
rect 294 2931 300 2932
rect 294 2927 295 2931
rect 299 2927 300 2931
rect 294 2926 300 2927
rect 154 2919 160 2920
rect 154 2915 155 2919
rect 159 2915 160 2919
rect 296 2915 298 2926
rect 111 2914 115 2915
rect 111 2909 115 2910
rect 143 2914 147 2915
rect 154 2914 160 2915
rect 295 2914 299 2915
rect 143 2909 147 2910
rect 295 2909 299 2910
rect 319 2914 323 2915
rect 319 2909 323 2910
rect 112 2885 114 2909
rect 144 2898 146 2909
rect 234 2907 240 2908
rect 234 2903 235 2907
rect 239 2903 240 2907
rect 234 2902 240 2903
rect 142 2897 148 2898
rect 142 2893 143 2897
rect 147 2893 148 2897
rect 142 2892 148 2893
rect 110 2884 116 2885
rect 110 2880 111 2884
rect 115 2880 116 2884
rect 236 2880 238 2902
rect 320 2898 322 2909
rect 356 2908 358 2942
rect 462 2931 468 2932
rect 462 2927 463 2931
rect 467 2927 468 2931
rect 462 2926 468 2927
rect 630 2931 636 2932
rect 630 2927 631 2931
rect 635 2927 636 2931
rect 630 2926 636 2927
rect 464 2915 466 2926
rect 475 2924 479 2925
rect 474 2919 480 2920
rect 474 2915 475 2919
rect 479 2915 480 2919
rect 632 2915 634 2926
rect 692 2925 694 2958
rect 790 2931 796 2932
rect 790 2927 791 2931
rect 795 2927 796 2931
rect 790 2926 796 2927
rect 934 2931 940 2932
rect 934 2927 935 2931
rect 939 2927 940 2931
rect 934 2926 940 2927
rect 691 2924 695 2925
rect 691 2919 695 2920
rect 792 2915 794 2926
rect 936 2915 938 2926
rect 948 2920 950 2994
rect 984 2983 986 3000
rect 983 2982 987 2983
rect 983 2977 987 2978
rect 1000 2964 1002 3050
rect 1088 3046 1090 3057
rect 1146 3055 1152 3056
rect 1146 3051 1147 3055
rect 1151 3051 1152 3055
rect 1146 3050 1152 3051
rect 1086 3045 1092 3046
rect 1086 3041 1087 3045
rect 1091 3041 1092 3045
rect 1086 3040 1092 3041
rect 1148 3032 1150 3050
rect 1184 3046 1186 3057
rect 1242 3055 1248 3056
rect 1242 3051 1243 3055
rect 1247 3051 1248 3055
rect 1242 3050 1248 3051
rect 1251 3052 1255 3053
rect 1182 3045 1188 3046
rect 1182 3041 1183 3045
rect 1187 3041 1188 3045
rect 1182 3040 1188 3041
rect 1244 3032 1246 3050
rect 1251 3047 1255 3048
rect 1146 3031 1152 3032
rect 1146 3027 1147 3031
rect 1151 3027 1152 3031
rect 1146 3026 1152 3027
rect 1242 3031 1248 3032
rect 1242 3027 1243 3031
rect 1247 3027 1248 3031
rect 1252 3028 1254 3047
rect 1288 3046 1290 3057
rect 1286 3045 1292 3046
rect 1286 3041 1287 3045
rect 1291 3041 1292 3045
rect 1286 3040 1292 3041
rect 1824 3033 1826 3057
rect 1864 3049 1866 3073
rect 1952 3062 1954 3073
rect 1964 3072 1966 3110
rect 2062 3099 2068 3100
rect 2062 3095 2063 3099
rect 2067 3095 2068 3099
rect 2062 3094 2068 3095
rect 2064 3079 2066 3094
rect 2124 3088 2126 3110
rect 2214 3099 2220 3100
rect 2214 3095 2215 3099
rect 2219 3095 2220 3099
rect 2214 3094 2220 3095
rect 2122 3087 2128 3088
rect 2122 3083 2123 3087
rect 2127 3083 2128 3087
rect 2122 3082 2128 3083
rect 2216 3079 2218 3094
rect 2276 3088 2278 3110
rect 2366 3099 2372 3100
rect 2366 3095 2367 3099
rect 2371 3095 2372 3099
rect 2366 3094 2372 3095
rect 2274 3087 2280 3088
rect 2274 3083 2275 3087
rect 2279 3083 2280 3087
rect 2274 3082 2280 3083
rect 2368 3079 2370 3094
rect 2428 3088 2430 3110
rect 2518 3099 2524 3100
rect 2518 3095 2519 3099
rect 2523 3095 2524 3099
rect 2518 3094 2524 3095
rect 2426 3087 2432 3088
rect 2426 3083 2427 3087
rect 2431 3083 2432 3087
rect 2426 3082 2432 3083
rect 2520 3079 2522 3094
rect 2532 3088 2534 3154
rect 2656 3151 2658 3160
rect 2808 3151 2810 3160
rect 2960 3151 2962 3160
rect 3112 3151 3114 3160
rect 3272 3151 3274 3160
rect 3576 3151 3578 3170
rect 2655 3150 2659 3151
rect 2655 3145 2659 3146
rect 2791 3150 2795 3151
rect 2791 3145 2795 3146
rect 2807 3150 2811 3151
rect 2807 3145 2811 3146
rect 2919 3150 2923 3151
rect 2919 3145 2923 3146
rect 2959 3150 2963 3151
rect 2959 3145 2963 3146
rect 3039 3150 3043 3151
rect 3039 3145 3043 3146
rect 3111 3150 3115 3151
rect 3111 3145 3115 3146
rect 3159 3150 3163 3151
rect 3159 3145 3163 3146
rect 3271 3150 3275 3151
rect 3271 3145 3275 3146
rect 3383 3150 3387 3151
rect 3383 3145 3387 3146
rect 3479 3150 3483 3151
rect 3479 3145 3483 3146
rect 3575 3150 3579 3151
rect 3575 3145 3579 3146
rect 2656 3140 2658 3145
rect 2792 3140 2794 3145
rect 2920 3140 2922 3145
rect 3040 3140 3042 3145
rect 3160 3140 3162 3145
rect 3272 3140 3274 3145
rect 3384 3140 3386 3145
rect 3480 3140 3482 3145
rect 2654 3139 2660 3140
rect 2654 3135 2655 3139
rect 2659 3135 2660 3139
rect 2654 3134 2660 3135
rect 2790 3139 2796 3140
rect 2790 3135 2791 3139
rect 2795 3135 2796 3139
rect 2790 3134 2796 3135
rect 2918 3139 2924 3140
rect 2918 3135 2919 3139
rect 2923 3135 2924 3139
rect 2918 3134 2924 3135
rect 3038 3139 3044 3140
rect 3038 3135 3039 3139
rect 3043 3135 3044 3139
rect 3038 3134 3044 3135
rect 3158 3139 3164 3140
rect 3158 3135 3159 3139
rect 3163 3135 3164 3139
rect 3158 3134 3164 3135
rect 3270 3139 3276 3140
rect 3270 3135 3271 3139
rect 3275 3135 3276 3139
rect 3270 3134 3276 3135
rect 3382 3139 3388 3140
rect 3382 3135 3383 3139
rect 3387 3135 3388 3139
rect 3382 3134 3388 3135
rect 3478 3139 3484 3140
rect 3478 3135 3479 3139
rect 3483 3135 3484 3139
rect 3478 3134 3484 3135
rect 3450 3131 3456 3132
rect 3450 3127 3451 3131
rect 3455 3127 3456 3131
rect 3576 3130 3578 3145
rect 3450 3126 3456 3127
rect 3574 3129 3580 3130
rect 3118 3115 3124 3116
rect 3118 3111 3119 3115
rect 3123 3111 3124 3115
rect 3118 3110 3124 3111
rect 2662 3099 2668 3100
rect 2662 3095 2663 3099
rect 2667 3095 2668 3099
rect 2662 3094 2668 3095
rect 2798 3099 2804 3100
rect 2798 3095 2799 3099
rect 2803 3095 2804 3099
rect 2798 3094 2804 3095
rect 2926 3099 2932 3100
rect 2926 3095 2927 3099
rect 2931 3095 2932 3099
rect 2926 3094 2932 3095
rect 3046 3099 3052 3100
rect 3046 3095 3047 3099
rect 3051 3095 3052 3099
rect 3046 3094 3052 3095
rect 2530 3087 2536 3088
rect 2530 3083 2531 3087
rect 2535 3083 2536 3087
rect 2530 3082 2536 3083
rect 2664 3079 2666 3094
rect 2670 3087 2676 3088
rect 2670 3083 2671 3087
rect 2675 3083 2676 3087
rect 2670 3082 2676 3083
rect 2063 3078 2067 3079
rect 2063 3073 2067 3074
rect 2079 3078 2083 3079
rect 2079 3073 2083 3074
rect 2215 3078 2219 3079
rect 2215 3073 2219 3074
rect 2367 3078 2371 3079
rect 2367 3073 2371 3074
rect 2519 3078 2523 3079
rect 2519 3073 2523 3074
rect 2527 3078 2531 3079
rect 2527 3073 2531 3074
rect 2663 3078 2667 3079
rect 2663 3073 2667 3074
rect 1962 3071 1968 3072
rect 1962 3067 1963 3071
rect 1967 3067 1968 3071
rect 1962 3066 1968 3067
rect 2042 3071 2048 3072
rect 2042 3067 2043 3071
rect 2047 3067 2048 3071
rect 2042 3066 2048 3067
rect 1950 3061 1956 3062
rect 1950 3057 1951 3061
rect 1955 3057 1956 3061
rect 1950 3056 1956 3057
rect 1862 3048 1868 3049
rect 2044 3048 2046 3066
rect 2080 3062 2082 3073
rect 2216 3062 2218 3073
rect 2368 3062 2370 3073
rect 2528 3062 2530 3073
rect 2078 3061 2084 3062
rect 2078 3057 2079 3061
rect 2083 3057 2084 3061
rect 2078 3056 2084 3057
rect 2214 3061 2220 3062
rect 2214 3057 2215 3061
rect 2219 3057 2220 3061
rect 2214 3056 2220 3057
rect 2366 3061 2372 3062
rect 2366 3057 2367 3061
rect 2371 3057 2372 3061
rect 2366 3056 2372 3057
rect 2526 3061 2532 3062
rect 2526 3057 2527 3061
rect 2531 3057 2532 3061
rect 2526 3056 2532 3057
rect 1862 3044 1863 3048
rect 1867 3044 1868 3048
rect 1862 3043 1868 3044
rect 2042 3047 2048 3048
rect 2042 3043 2043 3047
rect 2047 3043 2048 3047
rect 2672 3044 2674 3082
rect 2800 3079 2802 3094
rect 2928 3079 2930 3094
rect 3048 3079 3050 3094
rect 2679 3078 2683 3079
rect 2679 3073 2683 3074
rect 2799 3078 2803 3079
rect 2799 3073 2803 3074
rect 2831 3078 2835 3079
rect 2831 3073 2835 3074
rect 2927 3078 2931 3079
rect 2927 3073 2931 3074
rect 2975 3078 2979 3079
rect 2975 3073 2979 3074
rect 3047 3078 3051 3079
rect 3047 3073 3051 3074
rect 3111 3078 3115 3079
rect 3111 3073 3115 3074
rect 2680 3062 2682 3073
rect 2766 3071 2772 3072
rect 2766 3067 2767 3071
rect 2771 3067 2772 3071
rect 2766 3066 2772 3067
rect 2678 3061 2684 3062
rect 2678 3057 2679 3061
rect 2683 3057 2684 3061
rect 2678 3056 2684 3057
rect 2768 3044 2770 3066
rect 2832 3062 2834 3073
rect 2866 3071 2872 3072
rect 2866 3067 2867 3071
rect 2871 3067 2872 3071
rect 2866 3066 2872 3067
rect 2830 3061 2836 3062
rect 2830 3057 2831 3061
rect 2835 3057 2836 3061
rect 2830 3056 2836 3057
rect 2042 3042 2048 3043
rect 2670 3043 2676 3044
rect 2670 3039 2671 3043
rect 2675 3039 2676 3043
rect 2670 3038 2676 3039
rect 2766 3043 2772 3044
rect 2766 3039 2767 3043
rect 2771 3039 2772 3043
rect 2766 3038 2772 3039
rect 1822 3032 1828 3033
rect 1822 3028 1823 3032
rect 1827 3028 1828 3032
rect 1242 3026 1248 3027
rect 1250 3027 1256 3028
rect 1822 3027 1828 3028
rect 1862 3031 1868 3032
rect 1862 3027 1863 3031
rect 1867 3027 1868 3031
rect 1250 3023 1251 3027
rect 1255 3023 1256 3027
rect 1862 3026 1868 3027
rect 2594 3031 2600 3032
rect 2594 3027 2595 3031
rect 2599 3027 2600 3031
rect 2594 3026 2600 3027
rect 1250 3022 1256 3023
rect 1822 3015 1828 3016
rect 1822 3011 1823 3015
rect 1827 3011 1828 3015
rect 1822 3010 1828 3011
rect 1078 3005 1084 3006
rect 1078 3001 1079 3005
rect 1083 3001 1084 3005
rect 1078 3000 1084 3001
rect 1174 3005 1180 3006
rect 1174 3001 1175 3005
rect 1179 3001 1180 3005
rect 1174 3000 1180 3001
rect 1278 3005 1284 3006
rect 1278 3001 1279 3005
rect 1283 3001 1284 3005
rect 1278 3000 1284 3001
rect 1080 2983 1082 3000
rect 1176 2983 1178 3000
rect 1280 2983 1282 3000
rect 1824 2983 1826 3010
rect 1864 2999 1866 3026
rect 1942 3021 1948 3022
rect 1942 3017 1943 3021
rect 1947 3017 1948 3021
rect 1942 3016 1948 3017
rect 2070 3021 2076 3022
rect 2070 3017 2071 3021
rect 2075 3017 2076 3021
rect 2070 3016 2076 3017
rect 2206 3021 2212 3022
rect 2206 3017 2207 3021
rect 2211 3017 2212 3021
rect 2206 3016 2212 3017
rect 2358 3021 2364 3022
rect 2358 3017 2359 3021
rect 2363 3017 2364 3021
rect 2358 3016 2364 3017
rect 2518 3021 2524 3022
rect 2518 3017 2519 3021
rect 2523 3017 2524 3021
rect 2518 3016 2524 3017
rect 1944 2999 1946 3016
rect 2072 2999 2074 3016
rect 2208 2999 2210 3016
rect 2360 2999 2362 3016
rect 2520 2999 2522 3016
rect 1863 2998 1867 2999
rect 1863 2993 1867 2994
rect 1887 2998 1891 2999
rect 1887 2993 1891 2994
rect 1943 2998 1947 2999
rect 1943 2993 1947 2994
rect 1975 2998 1979 2999
rect 1975 2993 1979 2994
rect 2063 2998 2067 2999
rect 2063 2993 2067 2994
rect 2071 2998 2075 2999
rect 2071 2993 2075 2994
rect 2151 2998 2155 2999
rect 2151 2993 2155 2994
rect 2207 2998 2211 2999
rect 2207 2993 2211 2994
rect 2239 2998 2243 2999
rect 2239 2993 2243 2994
rect 2351 2998 2355 2999
rect 2351 2993 2355 2994
rect 2359 2998 2363 2999
rect 2359 2993 2363 2994
rect 2463 2998 2467 2999
rect 2463 2993 2467 2994
rect 2519 2998 2523 2999
rect 2519 2993 2523 2994
rect 2575 2998 2579 2999
rect 2575 2993 2579 2994
rect 1063 2982 1067 2983
rect 1063 2977 1067 2978
rect 1079 2982 1083 2983
rect 1079 2977 1083 2978
rect 1175 2982 1179 2983
rect 1175 2977 1179 2978
rect 1191 2982 1195 2983
rect 1191 2977 1195 2978
rect 1279 2982 1283 2983
rect 1279 2977 1283 2978
rect 1311 2982 1315 2983
rect 1311 2977 1315 2978
rect 1423 2982 1427 2983
rect 1423 2977 1427 2978
rect 1527 2982 1531 2983
rect 1527 2977 1531 2978
rect 1639 2982 1643 2983
rect 1639 2977 1643 2978
rect 1727 2982 1731 2983
rect 1727 2977 1731 2978
rect 1823 2982 1827 2983
rect 1864 2978 1866 2993
rect 1888 2988 1890 2993
rect 1976 2988 1978 2993
rect 2064 2988 2066 2993
rect 2152 2988 2154 2993
rect 2240 2988 2242 2993
rect 2352 2988 2354 2993
rect 2464 2988 2466 2993
rect 2576 2988 2578 2993
rect 1886 2987 1892 2988
rect 1886 2983 1887 2987
rect 1891 2983 1892 2987
rect 1886 2982 1892 2983
rect 1974 2987 1980 2988
rect 1974 2983 1975 2987
rect 1979 2983 1980 2987
rect 1974 2982 1980 2983
rect 2062 2987 2068 2988
rect 2062 2983 2063 2987
rect 2067 2983 2068 2987
rect 2062 2982 2068 2983
rect 2150 2987 2156 2988
rect 2150 2983 2151 2987
rect 2155 2983 2156 2987
rect 2150 2982 2156 2983
rect 2238 2987 2244 2988
rect 2238 2983 2239 2987
rect 2243 2983 2244 2987
rect 2238 2982 2244 2983
rect 2350 2987 2356 2988
rect 2350 2983 2351 2987
rect 2355 2983 2356 2987
rect 2350 2982 2356 2983
rect 2462 2987 2468 2988
rect 2462 2983 2463 2987
rect 2467 2983 2468 2987
rect 2462 2982 2468 2983
rect 2574 2987 2580 2988
rect 2574 2983 2575 2987
rect 2579 2983 2580 2987
rect 2574 2982 2580 2983
rect 1823 2977 1827 2978
rect 1862 2977 1868 2978
rect 1064 2972 1066 2977
rect 1192 2972 1194 2977
rect 1312 2972 1314 2977
rect 1424 2972 1426 2977
rect 1528 2972 1530 2977
rect 1640 2972 1642 2977
rect 1728 2972 1730 2977
rect 1062 2971 1068 2972
rect 1062 2967 1063 2971
rect 1067 2967 1068 2971
rect 1062 2966 1068 2967
rect 1190 2971 1196 2972
rect 1190 2967 1191 2971
rect 1195 2967 1196 2971
rect 1190 2966 1196 2967
rect 1310 2971 1316 2972
rect 1310 2967 1311 2971
rect 1315 2967 1316 2971
rect 1310 2966 1316 2967
rect 1422 2971 1428 2972
rect 1422 2967 1423 2971
rect 1427 2967 1428 2971
rect 1422 2966 1428 2967
rect 1526 2971 1532 2972
rect 1526 2967 1527 2971
rect 1531 2967 1532 2971
rect 1526 2966 1532 2967
rect 1638 2971 1644 2972
rect 1638 2967 1639 2971
rect 1643 2967 1644 2971
rect 1638 2966 1644 2967
rect 1726 2971 1732 2972
rect 1726 2967 1727 2971
rect 1731 2967 1732 2971
rect 1726 2966 1732 2967
rect 998 2963 1004 2964
rect 998 2959 999 2963
rect 1003 2959 1004 2963
rect 1824 2962 1826 2977
rect 1862 2973 1863 2977
rect 1867 2973 1868 2977
rect 1862 2972 1868 2973
rect 1870 2963 1876 2964
rect 998 2958 1004 2959
rect 1822 2961 1828 2962
rect 1822 2957 1823 2961
rect 1827 2957 1828 2961
rect 1822 2956 1828 2957
rect 1862 2960 1868 2961
rect 1862 2956 1863 2960
rect 1867 2956 1868 2960
rect 1870 2959 1871 2963
rect 1875 2959 1876 2963
rect 1870 2958 1876 2959
rect 1954 2963 1960 2964
rect 1954 2959 1955 2963
rect 1959 2959 1960 2963
rect 1954 2958 1960 2959
rect 2042 2963 2048 2964
rect 2042 2959 2043 2963
rect 2047 2959 2048 2963
rect 2042 2958 2048 2959
rect 2130 2963 2136 2964
rect 2130 2959 2131 2963
rect 2135 2959 2136 2963
rect 2130 2958 2136 2959
rect 2218 2963 2224 2964
rect 2218 2959 2219 2963
rect 2223 2959 2224 2963
rect 2218 2958 2224 2959
rect 2306 2963 2312 2964
rect 2306 2959 2307 2963
rect 2311 2959 2312 2963
rect 2306 2958 2312 2959
rect 2418 2963 2424 2964
rect 2418 2959 2419 2963
rect 2423 2959 2424 2963
rect 2418 2958 2424 2959
rect 2530 2963 2536 2964
rect 2530 2959 2531 2963
rect 2535 2959 2536 2963
rect 2530 2958 2536 2959
rect 1862 2955 1868 2956
rect 1406 2947 1412 2948
rect 1406 2943 1407 2947
rect 1411 2943 1412 2947
rect 1406 2942 1412 2943
rect 1414 2947 1420 2948
rect 1414 2943 1415 2947
rect 1419 2943 1420 2947
rect 1414 2942 1420 2943
rect 1490 2947 1496 2948
rect 1490 2943 1491 2947
rect 1495 2943 1496 2947
rect 1490 2942 1496 2943
rect 1594 2947 1600 2948
rect 1594 2943 1595 2947
rect 1599 2943 1600 2947
rect 1594 2942 1600 2943
rect 1822 2944 1828 2945
rect 1070 2931 1076 2932
rect 1070 2927 1071 2931
rect 1075 2927 1076 2931
rect 1070 2926 1076 2927
rect 1198 2931 1204 2932
rect 1198 2927 1199 2931
rect 1203 2927 1204 2931
rect 1198 2926 1204 2927
rect 1318 2931 1324 2932
rect 1318 2927 1319 2931
rect 1323 2927 1324 2931
rect 1318 2926 1324 2927
rect 946 2919 952 2920
rect 946 2915 947 2919
rect 951 2915 952 2919
rect 1072 2915 1074 2926
rect 1119 2924 1123 2925
rect 1118 2919 1124 2920
rect 1118 2915 1119 2919
rect 1123 2915 1124 2919
rect 1200 2915 1202 2926
rect 1320 2915 1322 2926
rect 463 2914 467 2915
rect 474 2914 480 2915
rect 519 2914 523 2915
rect 463 2909 467 2910
rect 519 2909 523 2910
rect 631 2914 635 2915
rect 631 2909 635 2910
rect 711 2914 715 2915
rect 711 2909 715 2910
rect 791 2914 795 2915
rect 791 2909 795 2910
rect 895 2914 899 2915
rect 895 2909 899 2910
rect 935 2914 939 2915
rect 946 2914 952 2915
rect 1071 2914 1075 2915
rect 1118 2914 1124 2915
rect 1199 2914 1203 2915
rect 935 2909 939 2910
rect 1071 2909 1075 2910
rect 1199 2909 1203 2910
rect 1239 2914 1243 2915
rect 1239 2909 1243 2910
rect 1319 2914 1323 2915
rect 1319 2909 1323 2910
rect 1399 2914 1403 2915
rect 1399 2909 1403 2910
rect 354 2907 360 2908
rect 354 2903 355 2907
rect 359 2903 360 2907
rect 354 2902 360 2903
rect 520 2898 522 2909
rect 712 2898 714 2909
rect 778 2907 784 2908
rect 778 2903 779 2907
rect 783 2903 784 2907
rect 778 2902 784 2903
rect 318 2897 324 2898
rect 318 2893 319 2897
rect 323 2893 324 2897
rect 318 2892 324 2893
rect 518 2897 524 2898
rect 518 2893 519 2897
rect 523 2893 524 2897
rect 518 2892 524 2893
rect 710 2897 716 2898
rect 710 2893 711 2897
rect 715 2893 716 2897
rect 710 2892 716 2893
rect 780 2880 782 2902
rect 896 2898 898 2909
rect 902 2907 908 2908
rect 902 2903 903 2907
rect 907 2903 908 2907
rect 902 2902 908 2903
rect 894 2897 900 2898
rect 894 2893 895 2897
rect 899 2893 900 2897
rect 894 2892 900 2893
rect 110 2879 116 2880
rect 234 2879 240 2880
rect 234 2875 235 2879
rect 239 2875 240 2879
rect 234 2874 240 2875
rect 778 2879 784 2880
rect 778 2875 779 2879
rect 783 2875 784 2879
rect 778 2874 784 2875
rect 110 2867 116 2868
rect 110 2863 111 2867
rect 115 2863 116 2867
rect 110 2862 116 2863
rect 112 2843 114 2862
rect 134 2857 140 2858
rect 134 2853 135 2857
rect 139 2853 140 2857
rect 134 2852 140 2853
rect 310 2857 316 2858
rect 310 2853 311 2857
rect 315 2853 316 2857
rect 310 2852 316 2853
rect 510 2857 516 2858
rect 510 2853 511 2857
rect 515 2853 516 2857
rect 510 2852 516 2853
rect 702 2857 708 2858
rect 702 2853 703 2857
rect 707 2853 708 2857
rect 702 2852 708 2853
rect 886 2857 892 2858
rect 886 2853 887 2857
rect 891 2853 892 2857
rect 886 2852 892 2853
rect 136 2843 138 2852
rect 178 2851 184 2852
rect 178 2847 179 2851
rect 183 2847 184 2851
rect 178 2846 184 2847
rect 111 2842 115 2843
rect 111 2837 115 2838
rect 135 2842 139 2843
rect 135 2837 139 2838
rect 159 2842 163 2843
rect 159 2837 163 2838
rect 112 2822 114 2837
rect 160 2832 162 2837
rect 158 2831 164 2832
rect 158 2827 159 2831
rect 163 2827 164 2831
rect 158 2826 164 2827
rect 110 2821 116 2822
rect 110 2817 111 2821
rect 115 2817 116 2821
rect 110 2816 116 2817
rect 110 2804 116 2805
rect 110 2800 111 2804
rect 115 2800 116 2804
rect 110 2799 116 2800
rect 112 2767 114 2799
rect 166 2791 172 2792
rect 166 2787 167 2791
rect 171 2787 172 2791
rect 166 2786 172 2787
rect 168 2767 170 2786
rect 180 2780 182 2846
rect 312 2843 314 2852
rect 512 2843 514 2852
rect 704 2843 706 2852
rect 888 2843 890 2852
rect 311 2842 315 2843
rect 311 2837 315 2838
rect 319 2842 323 2843
rect 319 2837 323 2838
rect 487 2842 491 2843
rect 487 2837 491 2838
rect 511 2842 515 2843
rect 511 2837 515 2838
rect 655 2842 659 2843
rect 655 2837 659 2838
rect 703 2842 707 2843
rect 703 2837 707 2838
rect 823 2842 827 2843
rect 823 2837 827 2838
rect 887 2842 891 2843
rect 887 2837 891 2838
rect 320 2832 322 2837
rect 488 2832 490 2837
rect 656 2832 658 2837
rect 824 2832 826 2837
rect 318 2831 324 2832
rect 318 2827 319 2831
rect 323 2827 324 2831
rect 318 2826 324 2827
rect 486 2831 492 2832
rect 486 2827 487 2831
rect 491 2827 492 2831
rect 486 2826 492 2827
rect 654 2831 660 2832
rect 654 2827 655 2831
rect 659 2827 660 2831
rect 654 2826 660 2827
rect 822 2831 828 2832
rect 822 2827 823 2831
rect 827 2827 828 2831
rect 822 2826 828 2827
rect 904 2824 906 2902
rect 1072 2898 1074 2909
rect 1118 2907 1124 2908
rect 1118 2903 1119 2907
rect 1123 2903 1124 2907
rect 1118 2902 1124 2903
rect 1162 2907 1168 2908
rect 1162 2903 1163 2907
rect 1167 2903 1168 2907
rect 1162 2902 1168 2903
rect 1070 2897 1076 2898
rect 1070 2893 1071 2897
rect 1075 2893 1076 2897
rect 1120 2893 1122 2902
rect 1070 2892 1076 2893
rect 1119 2892 1123 2893
rect 1119 2887 1123 2888
rect 1164 2884 1166 2902
rect 1240 2898 1242 2909
rect 1400 2898 1402 2909
rect 1408 2908 1410 2942
rect 1416 2925 1418 2942
rect 1430 2931 1436 2932
rect 1430 2927 1431 2931
rect 1435 2927 1436 2931
rect 1430 2926 1436 2927
rect 1415 2924 1419 2925
rect 1415 2919 1419 2920
rect 1432 2915 1434 2926
rect 1492 2920 1494 2942
rect 1534 2931 1540 2932
rect 1534 2927 1535 2931
rect 1539 2927 1540 2931
rect 1534 2926 1540 2927
rect 1490 2919 1496 2920
rect 1490 2915 1491 2919
rect 1495 2915 1496 2919
rect 1536 2915 1538 2926
rect 1596 2920 1598 2942
rect 1822 2940 1823 2944
rect 1827 2940 1828 2944
rect 1822 2939 1828 2940
rect 1646 2931 1652 2932
rect 1646 2927 1647 2931
rect 1651 2927 1652 2931
rect 1646 2926 1652 2927
rect 1734 2931 1740 2932
rect 1734 2927 1735 2931
rect 1739 2927 1740 2931
rect 1734 2926 1740 2927
rect 1594 2919 1600 2920
rect 1594 2915 1595 2919
rect 1599 2915 1600 2919
rect 1648 2915 1650 2926
rect 1736 2915 1738 2926
rect 1824 2915 1826 2939
rect 1864 2923 1866 2955
rect 1863 2922 1867 2923
rect 1872 2920 1874 2958
rect 1894 2947 1900 2948
rect 1894 2943 1895 2947
rect 1899 2943 1900 2947
rect 1894 2942 1900 2943
rect 1896 2923 1898 2942
rect 1956 2936 1958 2958
rect 1982 2947 1988 2948
rect 1982 2943 1983 2947
rect 1987 2943 1988 2947
rect 1982 2942 1988 2943
rect 1954 2935 1960 2936
rect 1954 2931 1955 2935
rect 1959 2931 1960 2935
rect 1954 2930 1960 2931
rect 1984 2923 1986 2942
rect 2044 2936 2046 2958
rect 2070 2947 2076 2948
rect 2070 2943 2071 2947
rect 2075 2943 2076 2947
rect 2070 2942 2076 2943
rect 2042 2935 2048 2936
rect 2042 2931 2043 2935
rect 2047 2931 2048 2935
rect 2042 2930 2048 2931
rect 2072 2923 2074 2942
rect 2132 2936 2134 2958
rect 2158 2947 2164 2948
rect 2158 2943 2159 2947
rect 2163 2943 2164 2947
rect 2158 2942 2164 2943
rect 2130 2935 2136 2936
rect 2130 2931 2131 2935
rect 2135 2931 2136 2935
rect 2130 2930 2136 2931
rect 2160 2923 2162 2942
rect 2220 2936 2222 2958
rect 2246 2947 2252 2948
rect 2246 2943 2247 2947
rect 2251 2943 2252 2947
rect 2246 2942 2252 2943
rect 2218 2935 2224 2936
rect 2218 2931 2219 2935
rect 2223 2931 2224 2935
rect 2218 2930 2224 2931
rect 2248 2923 2250 2942
rect 2308 2936 2310 2958
rect 2358 2947 2364 2948
rect 2358 2943 2359 2947
rect 2363 2943 2364 2947
rect 2358 2942 2364 2943
rect 2306 2935 2312 2936
rect 2306 2931 2307 2935
rect 2311 2931 2312 2935
rect 2306 2930 2312 2931
rect 2360 2923 2362 2942
rect 2420 2936 2422 2958
rect 2470 2947 2476 2948
rect 2470 2943 2471 2947
rect 2475 2943 2476 2947
rect 2470 2942 2476 2943
rect 2418 2935 2424 2936
rect 2418 2931 2419 2935
rect 2423 2931 2424 2935
rect 2418 2930 2424 2931
rect 2472 2923 2474 2942
rect 2532 2936 2534 2958
rect 2582 2947 2588 2948
rect 2582 2943 2583 2947
rect 2587 2943 2588 2947
rect 2582 2942 2588 2943
rect 2530 2935 2536 2936
rect 2530 2931 2531 2935
rect 2535 2931 2536 2935
rect 2530 2930 2536 2931
rect 2584 2923 2586 2942
rect 2596 2936 2598 3026
rect 2670 3021 2676 3022
rect 2670 3017 2671 3021
rect 2675 3017 2676 3021
rect 2670 3016 2676 3017
rect 2822 3021 2828 3022
rect 2822 3017 2823 3021
rect 2827 3017 2828 3021
rect 2822 3016 2828 3017
rect 2672 2999 2674 3016
rect 2706 3015 2712 3016
rect 2706 3011 2707 3015
rect 2711 3011 2712 3015
rect 2706 3010 2712 3011
rect 2671 2998 2675 2999
rect 2671 2993 2675 2994
rect 2687 2998 2691 2999
rect 2687 2993 2691 2994
rect 2688 2988 2690 2993
rect 2686 2987 2692 2988
rect 2686 2983 2687 2987
rect 2691 2983 2692 2987
rect 2686 2982 2692 2983
rect 2694 2947 2700 2948
rect 2694 2943 2695 2947
rect 2699 2943 2700 2947
rect 2694 2942 2700 2943
rect 2594 2935 2600 2936
rect 2594 2931 2595 2935
rect 2599 2931 2600 2935
rect 2594 2930 2600 2931
rect 2696 2923 2698 2942
rect 2708 2936 2710 3010
rect 2824 2999 2826 3016
rect 2799 2998 2803 2999
rect 2799 2993 2803 2994
rect 2823 2998 2827 2999
rect 2823 2993 2827 2994
rect 2800 2988 2802 2993
rect 2798 2987 2804 2988
rect 2798 2983 2799 2987
rect 2803 2983 2804 2987
rect 2798 2982 2804 2983
rect 2868 2980 2870 3066
rect 2976 3062 2978 3073
rect 3112 3062 3114 3073
rect 3120 3072 3122 3110
rect 3166 3099 3172 3100
rect 3166 3095 3167 3099
rect 3171 3095 3172 3099
rect 3166 3094 3172 3095
rect 3278 3099 3284 3100
rect 3278 3095 3279 3099
rect 3283 3095 3284 3099
rect 3278 3094 3284 3095
rect 3390 3099 3396 3100
rect 3390 3095 3391 3099
rect 3395 3095 3396 3099
rect 3390 3094 3396 3095
rect 3168 3079 3170 3094
rect 3178 3087 3184 3088
rect 3178 3083 3179 3087
rect 3183 3083 3184 3087
rect 3178 3082 3184 3083
rect 3167 3078 3171 3079
rect 3167 3073 3171 3074
rect 3118 3071 3124 3072
rect 3118 3067 3119 3071
rect 3123 3067 3124 3071
rect 3118 3066 3124 3067
rect 2974 3061 2980 3062
rect 2974 3057 2975 3061
rect 2979 3057 2980 3061
rect 2974 3056 2980 3057
rect 3110 3061 3116 3062
rect 3110 3057 3111 3061
rect 3115 3057 3116 3061
rect 3110 3056 3116 3057
rect 3180 3044 3182 3082
rect 3280 3079 3282 3094
rect 3392 3079 3394 3094
rect 3452 3080 3454 3126
rect 3574 3125 3575 3129
rect 3579 3125 3580 3129
rect 3574 3124 3580 3125
rect 3574 3112 3580 3113
rect 3574 3108 3575 3112
rect 3579 3108 3580 3112
rect 3574 3107 3580 3108
rect 3486 3099 3492 3100
rect 3486 3095 3487 3099
rect 3491 3095 3492 3099
rect 3486 3094 3492 3095
rect 3450 3079 3456 3080
rect 3488 3079 3490 3094
rect 3576 3079 3578 3107
rect 3239 3078 3243 3079
rect 3239 3073 3243 3074
rect 3279 3078 3283 3079
rect 3279 3073 3283 3074
rect 3375 3078 3379 3079
rect 3375 3073 3379 3074
rect 3391 3078 3395 3079
rect 3450 3075 3451 3079
rect 3455 3075 3456 3079
rect 3450 3074 3456 3075
rect 3487 3078 3491 3079
rect 3391 3073 3395 3074
rect 3487 3073 3491 3074
rect 3575 3078 3579 3079
rect 3575 3073 3579 3074
rect 3240 3062 3242 3073
rect 3358 3071 3364 3072
rect 3358 3067 3359 3071
rect 3363 3067 3364 3071
rect 3358 3066 3364 3067
rect 3238 3061 3244 3062
rect 3238 3057 3239 3061
rect 3243 3057 3244 3061
rect 3238 3056 3244 3057
rect 3178 3043 3184 3044
rect 3178 3039 3179 3043
rect 3183 3039 3184 3043
rect 3178 3038 3184 3039
rect 2966 3021 2972 3022
rect 2966 3017 2967 3021
rect 2971 3017 2972 3021
rect 2966 3016 2972 3017
rect 3102 3021 3108 3022
rect 3102 3017 3103 3021
rect 3107 3017 3108 3021
rect 3102 3016 3108 3017
rect 3230 3021 3236 3022
rect 3230 3017 3231 3021
rect 3235 3017 3236 3021
rect 3230 3016 3236 3017
rect 2968 2999 2970 3016
rect 3104 2999 3106 3016
rect 3232 2999 3234 3016
rect 2903 2998 2907 2999
rect 2903 2993 2907 2994
rect 2967 2998 2971 2999
rect 2967 2993 2971 2994
rect 3007 2998 3011 2999
rect 3007 2993 3011 2994
rect 3103 2998 3107 2999
rect 3103 2993 3107 2994
rect 3199 2998 3203 2999
rect 3199 2993 3203 2994
rect 3231 2998 3235 2999
rect 3231 2993 3235 2994
rect 3295 2998 3299 2999
rect 3295 2993 3299 2994
rect 2904 2988 2906 2993
rect 3008 2988 3010 2993
rect 3104 2988 3106 2993
rect 3200 2988 3202 2993
rect 3296 2988 3298 2993
rect 2902 2987 2908 2988
rect 2902 2983 2903 2987
rect 2907 2983 2908 2987
rect 2902 2982 2908 2983
rect 3006 2987 3012 2988
rect 3006 2983 3007 2987
rect 3011 2983 3012 2987
rect 3006 2982 3012 2983
rect 3102 2987 3108 2988
rect 3102 2983 3103 2987
rect 3107 2983 3108 2987
rect 3102 2982 3108 2983
rect 3198 2987 3204 2988
rect 3198 2983 3199 2987
rect 3203 2983 3204 2987
rect 3198 2982 3204 2983
rect 3294 2987 3300 2988
rect 3294 2983 3295 2987
rect 3299 2983 3300 2987
rect 3360 2987 3362 3066
rect 3376 3062 3378 3073
rect 3488 3062 3490 3073
rect 3374 3061 3380 3062
rect 3374 3057 3375 3061
rect 3379 3057 3380 3061
rect 3374 3056 3380 3057
rect 3486 3061 3492 3062
rect 3486 3057 3487 3061
rect 3491 3057 3492 3061
rect 3486 3056 3492 3057
rect 3576 3049 3578 3073
rect 3574 3048 3580 3049
rect 3574 3044 3575 3048
rect 3579 3044 3580 3048
rect 3574 3043 3580 3044
rect 3574 3031 3580 3032
rect 3574 3027 3575 3031
rect 3579 3027 3580 3031
rect 3574 3026 3580 3027
rect 3366 3021 3372 3022
rect 3366 3017 3367 3021
rect 3371 3017 3372 3021
rect 3366 3016 3372 3017
rect 3478 3021 3484 3022
rect 3478 3017 3479 3021
rect 3483 3017 3484 3021
rect 3478 3016 3484 3017
rect 3368 2999 3370 3016
rect 3480 2999 3482 3016
rect 3498 3015 3504 3016
rect 3498 3011 3499 3015
rect 3503 3011 3504 3015
rect 3498 3010 3504 3011
rect 3367 2998 3371 2999
rect 3367 2993 3371 2994
rect 3391 2998 3395 2999
rect 3391 2993 3395 2994
rect 3479 2998 3483 2999
rect 3479 2993 3483 2994
rect 3392 2988 3394 2993
rect 3480 2988 3482 2993
rect 3390 2987 3396 2988
rect 3360 2985 3366 2987
rect 3294 2982 3300 2983
rect 3364 2980 3366 2985
rect 3390 2983 3391 2987
rect 3395 2983 3396 2987
rect 3390 2982 3396 2983
rect 3478 2987 3484 2988
rect 3478 2983 3479 2987
rect 3483 2983 3484 2987
rect 3478 2982 3484 2983
rect 2866 2979 2872 2980
rect 2866 2975 2867 2979
rect 2871 2975 2872 2979
rect 2866 2974 2872 2975
rect 3362 2979 3368 2980
rect 3362 2975 3363 2979
rect 3367 2975 3368 2979
rect 3362 2974 3368 2975
rect 2806 2947 2812 2948
rect 2806 2943 2807 2947
rect 2811 2943 2812 2947
rect 2806 2942 2812 2943
rect 2910 2947 2916 2948
rect 2910 2943 2911 2947
rect 2915 2943 2916 2947
rect 2910 2942 2916 2943
rect 3014 2947 3020 2948
rect 3014 2943 3015 2947
rect 3019 2943 3020 2947
rect 3014 2942 3020 2943
rect 3110 2947 3116 2948
rect 3110 2943 3111 2947
rect 3115 2943 3116 2947
rect 3110 2942 3116 2943
rect 3206 2947 3212 2948
rect 3206 2943 3207 2947
rect 3211 2943 3212 2947
rect 3206 2942 3212 2943
rect 3302 2947 3308 2948
rect 3302 2943 3303 2947
rect 3307 2943 3308 2947
rect 3302 2942 3308 2943
rect 3398 2947 3404 2948
rect 3398 2943 3399 2947
rect 3403 2943 3404 2947
rect 3398 2942 3404 2943
rect 3486 2947 3492 2948
rect 3486 2943 3487 2947
rect 3491 2943 3492 2947
rect 3486 2942 3492 2943
rect 2706 2935 2712 2936
rect 2706 2931 2707 2935
rect 2711 2931 2712 2935
rect 2706 2930 2712 2931
rect 2808 2923 2810 2942
rect 2912 2923 2914 2942
rect 2954 2935 2960 2936
rect 2954 2931 2955 2935
rect 2959 2931 2960 2935
rect 2954 2930 2960 2931
rect 1895 2922 1899 2923
rect 1863 2917 1867 2918
rect 1870 2919 1876 2920
rect 1431 2914 1435 2915
rect 1490 2914 1496 2915
rect 1535 2914 1539 2915
rect 1431 2909 1435 2910
rect 1535 2909 1539 2910
rect 1551 2914 1555 2915
rect 1594 2914 1600 2915
rect 1647 2914 1651 2915
rect 1551 2909 1555 2910
rect 1647 2909 1651 2910
rect 1711 2914 1715 2915
rect 1711 2909 1715 2910
rect 1735 2914 1739 2915
rect 1735 2909 1739 2910
rect 1823 2914 1827 2915
rect 1823 2909 1827 2910
rect 1406 2907 1412 2908
rect 1406 2903 1407 2907
rect 1411 2903 1412 2907
rect 1406 2902 1412 2903
rect 1552 2898 1554 2909
rect 1651 2900 1655 2901
rect 1238 2897 1244 2898
rect 1238 2893 1239 2897
rect 1243 2893 1244 2897
rect 1238 2892 1244 2893
rect 1398 2897 1404 2898
rect 1398 2893 1399 2897
rect 1403 2893 1404 2897
rect 1398 2892 1404 2893
rect 1550 2897 1556 2898
rect 1550 2893 1551 2897
rect 1555 2893 1556 2897
rect 1712 2898 1714 2909
rect 1651 2895 1655 2896
rect 1710 2897 1716 2898
rect 1550 2892 1556 2893
rect 1162 2883 1168 2884
rect 1162 2879 1163 2883
rect 1167 2879 1168 2883
rect 1652 2880 1654 2895
rect 1710 2893 1711 2897
rect 1715 2893 1716 2897
rect 1710 2892 1716 2893
rect 1824 2885 1826 2909
rect 1864 2893 1866 2917
rect 1870 2915 1871 2919
rect 1875 2915 1876 2919
rect 1895 2917 1899 2918
rect 1983 2922 1987 2923
rect 1983 2917 1987 2918
rect 2071 2922 2075 2923
rect 2071 2917 2075 2918
rect 2159 2922 2163 2923
rect 2159 2917 2163 2918
rect 2247 2922 2251 2923
rect 2247 2917 2251 2918
rect 2359 2922 2363 2923
rect 2359 2917 2363 2918
rect 2471 2922 2475 2923
rect 2471 2917 2475 2918
rect 2583 2922 2587 2923
rect 2583 2917 2587 2918
rect 2695 2922 2699 2923
rect 2695 2917 2699 2918
rect 2807 2922 2811 2923
rect 2807 2917 2811 2918
rect 2895 2922 2899 2923
rect 2895 2917 2899 2918
rect 2911 2922 2915 2923
rect 2911 2917 2915 2918
rect 1870 2914 1876 2915
rect 2896 2906 2898 2917
rect 2894 2905 2900 2906
rect 2894 2901 2895 2905
rect 2899 2901 2900 2905
rect 2894 2900 2900 2901
rect 1862 2892 1868 2893
rect 2956 2892 2958 2930
rect 3016 2923 3018 2942
rect 3112 2923 3114 2942
rect 3208 2923 3210 2942
rect 3304 2923 3306 2942
rect 3400 2923 3402 2942
rect 3488 2923 3490 2942
rect 3500 2936 3502 3010
rect 3576 2999 3578 3026
rect 3575 2998 3579 2999
rect 3575 2993 3579 2994
rect 3576 2978 3578 2993
rect 3574 2977 3580 2978
rect 3574 2973 3575 2977
rect 3579 2973 3580 2977
rect 3574 2972 3580 2973
rect 3574 2960 3580 2961
rect 3574 2956 3575 2960
rect 3579 2956 3580 2960
rect 3574 2955 3580 2956
rect 3498 2935 3504 2936
rect 3498 2931 3499 2935
rect 3503 2931 3504 2935
rect 3498 2930 3504 2931
rect 3576 2923 3578 2955
rect 3015 2922 3019 2923
rect 3015 2917 3019 2918
rect 3111 2922 3115 2923
rect 3111 2917 3115 2918
rect 3199 2922 3203 2923
rect 3199 2917 3203 2918
rect 3207 2922 3211 2923
rect 3207 2917 3211 2918
rect 3303 2922 3307 2923
rect 3303 2917 3307 2918
rect 3399 2922 3403 2923
rect 3399 2917 3403 2918
rect 3487 2922 3491 2923
rect 3487 2917 3491 2918
rect 3575 2922 3579 2923
rect 3575 2917 3579 2918
rect 3162 2915 3168 2916
rect 3162 2911 3163 2915
rect 3167 2911 3168 2915
rect 3162 2910 3168 2911
rect 1862 2888 1863 2892
rect 1867 2888 1868 2892
rect 1862 2887 1868 2888
rect 2954 2891 2960 2892
rect 2954 2887 2955 2891
rect 2959 2887 2960 2891
rect 2954 2886 2960 2887
rect 1822 2884 1828 2885
rect 1822 2880 1823 2884
rect 1827 2880 1828 2884
rect 1162 2878 1168 2879
rect 1650 2879 1656 2880
rect 1822 2879 1828 2880
rect 1650 2875 1651 2879
rect 1655 2875 1656 2879
rect 1650 2874 1656 2875
rect 1862 2875 1868 2876
rect 1862 2871 1863 2875
rect 1867 2871 1868 2875
rect 1862 2870 1868 2871
rect 1822 2867 1828 2868
rect 1822 2863 1823 2867
rect 1827 2863 1828 2867
rect 1822 2862 1828 2863
rect 1062 2857 1068 2858
rect 1062 2853 1063 2857
rect 1067 2853 1068 2857
rect 1062 2852 1068 2853
rect 1230 2857 1236 2858
rect 1230 2853 1231 2857
rect 1235 2853 1236 2857
rect 1230 2852 1236 2853
rect 1390 2857 1396 2858
rect 1390 2853 1391 2857
rect 1395 2853 1396 2857
rect 1390 2852 1396 2853
rect 1542 2857 1548 2858
rect 1542 2853 1543 2857
rect 1547 2853 1548 2857
rect 1542 2852 1548 2853
rect 1702 2857 1708 2858
rect 1702 2853 1703 2857
rect 1707 2853 1708 2857
rect 1702 2852 1708 2853
rect 1064 2843 1066 2852
rect 1232 2843 1234 2852
rect 1290 2851 1296 2852
rect 1290 2847 1291 2851
rect 1295 2847 1296 2851
rect 1290 2846 1296 2847
rect 975 2842 979 2843
rect 975 2837 979 2838
rect 1063 2842 1067 2843
rect 1063 2837 1067 2838
rect 1127 2842 1131 2843
rect 1127 2837 1131 2838
rect 1231 2842 1235 2843
rect 1231 2837 1235 2838
rect 1271 2842 1275 2843
rect 1271 2837 1275 2838
rect 976 2832 978 2837
rect 1128 2832 1130 2837
rect 1272 2832 1274 2837
rect 974 2831 980 2832
rect 974 2827 975 2831
rect 979 2827 980 2831
rect 974 2826 980 2827
rect 1126 2831 1132 2832
rect 1126 2827 1127 2831
rect 1131 2827 1132 2831
rect 1126 2826 1132 2827
rect 1270 2831 1276 2832
rect 1270 2827 1271 2831
rect 1275 2827 1276 2831
rect 1270 2826 1276 2827
rect 902 2823 908 2824
rect 902 2819 903 2823
rect 907 2819 908 2823
rect 902 2818 908 2819
rect 250 2807 256 2808
rect 250 2803 251 2807
rect 255 2803 256 2807
rect 250 2802 256 2803
rect 386 2807 392 2808
rect 386 2803 387 2807
rect 391 2803 392 2807
rect 386 2802 392 2803
rect 252 2780 254 2802
rect 326 2791 332 2792
rect 326 2787 327 2791
rect 331 2787 332 2791
rect 326 2786 332 2787
rect 178 2779 184 2780
rect 178 2775 179 2779
rect 183 2775 184 2779
rect 178 2774 184 2775
rect 250 2779 256 2780
rect 250 2775 251 2779
rect 255 2775 256 2779
rect 250 2774 256 2775
rect 328 2767 330 2786
rect 111 2766 115 2767
rect 111 2761 115 2762
rect 167 2766 171 2767
rect 167 2761 171 2762
rect 207 2766 211 2767
rect 207 2761 211 2762
rect 327 2766 331 2767
rect 327 2761 331 2762
rect 335 2766 339 2767
rect 335 2761 339 2762
rect 112 2737 114 2761
rect 208 2750 210 2761
rect 302 2759 308 2760
rect 302 2755 303 2759
rect 307 2755 308 2759
rect 302 2754 308 2755
rect 206 2749 212 2750
rect 206 2745 207 2749
rect 211 2745 212 2749
rect 206 2744 212 2745
rect 110 2736 116 2737
rect 110 2732 111 2736
rect 115 2732 116 2736
rect 304 2732 306 2754
rect 336 2750 338 2761
rect 388 2760 390 2802
rect 494 2791 500 2792
rect 494 2787 495 2791
rect 499 2787 500 2791
rect 494 2786 500 2787
rect 662 2791 668 2792
rect 662 2787 663 2791
rect 667 2787 668 2791
rect 662 2786 668 2787
rect 830 2791 836 2792
rect 830 2787 831 2791
rect 835 2787 836 2791
rect 830 2786 836 2787
rect 982 2791 988 2792
rect 982 2787 983 2791
rect 987 2787 988 2791
rect 1134 2791 1140 2792
rect 982 2786 988 2787
rect 995 2788 999 2789
rect 496 2767 498 2786
rect 530 2779 536 2780
rect 530 2775 531 2779
rect 535 2775 536 2779
rect 530 2774 536 2775
rect 471 2766 475 2767
rect 471 2761 475 2762
rect 495 2766 499 2767
rect 495 2761 499 2762
rect 386 2759 392 2760
rect 386 2755 387 2759
rect 391 2755 392 2759
rect 386 2754 392 2755
rect 472 2750 474 2761
rect 334 2749 340 2750
rect 334 2745 335 2749
rect 339 2745 340 2749
rect 334 2744 340 2745
rect 470 2749 476 2750
rect 470 2745 471 2749
rect 475 2745 476 2749
rect 470 2744 476 2745
rect 532 2736 534 2774
rect 664 2767 666 2786
rect 832 2767 834 2786
rect 984 2767 986 2786
rect 1134 2787 1135 2791
rect 1139 2787 1140 2791
rect 1134 2786 1140 2787
rect 1278 2791 1284 2792
rect 1278 2787 1279 2791
rect 1283 2787 1284 2791
rect 1278 2786 1284 2787
rect 995 2783 999 2784
rect 996 2780 998 2783
rect 994 2779 1000 2780
rect 994 2775 995 2779
rect 999 2775 1000 2779
rect 994 2774 1000 2775
rect 1136 2767 1138 2786
rect 1280 2767 1282 2786
rect 1292 2780 1294 2846
rect 1392 2843 1394 2852
rect 1544 2843 1546 2852
rect 1704 2843 1706 2852
rect 1824 2843 1826 2862
rect 1864 2855 1866 2870
rect 2886 2865 2892 2866
rect 2886 2861 2887 2865
rect 2891 2861 2892 2865
rect 2886 2860 2892 2861
rect 2888 2855 2890 2860
rect 1863 2854 1867 2855
rect 1863 2849 1867 2850
rect 2831 2854 2835 2855
rect 2831 2849 2835 2850
rect 2887 2854 2891 2855
rect 2887 2849 2891 2850
rect 2919 2854 2923 2855
rect 2919 2849 2923 2850
rect 3007 2854 3011 2855
rect 3007 2849 3011 2850
rect 3095 2854 3099 2855
rect 3095 2849 3099 2850
rect 1391 2842 1395 2843
rect 1391 2837 1395 2838
rect 1415 2842 1419 2843
rect 1415 2837 1419 2838
rect 1543 2842 1547 2843
rect 1543 2837 1547 2838
rect 1559 2842 1563 2843
rect 1559 2837 1563 2838
rect 1703 2842 1707 2843
rect 1703 2837 1707 2838
rect 1823 2842 1827 2843
rect 1823 2837 1827 2838
rect 1416 2832 1418 2837
rect 1560 2832 1562 2837
rect 1414 2831 1420 2832
rect 1414 2827 1415 2831
rect 1419 2827 1420 2831
rect 1414 2826 1420 2827
rect 1558 2831 1564 2832
rect 1558 2827 1559 2831
rect 1563 2827 1564 2831
rect 1558 2826 1564 2827
rect 1482 2823 1488 2824
rect 1482 2819 1483 2823
rect 1487 2819 1488 2823
rect 1824 2822 1826 2837
rect 1864 2834 1866 2849
rect 2832 2844 2834 2849
rect 2920 2844 2922 2849
rect 3008 2844 3010 2849
rect 3096 2844 3098 2849
rect 2830 2843 2836 2844
rect 2830 2839 2831 2843
rect 2835 2839 2836 2843
rect 2830 2838 2836 2839
rect 2918 2843 2924 2844
rect 2918 2839 2919 2843
rect 2923 2839 2924 2843
rect 2918 2838 2924 2839
rect 3006 2843 3012 2844
rect 3006 2839 3007 2843
rect 3011 2839 3012 2843
rect 3006 2838 3012 2839
rect 3094 2843 3100 2844
rect 3094 2839 3095 2843
rect 3099 2839 3100 2843
rect 3094 2838 3100 2839
rect 3164 2836 3166 2910
rect 3200 2906 3202 2917
rect 3488 2906 3490 2917
rect 3198 2905 3204 2906
rect 3198 2901 3199 2905
rect 3203 2901 3204 2905
rect 3198 2900 3204 2901
rect 3486 2905 3492 2906
rect 3486 2901 3487 2905
rect 3491 2901 3492 2905
rect 3486 2900 3492 2901
rect 3576 2893 3578 2917
rect 3574 2892 3580 2893
rect 3574 2888 3575 2892
rect 3579 2888 3580 2892
rect 3574 2887 3580 2888
rect 3574 2875 3580 2876
rect 3574 2871 3575 2875
rect 3579 2871 3580 2875
rect 3574 2870 3580 2871
rect 3190 2865 3196 2866
rect 3190 2861 3191 2865
rect 3195 2861 3196 2865
rect 3190 2860 3196 2861
rect 3478 2865 3484 2866
rect 3478 2861 3479 2865
rect 3483 2861 3484 2865
rect 3478 2860 3484 2861
rect 3192 2855 3194 2860
rect 3480 2855 3482 2860
rect 3498 2859 3504 2860
rect 3498 2855 3499 2859
rect 3503 2855 3504 2859
rect 3576 2855 3578 2870
rect 3191 2854 3195 2855
rect 3191 2849 3195 2850
rect 3479 2854 3483 2855
rect 3498 2854 3504 2855
rect 3575 2854 3579 2855
rect 3479 2849 3483 2850
rect 3162 2835 3168 2836
rect 1862 2833 1868 2834
rect 1862 2829 1863 2833
rect 1867 2829 1868 2833
rect 3162 2831 3163 2835
rect 3167 2831 3168 2835
rect 3162 2830 3168 2831
rect 1862 2828 1868 2829
rect 1482 2818 1488 2819
rect 1822 2821 1828 2822
rect 1422 2791 1428 2792
rect 1422 2787 1423 2791
rect 1427 2787 1428 2791
rect 1484 2789 1486 2818
rect 1822 2817 1823 2821
rect 1827 2817 1828 2821
rect 2898 2819 2904 2820
rect 1822 2816 1828 2817
rect 1862 2816 1868 2817
rect 1862 2812 1863 2816
rect 1867 2812 1868 2816
rect 2898 2815 2899 2819
rect 2903 2815 2904 2819
rect 2898 2814 2904 2815
rect 2986 2819 2992 2820
rect 2986 2815 2987 2819
rect 2991 2815 2992 2819
rect 2986 2814 2992 2815
rect 3074 2819 3080 2820
rect 3074 2815 3075 2819
rect 3079 2815 3080 2819
rect 3074 2814 3080 2815
rect 1862 2811 1868 2812
rect 1822 2804 1828 2805
rect 1822 2800 1823 2804
rect 1827 2800 1828 2804
rect 1822 2799 1828 2800
rect 1566 2791 1572 2792
rect 1422 2786 1428 2787
rect 1483 2788 1487 2789
rect 1290 2779 1296 2780
rect 1290 2775 1291 2779
rect 1295 2775 1296 2779
rect 1290 2774 1296 2775
rect 1424 2767 1426 2786
rect 1566 2787 1567 2791
rect 1571 2787 1572 2791
rect 1566 2786 1572 2787
rect 1483 2783 1487 2784
rect 1568 2767 1570 2786
rect 1824 2767 1826 2799
rect 1864 2787 1866 2811
rect 2838 2803 2844 2804
rect 2838 2799 2839 2803
rect 2843 2799 2844 2803
rect 2838 2798 2844 2799
rect 2840 2787 2842 2798
rect 2900 2792 2902 2814
rect 2926 2803 2932 2804
rect 2926 2799 2927 2803
rect 2931 2799 2932 2803
rect 2926 2798 2932 2799
rect 2850 2791 2856 2792
rect 2850 2787 2851 2791
rect 2855 2787 2856 2791
rect 1863 2786 1867 2787
rect 1863 2781 1867 2782
rect 2671 2786 2675 2787
rect 2671 2781 2675 2782
rect 2807 2786 2811 2787
rect 2807 2781 2811 2782
rect 2839 2786 2843 2787
rect 2850 2786 2856 2787
rect 2898 2791 2904 2792
rect 2898 2787 2899 2791
rect 2903 2787 2904 2791
rect 2928 2787 2930 2798
rect 2988 2792 2990 2814
rect 3014 2803 3020 2804
rect 3014 2799 3015 2803
rect 3019 2799 3020 2803
rect 3014 2798 3020 2799
rect 2986 2791 2992 2792
rect 2986 2787 2987 2791
rect 2991 2787 2992 2791
rect 3016 2787 3018 2798
rect 3076 2792 3078 2814
rect 3102 2803 3108 2804
rect 3102 2799 3103 2803
rect 3107 2799 3108 2803
rect 3102 2798 3108 2799
rect 3074 2791 3080 2792
rect 3074 2787 3075 2791
rect 3079 2787 3080 2791
rect 3104 2787 3106 2798
rect 2898 2786 2904 2787
rect 2927 2786 2931 2787
rect 2839 2781 2843 2782
rect 607 2766 611 2767
rect 607 2761 611 2762
rect 663 2766 667 2767
rect 663 2761 667 2762
rect 751 2766 755 2767
rect 751 2761 755 2762
rect 831 2766 835 2767
rect 831 2761 835 2762
rect 887 2766 891 2767
rect 887 2761 891 2762
rect 983 2766 987 2767
rect 983 2761 987 2762
rect 1023 2766 1027 2767
rect 1023 2761 1027 2762
rect 1135 2766 1139 2767
rect 1135 2761 1139 2762
rect 1151 2766 1155 2767
rect 1151 2761 1155 2762
rect 1279 2766 1283 2767
rect 1279 2761 1283 2762
rect 1287 2766 1291 2767
rect 1287 2761 1291 2762
rect 1423 2766 1427 2767
rect 1423 2761 1427 2762
rect 1567 2766 1571 2767
rect 1567 2761 1571 2762
rect 1823 2766 1827 2767
rect 1823 2761 1827 2762
rect 608 2750 610 2761
rect 650 2759 656 2760
rect 650 2755 651 2759
rect 655 2755 656 2759
rect 650 2754 656 2755
rect 606 2749 612 2750
rect 606 2745 607 2749
rect 611 2745 612 2749
rect 606 2744 612 2745
rect 530 2735 536 2736
rect 110 2731 116 2732
rect 302 2731 308 2732
rect 302 2727 303 2731
rect 307 2727 308 2731
rect 530 2731 531 2735
rect 535 2731 536 2735
rect 530 2730 536 2731
rect 302 2726 308 2727
rect 110 2719 116 2720
rect 110 2715 111 2719
rect 115 2715 116 2719
rect 110 2714 116 2715
rect 112 2695 114 2714
rect 198 2709 204 2710
rect 198 2705 199 2709
rect 203 2705 204 2709
rect 198 2704 204 2705
rect 326 2709 332 2710
rect 326 2705 327 2709
rect 331 2705 332 2709
rect 326 2704 332 2705
rect 462 2709 468 2710
rect 462 2705 463 2709
rect 467 2705 468 2709
rect 462 2704 468 2705
rect 598 2709 604 2710
rect 598 2705 599 2709
rect 603 2705 604 2709
rect 598 2704 604 2705
rect 200 2695 202 2704
rect 234 2703 240 2704
rect 234 2699 235 2703
rect 239 2699 240 2703
rect 234 2698 240 2699
rect 111 2694 115 2695
rect 111 2689 115 2690
rect 199 2694 203 2695
rect 199 2689 203 2690
rect 215 2694 219 2695
rect 215 2689 219 2690
rect 112 2674 114 2689
rect 216 2684 218 2689
rect 214 2683 220 2684
rect 214 2679 215 2683
rect 219 2679 220 2683
rect 214 2678 220 2679
rect 110 2673 116 2674
rect 110 2669 111 2673
rect 115 2669 116 2673
rect 110 2668 116 2669
rect 110 2656 116 2657
rect 110 2652 111 2656
rect 115 2652 116 2656
rect 110 2651 116 2652
rect 112 2623 114 2651
rect 222 2643 228 2644
rect 222 2639 223 2643
rect 227 2639 228 2643
rect 222 2638 228 2639
rect 224 2623 226 2638
rect 236 2632 238 2698
rect 328 2695 330 2704
rect 464 2695 466 2704
rect 600 2695 602 2704
rect 327 2694 331 2695
rect 327 2689 331 2690
rect 335 2694 339 2695
rect 335 2689 339 2690
rect 463 2694 467 2695
rect 463 2689 467 2690
rect 583 2694 587 2695
rect 583 2689 587 2690
rect 599 2694 603 2695
rect 599 2689 603 2690
rect 336 2684 338 2689
rect 464 2684 466 2689
rect 584 2684 586 2689
rect 334 2683 340 2684
rect 334 2679 335 2683
rect 339 2679 340 2683
rect 334 2678 340 2679
rect 462 2683 468 2684
rect 462 2679 463 2683
rect 467 2679 468 2683
rect 462 2678 468 2679
rect 582 2683 588 2684
rect 582 2679 583 2683
rect 587 2679 588 2683
rect 582 2678 588 2679
rect 652 2676 654 2754
rect 752 2750 754 2761
rect 888 2750 890 2761
rect 1024 2750 1026 2761
rect 1152 2750 1154 2761
rect 1288 2750 1290 2761
rect 1424 2750 1426 2761
rect 750 2749 756 2750
rect 750 2745 751 2749
rect 755 2745 756 2749
rect 750 2744 756 2745
rect 886 2749 892 2750
rect 886 2745 887 2749
rect 891 2745 892 2749
rect 886 2744 892 2745
rect 1022 2749 1028 2750
rect 1022 2745 1023 2749
rect 1027 2745 1028 2749
rect 1022 2744 1028 2745
rect 1150 2749 1156 2750
rect 1150 2745 1151 2749
rect 1155 2745 1156 2749
rect 1150 2744 1156 2745
rect 1286 2749 1292 2750
rect 1286 2745 1287 2749
rect 1291 2745 1292 2749
rect 1286 2744 1292 2745
rect 1422 2749 1428 2750
rect 1422 2745 1423 2749
rect 1427 2745 1428 2749
rect 1422 2744 1428 2745
rect 1824 2737 1826 2761
rect 1864 2757 1866 2781
rect 2672 2770 2674 2781
rect 2734 2779 2740 2780
rect 2734 2775 2735 2779
rect 2739 2775 2740 2779
rect 2734 2774 2740 2775
rect 2670 2769 2676 2770
rect 2670 2765 2671 2769
rect 2675 2765 2676 2769
rect 2670 2764 2676 2765
rect 1862 2756 1868 2757
rect 1862 2752 1863 2756
rect 1867 2752 1868 2756
rect 1862 2751 1868 2752
rect 1862 2739 1868 2740
rect 1822 2736 1828 2737
rect 1822 2732 1823 2736
rect 1827 2732 1828 2736
rect 1862 2735 1863 2739
rect 1867 2735 1868 2739
rect 1862 2734 1868 2735
rect 1822 2731 1828 2732
rect 1822 2719 1828 2720
rect 1864 2719 1866 2734
rect 2736 2733 2738 2774
rect 2808 2770 2810 2781
rect 2806 2769 2812 2770
rect 2806 2765 2807 2769
rect 2811 2765 2812 2769
rect 2852 2765 2854 2786
rect 2927 2781 2931 2782
rect 2967 2786 2971 2787
rect 2986 2786 2992 2787
rect 3015 2786 3019 2787
rect 3074 2786 3080 2787
rect 3103 2786 3107 2787
rect 2967 2781 2971 2782
rect 3015 2781 3019 2782
rect 3103 2781 3107 2782
rect 3143 2786 3147 2787
rect 3143 2781 3147 2782
rect 3327 2786 3331 2787
rect 3327 2781 3331 2782
rect 3487 2786 3491 2787
rect 3487 2781 3491 2782
rect 2968 2770 2970 2781
rect 3144 2770 3146 2781
rect 3328 2770 3330 2781
rect 3488 2770 3490 2781
rect 3500 2780 3502 2854
rect 3575 2849 3579 2850
rect 3576 2834 3578 2849
rect 3574 2833 3580 2834
rect 3574 2829 3575 2833
rect 3579 2829 3580 2833
rect 3574 2828 3580 2829
rect 3574 2816 3580 2817
rect 3574 2812 3575 2816
rect 3579 2812 3580 2816
rect 3574 2811 3580 2812
rect 3576 2787 3578 2811
rect 3575 2786 3579 2787
rect 3575 2781 3579 2782
rect 3498 2779 3504 2780
rect 3498 2775 3499 2779
rect 3503 2775 3504 2779
rect 3498 2774 3504 2775
rect 2966 2769 2972 2770
rect 2966 2765 2967 2769
rect 2971 2765 2972 2769
rect 2806 2764 2812 2765
rect 2851 2764 2855 2765
rect 2966 2764 2972 2765
rect 3142 2769 3148 2770
rect 3142 2765 3143 2769
rect 3147 2765 3148 2769
rect 3326 2769 3332 2770
rect 3326 2765 3327 2769
rect 3331 2765 3332 2769
rect 3142 2764 3148 2765
rect 3259 2764 3263 2765
rect 3326 2764 3332 2765
rect 3486 2769 3492 2770
rect 3486 2765 3487 2769
rect 3491 2765 3492 2769
rect 3486 2764 3492 2765
rect 2851 2759 2855 2760
rect 3259 2759 3263 2760
rect 3260 2752 3262 2759
rect 3576 2757 3578 2781
rect 3574 2756 3580 2757
rect 3574 2752 3575 2756
rect 3579 2752 3580 2756
rect 3258 2751 3264 2752
rect 3574 2751 3580 2752
rect 3258 2747 3259 2751
rect 3263 2747 3264 2751
rect 3258 2746 3264 2747
rect 3574 2739 3580 2740
rect 3574 2735 3575 2739
rect 3579 2735 3580 2739
rect 3574 2734 3580 2735
rect 2735 2732 2739 2733
rect 2662 2729 2668 2730
rect 2662 2725 2663 2729
rect 2667 2725 2668 2729
rect 3363 2732 3367 2733
rect 2735 2727 2739 2728
rect 2798 2729 2804 2730
rect 2662 2724 2668 2725
rect 2798 2725 2799 2729
rect 2803 2725 2804 2729
rect 2798 2724 2804 2725
rect 2958 2729 2964 2730
rect 2958 2725 2959 2729
rect 2963 2725 2964 2729
rect 2958 2724 2964 2725
rect 3134 2729 3140 2730
rect 3134 2725 3135 2729
rect 3139 2725 3140 2729
rect 3134 2724 3140 2725
rect 3318 2729 3324 2730
rect 3318 2725 3319 2729
rect 3323 2725 3324 2729
rect 3363 2727 3367 2728
rect 3478 2729 3484 2730
rect 3318 2724 3324 2725
rect 2664 2719 2666 2724
rect 2800 2719 2802 2724
rect 2960 2719 2962 2724
rect 3136 2719 3138 2724
rect 3320 2719 3322 2724
rect 1822 2715 1823 2719
rect 1827 2715 1828 2719
rect 1822 2714 1828 2715
rect 1863 2718 1867 2719
rect 742 2709 748 2710
rect 742 2705 743 2709
rect 747 2705 748 2709
rect 742 2704 748 2705
rect 878 2709 884 2710
rect 878 2705 879 2709
rect 883 2705 884 2709
rect 878 2704 884 2705
rect 1014 2709 1020 2710
rect 1014 2705 1015 2709
rect 1019 2705 1020 2709
rect 1014 2704 1020 2705
rect 1142 2709 1148 2710
rect 1142 2705 1143 2709
rect 1147 2705 1148 2709
rect 1142 2704 1148 2705
rect 1278 2709 1284 2710
rect 1278 2705 1279 2709
rect 1283 2705 1284 2709
rect 1278 2704 1284 2705
rect 1414 2709 1420 2710
rect 1414 2705 1415 2709
rect 1419 2705 1420 2709
rect 1414 2704 1420 2705
rect 744 2695 746 2704
rect 880 2695 882 2704
rect 1016 2695 1018 2704
rect 1144 2695 1146 2704
rect 1178 2703 1184 2704
rect 1178 2699 1179 2703
rect 1183 2699 1184 2703
rect 1178 2698 1184 2699
rect 703 2694 707 2695
rect 703 2689 707 2690
rect 743 2694 747 2695
rect 743 2689 747 2690
rect 823 2694 827 2695
rect 823 2689 827 2690
rect 879 2694 883 2695
rect 879 2689 883 2690
rect 935 2694 939 2695
rect 935 2689 939 2690
rect 1015 2694 1019 2695
rect 1015 2689 1019 2690
rect 1047 2694 1051 2695
rect 1047 2689 1051 2690
rect 1143 2694 1147 2695
rect 1143 2689 1147 2690
rect 1159 2694 1163 2695
rect 1159 2689 1163 2690
rect 704 2684 706 2689
rect 824 2684 826 2689
rect 936 2684 938 2689
rect 1048 2684 1050 2689
rect 1160 2684 1162 2689
rect 702 2683 708 2684
rect 702 2679 703 2683
rect 707 2679 708 2683
rect 702 2678 708 2679
rect 822 2683 828 2684
rect 822 2679 823 2683
rect 827 2679 828 2683
rect 822 2678 828 2679
rect 934 2683 940 2684
rect 934 2679 935 2683
rect 939 2679 940 2683
rect 934 2678 940 2679
rect 1046 2683 1052 2684
rect 1046 2679 1047 2683
rect 1051 2679 1052 2683
rect 1046 2678 1052 2679
rect 1158 2683 1164 2684
rect 1158 2679 1159 2683
rect 1163 2679 1164 2683
rect 1158 2678 1164 2679
rect 650 2675 656 2676
rect 650 2671 651 2675
rect 655 2671 656 2675
rect 650 2670 656 2671
rect 814 2659 820 2660
rect 814 2655 815 2659
rect 819 2655 820 2659
rect 814 2654 820 2655
rect 1138 2659 1144 2660
rect 1138 2655 1139 2659
rect 1143 2655 1144 2659
rect 1138 2654 1144 2655
rect 342 2643 348 2644
rect 342 2639 343 2643
rect 347 2639 348 2643
rect 342 2638 348 2639
rect 470 2643 476 2644
rect 470 2639 471 2643
rect 475 2639 476 2643
rect 470 2638 476 2639
rect 590 2643 596 2644
rect 590 2639 591 2643
rect 595 2639 596 2643
rect 590 2638 596 2639
rect 710 2643 716 2644
rect 710 2639 711 2643
rect 715 2639 716 2643
rect 710 2638 716 2639
rect 234 2631 240 2632
rect 234 2627 235 2631
rect 239 2627 240 2631
rect 234 2626 240 2627
rect 344 2623 346 2638
rect 472 2623 474 2638
rect 592 2623 594 2638
rect 712 2623 714 2638
rect 111 2622 115 2623
rect 111 2617 115 2618
rect 223 2622 227 2623
rect 223 2617 227 2618
rect 343 2622 347 2623
rect 343 2617 347 2618
rect 471 2622 475 2623
rect 471 2617 475 2618
rect 559 2622 563 2623
rect 559 2617 563 2618
rect 591 2622 595 2623
rect 591 2617 595 2618
rect 647 2622 651 2623
rect 647 2617 651 2618
rect 711 2622 715 2623
rect 711 2617 715 2618
rect 735 2622 739 2623
rect 735 2617 739 2618
rect 112 2593 114 2617
rect 472 2606 474 2617
rect 482 2615 488 2616
rect 482 2611 483 2615
rect 487 2611 488 2615
rect 482 2610 488 2611
rect 470 2605 476 2606
rect 470 2601 471 2605
rect 475 2601 476 2605
rect 470 2600 476 2601
rect 110 2592 116 2593
rect 110 2588 111 2592
rect 115 2588 116 2592
rect 110 2587 116 2588
rect 110 2575 116 2576
rect 110 2571 111 2575
rect 115 2571 116 2575
rect 110 2570 116 2571
rect 112 2547 114 2570
rect 462 2565 468 2566
rect 462 2561 463 2565
rect 467 2561 468 2565
rect 462 2560 468 2561
rect 464 2547 466 2560
rect 111 2546 115 2547
rect 111 2541 115 2542
rect 463 2546 467 2547
rect 463 2541 467 2542
rect 112 2526 114 2541
rect 484 2528 486 2610
rect 560 2606 562 2617
rect 648 2606 650 2617
rect 736 2606 738 2617
rect 816 2616 818 2654
rect 830 2643 836 2644
rect 830 2639 831 2643
rect 835 2639 836 2643
rect 830 2638 836 2639
rect 942 2643 948 2644
rect 942 2639 943 2643
rect 947 2639 948 2643
rect 942 2638 948 2639
rect 1054 2643 1060 2644
rect 1054 2639 1055 2643
rect 1059 2639 1060 2643
rect 1054 2638 1060 2639
rect 832 2623 834 2638
rect 843 2636 847 2637
rect 842 2631 848 2632
rect 842 2627 843 2631
rect 847 2627 848 2631
rect 842 2626 848 2627
rect 944 2623 946 2638
rect 1056 2623 1058 2638
rect 823 2622 827 2623
rect 823 2617 827 2618
rect 831 2622 835 2623
rect 831 2617 835 2618
rect 911 2622 915 2623
rect 911 2617 915 2618
rect 943 2622 947 2623
rect 943 2617 947 2618
rect 999 2622 1003 2623
rect 999 2617 1003 2618
rect 1055 2622 1059 2623
rect 1055 2617 1059 2618
rect 1087 2622 1091 2623
rect 1087 2617 1091 2618
rect 814 2615 820 2616
rect 814 2611 815 2615
rect 819 2611 820 2615
rect 814 2610 820 2611
rect 824 2606 826 2617
rect 912 2606 914 2617
rect 1000 2606 1002 2617
rect 1088 2606 1090 2617
rect 1140 2616 1142 2654
rect 1166 2643 1172 2644
rect 1166 2639 1167 2643
rect 1171 2639 1172 2643
rect 1166 2638 1172 2639
rect 1168 2623 1170 2638
rect 1180 2632 1182 2698
rect 1280 2695 1282 2704
rect 1416 2695 1418 2704
rect 1824 2695 1826 2714
rect 1863 2713 1867 2714
rect 1887 2718 1891 2719
rect 1887 2713 1891 2714
rect 1975 2718 1979 2719
rect 1975 2713 1979 2714
rect 2063 2718 2067 2719
rect 2063 2713 2067 2714
rect 2151 2718 2155 2719
rect 2151 2713 2155 2714
rect 2239 2718 2243 2719
rect 2239 2713 2243 2714
rect 2327 2718 2331 2719
rect 2327 2713 2331 2714
rect 2415 2718 2419 2719
rect 2415 2713 2419 2714
rect 2503 2718 2507 2719
rect 2503 2713 2507 2714
rect 2591 2718 2595 2719
rect 2591 2713 2595 2714
rect 2663 2718 2667 2719
rect 2663 2713 2667 2714
rect 2679 2718 2683 2719
rect 2679 2713 2683 2714
rect 2767 2718 2771 2719
rect 2767 2713 2771 2714
rect 2799 2718 2803 2719
rect 2799 2713 2803 2714
rect 2855 2718 2859 2719
rect 2855 2713 2859 2714
rect 2943 2718 2947 2719
rect 2943 2713 2947 2714
rect 2959 2718 2963 2719
rect 2959 2713 2963 2714
rect 3031 2718 3035 2719
rect 3031 2713 3035 2714
rect 3119 2718 3123 2719
rect 3119 2713 3123 2714
rect 3135 2718 3139 2719
rect 3135 2713 3139 2714
rect 3207 2718 3211 2719
rect 3207 2713 3211 2714
rect 3295 2718 3299 2719
rect 3295 2713 3299 2714
rect 3319 2718 3323 2719
rect 3319 2713 3323 2714
rect 1864 2698 1866 2713
rect 1888 2708 1890 2713
rect 1976 2708 1978 2713
rect 2064 2708 2066 2713
rect 2152 2708 2154 2713
rect 2240 2708 2242 2713
rect 2328 2708 2330 2713
rect 2416 2708 2418 2713
rect 2504 2708 2506 2713
rect 2592 2708 2594 2713
rect 2680 2708 2682 2713
rect 2768 2708 2770 2713
rect 2856 2708 2858 2713
rect 2944 2708 2946 2713
rect 3032 2708 3034 2713
rect 3120 2708 3122 2713
rect 3208 2708 3210 2713
rect 3296 2708 3298 2713
rect 1886 2707 1892 2708
rect 1886 2703 1887 2707
rect 1891 2703 1892 2707
rect 1886 2702 1892 2703
rect 1974 2707 1980 2708
rect 1974 2703 1975 2707
rect 1979 2703 1980 2707
rect 1974 2702 1980 2703
rect 2062 2707 2068 2708
rect 2062 2703 2063 2707
rect 2067 2703 2068 2707
rect 2062 2702 2068 2703
rect 2150 2707 2156 2708
rect 2150 2703 2151 2707
rect 2155 2703 2156 2707
rect 2150 2702 2156 2703
rect 2238 2707 2244 2708
rect 2238 2703 2239 2707
rect 2243 2703 2244 2707
rect 2238 2702 2244 2703
rect 2326 2707 2332 2708
rect 2326 2703 2327 2707
rect 2331 2703 2332 2707
rect 2326 2702 2332 2703
rect 2414 2707 2420 2708
rect 2414 2703 2415 2707
rect 2419 2703 2420 2707
rect 2414 2702 2420 2703
rect 2502 2707 2508 2708
rect 2502 2703 2503 2707
rect 2507 2703 2508 2707
rect 2502 2702 2508 2703
rect 2590 2707 2596 2708
rect 2590 2703 2591 2707
rect 2595 2703 2596 2707
rect 2590 2702 2596 2703
rect 2678 2707 2684 2708
rect 2678 2703 2679 2707
rect 2683 2703 2684 2707
rect 2678 2702 2684 2703
rect 2766 2707 2772 2708
rect 2766 2703 2767 2707
rect 2771 2703 2772 2707
rect 2766 2702 2772 2703
rect 2854 2707 2860 2708
rect 2854 2703 2855 2707
rect 2859 2703 2860 2707
rect 2854 2702 2860 2703
rect 2942 2707 2948 2708
rect 2942 2703 2943 2707
rect 2947 2703 2948 2707
rect 2942 2702 2948 2703
rect 3030 2707 3036 2708
rect 3030 2703 3031 2707
rect 3035 2703 3036 2707
rect 3030 2702 3036 2703
rect 3118 2707 3124 2708
rect 3118 2703 3119 2707
rect 3123 2703 3124 2707
rect 3118 2702 3124 2703
rect 3206 2707 3212 2708
rect 3206 2703 3207 2707
rect 3211 2703 3212 2707
rect 3206 2702 3212 2703
rect 3294 2707 3300 2708
rect 3294 2703 3295 2707
rect 3299 2703 3300 2707
rect 3294 2702 3300 2703
rect 3364 2700 3366 2727
rect 3478 2725 3479 2729
rect 3483 2725 3484 2729
rect 3478 2724 3484 2725
rect 3480 2719 3482 2724
rect 3498 2723 3504 2724
rect 3498 2719 3499 2723
rect 3503 2719 3504 2723
rect 3576 2719 3578 2734
rect 3391 2718 3395 2719
rect 3391 2713 3395 2714
rect 3479 2718 3483 2719
rect 3498 2718 3504 2719
rect 3575 2718 3579 2719
rect 3479 2713 3483 2714
rect 3392 2708 3394 2713
rect 3480 2708 3482 2713
rect 3390 2707 3396 2708
rect 3390 2703 3391 2707
rect 3395 2703 3396 2707
rect 3390 2702 3396 2703
rect 3478 2707 3484 2708
rect 3478 2703 3479 2707
rect 3483 2703 3484 2707
rect 3478 2702 3484 2703
rect 3362 2699 3368 2700
rect 1862 2697 1868 2698
rect 1271 2694 1275 2695
rect 1271 2689 1275 2690
rect 1279 2694 1283 2695
rect 1279 2689 1283 2690
rect 1415 2694 1419 2695
rect 1415 2689 1419 2690
rect 1823 2694 1827 2695
rect 1862 2693 1863 2697
rect 1867 2693 1868 2697
rect 3362 2695 3363 2699
rect 3367 2695 3368 2699
rect 3362 2694 3368 2695
rect 1862 2692 1868 2693
rect 1823 2689 1827 2690
rect 1272 2684 1274 2689
rect 1270 2683 1276 2684
rect 1270 2679 1271 2683
rect 1275 2679 1276 2683
rect 1270 2678 1276 2679
rect 1226 2675 1232 2676
rect 1226 2671 1227 2675
rect 1231 2671 1232 2675
rect 1824 2674 1826 2689
rect 2042 2683 2048 2684
rect 1862 2680 1868 2681
rect 1862 2676 1863 2680
rect 1867 2676 1868 2680
rect 2042 2679 2043 2683
rect 2047 2679 2048 2683
rect 2042 2678 2048 2679
rect 3470 2683 3476 2684
rect 3470 2679 3471 2683
rect 3475 2679 3476 2683
rect 3470 2678 3476 2679
rect 1862 2675 1868 2676
rect 1226 2670 1232 2671
rect 1822 2673 1828 2674
rect 1228 2637 1230 2670
rect 1822 2669 1823 2673
rect 1827 2669 1828 2673
rect 1822 2668 1828 2669
rect 1822 2656 1828 2657
rect 1822 2652 1823 2656
rect 1827 2652 1828 2656
rect 1822 2651 1828 2652
rect 1278 2643 1284 2644
rect 1278 2639 1279 2643
rect 1283 2639 1284 2643
rect 1278 2638 1284 2639
rect 1227 2636 1231 2637
rect 1178 2631 1184 2632
rect 1227 2631 1231 2632
rect 1178 2627 1179 2631
rect 1183 2627 1184 2631
rect 1178 2626 1184 2627
rect 1280 2623 1282 2638
rect 1824 2623 1826 2651
rect 1864 2631 1866 2675
rect 1894 2667 1900 2668
rect 1894 2663 1895 2667
rect 1899 2663 1900 2667
rect 1894 2662 1900 2663
rect 1982 2667 1988 2668
rect 1982 2663 1983 2667
rect 1987 2663 1988 2667
rect 1982 2662 1988 2663
rect 1896 2631 1898 2662
rect 1950 2655 1956 2656
rect 1950 2651 1951 2655
rect 1955 2651 1956 2655
rect 1950 2650 1956 2651
rect 1863 2630 1867 2631
rect 1863 2625 1867 2626
rect 1895 2630 1899 2631
rect 1895 2625 1899 2626
rect 1167 2622 1171 2623
rect 1167 2617 1171 2618
rect 1175 2622 1179 2623
rect 1175 2617 1179 2618
rect 1263 2622 1267 2623
rect 1263 2617 1267 2618
rect 1279 2622 1283 2623
rect 1279 2617 1283 2618
rect 1823 2622 1827 2623
rect 1823 2617 1827 2618
rect 1138 2615 1144 2616
rect 1138 2611 1139 2615
rect 1143 2611 1144 2615
rect 1138 2610 1144 2611
rect 1176 2606 1178 2617
rect 1264 2606 1266 2617
rect 558 2605 564 2606
rect 558 2601 559 2605
rect 563 2601 564 2605
rect 558 2600 564 2601
rect 646 2605 652 2606
rect 646 2601 647 2605
rect 651 2601 652 2605
rect 646 2600 652 2601
rect 734 2605 740 2606
rect 734 2601 735 2605
rect 739 2601 740 2605
rect 734 2600 740 2601
rect 822 2605 828 2606
rect 822 2601 823 2605
rect 827 2601 828 2605
rect 822 2600 828 2601
rect 910 2605 916 2606
rect 910 2601 911 2605
rect 915 2601 916 2605
rect 910 2600 916 2601
rect 998 2605 1004 2606
rect 998 2601 999 2605
rect 1003 2601 1004 2605
rect 998 2600 1004 2601
rect 1086 2605 1092 2606
rect 1086 2601 1087 2605
rect 1091 2601 1092 2605
rect 1086 2600 1092 2601
rect 1174 2605 1180 2606
rect 1174 2601 1175 2605
rect 1179 2601 1180 2605
rect 1174 2600 1180 2601
rect 1262 2605 1268 2606
rect 1262 2601 1263 2605
rect 1267 2601 1268 2605
rect 1262 2600 1268 2601
rect 1824 2593 1826 2617
rect 1864 2601 1866 2625
rect 1862 2600 1868 2601
rect 1862 2596 1863 2600
rect 1867 2596 1868 2600
rect 1952 2597 1954 2650
rect 1984 2631 1986 2662
rect 2044 2656 2046 2678
rect 2070 2667 2076 2668
rect 2070 2663 2071 2667
rect 2075 2663 2076 2667
rect 2070 2662 2076 2663
rect 2158 2667 2164 2668
rect 2158 2663 2159 2667
rect 2163 2663 2164 2667
rect 2158 2662 2164 2663
rect 2246 2667 2252 2668
rect 2246 2663 2247 2667
rect 2251 2663 2252 2667
rect 2246 2662 2252 2663
rect 2334 2667 2340 2668
rect 2334 2663 2335 2667
rect 2339 2663 2340 2667
rect 2334 2662 2340 2663
rect 2422 2667 2428 2668
rect 2422 2663 2423 2667
rect 2427 2663 2428 2667
rect 2422 2662 2428 2663
rect 2510 2667 2516 2668
rect 2510 2663 2511 2667
rect 2515 2663 2516 2667
rect 2510 2662 2516 2663
rect 2598 2667 2604 2668
rect 2598 2663 2599 2667
rect 2603 2663 2604 2667
rect 2598 2662 2604 2663
rect 2686 2667 2692 2668
rect 2686 2663 2687 2667
rect 2691 2663 2692 2667
rect 2686 2662 2692 2663
rect 2774 2667 2780 2668
rect 2774 2663 2775 2667
rect 2779 2663 2780 2667
rect 2774 2662 2780 2663
rect 2862 2667 2868 2668
rect 2862 2663 2863 2667
rect 2867 2663 2868 2667
rect 2862 2662 2868 2663
rect 2950 2667 2956 2668
rect 2950 2663 2951 2667
rect 2955 2663 2956 2667
rect 2950 2662 2956 2663
rect 3038 2667 3044 2668
rect 3038 2663 3039 2667
rect 3043 2663 3044 2667
rect 3038 2662 3044 2663
rect 3126 2667 3132 2668
rect 3126 2663 3127 2667
rect 3131 2663 3132 2667
rect 3126 2662 3132 2663
rect 3214 2667 3220 2668
rect 3214 2663 3215 2667
rect 3219 2663 3220 2667
rect 3214 2662 3220 2663
rect 3302 2667 3308 2668
rect 3302 2663 3303 2667
rect 3307 2663 3308 2667
rect 3302 2662 3308 2663
rect 3398 2667 3404 2668
rect 3398 2663 3399 2667
rect 3403 2663 3404 2667
rect 3398 2662 3404 2663
rect 2042 2655 2048 2656
rect 2042 2651 2043 2655
rect 2047 2651 2048 2655
rect 2042 2650 2048 2651
rect 2072 2631 2074 2662
rect 2160 2631 2162 2662
rect 2248 2631 2250 2662
rect 2336 2631 2338 2662
rect 2424 2631 2426 2662
rect 2498 2631 2504 2632
rect 2512 2631 2514 2662
rect 2600 2631 2602 2662
rect 2688 2631 2690 2662
rect 2776 2631 2778 2662
rect 2864 2631 2866 2662
rect 2952 2631 2954 2662
rect 3040 2631 3042 2662
rect 3078 2631 3084 2632
rect 3128 2631 3130 2662
rect 3216 2631 3218 2662
rect 3304 2631 3306 2662
rect 3400 2631 3402 2662
rect 1983 2630 1987 2631
rect 1983 2625 1987 2626
rect 2071 2630 2075 2631
rect 2071 2625 2075 2626
rect 2159 2630 2163 2631
rect 2159 2625 2163 2626
rect 2247 2630 2251 2631
rect 2247 2625 2251 2626
rect 2279 2630 2283 2631
rect 2279 2625 2283 2626
rect 2335 2630 2339 2631
rect 2335 2625 2339 2626
rect 2415 2630 2419 2631
rect 2415 2625 2419 2626
rect 2423 2630 2427 2631
rect 2498 2627 2499 2631
rect 2503 2627 2504 2631
rect 2498 2626 2504 2627
rect 2511 2630 2515 2631
rect 2423 2625 2427 2626
rect 2160 2614 2162 2625
rect 2280 2614 2282 2625
rect 2416 2614 2418 2625
rect 2158 2613 2164 2614
rect 2158 2609 2159 2613
rect 2163 2609 2164 2613
rect 2158 2608 2164 2609
rect 2278 2613 2284 2614
rect 2278 2609 2279 2613
rect 2283 2609 2284 2613
rect 2278 2608 2284 2609
rect 2414 2613 2420 2614
rect 2414 2609 2415 2613
rect 2419 2609 2420 2613
rect 2414 2608 2420 2609
rect 1862 2595 1868 2596
rect 1951 2596 1955 2597
rect 1822 2592 1828 2593
rect 1822 2588 1823 2592
rect 1827 2588 1828 2592
rect 1951 2591 1955 2592
rect 1822 2587 1828 2588
rect 1862 2583 1868 2584
rect 1862 2579 1863 2583
rect 1867 2579 1868 2583
rect 1862 2578 1868 2579
rect 714 2575 720 2576
rect 714 2571 715 2575
rect 719 2571 720 2575
rect 714 2570 720 2571
rect 1822 2575 1828 2576
rect 1822 2571 1823 2575
rect 1827 2571 1828 2575
rect 1822 2570 1828 2571
rect 550 2565 556 2566
rect 550 2561 551 2565
rect 555 2561 556 2565
rect 550 2560 556 2561
rect 638 2565 644 2566
rect 638 2561 639 2565
rect 643 2561 644 2565
rect 638 2560 644 2561
rect 552 2547 554 2560
rect 640 2547 642 2560
rect 495 2546 499 2547
rect 495 2541 499 2542
rect 551 2546 555 2547
rect 551 2541 555 2542
rect 583 2546 587 2547
rect 583 2541 587 2542
rect 639 2546 643 2547
rect 639 2541 643 2542
rect 671 2546 675 2547
rect 671 2541 675 2542
rect 496 2536 498 2541
rect 584 2536 586 2541
rect 672 2536 674 2541
rect 494 2535 500 2536
rect 494 2531 495 2535
rect 499 2531 500 2535
rect 494 2530 500 2531
rect 582 2535 588 2536
rect 582 2531 583 2535
rect 587 2531 588 2535
rect 582 2530 588 2531
rect 670 2535 676 2536
rect 670 2531 671 2535
rect 675 2531 676 2535
rect 670 2530 676 2531
rect 482 2527 488 2528
rect 110 2525 116 2526
rect 110 2521 111 2525
rect 115 2521 116 2525
rect 482 2523 483 2527
rect 487 2523 488 2527
rect 482 2522 488 2523
rect 110 2520 116 2521
rect 562 2511 568 2512
rect 110 2508 116 2509
rect 110 2504 111 2508
rect 115 2504 116 2508
rect 562 2507 563 2511
rect 567 2507 568 2511
rect 562 2506 568 2507
rect 110 2503 116 2504
rect 112 2475 114 2503
rect 502 2495 508 2496
rect 502 2491 503 2495
rect 507 2491 508 2495
rect 502 2490 508 2491
rect 504 2475 506 2490
rect 564 2484 566 2506
rect 590 2495 596 2496
rect 590 2491 591 2495
rect 595 2491 596 2495
rect 590 2490 596 2491
rect 678 2495 684 2496
rect 678 2491 679 2495
rect 683 2491 684 2495
rect 678 2490 684 2491
rect 562 2483 568 2484
rect 562 2479 563 2483
rect 567 2479 568 2483
rect 562 2478 568 2479
rect 582 2483 588 2484
rect 582 2479 583 2483
rect 587 2479 588 2483
rect 582 2478 588 2479
rect 111 2474 115 2475
rect 111 2469 115 2470
rect 359 2474 363 2475
rect 359 2469 363 2470
rect 471 2474 475 2475
rect 471 2469 475 2470
rect 503 2474 507 2475
rect 503 2469 507 2470
rect 112 2445 114 2469
rect 360 2458 362 2469
rect 414 2463 420 2464
rect 414 2458 415 2463
rect 358 2457 364 2458
rect 358 2453 359 2457
rect 363 2453 364 2457
rect 419 2458 420 2463
rect 472 2458 474 2469
rect 415 2455 419 2456
rect 470 2457 476 2458
rect 358 2452 364 2453
rect 470 2453 471 2457
rect 475 2453 476 2457
rect 470 2452 476 2453
rect 110 2444 116 2445
rect 110 2440 111 2444
rect 115 2440 116 2444
rect 584 2440 586 2478
rect 592 2475 594 2490
rect 680 2475 682 2490
rect 716 2484 718 2570
rect 726 2565 732 2566
rect 726 2561 727 2565
rect 731 2561 732 2565
rect 726 2560 732 2561
rect 814 2565 820 2566
rect 814 2561 815 2565
rect 819 2561 820 2565
rect 814 2560 820 2561
rect 902 2565 908 2566
rect 902 2561 903 2565
rect 907 2561 908 2565
rect 902 2560 908 2561
rect 990 2565 996 2566
rect 990 2561 991 2565
rect 995 2561 996 2565
rect 990 2560 996 2561
rect 1078 2565 1084 2566
rect 1078 2561 1079 2565
rect 1083 2561 1084 2565
rect 1078 2560 1084 2561
rect 1166 2565 1172 2566
rect 1166 2561 1167 2565
rect 1171 2561 1172 2565
rect 1166 2560 1172 2561
rect 1254 2565 1260 2566
rect 1254 2561 1255 2565
rect 1259 2561 1260 2565
rect 1254 2560 1260 2561
rect 728 2547 730 2560
rect 816 2547 818 2560
rect 904 2547 906 2560
rect 954 2559 960 2560
rect 954 2555 955 2559
rect 959 2555 960 2559
rect 954 2554 960 2555
rect 727 2546 731 2547
rect 727 2541 731 2542
rect 759 2546 763 2547
rect 759 2541 763 2542
rect 815 2546 819 2547
rect 815 2541 819 2542
rect 847 2546 851 2547
rect 847 2541 851 2542
rect 903 2546 907 2547
rect 903 2541 907 2542
rect 935 2546 939 2547
rect 935 2541 939 2542
rect 760 2536 762 2541
rect 848 2536 850 2541
rect 936 2536 938 2541
rect 758 2535 764 2536
rect 758 2531 759 2535
rect 763 2531 764 2535
rect 758 2530 764 2531
rect 846 2535 852 2536
rect 846 2531 847 2535
rect 851 2531 852 2535
rect 846 2530 852 2531
rect 934 2535 940 2536
rect 934 2531 935 2535
rect 939 2531 940 2535
rect 934 2530 940 2531
rect 838 2527 844 2528
rect 838 2523 839 2527
rect 843 2523 844 2527
rect 838 2522 844 2523
rect 766 2495 772 2496
rect 766 2491 767 2495
rect 771 2491 772 2495
rect 766 2490 772 2491
rect 714 2483 720 2484
rect 714 2479 715 2483
rect 719 2479 720 2483
rect 714 2478 720 2479
rect 768 2475 770 2490
rect 591 2474 595 2475
rect 591 2469 595 2470
rect 679 2474 683 2475
rect 679 2469 683 2470
rect 719 2474 723 2475
rect 719 2469 723 2470
rect 767 2474 771 2475
rect 767 2469 771 2470
rect 592 2458 594 2469
rect 720 2458 722 2469
rect 840 2468 842 2522
rect 854 2495 860 2496
rect 854 2491 855 2495
rect 859 2491 860 2495
rect 854 2490 860 2491
rect 942 2495 948 2496
rect 942 2491 943 2495
rect 947 2491 948 2495
rect 942 2490 948 2491
rect 856 2475 858 2490
rect 944 2475 946 2490
rect 956 2484 958 2554
rect 992 2547 994 2560
rect 1080 2547 1082 2560
rect 1168 2547 1170 2560
rect 1256 2547 1258 2560
rect 1824 2547 1826 2570
rect 1864 2563 1866 2578
rect 2150 2573 2156 2574
rect 2150 2569 2151 2573
rect 2155 2569 2156 2573
rect 2150 2568 2156 2569
rect 2270 2573 2276 2574
rect 2270 2569 2271 2573
rect 2275 2569 2276 2573
rect 2270 2568 2276 2569
rect 2406 2573 2412 2574
rect 2406 2569 2407 2573
rect 2411 2569 2412 2573
rect 2406 2568 2412 2569
rect 2152 2563 2154 2568
rect 2272 2563 2274 2568
rect 2408 2563 2410 2568
rect 1863 2562 1867 2563
rect 1863 2557 1867 2558
rect 2103 2562 2107 2563
rect 2103 2557 2107 2558
rect 2151 2562 2155 2563
rect 2151 2557 2155 2558
rect 2199 2562 2203 2563
rect 2199 2557 2203 2558
rect 2271 2562 2275 2563
rect 2271 2557 2275 2558
rect 2311 2562 2315 2563
rect 2311 2557 2315 2558
rect 2407 2562 2411 2563
rect 2407 2557 2411 2558
rect 2431 2562 2435 2563
rect 2431 2557 2435 2558
rect 991 2546 995 2547
rect 991 2541 995 2542
rect 1023 2546 1027 2547
rect 1023 2541 1027 2542
rect 1079 2546 1083 2547
rect 1079 2541 1083 2542
rect 1111 2546 1115 2547
rect 1111 2541 1115 2542
rect 1167 2546 1171 2547
rect 1167 2541 1171 2542
rect 1199 2546 1203 2547
rect 1199 2541 1203 2542
rect 1255 2546 1259 2547
rect 1255 2541 1259 2542
rect 1287 2546 1291 2547
rect 1287 2541 1291 2542
rect 1823 2546 1827 2547
rect 1864 2542 1866 2557
rect 2104 2552 2106 2557
rect 2200 2552 2202 2557
rect 2312 2552 2314 2557
rect 2432 2552 2434 2557
rect 2102 2551 2108 2552
rect 2102 2547 2103 2551
rect 2107 2547 2108 2551
rect 2102 2546 2108 2547
rect 2198 2551 2204 2552
rect 2198 2547 2199 2551
rect 2203 2547 2204 2551
rect 2198 2546 2204 2547
rect 2310 2551 2316 2552
rect 2310 2547 2311 2551
rect 2315 2547 2316 2551
rect 2310 2546 2316 2547
rect 2430 2551 2436 2552
rect 2430 2547 2431 2551
rect 2435 2547 2436 2551
rect 2430 2546 2436 2547
rect 2500 2544 2502 2626
rect 2511 2625 2515 2626
rect 2551 2630 2555 2631
rect 2551 2625 2555 2626
rect 2599 2630 2603 2631
rect 2599 2625 2603 2626
rect 2687 2630 2691 2631
rect 2687 2625 2691 2626
rect 2695 2630 2699 2631
rect 2695 2625 2699 2626
rect 2775 2630 2779 2631
rect 2775 2625 2779 2626
rect 2847 2630 2851 2631
rect 2847 2625 2851 2626
rect 2863 2630 2867 2631
rect 2863 2625 2867 2626
rect 2951 2630 2955 2631
rect 2951 2625 2955 2626
rect 2999 2630 3003 2631
rect 2999 2625 3003 2626
rect 3039 2630 3043 2631
rect 3078 2627 3079 2631
rect 3083 2627 3084 2631
rect 3078 2626 3084 2627
rect 3127 2630 3131 2631
rect 3039 2625 3043 2626
rect 2552 2614 2554 2625
rect 2696 2614 2698 2625
rect 2848 2614 2850 2625
rect 3000 2614 3002 2625
rect 2550 2613 2556 2614
rect 2550 2609 2551 2613
rect 2555 2609 2556 2613
rect 2550 2608 2556 2609
rect 2694 2613 2700 2614
rect 2694 2609 2695 2613
rect 2699 2609 2700 2613
rect 2694 2608 2700 2609
rect 2846 2613 2852 2614
rect 2846 2609 2847 2613
rect 2851 2609 2852 2613
rect 2846 2608 2852 2609
rect 2998 2613 3004 2614
rect 2998 2609 2999 2613
rect 3003 2609 3004 2613
rect 2998 2608 3004 2609
rect 2643 2596 2647 2597
rect 3080 2596 3082 2626
rect 3127 2625 3131 2626
rect 3159 2630 3163 2631
rect 3159 2625 3163 2626
rect 3215 2630 3219 2631
rect 3215 2625 3219 2626
rect 3303 2630 3307 2631
rect 3303 2625 3307 2626
rect 3399 2630 3403 2631
rect 3399 2625 3403 2626
rect 3160 2614 3162 2625
rect 3166 2623 3172 2624
rect 3166 2619 3167 2623
rect 3171 2619 3172 2623
rect 3166 2618 3172 2619
rect 3158 2613 3164 2614
rect 3158 2609 3159 2613
rect 3163 2609 3164 2613
rect 3158 2608 3164 2609
rect 2642 2591 2643 2596
rect 2647 2591 2648 2596
rect 2642 2590 2648 2591
rect 3078 2595 3084 2596
rect 3078 2591 3079 2595
rect 3083 2591 3084 2595
rect 3078 2590 3084 2591
rect 2542 2573 2548 2574
rect 2542 2569 2543 2573
rect 2547 2569 2548 2573
rect 2542 2568 2548 2569
rect 2686 2573 2692 2574
rect 2686 2569 2687 2573
rect 2691 2569 2692 2573
rect 2686 2568 2692 2569
rect 2838 2573 2844 2574
rect 2838 2569 2839 2573
rect 2843 2569 2844 2573
rect 2838 2568 2844 2569
rect 2990 2573 2996 2574
rect 2990 2569 2991 2573
rect 2995 2569 2996 2573
rect 2990 2568 2996 2569
rect 3150 2573 3156 2574
rect 3150 2569 3151 2573
rect 3155 2569 3156 2573
rect 3150 2568 3156 2569
rect 2544 2563 2546 2568
rect 2688 2563 2690 2568
rect 2840 2563 2842 2568
rect 2992 2563 2994 2568
rect 3018 2567 3024 2568
rect 3018 2563 3019 2567
rect 3023 2563 3024 2567
rect 3152 2563 3154 2568
rect 2543 2562 2547 2563
rect 2543 2557 2547 2558
rect 2559 2562 2563 2563
rect 2559 2557 2563 2558
rect 2687 2562 2691 2563
rect 2687 2557 2691 2558
rect 2695 2562 2699 2563
rect 2695 2557 2699 2558
rect 2839 2562 2843 2563
rect 2839 2557 2843 2558
rect 2847 2562 2851 2563
rect 2847 2557 2851 2558
rect 2991 2562 2995 2563
rect 2991 2557 2995 2558
rect 2999 2562 3003 2563
rect 3018 2562 3024 2563
rect 3151 2562 3155 2563
rect 2999 2557 3003 2558
rect 2560 2552 2562 2557
rect 2696 2552 2698 2557
rect 2848 2552 2850 2557
rect 3000 2552 3002 2557
rect 2558 2551 2564 2552
rect 2558 2547 2559 2551
rect 2563 2547 2564 2551
rect 2558 2546 2564 2547
rect 2694 2551 2700 2552
rect 2694 2547 2695 2551
rect 2699 2547 2700 2551
rect 2694 2546 2700 2547
rect 2846 2551 2852 2552
rect 2846 2547 2847 2551
rect 2851 2547 2852 2551
rect 2846 2546 2852 2547
rect 2998 2551 3004 2552
rect 2998 2547 2999 2551
rect 3003 2547 3004 2551
rect 2998 2546 3004 2547
rect 2498 2543 2504 2544
rect 1823 2541 1827 2542
rect 1862 2541 1868 2542
rect 1024 2536 1026 2541
rect 1112 2536 1114 2541
rect 1200 2536 1202 2541
rect 1288 2536 1290 2541
rect 1022 2535 1028 2536
rect 1022 2531 1023 2535
rect 1027 2531 1028 2535
rect 1022 2530 1028 2531
rect 1110 2535 1116 2536
rect 1110 2531 1111 2535
rect 1115 2531 1116 2535
rect 1110 2530 1116 2531
rect 1198 2535 1204 2536
rect 1198 2531 1199 2535
rect 1203 2531 1204 2535
rect 1198 2530 1204 2531
rect 1286 2535 1292 2536
rect 1286 2531 1287 2535
rect 1291 2531 1292 2535
rect 1286 2530 1292 2531
rect 1266 2527 1272 2528
rect 1266 2523 1267 2527
rect 1271 2523 1272 2527
rect 1824 2526 1826 2541
rect 1862 2537 1863 2541
rect 1867 2537 1868 2541
rect 2498 2539 2499 2543
rect 2503 2539 2504 2543
rect 2498 2538 2504 2539
rect 1862 2536 1868 2537
rect 2626 2527 2632 2528
rect 1266 2522 1272 2523
rect 1822 2525 1828 2526
rect 1030 2495 1036 2496
rect 979 2492 983 2493
rect 1030 2491 1031 2495
rect 1035 2491 1036 2495
rect 1030 2490 1036 2491
rect 1118 2495 1124 2496
rect 1118 2491 1119 2495
rect 1123 2491 1124 2495
rect 1118 2490 1124 2491
rect 1206 2495 1212 2496
rect 1206 2491 1207 2495
rect 1211 2491 1212 2495
rect 1268 2493 1270 2522
rect 1822 2521 1823 2525
rect 1827 2521 1828 2525
rect 1822 2520 1828 2521
rect 1862 2524 1868 2525
rect 1862 2520 1863 2524
rect 1867 2520 1868 2524
rect 2626 2523 2627 2527
rect 2631 2523 2632 2527
rect 2626 2522 2632 2523
rect 2762 2527 2768 2528
rect 2762 2523 2763 2527
rect 2767 2523 2768 2527
rect 2762 2522 2768 2523
rect 2914 2527 2920 2528
rect 2914 2523 2915 2527
rect 2919 2523 2920 2527
rect 2914 2522 2920 2523
rect 1862 2519 1868 2520
rect 1822 2508 1828 2509
rect 1822 2504 1823 2508
rect 1827 2504 1828 2508
rect 1822 2503 1828 2504
rect 1294 2495 1300 2496
rect 1206 2490 1212 2491
rect 1267 2492 1271 2493
rect 979 2487 983 2488
rect 954 2483 960 2484
rect 954 2479 955 2483
rect 959 2479 960 2483
rect 954 2478 960 2479
rect 847 2474 851 2475
rect 847 2469 851 2470
rect 855 2474 859 2475
rect 855 2469 859 2470
rect 943 2474 947 2475
rect 943 2469 947 2470
rect 967 2474 971 2475
rect 967 2469 971 2470
rect 730 2467 736 2468
rect 730 2463 731 2467
rect 735 2463 736 2467
rect 730 2462 736 2463
rect 838 2467 844 2468
rect 838 2463 839 2467
rect 843 2463 844 2467
rect 838 2462 844 2463
rect 590 2457 596 2458
rect 590 2453 591 2457
rect 595 2453 596 2457
rect 590 2452 596 2453
rect 718 2457 724 2458
rect 718 2453 719 2457
rect 723 2453 724 2457
rect 718 2452 724 2453
rect 110 2439 116 2440
rect 582 2439 588 2440
rect 582 2435 583 2439
rect 587 2435 588 2439
rect 582 2434 588 2435
rect 110 2427 116 2428
rect 110 2423 111 2427
rect 115 2423 116 2427
rect 110 2422 116 2423
rect 112 2403 114 2422
rect 350 2417 356 2418
rect 350 2413 351 2417
rect 355 2413 356 2417
rect 350 2412 356 2413
rect 462 2417 468 2418
rect 462 2413 463 2417
rect 467 2413 468 2417
rect 462 2412 468 2413
rect 582 2417 588 2418
rect 582 2413 583 2417
rect 587 2413 588 2417
rect 582 2412 588 2413
rect 710 2417 716 2418
rect 710 2413 711 2417
rect 715 2413 716 2417
rect 710 2412 716 2413
rect 352 2403 354 2412
rect 464 2403 466 2412
rect 490 2411 496 2412
rect 490 2407 491 2411
rect 495 2407 496 2411
rect 490 2406 496 2407
rect 111 2402 115 2403
rect 111 2397 115 2398
rect 135 2402 139 2403
rect 135 2397 139 2398
rect 287 2402 291 2403
rect 287 2397 291 2398
rect 351 2402 355 2403
rect 351 2397 355 2398
rect 463 2402 467 2403
rect 463 2397 467 2398
rect 471 2402 475 2403
rect 471 2397 475 2398
rect 112 2382 114 2397
rect 136 2392 138 2397
rect 288 2392 290 2397
rect 472 2392 474 2397
rect 134 2391 140 2392
rect 134 2387 135 2391
rect 139 2387 140 2391
rect 134 2386 140 2387
rect 286 2391 292 2392
rect 286 2387 287 2391
rect 291 2387 292 2391
rect 286 2386 292 2387
rect 470 2391 476 2392
rect 470 2387 471 2391
rect 475 2387 476 2391
rect 470 2386 476 2387
rect 202 2383 208 2384
rect 110 2381 116 2382
rect 110 2377 111 2381
rect 115 2377 116 2381
rect 202 2379 203 2383
rect 207 2379 208 2383
rect 202 2378 208 2379
rect 110 2376 116 2377
rect 110 2364 116 2365
rect 110 2360 111 2364
rect 115 2360 116 2364
rect 110 2359 116 2360
rect 112 2331 114 2359
rect 142 2351 148 2352
rect 142 2347 143 2351
rect 147 2347 148 2351
rect 142 2346 148 2347
rect 144 2331 146 2346
rect 204 2340 206 2378
rect 362 2367 368 2368
rect 362 2363 363 2367
rect 367 2363 368 2367
rect 362 2362 368 2363
rect 294 2351 300 2352
rect 294 2347 295 2351
rect 299 2347 300 2351
rect 294 2346 300 2347
rect 202 2339 208 2340
rect 202 2335 203 2339
rect 207 2335 208 2339
rect 202 2334 208 2335
rect 296 2331 298 2346
rect 364 2340 366 2362
rect 478 2351 484 2352
rect 478 2347 479 2351
rect 483 2347 484 2351
rect 478 2346 484 2347
rect 362 2339 368 2340
rect 362 2335 363 2339
rect 367 2335 368 2339
rect 362 2334 368 2335
rect 480 2331 482 2346
rect 492 2340 494 2406
rect 584 2403 586 2412
rect 712 2403 714 2412
rect 583 2402 587 2403
rect 583 2397 587 2398
rect 663 2402 667 2403
rect 663 2397 667 2398
rect 711 2402 715 2403
rect 711 2397 715 2398
rect 664 2392 666 2397
rect 662 2391 668 2392
rect 662 2387 663 2391
rect 667 2387 668 2391
rect 662 2386 668 2387
rect 732 2384 734 2462
rect 787 2460 791 2461
rect 848 2458 850 2469
rect 968 2458 970 2469
rect 980 2468 982 2487
rect 1032 2475 1034 2490
rect 1120 2475 1122 2490
rect 1208 2475 1210 2490
rect 1294 2491 1295 2495
rect 1299 2491 1300 2495
rect 1294 2490 1300 2491
rect 1267 2487 1271 2488
rect 1296 2475 1298 2490
rect 1824 2475 1826 2503
rect 1864 2491 1866 2519
rect 2110 2511 2116 2512
rect 2110 2507 2111 2511
rect 2115 2507 2116 2511
rect 2110 2506 2116 2507
rect 2206 2511 2212 2512
rect 2206 2507 2207 2511
rect 2211 2507 2212 2511
rect 2206 2506 2212 2507
rect 2318 2511 2324 2512
rect 2318 2507 2319 2511
rect 2323 2507 2324 2511
rect 2318 2506 2324 2507
rect 2438 2511 2444 2512
rect 2438 2507 2439 2511
rect 2443 2507 2444 2511
rect 2438 2506 2444 2507
rect 2566 2511 2572 2512
rect 2566 2507 2567 2511
rect 2571 2507 2572 2511
rect 2566 2506 2572 2507
rect 2112 2491 2114 2506
rect 2208 2491 2210 2506
rect 2320 2491 2322 2506
rect 2440 2491 2442 2506
rect 2568 2491 2570 2506
rect 1863 2490 1867 2491
rect 1863 2485 1867 2486
rect 2087 2490 2091 2491
rect 2087 2485 2091 2486
rect 2111 2490 2115 2491
rect 2111 2485 2115 2486
rect 2183 2490 2187 2491
rect 2183 2485 2187 2486
rect 2207 2490 2211 2491
rect 2207 2485 2211 2486
rect 2287 2490 2291 2491
rect 2287 2485 2291 2486
rect 2319 2490 2323 2491
rect 2319 2485 2323 2486
rect 2407 2490 2411 2491
rect 2407 2485 2411 2486
rect 2439 2490 2443 2491
rect 2439 2485 2443 2486
rect 2543 2490 2547 2491
rect 2543 2485 2547 2486
rect 2567 2490 2571 2491
rect 2567 2485 2571 2486
rect 1031 2474 1035 2475
rect 1031 2469 1035 2470
rect 1087 2474 1091 2475
rect 1087 2469 1091 2470
rect 1119 2474 1123 2475
rect 1119 2469 1123 2470
rect 1207 2474 1211 2475
rect 1207 2469 1211 2470
rect 1295 2474 1299 2475
rect 1295 2469 1299 2470
rect 1335 2474 1339 2475
rect 1335 2469 1339 2470
rect 1463 2474 1467 2475
rect 1463 2469 1467 2470
rect 1823 2474 1827 2475
rect 1823 2469 1827 2470
rect 978 2467 984 2468
rect 978 2463 979 2467
rect 983 2463 984 2467
rect 978 2462 984 2463
rect 1088 2458 1090 2469
rect 1146 2467 1152 2468
rect 1146 2463 1147 2467
rect 1151 2463 1152 2467
rect 1146 2462 1152 2463
rect 787 2455 791 2456
rect 846 2457 852 2458
rect 788 2440 790 2455
rect 846 2453 847 2457
rect 851 2453 852 2457
rect 846 2452 852 2453
rect 966 2457 972 2458
rect 966 2453 967 2457
rect 971 2453 972 2457
rect 966 2452 972 2453
rect 1086 2457 1092 2458
rect 1086 2453 1087 2457
rect 1091 2453 1092 2457
rect 1086 2452 1092 2453
rect 1148 2444 1150 2462
rect 1208 2458 1210 2469
rect 1336 2458 1338 2469
rect 1464 2458 1466 2469
rect 1206 2457 1212 2458
rect 1206 2453 1207 2457
rect 1211 2453 1212 2457
rect 1206 2452 1212 2453
rect 1334 2457 1340 2458
rect 1334 2453 1335 2457
rect 1339 2453 1340 2457
rect 1334 2452 1340 2453
rect 1462 2457 1468 2458
rect 1462 2453 1463 2457
rect 1467 2453 1468 2457
rect 1462 2452 1468 2453
rect 1824 2445 1826 2469
rect 1864 2461 1866 2485
rect 2088 2474 2090 2485
rect 2098 2483 2104 2484
rect 2098 2479 2099 2483
rect 2103 2479 2104 2483
rect 2098 2478 2104 2479
rect 2086 2473 2092 2474
rect 2086 2469 2087 2473
rect 2091 2469 2092 2473
rect 2100 2469 2102 2478
rect 2184 2474 2186 2485
rect 2288 2474 2290 2485
rect 2408 2474 2410 2485
rect 2544 2474 2546 2485
rect 2628 2484 2630 2522
rect 2702 2511 2708 2512
rect 2702 2507 2703 2511
rect 2707 2507 2708 2511
rect 2702 2506 2708 2507
rect 2704 2491 2706 2506
rect 2764 2500 2766 2522
rect 2854 2511 2860 2512
rect 2854 2507 2855 2511
rect 2859 2507 2860 2511
rect 2854 2506 2860 2507
rect 2762 2499 2768 2500
rect 2762 2495 2763 2499
rect 2767 2495 2768 2499
rect 2762 2494 2768 2495
rect 2856 2491 2858 2506
rect 2916 2500 2918 2522
rect 3006 2511 3012 2512
rect 3006 2507 3007 2511
rect 3011 2507 3012 2511
rect 3006 2506 3012 2507
rect 2914 2499 2920 2500
rect 2914 2495 2915 2499
rect 2919 2495 2920 2499
rect 2914 2494 2920 2495
rect 3008 2491 3010 2506
rect 3020 2500 3022 2562
rect 3151 2557 3155 2558
rect 3159 2562 3163 2563
rect 3159 2557 3163 2558
rect 3160 2552 3162 2557
rect 3158 2551 3164 2552
rect 3158 2547 3159 2551
rect 3163 2547 3164 2551
rect 3158 2546 3164 2547
rect 3168 2540 3170 2618
rect 3327 2562 3331 2563
rect 3327 2557 3331 2558
rect 3328 2552 3330 2557
rect 3326 2551 3332 2552
rect 3326 2547 3327 2551
rect 3331 2547 3332 2551
rect 3326 2546 3332 2547
rect 3166 2539 3172 2540
rect 3166 2535 3167 2539
rect 3171 2535 3172 2539
rect 3166 2534 3172 2535
rect 3226 2527 3232 2528
rect 3226 2523 3227 2527
rect 3231 2523 3232 2527
rect 3226 2522 3232 2523
rect 3166 2511 3172 2512
rect 3166 2507 3167 2511
rect 3171 2507 3172 2511
rect 3166 2506 3172 2507
rect 3018 2499 3024 2500
rect 3018 2495 3019 2499
rect 3023 2495 3024 2499
rect 3018 2494 3024 2495
rect 3168 2491 3170 2506
rect 3228 2500 3230 2522
rect 3334 2511 3340 2512
rect 3334 2507 3335 2511
rect 3339 2507 3340 2511
rect 3334 2506 3340 2507
rect 3226 2499 3232 2500
rect 3226 2495 3227 2499
rect 3231 2495 3232 2499
rect 3226 2494 3232 2495
rect 3336 2491 3338 2506
rect 3472 2500 3474 2678
rect 3486 2667 3492 2668
rect 3486 2663 3487 2667
rect 3491 2663 3492 2667
rect 3486 2662 3492 2663
rect 3488 2631 3490 2662
rect 3500 2656 3502 2718
rect 3575 2713 3579 2714
rect 3576 2698 3578 2713
rect 3574 2697 3580 2698
rect 3574 2693 3575 2697
rect 3579 2693 3580 2697
rect 3574 2692 3580 2693
rect 3574 2680 3580 2681
rect 3574 2676 3575 2680
rect 3579 2676 3580 2680
rect 3574 2675 3580 2676
rect 3498 2655 3504 2656
rect 3498 2651 3499 2655
rect 3503 2651 3504 2655
rect 3498 2650 3504 2651
rect 3576 2631 3578 2675
rect 3487 2630 3491 2631
rect 3487 2625 3491 2626
rect 3575 2630 3579 2631
rect 3575 2625 3579 2626
rect 3576 2601 3578 2625
rect 3574 2600 3580 2601
rect 3574 2596 3575 2600
rect 3579 2596 3580 2600
rect 3574 2595 3580 2596
rect 3574 2583 3580 2584
rect 3574 2579 3575 2583
rect 3579 2579 3580 2583
rect 3574 2578 3580 2579
rect 3576 2563 3578 2578
rect 3479 2562 3483 2563
rect 3479 2557 3483 2558
rect 3575 2562 3579 2563
rect 3575 2557 3579 2558
rect 3480 2552 3482 2557
rect 3478 2551 3484 2552
rect 3478 2547 3479 2551
rect 3483 2547 3484 2551
rect 3478 2546 3484 2547
rect 3576 2542 3578 2557
rect 3574 2541 3580 2542
rect 3574 2537 3575 2541
rect 3579 2537 3580 2541
rect 3574 2536 3580 2537
rect 3574 2524 3580 2525
rect 3574 2520 3575 2524
rect 3579 2520 3580 2524
rect 3574 2519 3580 2520
rect 3486 2511 3492 2512
rect 3486 2507 3487 2511
rect 3491 2507 3492 2511
rect 3486 2506 3492 2507
rect 3354 2499 3360 2500
rect 3354 2495 3355 2499
rect 3359 2495 3360 2499
rect 3354 2494 3360 2495
rect 3470 2499 3476 2500
rect 3470 2495 3471 2499
rect 3475 2495 3476 2499
rect 3470 2494 3476 2495
rect 2703 2490 2707 2491
rect 2703 2485 2707 2486
rect 2855 2490 2859 2491
rect 2855 2485 2859 2486
rect 2887 2490 2891 2491
rect 2887 2485 2891 2486
rect 3007 2490 3011 2491
rect 3007 2485 3011 2486
rect 3087 2490 3091 2491
rect 3087 2485 3091 2486
rect 3167 2490 3171 2491
rect 3167 2485 3171 2486
rect 3295 2490 3299 2491
rect 3295 2485 3299 2486
rect 3335 2490 3339 2491
rect 3335 2485 3339 2486
rect 2622 2483 2630 2484
rect 2622 2479 2623 2483
rect 2627 2481 2630 2483
rect 2627 2479 2628 2481
rect 2622 2478 2628 2479
rect 2704 2474 2706 2485
rect 2888 2474 2890 2485
rect 3088 2474 3090 2485
rect 3296 2474 3298 2485
rect 3302 2483 3308 2484
rect 3302 2479 3303 2483
rect 3307 2479 3308 2483
rect 3302 2478 3308 2479
rect 2182 2473 2188 2474
rect 2182 2469 2183 2473
rect 2187 2469 2188 2473
rect 2086 2468 2092 2469
rect 2099 2468 2103 2469
rect 2182 2468 2188 2469
rect 2286 2473 2292 2474
rect 2286 2469 2287 2473
rect 2291 2469 2292 2473
rect 2406 2473 2412 2474
rect 2406 2469 2407 2473
rect 2411 2469 2412 2473
rect 2286 2468 2292 2469
rect 2379 2468 2383 2469
rect 2406 2468 2412 2469
rect 2542 2473 2548 2474
rect 2542 2469 2543 2473
rect 2547 2469 2548 2473
rect 2542 2468 2548 2469
rect 2702 2473 2708 2474
rect 2702 2469 2703 2473
rect 2707 2469 2708 2473
rect 2702 2468 2708 2469
rect 2886 2473 2892 2474
rect 2886 2469 2887 2473
rect 2891 2469 2892 2473
rect 2886 2468 2892 2469
rect 3086 2473 3092 2474
rect 3086 2469 3087 2473
rect 3091 2469 3092 2473
rect 3086 2468 3092 2469
rect 3294 2473 3300 2474
rect 3294 2469 3295 2473
rect 3299 2469 3300 2473
rect 3294 2468 3300 2469
rect 2099 2463 2103 2464
rect 2379 2463 2383 2464
rect 1862 2460 1868 2461
rect 1862 2456 1863 2460
rect 1867 2456 1868 2460
rect 1862 2455 1868 2456
rect 1822 2444 1828 2445
rect 1146 2443 1152 2444
rect 786 2439 792 2440
rect 786 2435 787 2439
rect 791 2435 792 2439
rect 1146 2439 1147 2443
rect 1151 2439 1152 2443
rect 1822 2440 1823 2444
rect 1827 2440 1828 2444
rect 1822 2439 1828 2440
rect 1862 2443 1868 2444
rect 1862 2439 1863 2443
rect 1867 2439 1868 2443
rect 1146 2438 1152 2439
rect 1862 2438 1868 2439
rect 786 2434 792 2435
rect 1402 2427 1408 2428
rect 1402 2423 1403 2427
rect 1407 2423 1408 2427
rect 1402 2422 1408 2423
rect 1822 2427 1828 2428
rect 1822 2423 1823 2427
rect 1827 2423 1828 2427
rect 1822 2422 1828 2423
rect 838 2417 844 2418
rect 838 2413 839 2417
rect 843 2413 844 2417
rect 838 2412 844 2413
rect 958 2417 964 2418
rect 958 2413 959 2417
rect 963 2413 964 2417
rect 958 2412 964 2413
rect 1078 2417 1084 2418
rect 1078 2413 1079 2417
rect 1083 2413 1084 2417
rect 1078 2412 1084 2413
rect 1198 2417 1204 2418
rect 1198 2413 1199 2417
rect 1203 2413 1204 2417
rect 1198 2412 1204 2413
rect 1326 2417 1332 2418
rect 1326 2413 1327 2417
rect 1331 2413 1332 2417
rect 1326 2412 1332 2413
rect 840 2403 842 2412
rect 960 2403 962 2412
rect 1080 2403 1082 2412
rect 1200 2403 1202 2412
rect 1328 2403 1330 2412
rect 839 2402 843 2403
rect 839 2397 843 2398
rect 847 2402 851 2403
rect 847 2397 851 2398
rect 959 2402 963 2403
rect 959 2397 963 2398
rect 1031 2402 1035 2403
rect 1031 2397 1035 2398
rect 1079 2402 1083 2403
rect 1079 2397 1083 2398
rect 1199 2402 1203 2403
rect 1199 2397 1203 2398
rect 1207 2402 1211 2403
rect 1207 2397 1211 2398
rect 1327 2402 1331 2403
rect 1327 2397 1331 2398
rect 1375 2402 1379 2403
rect 1375 2397 1379 2398
rect 848 2392 850 2397
rect 1032 2392 1034 2397
rect 1208 2392 1210 2397
rect 1376 2392 1378 2397
rect 846 2391 852 2392
rect 846 2387 847 2391
rect 851 2387 852 2391
rect 846 2386 852 2387
rect 1030 2391 1036 2392
rect 1030 2387 1031 2391
rect 1035 2387 1036 2391
rect 1030 2386 1036 2387
rect 1206 2391 1212 2392
rect 1206 2387 1207 2391
rect 1211 2387 1212 2391
rect 1206 2386 1212 2387
rect 1374 2391 1380 2392
rect 1374 2387 1375 2391
rect 1379 2387 1380 2391
rect 1374 2386 1380 2387
rect 730 2383 736 2384
rect 730 2379 731 2383
rect 735 2379 736 2383
rect 730 2378 736 2379
rect 730 2367 736 2368
rect 730 2363 731 2367
rect 735 2363 736 2367
rect 730 2362 736 2363
rect 670 2351 676 2352
rect 670 2347 671 2351
rect 675 2347 676 2351
rect 670 2346 676 2347
rect 490 2339 496 2340
rect 490 2335 491 2339
rect 495 2335 496 2339
rect 490 2334 496 2335
rect 672 2331 674 2346
rect 732 2340 734 2362
rect 854 2351 860 2352
rect 854 2347 855 2351
rect 859 2347 860 2351
rect 854 2346 860 2347
rect 1038 2351 1044 2352
rect 1038 2347 1039 2351
rect 1043 2347 1044 2351
rect 1214 2351 1220 2352
rect 1038 2346 1044 2347
rect 1095 2348 1099 2349
rect 730 2339 736 2340
rect 730 2335 731 2339
rect 735 2335 736 2339
rect 730 2334 736 2335
rect 846 2339 852 2340
rect 846 2335 847 2339
rect 851 2335 852 2339
rect 846 2334 852 2335
rect 111 2330 115 2331
rect 111 2325 115 2326
rect 143 2330 147 2331
rect 143 2325 147 2326
rect 295 2330 299 2331
rect 295 2325 299 2326
rect 479 2330 483 2331
rect 479 2325 483 2326
rect 671 2330 675 2331
rect 671 2325 675 2326
rect 112 2301 114 2325
rect 144 2314 146 2325
rect 226 2323 232 2324
rect 226 2319 227 2323
rect 231 2319 232 2323
rect 226 2318 232 2319
rect 142 2313 148 2314
rect 142 2309 143 2313
rect 147 2309 148 2313
rect 142 2308 148 2309
rect 110 2300 116 2301
rect 110 2296 111 2300
rect 115 2296 116 2300
rect 228 2296 230 2318
rect 296 2314 298 2325
rect 480 2314 482 2325
rect 490 2323 496 2324
rect 490 2319 491 2323
rect 495 2319 496 2323
rect 490 2318 496 2319
rect 294 2313 300 2314
rect 294 2309 295 2313
rect 299 2309 300 2313
rect 294 2308 300 2309
rect 478 2313 484 2314
rect 478 2309 479 2313
rect 483 2309 484 2313
rect 478 2308 484 2309
rect 110 2295 116 2296
rect 226 2295 232 2296
rect 226 2291 227 2295
rect 231 2291 232 2295
rect 226 2290 232 2291
rect 110 2283 116 2284
rect 110 2279 111 2283
rect 115 2279 116 2283
rect 110 2278 116 2279
rect 112 2255 114 2278
rect 134 2273 140 2274
rect 134 2269 135 2273
rect 139 2269 140 2273
rect 134 2268 140 2269
rect 286 2273 292 2274
rect 286 2269 287 2273
rect 291 2269 292 2273
rect 286 2268 292 2269
rect 470 2273 476 2274
rect 470 2269 471 2273
rect 475 2269 476 2273
rect 470 2268 476 2269
rect 136 2255 138 2268
rect 154 2267 160 2268
rect 154 2263 155 2267
rect 159 2263 160 2267
rect 154 2262 160 2263
rect 111 2254 115 2255
rect 111 2249 115 2250
rect 135 2254 139 2255
rect 135 2249 139 2250
rect 112 2234 114 2249
rect 136 2244 138 2249
rect 134 2243 140 2244
rect 134 2239 135 2243
rect 139 2239 140 2243
rect 134 2238 140 2239
rect 110 2233 116 2234
rect 110 2229 111 2233
rect 115 2229 116 2233
rect 110 2228 116 2229
rect 110 2216 116 2217
rect 110 2212 111 2216
rect 115 2212 116 2216
rect 110 2211 116 2212
rect 112 2183 114 2211
rect 142 2203 148 2204
rect 142 2199 143 2203
rect 147 2199 148 2203
rect 142 2198 148 2199
rect 144 2183 146 2198
rect 156 2192 158 2262
rect 288 2255 290 2268
rect 472 2255 474 2268
rect 255 2254 259 2255
rect 255 2249 259 2250
rect 287 2254 291 2255
rect 287 2249 291 2250
rect 407 2254 411 2255
rect 407 2249 411 2250
rect 471 2254 475 2255
rect 471 2249 475 2250
rect 256 2244 258 2249
rect 408 2244 410 2249
rect 254 2243 260 2244
rect 254 2239 255 2243
rect 259 2239 260 2243
rect 254 2238 260 2239
rect 406 2243 412 2244
rect 406 2239 407 2243
rect 411 2239 412 2243
rect 406 2238 412 2239
rect 492 2236 494 2318
rect 672 2314 674 2325
rect 670 2313 676 2314
rect 670 2309 671 2313
rect 675 2309 676 2313
rect 670 2308 676 2309
rect 848 2296 850 2334
rect 856 2331 858 2346
rect 1040 2331 1042 2346
rect 1214 2347 1215 2351
rect 1219 2347 1220 2351
rect 1214 2346 1220 2347
rect 1382 2351 1388 2352
rect 1382 2347 1383 2351
rect 1387 2347 1388 2351
rect 1404 2349 1406 2422
rect 1454 2417 1460 2418
rect 1454 2413 1455 2417
rect 1459 2413 1460 2417
rect 1454 2412 1460 2413
rect 1456 2403 1458 2412
rect 1824 2403 1826 2422
rect 1864 2419 1866 2438
rect 2078 2433 2084 2434
rect 2078 2429 2079 2433
rect 2083 2429 2084 2433
rect 2078 2428 2084 2429
rect 2174 2433 2180 2434
rect 2174 2429 2175 2433
rect 2179 2429 2180 2433
rect 2174 2428 2180 2429
rect 2278 2433 2284 2434
rect 2278 2429 2279 2433
rect 2283 2429 2284 2433
rect 2278 2428 2284 2429
rect 2080 2419 2082 2428
rect 2176 2419 2178 2428
rect 2280 2419 2282 2428
rect 1863 2418 1867 2419
rect 1863 2413 1867 2414
rect 1951 2418 1955 2419
rect 1951 2413 1955 2414
rect 2063 2418 2067 2419
rect 2063 2413 2067 2414
rect 2079 2418 2083 2419
rect 2079 2413 2083 2414
rect 2175 2418 2179 2419
rect 2175 2413 2179 2414
rect 2183 2418 2187 2419
rect 2183 2413 2187 2414
rect 2279 2418 2283 2419
rect 2279 2413 2283 2414
rect 2311 2418 2315 2419
rect 2311 2413 2315 2414
rect 1455 2402 1459 2403
rect 1455 2397 1459 2398
rect 1543 2402 1547 2403
rect 1543 2397 1547 2398
rect 1711 2402 1715 2403
rect 1711 2397 1715 2398
rect 1823 2402 1827 2403
rect 1864 2398 1866 2413
rect 1952 2408 1954 2413
rect 2064 2408 2066 2413
rect 2184 2408 2186 2413
rect 2312 2408 2314 2413
rect 1950 2407 1956 2408
rect 1950 2403 1951 2407
rect 1955 2403 1956 2407
rect 1950 2402 1956 2403
rect 2062 2407 2068 2408
rect 2062 2403 2063 2407
rect 2067 2403 2068 2407
rect 2062 2402 2068 2403
rect 2182 2407 2188 2408
rect 2182 2403 2183 2407
rect 2187 2403 2188 2407
rect 2182 2402 2188 2403
rect 2310 2407 2316 2408
rect 2310 2403 2311 2407
rect 2315 2403 2316 2407
rect 2310 2402 2316 2403
rect 2380 2400 2382 2463
rect 3304 2459 3306 2478
rect 3356 2460 3358 2494
rect 3488 2491 3490 2506
rect 3576 2491 3578 2519
rect 3487 2490 3491 2491
rect 3487 2485 3491 2486
rect 3575 2490 3579 2491
rect 3575 2485 3579 2486
rect 3488 2474 3490 2485
rect 3486 2473 3492 2474
rect 3486 2469 3487 2473
rect 3491 2469 3492 2473
rect 3486 2468 3492 2469
rect 3576 2461 3578 2485
rect 3574 2460 3580 2461
rect 3296 2457 3306 2459
rect 3354 2459 3360 2460
rect 2954 2443 2960 2444
rect 2954 2439 2955 2443
rect 2959 2439 2960 2443
rect 2954 2438 2960 2439
rect 2398 2433 2404 2434
rect 2398 2429 2399 2433
rect 2403 2429 2404 2433
rect 2398 2428 2404 2429
rect 2534 2433 2540 2434
rect 2534 2429 2535 2433
rect 2539 2429 2540 2433
rect 2534 2428 2540 2429
rect 2694 2433 2700 2434
rect 2694 2429 2695 2433
rect 2699 2429 2700 2433
rect 2694 2428 2700 2429
rect 2878 2433 2884 2434
rect 2878 2429 2879 2433
rect 2883 2429 2884 2433
rect 2878 2428 2884 2429
rect 2400 2419 2402 2428
rect 2536 2419 2538 2428
rect 2610 2419 2616 2420
rect 2696 2419 2698 2428
rect 2880 2419 2882 2428
rect 2956 2420 2958 2438
rect 3078 2433 3084 2434
rect 3078 2429 3079 2433
rect 3083 2429 3084 2433
rect 3078 2428 3084 2429
rect 3286 2433 3292 2434
rect 3286 2429 3287 2433
rect 3291 2429 3292 2433
rect 3286 2428 3292 2429
rect 2954 2419 2960 2420
rect 3080 2419 3082 2428
rect 3288 2419 3290 2428
rect 2399 2418 2403 2419
rect 2399 2413 2403 2414
rect 2447 2418 2451 2419
rect 2447 2413 2451 2414
rect 2535 2418 2539 2419
rect 2535 2413 2539 2414
rect 2591 2418 2595 2419
rect 2610 2415 2611 2419
rect 2615 2415 2616 2419
rect 2610 2414 2616 2415
rect 2695 2418 2699 2419
rect 2591 2413 2595 2414
rect 2448 2408 2450 2413
rect 2592 2408 2594 2413
rect 2446 2407 2452 2408
rect 2446 2403 2447 2407
rect 2451 2403 2452 2407
rect 2446 2402 2452 2403
rect 2590 2407 2596 2408
rect 2590 2403 2591 2407
rect 2595 2403 2596 2407
rect 2590 2402 2596 2403
rect 2378 2399 2384 2400
rect 1823 2397 1827 2398
rect 1862 2397 1868 2398
rect 1544 2392 1546 2397
rect 1712 2392 1714 2397
rect 1542 2391 1548 2392
rect 1542 2387 1543 2391
rect 1547 2387 1548 2391
rect 1542 2386 1548 2387
rect 1710 2391 1716 2392
rect 1710 2387 1711 2391
rect 1715 2387 1716 2391
rect 1710 2386 1716 2387
rect 1824 2382 1826 2397
rect 1862 2393 1863 2397
rect 1867 2393 1868 2397
rect 2378 2395 2379 2399
rect 2383 2395 2384 2399
rect 2378 2394 2384 2395
rect 1862 2392 1868 2393
rect 1822 2381 1828 2382
rect 1822 2377 1823 2381
rect 1827 2377 1828 2381
rect 1822 2376 1828 2377
rect 1862 2380 1868 2381
rect 1862 2376 1863 2380
rect 1867 2376 1868 2380
rect 1862 2375 1868 2376
rect 1778 2367 1784 2368
rect 1778 2363 1779 2367
rect 1783 2363 1784 2367
rect 1778 2362 1784 2363
rect 1822 2364 1828 2365
rect 1550 2351 1556 2352
rect 1382 2346 1388 2347
rect 1403 2348 1407 2349
rect 1095 2343 1099 2344
rect 1096 2340 1098 2343
rect 1094 2339 1100 2340
rect 1094 2335 1095 2339
rect 1099 2335 1100 2339
rect 1094 2334 1100 2335
rect 1216 2331 1218 2346
rect 1384 2331 1386 2346
rect 1550 2347 1551 2351
rect 1555 2347 1556 2351
rect 1550 2346 1556 2347
rect 1718 2351 1724 2352
rect 1718 2347 1719 2351
rect 1723 2347 1724 2351
rect 1718 2346 1724 2347
rect 1403 2343 1407 2344
rect 1552 2331 1554 2346
rect 1720 2331 1722 2346
rect 855 2330 859 2331
rect 855 2325 859 2326
rect 863 2330 867 2331
rect 863 2325 867 2326
rect 1039 2330 1043 2331
rect 1039 2325 1043 2326
rect 1055 2330 1059 2331
rect 1055 2325 1059 2326
rect 1215 2330 1219 2331
rect 1215 2325 1219 2326
rect 1231 2330 1235 2331
rect 1231 2325 1235 2326
rect 1383 2330 1387 2331
rect 1383 2325 1387 2326
rect 1407 2330 1411 2331
rect 1407 2325 1411 2326
rect 1551 2330 1555 2331
rect 1551 2325 1555 2326
rect 1583 2330 1587 2331
rect 1583 2325 1587 2326
rect 1719 2330 1723 2331
rect 1719 2325 1723 2326
rect 1735 2330 1739 2331
rect 1735 2325 1739 2326
rect 864 2314 866 2325
rect 1056 2314 1058 2325
rect 1150 2323 1156 2324
rect 1150 2319 1151 2323
rect 1155 2319 1156 2323
rect 1150 2318 1156 2319
rect 862 2313 868 2314
rect 862 2309 863 2313
rect 867 2309 868 2313
rect 862 2308 868 2309
rect 1054 2313 1060 2314
rect 1054 2309 1055 2313
rect 1059 2309 1060 2313
rect 1054 2308 1060 2309
rect 1152 2301 1154 2318
rect 1232 2314 1234 2325
rect 1408 2314 1410 2325
rect 1584 2314 1586 2325
rect 1650 2323 1656 2324
rect 1650 2319 1651 2323
rect 1655 2319 1656 2323
rect 1650 2318 1656 2319
rect 1230 2313 1236 2314
rect 1230 2309 1231 2313
rect 1235 2309 1236 2313
rect 1230 2308 1236 2309
rect 1406 2313 1412 2314
rect 1406 2309 1407 2313
rect 1411 2309 1412 2313
rect 1406 2308 1412 2309
rect 1582 2313 1588 2314
rect 1582 2309 1583 2313
rect 1587 2309 1588 2313
rect 1582 2308 1588 2309
rect 1151 2300 1155 2301
rect 1339 2300 1343 2301
rect 1652 2296 1654 2318
rect 1736 2314 1738 2325
rect 1780 2324 1782 2362
rect 1822 2360 1823 2364
rect 1827 2360 1828 2364
rect 1822 2359 1828 2360
rect 1824 2331 1826 2359
rect 1864 2343 1866 2375
rect 1958 2367 1964 2368
rect 1958 2363 1959 2367
rect 1963 2363 1964 2367
rect 1958 2362 1964 2363
rect 2070 2367 2076 2368
rect 2070 2363 2071 2367
rect 2075 2363 2076 2367
rect 2070 2362 2076 2363
rect 2190 2367 2196 2368
rect 2190 2363 2191 2367
rect 2195 2363 2196 2367
rect 2190 2362 2196 2363
rect 2318 2367 2324 2368
rect 2318 2363 2319 2367
rect 2323 2363 2324 2367
rect 2318 2362 2324 2363
rect 2454 2367 2460 2368
rect 2454 2363 2455 2367
rect 2459 2363 2460 2367
rect 2454 2362 2460 2363
rect 2598 2367 2604 2368
rect 2598 2363 2599 2367
rect 2603 2363 2604 2367
rect 2598 2362 2604 2363
rect 1960 2343 1962 2362
rect 2046 2355 2052 2356
rect 2046 2351 2047 2355
rect 2051 2351 2052 2355
rect 2046 2350 2052 2351
rect 1863 2342 1867 2343
rect 1863 2337 1867 2338
rect 1895 2342 1899 2343
rect 1895 2337 1899 2338
rect 1959 2342 1963 2343
rect 1959 2337 1963 2338
rect 2007 2342 2011 2343
rect 2007 2337 2011 2338
rect 1823 2330 1827 2331
rect 1823 2325 1827 2326
rect 1778 2323 1784 2324
rect 1778 2319 1779 2323
rect 1783 2319 1784 2323
rect 1778 2318 1784 2319
rect 1734 2313 1740 2314
rect 1734 2309 1735 2313
rect 1739 2309 1740 2313
rect 1734 2308 1740 2309
rect 1824 2301 1826 2325
rect 1864 2313 1866 2337
rect 1896 2326 1898 2337
rect 1950 2335 1956 2336
rect 1950 2331 1951 2335
rect 1955 2331 1956 2335
rect 1950 2330 1956 2331
rect 1894 2325 1900 2326
rect 1894 2321 1895 2325
rect 1899 2321 1900 2325
rect 1894 2320 1900 2321
rect 1862 2312 1868 2313
rect 1862 2308 1863 2312
rect 1867 2308 1868 2312
rect 1862 2307 1868 2308
rect 1822 2300 1828 2301
rect 1822 2296 1823 2300
rect 1827 2296 1828 2300
rect 846 2295 852 2296
rect 1151 2295 1155 2296
rect 1338 2295 1344 2296
rect 846 2291 847 2295
rect 851 2291 852 2295
rect 846 2290 852 2291
rect 1338 2291 1339 2295
rect 1343 2291 1344 2295
rect 1338 2290 1344 2291
rect 1650 2295 1656 2296
rect 1822 2295 1828 2296
rect 1862 2295 1868 2296
rect 1650 2291 1651 2295
rect 1655 2291 1656 2295
rect 1650 2290 1656 2291
rect 1862 2291 1863 2295
rect 1867 2291 1868 2295
rect 1862 2290 1868 2291
rect 1318 2283 1324 2284
rect 1318 2279 1319 2283
rect 1323 2279 1324 2283
rect 1318 2278 1324 2279
rect 1822 2283 1828 2284
rect 1822 2279 1823 2283
rect 1827 2279 1828 2283
rect 1822 2278 1828 2279
rect 662 2273 668 2274
rect 662 2269 663 2273
rect 667 2269 668 2273
rect 662 2268 668 2269
rect 854 2273 860 2274
rect 854 2269 855 2273
rect 859 2269 860 2273
rect 854 2268 860 2269
rect 1046 2273 1052 2274
rect 1046 2269 1047 2273
rect 1051 2269 1052 2273
rect 1046 2268 1052 2269
rect 1222 2273 1228 2274
rect 1222 2269 1223 2273
rect 1227 2269 1228 2273
rect 1222 2268 1228 2269
rect 664 2255 666 2268
rect 856 2255 858 2268
rect 1048 2255 1050 2268
rect 1224 2255 1226 2268
rect 559 2254 563 2255
rect 559 2249 563 2250
rect 663 2254 667 2255
rect 663 2249 667 2250
rect 719 2254 723 2255
rect 719 2249 723 2250
rect 855 2254 859 2255
rect 855 2249 859 2250
rect 871 2254 875 2255
rect 871 2249 875 2250
rect 1015 2254 1019 2255
rect 1015 2249 1019 2250
rect 1047 2254 1051 2255
rect 1047 2249 1051 2250
rect 1159 2254 1163 2255
rect 1159 2249 1163 2250
rect 1223 2254 1227 2255
rect 1223 2249 1227 2250
rect 1303 2254 1307 2255
rect 1303 2249 1307 2250
rect 560 2244 562 2249
rect 720 2244 722 2249
rect 872 2244 874 2249
rect 1016 2244 1018 2249
rect 1160 2244 1162 2249
rect 1304 2244 1306 2249
rect 558 2243 564 2244
rect 558 2239 559 2243
rect 563 2239 564 2243
rect 558 2238 564 2239
rect 718 2243 724 2244
rect 718 2239 719 2243
rect 723 2239 724 2243
rect 718 2238 724 2239
rect 870 2243 876 2244
rect 870 2239 871 2243
rect 875 2239 876 2243
rect 870 2238 876 2239
rect 1014 2243 1020 2244
rect 1014 2239 1015 2243
rect 1019 2239 1020 2243
rect 1014 2238 1020 2239
rect 1158 2243 1164 2244
rect 1158 2239 1159 2243
rect 1163 2239 1164 2243
rect 1158 2238 1164 2239
rect 1302 2243 1308 2244
rect 1302 2239 1303 2243
rect 1307 2239 1308 2243
rect 1302 2238 1308 2239
rect 374 2235 380 2236
rect 374 2231 375 2235
rect 379 2231 380 2235
rect 374 2230 380 2231
rect 490 2235 496 2236
rect 490 2231 491 2235
rect 495 2231 496 2235
rect 490 2230 496 2231
rect 262 2203 268 2204
rect 262 2199 263 2203
rect 267 2199 268 2203
rect 262 2198 268 2199
rect 154 2191 160 2192
rect 154 2187 155 2191
rect 159 2187 160 2191
rect 154 2186 160 2187
rect 264 2183 266 2198
rect 376 2184 378 2230
rect 626 2219 632 2220
rect 626 2215 627 2219
rect 631 2215 632 2219
rect 626 2214 632 2215
rect 1082 2219 1088 2220
rect 1082 2215 1083 2219
rect 1087 2215 1088 2219
rect 1082 2214 1088 2215
rect 1098 2219 1104 2220
rect 1098 2215 1099 2219
rect 1103 2215 1104 2219
rect 1098 2214 1104 2215
rect 414 2203 420 2204
rect 414 2199 415 2203
rect 419 2199 420 2203
rect 414 2198 420 2199
rect 566 2203 572 2204
rect 566 2199 567 2203
rect 571 2199 572 2203
rect 566 2198 572 2199
rect 374 2183 380 2184
rect 416 2183 418 2198
rect 568 2183 570 2198
rect 628 2192 630 2214
rect 726 2203 732 2204
rect 726 2199 727 2203
rect 731 2199 732 2203
rect 726 2198 732 2199
rect 878 2203 884 2204
rect 878 2199 879 2203
rect 883 2199 884 2203
rect 878 2198 884 2199
rect 1022 2203 1028 2204
rect 1022 2199 1023 2203
rect 1027 2199 1028 2203
rect 1022 2198 1028 2199
rect 626 2191 632 2192
rect 626 2187 627 2191
rect 631 2187 632 2191
rect 626 2186 632 2187
rect 728 2183 730 2198
rect 880 2183 882 2198
rect 891 2196 895 2197
rect 890 2191 896 2192
rect 890 2187 891 2191
rect 895 2187 896 2191
rect 890 2186 896 2187
rect 898 2183 904 2184
rect 1024 2183 1026 2198
rect 111 2182 115 2183
rect 111 2177 115 2178
rect 143 2182 147 2183
rect 143 2177 147 2178
rect 215 2182 219 2183
rect 215 2177 219 2178
rect 263 2182 267 2183
rect 263 2177 267 2178
rect 311 2182 315 2183
rect 374 2179 375 2183
rect 379 2179 380 2183
rect 374 2178 380 2179
rect 415 2182 419 2183
rect 311 2177 315 2178
rect 415 2177 419 2178
rect 519 2182 523 2183
rect 519 2177 523 2178
rect 567 2182 571 2183
rect 567 2177 571 2178
rect 623 2182 627 2183
rect 623 2177 627 2178
rect 727 2182 731 2183
rect 727 2177 731 2178
rect 831 2182 835 2183
rect 831 2177 835 2178
rect 879 2182 883 2183
rect 898 2179 899 2183
rect 903 2179 904 2183
rect 898 2178 904 2179
rect 943 2182 947 2183
rect 879 2177 883 2178
rect 112 2153 114 2177
rect 216 2166 218 2177
rect 312 2166 314 2177
rect 416 2166 418 2177
rect 490 2167 496 2168
rect 214 2165 220 2166
rect 214 2161 215 2165
rect 219 2161 220 2165
rect 214 2160 220 2161
rect 310 2165 316 2166
rect 310 2161 311 2165
rect 315 2161 316 2165
rect 310 2160 316 2161
rect 414 2165 420 2166
rect 414 2161 415 2165
rect 419 2161 420 2165
rect 490 2163 491 2167
rect 495 2163 496 2167
rect 520 2166 522 2177
rect 624 2166 626 2177
rect 728 2166 730 2177
rect 832 2166 834 2177
rect 490 2162 496 2163
rect 518 2165 524 2166
rect 414 2160 420 2161
rect 110 2152 116 2153
rect 110 2148 111 2152
rect 115 2148 116 2152
rect 110 2147 116 2148
rect 110 2135 116 2136
rect 110 2131 111 2135
rect 115 2131 116 2135
rect 110 2130 116 2131
rect 112 2107 114 2130
rect 206 2125 212 2126
rect 206 2121 207 2125
rect 211 2121 212 2125
rect 206 2120 212 2121
rect 302 2125 308 2126
rect 302 2121 303 2125
rect 307 2121 308 2125
rect 302 2120 308 2121
rect 406 2125 412 2126
rect 406 2121 407 2125
rect 411 2121 412 2125
rect 406 2120 412 2121
rect 208 2107 210 2120
rect 304 2107 306 2120
rect 338 2119 344 2120
rect 338 2115 339 2119
rect 343 2115 344 2119
rect 338 2114 344 2115
rect 111 2106 115 2107
rect 111 2101 115 2102
rect 207 2106 211 2107
rect 207 2101 211 2102
rect 303 2106 307 2107
rect 303 2101 307 2102
rect 319 2106 323 2107
rect 319 2101 323 2102
rect 112 2086 114 2101
rect 320 2096 322 2101
rect 318 2095 324 2096
rect 318 2091 319 2095
rect 323 2091 324 2095
rect 318 2090 324 2091
rect 110 2085 116 2086
rect 110 2081 111 2085
rect 115 2081 116 2085
rect 110 2080 116 2081
rect 110 2068 116 2069
rect 110 2064 111 2068
rect 115 2064 116 2068
rect 110 2063 116 2064
rect 112 2031 114 2063
rect 326 2055 332 2056
rect 326 2051 327 2055
rect 331 2051 332 2055
rect 326 2050 332 2051
rect 328 2031 330 2050
rect 340 2044 342 2114
rect 408 2107 410 2120
rect 407 2106 411 2107
rect 407 2101 411 2102
rect 423 2106 427 2107
rect 423 2101 427 2102
rect 424 2096 426 2101
rect 422 2095 428 2096
rect 422 2091 423 2095
rect 427 2091 428 2095
rect 422 2090 428 2091
rect 492 2088 494 2162
rect 518 2161 519 2165
rect 523 2161 524 2165
rect 518 2160 524 2161
rect 622 2165 628 2166
rect 622 2161 623 2165
rect 627 2161 628 2165
rect 622 2160 628 2161
rect 726 2165 732 2166
rect 726 2161 727 2165
rect 731 2161 732 2165
rect 726 2160 732 2161
rect 830 2165 836 2166
rect 830 2161 831 2165
rect 835 2161 836 2165
rect 830 2160 836 2161
rect 900 2148 902 2178
rect 943 2177 947 2178
rect 1023 2182 1027 2183
rect 1023 2177 1027 2178
rect 1055 2182 1059 2183
rect 1055 2177 1059 2178
rect 944 2166 946 2177
rect 1056 2166 1058 2177
rect 1084 2176 1086 2214
rect 1100 2197 1102 2214
rect 1166 2203 1172 2204
rect 1166 2199 1167 2203
rect 1171 2199 1172 2203
rect 1166 2198 1172 2199
rect 1310 2203 1316 2204
rect 1310 2199 1311 2203
rect 1315 2199 1316 2203
rect 1310 2198 1316 2199
rect 1099 2196 1103 2197
rect 1099 2191 1103 2192
rect 1168 2183 1170 2198
rect 1191 2196 1195 2197
rect 1190 2191 1196 2192
rect 1190 2187 1191 2191
rect 1195 2187 1196 2191
rect 1190 2186 1196 2187
rect 1312 2183 1314 2198
rect 1320 2192 1322 2278
rect 1398 2273 1404 2274
rect 1398 2269 1399 2273
rect 1403 2269 1404 2273
rect 1398 2268 1404 2269
rect 1574 2273 1580 2274
rect 1574 2269 1575 2273
rect 1579 2269 1580 2273
rect 1574 2268 1580 2269
rect 1726 2273 1732 2274
rect 1726 2269 1727 2273
rect 1731 2269 1732 2273
rect 1726 2268 1732 2269
rect 1400 2255 1402 2268
rect 1576 2255 1578 2268
rect 1728 2255 1730 2268
rect 1824 2255 1826 2278
rect 1864 2271 1866 2290
rect 1886 2285 1892 2286
rect 1886 2281 1887 2285
rect 1891 2281 1892 2285
rect 1886 2280 1892 2281
rect 1888 2271 1890 2280
rect 1863 2270 1867 2271
rect 1863 2265 1867 2266
rect 1887 2270 1891 2271
rect 1887 2265 1891 2266
rect 1399 2254 1403 2255
rect 1399 2249 1403 2250
rect 1455 2254 1459 2255
rect 1455 2249 1459 2250
rect 1575 2254 1579 2255
rect 1575 2249 1579 2250
rect 1727 2254 1731 2255
rect 1727 2249 1731 2250
rect 1823 2254 1827 2255
rect 1864 2250 1866 2265
rect 1888 2260 1890 2265
rect 1886 2259 1892 2260
rect 1886 2255 1887 2259
rect 1891 2255 1892 2259
rect 1886 2254 1892 2255
rect 1952 2253 1954 2330
rect 2008 2326 2010 2337
rect 2006 2325 2012 2326
rect 2048 2325 2050 2350
rect 2072 2343 2074 2362
rect 2192 2343 2194 2362
rect 2320 2343 2322 2362
rect 2456 2343 2458 2362
rect 2600 2343 2602 2362
rect 2612 2356 2614 2414
rect 2695 2413 2699 2414
rect 2751 2418 2755 2419
rect 2751 2413 2755 2414
rect 2879 2418 2883 2419
rect 2879 2413 2883 2414
rect 2927 2418 2931 2419
rect 2954 2415 2955 2419
rect 2959 2415 2960 2419
rect 2954 2414 2960 2415
rect 3079 2418 3083 2419
rect 2927 2413 2931 2414
rect 3079 2413 3083 2414
rect 3111 2418 3115 2419
rect 3111 2413 3115 2414
rect 3287 2418 3291 2419
rect 3287 2413 3291 2414
rect 2752 2408 2754 2413
rect 2928 2408 2930 2413
rect 3112 2408 3114 2413
rect 2750 2407 2756 2408
rect 2750 2403 2751 2407
rect 2755 2403 2756 2407
rect 2750 2402 2756 2403
rect 2926 2407 2932 2408
rect 2926 2403 2927 2407
rect 2931 2403 2932 2407
rect 2926 2402 2932 2403
rect 3110 2407 3116 2408
rect 3110 2403 3111 2407
rect 3115 2403 3116 2407
rect 3110 2402 3116 2403
rect 3296 2400 3298 2457
rect 3354 2455 3355 2459
rect 3359 2455 3360 2459
rect 3574 2456 3575 2460
rect 3579 2456 3580 2460
rect 3574 2455 3580 2456
rect 3354 2454 3360 2455
rect 3574 2443 3580 2444
rect 3574 2439 3575 2443
rect 3579 2439 3580 2443
rect 3574 2438 3580 2439
rect 3478 2433 3484 2434
rect 3478 2429 3479 2433
rect 3483 2429 3484 2433
rect 3478 2428 3484 2429
rect 3480 2419 3482 2428
rect 3498 2427 3504 2428
rect 3498 2423 3499 2427
rect 3503 2423 3504 2427
rect 3498 2422 3504 2423
rect 3303 2418 3307 2419
rect 3303 2413 3307 2414
rect 3479 2418 3483 2419
rect 3479 2413 3483 2414
rect 3304 2408 3306 2413
rect 3480 2408 3482 2413
rect 3302 2407 3308 2408
rect 3302 2403 3303 2407
rect 3307 2403 3308 2407
rect 3302 2402 3308 2403
rect 3478 2407 3484 2408
rect 3478 2403 3479 2407
rect 3483 2403 3484 2407
rect 3478 2402 3484 2403
rect 3018 2399 3024 2400
rect 3018 2395 3019 2399
rect 3023 2395 3024 2399
rect 3018 2394 3024 2395
rect 3294 2399 3300 2400
rect 3294 2395 3295 2399
rect 3299 2395 3300 2399
rect 3294 2394 3300 2395
rect 2758 2367 2764 2368
rect 2758 2363 2759 2367
rect 2763 2363 2764 2367
rect 2758 2362 2764 2363
rect 2934 2367 2940 2368
rect 2934 2363 2935 2367
rect 2939 2363 2940 2367
rect 2934 2362 2940 2363
rect 2610 2355 2616 2356
rect 2610 2351 2611 2355
rect 2615 2351 2616 2355
rect 2610 2350 2616 2351
rect 2760 2343 2762 2362
rect 2936 2343 2938 2362
rect 3020 2344 3022 2394
rect 3118 2367 3124 2368
rect 3118 2363 3119 2367
rect 3123 2363 3124 2367
rect 3118 2362 3124 2363
rect 3310 2367 3316 2368
rect 3310 2363 3311 2367
rect 3315 2363 3316 2367
rect 3310 2362 3316 2363
rect 3486 2367 3492 2368
rect 3486 2363 3487 2367
rect 3491 2363 3492 2367
rect 3486 2362 3492 2363
rect 3018 2343 3024 2344
rect 3120 2343 3122 2362
rect 3312 2343 3314 2362
rect 3488 2343 3490 2362
rect 3500 2356 3502 2422
rect 3576 2419 3578 2438
rect 3575 2418 3579 2419
rect 3575 2413 3579 2414
rect 3576 2398 3578 2413
rect 3574 2397 3580 2398
rect 3574 2393 3575 2397
rect 3579 2393 3580 2397
rect 3574 2392 3580 2393
rect 3574 2380 3580 2381
rect 3574 2376 3575 2380
rect 3579 2376 3580 2380
rect 3574 2375 3580 2376
rect 3498 2355 3504 2356
rect 3498 2351 3499 2355
rect 3503 2351 3504 2355
rect 3498 2350 3504 2351
rect 3576 2343 3578 2375
rect 2071 2342 2075 2343
rect 2071 2337 2075 2338
rect 2159 2342 2163 2343
rect 2159 2337 2163 2338
rect 2191 2342 2195 2343
rect 2191 2337 2195 2338
rect 2311 2342 2315 2343
rect 2311 2337 2315 2338
rect 2319 2342 2323 2343
rect 2319 2337 2323 2338
rect 2455 2342 2459 2343
rect 2455 2337 2459 2338
rect 2463 2342 2467 2343
rect 2463 2337 2467 2338
rect 2599 2342 2603 2343
rect 2599 2337 2603 2338
rect 2615 2342 2619 2343
rect 2615 2337 2619 2338
rect 2759 2342 2763 2343
rect 2759 2337 2763 2338
rect 2775 2342 2779 2343
rect 2775 2337 2779 2338
rect 2935 2342 2939 2343
rect 2935 2337 2939 2338
rect 2943 2342 2947 2343
rect 3018 2339 3019 2343
rect 3023 2339 3024 2343
rect 3018 2338 3024 2339
rect 3111 2342 3115 2343
rect 2943 2337 2947 2338
rect 3111 2337 3115 2338
rect 3119 2342 3123 2343
rect 3119 2337 3123 2338
rect 3287 2342 3291 2343
rect 3287 2337 3291 2338
rect 3311 2342 3315 2343
rect 3311 2337 3315 2338
rect 3471 2342 3475 2343
rect 3471 2337 3475 2338
rect 3487 2342 3491 2343
rect 3487 2337 3491 2338
rect 3575 2342 3579 2343
rect 3575 2337 3579 2338
rect 2160 2326 2162 2337
rect 2312 2326 2314 2337
rect 2464 2326 2466 2337
rect 2616 2326 2618 2337
rect 2776 2326 2778 2337
rect 2874 2335 2880 2336
rect 2874 2331 2875 2335
rect 2879 2331 2880 2335
rect 2874 2330 2880 2331
rect 2158 2325 2164 2326
rect 2006 2321 2007 2325
rect 2011 2321 2012 2325
rect 2006 2320 2012 2321
rect 2047 2324 2051 2325
rect 2158 2321 2159 2325
rect 2163 2321 2164 2325
rect 2158 2320 2164 2321
rect 2310 2325 2316 2326
rect 2462 2325 2468 2326
rect 2310 2321 2311 2325
rect 2315 2321 2316 2325
rect 2310 2320 2316 2321
rect 2403 2324 2407 2325
rect 2462 2321 2463 2325
rect 2467 2321 2468 2325
rect 2462 2320 2468 2321
rect 2614 2325 2620 2326
rect 2614 2321 2615 2325
rect 2619 2321 2620 2325
rect 2614 2320 2620 2321
rect 2774 2325 2780 2326
rect 2774 2321 2775 2325
rect 2779 2321 2780 2325
rect 2774 2320 2780 2321
rect 2047 2319 2051 2320
rect 2403 2319 2407 2320
rect 2404 2308 2406 2319
rect 2876 2312 2878 2330
rect 2944 2326 2946 2337
rect 3112 2326 3114 2337
rect 3288 2326 3290 2337
rect 3472 2326 3474 2337
rect 2942 2325 2948 2326
rect 2942 2321 2943 2325
rect 2947 2321 2948 2325
rect 2942 2320 2948 2321
rect 3110 2325 3116 2326
rect 3110 2321 3111 2325
rect 3115 2321 3116 2325
rect 3110 2320 3116 2321
rect 3286 2325 3292 2326
rect 3286 2321 3287 2325
rect 3291 2321 3292 2325
rect 3286 2320 3292 2321
rect 3470 2325 3476 2326
rect 3470 2321 3471 2325
rect 3475 2321 3476 2325
rect 3470 2320 3476 2321
rect 3576 2313 3578 2337
rect 3574 2312 3580 2313
rect 2874 2311 2880 2312
rect 2402 2307 2408 2308
rect 2402 2303 2403 2307
rect 2407 2303 2408 2307
rect 2874 2307 2875 2311
rect 2879 2307 2880 2311
rect 3574 2308 3575 2312
rect 3579 2308 3580 2312
rect 3574 2307 3580 2308
rect 2874 2306 2880 2307
rect 2402 2302 2408 2303
rect 3574 2295 3580 2296
rect 3574 2291 3575 2295
rect 3579 2291 3580 2295
rect 3574 2290 3580 2291
rect 1998 2285 2004 2286
rect 1998 2281 1999 2285
rect 2003 2281 2004 2285
rect 1998 2280 2004 2281
rect 2150 2285 2156 2286
rect 2150 2281 2151 2285
rect 2155 2281 2156 2285
rect 2150 2280 2156 2281
rect 2302 2285 2308 2286
rect 2302 2281 2303 2285
rect 2307 2281 2308 2285
rect 2302 2280 2308 2281
rect 2454 2285 2460 2286
rect 2454 2281 2455 2285
rect 2459 2281 2460 2285
rect 2454 2280 2460 2281
rect 2606 2285 2612 2286
rect 2606 2281 2607 2285
rect 2611 2281 2612 2285
rect 2606 2280 2612 2281
rect 2766 2285 2772 2286
rect 2766 2281 2767 2285
rect 2771 2281 2772 2285
rect 2766 2280 2772 2281
rect 2934 2285 2940 2286
rect 2934 2281 2935 2285
rect 2939 2281 2940 2285
rect 2934 2280 2940 2281
rect 3102 2285 3108 2286
rect 3102 2281 3103 2285
rect 3107 2281 3108 2285
rect 3102 2280 3108 2281
rect 3278 2285 3284 2286
rect 3278 2281 3279 2285
rect 3283 2281 3284 2285
rect 3278 2280 3284 2281
rect 3462 2285 3468 2286
rect 3462 2281 3463 2285
rect 3467 2281 3468 2285
rect 3462 2280 3468 2281
rect 2000 2271 2002 2280
rect 2152 2271 2154 2280
rect 2304 2271 2306 2280
rect 2456 2271 2458 2280
rect 2608 2271 2610 2280
rect 2768 2271 2770 2280
rect 2798 2279 2804 2280
rect 2798 2275 2799 2279
rect 2803 2275 2804 2279
rect 2798 2274 2804 2275
rect 1999 2270 2003 2271
rect 1999 2265 2003 2266
rect 2023 2270 2027 2271
rect 2023 2265 2027 2266
rect 2151 2270 2155 2271
rect 2151 2265 2155 2266
rect 2199 2270 2203 2271
rect 2199 2265 2203 2266
rect 2303 2270 2307 2271
rect 2303 2265 2307 2266
rect 2383 2270 2387 2271
rect 2383 2265 2387 2266
rect 2455 2270 2459 2271
rect 2455 2265 2459 2266
rect 2567 2270 2571 2271
rect 2567 2265 2571 2266
rect 2607 2270 2611 2271
rect 2607 2265 2611 2266
rect 2743 2270 2747 2271
rect 2743 2265 2747 2266
rect 2767 2270 2771 2271
rect 2767 2265 2771 2266
rect 2024 2260 2026 2265
rect 2200 2260 2202 2265
rect 2384 2260 2386 2265
rect 2568 2260 2570 2265
rect 2744 2260 2746 2265
rect 2022 2259 2028 2260
rect 2022 2255 2023 2259
rect 2027 2255 2028 2259
rect 2022 2254 2028 2255
rect 2198 2259 2204 2260
rect 2198 2255 2199 2259
rect 2203 2255 2204 2259
rect 2198 2254 2204 2255
rect 2382 2259 2388 2260
rect 2382 2255 2383 2259
rect 2387 2255 2388 2259
rect 2382 2254 2388 2255
rect 2566 2259 2572 2260
rect 2566 2255 2567 2259
rect 2571 2255 2572 2259
rect 2566 2254 2572 2255
rect 2742 2259 2748 2260
rect 2742 2255 2743 2259
rect 2747 2255 2748 2259
rect 2742 2254 2748 2255
rect 1951 2252 1955 2253
rect 2479 2252 2483 2253
rect 1823 2249 1827 2250
rect 1862 2249 1868 2250
rect 1456 2244 1458 2249
rect 1454 2243 1460 2244
rect 1454 2239 1455 2243
rect 1459 2239 1460 2243
rect 1454 2238 1460 2239
rect 1398 2235 1404 2236
rect 1398 2231 1399 2235
rect 1403 2231 1404 2235
rect 1824 2234 1826 2249
rect 1862 2245 1863 2249
rect 1867 2245 1868 2249
rect 1951 2247 1955 2248
rect 2478 2247 2479 2252
rect 2483 2247 2484 2252
rect 2478 2246 2484 2247
rect 1862 2244 1868 2245
rect 1398 2230 1404 2231
rect 1822 2233 1828 2234
rect 1400 2197 1402 2230
rect 1822 2229 1823 2233
rect 1827 2229 1828 2233
rect 1822 2228 1828 2229
rect 1862 2232 1868 2233
rect 1862 2228 1863 2232
rect 1867 2228 1868 2232
rect 1862 2227 1868 2228
rect 1822 2216 1828 2217
rect 1822 2212 1823 2216
rect 1827 2212 1828 2216
rect 1822 2211 1828 2212
rect 1462 2203 1468 2204
rect 1462 2199 1463 2203
rect 1467 2199 1468 2203
rect 1462 2198 1468 2199
rect 1399 2196 1403 2197
rect 1318 2191 1324 2192
rect 1399 2191 1403 2192
rect 1318 2187 1319 2191
rect 1323 2187 1324 2191
rect 1318 2186 1324 2187
rect 1464 2183 1466 2198
rect 1824 2183 1826 2211
rect 1864 2199 1866 2227
rect 1894 2219 1900 2220
rect 1894 2215 1895 2219
rect 1899 2215 1900 2219
rect 1894 2214 1900 2215
rect 2030 2219 2036 2220
rect 2030 2215 2031 2219
rect 2035 2215 2036 2219
rect 2030 2214 2036 2215
rect 2206 2219 2212 2220
rect 2206 2215 2207 2219
rect 2211 2215 2212 2219
rect 2206 2214 2212 2215
rect 2390 2219 2396 2220
rect 2390 2215 2391 2219
rect 2395 2215 2396 2219
rect 2390 2214 2396 2215
rect 2574 2219 2580 2220
rect 2574 2215 2575 2219
rect 2579 2215 2580 2219
rect 2574 2214 2580 2215
rect 2750 2219 2756 2220
rect 2750 2215 2751 2219
rect 2755 2215 2756 2219
rect 2750 2214 2756 2215
rect 1896 2199 1898 2214
rect 2006 2207 2012 2208
rect 2006 2203 2007 2207
rect 2011 2203 2012 2207
rect 2006 2202 2012 2203
rect 1863 2198 1867 2199
rect 1863 2193 1867 2194
rect 1895 2198 1899 2199
rect 1895 2193 1899 2194
rect 1167 2182 1171 2183
rect 1167 2177 1171 2178
rect 1311 2182 1315 2183
rect 1311 2177 1315 2178
rect 1463 2182 1467 2183
rect 1463 2177 1467 2178
rect 1823 2182 1827 2183
rect 1823 2177 1827 2178
rect 1082 2175 1088 2176
rect 1082 2171 1083 2175
rect 1087 2171 1088 2175
rect 1082 2170 1088 2171
rect 1168 2166 1170 2177
rect 942 2165 948 2166
rect 942 2161 943 2165
rect 947 2161 948 2165
rect 942 2160 948 2161
rect 1054 2165 1060 2166
rect 1054 2161 1055 2165
rect 1059 2161 1060 2165
rect 1054 2160 1060 2161
rect 1166 2165 1172 2166
rect 1166 2161 1167 2165
rect 1171 2161 1172 2165
rect 1166 2160 1172 2161
rect 1824 2153 1826 2177
rect 1864 2169 1866 2193
rect 1896 2182 1898 2193
rect 1894 2181 1900 2182
rect 2008 2181 2010 2202
rect 2032 2199 2034 2214
rect 2208 2199 2210 2214
rect 2392 2199 2394 2214
rect 2576 2199 2578 2214
rect 2752 2199 2754 2214
rect 2771 2212 2775 2213
rect 2800 2208 2802 2274
rect 2936 2271 2938 2280
rect 3104 2271 3106 2280
rect 3280 2271 3282 2280
rect 3464 2271 3466 2280
rect 3498 2279 3504 2280
rect 3498 2275 3499 2279
rect 3503 2275 3504 2279
rect 3498 2274 3504 2275
rect 2911 2270 2915 2271
rect 2911 2265 2915 2266
rect 2935 2270 2939 2271
rect 2935 2265 2939 2266
rect 3079 2270 3083 2271
rect 3079 2265 3083 2266
rect 3103 2270 3107 2271
rect 3103 2265 3107 2266
rect 3239 2270 3243 2271
rect 3239 2265 3243 2266
rect 3279 2270 3283 2271
rect 3279 2265 3283 2266
rect 3407 2270 3411 2271
rect 3407 2265 3411 2266
rect 3463 2270 3467 2271
rect 3463 2265 3467 2266
rect 2912 2260 2914 2265
rect 3080 2260 3082 2265
rect 3240 2260 3242 2265
rect 3408 2260 3410 2265
rect 2910 2259 2916 2260
rect 2910 2255 2911 2259
rect 2915 2255 2916 2259
rect 2910 2254 2916 2255
rect 3078 2259 3084 2260
rect 3078 2255 3079 2259
rect 3083 2255 3084 2259
rect 3078 2254 3084 2255
rect 3238 2259 3244 2260
rect 3238 2255 3239 2259
rect 3243 2255 3244 2259
rect 3238 2254 3244 2255
rect 3406 2259 3412 2260
rect 3406 2255 3407 2259
rect 3411 2255 3412 2259
rect 3406 2254 3412 2255
rect 3146 2251 3152 2252
rect 3146 2247 3147 2251
rect 3151 2247 3152 2251
rect 3146 2246 3152 2247
rect 2918 2219 2924 2220
rect 2918 2215 2919 2219
rect 2923 2215 2924 2219
rect 2918 2214 2924 2215
rect 3086 2219 3092 2220
rect 3086 2215 3087 2219
rect 3091 2215 3092 2219
rect 3086 2214 3092 2215
rect 2771 2207 2775 2208
rect 2798 2207 2804 2208
rect 2031 2198 2035 2199
rect 2031 2193 2035 2194
rect 2039 2198 2043 2199
rect 2039 2193 2043 2194
rect 2207 2198 2211 2199
rect 2207 2193 2211 2194
rect 2215 2198 2219 2199
rect 2215 2193 2219 2194
rect 2391 2198 2395 2199
rect 2391 2193 2395 2194
rect 2399 2198 2403 2199
rect 2399 2193 2403 2194
rect 2575 2198 2579 2199
rect 2575 2193 2579 2194
rect 2583 2198 2587 2199
rect 2583 2193 2587 2194
rect 2751 2198 2755 2199
rect 2751 2193 2755 2194
rect 2759 2198 2763 2199
rect 2759 2193 2763 2194
rect 2040 2182 2042 2193
rect 2216 2182 2218 2193
rect 2400 2182 2402 2193
rect 2584 2182 2586 2193
rect 2760 2182 2762 2193
rect 2772 2192 2774 2207
rect 2798 2203 2799 2207
rect 2803 2203 2804 2207
rect 2798 2202 2804 2203
rect 2920 2199 2922 2214
rect 3088 2199 3090 2214
rect 3148 2213 3150 2246
rect 3246 2219 3252 2220
rect 3246 2215 3247 2219
rect 3251 2215 3252 2219
rect 3246 2214 3252 2215
rect 3414 2219 3420 2220
rect 3414 2215 3415 2219
rect 3419 2215 3420 2219
rect 3414 2214 3420 2215
rect 3147 2212 3151 2213
rect 3147 2207 3151 2208
rect 3248 2199 3250 2214
rect 3416 2199 3418 2214
rect 3426 2207 3432 2208
rect 3426 2203 3427 2207
rect 3431 2203 3432 2207
rect 3426 2202 3432 2203
rect 2919 2198 2923 2199
rect 2919 2193 2923 2194
rect 3071 2198 3075 2199
rect 3071 2193 3075 2194
rect 3087 2198 3091 2199
rect 3087 2193 3091 2194
rect 3215 2198 3219 2199
rect 3215 2193 3219 2194
rect 3247 2198 3251 2199
rect 3247 2193 3251 2194
rect 3359 2198 3363 2199
rect 3359 2193 3363 2194
rect 3415 2198 3419 2199
rect 3415 2193 3419 2194
rect 2770 2191 2776 2192
rect 2770 2187 2771 2191
rect 2775 2187 2776 2191
rect 2770 2186 2776 2187
rect 2920 2182 2922 2193
rect 3072 2182 3074 2193
rect 3216 2182 3218 2193
rect 3360 2182 3362 2193
rect 2038 2181 2044 2182
rect 1894 2177 1895 2181
rect 1899 2177 1900 2181
rect 1894 2176 1900 2177
rect 2007 2180 2011 2181
rect 2038 2177 2039 2181
rect 2043 2177 2044 2181
rect 2038 2176 2044 2177
rect 2214 2181 2220 2182
rect 2214 2177 2215 2181
rect 2219 2177 2220 2181
rect 2214 2176 2220 2177
rect 2398 2181 2404 2182
rect 2582 2181 2588 2182
rect 2398 2177 2399 2181
rect 2403 2177 2404 2181
rect 2398 2176 2404 2177
rect 2507 2180 2511 2181
rect 2582 2177 2583 2181
rect 2587 2177 2588 2181
rect 2582 2176 2588 2177
rect 2758 2181 2764 2182
rect 2758 2177 2759 2181
rect 2763 2177 2764 2181
rect 2758 2176 2764 2177
rect 2918 2181 2924 2182
rect 2918 2177 2919 2181
rect 2923 2177 2924 2181
rect 2918 2176 2924 2177
rect 3070 2181 3076 2182
rect 3070 2177 3071 2181
rect 3075 2177 3076 2181
rect 3070 2176 3076 2177
rect 3214 2181 3220 2182
rect 3214 2177 3215 2181
rect 3219 2177 3220 2181
rect 3214 2176 3220 2177
rect 3358 2181 3364 2182
rect 3358 2177 3359 2181
rect 3363 2177 3364 2181
rect 3358 2176 3364 2177
rect 2007 2175 2011 2176
rect 2507 2175 2511 2176
rect 1862 2168 1868 2169
rect 1862 2164 1863 2168
rect 1867 2164 1868 2168
rect 2508 2164 2510 2175
rect 1862 2163 1868 2164
rect 2506 2163 2512 2164
rect 2506 2159 2507 2163
rect 2511 2159 2512 2163
rect 2506 2158 2512 2159
rect 1822 2152 1828 2153
rect 1822 2148 1823 2152
rect 1827 2148 1828 2152
rect 898 2147 904 2148
rect 1822 2147 1828 2148
rect 1862 2151 1868 2152
rect 1862 2147 1863 2151
rect 1867 2147 1868 2151
rect 898 2143 899 2147
rect 903 2143 904 2147
rect 1862 2146 1868 2147
rect 3334 2151 3340 2152
rect 3334 2147 3335 2151
rect 3339 2147 3340 2151
rect 3334 2146 3340 2147
rect 898 2142 904 2143
rect 1822 2135 1828 2136
rect 1822 2131 1823 2135
rect 1827 2131 1828 2135
rect 1822 2130 1828 2131
rect 510 2125 516 2126
rect 510 2121 511 2125
rect 515 2121 516 2125
rect 510 2120 516 2121
rect 614 2125 620 2126
rect 614 2121 615 2125
rect 619 2121 620 2125
rect 614 2120 620 2121
rect 718 2125 724 2126
rect 718 2121 719 2125
rect 723 2121 724 2125
rect 718 2120 724 2121
rect 822 2125 828 2126
rect 822 2121 823 2125
rect 827 2121 828 2125
rect 822 2120 828 2121
rect 934 2125 940 2126
rect 934 2121 935 2125
rect 939 2121 940 2125
rect 934 2120 940 2121
rect 1046 2125 1052 2126
rect 1046 2121 1047 2125
rect 1051 2121 1052 2125
rect 1046 2120 1052 2121
rect 1158 2125 1164 2126
rect 1158 2121 1159 2125
rect 1163 2121 1164 2125
rect 1158 2120 1164 2121
rect 512 2107 514 2120
rect 616 2107 618 2120
rect 720 2107 722 2120
rect 824 2107 826 2120
rect 850 2119 856 2120
rect 850 2115 851 2119
rect 855 2115 856 2119
rect 850 2114 856 2115
rect 511 2106 515 2107
rect 511 2101 515 2102
rect 527 2106 531 2107
rect 527 2101 531 2102
rect 615 2106 619 2107
rect 615 2101 619 2102
rect 631 2106 635 2107
rect 631 2101 635 2102
rect 719 2106 723 2107
rect 719 2101 723 2102
rect 735 2106 739 2107
rect 735 2101 739 2102
rect 823 2106 827 2107
rect 823 2101 827 2102
rect 831 2106 835 2107
rect 831 2101 835 2102
rect 528 2096 530 2101
rect 632 2096 634 2101
rect 736 2096 738 2101
rect 832 2096 834 2101
rect 526 2095 532 2096
rect 526 2091 527 2095
rect 531 2091 532 2095
rect 526 2090 532 2091
rect 630 2095 636 2096
rect 630 2091 631 2095
rect 635 2091 636 2095
rect 630 2090 636 2091
rect 734 2095 740 2096
rect 734 2091 735 2095
rect 739 2091 740 2095
rect 734 2090 740 2091
rect 830 2095 836 2096
rect 830 2091 831 2095
rect 835 2091 836 2095
rect 830 2090 836 2091
rect 490 2087 496 2088
rect 490 2083 491 2087
rect 495 2083 496 2087
rect 490 2082 496 2083
rect 430 2055 436 2056
rect 430 2051 431 2055
rect 435 2051 436 2055
rect 430 2050 436 2051
rect 534 2055 540 2056
rect 534 2051 535 2055
rect 539 2051 540 2055
rect 534 2050 540 2051
rect 638 2055 644 2056
rect 638 2051 639 2055
rect 643 2051 644 2055
rect 638 2050 644 2051
rect 742 2055 748 2056
rect 742 2051 743 2055
rect 747 2051 748 2055
rect 742 2050 748 2051
rect 838 2055 844 2056
rect 838 2051 839 2055
rect 843 2051 844 2055
rect 838 2050 844 2051
rect 338 2043 344 2044
rect 338 2039 339 2043
rect 343 2039 344 2043
rect 338 2038 344 2039
rect 432 2031 434 2050
rect 536 2031 538 2050
rect 640 2031 642 2050
rect 744 2031 746 2050
rect 790 2043 796 2044
rect 790 2039 791 2043
rect 795 2039 796 2043
rect 790 2038 796 2039
rect 111 2030 115 2031
rect 111 2025 115 2026
rect 215 2030 219 2031
rect 215 2025 219 2026
rect 327 2030 331 2031
rect 327 2025 331 2026
rect 391 2030 395 2031
rect 391 2025 395 2026
rect 431 2030 435 2031
rect 431 2025 435 2026
rect 535 2030 539 2031
rect 535 2025 539 2026
rect 559 2030 563 2031
rect 559 2025 563 2026
rect 639 2030 643 2031
rect 639 2025 643 2026
rect 719 2030 723 2031
rect 719 2025 723 2026
rect 743 2030 747 2031
rect 743 2025 747 2026
rect 112 2001 114 2025
rect 216 2014 218 2025
rect 392 2014 394 2025
rect 560 2014 562 2025
rect 614 2023 620 2024
rect 614 2019 615 2023
rect 619 2019 620 2023
rect 614 2018 620 2019
rect 650 2023 656 2024
rect 650 2019 651 2023
rect 655 2019 656 2023
rect 650 2018 656 2019
rect 214 2013 220 2014
rect 214 2009 215 2013
rect 219 2009 220 2013
rect 214 2008 220 2009
rect 390 2013 396 2014
rect 390 2009 391 2013
rect 395 2009 396 2013
rect 390 2008 396 2009
rect 558 2013 564 2014
rect 558 2009 559 2013
rect 563 2009 564 2013
rect 558 2008 564 2009
rect 110 2000 116 2001
rect 110 1996 111 2000
rect 115 1996 116 2000
rect 110 1995 116 1996
rect 110 1983 116 1984
rect 110 1979 111 1983
rect 115 1979 116 1983
rect 110 1978 116 1979
rect 154 1983 160 1984
rect 154 1979 155 1983
rect 159 1979 160 1983
rect 154 1978 160 1979
rect 112 1955 114 1978
rect 111 1954 115 1955
rect 111 1949 115 1950
rect 135 1954 139 1955
rect 135 1949 139 1950
rect 112 1934 114 1949
rect 136 1944 138 1949
rect 134 1943 140 1944
rect 134 1939 135 1943
rect 139 1939 140 1943
rect 134 1938 140 1939
rect 110 1933 116 1934
rect 110 1929 111 1933
rect 115 1929 116 1933
rect 110 1928 116 1929
rect 110 1916 116 1917
rect 110 1912 111 1916
rect 115 1912 116 1916
rect 110 1911 116 1912
rect 112 1879 114 1911
rect 142 1903 148 1904
rect 142 1899 143 1903
rect 147 1899 148 1903
rect 142 1898 148 1899
rect 144 1879 146 1898
rect 156 1892 158 1978
rect 206 1973 212 1974
rect 206 1969 207 1973
rect 211 1969 212 1973
rect 206 1968 212 1969
rect 382 1973 388 1974
rect 382 1969 383 1973
rect 387 1969 388 1973
rect 382 1968 388 1969
rect 550 1973 556 1974
rect 550 1969 551 1973
rect 555 1969 556 1973
rect 550 1968 556 1969
rect 208 1955 210 1968
rect 384 1955 386 1968
rect 552 1955 554 1968
rect 207 1954 211 1955
rect 207 1949 211 1950
rect 311 1954 315 1955
rect 311 1949 315 1950
rect 383 1954 387 1955
rect 383 1949 387 1950
rect 519 1954 523 1955
rect 519 1949 523 1950
rect 551 1954 555 1955
rect 551 1949 555 1950
rect 312 1944 314 1949
rect 520 1944 522 1949
rect 310 1943 316 1944
rect 310 1939 311 1943
rect 315 1939 316 1943
rect 310 1938 316 1939
rect 518 1943 524 1944
rect 518 1939 519 1943
rect 523 1939 524 1943
rect 518 1938 524 1939
rect 616 1936 618 2018
rect 652 2000 654 2018
rect 720 2014 722 2025
rect 782 2023 788 2024
rect 782 2019 783 2023
rect 787 2019 788 2023
rect 782 2018 788 2019
rect 718 2013 724 2014
rect 718 2009 719 2013
rect 723 2009 724 2013
rect 718 2008 724 2009
rect 784 2000 786 2018
rect 650 1999 656 2000
rect 650 1995 651 1999
rect 655 1995 656 1999
rect 650 1994 656 1995
rect 782 1999 788 2000
rect 782 1995 783 1999
rect 787 1995 788 1999
rect 792 1996 794 2038
rect 840 2031 842 2050
rect 852 2044 854 2114
rect 936 2107 938 2120
rect 1048 2107 1050 2120
rect 1160 2107 1162 2120
rect 1824 2107 1826 2130
rect 1864 2127 1866 2146
rect 1886 2141 1892 2142
rect 1886 2137 1887 2141
rect 1891 2137 1892 2141
rect 1886 2136 1892 2137
rect 2030 2141 2036 2142
rect 2030 2137 2031 2141
rect 2035 2137 2036 2141
rect 2030 2136 2036 2137
rect 2206 2141 2212 2142
rect 2206 2137 2207 2141
rect 2211 2137 2212 2141
rect 2206 2136 2212 2137
rect 2390 2141 2396 2142
rect 2390 2137 2391 2141
rect 2395 2137 2396 2141
rect 2390 2136 2396 2137
rect 2574 2141 2580 2142
rect 2574 2137 2575 2141
rect 2579 2137 2580 2141
rect 2574 2136 2580 2137
rect 2750 2141 2756 2142
rect 2750 2137 2751 2141
rect 2755 2137 2756 2141
rect 2750 2136 2756 2137
rect 2910 2141 2916 2142
rect 2910 2137 2911 2141
rect 2915 2137 2916 2141
rect 2910 2136 2916 2137
rect 3062 2141 3068 2142
rect 3062 2137 3063 2141
rect 3067 2137 3068 2141
rect 3062 2136 3068 2137
rect 3206 2141 3212 2142
rect 3206 2137 3207 2141
rect 3211 2137 3212 2141
rect 3206 2136 3212 2137
rect 1888 2127 1890 2136
rect 2032 2127 2034 2136
rect 2208 2127 2210 2136
rect 2392 2127 2394 2136
rect 2576 2127 2578 2136
rect 2752 2127 2754 2136
rect 2912 2127 2914 2136
rect 3064 2127 3066 2136
rect 3208 2127 3210 2136
rect 1863 2126 1867 2127
rect 1863 2121 1867 2122
rect 1887 2126 1891 2127
rect 1887 2121 1891 2122
rect 2023 2126 2027 2127
rect 2023 2121 2027 2122
rect 2031 2126 2035 2127
rect 2031 2121 2035 2122
rect 2199 2126 2203 2127
rect 2199 2121 2203 2122
rect 2207 2126 2211 2127
rect 2207 2121 2211 2122
rect 2375 2126 2379 2127
rect 2375 2121 2379 2122
rect 2391 2126 2395 2127
rect 2391 2121 2395 2122
rect 2551 2126 2555 2127
rect 2551 2121 2555 2122
rect 2575 2126 2579 2127
rect 2575 2121 2579 2122
rect 2719 2126 2723 2127
rect 2719 2121 2723 2122
rect 2751 2126 2755 2127
rect 2751 2121 2755 2122
rect 2879 2126 2883 2127
rect 2879 2121 2883 2122
rect 2911 2126 2915 2127
rect 2911 2121 2915 2122
rect 3031 2126 3035 2127
rect 3031 2121 3035 2122
rect 3063 2126 3067 2127
rect 3063 2121 3067 2122
rect 3175 2126 3179 2127
rect 3175 2121 3179 2122
rect 3207 2126 3211 2127
rect 3207 2121 3211 2122
rect 3319 2126 3323 2127
rect 3319 2121 3323 2122
rect 927 2106 931 2107
rect 927 2101 931 2102
rect 935 2106 939 2107
rect 935 2101 939 2102
rect 1031 2106 1035 2107
rect 1031 2101 1035 2102
rect 1047 2106 1051 2107
rect 1047 2101 1051 2102
rect 1135 2106 1139 2107
rect 1135 2101 1139 2102
rect 1159 2106 1163 2107
rect 1159 2101 1163 2102
rect 1239 2106 1243 2107
rect 1239 2101 1243 2102
rect 1823 2106 1827 2107
rect 1864 2106 1866 2121
rect 1888 2116 1890 2121
rect 2024 2116 2026 2121
rect 2200 2116 2202 2121
rect 2376 2116 2378 2121
rect 2552 2116 2554 2121
rect 2720 2116 2722 2121
rect 2880 2116 2882 2121
rect 3032 2116 3034 2121
rect 3176 2116 3178 2121
rect 3320 2116 3322 2121
rect 1886 2115 1892 2116
rect 1886 2111 1887 2115
rect 1891 2111 1892 2115
rect 1886 2110 1892 2111
rect 2022 2115 2028 2116
rect 2022 2111 2023 2115
rect 2027 2111 2028 2115
rect 2022 2110 2028 2111
rect 2198 2115 2204 2116
rect 2198 2111 2199 2115
rect 2203 2111 2204 2115
rect 2198 2110 2204 2111
rect 2374 2115 2380 2116
rect 2374 2111 2375 2115
rect 2379 2111 2380 2115
rect 2374 2110 2380 2111
rect 2550 2115 2556 2116
rect 2550 2111 2551 2115
rect 2555 2111 2556 2115
rect 2550 2110 2556 2111
rect 2718 2115 2724 2116
rect 2718 2111 2719 2115
rect 2723 2111 2724 2115
rect 2718 2110 2724 2111
rect 2878 2115 2884 2116
rect 2878 2111 2879 2115
rect 2883 2111 2884 2115
rect 2878 2110 2884 2111
rect 3030 2115 3036 2116
rect 3030 2111 3031 2115
rect 3035 2111 3036 2115
rect 3030 2110 3036 2111
rect 3174 2115 3180 2116
rect 3174 2111 3175 2115
rect 3179 2111 3180 2115
rect 3174 2110 3180 2111
rect 3318 2115 3324 2116
rect 3318 2111 3319 2115
rect 3323 2111 3324 2115
rect 3318 2110 3324 2111
rect 2478 2107 2484 2108
rect 1823 2101 1827 2102
rect 1862 2105 1868 2106
rect 1862 2101 1863 2105
rect 1867 2101 1868 2105
rect 2478 2103 2479 2107
rect 2483 2103 2484 2107
rect 2478 2102 2484 2103
rect 928 2096 930 2101
rect 1032 2096 1034 2101
rect 1136 2096 1138 2101
rect 1240 2096 1242 2101
rect 926 2095 932 2096
rect 926 2091 927 2095
rect 931 2091 932 2095
rect 926 2090 932 2091
rect 1030 2095 1036 2096
rect 1030 2091 1031 2095
rect 1035 2091 1036 2095
rect 1030 2090 1036 2091
rect 1134 2095 1140 2096
rect 1134 2091 1135 2095
rect 1139 2091 1140 2095
rect 1134 2090 1140 2091
rect 1238 2095 1244 2096
rect 1238 2091 1239 2095
rect 1243 2091 1244 2095
rect 1238 2090 1244 2091
rect 1824 2086 1826 2101
rect 1862 2100 1868 2101
rect 1954 2091 1960 2092
rect 1862 2088 1868 2089
rect 1822 2085 1828 2086
rect 1822 2081 1823 2085
rect 1827 2081 1828 2085
rect 1862 2084 1863 2088
rect 1867 2084 1868 2088
rect 1954 2087 1955 2091
rect 1959 2087 1960 2091
rect 1954 2086 1960 2087
rect 1862 2083 1868 2084
rect 1822 2080 1828 2081
rect 1206 2071 1212 2072
rect 1206 2067 1207 2071
rect 1211 2067 1212 2071
rect 1206 2066 1212 2067
rect 1214 2071 1220 2072
rect 1214 2067 1215 2071
rect 1219 2067 1220 2071
rect 1214 2066 1220 2067
rect 1822 2068 1828 2069
rect 934 2055 940 2056
rect 934 2051 935 2055
rect 939 2051 940 2055
rect 934 2050 940 2051
rect 1038 2055 1044 2056
rect 1038 2051 1039 2055
rect 1043 2051 1044 2055
rect 1038 2050 1044 2051
rect 1142 2055 1148 2056
rect 1142 2051 1143 2055
rect 1147 2051 1148 2055
rect 1142 2050 1148 2051
rect 850 2043 856 2044
rect 850 2039 851 2043
rect 855 2039 856 2043
rect 850 2038 856 2039
rect 936 2031 938 2050
rect 1040 2031 1042 2050
rect 1144 2031 1146 2050
rect 1208 2044 1210 2066
rect 1206 2043 1212 2044
rect 1206 2039 1207 2043
rect 1211 2039 1212 2043
rect 1206 2038 1212 2039
rect 1216 2032 1218 2066
rect 1822 2064 1823 2068
rect 1827 2064 1828 2068
rect 1822 2063 1828 2064
rect 1246 2055 1252 2056
rect 1246 2051 1247 2055
rect 1251 2051 1252 2055
rect 1246 2050 1252 2051
rect 1214 2031 1220 2032
rect 1248 2031 1250 2050
rect 1824 2031 1826 2063
rect 1864 2051 1866 2083
rect 1894 2075 1900 2076
rect 1894 2071 1895 2075
rect 1899 2071 1900 2075
rect 1894 2070 1900 2071
rect 1896 2051 1898 2070
rect 1956 2064 1958 2086
rect 2030 2075 2036 2076
rect 2030 2071 2031 2075
rect 2035 2071 2036 2075
rect 2030 2070 2036 2071
rect 2206 2075 2212 2076
rect 2206 2071 2207 2075
rect 2211 2071 2212 2075
rect 2206 2070 2212 2071
rect 2382 2075 2388 2076
rect 2382 2071 2383 2075
rect 2387 2071 2388 2075
rect 2382 2070 2388 2071
rect 1954 2063 1960 2064
rect 1954 2059 1955 2063
rect 1959 2059 1960 2063
rect 1954 2058 1960 2059
rect 2032 2051 2034 2070
rect 2039 2068 2043 2069
rect 2038 2063 2044 2064
rect 2038 2059 2039 2063
rect 2043 2059 2044 2063
rect 2038 2058 2044 2059
rect 2208 2051 2210 2070
rect 2214 2063 2220 2064
rect 2214 2059 2215 2063
rect 2219 2059 2220 2063
rect 2214 2058 2220 2059
rect 1863 2050 1867 2051
rect 1863 2045 1867 2046
rect 1895 2050 1899 2051
rect 1895 2045 1899 2046
rect 2015 2050 2019 2051
rect 2015 2045 2019 2046
rect 2031 2050 2035 2051
rect 2031 2045 2035 2046
rect 2151 2050 2155 2051
rect 2151 2045 2155 2046
rect 2207 2050 2211 2051
rect 2207 2045 2211 2046
rect 839 2030 843 2031
rect 839 2025 843 2026
rect 863 2030 867 2031
rect 863 2025 867 2026
rect 935 2030 939 2031
rect 935 2025 939 2026
rect 999 2030 1003 2031
rect 999 2025 1003 2026
rect 1039 2030 1043 2031
rect 1039 2025 1043 2026
rect 1127 2030 1131 2031
rect 1127 2025 1131 2026
rect 1143 2030 1147 2031
rect 1214 2027 1215 2031
rect 1219 2027 1220 2031
rect 1214 2026 1220 2027
rect 1247 2030 1251 2031
rect 1143 2025 1147 2026
rect 1247 2025 1251 2026
rect 1367 2030 1371 2031
rect 1367 2025 1371 2026
rect 1495 2030 1499 2031
rect 1495 2025 1499 2026
rect 1823 2030 1827 2031
rect 1823 2025 1827 2026
rect 864 2014 866 2025
rect 1000 2014 1002 2025
rect 1074 2023 1080 2024
rect 1074 2019 1075 2023
rect 1079 2019 1080 2023
rect 1074 2018 1080 2019
rect 862 2013 868 2014
rect 862 2009 863 2013
rect 867 2009 868 2013
rect 862 2008 868 2009
rect 998 2013 1004 2014
rect 998 2009 999 2013
rect 1003 2009 1004 2013
rect 998 2008 1004 2009
rect 1076 2000 1078 2018
rect 1128 2014 1130 2025
rect 1248 2014 1250 2025
rect 1318 2023 1324 2024
rect 1318 2019 1319 2023
rect 1323 2019 1324 2023
rect 1318 2018 1324 2019
rect 1126 2013 1132 2014
rect 1126 2009 1127 2013
rect 1131 2009 1132 2013
rect 1126 2008 1132 2009
rect 1246 2013 1252 2014
rect 1246 2009 1247 2013
rect 1251 2009 1252 2013
rect 1246 2008 1252 2009
rect 1320 2000 1322 2018
rect 1368 2014 1370 2025
rect 1442 2023 1448 2024
rect 1442 2019 1443 2023
rect 1447 2019 1448 2023
rect 1442 2018 1448 2019
rect 1366 2013 1372 2014
rect 1366 2009 1367 2013
rect 1371 2009 1372 2013
rect 1366 2008 1372 2009
rect 1444 2000 1446 2018
rect 1496 2014 1498 2025
rect 1494 2013 1500 2014
rect 1494 2009 1495 2013
rect 1499 2009 1500 2013
rect 1494 2008 1500 2009
rect 1824 2001 1826 2025
rect 1864 2021 1866 2045
rect 1896 2034 1898 2045
rect 1958 2043 1964 2044
rect 1958 2039 1959 2043
rect 1963 2039 1964 2043
rect 1958 2038 1964 2039
rect 1894 2033 1900 2034
rect 1894 2029 1895 2033
rect 1899 2029 1900 2033
rect 1894 2028 1900 2029
rect 1862 2020 1868 2021
rect 1960 2020 1962 2038
rect 2016 2034 2018 2045
rect 2090 2043 2096 2044
rect 2090 2039 2091 2043
rect 2095 2039 2096 2043
rect 2090 2038 2096 2039
rect 2014 2033 2020 2034
rect 2006 2031 2012 2032
rect 2006 2026 2007 2031
rect 2011 2026 2012 2031
rect 2014 2029 2015 2033
rect 2019 2029 2020 2033
rect 2014 2028 2020 2029
rect 2007 2023 2011 2024
rect 2092 2020 2094 2038
rect 2152 2034 2154 2045
rect 2150 2033 2156 2034
rect 2150 2029 2151 2033
rect 2155 2029 2156 2033
rect 2150 2028 2156 2029
rect 2216 2020 2218 2058
rect 2384 2051 2386 2070
rect 2480 2069 2482 2102
rect 2618 2091 2624 2092
rect 2618 2087 2619 2091
rect 2623 2087 2624 2091
rect 2618 2086 2624 2087
rect 2790 2091 2796 2092
rect 2790 2087 2791 2091
rect 2795 2087 2796 2091
rect 2790 2086 2796 2087
rect 2946 2091 2952 2092
rect 2946 2087 2947 2091
rect 2951 2087 2952 2091
rect 2946 2086 2952 2087
rect 3098 2091 3104 2092
rect 3098 2087 3099 2091
rect 3103 2087 3104 2091
rect 3098 2086 3104 2087
rect 3242 2091 3248 2092
rect 3242 2087 3243 2091
rect 3247 2087 3248 2091
rect 3242 2086 3248 2087
rect 2558 2075 2564 2076
rect 2558 2071 2559 2075
rect 2563 2071 2564 2075
rect 2558 2070 2564 2071
rect 2479 2068 2483 2069
rect 2479 2063 2483 2064
rect 2560 2051 2562 2070
rect 2295 2050 2299 2051
rect 2295 2045 2299 2046
rect 2383 2050 2387 2051
rect 2383 2045 2387 2046
rect 2439 2050 2443 2051
rect 2439 2045 2443 2046
rect 2559 2050 2563 2051
rect 2559 2045 2563 2046
rect 2591 2050 2595 2051
rect 2591 2045 2595 2046
rect 2296 2034 2298 2045
rect 2362 2043 2368 2044
rect 2362 2039 2363 2043
rect 2367 2039 2368 2043
rect 2362 2038 2368 2039
rect 2294 2033 2300 2034
rect 2294 2029 2295 2033
rect 2299 2029 2300 2033
rect 2223 2028 2227 2029
rect 2294 2028 2300 2029
rect 2223 2023 2227 2024
rect 1862 2016 1863 2020
rect 1867 2016 1868 2020
rect 1862 2015 1868 2016
rect 1958 2019 1964 2020
rect 1958 2015 1959 2019
rect 1963 2015 1964 2019
rect 1958 2014 1964 2015
rect 2090 2019 2096 2020
rect 2090 2015 2091 2019
rect 2095 2015 2096 2019
rect 2090 2014 2096 2015
rect 2214 2019 2220 2020
rect 2214 2015 2215 2019
rect 2219 2015 2220 2019
rect 2224 2016 2226 2023
rect 2364 2016 2366 2038
rect 2440 2034 2442 2045
rect 2450 2043 2456 2044
rect 2450 2039 2451 2043
rect 2455 2039 2456 2043
rect 2450 2038 2456 2039
rect 2438 2033 2444 2034
rect 2438 2029 2439 2033
rect 2443 2029 2444 2033
rect 2438 2028 2444 2029
rect 2214 2014 2220 2015
rect 2222 2015 2228 2016
rect 2222 2011 2223 2015
rect 2227 2011 2228 2015
rect 2222 2010 2228 2011
rect 2362 2015 2368 2016
rect 2362 2011 2363 2015
rect 2367 2011 2368 2015
rect 2362 2010 2368 2011
rect 1862 2003 1868 2004
rect 1822 2000 1828 2001
rect 1074 1999 1080 2000
rect 782 1994 788 1995
rect 790 1995 796 1996
rect 790 1991 791 1995
rect 795 1991 796 1995
rect 1074 1995 1075 1999
rect 1079 1995 1080 1999
rect 1074 1994 1080 1995
rect 1318 1999 1324 2000
rect 1318 1995 1319 1999
rect 1323 1995 1324 1999
rect 1318 1994 1324 1995
rect 1442 1999 1448 2000
rect 1442 1995 1443 1999
rect 1447 1995 1448 1999
rect 1822 1996 1823 2000
rect 1827 1996 1828 2000
rect 1862 1999 1863 2003
rect 1867 1999 1868 2003
rect 1862 1998 1868 1999
rect 1822 1995 1828 1996
rect 1442 1994 1448 1995
rect 790 1990 796 1991
rect 1822 1983 1828 1984
rect 1822 1979 1823 1983
rect 1827 1979 1828 1983
rect 1864 1979 1866 1998
rect 1886 1993 1892 1994
rect 1886 1989 1887 1993
rect 1891 1989 1892 1993
rect 1886 1988 1892 1989
rect 2006 1993 2012 1994
rect 2006 1989 2007 1993
rect 2011 1989 2012 1993
rect 2006 1988 2012 1989
rect 2142 1993 2148 1994
rect 2142 1989 2143 1993
rect 2147 1989 2148 1993
rect 2142 1988 2148 1989
rect 2286 1993 2292 1994
rect 2286 1989 2287 1993
rect 2291 1989 2292 1993
rect 2286 1988 2292 1989
rect 2430 1993 2436 1994
rect 2430 1989 2431 1993
rect 2435 1989 2436 1993
rect 2430 1988 2436 1989
rect 1888 1979 1890 1988
rect 2008 1979 2010 1988
rect 2144 1979 2146 1988
rect 2288 1979 2290 1988
rect 2432 1979 2434 1988
rect 1822 1978 1828 1979
rect 1863 1978 1867 1979
rect 710 1973 716 1974
rect 710 1969 711 1973
rect 715 1969 716 1973
rect 710 1968 716 1969
rect 854 1973 860 1974
rect 854 1969 855 1973
rect 859 1969 860 1973
rect 854 1968 860 1969
rect 990 1973 996 1974
rect 990 1969 991 1973
rect 995 1969 996 1973
rect 990 1968 996 1969
rect 1118 1973 1124 1974
rect 1118 1969 1119 1973
rect 1123 1969 1124 1973
rect 1118 1968 1124 1969
rect 1238 1973 1244 1974
rect 1238 1969 1239 1973
rect 1243 1969 1244 1973
rect 1238 1968 1244 1969
rect 1358 1973 1364 1974
rect 1358 1969 1359 1973
rect 1363 1969 1364 1973
rect 1358 1968 1364 1969
rect 1486 1973 1492 1974
rect 1486 1969 1487 1973
rect 1491 1969 1492 1973
rect 1486 1968 1492 1969
rect 712 1955 714 1968
rect 856 1955 858 1968
rect 992 1955 994 1968
rect 1120 1955 1122 1968
rect 1134 1967 1140 1968
rect 1134 1963 1135 1967
rect 1139 1963 1140 1967
rect 1134 1962 1140 1963
rect 711 1954 715 1955
rect 711 1949 715 1950
rect 719 1954 723 1955
rect 719 1949 723 1950
rect 855 1954 859 1955
rect 855 1949 859 1950
rect 911 1954 915 1955
rect 911 1949 915 1950
rect 991 1954 995 1955
rect 991 1949 995 1950
rect 1095 1954 1099 1955
rect 1095 1949 1099 1950
rect 1119 1954 1123 1955
rect 1119 1949 1123 1950
rect 720 1944 722 1949
rect 912 1944 914 1949
rect 1096 1944 1098 1949
rect 718 1943 724 1944
rect 718 1939 719 1943
rect 723 1939 724 1943
rect 718 1938 724 1939
rect 910 1943 916 1944
rect 910 1939 911 1943
rect 915 1939 916 1943
rect 910 1938 916 1939
rect 1094 1943 1100 1944
rect 1094 1939 1095 1943
rect 1099 1939 1100 1943
rect 1094 1938 1100 1939
rect 378 1935 384 1936
rect 378 1931 379 1935
rect 383 1931 384 1935
rect 378 1930 384 1931
rect 614 1935 620 1936
rect 614 1931 615 1935
rect 619 1931 620 1935
rect 614 1930 620 1931
rect 242 1919 248 1920
rect 242 1915 243 1919
rect 247 1915 248 1919
rect 242 1914 248 1915
rect 244 1892 246 1914
rect 318 1903 324 1904
rect 318 1899 319 1903
rect 323 1899 324 1903
rect 318 1898 324 1899
rect 154 1891 160 1892
rect 154 1887 155 1891
rect 159 1887 160 1891
rect 154 1886 160 1887
rect 242 1891 248 1892
rect 242 1887 243 1891
rect 247 1887 248 1891
rect 242 1886 248 1887
rect 320 1879 322 1898
rect 111 1878 115 1879
rect 111 1873 115 1874
rect 143 1878 147 1879
rect 143 1873 147 1874
rect 311 1878 315 1879
rect 311 1873 315 1874
rect 319 1878 323 1879
rect 319 1873 323 1874
rect 112 1849 114 1873
rect 144 1862 146 1873
rect 234 1871 240 1872
rect 234 1867 235 1871
rect 239 1867 240 1871
rect 234 1866 240 1867
rect 142 1861 148 1862
rect 142 1857 143 1861
rect 147 1857 148 1861
rect 142 1856 148 1857
rect 110 1848 116 1849
rect 110 1844 111 1848
rect 115 1844 116 1848
rect 236 1844 238 1866
rect 312 1862 314 1873
rect 380 1872 382 1930
rect 786 1919 792 1920
rect 786 1915 787 1919
rect 791 1915 792 1919
rect 786 1914 792 1915
rect 526 1903 532 1904
rect 526 1899 527 1903
rect 531 1899 532 1903
rect 526 1898 532 1899
rect 726 1903 732 1904
rect 726 1899 727 1903
rect 731 1899 732 1903
rect 726 1898 732 1899
rect 528 1879 530 1898
rect 728 1879 730 1898
rect 788 1892 790 1914
rect 918 1903 924 1904
rect 918 1899 919 1903
rect 923 1899 924 1903
rect 918 1898 924 1899
rect 1102 1903 1108 1904
rect 1102 1899 1103 1903
rect 1107 1899 1108 1903
rect 1102 1898 1108 1899
rect 786 1891 792 1892
rect 786 1887 787 1891
rect 791 1887 792 1891
rect 786 1886 792 1887
rect 920 1879 922 1898
rect 946 1891 952 1892
rect 946 1887 947 1891
rect 951 1887 952 1891
rect 946 1886 952 1887
rect 511 1878 515 1879
rect 511 1873 515 1874
rect 527 1878 531 1879
rect 527 1873 531 1874
rect 703 1878 707 1879
rect 703 1873 707 1874
rect 727 1878 731 1879
rect 727 1873 731 1874
rect 887 1878 891 1879
rect 887 1873 891 1874
rect 919 1878 923 1879
rect 919 1873 923 1874
rect 378 1871 384 1872
rect 378 1867 379 1871
rect 383 1867 384 1871
rect 378 1866 384 1867
rect 512 1862 514 1873
rect 634 1863 640 1864
rect 310 1861 316 1862
rect 310 1857 311 1861
rect 315 1857 316 1861
rect 310 1856 316 1857
rect 510 1861 516 1862
rect 510 1857 511 1861
rect 515 1857 516 1861
rect 634 1859 635 1863
rect 639 1859 640 1863
rect 704 1862 706 1873
rect 888 1862 890 1873
rect 634 1858 640 1859
rect 702 1861 708 1862
rect 510 1856 516 1857
rect 110 1843 116 1844
rect 234 1843 240 1844
rect 234 1839 235 1843
rect 239 1839 240 1843
rect 234 1838 240 1839
rect 110 1831 116 1832
rect 110 1827 111 1831
rect 115 1827 116 1831
rect 110 1826 116 1827
rect 112 1803 114 1826
rect 134 1821 140 1822
rect 134 1817 135 1821
rect 139 1817 140 1821
rect 134 1816 140 1817
rect 302 1821 308 1822
rect 302 1817 303 1821
rect 307 1817 308 1821
rect 302 1816 308 1817
rect 502 1821 508 1822
rect 502 1817 503 1821
rect 507 1817 508 1821
rect 502 1816 508 1817
rect 136 1803 138 1816
rect 154 1815 160 1816
rect 154 1811 155 1815
rect 159 1811 160 1815
rect 154 1810 160 1811
rect 111 1802 115 1803
rect 111 1797 115 1798
rect 135 1802 139 1803
rect 135 1797 139 1798
rect 112 1782 114 1797
rect 136 1792 138 1797
rect 134 1791 140 1792
rect 134 1787 135 1791
rect 139 1787 140 1791
rect 134 1786 140 1787
rect 110 1781 116 1782
rect 110 1777 111 1781
rect 115 1777 116 1781
rect 110 1776 116 1777
rect 110 1764 116 1765
rect 110 1760 111 1764
rect 115 1760 116 1764
rect 110 1759 116 1760
rect 112 1735 114 1759
rect 142 1751 148 1752
rect 142 1747 143 1751
rect 147 1747 148 1751
rect 142 1746 148 1747
rect 144 1735 146 1746
rect 156 1740 158 1810
rect 304 1803 306 1816
rect 504 1803 506 1816
rect 263 1802 267 1803
rect 263 1797 267 1798
rect 303 1802 307 1803
rect 303 1797 307 1798
rect 415 1802 419 1803
rect 415 1797 419 1798
rect 503 1802 507 1803
rect 503 1797 507 1798
rect 567 1802 571 1803
rect 567 1797 571 1798
rect 264 1792 266 1797
rect 416 1792 418 1797
rect 568 1792 570 1797
rect 262 1791 268 1792
rect 262 1787 263 1791
rect 267 1787 268 1791
rect 262 1786 268 1787
rect 414 1791 420 1792
rect 414 1787 415 1791
rect 419 1787 420 1791
rect 414 1786 420 1787
rect 566 1791 572 1792
rect 566 1787 567 1791
rect 571 1787 572 1791
rect 566 1786 572 1787
rect 636 1784 638 1858
rect 702 1857 703 1861
rect 707 1857 708 1861
rect 702 1856 708 1857
rect 886 1861 892 1862
rect 886 1857 887 1861
rect 891 1857 892 1861
rect 886 1856 892 1857
rect 948 1848 950 1886
rect 1104 1879 1106 1898
rect 1136 1892 1138 1962
rect 1240 1955 1242 1968
rect 1360 1955 1362 1968
rect 1488 1955 1490 1968
rect 1824 1955 1826 1978
rect 1863 1973 1867 1974
rect 1887 1978 1891 1979
rect 1887 1973 1891 1974
rect 2007 1978 2011 1979
rect 2007 1973 2011 1974
rect 2023 1978 2027 1979
rect 2023 1973 2027 1974
rect 2111 1978 2115 1979
rect 2111 1973 2115 1974
rect 2143 1978 2147 1979
rect 2143 1973 2147 1974
rect 2199 1978 2203 1979
rect 2199 1973 2203 1974
rect 2287 1978 2291 1979
rect 2287 1973 2291 1974
rect 2383 1978 2387 1979
rect 2383 1973 2387 1974
rect 2431 1978 2435 1979
rect 2431 1973 2435 1974
rect 1864 1958 1866 1973
rect 2024 1968 2026 1973
rect 2112 1968 2114 1973
rect 2200 1968 2202 1973
rect 2288 1968 2290 1973
rect 2384 1968 2386 1973
rect 2022 1967 2028 1968
rect 2022 1963 2023 1967
rect 2027 1963 2028 1967
rect 2022 1962 2028 1963
rect 2110 1967 2116 1968
rect 2110 1963 2111 1967
rect 2115 1963 2116 1967
rect 2110 1962 2116 1963
rect 2198 1967 2204 1968
rect 2198 1963 2199 1967
rect 2203 1963 2204 1967
rect 2198 1962 2204 1963
rect 2286 1967 2292 1968
rect 2286 1963 2287 1967
rect 2291 1963 2292 1967
rect 2286 1962 2292 1963
rect 2382 1967 2388 1968
rect 2382 1963 2383 1967
rect 2387 1963 2388 1967
rect 2382 1962 2388 1963
rect 2452 1960 2454 2038
rect 2592 2034 2594 2045
rect 2620 2044 2622 2086
rect 2726 2075 2732 2076
rect 2726 2071 2727 2075
rect 2731 2071 2732 2075
rect 2726 2070 2732 2071
rect 2728 2051 2730 2070
rect 2792 2064 2794 2086
rect 2886 2075 2892 2076
rect 2886 2071 2887 2075
rect 2891 2071 2892 2075
rect 2886 2070 2892 2071
rect 2790 2063 2796 2064
rect 2790 2059 2791 2063
rect 2795 2059 2796 2063
rect 2790 2058 2796 2059
rect 2888 2051 2890 2070
rect 2948 2064 2950 2086
rect 3038 2075 3044 2076
rect 3038 2071 3039 2075
rect 3043 2071 3044 2075
rect 3038 2070 3044 2071
rect 2946 2063 2952 2064
rect 2946 2059 2947 2063
rect 2951 2059 2952 2063
rect 2946 2058 2952 2059
rect 3040 2051 3042 2070
rect 3100 2064 3102 2086
rect 3182 2075 3188 2076
rect 3182 2071 3183 2075
rect 3187 2071 3188 2075
rect 3182 2070 3188 2071
rect 3098 2063 3104 2064
rect 3098 2059 3099 2063
rect 3103 2059 3104 2063
rect 3098 2058 3104 2059
rect 3184 2051 3186 2070
rect 3244 2064 3246 2086
rect 3326 2075 3332 2076
rect 3326 2071 3327 2075
rect 3331 2071 3332 2075
rect 3326 2070 3332 2071
rect 3242 2063 3248 2064
rect 3242 2059 3243 2063
rect 3247 2059 3248 2063
rect 3242 2058 3248 2059
rect 3328 2051 3330 2070
rect 3336 2064 3338 2146
rect 3350 2141 3356 2142
rect 3350 2137 3351 2141
rect 3355 2137 3356 2141
rect 3350 2136 3356 2137
rect 3352 2127 3354 2136
rect 3351 2126 3355 2127
rect 3351 2121 3355 2122
rect 3428 2108 3430 2202
rect 3487 2198 3491 2199
rect 3487 2193 3491 2194
rect 3488 2182 3490 2193
rect 3500 2192 3502 2274
rect 3576 2271 3578 2290
rect 3575 2270 3579 2271
rect 3575 2265 3579 2266
rect 3576 2250 3578 2265
rect 3574 2249 3580 2250
rect 3574 2245 3575 2249
rect 3579 2245 3580 2249
rect 3574 2244 3580 2245
rect 3574 2232 3580 2233
rect 3574 2228 3575 2232
rect 3579 2228 3580 2232
rect 3574 2227 3580 2228
rect 3576 2199 3578 2227
rect 3575 2198 3579 2199
rect 3575 2193 3579 2194
rect 3498 2191 3504 2192
rect 3498 2187 3499 2191
rect 3503 2187 3504 2191
rect 3498 2186 3504 2187
rect 3486 2181 3492 2182
rect 3486 2177 3487 2181
rect 3491 2177 3492 2181
rect 3486 2176 3492 2177
rect 3576 2169 3578 2193
rect 3574 2168 3580 2169
rect 3574 2164 3575 2168
rect 3579 2164 3580 2168
rect 3574 2163 3580 2164
rect 3574 2151 3580 2152
rect 3574 2147 3575 2151
rect 3579 2147 3580 2151
rect 3574 2146 3580 2147
rect 3478 2141 3484 2142
rect 3478 2137 3479 2141
rect 3483 2137 3484 2141
rect 3478 2136 3484 2137
rect 3480 2127 3482 2136
rect 3498 2135 3504 2136
rect 3498 2131 3499 2135
rect 3503 2131 3504 2135
rect 3498 2130 3504 2131
rect 3471 2126 3475 2127
rect 3471 2121 3475 2122
rect 3479 2126 3483 2127
rect 3479 2121 3483 2122
rect 3472 2116 3474 2121
rect 3470 2115 3476 2116
rect 3470 2111 3471 2115
rect 3475 2111 3476 2115
rect 3470 2110 3476 2111
rect 3426 2107 3432 2108
rect 3426 2103 3427 2107
rect 3431 2103 3432 2107
rect 3426 2102 3432 2103
rect 3478 2075 3484 2076
rect 3478 2071 3479 2075
rect 3483 2071 3484 2075
rect 3478 2070 3484 2071
rect 3334 2063 3340 2064
rect 3334 2059 3335 2063
rect 3339 2059 3340 2063
rect 3334 2058 3340 2059
rect 3470 2063 3476 2064
rect 3470 2059 3471 2063
rect 3475 2059 3476 2063
rect 3470 2058 3476 2059
rect 2727 2050 2731 2051
rect 2727 2045 2731 2046
rect 2759 2050 2763 2051
rect 2759 2045 2763 2046
rect 2887 2050 2891 2051
rect 2887 2045 2891 2046
rect 2935 2050 2939 2051
rect 2935 2045 2939 2046
rect 3039 2050 3043 2051
rect 3039 2045 3043 2046
rect 3119 2050 3123 2051
rect 3119 2045 3123 2046
rect 3183 2050 3187 2051
rect 3183 2045 3187 2046
rect 3311 2050 3315 2051
rect 3311 2045 3315 2046
rect 3327 2050 3331 2051
rect 3327 2045 3331 2046
rect 2618 2043 2624 2044
rect 2618 2039 2619 2043
rect 2623 2039 2624 2043
rect 2618 2038 2624 2039
rect 2682 2043 2688 2044
rect 2682 2039 2683 2043
rect 2687 2039 2688 2043
rect 2682 2038 2688 2039
rect 2590 2033 2596 2034
rect 2590 2029 2591 2033
rect 2595 2029 2596 2033
rect 2590 2028 2596 2029
rect 2684 2020 2686 2038
rect 2760 2034 2762 2045
rect 2870 2043 2876 2044
rect 2870 2039 2871 2043
rect 2875 2039 2876 2043
rect 2870 2038 2876 2039
rect 2758 2033 2764 2034
rect 2758 2029 2759 2033
rect 2763 2029 2764 2033
rect 2758 2028 2764 2029
rect 2872 2020 2874 2038
rect 2936 2034 2938 2045
rect 3120 2034 3122 2045
rect 3222 2043 3228 2044
rect 3222 2039 3223 2043
rect 3227 2039 3228 2043
rect 3222 2038 3228 2039
rect 2934 2033 2940 2034
rect 2934 2029 2935 2033
rect 2939 2029 2940 2033
rect 2934 2028 2940 2029
rect 3118 2033 3124 2034
rect 3118 2029 3119 2033
rect 3123 2029 3124 2033
rect 3118 2028 3124 2029
rect 3224 2020 3226 2038
rect 3312 2034 3314 2045
rect 3310 2033 3316 2034
rect 3310 2029 3311 2033
rect 3315 2029 3316 2033
rect 3310 2028 3316 2029
rect 2682 2019 2688 2020
rect 2682 2015 2683 2019
rect 2687 2015 2688 2019
rect 2682 2014 2688 2015
rect 2870 2019 2876 2020
rect 2870 2015 2871 2019
rect 2875 2015 2876 2019
rect 2870 2014 2876 2015
rect 3222 2019 3228 2020
rect 3222 2015 3223 2019
rect 3227 2015 3228 2019
rect 3222 2014 3228 2015
rect 3310 2003 3316 2004
rect 3310 1999 3311 2003
rect 3315 1999 3316 2003
rect 3310 1998 3316 1999
rect 2582 1993 2588 1994
rect 2582 1989 2583 1993
rect 2587 1989 2588 1993
rect 2582 1988 2588 1989
rect 2750 1993 2756 1994
rect 2750 1989 2751 1993
rect 2755 1989 2756 1993
rect 2750 1988 2756 1989
rect 2926 1993 2932 1994
rect 2926 1989 2927 1993
rect 2931 1989 2932 1993
rect 2926 1988 2932 1989
rect 3110 1993 3116 1994
rect 3110 1989 3111 1993
rect 3115 1989 3116 1993
rect 3110 1988 3116 1989
rect 3302 1993 3308 1994
rect 3302 1989 3303 1993
rect 3307 1989 3308 1993
rect 3302 1988 3308 1989
rect 2584 1979 2586 1988
rect 2752 1979 2754 1988
rect 2928 1979 2930 1988
rect 3112 1979 3114 1988
rect 3304 1979 3306 1988
rect 2503 1978 2507 1979
rect 2503 1973 2507 1974
rect 2583 1978 2587 1979
rect 2583 1973 2587 1974
rect 2655 1978 2659 1979
rect 2655 1973 2659 1974
rect 2751 1978 2755 1979
rect 2751 1973 2755 1974
rect 2839 1978 2843 1979
rect 2839 1973 2843 1974
rect 2927 1978 2931 1979
rect 2927 1973 2931 1974
rect 3047 1978 3051 1979
rect 3047 1973 3051 1974
rect 3111 1978 3115 1979
rect 3111 1973 3115 1974
rect 3271 1978 3275 1979
rect 3271 1973 3275 1974
rect 3303 1978 3307 1979
rect 3303 1973 3307 1974
rect 2504 1968 2506 1973
rect 2656 1968 2658 1973
rect 2840 1968 2842 1973
rect 3048 1968 3050 1973
rect 3272 1968 3274 1973
rect 2502 1967 2508 1968
rect 2502 1963 2503 1967
rect 2507 1963 2508 1967
rect 2502 1962 2508 1963
rect 2654 1967 2660 1968
rect 2654 1963 2655 1967
rect 2659 1963 2660 1967
rect 2654 1962 2660 1963
rect 2838 1967 2844 1968
rect 2838 1963 2839 1967
rect 2843 1963 2844 1967
rect 2838 1962 2844 1963
rect 3046 1967 3052 1968
rect 3046 1963 3047 1967
rect 3051 1963 3052 1967
rect 3046 1962 3052 1963
rect 3270 1967 3276 1968
rect 3270 1963 3271 1967
rect 3275 1963 3276 1967
rect 3270 1962 3276 1963
rect 2450 1959 2456 1960
rect 1862 1957 1868 1958
rect 1239 1954 1243 1955
rect 1239 1949 1243 1950
rect 1263 1954 1267 1955
rect 1263 1949 1267 1950
rect 1359 1954 1363 1955
rect 1359 1949 1363 1950
rect 1423 1954 1427 1955
rect 1423 1949 1427 1950
rect 1487 1954 1491 1955
rect 1487 1949 1491 1950
rect 1583 1954 1587 1955
rect 1583 1949 1587 1950
rect 1727 1954 1731 1955
rect 1727 1949 1731 1950
rect 1823 1954 1827 1955
rect 1862 1953 1863 1957
rect 1867 1953 1868 1957
rect 2450 1955 2451 1959
rect 2455 1955 2456 1959
rect 2450 1954 2456 1955
rect 2570 1959 2576 1960
rect 2570 1955 2571 1959
rect 2575 1955 2576 1959
rect 2570 1954 2576 1955
rect 1862 1952 1868 1953
rect 1823 1949 1827 1950
rect 1264 1944 1266 1949
rect 1424 1944 1426 1949
rect 1584 1944 1586 1949
rect 1728 1944 1730 1949
rect 1262 1943 1268 1944
rect 1262 1939 1263 1943
rect 1267 1939 1268 1943
rect 1262 1938 1268 1939
rect 1422 1943 1428 1944
rect 1422 1939 1423 1943
rect 1427 1939 1428 1943
rect 1422 1938 1428 1939
rect 1582 1943 1588 1944
rect 1582 1939 1583 1943
rect 1587 1939 1588 1943
rect 1582 1938 1588 1939
rect 1726 1943 1732 1944
rect 1726 1939 1727 1943
rect 1731 1939 1732 1943
rect 1726 1938 1732 1939
rect 1718 1935 1724 1936
rect 1718 1931 1719 1935
rect 1723 1931 1724 1935
rect 1824 1934 1826 1949
rect 1862 1940 1868 1941
rect 1862 1936 1863 1940
rect 1867 1936 1868 1940
rect 1862 1935 1868 1936
rect 1718 1930 1724 1931
rect 1822 1933 1828 1934
rect 1270 1903 1276 1904
rect 1270 1899 1271 1903
rect 1275 1899 1276 1903
rect 1270 1898 1276 1899
rect 1430 1903 1436 1904
rect 1430 1899 1431 1903
rect 1435 1899 1436 1903
rect 1430 1898 1436 1899
rect 1590 1903 1596 1904
rect 1590 1899 1591 1903
rect 1595 1899 1596 1903
rect 1590 1898 1596 1899
rect 1134 1891 1140 1892
rect 1134 1887 1135 1891
rect 1139 1887 1140 1891
rect 1134 1886 1140 1887
rect 1272 1879 1274 1898
rect 1432 1879 1434 1898
rect 1592 1879 1594 1898
rect 1063 1878 1067 1879
rect 1063 1873 1067 1874
rect 1103 1878 1107 1879
rect 1103 1873 1107 1874
rect 1231 1878 1235 1879
rect 1231 1873 1235 1874
rect 1271 1878 1275 1879
rect 1271 1873 1275 1874
rect 1391 1878 1395 1879
rect 1391 1873 1395 1874
rect 1431 1878 1435 1879
rect 1431 1873 1435 1874
rect 1551 1878 1555 1879
rect 1551 1873 1555 1874
rect 1591 1878 1595 1879
rect 1591 1873 1595 1874
rect 1711 1878 1715 1879
rect 1711 1873 1715 1874
rect 1064 1862 1066 1873
rect 1134 1871 1140 1872
rect 1134 1866 1135 1871
rect 1139 1866 1140 1871
rect 1135 1863 1139 1864
rect 1232 1862 1234 1873
rect 1299 1868 1303 1869
rect 1299 1863 1303 1864
rect 1062 1861 1068 1862
rect 1062 1857 1063 1861
rect 1067 1857 1068 1861
rect 1062 1856 1068 1857
rect 1230 1861 1236 1862
rect 1230 1857 1231 1861
rect 1235 1857 1236 1861
rect 1230 1856 1236 1857
rect 946 1847 952 1848
rect 946 1843 947 1847
rect 951 1843 952 1847
rect 1300 1844 1302 1863
rect 1392 1862 1394 1873
rect 1552 1862 1554 1873
rect 1712 1862 1714 1873
rect 1720 1872 1722 1930
rect 1822 1929 1823 1933
rect 1827 1929 1828 1933
rect 1822 1928 1828 1929
rect 1822 1916 1828 1917
rect 1822 1912 1823 1916
rect 1827 1912 1828 1916
rect 1822 1911 1828 1912
rect 1734 1903 1740 1904
rect 1734 1899 1735 1903
rect 1739 1899 1740 1903
rect 1734 1898 1740 1899
rect 1736 1879 1738 1898
rect 1824 1879 1826 1911
rect 1864 1903 1866 1935
rect 2030 1927 2036 1928
rect 2030 1923 2031 1927
rect 2035 1923 2036 1927
rect 2030 1922 2036 1923
rect 2118 1927 2124 1928
rect 2118 1923 2119 1927
rect 2123 1923 2124 1927
rect 2118 1922 2124 1923
rect 2206 1927 2212 1928
rect 2206 1923 2207 1927
rect 2211 1923 2212 1927
rect 2206 1922 2212 1923
rect 2294 1927 2300 1928
rect 2294 1923 2295 1927
rect 2299 1923 2300 1927
rect 2294 1922 2300 1923
rect 2390 1927 2396 1928
rect 2390 1923 2391 1927
rect 2395 1923 2396 1927
rect 2390 1922 2396 1923
rect 2510 1927 2516 1928
rect 2510 1923 2511 1927
rect 2515 1923 2516 1927
rect 2510 1922 2516 1923
rect 2032 1903 2034 1922
rect 2042 1915 2048 1916
rect 2042 1911 2043 1915
rect 2047 1911 2048 1915
rect 2042 1910 2048 1911
rect 1863 1902 1867 1903
rect 1863 1897 1867 1898
rect 2031 1902 2035 1903
rect 2031 1897 2035 1898
rect 1735 1878 1739 1879
rect 1735 1873 1739 1874
rect 1823 1878 1827 1879
rect 1823 1873 1827 1874
rect 1864 1873 1866 1897
rect 1718 1871 1724 1872
rect 1718 1867 1719 1871
rect 1723 1867 1724 1871
rect 1718 1866 1724 1867
rect 1390 1861 1396 1862
rect 1390 1857 1391 1861
rect 1395 1857 1396 1861
rect 1390 1856 1396 1857
rect 1550 1861 1556 1862
rect 1550 1857 1551 1861
rect 1555 1857 1556 1861
rect 1550 1856 1556 1857
rect 1710 1861 1716 1862
rect 1710 1857 1711 1861
rect 1715 1857 1716 1861
rect 1710 1856 1716 1857
rect 1824 1849 1826 1873
rect 1862 1872 1868 1873
rect 1862 1868 1863 1872
rect 1867 1868 1868 1872
rect 2044 1868 2046 1910
rect 2120 1903 2122 1922
rect 2208 1903 2210 1922
rect 2296 1903 2298 1922
rect 2392 1903 2394 1922
rect 2512 1903 2514 1922
rect 2572 1916 2574 1954
rect 2646 1943 2652 1944
rect 2646 1939 2647 1943
rect 2651 1939 2652 1943
rect 2646 1938 2652 1939
rect 2722 1943 2728 1944
rect 2722 1939 2723 1943
rect 2727 1939 2728 1943
rect 2722 1938 2728 1939
rect 2906 1943 2912 1944
rect 2906 1939 2907 1943
rect 2911 1939 2912 1943
rect 2906 1938 2912 1939
rect 3114 1943 3120 1944
rect 3114 1939 3115 1943
rect 3119 1939 3120 1943
rect 3114 1938 3120 1939
rect 2570 1915 2576 1916
rect 2570 1911 2571 1915
rect 2575 1911 2576 1915
rect 2570 1910 2576 1911
rect 2119 1902 2123 1903
rect 2119 1897 2123 1898
rect 2175 1902 2179 1903
rect 2175 1897 2179 1898
rect 2207 1902 2211 1903
rect 2207 1897 2211 1898
rect 2263 1902 2267 1903
rect 2263 1897 2267 1898
rect 2295 1902 2299 1903
rect 2295 1897 2299 1898
rect 2351 1902 2355 1903
rect 2351 1897 2355 1898
rect 2391 1902 2395 1903
rect 2391 1897 2395 1898
rect 2439 1902 2443 1903
rect 2439 1897 2443 1898
rect 2511 1902 2515 1903
rect 2511 1897 2515 1898
rect 2527 1902 2531 1903
rect 2527 1897 2531 1898
rect 2639 1902 2643 1903
rect 2639 1897 2643 1898
rect 2176 1886 2178 1897
rect 2242 1895 2248 1896
rect 2242 1891 2243 1895
rect 2247 1891 2248 1895
rect 2242 1890 2248 1891
rect 2174 1885 2180 1886
rect 2174 1881 2175 1885
rect 2179 1881 2180 1885
rect 2174 1880 2180 1881
rect 2244 1868 2246 1890
rect 2264 1886 2266 1897
rect 2330 1895 2336 1896
rect 2330 1891 2331 1895
rect 2335 1891 2336 1895
rect 2330 1890 2336 1891
rect 2262 1885 2268 1886
rect 2262 1881 2263 1885
rect 2267 1881 2268 1885
rect 2262 1880 2268 1881
rect 2332 1868 2334 1890
rect 2352 1886 2354 1897
rect 2418 1895 2424 1896
rect 2418 1891 2419 1895
rect 2423 1891 2424 1895
rect 2418 1890 2424 1891
rect 2350 1885 2356 1886
rect 2350 1881 2351 1885
rect 2355 1881 2356 1885
rect 2350 1880 2356 1881
rect 2420 1868 2422 1890
rect 2440 1886 2442 1897
rect 2528 1886 2530 1897
rect 2534 1895 2540 1896
rect 2534 1891 2535 1895
rect 2539 1891 2540 1895
rect 2534 1890 2540 1891
rect 2438 1885 2444 1886
rect 2438 1881 2439 1885
rect 2443 1881 2444 1885
rect 2438 1880 2444 1881
rect 2526 1885 2532 1886
rect 2526 1881 2527 1885
rect 2531 1881 2532 1885
rect 2526 1880 2532 1881
rect 1862 1867 1868 1868
rect 2042 1867 2048 1868
rect 2042 1863 2043 1867
rect 2047 1863 2048 1867
rect 2042 1862 2048 1863
rect 2242 1867 2248 1868
rect 2242 1863 2243 1867
rect 2247 1863 2248 1867
rect 2242 1862 2248 1863
rect 2330 1867 2336 1868
rect 2330 1863 2331 1867
rect 2335 1863 2336 1867
rect 2330 1862 2336 1863
rect 2418 1867 2424 1868
rect 2418 1863 2419 1867
rect 2423 1863 2424 1867
rect 2418 1862 2424 1863
rect 1862 1855 1868 1856
rect 1862 1851 1863 1855
rect 1867 1851 1868 1855
rect 1862 1850 1868 1851
rect 1822 1848 1828 1849
rect 1822 1844 1823 1848
rect 1827 1844 1828 1848
rect 946 1842 952 1843
rect 1298 1843 1304 1844
rect 1822 1843 1828 1844
rect 1298 1839 1299 1843
rect 1303 1839 1304 1843
rect 1298 1838 1304 1839
rect 1298 1831 1304 1832
rect 1298 1827 1299 1831
rect 1303 1827 1304 1831
rect 1298 1826 1304 1827
rect 1822 1831 1828 1832
rect 1864 1831 1866 1850
rect 2166 1845 2172 1846
rect 2166 1841 2167 1845
rect 2171 1841 2172 1845
rect 2166 1840 2172 1841
rect 2254 1845 2260 1846
rect 2254 1841 2255 1845
rect 2259 1841 2260 1845
rect 2254 1840 2260 1841
rect 2342 1845 2348 1846
rect 2342 1841 2343 1845
rect 2347 1841 2348 1845
rect 2342 1840 2348 1841
rect 2430 1845 2436 1846
rect 2430 1841 2431 1845
rect 2435 1841 2436 1845
rect 2430 1840 2436 1841
rect 2518 1845 2524 1846
rect 2518 1841 2519 1845
rect 2523 1841 2524 1845
rect 2518 1840 2524 1841
rect 2168 1831 2170 1840
rect 2256 1831 2258 1840
rect 2344 1831 2346 1840
rect 2432 1831 2434 1840
rect 2520 1831 2522 1840
rect 1822 1827 1823 1831
rect 1827 1827 1828 1831
rect 1822 1826 1828 1827
rect 1863 1830 1867 1831
rect 694 1821 700 1822
rect 694 1817 695 1821
rect 699 1817 700 1821
rect 694 1816 700 1817
rect 878 1821 884 1822
rect 878 1817 879 1821
rect 883 1817 884 1821
rect 878 1816 884 1817
rect 1054 1821 1060 1822
rect 1054 1817 1055 1821
rect 1059 1817 1060 1821
rect 1054 1816 1060 1817
rect 1222 1821 1228 1822
rect 1222 1817 1223 1821
rect 1227 1817 1228 1821
rect 1222 1816 1228 1817
rect 696 1803 698 1816
rect 880 1803 882 1816
rect 1056 1803 1058 1816
rect 1224 1803 1226 1816
rect 695 1802 699 1803
rect 695 1797 699 1798
rect 719 1802 723 1803
rect 719 1797 723 1798
rect 863 1802 867 1803
rect 863 1797 867 1798
rect 879 1802 883 1803
rect 879 1797 883 1798
rect 1007 1802 1011 1803
rect 1007 1797 1011 1798
rect 1055 1802 1059 1803
rect 1055 1797 1059 1798
rect 1143 1802 1147 1803
rect 1143 1797 1147 1798
rect 1223 1802 1227 1803
rect 1223 1797 1227 1798
rect 1279 1802 1283 1803
rect 1279 1797 1283 1798
rect 720 1792 722 1797
rect 864 1792 866 1797
rect 1008 1792 1010 1797
rect 1144 1792 1146 1797
rect 1280 1792 1282 1797
rect 718 1791 724 1792
rect 718 1787 719 1791
rect 723 1787 724 1791
rect 718 1786 724 1787
rect 862 1791 868 1792
rect 862 1787 863 1791
rect 867 1787 868 1791
rect 862 1786 868 1787
rect 1006 1791 1012 1792
rect 1006 1787 1007 1791
rect 1011 1787 1012 1791
rect 1006 1786 1012 1787
rect 1142 1791 1148 1792
rect 1142 1787 1143 1791
rect 1147 1787 1148 1791
rect 1142 1786 1148 1787
rect 1278 1791 1284 1792
rect 1278 1787 1279 1791
rect 1283 1787 1284 1791
rect 1278 1786 1284 1787
rect 634 1783 640 1784
rect 634 1779 635 1783
rect 639 1779 640 1783
rect 634 1778 640 1779
rect 330 1767 336 1768
rect 330 1763 331 1767
rect 335 1763 336 1767
rect 330 1762 336 1763
rect 786 1767 792 1768
rect 786 1763 787 1767
rect 791 1763 792 1767
rect 786 1762 792 1763
rect 930 1767 936 1768
rect 930 1763 931 1767
rect 935 1763 936 1767
rect 930 1762 936 1763
rect 1074 1767 1080 1768
rect 1074 1763 1075 1767
rect 1079 1763 1080 1767
rect 1074 1762 1080 1763
rect 270 1751 276 1752
rect 270 1747 271 1751
rect 275 1747 276 1751
rect 270 1746 276 1747
rect 154 1739 160 1740
rect 154 1735 155 1739
rect 159 1735 160 1739
rect 272 1735 274 1746
rect 111 1734 115 1735
rect 111 1729 115 1730
rect 143 1734 147 1735
rect 154 1734 160 1735
rect 271 1734 275 1735
rect 143 1729 147 1730
rect 271 1729 275 1730
rect 279 1734 283 1735
rect 279 1729 283 1730
rect 112 1705 114 1729
rect 144 1718 146 1729
rect 218 1727 224 1728
rect 218 1723 219 1727
rect 223 1723 224 1727
rect 218 1722 224 1723
rect 142 1717 148 1718
rect 142 1713 143 1717
rect 147 1713 148 1717
rect 142 1712 148 1713
rect 110 1704 116 1705
rect 110 1700 111 1704
rect 115 1700 116 1704
rect 220 1700 222 1722
rect 280 1718 282 1729
rect 332 1728 334 1762
rect 422 1751 428 1752
rect 422 1747 423 1751
rect 427 1747 428 1751
rect 422 1746 428 1747
rect 574 1751 580 1752
rect 574 1747 575 1751
rect 579 1747 580 1751
rect 574 1746 580 1747
rect 726 1751 732 1752
rect 726 1747 727 1751
rect 731 1747 732 1751
rect 726 1746 732 1747
rect 414 1739 420 1740
rect 414 1735 415 1739
rect 419 1735 420 1739
rect 424 1735 426 1746
rect 576 1735 578 1746
rect 728 1735 730 1746
rect 414 1734 420 1735
rect 423 1734 427 1735
rect 330 1727 336 1728
rect 330 1723 331 1727
rect 335 1723 336 1727
rect 330 1722 336 1723
rect 278 1717 284 1718
rect 278 1713 279 1717
rect 283 1713 284 1717
rect 278 1712 284 1713
rect 416 1700 418 1734
rect 423 1729 427 1730
rect 431 1734 435 1735
rect 431 1729 435 1730
rect 575 1734 579 1735
rect 575 1729 579 1730
rect 583 1734 587 1735
rect 583 1729 587 1730
rect 727 1734 731 1735
rect 727 1729 731 1730
rect 432 1718 434 1729
rect 498 1727 504 1728
rect 498 1723 499 1727
rect 503 1723 504 1727
rect 498 1722 504 1723
rect 430 1717 436 1718
rect 430 1713 431 1717
rect 435 1713 436 1717
rect 430 1712 436 1713
rect 500 1700 502 1722
rect 584 1718 586 1729
rect 728 1718 730 1729
rect 788 1728 790 1762
rect 870 1751 876 1752
rect 870 1747 871 1751
rect 875 1747 876 1751
rect 870 1746 876 1747
rect 872 1735 874 1746
rect 932 1740 934 1762
rect 1014 1751 1020 1752
rect 1014 1747 1015 1751
rect 1019 1747 1020 1751
rect 1014 1746 1020 1747
rect 930 1739 936 1740
rect 930 1735 931 1739
rect 935 1735 936 1739
rect 1016 1735 1018 1746
rect 1076 1740 1078 1762
rect 1150 1751 1156 1752
rect 1150 1747 1151 1751
rect 1155 1747 1156 1751
rect 1150 1746 1156 1747
rect 1286 1751 1292 1752
rect 1286 1747 1287 1751
rect 1291 1747 1292 1751
rect 1286 1746 1292 1747
rect 1074 1739 1080 1740
rect 1074 1735 1075 1739
rect 1079 1735 1080 1739
rect 1152 1735 1154 1746
rect 1288 1735 1290 1746
rect 1300 1740 1302 1826
rect 1382 1821 1388 1822
rect 1382 1817 1383 1821
rect 1387 1817 1388 1821
rect 1382 1816 1388 1817
rect 1542 1821 1548 1822
rect 1542 1817 1543 1821
rect 1547 1817 1548 1821
rect 1542 1816 1548 1817
rect 1702 1821 1708 1822
rect 1702 1817 1703 1821
rect 1707 1817 1708 1821
rect 1702 1816 1708 1817
rect 1384 1803 1386 1816
rect 1544 1803 1546 1816
rect 1704 1803 1706 1816
rect 1824 1803 1826 1826
rect 1863 1825 1867 1826
rect 2167 1830 2171 1831
rect 2167 1825 2171 1826
rect 2255 1830 2259 1831
rect 2255 1825 2259 1826
rect 2319 1830 2323 1831
rect 2319 1825 2323 1826
rect 2343 1830 2347 1831
rect 2343 1825 2347 1826
rect 2431 1830 2435 1831
rect 2431 1825 2435 1826
rect 2439 1830 2443 1831
rect 2439 1825 2443 1826
rect 2519 1830 2523 1831
rect 2519 1825 2523 1826
rect 1864 1810 1866 1825
rect 2320 1820 2322 1825
rect 2440 1820 2442 1825
rect 2318 1819 2324 1820
rect 2318 1815 2319 1819
rect 2323 1815 2324 1819
rect 2318 1814 2324 1815
rect 2438 1819 2444 1820
rect 2438 1815 2439 1819
rect 2443 1815 2444 1819
rect 2438 1814 2444 1815
rect 2536 1812 2538 1890
rect 2640 1886 2642 1897
rect 2648 1896 2650 1938
rect 2662 1927 2668 1928
rect 2662 1923 2663 1927
rect 2667 1923 2668 1927
rect 2662 1922 2668 1923
rect 2664 1903 2666 1922
rect 2724 1916 2726 1938
rect 2846 1927 2852 1928
rect 2846 1923 2847 1927
rect 2851 1923 2852 1927
rect 2846 1922 2852 1923
rect 2722 1915 2728 1916
rect 2722 1911 2723 1915
rect 2727 1911 2728 1915
rect 2722 1910 2728 1911
rect 2848 1903 2850 1922
rect 2908 1916 2910 1938
rect 3054 1927 3060 1928
rect 3054 1923 3055 1927
rect 3059 1923 3060 1927
rect 3054 1922 3060 1923
rect 2906 1915 2912 1916
rect 2906 1911 2907 1915
rect 2911 1911 2912 1915
rect 2906 1910 2912 1911
rect 3056 1903 3058 1922
rect 3116 1916 3118 1938
rect 3278 1927 3284 1928
rect 3278 1923 3279 1927
rect 3283 1923 3284 1927
rect 3278 1922 3284 1923
rect 3114 1915 3120 1916
rect 3114 1911 3115 1915
rect 3119 1911 3120 1915
rect 3114 1910 3120 1911
rect 3280 1903 3282 1922
rect 3312 1916 3314 1998
rect 3310 1915 3316 1916
rect 3310 1911 3311 1915
rect 3315 1911 3316 1915
rect 3310 1910 3316 1911
rect 2663 1902 2667 1903
rect 2663 1897 2667 1898
rect 2775 1902 2779 1903
rect 2775 1897 2779 1898
rect 2847 1902 2851 1903
rect 2847 1897 2851 1898
rect 2935 1902 2939 1903
rect 2935 1897 2939 1898
rect 3055 1902 3059 1903
rect 3055 1897 3059 1898
rect 3119 1902 3123 1903
rect 3119 1897 3123 1898
rect 3279 1902 3283 1903
rect 3279 1897 3283 1898
rect 3311 1902 3315 1903
rect 3311 1897 3315 1898
rect 2646 1895 2652 1896
rect 2646 1891 2647 1895
rect 2651 1891 2652 1895
rect 2646 1890 2652 1891
rect 2776 1886 2778 1897
rect 2890 1895 2896 1896
rect 2890 1891 2891 1895
rect 2895 1891 2896 1895
rect 2890 1890 2896 1891
rect 2638 1885 2644 1886
rect 2638 1881 2639 1885
rect 2643 1881 2644 1885
rect 2638 1880 2644 1881
rect 2774 1885 2780 1886
rect 2774 1881 2775 1885
rect 2779 1881 2780 1885
rect 2774 1880 2780 1881
rect 2892 1872 2894 1890
rect 2936 1886 2938 1897
rect 3120 1886 3122 1897
rect 3312 1886 3314 1897
rect 2934 1885 2940 1886
rect 2934 1881 2935 1885
rect 2939 1881 2940 1885
rect 2934 1880 2940 1881
rect 3118 1885 3124 1886
rect 3118 1881 3119 1885
rect 3123 1881 3124 1885
rect 3118 1880 3124 1881
rect 3310 1885 3316 1886
rect 3310 1881 3311 1885
rect 3315 1881 3316 1885
rect 3310 1880 3316 1881
rect 2890 1871 2896 1872
rect 2890 1867 2891 1871
rect 2895 1867 2896 1871
rect 2890 1866 2896 1867
rect 3198 1855 3204 1856
rect 3198 1851 3199 1855
rect 3203 1851 3204 1855
rect 3198 1850 3204 1851
rect 2630 1845 2636 1846
rect 2630 1841 2631 1845
rect 2635 1841 2636 1845
rect 2630 1840 2636 1841
rect 2766 1845 2772 1846
rect 2766 1841 2767 1845
rect 2771 1841 2772 1845
rect 2766 1840 2772 1841
rect 2926 1845 2932 1846
rect 2926 1841 2927 1845
rect 2931 1841 2932 1845
rect 2926 1840 2932 1841
rect 3110 1845 3116 1846
rect 3110 1841 3111 1845
rect 3115 1841 3116 1845
rect 3110 1840 3116 1841
rect 2632 1831 2634 1840
rect 2768 1831 2770 1840
rect 2928 1831 2930 1840
rect 3112 1831 3114 1840
rect 2559 1830 2563 1831
rect 2559 1825 2563 1826
rect 2631 1830 2635 1831
rect 2631 1825 2635 1826
rect 2679 1830 2683 1831
rect 2679 1825 2683 1826
rect 2767 1830 2771 1831
rect 2767 1825 2771 1826
rect 2799 1830 2803 1831
rect 2799 1825 2803 1826
rect 2919 1830 2923 1831
rect 2919 1825 2923 1826
rect 2927 1830 2931 1831
rect 2927 1825 2931 1826
rect 3047 1830 3051 1831
rect 3047 1825 3051 1826
rect 3111 1830 3115 1831
rect 3111 1825 3115 1826
rect 3183 1830 3187 1831
rect 3183 1825 3187 1826
rect 2560 1820 2562 1825
rect 2680 1820 2682 1825
rect 2800 1820 2802 1825
rect 2920 1820 2922 1825
rect 3048 1820 3050 1825
rect 3184 1820 3186 1825
rect 2558 1819 2564 1820
rect 2558 1815 2559 1819
rect 2563 1815 2564 1819
rect 2558 1814 2564 1815
rect 2678 1819 2684 1820
rect 2678 1815 2679 1819
rect 2683 1815 2684 1819
rect 2678 1814 2684 1815
rect 2798 1819 2804 1820
rect 2798 1815 2799 1819
rect 2803 1815 2804 1819
rect 2798 1814 2804 1815
rect 2918 1819 2924 1820
rect 2918 1815 2919 1819
rect 2923 1815 2924 1819
rect 2918 1814 2924 1815
rect 3046 1819 3052 1820
rect 3046 1815 3047 1819
rect 3051 1815 3052 1819
rect 3046 1814 3052 1815
rect 3182 1819 3188 1820
rect 3182 1815 3183 1819
rect 3187 1815 3188 1819
rect 3182 1814 3188 1815
rect 2534 1811 2540 1812
rect 1862 1809 1868 1810
rect 1862 1805 1863 1809
rect 1867 1805 1868 1809
rect 2534 1807 2535 1811
rect 2539 1807 2540 1811
rect 2534 1806 2540 1807
rect 1862 1804 1868 1805
rect 1383 1802 1387 1803
rect 1383 1797 1387 1798
rect 1423 1802 1427 1803
rect 1423 1797 1427 1798
rect 1543 1802 1547 1803
rect 1543 1797 1547 1798
rect 1703 1802 1707 1803
rect 1703 1797 1707 1798
rect 1823 1802 1827 1803
rect 1823 1797 1827 1798
rect 1424 1792 1426 1797
rect 1422 1791 1428 1792
rect 1422 1787 1423 1791
rect 1427 1787 1428 1791
rect 1422 1786 1428 1787
rect 1346 1783 1352 1784
rect 1346 1779 1347 1783
rect 1351 1779 1352 1783
rect 1824 1782 1826 1797
rect 2506 1795 2512 1796
rect 1862 1792 1868 1793
rect 1862 1788 1863 1792
rect 1867 1788 1868 1792
rect 2506 1791 2507 1795
rect 2511 1791 2512 1795
rect 2506 1790 2512 1791
rect 2626 1795 2632 1796
rect 2626 1791 2627 1795
rect 2631 1791 2632 1795
rect 2626 1790 2632 1791
rect 1862 1787 1868 1788
rect 1346 1778 1352 1779
rect 1822 1781 1828 1782
rect 1298 1739 1304 1740
rect 1298 1735 1299 1739
rect 1303 1735 1304 1739
rect 863 1734 867 1735
rect 863 1729 867 1730
rect 871 1734 875 1735
rect 930 1734 936 1735
rect 991 1734 995 1735
rect 871 1729 875 1730
rect 991 1729 995 1730
rect 1015 1734 1019 1735
rect 1074 1734 1080 1735
rect 1127 1734 1131 1735
rect 1015 1729 1019 1730
rect 1127 1729 1131 1730
rect 1151 1734 1155 1735
rect 1151 1729 1155 1730
rect 1263 1734 1267 1735
rect 1263 1729 1267 1730
rect 1287 1734 1291 1735
rect 1298 1734 1304 1735
rect 1348 1732 1350 1778
rect 1822 1777 1823 1781
rect 1827 1777 1828 1781
rect 1822 1776 1828 1777
rect 1822 1764 1828 1765
rect 1822 1760 1823 1764
rect 1827 1760 1828 1764
rect 1822 1759 1828 1760
rect 1430 1751 1436 1752
rect 1430 1747 1431 1751
rect 1435 1747 1436 1751
rect 1430 1746 1436 1747
rect 1432 1735 1434 1746
rect 1824 1735 1826 1759
rect 1864 1755 1866 1787
rect 2326 1779 2332 1780
rect 2326 1775 2327 1779
rect 2331 1775 2332 1779
rect 2326 1774 2332 1775
rect 2446 1779 2452 1780
rect 2446 1775 2447 1779
rect 2451 1775 2452 1779
rect 2446 1774 2452 1775
rect 2328 1755 2330 1774
rect 2448 1755 2450 1774
rect 2508 1760 2510 1790
rect 2566 1779 2572 1780
rect 2566 1775 2567 1779
rect 2571 1775 2572 1779
rect 2566 1774 2572 1775
rect 2506 1759 2512 1760
rect 2506 1755 2507 1759
rect 2511 1755 2512 1759
rect 2568 1755 2570 1774
rect 2628 1768 2630 1790
rect 2686 1779 2692 1780
rect 2686 1775 2687 1779
rect 2691 1775 2692 1779
rect 2686 1774 2692 1775
rect 2806 1779 2812 1780
rect 2806 1775 2807 1779
rect 2811 1775 2812 1779
rect 2806 1774 2812 1775
rect 2926 1779 2932 1780
rect 2926 1775 2927 1779
rect 2931 1775 2932 1779
rect 2926 1774 2932 1775
rect 3054 1779 3060 1780
rect 3054 1775 3055 1779
rect 3059 1775 3060 1779
rect 3054 1774 3060 1775
rect 3190 1779 3196 1780
rect 3190 1775 3191 1779
rect 3195 1775 3196 1779
rect 3190 1774 3196 1775
rect 2626 1767 2632 1768
rect 2626 1763 2627 1767
rect 2631 1763 2632 1767
rect 2626 1762 2632 1763
rect 2688 1755 2690 1774
rect 2722 1767 2728 1768
rect 2722 1763 2723 1767
rect 2727 1763 2728 1767
rect 2722 1762 2728 1763
rect 1863 1754 1867 1755
rect 1863 1749 1867 1750
rect 2295 1754 2299 1755
rect 2295 1749 2299 1750
rect 2327 1754 2331 1755
rect 2327 1749 2331 1750
rect 2407 1754 2411 1755
rect 2407 1749 2411 1750
rect 2447 1754 2451 1755
rect 2506 1754 2512 1755
rect 2527 1754 2531 1755
rect 2447 1749 2451 1750
rect 2527 1749 2531 1750
rect 2567 1754 2571 1755
rect 2567 1749 2571 1750
rect 2655 1754 2659 1755
rect 2655 1749 2659 1750
rect 2687 1754 2691 1755
rect 2687 1749 2691 1750
rect 1431 1734 1435 1735
rect 1287 1729 1291 1730
rect 1346 1731 1352 1732
rect 786 1727 792 1728
rect 786 1723 787 1727
rect 791 1723 792 1727
rect 786 1722 792 1723
rect 864 1718 866 1729
rect 992 1718 994 1729
rect 1128 1718 1130 1729
rect 1264 1718 1266 1729
rect 1346 1727 1347 1731
rect 1351 1727 1352 1731
rect 1431 1729 1435 1730
rect 1823 1734 1827 1735
rect 1823 1729 1827 1730
rect 1346 1726 1352 1727
rect 582 1717 588 1718
rect 582 1713 583 1717
rect 587 1713 588 1717
rect 582 1712 588 1713
rect 726 1717 732 1718
rect 726 1713 727 1717
rect 731 1713 732 1717
rect 726 1712 732 1713
rect 862 1717 868 1718
rect 862 1713 863 1717
rect 867 1713 868 1717
rect 862 1712 868 1713
rect 990 1717 996 1718
rect 990 1713 991 1717
rect 995 1713 996 1717
rect 990 1712 996 1713
rect 1126 1717 1132 1718
rect 1126 1713 1127 1717
rect 1131 1713 1132 1717
rect 1126 1712 1132 1713
rect 1262 1717 1268 1718
rect 1262 1713 1263 1717
rect 1267 1713 1268 1717
rect 1262 1712 1268 1713
rect 1824 1705 1826 1729
rect 1864 1725 1866 1749
rect 2296 1738 2298 1749
rect 2306 1747 2312 1748
rect 2306 1743 2307 1747
rect 2311 1743 2312 1747
rect 2306 1742 2312 1743
rect 2294 1737 2300 1738
rect 2294 1733 2295 1737
rect 2299 1733 2300 1737
rect 2294 1732 2300 1733
rect 1862 1724 1868 1725
rect 1862 1720 1863 1724
rect 1867 1720 1868 1724
rect 1862 1719 1868 1720
rect 1862 1707 1868 1708
rect 1822 1704 1828 1705
rect 1822 1700 1823 1704
rect 1827 1700 1828 1704
rect 1862 1703 1863 1707
rect 1867 1703 1868 1707
rect 1862 1702 1868 1703
rect 110 1699 116 1700
rect 218 1699 224 1700
rect 218 1695 219 1699
rect 223 1695 224 1699
rect 218 1694 224 1695
rect 414 1699 420 1700
rect 414 1695 415 1699
rect 419 1695 420 1699
rect 414 1694 420 1695
rect 498 1699 504 1700
rect 1822 1699 1828 1700
rect 498 1695 499 1699
rect 503 1695 504 1699
rect 498 1694 504 1695
rect 110 1687 116 1688
rect 110 1683 111 1687
rect 115 1683 116 1687
rect 110 1682 116 1683
rect 1210 1687 1216 1688
rect 1210 1683 1211 1687
rect 1215 1683 1216 1687
rect 1210 1682 1216 1683
rect 1822 1687 1828 1688
rect 1822 1683 1823 1687
rect 1827 1683 1828 1687
rect 1864 1683 1866 1702
rect 2286 1697 2292 1698
rect 2286 1693 2287 1697
rect 2291 1693 2292 1697
rect 2286 1692 2292 1693
rect 2288 1683 2290 1692
rect 1822 1682 1828 1683
rect 1863 1682 1867 1683
rect 112 1667 114 1682
rect 134 1677 140 1678
rect 134 1673 135 1677
rect 139 1673 140 1677
rect 134 1672 140 1673
rect 270 1677 276 1678
rect 270 1673 271 1677
rect 275 1673 276 1677
rect 270 1672 276 1673
rect 422 1677 428 1678
rect 422 1673 423 1677
rect 427 1673 428 1677
rect 422 1672 428 1673
rect 574 1677 580 1678
rect 574 1673 575 1677
rect 579 1673 580 1677
rect 574 1672 580 1673
rect 718 1677 724 1678
rect 718 1673 719 1677
rect 723 1673 724 1677
rect 718 1672 724 1673
rect 854 1677 860 1678
rect 854 1673 855 1677
rect 859 1673 860 1677
rect 854 1672 860 1673
rect 982 1677 988 1678
rect 982 1673 983 1677
rect 987 1673 988 1677
rect 982 1672 988 1673
rect 1118 1677 1124 1678
rect 1118 1673 1119 1677
rect 1123 1673 1124 1677
rect 1118 1672 1124 1673
rect 136 1667 138 1672
rect 154 1671 160 1672
rect 154 1667 155 1671
rect 159 1667 160 1671
rect 272 1667 274 1672
rect 424 1667 426 1672
rect 576 1667 578 1672
rect 720 1667 722 1672
rect 856 1667 858 1672
rect 984 1667 986 1672
rect 1120 1667 1122 1672
rect 111 1666 115 1667
rect 111 1661 115 1662
rect 135 1666 139 1667
rect 154 1666 160 1667
rect 263 1666 267 1667
rect 135 1661 139 1662
rect 112 1646 114 1661
rect 136 1656 138 1661
rect 134 1655 140 1656
rect 134 1651 135 1655
rect 139 1651 140 1655
rect 134 1650 140 1651
rect 110 1645 116 1646
rect 110 1641 111 1645
rect 115 1641 116 1645
rect 110 1640 116 1641
rect 110 1628 116 1629
rect 110 1624 111 1628
rect 115 1624 116 1628
rect 110 1623 116 1624
rect 112 1595 114 1623
rect 142 1615 148 1616
rect 142 1611 143 1615
rect 147 1611 148 1615
rect 142 1610 148 1611
rect 144 1595 146 1610
rect 156 1604 158 1666
rect 263 1661 267 1662
rect 271 1666 275 1667
rect 271 1661 275 1662
rect 423 1666 427 1667
rect 423 1661 427 1662
rect 575 1666 579 1667
rect 575 1661 579 1662
rect 719 1666 723 1667
rect 719 1661 723 1662
rect 727 1666 731 1667
rect 727 1661 731 1662
rect 855 1666 859 1667
rect 855 1661 859 1662
rect 871 1666 875 1667
rect 871 1661 875 1662
rect 983 1666 987 1667
rect 983 1661 987 1662
rect 1007 1666 1011 1667
rect 1007 1661 1011 1662
rect 1119 1666 1123 1667
rect 1119 1661 1123 1662
rect 1143 1666 1147 1667
rect 1143 1661 1147 1662
rect 264 1656 266 1661
rect 424 1656 426 1661
rect 576 1656 578 1661
rect 728 1656 730 1661
rect 872 1656 874 1661
rect 1008 1656 1010 1661
rect 1144 1656 1146 1661
rect 262 1655 268 1656
rect 262 1651 263 1655
rect 267 1651 268 1655
rect 262 1650 268 1651
rect 422 1655 428 1656
rect 422 1651 423 1655
rect 427 1651 428 1655
rect 422 1650 428 1651
rect 574 1655 580 1656
rect 574 1651 575 1655
rect 579 1651 580 1655
rect 574 1650 580 1651
rect 726 1655 732 1656
rect 726 1651 727 1655
rect 731 1651 732 1655
rect 726 1650 732 1651
rect 870 1655 876 1656
rect 870 1651 871 1655
rect 875 1651 876 1655
rect 870 1650 876 1651
rect 1006 1655 1012 1656
rect 1006 1651 1007 1655
rect 1011 1651 1012 1655
rect 1006 1650 1012 1651
rect 1142 1655 1148 1656
rect 1142 1651 1143 1655
rect 1147 1651 1148 1655
rect 1142 1650 1148 1651
rect 202 1647 208 1648
rect 202 1643 203 1647
rect 207 1643 208 1647
rect 202 1642 208 1643
rect 154 1603 160 1604
rect 154 1599 155 1603
rect 159 1599 160 1603
rect 154 1598 160 1599
rect 111 1594 115 1595
rect 111 1589 115 1590
rect 143 1594 147 1595
rect 143 1589 147 1590
rect 167 1594 171 1595
rect 167 1589 171 1590
rect 112 1565 114 1589
rect 168 1578 170 1589
rect 204 1588 206 1642
rect 642 1631 648 1632
rect 642 1627 643 1631
rect 647 1627 648 1631
rect 1098 1631 1104 1632
rect 642 1626 648 1627
rect 1023 1628 1027 1629
rect 270 1615 276 1616
rect 270 1611 271 1615
rect 275 1611 276 1615
rect 270 1610 276 1611
rect 430 1615 436 1616
rect 430 1611 431 1615
rect 435 1611 436 1615
rect 582 1615 588 1616
rect 430 1610 436 1611
rect 443 1612 447 1613
rect 272 1595 274 1610
rect 432 1595 434 1610
rect 582 1611 583 1615
rect 587 1611 588 1615
rect 644 1613 646 1626
rect 1098 1627 1099 1631
rect 1103 1627 1104 1631
rect 1098 1626 1104 1627
rect 1023 1623 1027 1624
rect 734 1615 740 1616
rect 582 1610 588 1611
rect 643 1612 647 1613
rect 443 1607 447 1608
rect 444 1604 446 1607
rect 442 1603 448 1604
rect 442 1599 443 1603
rect 447 1599 448 1603
rect 442 1598 448 1599
rect 584 1595 586 1610
rect 734 1611 735 1615
rect 739 1611 740 1615
rect 734 1610 740 1611
rect 878 1615 884 1616
rect 878 1611 879 1615
rect 883 1611 884 1615
rect 1014 1615 1020 1616
rect 878 1610 884 1611
rect 891 1612 895 1613
rect 643 1607 647 1608
rect 736 1595 738 1610
rect 742 1603 748 1604
rect 742 1599 743 1603
rect 747 1599 748 1603
rect 742 1598 748 1599
rect 271 1594 275 1595
rect 271 1589 275 1590
rect 335 1594 339 1595
rect 335 1589 339 1590
rect 431 1594 435 1595
rect 431 1589 435 1590
rect 511 1594 515 1595
rect 511 1589 515 1590
rect 583 1594 587 1595
rect 583 1589 587 1590
rect 679 1594 683 1595
rect 679 1589 683 1590
rect 735 1594 739 1595
rect 735 1589 739 1590
rect 202 1587 208 1588
rect 202 1583 203 1587
rect 207 1583 208 1587
rect 202 1582 208 1583
rect 336 1578 338 1589
rect 512 1578 514 1589
rect 680 1578 682 1589
rect 166 1577 172 1578
rect 166 1573 167 1577
rect 171 1573 172 1577
rect 166 1572 172 1573
rect 334 1577 340 1578
rect 334 1573 335 1577
rect 339 1573 340 1577
rect 334 1572 340 1573
rect 510 1577 516 1578
rect 510 1573 511 1577
rect 515 1573 516 1577
rect 510 1572 516 1573
rect 678 1577 684 1578
rect 678 1573 679 1577
rect 683 1573 684 1577
rect 678 1572 684 1573
rect 110 1564 116 1565
rect 744 1564 746 1598
rect 750 1595 756 1596
rect 880 1595 882 1610
rect 1014 1611 1015 1615
rect 1019 1611 1020 1615
rect 1014 1610 1020 1611
rect 891 1607 895 1608
rect 892 1604 894 1607
rect 890 1603 896 1604
rect 890 1599 891 1603
rect 895 1599 896 1603
rect 890 1598 896 1599
rect 1016 1595 1018 1610
rect 750 1591 751 1595
rect 755 1591 756 1595
rect 750 1590 756 1591
rect 847 1594 851 1595
rect 110 1560 111 1564
rect 115 1560 116 1564
rect 110 1559 116 1560
rect 742 1563 748 1564
rect 742 1559 743 1563
rect 747 1559 748 1563
rect 752 1560 754 1590
rect 847 1589 851 1590
rect 879 1594 883 1595
rect 879 1589 883 1590
rect 999 1594 1003 1595
rect 999 1589 1003 1590
rect 1015 1594 1019 1595
rect 1015 1589 1019 1590
rect 848 1578 850 1589
rect 858 1587 864 1588
rect 858 1583 859 1587
rect 863 1583 864 1587
rect 858 1582 864 1583
rect 846 1577 852 1578
rect 846 1573 847 1577
rect 851 1573 852 1577
rect 846 1572 852 1573
rect 742 1558 748 1559
rect 750 1559 756 1560
rect 750 1555 751 1559
rect 755 1555 756 1559
rect 750 1554 756 1555
rect 110 1547 116 1548
rect 110 1543 111 1547
rect 115 1543 116 1547
rect 110 1542 116 1543
rect 406 1547 412 1548
rect 406 1543 407 1547
rect 411 1543 412 1547
rect 406 1542 412 1543
rect 112 1523 114 1542
rect 158 1537 164 1538
rect 158 1533 159 1537
rect 163 1533 164 1537
rect 158 1532 164 1533
rect 326 1537 332 1538
rect 326 1533 327 1537
rect 331 1533 332 1537
rect 326 1532 332 1533
rect 160 1523 162 1532
rect 328 1523 330 1532
rect 111 1522 115 1523
rect 111 1517 115 1518
rect 159 1522 163 1523
rect 159 1517 163 1518
rect 215 1522 219 1523
rect 215 1517 219 1518
rect 327 1522 331 1523
rect 327 1517 331 1518
rect 391 1522 395 1523
rect 391 1517 395 1518
rect 112 1502 114 1517
rect 216 1512 218 1517
rect 392 1512 394 1517
rect 214 1511 220 1512
rect 214 1507 215 1511
rect 219 1507 220 1511
rect 214 1506 220 1507
rect 390 1511 396 1512
rect 390 1507 391 1511
rect 395 1507 396 1511
rect 390 1506 396 1507
rect 110 1501 116 1502
rect 110 1497 111 1501
rect 115 1497 116 1501
rect 110 1496 116 1497
rect 282 1487 288 1488
rect 110 1484 116 1485
rect 110 1480 111 1484
rect 115 1480 116 1484
rect 282 1483 283 1487
rect 287 1483 288 1487
rect 282 1482 288 1483
rect 290 1487 296 1488
rect 290 1483 291 1487
rect 295 1483 296 1487
rect 290 1482 296 1483
rect 110 1479 116 1480
rect 112 1451 114 1479
rect 222 1471 228 1472
rect 222 1467 223 1471
rect 227 1467 228 1471
rect 222 1466 228 1467
rect 224 1451 226 1466
rect 111 1450 115 1451
rect 111 1445 115 1446
rect 223 1450 227 1451
rect 223 1445 227 1446
rect 255 1450 259 1451
rect 255 1445 259 1446
rect 112 1421 114 1445
rect 256 1434 258 1445
rect 284 1444 286 1482
rect 292 1460 294 1482
rect 398 1471 404 1472
rect 398 1467 399 1471
rect 403 1467 404 1471
rect 398 1466 404 1467
rect 290 1459 296 1460
rect 290 1455 291 1459
rect 295 1455 296 1459
rect 290 1454 296 1455
rect 400 1451 402 1466
rect 408 1460 410 1542
rect 502 1537 508 1538
rect 502 1533 503 1537
rect 507 1533 508 1537
rect 502 1532 508 1533
rect 670 1537 676 1538
rect 670 1533 671 1537
rect 675 1533 676 1537
rect 670 1532 676 1533
rect 838 1537 844 1538
rect 838 1533 839 1537
rect 843 1533 844 1537
rect 838 1532 844 1533
rect 504 1523 506 1532
rect 672 1523 674 1532
rect 840 1523 842 1532
rect 503 1522 507 1523
rect 503 1517 507 1518
rect 575 1522 579 1523
rect 575 1517 579 1518
rect 671 1522 675 1523
rect 671 1517 675 1518
rect 759 1522 763 1523
rect 759 1517 763 1518
rect 839 1522 843 1523
rect 839 1517 843 1518
rect 576 1512 578 1517
rect 760 1512 762 1517
rect 574 1511 580 1512
rect 574 1507 575 1511
rect 579 1507 580 1511
rect 574 1506 580 1507
rect 758 1511 764 1512
rect 758 1507 759 1511
rect 763 1507 764 1511
rect 758 1506 764 1507
rect 860 1504 862 1582
rect 1000 1578 1002 1589
rect 1024 1588 1026 1623
rect 1100 1604 1102 1626
rect 1150 1615 1156 1616
rect 1150 1611 1151 1615
rect 1155 1611 1156 1615
rect 1212 1613 1214 1682
rect 1254 1677 1260 1678
rect 1254 1673 1255 1677
rect 1259 1673 1260 1677
rect 1254 1672 1260 1673
rect 1256 1667 1258 1672
rect 1824 1667 1826 1682
rect 1863 1677 1867 1678
rect 2143 1682 2147 1683
rect 2143 1677 2147 1678
rect 2247 1682 2251 1683
rect 2247 1677 2251 1678
rect 2287 1682 2291 1683
rect 2308 1680 2310 1742
rect 2408 1738 2410 1749
rect 2528 1738 2530 1749
rect 2656 1738 2658 1749
rect 2714 1747 2720 1748
rect 2714 1743 2715 1747
rect 2719 1743 2720 1747
rect 2714 1742 2720 1743
rect 2406 1737 2412 1738
rect 2406 1733 2407 1737
rect 2411 1733 2412 1737
rect 2406 1732 2412 1733
rect 2526 1737 2532 1738
rect 2526 1733 2527 1737
rect 2531 1733 2532 1737
rect 2526 1732 2532 1733
rect 2654 1737 2660 1738
rect 2654 1733 2655 1737
rect 2659 1733 2660 1737
rect 2654 1732 2660 1733
rect 2716 1724 2718 1742
rect 2714 1723 2720 1724
rect 2714 1719 2715 1723
rect 2719 1719 2720 1723
rect 2724 1720 2726 1762
rect 2808 1755 2810 1774
rect 2819 1772 2823 1773
rect 2818 1767 2824 1768
rect 2818 1763 2819 1767
rect 2823 1763 2824 1767
rect 2818 1762 2824 1763
rect 2928 1755 2930 1774
rect 3056 1755 3058 1774
rect 3192 1755 3194 1774
rect 3200 1773 3202 1850
rect 3302 1845 3308 1846
rect 3302 1841 3303 1845
rect 3307 1841 3308 1845
rect 3302 1840 3308 1841
rect 3304 1831 3306 1840
rect 3303 1830 3307 1831
rect 3303 1825 3307 1826
rect 3319 1830 3323 1831
rect 3319 1825 3323 1826
rect 3463 1830 3467 1831
rect 3463 1825 3467 1826
rect 3320 1820 3322 1825
rect 3464 1820 3466 1825
rect 3318 1819 3324 1820
rect 3318 1815 3319 1819
rect 3323 1815 3324 1819
rect 3318 1814 3324 1815
rect 3462 1819 3468 1820
rect 3462 1815 3463 1819
rect 3467 1815 3468 1819
rect 3462 1814 3468 1815
rect 3472 1808 3474 2058
rect 3480 2051 3482 2070
rect 3479 2050 3483 2051
rect 3479 2045 3483 2046
rect 3487 2050 3491 2051
rect 3487 2045 3491 2046
rect 3488 2034 3490 2045
rect 3500 2044 3502 2130
rect 3576 2127 3578 2146
rect 3575 2126 3579 2127
rect 3575 2121 3579 2122
rect 3576 2106 3578 2121
rect 3574 2105 3580 2106
rect 3574 2101 3575 2105
rect 3579 2101 3580 2105
rect 3574 2100 3580 2101
rect 3574 2088 3580 2089
rect 3574 2084 3575 2088
rect 3579 2084 3580 2088
rect 3574 2083 3580 2084
rect 3576 2051 3578 2083
rect 3575 2050 3579 2051
rect 3575 2045 3579 2046
rect 3498 2043 3504 2044
rect 3498 2039 3499 2043
rect 3503 2039 3504 2043
rect 3498 2038 3504 2039
rect 3486 2033 3492 2034
rect 3486 2029 3487 2033
rect 3491 2029 3492 2033
rect 3486 2028 3492 2029
rect 3576 2021 3578 2045
rect 3574 2020 3580 2021
rect 3574 2016 3575 2020
rect 3579 2016 3580 2020
rect 3574 2015 3580 2016
rect 3574 2003 3580 2004
rect 3574 1999 3575 2003
rect 3579 1999 3580 2003
rect 3574 1998 3580 1999
rect 3478 1993 3484 1994
rect 3478 1989 3479 1993
rect 3483 1989 3484 1993
rect 3478 1988 3484 1989
rect 3480 1979 3482 1988
rect 3526 1987 3532 1988
rect 3526 1983 3527 1987
rect 3531 1983 3532 1987
rect 3526 1982 3532 1983
rect 3479 1978 3483 1979
rect 3479 1973 3483 1974
rect 3480 1968 3482 1973
rect 3478 1967 3484 1968
rect 3478 1963 3479 1967
rect 3483 1963 3484 1967
rect 3478 1962 3484 1963
rect 3486 1927 3492 1928
rect 3486 1923 3487 1927
rect 3491 1923 3492 1927
rect 3486 1922 3492 1923
rect 3488 1903 3490 1922
rect 3528 1916 3530 1982
rect 3576 1979 3578 1998
rect 3575 1978 3579 1979
rect 3575 1973 3579 1974
rect 3576 1958 3578 1973
rect 3574 1957 3580 1958
rect 3574 1953 3575 1957
rect 3579 1953 3580 1957
rect 3574 1952 3580 1953
rect 3574 1940 3580 1941
rect 3574 1936 3575 1940
rect 3579 1936 3580 1940
rect 3574 1935 3580 1936
rect 3526 1915 3532 1916
rect 3526 1911 3527 1915
rect 3531 1911 3532 1915
rect 3526 1910 3532 1911
rect 3576 1903 3578 1935
rect 3487 1902 3491 1903
rect 3487 1897 3491 1898
rect 3575 1902 3579 1903
rect 3575 1897 3579 1898
rect 3488 1886 3490 1897
rect 3486 1885 3492 1886
rect 3486 1881 3487 1885
rect 3491 1881 3492 1885
rect 3486 1880 3492 1881
rect 3576 1873 3578 1897
rect 3574 1872 3580 1873
rect 3574 1868 3575 1872
rect 3579 1868 3580 1872
rect 3574 1867 3580 1868
rect 3574 1855 3580 1856
rect 3574 1851 3575 1855
rect 3579 1851 3580 1855
rect 3574 1850 3580 1851
rect 3478 1845 3484 1846
rect 3478 1841 3479 1845
rect 3483 1841 3484 1845
rect 3478 1840 3484 1841
rect 3480 1831 3482 1840
rect 3498 1839 3504 1840
rect 3498 1835 3499 1839
rect 3503 1835 3504 1839
rect 3498 1834 3504 1835
rect 3479 1830 3483 1831
rect 3479 1825 3483 1826
rect 3470 1807 3476 1808
rect 3470 1803 3471 1807
rect 3475 1803 3476 1807
rect 3470 1802 3476 1803
rect 3390 1795 3396 1796
rect 3390 1791 3391 1795
rect 3395 1791 3396 1795
rect 3390 1790 3396 1791
rect 3326 1779 3332 1780
rect 3326 1775 3327 1779
rect 3331 1775 3332 1779
rect 3326 1774 3332 1775
rect 3199 1772 3203 1773
rect 3199 1767 3203 1768
rect 3328 1755 3330 1774
rect 2775 1754 2779 1755
rect 2775 1749 2779 1750
rect 2807 1754 2811 1755
rect 2807 1749 2811 1750
rect 2895 1754 2899 1755
rect 2895 1749 2899 1750
rect 2927 1754 2931 1755
rect 2927 1749 2931 1750
rect 3015 1754 3019 1755
rect 3015 1749 3019 1750
rect 3055 1754 3059 1755
rect 3055 1749 3059 1750
rect 3135 1754 3139 1755
rect 3135 1749 3139 1750
rect 3191 1754 3195 1755
rect 3191 1749 3195 1750
rect 3255 1754 3259 1755
rect 3255 1749 3259 1750
rect 3327 1754 3331 1755
rect 3327 1749 3331 1750
rect 3383 1754 3387 1755
rect 3383 1749 3387 1750
rect 2776 1738 2778 1749
rect 2896 1738 2898 1749
rect 2966 1747 2972 1748
rect 2966 1743 2967 1747
rect 2971 1743 2972 1747
rect 2966 1742 2972 1743
rect 2774 1737 2780 1738
rect 2774 1733 2775 1737
rect 2779 1733 2780 1737
rect 2774 1732 2780 1733
rect 2894 1737 2900 1738
rect 2894 1733 2895 1737
rect 2899 1733 2900 1737
rect 2894 1732 2900 1733
rect 2968 1720 2970 1742
rect 3016 1738 3018 1749
rect 3042 1747 3048 1748
rect 3042 1743 3043 1747
rect 3047 1743 3048 1747
rect 3042 1742 3048 1743
rect 3014 1737 3020 1738
rect 3014 1733 3015 1737
rect 3019 1733 3020 1737
rect 3014 1732 3020 1733
rect 2714 1718 2720 1719
rect 2722 1719 2728 1720
rect 2722 1715 2723 1719
rect 2727 1715 2728 1719
rect 2722 1714 2728 1715
rect 2966 1719 2972 1720
rect 2966 1715 2967 1719
rect 2971 1715 2972 1719
rect 2966 1714 2972 1715
rect 2854 1707 2860 1708
rect 2854 1703 2855 1707
rect 2859 1703 2860 1707
rect 2854 1702 2860 1703
rect 2398 1697 2404 1698
rect 2398 1693 2399 1697
rect 2403 1693 2404 1697
rect 2398 1692 2404 1693
rect 2518 1697 2524 1698
rect 2518 1693 2519 1697
rect 2523 1693 2524 1697
rect 2518 1692 2524 1693
rect 2646 1697 2652 1698
rect 2646 1693 2647 1697
rect 2651 1693 2652 1697
rect 2646 1692 2652 1693
rect 2766 1697 2772 1698
rect 2766 1693 2767 1697
rect 2771 1693 2772 1697
rect 2766 1692 2772 1693
rect 2400 1683 2402 1692
rect 2520 1683 2522 1692
rect 2648 1683 2650 1692
rect 2768 1683 2770 1692
rect 2367 1682 2371 1683
rect 2287 1677 2291 1678
rect 2306 1679 2312 1680
rect 1255 1666 1259 1667
rect 1255 1661 1259 1662
rect 1279 1666 1283 1667
rect 1279 1661 1283 1662
rect 1415 1666 1419 1667
rect 1415 1661 1419 1662
rect 1823 1666 1827 1667
rect 1864 1662 1866 1677
rect 2144 1672 2146 1677
rect 2248 1672 2250 1677
rect 2306 1675 2307 1679
rect 2311 1675 2312 1679
rect 2367 1677 2371 1678
rect 2399 1682 2403 1683
rect 2399 1677 2403 1678
rect 2503 1682 2507 1683
rect 2503 1677 2507 1678
rect 2519 1682 2523 1683
rect 2519 1677 2523 1678
rect 2647 1682 2651 1683
rect 2647 1677 2651 1678
rect 2767 1682 2771 1683
rect 2767 1677 2771 1678
rect 2807 1682 2811 1683
rect 2807 1677 2811 1678
rect 2306 1674 2312 1675
rect 2368 1672 2370 1677
rect 2504 1672 2506 1677
rect 2648 1672 2650 1677
rect 2808 1672 2810 1677
rect 2142 1671 2148 1672
rect 2142 1667 2143 1671
rect 2147 1667 2148 1671
rect 2142 1666 2148 1667
rect 2246 1671 2252 1672
rect 2246 1667 2247 1671
rect 2251 1667 2252 1671
rect 2246 1666 2252 1667
rect 2366 1671 2372 1672
rect 2366 1667 2367 1671
rect 2371 1667 2372 1671
rect 2366 1666 2372 1667
rect 2502 1671 2508 1672
rect 2502 1667 2503 1671
rect 2507 1667 2508 1671
rect 2502 1666 2508 1667
rect 2646 1671 2652 1672
rect 2646 1667 2647 1671
rect 2651 1667 2652 1671
rect 2646 1666 2652 1667
rect 2806 1671 2812 1672
rect 2806 1667 2807 1671
rect 2811 1667 2812 1671
rect 2806 1666 2812 1667
rect 1823 1661 1827 1662
rect 1862 1661 1868 1662
rect 1280 1656 1282 1661
rect 1416 1656 1418 1661
rect 1278 1655 1284 1656
rect 1278 1651 1279 1655
rect 1283 1651 1284 1655
rect 1278 1650 1284 1651
rect 1414 1655 1420 1656
rect 1414 1651 1415 1655
rect 1419 1651 1420 1655
rect 1414 1650 1420 1651
rect 1346 1647 1352 1648
rect 1346 1643 1347 1647
rect 1351 1643 1352 1647
rect 1824 1646 1826 1661
rect 1862 1657 1863 1661
rect 1867 1657 1868 1661
rect 1862 1656 1868 1657
rect 1346 1642 1352 1643
rect 1822 1645 1828 1646
rect 1348 1629 1350 1642
rect 1822 1641 1823 1645
rect 1827 1641 1828 1645
rect 1822 1640 1828 1641
rect 1862 1644 1868 1645
rect 1862 1640 1863 1644
rect 1867 1640 1868 1644
rect 1862 1639 1868 1640
rect 1347 1628 1351 1629
rect 1347 1623 1351 1624
rect 1822 1628 1828 1629
rect 1822 1624 1823 1628
rect 1827 1624 1828 1628
rect 1822 1623 1828 1624
rect 1286 1615 1292 1616
rect 1150 1610 1156 1611
rect 1211 1612 1215 1613
rect 1098 1603 1104 1604
rect 1098 1599 1099 1603
rect 1103 1599 1104 1603
rect 1098 1598 1104 1599
rect 1152 1595 1154 1610
rect 1286 1611 1287 1615
rect 1291 1611 1292 1615
rect 1286 1610 1292 1611
rect 1422 1615 1428 1616
rect 1422 1611 1423 1615
rect 1427 1611 1428 1615
rect 1422 1610 1428 1611
rect 1211 1607 1215 1608
rect 1288 1595 1290 1610
rect 1424 1595 1426 1610
rect 1824 1595 1826 1623
rect 1864 1615 1866 1639
rect 2150 1631 2156 1632
rect 2150 1627 2151 1631
rect 2155 1627 2156 1631
rect 2150 1626 2156 1627
rect 2254 1631 2260 1632
rect 2254 1627 2255 1631
rect 2259 1627 2260 1631
rect 2254 1626 2260 1627
rect 2374 1631 2380 1632
rect 2374 1627 2375 1631
rect 2379 1627 2380 1631
rect 2374 1626 2380 1627
rect 2510 1631 2516 1632
rect 2510 1627 2511 1631
rect 2515 1627 2516 1631
rect 2510 1626 2516 1627
rect 2654 1631 2660 1632
rect 2654 1627 2655 1631
rect 2659 1627 2660 1631
rect 2654 1626 2660 1627
rect 2814 1631 2820 1632
rect 2814 1627 2815 1631
rect 2819 1627 2820 1631
rect 2814 1626 2820 1627
rect 2152 1615 2154 1626
rect 2226 1619 2232 1620
rect 2226 1615 2227 1619
rect 2231 1615 2232 1619
rect 2256 1615 2258 1626
rect 2376 1615 2378 1626
rect 2512 1615 2514 1626
rect 2656 1615 2658 1626
rect 2816 1615 2818 1626
rect 2856 1620 2858 1702
rect 2886 1697 2892 1698
rect 2886 1693 2887 1697
rect 2891 1693 2892 1697
rect 2886 1692 2892 1693
rect 3006 1697 3012 1698
rect 3006 1693 3007 1697
rect 3011 1693 3012 1697
rect 3006 1692 3012 1693
rect 2888 1683 2890 1692
rect 3008 1683 3010 1692
rect 2887 1682 2891 1683
rect 2887 1677 2891 1678
rect 2975 1682 2979 1683
rect 2975 1677 2979 1678
rect 3007 1682 3011 1683
rect 3007 1677 3011 1678
rect 2976 1672 2978 1677
rect 2974 1671 2980 1672
rect 2974 1667 2975 1671
rect 2979 1667 2980 1671
rect 2974 1666 2980 1667
rect 3044 1664 3046 1742
rect 3136 1738 3138 1749
rect 3256 1738 3258 1749
rect 3384 1738 3386 1749
rect 3392 1748 3394 1790
rect 3470 1779 3476 1780
rect 3470 1775 3471 1779
rect 3475 1775 3476 1779
rect 3470 1774 3476 1775
rect 3462 1767 3468 1768
rect 3462 1763 3463 1767
rect 3467 1763 3468 1767
rect 3462 1762 3468 1763
rect 3390 1747 3396 1748
rect 3390 1743 3391 1747
rect 3395 1743 3396 1747
rect 3390 1742 3396 1743
rect 3134 1737 3140 1738
rect 3134 1733 3135 1737
rect 3139 1733 3140 1737
rect 3134 1732 3140 1733
rect 3254 1737 3260 1738
rect 3254 1733 3255 1737
rect 3259 1733 3260 1737
rect 3254 1732 3260 1733
rect 3382 1737 3388 1738
rect 3382 1733 3383 1737
rect 3387 1733 3388 1737
rect 3382 1732 3388 1733
rect 3334 1707 3340 1708
rect 3334 1703 3335 1707
rect 3339 1703 3340 1707
rect 3334 1702 3340 1703
rect 3126 1697 3132 1698
rect 3126 1693 3127 1697
rect 3131 1693 3132 1697
rect 3126 1692 3132 1693
rect 3246 1697 3252 1698
rect 3246 1693 3247 1697
rect 3251 1693 3252 1697
rect 3246 1692 3252 1693
rect 3128 1683 3130 1692
rect 3248 1683 3250 1692
rect 3127 1682 3131 1683
rect 3127 1677 3131 1678
rect 3143 1682 3147 1683
rect 3143 1677 3147 1678
rect 3247 1682 3251 1683
rect 3247 1677 3251 1678
rect 3319 1682 3323 1683
rect 3319 1677 3323 1678
rect 3144 1672 3146 1677
rect 3320 1672 3322 1677
rect 3142 1671 3148 1672
rect 3142 1667 3143 1671
rect 3147 1667 3148 1671
rect 3142 1666 3148 1667
rect 3318 1671 3324 1672
rect 3318 1667 3319 1671
rect 3323 1667 3324 1671
rect 3318 1666 3324 1667
rect 2954 1663 2960 1664
rect 2954 1659 2955 1663
rect 2959 1659 2960 1663
rect 2954 1658 2960 1659
rect 3042 1663 3048 1664
rect 3042 1659 3043 1663
rect 3047 1659 3048 1663
rect 3042 1658 3048 1659
rect 2854 1619 2860 1620
rect 2854 1615 2855 1619
rect 2859 1615 2860 1619
rect 1863 1614 1867 1615
rect 1863 1609 1867 1610
rect 2007 1614 2011 1615
rect 2007 1609 2011 1610
rect 2103 1614 2107 1615
rect 2103 1609 2107 1610
rect 2151 1614 2155 1615
rect 2151 1609 2155 1610
rect 2207 1614 2211 1615
rect 2226 1614 2232 1615
rect 2255 1614 2259 1615
rect 2207 1609 2211 1610
rect 1151 1594 1155 1595
rect 1151 1589 1155 1590
rect 1287 1594 1291 1595
rect 1287 1589 1291 1590
rect 1295 1594 1299 1595
rect 1295 1589 1299 1590
rect 1423 1594 1427 1595
rect 1423 1589 1427 1590
rect 1439 1594 1443 1595
rect 1439 1589 1443 1590
rect 1583 1594 1587 1595
rect 1583 1589 1587 1590
rect 1823 1594 1827 1595
rect 1823 1589 1827 1590
rect 1022 1587 1028 1588
rect 1022 1583 1023 1587
rect 1027 1583 1028 1587
rect 1022 1582 1028 1583
rect 1152 1578 1154 1589
rect 1296 1578 1298 1589
rect 1440 1578 1442 1589
rect 1584 1578 1586 1589
rect 998 1577 1004 1578
rect 998 1573 999 1577
rect 1003 1573 1004 1577
rect 998 1572 1004 1573
rect 1150 1577 1156 1578
rect 1150 1573 1151 1577
rect 1155 1573 1156 1577
rect 1150 1572 1156 1573
rect 1294 1577 1300 1578
rect 1294 1573 1295 1577
rect 1299 1573 1300 1577
rect 1294 1572 1300 1573
rect 1438 1577 1444 1578
rect 1438 1573 1439 1577
rect 1443 1573 1444 1577
rect 1438 1572 1444 1573
rect 1582 1577 1588 1578
rect 1582 1573 1583 1577
rect 1587 1573 1588 1577
rect 1582 1572 1588 1573
rect 1824 1565 1826 1589
rect 1864 1585 1866 1609
rect 2008 1598 2010 1609
rect 2018 1607 2024 1608
rect 2018 1602 2019 1607
rect 2023 1602 2024 1607
rect 2019 1599 2023 1600
rect 2104 1598 2106 1609
rect 2208 1598 2210 1609
rect 2006 1597 2012 1598
rect 2006 1593 2007 1597
rect 2011 1593 2012 1597
rect 2006 1592 2012 1593
rect 2102 1597 2108 1598
rect 2102 1593 2103 1597
rect 2107 1593 2108 1597
rect 2102 1592 2108 1593
rect 2206 1597 2212 1598
rect 2206 1593 2207 1597
rect 2211 1593 2212 1597
rect 2206 1592 2212 1593
rect 1862 1584 1868 1585
rect 1862 1580 1863 1584
rect 1867 1580 1868 1584
rect 1862 1579 1868 1580
rect 1862 1567 1868 1568
rect 1822 1564 1828 1565
rect 1822 1560 1823 1564
rect 1827 1560 1828 1564
rect 1862 1563 1863 1567
rect 1867 1563 1868 1567
rect 1862 1562 1868 1563
rect 1822 1559 1828 1560
rect 1518 1547 1524 1548
rect 1518 1543 1519 1547
rect 1523 1543 1524 1547
rect 1518 1542 1524 1543
rect 1822 1547 1828 1548
rect 1822 1543 1823 1547
rect 1827 1543 1828 1547
rect 1822 1542 1828 1543
rect 990 1537 996 1538
rect 990 1533 991 1537
rect 995 1533 996 1537
rect 990 1532 996 1533
rect 1142 1537 1148 1538
rect 1142 1533 1143 1537
rect 1147 1533 1148 1537
rect 1142 1532 1148 1533
rect 1286 1537 1292 1538
rect 1286 1533 1287 1537
rect 1291 1533 1292 1537
rect 1286 1532 1292 1533
rect 1430 1537 1436 1538
rect 1430 1533 1431 1537
rect 1435 1533 1436 1537
rect 1430 1532 1436 1533
rect 992 1523 994 1532
rect 1144 1523 1146 1532
rect 1288 1523 1290 1532
rect 1432 1523 1434 1532
rect 935 1522 939 1523
rect 935 1517 939 1518
rect 991 1522 995 1523
rect 991 1517 995 1518
rect 1095 1522 1099 1523
rect 1095 1517 1099 1518
rect 1143 1522 1147 1523
rect 1143 1517 1147 1518
rect 1255 1522 1259 1523
rect 1255 1517 1259 1518
rect 1287 1522 1291 1523
rect 1287 1517 1291 1518
rect 1407 1522 1411 1523
rect 1407 1517 1411 1518
rect 1431 1522 1435 1523
rect 1431 1517 1435 1518
rect 936 1512 938 1517
rect 1096 1512 1098 1517
rect 1256 1512 1258 1517
rect 1408 1512 1410 1517
rect 934 1511 940 1512
rect 934 1507 935 1511
rect 939 1507 940 1511
rect 934 1506 940 1507
rect 1094 1511 1100 1512
rect 1094 1507 1095 1511
rect 1099 1507 1100 1511
rect 1094 1506 1100 1507
rect 1254 1511 1260 1512
rect 1254 1507 1255 1511
rect 1259 1507 1260 1511
rect 1254 1506 1260 1507
rect 1406 1511 1412 1512
rect 1406 1507 1407 1511
rect 1411 1507 1412 1511
rect 1406 1506 1412 1507
rect 858 1503 864 1504
rect 858 1499 859 1503
rect 863 1499 864 1503
rect 858 1498 864 1499
rect 582 1471 588 1472
rect 582 1467 583 1471
rect 587 1467 588 1471
rect 582 1466 588 1467
rect 766 1471 772 1472
rect 766 1467 767 1471
rect 771 1467 772 1471
rect 766 1466 772 1467
rect 942 1471 948 1472
rect 942 1467 943 1471
rect 947 1467 948 1471
rect 942 1466 948 1467
rect 1102 1471 1108 1472
rect 1102 1467 1103 1471
rect 1107 1467 1108 1471
rect 1262 1471 1268 1472
rect 1102 1466 1108 1467
rect 1115 1468 1119 1469
rect 406 1459 412 1460
rect 406 1455 407 1459
rect 411 1455 412 1459
rect 406 1454 412 1455
rect 584 1451 586 1466
rect 738 1459 744 1460
rect 738 1455 739 1459
rect 743 1455 744 1459
rect 738 1454 744 1455
rect 383 1450 387 1451
rect 383 1445 387 1446
rect 399 1450 403 1451
rect 399 1445 403 1446
rect 519 1450 523 1451
rect 519 1445 523 1446
rect 583 1450 587 1451
rect 583 1445 587 1446
rect 671 1450 675 1451
rect 671 1445 675 1446
rect 282 1443 288 1444
rect 282 1439 283 1443
rect 287 1439 288 1443
rect 282 1438 288 1439
rect 330 1443 336 1444
rect 330 1439 331 1443
rect 335 1439 336 1443
rect 330 1438 336 1439
rect 254 1433 260 1434
rect 254 1429 255 1433
rect 259 1429 260 1433
rect 254 1428 260 1429
rect 110 1420 116 1421
rect 332 1420 334 1438
rect 384 1434 386 1445
rect 520 1434 522 1445
rect 672 1434 674 1445
rect 690 1443 696 1444
rect 690 1439 691 1443
rect 695 1439 696 1443
rect 690 1438 696 1439
rect 382 1433 388 1434
rect 382 1429 383 1433
rect 387 1429 388 1433
rect 382 1428 388 1429
rect 518 1433 524 1434
rect 518 1429 519 1433
rect 523 1429 524 1433
rect 518 1428 524 1429
rect 670 1433 676 1434
rect 670 1429 671 1433
rect 675 1429 676 1433
rect 670 1428 676 1429
rect 110 1416 111 1420
rect 115 1416 116 1420
rect 110 1415 116 1416
rect 330 1419 336 1420
rect 330 1415 331 1419
rect 335 1415 336 1419
rect 330 1414 336 1415
rect 110 1403 116 1404
rect 110 1399 111 1403
rect 115 1399 116 1403
rect 110 1398 116 1399
rect 112 1383 114 1398
rect 246 1393 252 1394
rect 246 1389 247 1393
rect 251 1389 252 1393
rect 246 1388 252 1389
rect 374 1393 380 1394
rect 374 1389 375 1393
rect 379 1389 380 1393
rect 374 1388 380 1389
rect 510 1393 516 1394
rect 510 1389 511 1393
rect 515 1389 516 1393
rect 510 1388 516 1389
rect 662 1393 668 1394
rect 662 1389 663 1393
rect 667 1389 668 1393
rect 662 1388 668 1389
rect 248 1383 250 1388
rect 376 1383 378 1388
rect 512 1383 514 1388
rect 542 1387 548 1388
rect 542 1383 543 1387
rect 547 1383 548 1387
rect 664 1383 666 1388
rect 111 1382 115 1383
rect 111 1377 115 1378
rect 247 1382 251 1383
rect 247 1377 251 1378
rect 351 1382 355 1383
rect 351 1377 355 1378
rect 375 1382 379 1383
rect 375 1377 379 1378
rect 439 1382 443 1383
rect 439 1377 443 1378
rect 511 1382 515 1383
rect 511 1377 515 1378
rect 527 1382 531 1383
rect 542 1382 548 1383
rect 623 1382 627 1383
rect 527 1377 531 1378
rect 112 1362 114 1377
rect 352 1372 354 1377
rect 440 1372 442 1377
rect 528 1372 530 1377
rect 350 1371 356 1372
rect 350 1367 351 1371
rect 355 1367 356 1371
rect 350 1366 356 1367
rect 438 1371 444 1372
rect 438 1367 439 1371
rect 443 1367 444 1371
rect 438 1366 444 1367
rect 526 1371 532 1372
rect 526 1367 527 1371
rect 531 1367 532 1371
rect 526 1366 532 1367
rect 110 1361 116 1362
rect 110 1357 111 1361
rect 115 1357 116 1361
rect 110 1356 116 1357
rect 367 1348 371 1349
rect 515 1348 519 1349
rect 110 1344 116 1345
rect 110 1340 111 1344
rect 115 1340 116 1344
rect 367 1343 371 1344
rect 506 1347 512 1348
rect 506 1343 507 1347
rect 511 1343 512 1347
rect 110 1339 116 1340
rect 112 1315 114 1339
rect 358 1331 364 1332
rect 358 1327 359 1331
rect 363 1327 364 1331
rect 358 1326 364 1327
rect 360 1315 362 1326
rect 368 1320 370 1343
rect 506 1342 512 1343
rect 514 1343 515 1348
rect 519 1343 520 1348
rect 514 1342 520 1343
rect 446 1331 452 1332
rect 446 1327 447 1331
rect 451 1327 452 1331
rect 446 1326 452 1327
rect 366 1319 372 1320
rect 366 1315 367 1319
rect 371 1315 372 1319
rect 448 1315 450 1326
rect 111 1314 115 1315
rect 111 1309 115 1310
rect 359 1314 363 1315
rect 366 1314 372 1315
rect 447 1314 451 1315
rect 359 1309 363 1310
rect 447 1309 451 1310
rect 455 1314 459 1315
rect 455 1309 459 1310
rect 112 1285 114 1309
rect 456 1298 458 1309
rect 508 1308 510 1342
rect 534 1331 540 1332
rect 534 1327 535 1331
rect 539 1327 540 1331
rect 534 1326 540 1327
rect 536 1315 538 1326
rect 544 1324 546 1382
rect 623 1377 627 1378
rect 663 1382 667 1383
rect 663 1377 667 1378
rect 624 1372 626 1377
rect 622 1371 628 1372
rect 622 1367 623 1371
rect 627 1367 628 1371
rect 622 1366 628 1367
rect 692 1364 694 1438
rect 740 1404 742 1454
rect 768 1451 770 1466
rect 944 1451 946 1466
rect 1104 1451 1106 1466
rect 1262 1467 1263 1471
rect 1267 1467 1268 1471
rect 1262 1466 1268 1467
rect 1414 1471 1420 1472
rect 1414 1467 1415 1471
rect 1419 1467 1420 1471
rect 1520 1469 1522 1542
rect 1574 1537 1580 1538
rect 1574 1533 1575 1537
rect 1579 1533 1580 1537
rect 1574 1532 1580 1533
rect 1576 1523 1578 1532
rect 1824 1523 1826 1542
rect 1864 1539 1866 1562
rect 1998 1557 2004 1558
rect 1998 1553 1999 1557
rect 2003 1553 2004 1557
rect 1998 1552 2004 1553
rect 2094 1557 2100 1558
rect 2094 1553 2095 1557
rect 2099 1553 2100 1557
rect 2094 1552 2100 1553
rect 2198 1557 2204 1558
rect 2198 1553 2199 1557
rect 2203 1553 2204 1557
rect 2198 1552 2204 1553
rect 2228 1552 2230 1614
rect 2255 1609 2259 1610
rect 2327 1614 2331 1615
rect 2327 1609 2331 1610
rect 2375 1614 2379 1615
rect 2375 1609 2379 1610
rect 2463 1614 2467 1615
rect 2463 1609 2467 1610
rect 2511 1614 2515 1615
rect 2511 1609 2515 1610
rect 2607 1614 2611 1615
rect 2607 1609 2611 1610
rect 2655 1614 2659 1615
rect 2655 1609 2659 1610
rect 2767 1614 2771 1615
rect 2767 1609 2771 1610
rect 2815 1614 2819 1615
rect 2854 1614 2860 1615
rect 2943 1614 2947 1615
rect 2815 1609 2819 1610
rect 2943 1609 2947 1610
rect 2307 1604 2311 1605
rect 2307 1599 2311 1600
rect 2000 1539 2002 1552
rect 2096 1539 2098 1552
rect 2200 1539 2202 1552
rect 2226 1551 2232 1552
rect 2226 1547 2227 1551
rect 2231 1547 2232 1551
rect 2226 1546 2232 1547
rect 1863 1538 1867 1539
rect 1863 1533 1867 1534
rect 1887 1538 1891 1539
rect 1887 1533 1891 1534
rect 1975 1538 1979 1539
rect 1975 1533 1979 1534
rect 1999 1538 2003 1539
rect 1999 1533 2003 1534
rect 2095 1538 2099 1539
rect 2095 1533 2099 1534
rect 2103 1538 2107 1539
rect 2103 1533 2107 1534
rect 2199 1538 2203 1539
rect 2199 1533 2203 1534
rect 2239 1538 2243 1539
rect 2239 1533 2243 1534
rect 1559 1522 1563 1523
rect 1559 1517 1563 1518
rect 1575 1522 1579 1523
rect 1575 1517 1579 1518
rect 1711 1522 1715 1523
rect 1711 1517 1715 1518
rect 1823 1522 1827 1523
rect 1864 1518 1866 1533
rect 1888 1528 1890 1533
rect 1976 1528 1978 1533
rect 2104 1528 2106 1533
rect 2240 1528 2242 1533
rect 1886 1527 1892 1528
rect 1886 1523 1887 1527
rect 1891 1523 1892 1527
rect 1886 1522 1892 1523
rect 1974 1527 1980 1528
rect 1974 1523 1975 1527
rect 1979 1523 1980 1527
rect 1974 1522 1980 1523
rect 2102 1527 2108 1528
rect 2102 1523 2103 1527
rect 2107 1523 2108 1527
rect 2102 1522 2108 1523
rect 2238 1527 2244 1528
rect 2238 1523 2239 1527
rect 2243 1523 2244 1527
rect 2238 1522 2244 1523
rect 2308 1520 2310 1599
rect 2328 1598 2330 1609
rect 2464 1598 2466 1609
rect 2608 1598 2610 1609
rect 2768 1598 2770 1609
rect 2944 1598 2946 1609
rect 2956 1608 2958 1658
rect 2966 1647 2972 1648
rect 2966 1643 2967 1647
rect 2971 1643 2972 1647
rect 2966 1642 2972 1643
rect 2968 1620 2970 1642
rect 2982 1631 2988 1632
rect 2982 1627 2983 1631
rect 2987 1627 2988 1631
rect 2982 1626 2988 1627
rect 3150 1631 3156 1632
rect 3150 1627 3151 1631
rect 3155 1627 3156 1631
rect 3150 1626 3156 1627
rect 3326 1631 3332 1632
rect 3326 1627 3327 1631
rect 3331 1627 3332 1631
rect 3326 1626 3332 1627
rect 2966 1619 2972 1620
rect 2966 1615 2967 1619
rect 2971 1615 2972 1619
rect 2984 1615 2986 1626
rect 3152 1615 3154 1626
rect 3186 1619 3192 1620
rect 3186 1615 3187 1619
rect 3191 1615 3192 1619
rect 3328 1615 3330 1626
rect 3336 1620 3338 1702
rect 3374 1697 3380 1698
rect 3374 1693 3375 1697
rect 3379 1693 3380 1697
rect 3374 1692 3380 1693
rect 3376 1683 3378 1692
rect 3375 1682 3379 1683
rect 3375 1677 3379 1678
rect 3446 1647 3452 1648
rect 3446 1643 3447 1647
rect 3451 1643 3452 1647
rect 3446 1642 3452 1643
rect 3334 1619 3340 1620
rect 3334 1615 3335 1619
rect 3339 1615 3340 1619
rect 2966 1614 2972 1615
rect 2983 1614 2987 1615
rect 2983 1609 2987 1610
rect 3127 1614 3131 1615
rect 3127 1609 3131 1610
rect 3151 1614 3155 1615
rect 3186 1614 3192 1615
rect 3319 1614 3323 1615
rect 3151 1609 3155 1610
rect 2954 1607 2960 1608
rect 2954 1603 2955 1607
rect 2959 1603 2960 1607
rect 2954 1602 2960 1603
rect 3128 1598 3130 1609
rect 2326 1597 2332 1598
rect 2326 1593 2327 1597
rect 2331 1593 2332 1597
rect 2326 1592 2332 1593
rect 2462 1597 2468 1598
rect 2462 1593 2463 1597
rect 2467 1593 2468 1597
rect 2462 1592 2468 1593
rect 2606 1597 2612 1598
rect 2606 1593 2607 1597
rect 2611 1593 2612 1597
rect 2606 1592 2612 1593
rect 2766 1597 2772 1598
rect 2766 1593 2767 1597
rect 2771 1593 2772 1597
rect 2766 1592 2772 1593
rect 2942 1597 2948 1598
rect 2942 1593 2943 1597
rect 2947 1593 2948 1597
rect 2942 1592 2948 1593
rect 3126 1597 3132 1598
rect 3126 1593 3127 1597
rect 3131 1593 3132 1597
rect 3126 1592 3132 1593
rect 3188 1584 3190 1614
rect 3319 1609 3323 1610
rect 3327 1614 3331 1615
rect 3334 1614 3340 1615
rect 3327 1609 3331 1610
rect 3320 1598 3322 1609
rect 3326 1603 3332 1604
rect 3326 1599 3327 1603
rect 3331 1599 3332 1603
rect 3326 1598 3332 1599
rect 3318 1597 3324 1598
rect 3318 1593 3319 1597
rect 3323 1593 3324 1597
rect 3318 1592 3324 1593
rect 3186 1583 3192 1584
rect 3186 1579 3187 1583
rect 3191 1579 3192 1583
rect 3186 1578 3192 1579
rect 2726 1567 2732 1568
rect 2726 1563 2727 1567
rect 2731 1563 2732 1567
rect 2726 1562 2732 1563
rect 2318 1557 2324 1558
rect 2318 1553 2319 1557
rect 2323 1553 2324 1557
rect 2318 1552 2324 1553
rect 2454 1557 2460 1558
rect 2454 1553 2455 1557
rect 2459 1553 2460 1557
rect 2454 1552 2460 1553
rect 2598 1557 2604 1558
rect 2598 1553 2599 1557
rect 2603 1553 2604 1557
rect 2598 1552 2604 1553
rect 2320 1539 2322 1552
rect 2456 1539 2458 1552
rect 2600 1539 2602 1552
rect 2319 1538 2323 1539
rect 2319 1533 2323 1534
rect 2383 1538 2387 1539
rect 2383 1533 2387 1534
rect 2455 1538 2459 1539
rect 2455 1533 2459 1534
rect 2543 1538 2547 1539
rect 2543 1533 2547 1534
rect 2599 1538 2603 1539
rect 2599 1533 2603 1534
rect 2711 1538 2715 1539
rect 2711 1533 2715 1534
rect 2384 1528 2386 1533
rect 2544 1528 2546 1533
rect 2712 1528 2714 1533
rect 2382 1527 2388 1528
rect 2382 1523 2383 1527
rect 2387 1523 2388 1527
rect 2382 1522 2388 1523
rect 2542 1527 2548 1528
rect 2542 1523 2543 1527
rect 2547 1523 2548 1527
rect 2542 1522 2548 1523
rect 2710 1527 2716 1528
rect 2710 1523 2711 1527
rect 2715 1523 2716 1527
rect 2710 1522 2716 1523
rect 2306 1519 2312 1520
rect 1823 1517 1827 1518
rect 1862 1517 1868 1518
rect 1560 1512 1562 1517
rect 1712 1512 1714 1517
rect 1558 1511 1564 1512
rect 1558 1507 1559 1511
rect 1563 1507 1564 1511
rect 1558 1506 1564 1507
rect 1710 1511 1716 1512
rect 1710 1507 1711 1511
rect 1715 1507 1716 1511
rect 1710 1506 1716 1507
rect 1626 1503 1632 1504
rect 1626 1499 1627 1503
rect 1631 1499 1632 1503
rect 1824 1502 1826 1517
rect 1862 1513 1863 1517
rect 1867 1513 1868 1517
rect 2306 1515 2307 1519
rect 2311 1515 2312 1519
rect 2306 1514 2312 1515
rect 1862 1512 1868 1513
rect 2042 1503 2048 1504
rect 1626 1498 1632 1499
rect 1822 1501 1828 1502
rect 1566 1471 1572 1472
rect 1414 1466 1420 1467
rect 1519 1468 1523 1469
rect 1115 1463 1119 1464
rect 1116 1460 1118 1463
rect 1114 1459 1120 1460
rect 1114 1455 1115 1459
rect 1119 1455 1120 1459
rect 1114 1454 1120 1455
rect 1264 1451 1266 1466
rect 1416 1451 1418 1466
rect 1566 1467 1567 1471
rect 1571 1467 1572 1471
rect 1566 1466 1572 1467
rect 1519 1463 1523 1464
rect 1568 1451 1570 1466
rect 1628 1452 1630 1498
rect 1822 1497 1823 1501
rect 1827 1497 1828 1501
rect 1822 1496 1828 1497
rect 1862 1500 1868 1501
rect 1862 1496 1863 1500
rect 1867 1496 1868 1500
rect 2042 1499 2043 1503
rect 2047 1499 2048 1503
rect 2042 1498 2048 1499
rect 2610 1503 2616 1504
rect 2610 1499 2611 1503
rect 2615 1499 2616 1503
rect 2610 1498 2616 1499
rect 1862 1495 1868 1496
rect 1822 1484 1828 1485
rect 1822 1480 1823 1484
rect 1827 1480 1828 1484
rect 1822 1479 1828 1480
rect 1718 1471 1724 1472
rect 1718 1467 1719 1471
rect 1723 1467 1724 1471
rect 1718 1466 1724 1467
rect 1626 1451 1632 1452
rect 1720 1451 1722 1466
rect 1824 1451 1826 1479
rect 1864 1467 1866 1495
rect 1894 1487 1900 1488
rect 1894 1483 1895 1487
rect 1899 1483 1900 1487
rect 1894 1482 1900 1483
rect 1982 1487 1988 1488
rect 1982 1483 1983 1487
rect 1987 1483 1988 1487
rect 1982 1482 1988 1483
rect 1896 1467 1898 1482
rect 1950 1475 1956 1476
rect 1950 1471 1951 1475
rect 1955 1471 1956 1475
rect 1950 1470 1956 1471
rect 1863 1466 1867 1467
rect 1863 1461 1867 1462
rect 1895 1466 1899 1467
rect 1895 1461 1899 1462
rect 767 1450 771 1451
rect 767 1445 771 1446
rect 831 1450 835 1451
rect 831 1445 835 1446
rect 943 1450 947 1451
rect 943 1445 947 1446
rect 991 1450 995 1451
rect 991 1445 995 1446
rect 1103 1450 1107 1451
rect 1103 1445 1107 1446
rect 1143 1450 1147 1451
rect 1143 1445 1147 1446
rect 1263 1450 1267 1451
rect 1263 1445 1267 1446
rect 1295 1450 1299 1451
rect 1295 1445 1299 1446
rect 1415 1450 1419 1451
rect 1415 1445 1419 1446
rect 1447 1450 1451 1451
rect 1447 1445 1451 1446
rect 1567 1450 1571 1451
rect 1567 1445 1571 1446
rect 1599 1450 1603 1451
rect 1626 1447 1627 1451
rect 1631 1447 1632 1451
rect 1626 1446 1632 1447
rect 1719 1450 1723 1451
rect 1599 1445 1603 1446
rect 1719 1445 1723 1446
rect 1735 1450 1739 1451
rect 1735 1445 1739 1446
rect 1823 1450 1827 1451
rect 1823 1445 1827 1446
rect 832 1434 834 1445
rect 992 1434 994 1445
rect 1144 1434 1146 1445
rect 1202 1443 1208 1444
rect 1202 1439 1203 1443
rect 1207 1439 1208 1443
rect 1202 1438 1208 1439
rect 830 1433 836 1434
rect 830 1429 831 1433
rect 835 1429 836 1433
rect 830 1428 836 1429
rect 990 1433 996 1434
rect 990 1429 991 1433
rect 995 1429 996 1433
rect 990 1428 996 1429
rect 1142 1433 1148 1434
rect 1142 1429 1143 1433
rect 1147 1429 1148 1433
rect 1142 1428 1148 1429
rect 738 1403 744 1404
rect 738 1399 739 1403
rect 743 1399 744 1403
rect 738 1398 744 1399
rect 898 1403 904 1404
rect 898 1399 899 1403
rect 903 1399 904 1403
rect 898 1398 904 1399
rect 822 1393 828 1394
rect 822 1389 823 1393
rect 827 1389 828 1393
rect 822 1388 828 1389
rect 824 1383 826 1388
rect 727 1382 731 1383
rect 727 1377 731 1378
rect 823 1382 827 1383
rect 823 1377 827 1378
rect 847 1382 851 1383
rect 847 1377 851 1378
rect 728 1372 730 1377
rect 848 1372 850 1377
rect 726 1371 732 1372
rect 726 1367 727 1371
rect 731 1367 732 1371
rect 726 1366 732 1367
rect 846 1371 852 1372
rect 846 1367 847 1371
rect 851 1367 852 1371
rect 846 1366 852 1367
rect 690 1363 696 1364
rect 690 1359 691 1363
rect 695 1359 696 1363
rect 690 1358 696 1359
rect 794 1347 800 1348
rect 794 1343 795 1347
rect 799 1343 800 1347
rect 794 1342 800 1343
rect 630 1331 636 1332
rect 630 1327 631 1331
rect 635 1327 636 1331
rect 630 1326 636 1327
rect 734 1331 740 1332
rect 734 1327 735 1331
rect 739 1327 740 1331
rect 734 1326 740 1327
rect 542 1323 548 1324
rect 542 1319 543 1323
rect 547 1319 548 1323
rect 542 1318 548 1319
rect 632 1315 634 1326
rect 736 1315 738 1326
rect 796 1320 798 1342
rect 854 1331 860 1332
rect 854 1327 855 1331
rect 859 1327 860 1331
rect 854 1326 860 1327
rect 794 1319 800 1320
rect 794 1315 795 1319
rect 799 1315 800 1319
rect 856 1315 858 1326
rect 900 1320 902 1398
rect 982 1393 988 1394
rect 982 1389 983 1393
rect 987 1389 988 1393
rect 982 1388 988 1389
rect 1134 1393 1140 1394
rect 1134 1389 1135 1393
rect 1139 1389 1140 1393
rect 1134 1388 1140 1389
rect 984 1383 986 1388
rect 1136 1383 1138 1388
rect 983 1382 987 1383
rect 983 1377 987 1378
rect 1127 1382 1131 1383
rect 1127 1377 1131 1378
rect 1135 1382 1139 1383
rect 1135 1377 1139 1378
rect 984 1372 986 1377
rect 1128 1372 1130 1377
rect 982 1371 988 1372
rect 982 1367 983 1371
rect 987 1367 988 1371
rect 982 1366 988 1367
rect 1126 1371 1132 1372
rect 1126 1367 1127 1371
rect 1131 1367 1132 1371
rect 1126 1366 1132 1367
rect 1204 1364 1206 1438
rect 1296 1434 1298 1445
rect 1448 1434 1450 1445
rect 1600 1434 1602 1445
rect 1678 1443 1684 1444
rect 1678 1439 1679 1443
rect 1683 1439 1684 1443
rect 1678 1438 1684 1439
rect 1294 1433 1300 1434
rect 1294 1429 1295 1433
rect 1299 1429 1300 1433
rect 1294 1428 1300 1429
rect 1446 1433 1452 1434
rect 1446 1429 1447 1433
rect 1451 1429 1452 1433
rect 1446 1428 1452 1429
rect 1598 1433 1604 1434
rect 1598 1429 1599 1433
rect 1603 1429 1604 1433
rect 1598 1428 1604 1429
rect 1286 1393 1292 1394
rect 1286 1389 1287 1393
rect 1291 1389 1292 1393
rect 1286 1388 1292 1389
rect 1438 1393 1444 1394
rect 1438 1389 1439 1393
rect 1443 1389 1444 1393
rect 1438 1388 1444 1389
rect 1590 1393 1596 1394
rect 1590 1389 1591 1393
rect 1595 1389 1596 1393
rect 1590 1388 1596 1389
rect 1288 1383 1290 1388
rect 1440 1383 1442 1388
rect 1592 1383 1594 1388
rect 1279 1382 1283 1383
rect 1279 1377 1283 1378
rect 1287 1382 1291 1383
rect 1287 1377 1291 1378
rect 1431 1382 1435 1383
rect 1431 1377 1435 1378
rect 1439 1382 1443 1383
rect 1439 1377 1443 1378
rect 1591 1382 1595 1383
rect 1591 1377 1595 1378
rect 1280 1372 1282 1377
rect 1432 1372 1434 1377
rect 1592 1372 1594 1377
rect 1278 1371 1284 1372
rect 1278 1367 1279 1371
rect 1283 1367 1284 1371
rect 1278 1366 1284 1367
rect 1430 1371 1436 1372
rect 1430 1367 1431 1371
rect 1435 1367 1436 1371
rect 1430 1366 1436 1367
rect 1590 1371 1596 1372
rect 1590 1367 1591 1371
rect 1595 1367 1596 1371
rect 1590 1366 1596 1367
rect 1680 1364 1682 1438
rect 1736 1434 1738 1445
rect 1734 1433 1740 1434
rect 1734 1429 1735 1433
rect 1739 1429 1740 1433
rect 1734 1428 1740 1429
rect 1824 1421 1826 1445
rect 1864 1437 1866 1461
rect 1896 1450 1898 1461
rect 1894 1449 1900 1450
rect 1894 1445 1895 1449
rect 1899 1445 1900 1449
rect 1894 1444 1900 1445
rect 1952 1437 1954 1470
rect 1984 1467 1986 1482
rect 2044 1476 2046 1498
rect 2110 1487 2116 1488
rect 2110 1483 2111 1487
rect 2115 1483 2116 1487
rect 2110 1482 2116 1483
rect 2246 1487 2252 1488
rect 2246 1483 2247 1487
rect 2251 1483 2252 1487
rect 2246 1482 2252 1483
rect 2390 1487 2396 1488
rect 2390 1483 2391 1487
rect 2395 1483 2396 1487
rect 2390 1482 2396 1483
rect 2550 1487 2556 1488
rect 2550 1483 2551 1487
rect 2555 1483 2556 1487
rect 2550 1482 2556 1483
rect 2042 1475 2048 1476
rect 2042 1471 2043 1475
rect 2047 1471 2048 1475
rect 2042 1470 2048 1471
rect 2112 1467 2114 1482
rect 2248 1467 2250 1482
rect 2392 1467 2394 1482
rect 2552 1467 2554 1482
rect 2612 1476 2614 1498
rect 2718 1487 2724 1488
rect 2718 1483 2719 1487
rect 2723 1483 2724 1487
rect 2718 1482 2724 1483
rect 2610 1475 2616 1476
rect 2610 1471 2611 1475
rect 2615 1471 2616 1475
rect 2610 1470 2616 1471
rect 2720 1467 2722 1482
rect 2728 1476 2730 1562
rect 2758 1557 2764 1558
rect 2758 1553 2759 1557
rect 2763 1553 2764 1557
rect 2758 1552 2764 1553
rect 2934 1557 2940 1558
rect 2934 1553 2935 1557
rect 2939 1553 2940 1557
rect 2934 1552 2940 1553
rect 3118 1557 3124 1558
rect 3118 1553 3119 1557
rect 3123 1553 3124 1557
rect 3118 1552 3124 1553
rect 3310 1557 3316 1558
rect 3310 1553 3311 1557
rect 3315 1553 3316 1557
rect 3310 1552 3316 1553
rect 2760 1539 2762 1552
rect 2936 1539 2938 1552
rect 3120 1539 3122 1552
rect 3312 1539 3314 1552
rect 2759 1538 2763 1539
rect 2759 1533 2763 1534
rect 2879 1538 2883 1539
rect 2879 1533 2883 1534
rect 2935 1538 2939 1539
rect 2935 1533 2939 1534
rect 3055 1538 3059 1539
rect 3055 1533 3059 1534
rect 3119 1538 3123 1539
rect 3119 1533 3123 1534
rect 3239 1538 3243 1539
rect 3239 1533 3243 1534
rect 3311 1538 3315 1539
rect 3311 1533 3315 1534
rect 2880 1528 2882 1533
rect 3056 1528 3058 1533
rect 3240 1528 3242 1533
rect 2878 1527 2884 1528
rect 2878 1523 2879 1527
rect 2883 1523 2884 1527
rect 2878 1522 2884 1523
rect 3054 1527 3060 1528
rect 3054 1523 3055 1527
rect 3059 1523 3060 1527
rect 3054 1522 3060 1523
rect 3238 1527 3244 1528
rect 3238 1523 3239 1527
rect 3243 1523 3244 1527
rect 3238 1522 3244 1523
rect 3328 1520 3330 1598
rect 3431 1538 3435 1539
rect 3431 1533 3435 1534
rect 3432 1528 3434 1533
rect 3430 1527 3436 1528
rect 3430 1523 3431 1527
rect 3435 1523 3436 1527
rect 3430 1522 3436 1523
rect 3326 1519 3332 1520
rect 3326 1515 3327 1519
rect 3331 1515 3332 1519
rect 3326 1514 3332 1515
rect 3122 1503 3128 1504
rect 3122 1499 3123 1503
rect 3127 1499 3128 1503
rect 3122 1498 3128 1499
rect 2886 1487 2892 1488
rect 2886 1483 2887 1487
rect 2891 1483 2892 1487
rect 2886 1482 2892 1483
rect 3062 1487 3068 1488
rect 3062 1483 3063 1487
rect 3067 1483 3068 1487
rect 3062 1482 3068 1483
rect 2726 1475 2732 1476
rect 2726 1471 2727 1475
rect 2731 1471 2732 1475
rect 2726 1470 2732 1471
rect 2826 1475 2832 1476
rect 2826 1471 2827 1475
rect 2831 1471 2832 1475
rect 2826 1470 2832 1471
rect 1983 1466 1987 1467
rect 1983 1461 1987 1462
rect 2023 1466 2027 1467
rect 2023 1461 2027 1462
rect 2111 1466 2115 1467
rect 2111 1461 2115 1462
rect 2175 1466 2179 1467
rect 2175 1461 2179 1462
rect 2247 1466 2251 1467
rect 2247 1461 2251 1462
rect 2319 1466 2323 1467
rect 2319 1461 2323 1462
rect 2391 1466 2395 1467
rect 2391 1461 2395 1462
rect 2463 1466 2467 1467
rect 2463 1461 2467 1462
rect 2551 1466 2555 1467
rect 2551 1461 2555 1462
rect 2615 1466 2619 1467
rect 2615 1461 2619 1462
rect 2719 1466 2723 1467
rect 2719 1461 2723 1462
rect 2767 1466 2771 1467
rect 2767 1461 2771 1462
rect 2024 1450 2026 1461
rect 2176 1450 2178 1461
rect 2234 1459 2240 1460
rect 2234 1455 2235 1459
rect 2239 1455 2240 1459
rect 2234 1454 2240 1455
rect 2022 1449 2028 1450
rect 2022 1445 2023 1449
rect 2027 1445 2028 1449
rect 2022 1444 2028 1445
rect 2174 1449 2180 1450
rect 2174 1445 2175 1449
rect 2179 1445 2180 1449
rect 2174 1444 2180 1445
rect 1862 1436 1868 1437
rect 1862 1432 1863 1436
rect 1867 1432 1868 1436
rect 1862 1431 1868 1432
rect 1951 1436 1955 1437
rect 2236 1436 2238 1454
rect 2320 1450 2322 1461
rect 2464 1450 2466 1461
rect 2518 1459 2524 1460
rect 2518 1455 2519 1459
rect 2523 1455 2524 1459
rect 2518 1454 2524 1455
rect 2318 1449 2324 1450
rect 2318 1445 2319 1449
rect 2323 1445 2324 1449
rect 2318 1444 2324 1445
rect 2462 1449 2468 1450
rect 2462 1445 2463 1449
rect 2467 1445 2468 1449
rect 2462 1444 2468 1445
rect 2243 1436 2247 1437
rect 1951 1431 1955 1432
rect 2234 1435 2240 1436
rect 2234 1431 2235 1435
rect 2239 1431 2240 1435
rect 2234 1430 2240 1431
rect 2242 1431 2248 1432
rect 2242 1427 2243 1431
rect 2247 1427 2248 1431
rect 2242 1426 2248 1427
rect 1822 1420 1828 1421
rect 1822 1416 1823 1420
rect 1827 1416 1828 1420
rect 1822 1415 1828 1416
rect 1862 1419 1868 1420
rect 1862 1415 1863 1419
rect 1867 1415 1868 1419
rect 1862 1414 1868 1415
rect 2378 1415 2384 1416
rect 1718 1403 1724 1404
rect 1718 1399 1719 1403
rect 1723 1399 1724 1403
rect 1718 1398 1724 1399
rect 1822 1403 1828 1404
rect 1822 1399 1823 1403
rect 1827 1399 1828 1403
rect 1822 1398 1828 1399
rect 1202 1363 1208 1364
rect 1202 1359 1203 1363
rect 1207 1359 1208 1363
rect 1202 1358 1208 1359
rect 1678 1363 1684 1364
rect 1678 1359 1679 1363
rect 1683 1359 1684 1363
rect 1678 1358 1684 1359
rect 1451 1332 1455 1333
rect 990 1331 996 1332
rect 990 1327 991 1331
rect 995 1327 996 1331
rect 990 1326 996 1327
rect 1134 1331 1140 1332
rect 1134 1327 1135 1331
rect 1139 1327 1140 1331
rect 1134 1326 1140 1327
rect 1286 1331 1292 1332
rect 1286 1327 1287 1331
rect 1291 1327 1292 1331
rect 1286 1326 1292 1327
rect 1438 1331 1444 1332
rect 1438 1327 1439 1331
rect 1443 1327 1444 1331
rect 1451 1327 1455 1328
rect 1598 1331 1604 1332
rect 1598 1327 1599 1331
rect 1603 1327 1604 1331
rect 1438 1326 1444 1327
rect 898 1319 904 1320
rect 898 1315 899 1319
rect 903 1315 904 1319
rect 992 1315 994 1326
rect 1026 1319 1032 1320
rect 1026 1315 1027 1319
rect 1031 1315 1032 1319
rect 1136 1315 1138 1326
rect 1288 1315 1290 1326
rect 1440 1315 1442 1326
rect 1452 1320 1454 1327
rect 1598 1326 1604 1327
rect 1450 1319 1456 1320
rect 1450 1315 1451 1319
rect 1455 1315 1456 1319
rect 1600 1315 1602 1326
rect 1720 1320 1722 1398
rect 1726 1393 1732 1394
rect 1726 1389 1727 1393
rect 1731 1389 1732 1393
rect 1726 1388 1732 1389
rect 1728 1383 1730 1388
rect 1824 1383 1826 1398
rect 1864 1387 1866 1414
rect 2378 1411 2379 1415
rect 2383 1411 2384 1415
rect 2378 1410 2384 1411
rect 1886 1409 1892 1410
rect 1886 1405 1887 1409
rect 1891 1405 1892 1409
rect 1886 1404 1892 1405
rect 2014 1409 2020 1410
rect 2014 1405 2015 1409
rect 2019 1405 2020 1409
rect 2014 1404 2020 1405
rect 2166 1409 2172 1410
rect 2166 1405 2167 1409
rect 2171 1405 2172 1409
rect 2166 1404 2172 1405
rect 2310 1409 2316 1410
rect 2310 1405 2311 1409
rect 2315 1405 2316 1409
rect 2310 1404 2316 1405
rect 1888 1387 1890 1404
rect 2016 1387 2018 1404
rect 2168 1387 2170 1404
rect 2312 1387 2314 1404
rect 1863 1386 1867 1387
rect 1727 1382 1731 1383
rect 1727 1377 1731 1378
rect 1823 1382 1827 1383
rect 1863 1381 1867 1382
rect 1887 1386 1891 1387
rect 1887 1381 1891 1382
rect 2015 1386 2019 1387
rect 2015 1381 2019 1382
rect 2143 1386 2147 1387
rect 2143 1381 2147 1382
rect 2167 1386 2171 1387
rect 2167 1381 2171 1382
rect 2311 1386 2315 1387
rect 2311 1381 2315 1382
rect 1823 1377 1827 1378
rect 1728 1372 1730 1377
rect 1726 1371 1732 1372
rect 1726 1367 1727 1371
rect 1731 1367 1732 1371
rect 1726 1366 1732 1367
rect 1824 1362 1826 1377
rect 1864 1366 1866 1381
rect 1888 1376 1890 1381
rect 2144 1376 2146 1381
rect 1886 1375 1892 1376
rect 1886 1371 1887 1375
rect 1891 1371 1892 1375
rect 1886 1370 1892 1371
rect 2142 1375 2148 1376
rect 2142 1371 2143 1375
rect 2147 1371 2148 1375
rect 2142 1370 2148 1371
rect 1862 1365 1868 1366
rect 1822 1361 1828 1362
rect 1822 1357 1823 1361
rect 1827 1357 1828 1361
rect 1862 1361 1863 1365
rect 1867 1361 1868 1365
rect 1862 1360 1868 1361
rect 1822 1356 1828 1357
rect 1870 1351 1876 1352
rect 1862 1348 1868 1349
rect 1822 1344 1828 1345
rect 1822 1340 1823 1344
rect 1827 1340 1828 1344
rect 1862 1344 1863 1348
rect 1867 1344 1868 1348
rect 1870 1347 1871 1351
rect 1875 1347 1876 1351
rect 1870 1346 1876 1347
rect 1862 1343 1868 1344
rect 1822 1339 1828 1340
rect 1734 1331 1740 1332
rect 1734 1327 1735 1331
rect 1739 1327 1740 1331
rect 1734 1326 1740 1327
rect 1718 1319 1724 1320
rect 1718 1315 1719 1319
rect 1723 1315 1724 1319
rect 1736 1315 1738 1326
rect 1824 1315 1826 1339
rect 1864 1319 1866 1343
rect 1872 1333 1874 1346
rect 1894 1335 1900 1336
rect 1871 1332 1875 1333
rect 1894 1331 1895 1335
rect 1899 1331 1900 1335
rect 1894 1330 1900 1331
rect 2150 1335 2156 1336
rect 2150 1331 2151 1335
rect 2155 1331 2156 1335
rect 2150 1330 2156 1331
rect 1871 1327 1875 1328
rect 1896 1319 1898 1330
rect 1906 1323 1912 1324
rect 1906 1319 1907 1323
rect 1911 1319 1912 1323
rect 2152 1319 2154 1330
rect 2380 1324 2382 1410
rect 2454 1409 2460 1410
rect 2454 1405 2455 1409
rect 2459 1405 2460 1409
rect 2454 1404 2460 1405
rect 2456 1387 2458 1404
rect 2391 1386 2395 1387
rect 2391 1381 2395 1382
rect 2455 1386 2459 1387
rect 2455 1381 2459 1382
rect 2392 1376 2394 1381
rect 2390 1375 2396 1376
rect 2390 1371 2391 1375
rect 2395 1371 2396 1375
rect 2390 1370 2396 1371
rect 2520 1368 2522 1454
rect 2616 1450 2618 1461
rect 2768 1450 2770 1461
rect 2614 1449 2620 1450
rect 2614 1445 2615 1449
rect 2619 1445 2620 1449
rect 2614 1444 2620 1445
rect 2766 1449 2772 1450
rect 2766 1445 2767 1449
rect 2771 1445 2772 1449
rect 2766 1444 2772 1445
rect 2828 1436 2830 1470
rect 2888 1467 2890 1482
rect 3064 1467 3066 1482
rect 2887 1466 2891 1467
rect 2887 1461 2891 1462
rect 2935 1466 2939 1467
rect 2935 1461 2939 1462
rect 3063 1466 3067 1467
rect 3063 1461 3067 1462
rect 3103 1466 3107 1467
rect 3103 1461 3107 1462
rect 2936 1450 2938 1461
rect 3104 1450 3106 1461
rect 3124 1460 3126 1498
rect 3246 1487 3252 1488
rect 3246 1483 3247 1487
rect 3251 1483 3252 1487
rect 3246 1482 3252 1483
rect 3438 1487 3444 1488
rect 3438 1483 3439 1487
rect 3443 1483 3444 1487
rect 3438 1482 3444 1483
rect 3248 1467 3250 1482
rect 3440 1467 3442 1482
rect 3448 1476 3450 1642
rect 3464 1580 3466 1762
rect 3472 1755 3474 1774
rect 3471 1754 3475 1755
rect 3471 1749 3475 1750
rect 3487 1754 3491 1755
rect 3487 1749 3491 1750
rect 3488 1738 3490 1749
rect 3500 1748 3502 1834
rect 3576 1831 3578 1850
rect 3575 1830 3579 1831
rect 3575 1825 3579 1826
rect 3576 1810 3578 1825
rect 3574 1809 3580 1810
rect 3574 1805 3575 1809
rect 3579 1805 3580 1809
rect 3574 1804 3580 1805
rect 3574 1792 3580 1793
rect 3574 1788 3575 1792
rect 3579 1788 3580 1792
rect 3574 1787 3580 1788
rect 3576 1755 3578 1787
rect 3575 1754 3579 1755
rect 3575 1749 3579 1750
rect 3498 1747 3504 1748
rect 3498 1743 3499 1747
rect 3503 1743 3504 1747
rect 3498 1742 3504 1743
rect 3486 1737 3492 1738
rect 3486 1733 3487 1737
rect 3491 1733 3492 1737
rect 3486 1732 3492 1733
rect 3576 1725 3578 1749
rect 3574 1724 3580 1725
rect 3574 1720 3575 1724
rect 3579 1720 3580 1724
rect 3574 1719 3580 1720
rect 3574 1707 3580 1708
rect 3574 1703 3575 1707
rect 3579 1703 3580 1707
rect 3574 1702 3580 1703
rect 3478 1697 3484 1698
rect 3478 1693 3479 1697
rect 3483 1693 3484 1697
rect 3478 1692 3484 1693
rect 3480 1683 3482 1692
rect 3498 1691 3504 1692
rect 3498 1687 3499 1691
rect 3503 1687 3504 1691
rect 3498 1686 3504 1687
rect 3479 1682 3483 1683
rect 3479 1677 3483 1678
rect 3480 1672 3482 1677
rect 3478 1671 3484 1672
rect 3478 1667 3479 1671
rect 3483 1667 3484 1671
rect 3478 1666 3484 1667
rect 3486 1631 3492 1632
rect 3486 1627 3487 1631
rect 3491 1627 3492 1631
rect 3486 1626 3492 1627
rect 3488 1615 3490 1626
rect 3500 1620 3502 1686
rect 3576 1683 3578 1702
rect 3575 1682 3579 1683
rect 3575 1677 3579 1678
rect 3576 1662 3578 1677
rect 3574 1661 3580 1662
rect 3574 1657 3575 1661
rect 3579 1657 3580 1661
rect 3574 1656 3580 1657
rect 3574 1644 3580 1645
rect 3574 1640 3575 1644
rect 3579 1640 3580 1644
rect 3574 1639 3580 1640
rect 3498 1619 3504 1620
rect 3498 1615 3499 1619
rect 3503 1615 3504 1619
rect 3576 1615 3578 1639
rect 3487 1614 3491 1615
rect 3498 1614 3504 1615
rect 3575 1614 3579 1615
rect 3487 1609 3491 1610
rect 3575 1609 3579 1610
rect 3488 1598 3490 1609
rect 3486 1597 3492 1598
rect 3486 1593 3487 1597
rect 3491 1593 3492 1597
rect 3486 1592 3492 1593
rect 3576 1585 3578 1609
rect 3574 1584 3580 1585
rect 3574 1580 3575 1584
rect 3579 1580 3580 1584
rect 3462 1579 3468 1580
rect 3574 1579 3580 1580
rect 3462 1575 3463 1579
rect 3467 1575 3468 1579
rect 3462 1574 3468 1575
rect 3574 1567 3580 1568
rect 3574 1563 3575 1567
rect 3579 1563 3580 1567
rect 3574 1562 3580 1563
rect 3478 1557 3484 1558
rect 3478 1553 3479 1557
rect 3483 1553 3484 1557
rect 3478 1552 3484 1553
rect 3480 1539 3482 1552
rect 3576 1539 3578 1562
rect 3479 1538 3483 1539
rect 3479 1533 3483 1534
rect 3575 1538 3579 1539
rect 3575 1533 3579 1534
rect 3576 1518 3578 1533
rect 3574 1517 3580 1518
rect 3574 1513 3575 1517
rect 3579 1513 3580 1517
rect 3574 1512 3580 1513
rect 3498 1503 3504 1504
rect 3498 1499 3499 1503
rect 3503 1499 3504 1503
rect 3498 1498 3504 1499
rect 3574 1500 3580 1501
rect 3446 1475 3452 1476
rect 3446 1471 3447 1475
rect 3451 1471 3452 1475
rect 3446 1470 3452 1471
rect 3247 1466 3251 1467
rect 3247 1461 3251 1462
rect 3279 1466 3283 1467
rect 3279 1461 3283 1462
rect 3439 1466 3443 1467
rect 3439 1461 3443 1462
rect 3463 1466 3467 1467
rect 3463 1461 3467 1462
rect 3122 1459 3128 1460
rect 3122 1455 3123 1459
rect 3127 1455 3128 1459
rect 3122 1454 3128 1455
rect 3280 1450 3282 1461
rect 3464 1450 3466 1461
rect 3500 1460 3502 1498
rect 3574 1496 3575 1500
rect 3579 1496 3580 1500
rect 3574 1495 3580 1496
rect 3576 1467 3578 1495
rect 3575 1466 3579 1467
rect 3575 1461 3579 1462
rect 3498 1459 3504 1460
rect 3498 1455 3499 1459
rect 3503 1455 3504 1459
rect 3498 1454 3504 1455
rect 2934 1449 2940 1450
rect 2934 1445 2935 1449
rect 2939 1445 2940 1449
rect 2934 1444 2940 1445
rect 3102 1449 3108 1450
rect 3102 1445 3103 1449
rect 3107 1445 3108 1449
rect 3102 1444 3108 1445
rect 3278 1449 3284 1450
rect 3278 1445 3279 1449
rect 3283 1445 3284 1449
rect 3278 1444 3284 1445
rect 3462 1449 3468 1450
rect 3462 1445 3463 1449
rect 3467 1445 3468 1449
rect 3462 1444 3468 1445
rect 3576 1437 3578 1461
rect 3574 1436 3580 1437
rect 2826 1435 2832 1436
rect 2826 1431 2827 1435
rect 2831 1431 2832 1435
rect 3574 1432 3575 1436
rect 3579 1432 3580 1436
rect 3574 1431 3580 1432
rect 2826 1430 2832 1431
rect 2866 1419 2872 1420
rect 2866 1415 2867 1419
rect 2871 1415 2872 1419
rect 2866 1414 2872 1415
rect 3574 1419 3580 1420
rect 3574 1415 3575 1419
rect 3579 1415 3580 1419
rect 3574 1414 3580 1415
rect 2606 1409 2612 1410
rect 2606 1405 2607 1409
rect 2611 1405 2612 1409
rect 2606 1404 2612 1405
rect 2758 1409 2764 1410
rect 2758 1405 2759 1409
rect 2763 1405 2764 1409
rect 2758 1404 2764 1405
rect 2608 1387 2610 1404
rect 2760 1387 2762 1404
rect 2607 1386 2611 1387
rect 2607 1381 2611 1382
rect 2623 1386 2627 1387
rect 2623 1381 2627 1382
rect 2759 1386 2763 1387
rect 2759 1381 2763 1382
rect 2847 1386 2851 1387
rect 2847 1381 2851 1382
rect 2624 1376 2626 1381
rect 2848 1376 2850 1381
rect 2622 1375 2628 1376
rect 2622 1371 2623 1375
rect 2627 1371 2628 1375
rect 2622 1370 2628 1371
rect 2846 1375 2852 1376
rect 2846 1371 2847 1375
rect 2851 1371 2852 1375
rect 2846 1370 2852 1371
rect 2518 1367 2524 1368
rect 2518 1363 2519 1367
rect 2523 1363 2524 1367
rect 2518 1362 2524 1363
rect 2462 1351 2468 1352
rect 2462 1347 2463 1351
rect 2467 1347 2468 1351
rect 2462 1346 2468 1347
rect 2398 1335 2404 1336
rect 2398 1331 2399 1335
rect 2403 1331 2404 1335
rect 2398 1330 2404 1331
rect 2378 1323 2384 1324
rect 2378 1319 2379 1323
rect 2383 1319 2384 1323
rect 2400 1319 2402 1330
rect 2464 1324 2466 1346
rect 2630 1335 2636 1336
rect 2630 1331 2631 1335
rect 2635 1331 2636 1335
rect 2630 1330 2636 1331
rect 2854 1335 2860 1336
rect 2854 1331 2855 1335
rect 2859 1331 2860 1335
rect 2854 1330 2860 1331
rect 2462 1323 2468 1324
rect 2462 1319 2463 1323
rect 2467 1319 2468 1323
rect 2632 1319 2634 1330
rect 2682 1323 2688 1324
rect 2682 1319 2683 1323
rect 2687 1319 2688 1323
rect 2856 1319 2858 1330
rect 2868 1324 2870 1414
rect 2926 1409 2932 1410
rect 2926 1405 2927 1409
rect 2931 1405 2932 1409
rect 2926 1404 2932 1405
rect 3094 1409 3100 1410
rect 3094 1405 3095 1409
rect 3099 1405 3100 1409
rect 3094 1404 3100 1405
rect 3270 1409 3276 1410
rect 3270 1405 3271 1409
rect 3275 1405 3276 1409
rect 3270 1404 3276 1405
rect 3454 1409 3460 1410
rect 3454 1405 3455 1409
rect 3459 1405 3460 1409
rect 3454 1404 3460 1405
rect 2928 1387 2930 1404
rect 3096 1387 3098 1404
rect 3272 1387 3274 1404
rect 3456 1387 3458 1404
rect 3498 1403 3504 1404
rect 3498 1399 3499 1403
rect 3503 1399 3504 1403
rect 3498 1398 3504 1399
rect 2927 1386 2931 1387
rect 2927 1381 2931 1382
rect 3063 1386 3067 1387
rect 3063 1381 3067 1382
rect 3095 1386 3099 1387
rect 3095 1381 3099 1382
rect 3271 1386 3275 1387
rect 3271 1381 3275 1382
rect 3455 1386 3459 1387
rect 3455 1381 3459 1382
rect 3479 1386 3483 1387
rect 3479 1381 3483 1382
rect 3064 1376 3066 1381
rect 3272 1376 3274 1381
rect 3480 1376 3482 1381
rect 3062 1375 3068 1376
rect 3062 1371 3063 1375
rect 3067 1371 3068 1375
rect 3062 1370 3068 1371
rect 3270 1375 3276 1376
rect 3270 1371 3271 1375
rect 3275 1371 3276 1375
rect 3270 1370 3276 1371
rect 3478 1375 3484 1376
rect 3478 1371 3479 1375
rect 3483 1371 3484 1375
rect 3478 1370 3484 1371
rect 2970 1367 2976 1368
rect 2970 1363 2971 1367
rect 2975 1363 2976 1367
rect 2970 1362 2976 1363
rect 2866 1323 2872 1324
rect 2866 1319 2867 1323
rect 2871 1319 2872 1323
rect 1863 1318 1867 1319
rect 535 1314 539 1315
rect 535 1309 539 1310
rect 543 1314 547 1315
rect 543 1309 547 1310
rect 631 1314 635 1315
rect 631 1309 635 1310
rect 719 1314 723 1315
rect 719 1309 723 1310
rect 735 1314 739 1315
rect 794 1314 800 1315
rect 831 1314 835 1315
rect 735 1309 739 1310
rect 831 1309 835 1310
rect 855 1314 859 1315
rect 898 1314 904 1315
rect 967 1314 971 1315
rect 855 1309 859 1310
rect 967 1309 971 1310
rect 991 1314 995 1315
rect 1026 1314 1032 1315
rect 1135 1314 1139 1315
rect 991 1309 995 1310
rect 506 1307 512 1308
rect 506 1303 507 1307
rect 511 1303 512 1307
rect 506 1302 512 1303
rect 544 1298 546 1309
rect 632 1298 634 1309
rect 720 1298 722 1309
rect 832 1298 834 1309
rect 968 1298 970 1309
rect 454 1297 460 1298
rect 454 1293 455 1297
rect 459 1293 460 1297
rect 454 1292 460 1293
rect 542 1297 548 1298
rect 542 1293 543 1297
rect 547 1293 548 1297
rect 542 1292 548 1293
rect 630 1297 636 1298
rect 630 1293 631 1297
rect 635 1293 636 1297
rect 630 1292 636 1293
rect 718 1297 724 1298
rect 718 1293 719 1297
rect 723 1293 724 1297
rect 718 1292 724 1293
rect 830 1297 836 1298
rect 830 1293 831 1297
rect 835 1293 836 1297
rect 830 1292 836 1293
rect 966 1297 972 1298
rect 966 1293 967 1297
rect 971 1293 972 1297
rect 966 1292 972 1293
rect 110 1284 116 1285
rect 1028 1284 1030 1314
rect 1135 1309 1139 1310
rect 1287 1314 1291 1315
rect 1287 1309 1291 1310
rect 1327 1314 1331 1315
rect 1327 1309 1331 1310
rect 1439 1314 1443 1315
rect 1450 1314 1456 1315
rect 1535 1314 1539 1315
rect 1439 1309 1443 1310
rect 1535 1309 1539 1310
rect 1599 1314 1603 1315
rect 1718 1314 1724 1315
rect 1735 1314 1739 1315
rect 1599 1309 1603 1310
rect 1735 1309 1739 1310
rect 1823 1314 1827 1315
rect 1863 1313 1867 1314
rect 1895 1318 1899 1319
rect 1906 1318 1912 1319
rect 1927 1318 1931 1319
rect 1895 1313 1899 1314
rect 1823 1309 1827 1310
rect 1058 1307 1064 1308
rect 1058 1303 1059 1307
rect 1063 1303 1064 1307
rect 1058 1302 1064 1303
rect 110 1280 111 1284
rect 115 1280 116 1284
rect 110 1279 116 1280
rect 1026 1283 1032 1284
rect 1026 1279 1027 1283
rect 1031 1279 1032 1283
rect 1060 1280 1062 1302
rect 1136 1298 1138 1309
rect 1230 1307 1236 1308
rect 1230 1303 1231 1307
rect 1235 1303 1236 1307
rect 1230 1302 1236 1303
rect 1134 1297 1140 1298
rect 1134 1293 1135 1297
rect 1139 1293 1140 1297
rect 1134 1292 1140 1293
rect 1232 1280 1234 1302
rect 1328 1298 1330 1309
rect 1394 1307 1400 1308
rect 1394 1303 1395 1307
rect 1399 1303 1400 1307
rect 1394 1302 1400 1303
rect 1326 1297 1332 1298
rect 1326 1293 1327 1297
rect 1331 1293 1332 1297
rect 1326 1292 1332 1293
rect 1396 1280 1398 1302
rect 1536 1298 1538 1309
rect 1542 1307 1548 1308
rect 1542 1303 1543 1307
rect 1547 1303 1548 1307
rect 1542 1302 1548 1303
rect 1534 1297 1540 1298
rect 1534 1293 1535 1297
rect 1539 1293 1540 1297
rect 1534 1292 1540 1293
rect 1026 1278 1032 1279
rect 1058 1279 1064 1280
rect 1058 1275 1059 1279
rect 1063 1275 1064 1279
rect 1058 1274 1064 1275
rect 1230 1279 1236 1280
rect 1230 1275 1231 1279
rect 1235 1275 1236 1279
rect 1230 1274 1236 1275
rect 1394 1279 1400 1280
rect 1394 1275 1395 1279
rect 1399 1275 1400 1279
rect 1394 1274 1400 1275
rect 110 1267 116 1268
rect 110 1263 111 1267
rect 115 1263 116 1267
rect 110 1262 116 1263
rect 830 1267 836 1268
rect 830 1263 831 1267
rect 835 1263 836 1267
rect 830 1262 836 1263
rect 112 1247 114 1262
rect 446 1257 452 1258
rect 446 1253 447 1257
rect 451 1253 452 1257
rect 446 1252 452 1253
rect 534 1257 540 1258
rect 534 1253 535 1257
rect 539 1253 540 1257
rect 534 1252 540 1253
rect 622 1257 628 1258
rect 622 1253 623 1257
rect 627 1253 628 1257
rect 622 1252 628 1253
rect 710 1257 716 1258
rect 710 1253 711 1257
rect 715 1253 716 1257
rect 710 1252 716 1253
rect 822 1257 828 1258
rect 822 1253 823 1257
rect 827 1253 828 1257
rect 822 1252 828 1253
rect 448 1247 450 1252
rect 536 1247 538 1252
rect 624 1247 626 1252
rect 712 1247 714 1252
rect 824 1247 826 1252
rect 111 1246 115 1247
rect 111 1241 115 1242
rect 447 1246 451 1247
rect 447 1241 451 1242
rect 535 1246 539 1247
rect 535 1241 539 1242
rect 543 1246 547 1247
rect 543 1241 547 1242
rect 623 1246 627 1247
rect 623 1241 627 1242
rect 631 1246 635 1247
rect 631 1241 635 1242
rect 711 1246 715 1247
rect 711 1241 715 1242
rect 719 1246 723 1247
rect 719 1241 723 1242
rect 807 1246 811 1247
rect 807 1241 811 1242
rect 823 1246 827 1247
rect 823 1241 827 1242
rect 112 1226 114 1241
rect 544 1236 546 1241
rect 632 1236 634 1241
rect 720 1236 722 1241
rect 808 1236 810 1241
rect 542 1235 548 1236
rect 542 1231 543 1235
rect 547 1231 548 1235
rect 542 1230 548 1231
rect 630 1235 636 1236
rect 630 1231 631 1235
rect 635 1231 636 1235
rect 630 1230 636 1231
rect 718 1235 724 1236
rect 718 1231 719 1235
rect 723 1231 724 1235
rect 718 1230 724 1231
rect 806 1235 812 1236
rect 806 1231 807 1235
rect 811 1231 812 1235
rect 806 1230 812 1231
rect 698 1227 704 1228
rect 110 1225 116 1226
rect 110 1221 111 1225
rect 115 1221 116 1225
rect 698 1223 699 1227
rect 703 1223 704 1227
rect 698 1222 704 1223
rect 110 1220 116 1221
rect 110 1208 116 1209
rect 110 1204 111 1208
rect 115 1204 116 1208
rect 110 1203 116 1204
rect 112 1171 114 1203
rect 550 1195 556 1196
rect 550 1191 551 1195
rect 555 1191 556 1195
rect 550 1190 556 1191
rect 638 1195 644 1196
rect 638 1191 639 1195
rect 643 1191 644 1195
rect 638 1190 644 1191
rect 552 1171 554 1190
rect 640 1171 642 1190
rect 700 1176 702 1222
rect 726 1195 732 1196
rect 726 1191 727 1195
rect 731 1191 732 1195
rect 726 1190 732 1191
rect 814 1195 820 1196
rect 814 1191 815 1195
rect 819 1191 820 1195
rect 814 1190 820 1191
rect 698 1175 704 1176
rect 698 1171 699 1175
rect 703 1171 704 1175
rect 728 1171 730 1190
rect 816 1171 818 1190
rect 832 1188 834 1262
rect 958 1257 964 1258
rect 958 1253 959 1257
rect 963 1253 964 1257
rect 958 1252 964 1253
rect 1126 1257 1132 1258
rect 1126 1253 1127 1257
rect 1131 1253 1132 1257
rect 1126 1252 1132 1253
rect 1318 1257 1324 1258
rect 1318 1253 1319 1257
rect 1323 1253 1324 1257
rect 1318 1252 1324 1253
rect 1526 1257 1532 1258
rect 1526 1253 1527 1257
rect 1531 1253 1532 1257
rect 1526 1252 1532 1253
rect 960 1247 962 1252
rect 1128 1247 1130 1252
rect 1320 1247 1322 1252
rect 1528 1247 1530 1252
rect 895 1246 899 1247
rect 895 1241 899 1242
rect 959 1246 963 1247
rect 959 1241 963 1242
rect 991 1246 995 1247
rect 991 1241 995 1242
rect 1095 1246 1099 1247
rect 1095 1241 1099 1242
rect 1127 1246 1131 1247
rect 1127 1241 1131 1242
rect 1207 1246 1211 1247
rect 1207 1241 1211 1242
rect 1319 1246 1323 1247
rect 1319 1241 1323 1242
rect 1335 1246 1339 1247
rect 1335 1241 1339 1242
rect 1471 1246 1475 1247
rect 1471 1241 1475 1242
rect 1527 1246 1531 1247
rect 1527 1241 1531 1242
rect 896 1236 898 1241
rect 992 1236 994 1241
rect 1096 1236 1098 1241
rect 1208 1236 1210 1241
rect 1336 1236 1338 1241
rect 1472 1236 1474 1241
rect 894 1235 900 1236
rect 894 1231 895 1235
rect 899 1231 900 1235
rect 894 1230 900 1231
rect 990 1235 996 1236
rect 990 1231 991 1235
rect 995 1231 996 1235
rect 990 1230 996 1231
rect 1094 1235 1100 1236
rect 1094 1231 1095 1235
rect 1099 1231 1100 1235
rect 1094 1230 1100 1231
rect 1206 1235 1212 1236
rect 1206 1231 1207 1235
rect 1211 1231 1212 1235
rect 1206 1230 1212 1231
rect 1334 1235 1340 1236
rect 1334 1231 1335 1235
rect 1339 1231 1340 1235
rect 1334 1230 1340 1231
rect 1470 1235 1476 1236
rect 1470 1231 1471 1235
rect 1475 1231 1476 1235
rect 1470 1230 1476 1231
rect 1544 1228 1546 1302
rect 1736 1298 1738 1309
rect 1734 1297 1740 1298
rect 1734 1293 1735 1297
rect 1739 1293 1740 1297
rect 1734 1292 1740 1293
rect 1824 1285 1826 1309
rect 1864 1289 1866 1313
rect 1862 1288 1868 1289
rect 1822 1284 1828 1285
rect 1822 1280 1823 1284
rect 1827 1280 1828 1284
rect 1862 1284 1863 1288
rect 1867 1284 1868 1288
rect 1908 1284 1910 1318
rect 1927 1313 1931 1314
rect 2111 1318 2115 1319
rect 2111 1313 2115 1314
rect 2151 1318 2155 1319
rect 2151 1313 2155 1314
rect 2287 1318 2291 1319
rect 2378 1318 2384 1319
rect 2399 1318 2403 1319
rect 2287 1313 2291 1314
rect 2399 1313 2403 1314
rect 2455 1318 2459 1319
rect 2462 1318 2468 1319
rect 2623 1318 2627 1319
rect 2455 1313 2459 1314
rect 2623 1313 2627 1314
rect 2631 1318 2635 1319
rect 2682 1318 2688 1319
rect 2791 1318 2795 1319
rect 2631 1313 2635 1314
rect 1928 1302 1930 1313
rect 2030 1311 2036 1312
rect 2030 1307 2031 1311
rect 2035 1307 2036 1311
rect 2030 1306 2036 1307
rect 1926 1301 1932 1302
rect 1926 1297 1927 1301
rect 1931 1297 1932 1301
rect 1926 1296 1932 1297
rect 2032 1284 2034 1306
rect 2112 1302 2114 1313
rect 2230 1311 2236 1312
rect 2230 1307 2231 1311
rect 2235 1307 2236 1311
rect 2230 1306 2236 1307
rect 2110 1301 2116 1302
rect 2110 1297 2111 1301
rect 2115 1297 2116 1301
rect 2110 1296 2116 1297
rect 1862 1283 1868 1284
rect 1906 1283 1912 1284
rect 1822 1279 1828 1280
rect 1906 1279 1907 1283
rect 1911 1279 1912 1283
rect 1906 1278 1912 1279
rect 2030 1283 2036 1284
rect 2030 1279 2031 1283
rect 2035 1279 2036 1283
rect 2030 1278 2036 1279
rect 1862 1271 1868 1272
rect 1626 1267 1632 1268
rect 1626 1263 1627 1267
rect 1631 1263 1632 1267
rect 1626 1262 1632 1263
rect 1822 1267 1828 1268
rect 1822 1263 1823 1267
rect 1827 1263 1828 1267
rect 1862 1267 1863 1271
rect 1867 1267 1868 1271
rect 1862 1266 1868 1267
rect 1822 1262 1828 1263
rect 1607 1246 1611 1247
rect 1607 1241 1611 1242
rect 1608 1236 1610 1241
rect 1606 1235 1612 1236
rect 1606 1231 1607 1235
rect 1611 1231 1612 1235
rect 1606 1230 1612 1231
rect 874 1227 880 1228
rect 874 1223 875 1227
rect 879 1223 880 1227
rect 874 1222 880 1223
rect 1542 1227 1548 1228
rect 1542 1223 1543 1227
rect 1547 1223 1548 1227
rect 1542 1222 1548 1223
rect 826 1187 834 1188
rect 826 1183 827 1187
rect 831 1184 834 1187
rect 831 1183 832 1184
rect 826 1182 832 1183
rect 876 1176 878 1222
rect 902 1195 908 1196
rect 902 1191 903 1195
rect 907 1191 908 1195
rect 902 1190 908 1191
rect 998 1195 1004 1196
rect 998 1191 999 1195
rect 1003 1191 1004 1195
rect 998 1190 1004 1191
rect 1102 1195 1108 1196
rect 1102 1191 1103 1195
rect 1107 1191 1108 1195
rect 1102 1190 1108 1191
rect 1214 1195 1220 1196
rect 1214 1191 1215 1195
rect 1219 1191 1220 1195
rect 1214 1190 1220 1191
rect 1342 1195 1348 1196
rect 1342 1191 1343 1195
rect 1347 1191 1348 1195
rect 1342 1190 1348 1191
rect 1478 1195 1484 1196
rect 1478 1191 1479 1195
rect 1483 1191 1484 1195
rect 1478 1190 1484 1191
rect 1614 1195 1620 1196
rect 1614 1191 1615 1195
rect 1619 1191 1620 1195
rect 1614 1190 1620 1191
rect 874 1175 880 1176
rect 874 1171 875 1175
rect 879 1171 880 1175
rect 904 1171 906 1190
rect 1000 1171 1002 1190
rect 1010 1183 1016 1184
rect 1010 1179 1011 1183
rect 1015 1179 1016 1183
rect 1010 1178 1016 1179
rect 111 1170 115 1171
rect 111 1165 115 1166
rect 359 1170 363 1171
rect 359 1165 363 1166
rect 471 1170 475 1171
rect 471 1165 475 1166
rect 551 1170 555 1171
rect 551 1165 555 1166
rect 591 1170 595 1171
rect 591 1165 595 1166
rect 639 1170 643 1171
rect 698 1170 704 1171
rect 711 1170 715 1171
rect 639 1165 643 1166
rect 711 1165 715 1166
rect 727 1170 731 1171
rect 727 1165 731 1166
rect 815 1170 819 1171
rect 815 1165 819 1166
rect 831 1170 835 1171
rect 874 1170 880 1171
rect 903 1170 907 1171
rect 831 1165 835 1166
rect 903 1165 907 1166
rect 951 1170 955 1171
rect 951 1165 955 1166
rect 999 1170 1003 1171
rect 999 1165 1003 1166
rect 112 1141 114 1165
rect 360 1154 362 1165
rect 414 1163 420 1164
rect 414 1159 415 1163
rect 419 1159 420 1163
rect 414 1158 420 1159
rect 358 1153 364 1154
rect 358 1149 359 1153
rect 363 1149 364 1153
rect 358 1148 364 1149
rect 416 1141 418 1158
rect 472 1154 474 1165
rect 592 1154 594 1165
rect 712 1154 714 1165
rect 770 1163 776 1164
rect 770 1159 771 1163
rect 775 1159 776 1163
rect 770 1158 776 1159
rect 470 1153 476 1154
rect 470 1149 471 1153
rect 475 1149 476 1153
rect 470 1148 476 1149
rect 590 1153 596 1154
rect 590 1149 591 1153
rect 595 1149 596 1153
rect 590 1148 596 1149
rect 710 1153 716 1154
rect 710 1149 711 1153
rect 715 1149 716 1153
rect 710 1148 716 1149
rect 110 1140 116 1141
rect 110 1136 111 1140
rect 115 1136 116 1140
rect 110 1135 116 1136
rect 415 1140 419 1141
rect 772 1140 774 1158
rect 832 1154 834 1165
rect 952 1154 954 1165
rect 830 1153 836 1154
rect 830 1149 831 1153
rect 835 1149 836 1153
rect 830 1148 836 1149
rect 950 1153 956 1154
rect 950 1149 951 1153
rect 955 1149 956 1153
rect 950 1148 956 1149
rect 779 1140 783 1141
rect 1012 1140 1014 1178
rect 1104 1171 1106 1190
rect 1216 1171 1218 1190
rect 1344 1171 1346 1190
rect 1480 1171 1482 1190
rect 1616 1171 1618 1190
rect 1628 1184 1630 1262
rect 1726 1257 1732 1258
rect 1726 1253 1727 1257
rect 1731 1253 1732 1257
rect 1726 1252 1732 1253
rect 1728 1247 1730 1252
rect 1824 1247 1826 1262
rect 1727 1246 1731 1247
rect 1727 1241 1731 1242
rect 1823 1246 1827 1247
rect 1864 1243 1866 1266
rect 1918 1261 1924 1262
rect 1918 1257 1919 1261
rect 1923 1257 1924 1261
rect 1918 1256 1924 1257
rect 2102 1261 2108 1262
rect 2102 1257 2103 1261
rect 2107 1257 2108 1261
rect 2102 1256 2108 1257
rect 1920 1243 1922 1256
rect 2104 1243 2106 1256
rect 1823 1241 1827 1242
rect 1863 1242 1867 1243
rect 1728 1236 1730 1241
rect 1726 1235 1732 1236
rect 1726 1231 1727 1235
rect 1731 1231 1732 1235
rect 1726 1230 1732 1231
rect 1824 1226 1826 1241
rect 1863 1237 1867 1238
rect 1919 1242 1923 1243
rect 1919 1237 1923 1238
rect 2103 1242 2107 1243
rect 2103 1237 2107 1238
rect 2143 1242 2147 1243
rect 2143 1237 2147 1238
rect 1822 1225 1828 1226
rect 1822 1221 1823 1225
rect 1827 1221 1828 1225
rect 1864 1222 1866 1237
rect 2144 1232 2146 1237
rect 2142 1231 2148 1232
rect 2142 1227 2143 1231
rect 2147 1227 2148 1231
rect 2142 1226 2148 1227
rect 2232 1224 2234 1306
rect 2288 1302 2290 1313
rect 2456 1302 2458 1313
rect 2624 1302 2626 1313
rect 2286 1301 2292 1302
rect 2286 1297 2287 1301
rect 2291 1297 2292 1301
rect 2286 1296 2292 1297
rect 2454 1301 2460 1302
rect 2454 1297 2455 1301
rect 2459 1297 2460 1301
rect 2454 1296 2460 1297
rect 2622 1301 2628 1302
rect 2622 1297 2623 1301
rect 2627 1297 2628 1301
rect 2622 1296 2628 1297
rect 2684 1288 2686 1318
rect 2791 1313 2795 1314
rect 2855 1318 2859 1319
rect 2866 1318 2872 1319
rect 2959 1318 2963 1319
rect 2855 1313 2859 1314
rect 2959 1313 2963 1314
rect 2718 1311 2724 1312
rect 2718 1307 2719 1311
rect 2723 1307 2724 1311
rect 2718 1306 2724 1307
rect 2682 1287 2688 1288
rect 2682 1283 2683 1287
rect 2687 1283 2688 1287
rect 2720 1284 2722 1306
rect 2792 1302 2794 1313
rect 2814 1311 2820 1312
rect 2814 1307 2815 1311
rect 2819 1307 2820 1311
rect 2814 1306 2820 1307
rect 2790 1301 2796 1302
rect 2790 1297 2791 1301
rect 2795 1297 2796 1301
rect 2790 1296 2796 1297
rect 2682 1282 2688 1283
rect 2718 1283 2724 1284
rect 2718 1279 2719 1283
rect 2723 1279 2724 1283
rect 2718 1278 2724 1279
rect 2278 1261 2284 1262
rect 2278 1257 2279 1261
rect 2283 1257 2284 1261
rect 2278 1256 2284 1257
rect 2446 1261 2452 1262
rect 2446 1257 2447 1261
rect 2451 1257 2452 1261
rect 2446 1256 2452 1257
rect 2614 1261 2620 1262
rect 2614 1257 2615 1261
rect 2619 1257 2620 1261
rect 2614 1256 2620 1257
rect 2782 1261 2788 1262
rect 2782 1257 2783 1261
rect 2787 1257 2788 1261
rect 2782 1256 2788 1257
rect 2280 1243 2282 1256
rect 2448 1243 2450 1256
rect 2506 1255 2512 1256
rect 2506 1251 2507 1255
rect 2511 1251 2512 1255
rect 2506 1250 2512 1251
rect 2279 1242 2283 1243
rect 2279 1237 2283 1238
rect 2319 1242 2323 1243
rect 2319 1237 2323 1238
rect 2447 1242 2451 1243
rect 2447 1237 2451 1238
rect 2487 1242 2491 1243
rect 2487 1237 2491 1238
rect 2320 1232 2322 1237
rect 2488 1232 2490 1237
rect 2318 1231 2324 1232
rect 2318 1227 2319 1231
rect 2323 1227 2324 1231
rect 2318 1226 2324 1227
rect 2486 1231 2492 1232
rect 2486 1227 2487 1231
rect 2491 1227 2492 1231
rect 2486 1226 2492 1227
rect 2230 1223 2236 1224
rect 1822 1220 1828 1221
rect 1862 1221 1868 1222
rect 1862 1217 1863 1221
rect 1867 1217 1868 1221
rect 2230 1219 2231 1223
rect 2235 1219 2236 1223
rect 2230 1218 2236 1219
rect 1862 1216 1868 1217
rect 1814 1211 1820 1212
rect 1814 1207 1815 1211
rect 1819 1207 1820 1211
rect 1814 1206 1820 1207
rect 1822 1208 1828 1209
rect 1734 1195 1740 1196
rect 1734 1191 1735 1195
rect 1739 1191 1740 1195
rect 1734 1190 1740 1191
rect 1626 1183 1632 1184
rect 1626 1179 1627 1183
rect 1631 1179 1632 1183
rect 1626 1178 1632 1179
rect 1736 1171 1738 1190
rect 1063 1170 1067 1171
rect 1063 1165 1067 1166
rect 1103 1170 1107 1171
rect 1103 1165 1107 1166
rect 1183 1170 1187 1171
rect 1183 1165 1187 1166
rect 1215 1170 1219 1171
rect 1215 1165 1219 1166
rect 1303 1170 1307 1171
rect 1303 1165 1307 1166
rect 1343 1170 1347 1171
rect 1343 1165 1347 1166
rect 1423 1170 1427 1171
rect 1423 1165 1427 1166
rect 1479 1170 1483 1171
rect 1479 1165 1483 1166
rect 1615 1170 1619 1171
rect 1615 1165 1619 1166
rect 1735 1170 1739 1171
rect 1816 1168 1818 1206
rect 1822 1204 1823 1208
rect 1827 1204 1828 1208
rect 2210 1207 2216 1208
rect 1822 1203 1828 1204
rect 1862 1204 1868 1205
rect 1824 1171 1826 1203
rect 1862 1200 1863 1204
rect 1867 1200 1868 1204
rect 2210 1203 2211 1207
rect 2215 1203 2216 1207
rect 2210 1202 2216 1203
rect 1862 1199 1868 1200
rect 1864 1175 1866 1199
rect 2150 1191 2156 1192
rect 2150 1187 2151 1191
rect 2155 1187 2156 1191
rect 2150 1186 2156 1187
rect 2152 1175 2154 1186
rect 2212 1180 2214 1202
rect 2326 1191 2332 1192
rect 2326 1187 2327 1191
rect 2331 1187 2332 1191
rect 2326 1186 2332 1187
rect 2494 1191 2500 1192
rect 2494 1187 2495 1191
rect 2499 1187 2500 1191
rect 2494 1186 2500 1187
rect 2210 1179 2216 1180
rect 2210 1175 2211 1179
rect 2215 1175 2216 1179
rect 2328 1175 2330 1186
rect 2354 1179 2360 1180
rect 2354 1175 2355 1179
rect 2359 1175 2360 1179
rect 2496 1175 2498 1186
rect 2508 1180 2510 1250
rect 2616 1243 2618 1256
rect 2784 1243 2786 1256
rect 2615 1242 2619 1243
rect 2615 1237 2619 1238
rect 2655 1242 2659 1243
rect 2655 1237 2659 1238
rect 2783 1242 2787 1243
rect 2783 1237 2787 1238
rect 2656 1232 2658 1237
rect 2654 1231 2660 1232
rect 2654 1227 2655 1231
rect 2659 1227 2660 1231
rect 2654 1226 2660 1227
rect 2816 1224 2818 1306
rect 2960 1302 2962 1313
rect 2972 1312 2974 1362
rect 3070 1335 3076 1336
rect 3070 1331 3071 1335
rect 3075 1331 3076 1335
rect 3070 1330 3076 1331
rect 3278 1335 3284 1336
rect 3278 1331 3279 1335
rect 3283 1331 3284 1335
rect 3278 1330 3284 1331
rect 3486 1335 3492 1336
rect 3486 1331 3487 1335
rect 3491 1331 3492 1335
rect 3486 1330 3492 1331
rect 3072 1319 3074 1330
rect 3280 1319 3282 1330
rect 3418 1323 3424 1324
rect 3418 1319 3419 1323
rect 3423 1319 3424 1323
rect 3488 1319 3490 1330
rect 3500 1324 3502 1398
rect 3576 1387 3578 1414
rect 3575 1386 3579 1387
rect 3575 1381 3579 1382
rect 3576 1366 3578 1381
rect 3574 1365 3580 1366
rect 3574 1361 3575 1365
rect 3579 1361 3580 1365
rect 3574 1360 3580 1361
rect 3574 1348 3580 1349
rect 3574 1344 3575 1348
rect 3579 1344 3580 1348
rect 3574 1343 3580 1344
rect 3498 1323 3504 1324
rect 3498 1319 3499 1323
rect 3503 1319 3504 1323
rect 3576 1319 3578 1343
rect 3071 1318 3075 1319
rect 3071 1313 3075 1314
rect 3135 1318 3139 1319
rect 3135 1313 3139 1314
rect 3279 1318 3283 1319
rect 3279 1313 3283 1314
rect 3319 1318 3323 1319
rect 3418 1318 3424 1319
rect 3487 1318 3491 1319
rect 3498 1318 3504 1319
rect 3575 1318 3579 1319
rect 3319 1313 3323 1314
rect 2970 1311 2976 1312
rect 2970 1307 2971 1311
rect 2975 1307 2976 1311
rect 2970 1306 2976 1307
rect 3136 1302 3138 1313
rect 3320 1302 3322 1313
rect 2958 1301 2964 1302
rect 2958 1297 2959 1301
rect 2963 1297 2964 1301
rect 2958 1296 2964 1297
rect 3134 1301 3140 1302
rect 3134 1297 3135 1301
rect 3139 1297 3140 1301
rect 3134 1296 3140 1297
rect 3318 1301 3324 1302
rect 3318 1297 3319 1301
rect 3323 1297 3324 1301
rect 3318 1296 3324 1297
rect 2950 1261 2956 1262
rect 2950 1257 2951 1261
rect 2955 1257 2956 1261
rect 2950 1256 2956 1257
rect 3126 1261 3132 1262
rect 3126 1257 3127 1261
rect 3131 1257 3132 1261
rect 3126 1256 3132 1257
rect 3310 1261 3316 1262
rect 3310 1257 3311 1261
rect 3315 1257 3316 1261
rect 3310 1256 3316 1257
rect 2952 1243 2954 1256
rect 3128 1243 3130 1256
rect 3312 1243 3314 1256
rect 3346 1255 3352 1256
rect 3346 1251 3347 1255
rect 3351 1251 3352 1255
rect 3346 1250 3352 1251
rect 2823 1242 2827 1243
rect 2823 1237 2827 1238
rect 2951 1242 2955 1243
rect 2951 1237 2955 1238
rect 2991 1242 2995 1243
rect 2991 1237 2995 1238
rect 3127 1242 3131 1243
rect 3127 1237 3131 1238
rect 3159 1242 3163 1243
rect 3159 1237 3163 1238
rect 3311 1242 3315 1243
rect 3311 1237 3315 1238
rect 3327 1242 3331 1243
rect 3327 1237 3331 1238
rect 2824 1232 2826 1237
rect 2992 1232 2994 1237
rect 3160 1232 3162 1237
rect 3328 1232 3330 1237
rect 2822 1231 2828 1232
rect 2822 1227 2823 1231
rect 2827 1227 2828 1231
rect 2822 1226 2828 1227
rect 2990 1231 2996 1232
rect 2990 1227 2991 1231
rect 2995 1227 2996 1231
rect 2990 1226 2996 1227
rect 3158 1231 3164 1232
rect 3158 1227 3159 1231
rect 3163 1227 3164 1231
rect 3158 1226 3164 1227
rect 3326 1231 3332 1232
rect 3326 1227 3327 1231
rect 3331 1227 3332 1231
rect 3326 1226 3332 1227
rect 2814 1223 2820 1224
rect 2814 1219 2815 1223
rect 2819 1219 2820 1223
rect 2814 1218 2820 1219
rect 3058 1223 3064 1224
rect 3058 1219 3059 1223
rect 3063 1219 3064 1223
rect 3058 1218 3064 1219
rect 2798 1207 2804 1208
rect 2798 1203 2799 1207
rect 2803 1203 2804 1207
rect 2798 1202 2804 1203
rect 2662 1191 2668 1192
rect 2662 1187 2663 1191
rect 2667 1187 2668 1191
rect 2662 1186 2668 1187
rect 2506 1179 2512 1180
rect 2506 1175 2507 1179
rect 2511 1175 2512 1179
rect 2664 1175 2666 1186
rect 2800 1180 2802 1202
rect 2830 1191 2836 1192
rect 2830 1187 2831 1191
rect 2835 1187 2836 1191
rect 2830 1186 2836 1187
rect 2998 1191 3004 1192
rect 2998 1187 2999 1191
rect 3003 1187 3004 1191
rect 2998 1186 3004 1187
rect 2682 1179 2688 1180
rect 2682 1175 2683 1179
rect 2687 1175 2688 1179
rect 2798 1179 2804 1180
rect 2798 1175 2799 1179
rect 2803 1175 2804 1179
rect 2832 1175 2834 1186
rect 3000 1175 3002 1186
rect 3060 1180 3062 1218
rect 3150 1207 3156 1208
rect 3150 1203 3151 1207
rect 3155 1203 3156 1207
rect 3150 1202 3156 1203
rect 3226 1207 3232 1208
rect 3226 1203 3227 1207
rect 3231 1203 3232 1207
rect 3226 1202 3232 1203
rect 3058 1179 3064 1180
rect 3058 1175 3059 1179
rect 3063 1175 3064 1179
rect 1863 1174 1867 1175
rect 1823 1170 1827 1171
rect 1735 1165 1739 1166
rect 1814 1167 1820 1168
rect 1018 1163 1024 1164
rect 1018 1159 1019 1163
rect 1023 1159 1024 1163
rect 1018 1158 1024 1159
rect 415 1135 419 1136
rect 770 1139 776 1140
rect 770 1135 771 1139
rect 775 1135 776 1139
rect 1010 1139 1016 1140
rect 770 1134 776 1135
rect 778 1135 784 1136
rect 778 1131 779 1135
rect 783 1131 784 1135
rect 1010 1135 1011 1139
rect 1015 1135 1016 1139
rect 1020 1136 1022 1158
rect 1064 1154 1066 1165
rect 1134 1163 1140 1164
rect 1134 1159 1135 1163
rect 1139 1159 1140 1163
rect 1134 1158 1140 1159
rect 1062 1153 1068 1154
rect 1062 1149 1063 1153
rect 1067 1149 1068 1153
rect 1062 1148 1068 1149
rect 1136 1136 1138 1158
rect 1184 1154 1186 1165
rect 1304 1154 1306 1165
rect 1322 1163 1328 1164
rect 1322 1159 1323 1163
rect 1327 1159 1328 1163
rect 1322 1158 1328 1159
rect 1182 1153 1188 1154
rect 1182 1149 1183 1153
rect 1187 1149 1188 1153
rect 1182 1148 1188 1149
rect 1302 1153 1308 1154
rect 1302 1149 1303 1153
rect 1307 1149 1308 1153
rect 1302 1148 1308 1149
rect 1010 1134 1016 1135
rect 1018 1135 1024 1136
rect 778 1130 784 1131
rect 1018 1131 1019 1135
rect 1023 1131 1024 1135
rect 1018 1130 1024 1131
rect 1134 1135 1140 1136
rect 1134 1131 1135 1135
rect 1139 1131 1140 1135
rect 1134 1130 1140 1131
rect 110 1123 116 1124
rect 110 1119 111 1123
rect 115 1119 116 1123
rect 110 1118 116 1119
rect 112 1099 114 1118
rect 350 1113 356 1114
rect 350 1109 351 1113
rect 355 1109 356 1113
rect 350 1108 356 1109
rect 462 1113 468 1114
rect 462 1109 463 1113
rect 467 1109 468 1113
rect 462 1108 468 1109
rect 582 1113 588 1114
rect 582 1109 583 1113
rect 587 1109 588 1113
rect 582 1108 588 1109
rect 702 1113 708 1114
rect 702 1109 703 1113
rect 707 1109 708 1113
rect 702 1108 708 1109
rect 822 1113 828 1114
rect 822 1109 823 1113
rect 827 1109 828 1113
rect 822 1108 828 1109
rect 942 1113 948 1114
rect 942 1109 943 1113
rect 947 1109 948 1113
rect 942 1108 948 1109
rect 1054 1113 1060 1114
rect 1054 1109 1055 1113
rect 1059 1109 1060 1113
rect 1054 1108 1060 1109
rect 1174 1113 1180 1114
rect 1174 1109 1175 1113
rect 1179 1109 1180 1113
rect 1174 1108 1180 1109
rect 1294 1113 1300 1114
rect 1294 1109 1295 1113
rect 1299 1109 1300 1113
rect 1294 1108 1300 1109
rect 352 1099 354 1108
rect 464 1099 466 1108
rect 584 1099 586 1108
rect 630 1107 636 1108
rect 630 1103 631 1107
rect 635 1103 636 1107
rect 630 1102 636 1103
rect 111 1098 115 1099
rect 111 1093 115 1094
rect 143 1098 147 1099
rect 143 1093 147 1094
rect 287 1098 291 1099
rect 287 1093 291 1094
rect 351 1098 355 1099
rect 351 1093 355 1094
rect 447 1098 451 1099
rect 447 1093 451 1094
rect 463 1098 467 1099
rect 463 1093 467 1094
rect 583 1098 587 1099
rect 583 1093 587 1094
rect 615 1098 619 1099
rect 615 1093 619 1094
rect 112 1078 114 1093
rect 144 1088 146 1093
rect 288 1088 290 1093
rect 448 1088 450 1093
rect 616 1088 618 1093
rect 142 1087 148 1088
rect 142 1083 143 1087
rect 147 1083 148 1087
rect 142 1082 148 1083
rect 286 1087 292 1088
rect 286 1083 287 1087
rect 291 1083 292 1087
rect 286 1082 292 1083
rect 446 1087 452 1088
rect 446 1083 447 1087
rect 451 1083 452 1087
rect 446 1082 452 1083
rect 614 1087 620 1088
rect 614 1083 615 1087
rect 619 1083 620 1087
rect 614 1082 620 1083
rect 110 1077 116 1078
rect 110 1073 111 1077
rect 115 1073 116 1077
rect 110 1072 116 1073
rect 514 1063 520 1064
rect 110 1060 116 1061
rect 110 1056 111 1060
rect 115 1056 116 1060
rect 514 1059 515 1063
rect 519 1059 520 1063
rect 514 1058 520 1059
rect 110 1055 116 1056
rect 112 1027 114 1055
rect 150 1047 156 1048
rect 150 1043 151 1047
rect 155 1043 156 1047
rect 294 1047 300 1048
rect 150 1042 156 1043
rect 163 1044 167 1045
rect 152 1027 154 1042
rect 294 1043 295 1047
rect 299 1043 300 1047
rect 294 1042 300 1043
rect 454 1047 460 1048
rect 454 1043 455 1047
rect 459 1043 460 1047
rect 454 1042 460 1043
rect 163 1039 167 1040
rect 164 1036 166 1039
rect 162 1035 168 1036
rect 162 1031 163 1035
rect 167 1031 168 1035
rect 162 1030 168 1031
rect 296 1027 298 1042
rect 456 1027 458 1042
rect 111 1026 115 1027
rect 111 1021 115 1022
rect 143 1026 147 1027
rect 143 1021 147 1022
rect 151 1026 155 1027
rect 151 1021 155 1022
rect 287 1026 291 1027
rect 287 1021 291 1022
rect 295 1026 299 1027
rect 295 1021 299 1022
rect 455 1026 459 1027
rect 455 1021 459 1022
rect 471 1026 475 1027
rect 471 1021 475 1022
rect 112 997 114 1021
rect 144 1010 146 1021
rect 246 1019 252 1020
rect 246 1015 247 1019
rect 251 1015 252 1019
rect 246 1014 252 1015
rect 142 1009 148 1010
rect 142 1005 143 1009
rect 147 1005 148 1009
rect 142 1004 148 1005
rect 248 997 250 1014
rect 288 1010 290 1021
rect 472 1010 474 1021
rect 516 1020 518 1058
rect 622 1047 628 1048
rect 622 1043 623 1047
rect 627 1043 628 1047
rect 622 1042 628 1043
rect 624 1027 626 1042
rect 632 1036 634 1102
rect 704 1099 706 1108
rect 824 1099 826 1108
rect 944 1099 946 1108
rect 1056 1099 1058 1108
rect 1176 1099 1178 1108
rect 1296 1099 1298 1108
rect 703 1098 707 1099
rect 703 1093 707 1094
rect 783 1098 787 1099
rect 783 1093 787 1094
rect 823 1098 827 1099
rect 823 1093 827 1094
rect 943 1098 947 1099
rect 943 1093 947 1094
rect 1055 1098 1059 1099
rect 1055 1093 1059 1094
rect 1103 1098 1107 1099
rect 1103 1093 1107 1094
rect 1175 1098 1179 1099
rect 1175 1093 1179 1094
rect 1255 1098 1259 1099
rect 1255 1093 1259 1094
rect 1295 1098 1299 1099
rect 1295 1093 1299 1094
rect 784 1088 786 1093
rect 944 1088 946 1093
rect 1104 1088 1106 1093
rect 1256 1088 1258 1093
rect 782 1087 788 1088
rect 782 1083 783 1087
rect 787 1083 788 1087
rect 782 1082 788 1083
rect 942 1087 948 1088
rect 942 1083 943 1087
rect 947 1083 948 1087
rect 942 1082 948 1083
rect 1102 1087 1108 1088
rect 1102 1083 1103 1087
rect 1107 1083 1108 1087
rect 1102 1082 1108 1083
rect 1254 1087 1260 1088
rect 1254 1083 1255 1087
rect 1259 1083 1260 1087
rect 1254 1082 1260 1083
rect 1324 1080 1326 1158
rect 1424 1154 1426 1165
rect 1814 1163 1815 1167
rect 1819 1163 1820 1167
rect 1863 1169 1867 1170
rect 1895 1174 1899 1175
rect 1895 1169 1899 1170
rect 2007 1174 2011 1175
rect 2007 1169 2011 1170
rect 2143 1174 2147 1175
rect 2143 1169 2147 1170
rect 2151 1174 2155 1175
rect 2210 1174 2216 1175
rect 2295 1174 2299 1175
rect 2151 1169 2155 1170
rect 2295 1169 2299 1170
rect 2327 1174 2331 1175
rect 2354 1174 2360 1175
rect 2455 1174 2459 1175
rect 2327 1169 2331 1170
rect 1823 1165 1827 1166
rect 1814 1162 1820 1163
rect 1422 1153 1428 1154
rect 1422 1149 1423 1153
rect 1427 1149 1428 1153
rect 1422 1148 1428 1149
rect 1824 1141 1826 1165
rect 1864 1145 1866 1169
rect 1896 1158 1898 1169
rect 2008 1158 2010 1169
rect 2144 1158 2146 1169
rect 2296 1158 2298 1169
rect 2302 1167 2308 1168
rect 2302 1163 2303 1167
rect 2307 1163 2308 1167
rect 2302 1162 2308 1163
rect 1894 1157 1900 1158
rect 1894 1153 1895 1157
rect 1899 1153 1900 1157
rect 1894 1152 1900 1153
rect 2006 1157 2012 1158
rect 2006 1153 2007 1157
rect 2011 1153 2012 1157
rect 2006 1152 2012 1153
rect 2142 1157 2148 1158
rect 2142 1153 2143 1157
rect 2147 1153 2148 1157
rect 2142 1152 2148 1153
rect 2294 1157 2300 1158
rect 2294 1153 2295 1157
rect 2299 1153 2300 1157
rect 2294 1152 2300 1153
rect 1862 1144 1868 1145
rect 1822 1140 1828 1141
rect 1822 1136 1823 1140
rect 1827 1136 1828 1140
rect 1862 1140 1863 1144
rect 1867 1140 1868 1144
rect 1862 1139 1868 1140
rect 1822 1135 1828 1136
rect 1862 1127 1868 1128
rect 1822 1123 1828 1124
rect 1822 1119 1823 1123
rect 1827 1119 1828 1123
rect 1862 1123 1863 1127
rect 1867 1123 1868 1127
rect 1862 1122 1868 1123
rect 2074 1127 2080 1128
rect 2074 1123 2075 1127
rect 2079 1123 2080 1127
rect 2074 1122 2080 1123
rect 1822 1118 1828 1119
rect 1414 1113 1420 1114
rect 1414 1109 1415 1113
rect 1419 1109 1420 1113
rect 1414 1108 1420 1109
rect 1416 1099 1418 1108
rect 1824 1099 1826 1118
rect 1864 1099 1866 1122
rect 1886 1117 1892 1118
rect 1886 1113 1887 1117
rect 1891 1113 1892 1117
rect 1886 1112 1892 1113
rect 1998 1117 2004 1118
rect 1998 1113 1999 1117
rect 2003 1113 2004 1117
rect 1998 1112 2004 1113
rect 1888 1099 1890 1112
rect 2000 1099 2002 1112
rect 1407 1098 1411 1099
rect 1407 1093 1411 1094
rect 1415 1098 1419 1099
rect 1415 1093 1419 1094
rect 1559 1098 1563 1099
rect 1559 1093 1563 1094
rect 1823 1098 1827 1099
rect 1823 1093 1827 1094
rect 1863 1098 1867 1099
rect 1863 1093 1867 1094
rect 1887 1098 1891 1099
rect 1887 1093 1891 1094
rect 1895 1098 1899 1099
rect 1895 1093 1899 1094
rect 1999 1098 2003 1099
rect 1999 1093 2003 1094
rect 2047 1098 2051 1099
rect 2047 1093 2051 1094
rect 1408 1088 1410 1093
rect 1560 1088 1562 1093
rect 1406 1087 1412 1088
rect 1406 1083 1407 1087
rect 1411 1083 1412 1087
rect 1406 1082 1412 1083
rect 1558 1087 1564 1088
rect 1558 1083 1559 1087
rect 1563 1083 1564 1087
rect 1558 1082 1564 1083
rect 682 1079 688 1080
rect 682 1075 683 1079
rect 687 1075 688 1079
rect 682 1074 688 1075
rect 1322 1079 1328 1080
rect 1322 1075 1323 1079
rect 1327 1075 1328 1079
rect 1322 1074 1328 1075
rect 1474 1079 1480 1080
rect 1474 1075 1475 1079
rect 1479 1075 1480 1079
rect 1824 1078 1826 1093
rect 1864 1078 1866 1093
rect 1896 1088 1898 1093
rect 2048 1088 2050 1093
rect 1894 1087 1900 1088
rect 1894 1083 1895 1087
rect 1899 1083 1900 1087
rect 1894 1082 1900 1083
rect 2046 1087 2052 1088
rect 2046 1083 2047 1087
rect 2051 1083 2052 1087
rect 2046 1082 2052 1083
rect 1474 1074 1480 1075
rect 1822 1077 1828 1078
rect 684 1045 686 1074
rect 1242 1063 1248 1064
rect 1242 1059 1243 1063
rect 1247 1059 1248 1063
rect 1242 1058 1248 1059
rect 790 1047 796 1048
rect 683 1044 687 1045
rect 790 1043 791 1047
rect 795 1043 796 1047
rect 790 1042 796 1043
rect 950 1047 956 1048
rect 950 1043 951 1047
rect 955 1043 956 1047
rect 1110 1047 1116 1048
rect 950 1042 956 1043
rect 959 1044 963 1045
rect 683 1039 687 1040
rect 630 1035 636 1036
rect 630 1031 631 1035
rect 635 1031 636 1035
rect 630 1030 636 1031
rect 792 1027 794 1042
rect 952 1027 954 1042
rect 1110 1043 1111 1047
rect 1115 1043 1116 1047
rect 1110 1042 1116 1043
rect 959 1039 963 1040
rect 960 1036 962 1039
rect 958 1035 964 1036
rect 958 1031 959 1035
rect 963 1031 964 1035
rect 958 1030 964 1031
rect 1112 1027 1114 1042
rect 1244 1036 1246 1058
rect 1262 1047 1268 1048
rect 1262 1043 1263 1047
rect 1267 1043 1268 1047
rect 1262 1042 1268 1043
rect 1414 1047 1420 1048
rect 1414 1043 1415 1047
rect 1419 1043 1420 1047
rect 1476 1045 1478 1074
rect 1822 1073 1823 1077
rect 1827 1073 1828 1077
rect 1822 1072 1828 1073
rect 1862 1077 1868 1078
rect 1862 1073 1863 1077
rect 1867 1073 1868 1077
rect 1862 1072 1868 1073
rect 1982 1063 1988 1064
rect 1822 1060 1828 1061
rect 1822 1056 1823 1060
rect 1827 1056 1828 1060
rect 1822 1055 1828 1056
rect 1862 1060 1868 1061
rect 1862 1056 1863 1060
rect 1867 1056 1868 1060
rect 1982 1059 1983 1063
rect 1987 1059 1988 1063
rect 1982 1058 1988 1059
rect 1990 1063 1996 1064
rect 1990 1059 1991 1063
rect 1995 1059 1996 1063
rect 1990 1058 1996 1059
rect 1862 1055 1868 1056
rect 1566 1047 1572 1048
rect 1414 1042 1420 1043
rect 1475 1044 1479 1045
rect 1242 1035 1248 1036
rect 1242 1031 1243 1035
rect 1247 1031 1248 1035
rect 1242 1030 1248 1031
rect 1264 1027 1266 1042
rect 1416 1027 1418 1042
rect 1566 1043 1567 1047
rect 1571 1043 1572 1047
rect 1566 1042 1572 1043
rect 1475 1039 1479 1040
rect 1434 1035 1440 1036
rect 1434 1031 1435 1035
rect 1439 1031 1440 1035
rect 1434 1030 1440 1031
rect 623 1026 627 1027
rect 623 1021 627 1022
rect 663 1026 667 1027
rect 663 1021 667 1022
rect 791 1026 795 1027
rect 791 1021 795 1022
rect 847 1026 851 1027
rect 847 1021 851 1022
rect 951 1026 955 1027
rect 951 1021 955 1022
rect 1031 1026 1035 1027
rect 1031 1021 1035 1022
rect 1111 1026 1115 1027
rect 1111 1021 1115 1022
rect 1207 1026 1211 1027
rect 1207 1021 1211 1022
rect 1263 1026 1267 1027
rect 1263 1021 1267 1022
rect 1375 1026 1379 1027
rect 1375 1021 1379 1022
rect 1415 1026 1419 1027
rect 1415 1021 1419 1022
rect 514 1019 520 1020
rect 514 1015 515 1019
rect 519 1015 520 1019
rect 514 1014 520 1015
rect 664 1010 666 1021
rect 848 1010 850 1021
rect 1032 1010 1034 1021
rect 1118 1019 1124 1020
rect 1118 1015 1119 1019
rect 1123 1015 1124 1019
rect 1118 1014 1124 1015
rect 286 1009 292 1010
rect 286 1005 287 1009
rect 291 1005 292 1009
rect 286 1004 292 1005
rect 470 1009 476 1010
rect 470 1005 471 1009
rect 475 1005 476 1009
rect 470 1004 476 1005
rect 662 1009 668 1010
rect 662 1005 663 1009
rect 667 1005 668 1009
rect 662 1004 668 1005
rect 846 1009 852 1010
rect 846 1005 847 1009
rect 851 1005 852 1009
rect 846 1004 852 1005
rect 1030 1009 1036 1010
rect 1030 1005 1031 1009
rect 1035 1005 1036 1009
rect 1030 1004 1036 1005
rect 1120 997 1122 1014
rect 1208 1010 1210 1021
rect 1376 1010 1378 1021
rect 1206 1009 1212 1010
rect 1206 1005 1207 1009
rect 1211 1005 1212 1009
rect 1206 1004 1212 1005
rect 1374 1009 1380 1010
rect 1374 1005 1375 1009
rect 1379 1005 1380 1009
rect 1374 1004 1380 1005
rect 110 996 116 997
rect 110 992 111 996
rect 115 992 116 996
rect 110 991 116 992
rect 247 996 251 997
rect 771 996 775 997
rect 1119 996 1123 997
rect 1436 996 1438 1030
rect 1568 1027 1570 1042
rect 1824 1027 1826 1055
rect 1864 1027 1866 1055
rect 1902 1047 1908 1048
rect 1902 1043 1903 1047
rect 1907 1043 1908 1047
rect 1902 1042 1908 1043
rect 1904 1027 1906 1042
rect 1543 1026 1547 1027
rect 1543 1021 1547 1022
rect 1567 1026 1571 1027
rect 1567 1021 1571 1022
rect 1711 1026 1715 1027
rect 1711 1021 1715 1022
rect 1823 1026 1827 1027
rect 1823 1021 1827 1022
rect 1863 1026 1867 1027
rect 1863 1021 1867 1022
rect 1903 1026 1907 1027
rect 1903 1021 1907 1022
rect 1975 1026 1979 1027
rect 1975 1021 1979 1022
rect 1544 1010 1546 1021
rect 1610 1019 1616 1020
rect 1610 1015 1611 1019
rect 1615 1015 1616 1019
rect 1610 1014 1616 1015
rect 1542 1009 1548 1010
rect 1542 1005 1543 1009
rect 1547 1005 1548 1009
rect 1542 1004 1548 1005
rect 1459 996 1463 997
rect 247 991 251 992
rect 770 991 776 992
rect 1119 991 1123 992
rect 1434 995 1440 996
rect 1434 991 1435 995
rect 1439 991 1440 995
rect 1612 992 1614 1014
rect 1712 1010 1714 1021
rect 1718 1019 1724 1020
rect 1718 1015 1719 1019
rect 1723 1015 1724 1019
rect 1718 1014 1724 1015
rect 1710 1009 1716 1010
rect 1710 1005 1711 1009
rect 1715 1005 1716 1009
rect 1710 1004 1716 1005
rect 770 987 771 991
rect 775 987 776 991
rect 1434 990 1440 991
rect 1458 991 1464 992
rect 770 986 776 987
rect 1458 987 1459 991
rect 1463 987 1464 991
rect 1458 986 1464 987
rect 1610 991 1616 992
rect 1610 987 1611 991
rect 1615 987 1616 991
rect 1610 986 1616 987
rect 110 979 116 980
rect 110 975 111 979
rect 115 975 116 979
rect 110 974 116 975
rect 112 955 114 974
rect 134 969 140 970
rect 134 965 135 969
rect 139 965 140 969
rect 134 964 140 965
rect 278 969 284 970
rect 278 965 279 969
rect 283 965 284 969
rect 278 964 284 965
rect 462 969 468 970
rect 462 965 463 969
rect 467 965 468 969
rect 462 964 468 965
rect 654 969 660 970
rect 654 965 655 969
rect 659 965 660 969
rect 654 964 660 965
rect 838 969 844 970
rect 838 965 839 969
rect 843 965 844 969
rect 838 964 844 965
rect 1022 969 1028 970
rect 1022 965 1023 969
rect 1027 965 1028 969
rect 1022 964 1028 965
rect 1198 969 1204 970
rect 1198 965 1199 969
rect 1203 965 1204 969
rect 1198 964 1204 965
rect 1366 969 1372 970
rect 1366 965 1367 969
rect 1371 965 1372 969
rect 1366 964 1372 965
rect 1534 969 1540 970
rect 1534 965 1535 969
rect 1539 965 1540 969
rect 1534 964 1540 965
rect 1702 969 1708 970
rect 1702 965 1703 969
rect 1707 965 1708 969
rect 1702 964 1708 965
rect 136 955 138 964
rect 280 955 282 964
rect 464 955 466 964
rect 656 955 658 964
rect 840 955 842 964
rect 1024 955 1026 964
rect 1200 955 1202 964
rect 1368 955 1370 964
rect 1536 955 1538 964
rect 1704 955 1706 964
rect 111 954 115 955
rect 111 949 115 950
rect 135 954 139 955
rect 135 949 139 950
rect 279 954 283 955
rect 279 949 283 950
rect 287 954 291 955
rect 287 949 291 950
rect 463 954 467 955
rect 463 949 467 950
rect 471 954 475 955
rect 471 949 475 950
rect 655 954 659 955
rect 655 949 659 950
rect 663 954 667 955
rect 663 949 667 950
rect 839 954 843 955
rect 839 949 843 950
rect 855 954 859 955
rect 855 949 859 950
rect 1023 954 1027 955
rect 1023 949 1027 950
rect 1047 954 1051 955
rect 1047 949 1051 950
rect 1199 954 1203 955
rect 1199 949 1203 950
rect 1223 954 1227 955
rect 1223 949 1227 950
rect 1367 954 1371 955
rect 1367 949 1371 950
rect 1399 954 1403 955
rect 1399 949 1403 950
rect 1535 954 1539 955
rect 1535 949 1539 950
rect 1575 954 1579 955
rect 1575 949 1579 950
rect 1703 954 1707 955
rect 1703 949 1707 950
rect 112 934 114 949
rect 136 944 138 949
rect 288 944 290 949
rect 472 944 474 949
rect 664 944 666 949
rect 856 944 858 949
rect 1048 944 1050 949
rect 1224 944 1226 949
rect 1400 944 1402 949
rect 1576 944 1578 949
rect 134 943 140 944
rect 134 939 135 943
rect 139 939 140 943
rect 134 938 140 939
rect 286 943 292 944
rect 286 939 287 943
rect 291 939 292 943
rect 286 938 292 939
rect 470 943 476 944
rect 470 939 471 943
rect 475 939 476 943
rect 470 938 476 939
rect 662 943 668 944
rect 662 939 663 943
rect 667 939 668 943
rect 662 938 668 939
rect 854 943 860 944
rect 854 939 855 943
rect 859 939 860 943
rect 854 938 860 939
rect 1046 943 1052 944
rect 1046 939 1047 943
rect 1051 939 1052 943
rect 1046 938 1052 939
rect 1222 943 1228 944
rect 1222 939 1223 943
rect 1227 939 1228 943
rect 1222 938 1228 939
rect 1398 943 1404 944
rect 1398 939 1399 943
rect 1403 939 1404 943
rect 1398 938 1404 939
rect 1574 943 1580 944
rect 1574 939 1575 943
rect 1579 939 1580 943
rect 1574 938 1580 939
rect 1720 936 1722 1014
rect 1824 997 1826 1021
rect 1864 997 1866 1021
rect 1976 1010 1978 1021
rect 1984 1020 1986 1058
rect 1992 1036 1994 1058
rect 2054 1047 2060 1048
rect 2054 1043 2055 1047
rect 2059 1043 2060 1047
rect 2054 1042 2060 1043
rect 1990 1035 1996 1036
rect 1990 1031 1991 1035
rect 1995 1031 1996 1035
rect 1990 1030 1996 1031
rect 2056 1027 2058 1042
rect 2076 1036 2078 1122
rect 2134 1117 2140 1118
rect 2134 1113 2135 1117
rect 2139 1113 2140 1117
rect 2134 1112 2140 1113
rect 2286 1117 2292 1118
rect 2286 1113 2287 1117
rect 2291 1113 2292 1117
rect 2286 1112 2292 1113
rect 2136 1099 2138 1112
rect 2288 1099 2290 1112
rect 2135 1098 2139 1099
rect 2135 1093 2139 1094
rect 2215 1098 2219 1099
rect 2215 1093 2219 1094
rect 2287 1098 2291 1099
rect 2287 1093 2291 1094
rect 2216 1088 2218 1093
rect 2214 1087 2220 1088
rect 2214 1083 2215 1087
rect 2219 1083 2220 1087
rect 2214 1082 2220 1083
rect 2304 1080 2306 1162
rect 2356 1144 2358 1174
rect 2455 1169 2459 1170
rect 2495 1174 2499 1175
rect 2506 1174 2512 1175
rect 2623 1174 2627 1175
rect 2495 1169 2499 1170
rect 2623 1169 2627 1170
rect 2663 1174 2667 1175
rect 2682 1174 2688 1175
rect 2791 1174 2795 1175
rect 2798 1174 2804 1175
rect 2831 1174 2835 1175
rect 2663 1169 2667 1170
rect 2456 1158 2458 1169
rect 2624 1158 2626 1169
rect 2634 1167 2640 1168
rect 2634 1163 2635 1167
rect 2639 1163 2640 1167
rect 2634 1162 2640 1163
rect 2454 1157 2460 1158
rect 2454 1153 2455 1157
rect 2459 1153 2460 1157
rect 2454 1152 2460 1153
rect 2622 1157 2628 1158
rect 2622 1153 2623 1157
rect 2627 1153 2628 1157
rect 2622 1152 2628 1153
rect 2354 1143 2360 1144
rect 2354 1139 2355 1143
rect 2359 1139 2360 1143
rect 2354 1138 2360 1139
rect 2582 1127 2588 1128
rect 2582 1123 2583 1127
rect 2587 1123 2588 1127
rect 2582 1122 2588 1123
rect 2446 1117 2452 1118
rect 2446 1113 2447 1117
rect 2451 1113 2452 1117
rect 2446 1112 2452 1113
rect 2448 1099 2450 1112
rect 2391 1098 2395 1099
rect 2391 1093 2395 1094
rect 2447 1098 2451 1099
rect 2447 1093 2451 1094
rect 2567 1098 2571 1099
rect 2567 1093 2571 1094
rect 2392 1088 2394 1093
rect 2568 1088 2570 1093
rect 2390 1087 2396 1088
rect 2390 1083 2391 1087
rect 2395 1083 2396 1087
rect 2390 1082 2396 1083
rect 2566 1087 2572 1088
rect 2566 1083 2567 1087
rect 2571 1083 2572 1087
rect 2566 1082 2572 1083
rect 2302 1079 2308 1080
rect 2302 1075 2303 1079
rect 2307 1075 2308 1079
rect 2302 1074 2308 1075
rect 2282 1063 2288 1064
rect 2282 1059 2283 1063
rect 2287 1059 2288 1063
rect 2282 1058 2288 1059
rect 2506 1063 2512 1064
rect 2506 1059 2507 1063
rect 2511 1059 2512 1063
rect 2506 1058 2512 1059
rect 2222 1047 2228 1048
rect 2222 1043 2223 1047
rect 2227 1043 2228 1047
rect 2222 1042 2228 1043
rect 2074 1035 2080 1036
rect 2074 1031 2075 1035
rect 2079 1031 2080 1035
rect 2074 1030 2080 1031
rect 2224 1027 2226 1042
rect 2284 1036 2286 1058
rect 2398 1047 2404 1048
rect 2398 1043 2399 1047
rect 2403 1043 2404 1047
rect 2398 1042 2404 1043
rect 2282 1035 2288 1036
rect 2282 1031 2283 1035
rect 2287 1031 2288 1035
rect 2282 1030 2288 1031
rect 2400 1027 2402 1042
rect 2418 1035 2424 1036
rect 2418 1031 2419 1035
rect 2423 1031 2424 1035
rect 2418 1030 2424 1031
rect 2055 1026 2059 1027
rect 2055 1021 2059 1022
rect 2095 1026 2099 1027
rect 2095 1021 2099 1022
rect 2223 1026 2227 1027
rect 2223 1021 2227 1022
rect 2359 1026 2363 1027
rect 2359 1021 2363 1022
rect 2399 1026 2403 1027
rect 2399 1021 2403 1022
rect 1982 1019 1988 1020
rect 1982 1015 1983 1019
rect 1987 1015 1988 1019
rect 1982 1014 1988 1015
rect 2066 1019 2072 1020
rect 2066 1015 2067 1019
rect 2071 1015 2072 1019
rect 2066 1014 2072 1015
rect 1974 1009 1980 1010
rect 1974 1005 1975 1009
rect 1979 1005 1980 1009
rect 1974 1004 1980 1005
rect 1822 996 1828 997
rect 1822 992 1823 996
rect 1827 992 1828 996
rect 1822 991 1828 992
rect 1862 996 1868 997
rect 2068 996 2070 1014
rect 2096 1010 2098 1021
rect 2224 1010 2226 1021
rect 2360 1010 2362 1021
rect 2094 1009 2100 1010
rect 2094 1005 2095 1009
rect 2099 1005 2100 1009
rect 2094 1004 2100 1005
rect 2222 1009 2228 1010
rect 2222 1005 2223 1009
rect 2227 1005 2228 1009
rect 2222 1004 2228 1005
rect 2358 1009 2364 1010
rect 2358 1005 2359 1009
rect 2363 1005 2364 1009
rect 2358 1004 2364 1005
rect 2420 996 2422 1030
rect 2495 1026 2499 1027
rect 2495 1021 2499 1022
rect 2496 1010 2498 1021
rect 2508 1020 2510 1058
rect 2574 1047 2580 1048
rect 2574 1043 2575 1047
rect 2579 1043 2580 1047
rect 2574 1042 2580 1043
rect 2576 1027 2578 1042
rect 2584 1036 2586 1122
rect 2614 1117 2620 1118
rect 2614 1113 2615 1117
rect 2619 1113 2620 1117
rect 2614 1112 2620 1113
rect 2636 1112 2638 1162
rect 2684 1144 2686 1174
rect 2791 1169 2795 1170
rect 2831 1169 2835 1170
rect 2967 1174 2971 1175
rect 2967 1169 2971 1170
rect 2999 1174 3003 1175
rect 3058 1174 3064 1175
rect 3143 1174 3147 1175
rect 2999 1169 3003 1170
rect 3143 1169 3147 1170
rect 2792 1158 2794 1169
rect 2802 1167 2808 1168
rect 2802 1163 2803 1167
rect 2807 1163 2808 1167
rect 2802 1162 2808 1163
rect 2790 1157 2796 1158
rect 2790 1153 2791 1157
rect 2795 1153 2796 1157
rect 2790 1152 2796 1153
rect 2682 1143 2688 1144
rect 2682 1139 2683 1143
rect 2687 1139 2688 1143
rect 2682 1138 2688 1139
rect 2782 1117 2788 1118
rect 2782 1113 2783 1117
rect 2787 1113 2788 1117
rect 2782 1112 2788 1113
rect 2616 1099 2618 1112
rect 2634 1111 2640 1112
rect 2634 1107 2635 1111
rect 2639 1107 2640 1111
rect 2634 1106 2640 1107
rect 2784 1099 2786 1112
rect 2615 1098 2619 1099
rect 2615 1093 2619 1094
rect 2735 1098 2739 1099
rect 2735 1093 2739 1094
rect 2783 1098 2787 1099
rect 2783 1093 2787 1094
rect 2736 1088 2738 1093
rect 2734 1087 2740 1088
rect 2734 1083 2735 1087
rect 2739 1083 2740 1087
rect 2734 1082 2740 1083
rect 2804 1080 2806 1162
rect 2968 1158 2970 1169
rect 3144 1158 3146 1169
rect 3152 1168 3154 1202
rect 3166 1191 3172 1192
rect 3166 1187 3167 1191
rect 3171 1187 3172 1191
rect 3166 1186 3172 1187
rect 3168 1175 3170 1186
rect 3228 1180 3230 1202
rect 3334 1191 3340 1192
rect 3334 1187 3335 1191
rect 3339 1187 3340 1191
rect 3334 1186 3340 1187
rect 3226 1179 3232 1180
rect 3226 1175 3227 1179
rect 3231 1175 3232 1179
rect 3336 1175 3338 1186
rect 3348 1180 3350 1250
rect 3346 1179 3352 1180
rect 3346 1175 3347 1179
rect 3351 1175 3352 1179
rect 3167 1174 3171 1175
rect 3226 1174 3232 1175
rect 3327 1174 3331 1175
rect 3167 1169 3171 1170
rect 3327 1169 3331 1170
rect 3335 1174 3339 1175
rect 3346 1174 3352 1175
rect 3335 1169 3339 1170
rect 3150 1167 3156 1168
rect 3150 1163 3151 1167
rect 3155 1163 3156 1167
rect 3150 1162 3156 1163
rect 3328 1158 3330 1169
rect 2966 1157 2972 1158
rect 2966 1153 2967 1157
rect 2971 1153 2972 1157
rect 2966 1152 2972 1153
rect 3142 1157 3148 1158
rect 3142 1153 3143 1157
rect 3147 1153 3148 1157
rect 3142 1152 3148 1153
rect 3326 1157 3332 1158
rect 3326 1153 3327 1157
rect 3331 1153 3332 1157
rect 3326 1152 3332 1153
rect 2958 1117 2964 1118
rect 2958 1113 2959 1117
rect 2963 1113 2964 1117
rect 2958 1112 2964 1113
rect 3134 1117 3140 1118
rect 3134 1113 3135 1117
rect 3139 1113 3140 1117
rect 3134 1112 3140 1113
rect 3318 1117 3324 1118
rect 3318 1113 3319 1117
rect 3323 1113 3324 1117
rect 3318 1112 3324 1113
rect 2960 1099 2962 1112
rect 3136 1099 3138 1112
rect 3320 1099 3322 1112
rect 3366 1111 3372 1112
rect 3366 1107 3367 1111
rect 3371 1107 3372 1111
rect 3366 1106 3372 1107
rect 2895 1098 2899 1099
rect 2895 1093 2899 1094
rect 2959 1098 2963 1099
rect 2959 1093 2963 1094
rect 3047 1098 3051 1099
rect 3047 1093 3051 1094
rect 3135 1098 3139 1099
rect 3135 1093 3139 1094
rect 3199 1098 3203 1099
rect 3199 1093 3203 1094
rect 3319 1098 3323 1099
rect 3319 1093 3323 1094
rect 3351 1098 3355 1099
rect 3351 1093 3355 1094
rect 2896 1088 2898 1093
rect 3048 1088 3050 1093
rect 3200 1088 3202 1093
rect 3352 1088 3354 1093
rect 2894 1087 2900 1088
rect 2894 1083 2895 1087
rect 2899 1083 2900 1087
rect 2894 1082 2900 1083
rect 3046 1087 3052 1088
rect 3046 1083 3047 1087
rect 3051 1083 3052 1087
rect 3046 1082 3052 1083
rect 3198 1087 3204 1088
rect 3198 1083 3199 1087
rect 3203 1083 3204 1087
rect 3198 1082 3204 1083
rect 3350 1087 3356 1088
rect 3350 1083 3351 1087
rect 3355 1083 3356 1087
rect 3350 1082 3356 1083
rect 2802 1079 2808 1080
rect 2802 1075 2803 1079
rect 2807 1075 2808 1079
rect 2802 1074 2808 1075
rect 2802 1063 2808 1064
rect 2802 1059 2803 1063
rect 2807 1059 2808 1063
rect 2802 1058 2808 1059
rect 2962 1063 2968 1064
rect 2962 1059 2963 1063
rect 2967 1059 2968 1063
rect 2962 1058 2968 1059
rect 3114 1063 3120 1064
rect 3114 1059 3115 1063
rect 3119 1059 3120 1063
rect 3114 1058 3120 1059
rect 3266 1063 3272 1064
rect 3266 1059 3267 1063
rect 3271 1059 3272 1063
rect 3266 1058 3272 1059
rect 2742 1047 2748 1048
rect 2742 1043 2743 1047
rect 2747 1043 2748 1047
rect 2742 1042 2748 1043
rect 2582 1035 2588 1036
rect 2582 1031 2583 1035
rect 2587 1031 2588 1035
rect 2582 1030 2588 1031
rect 2744 1027 2746 1042
rect 2575 1026 2579 1027
rect 2575 1021 2579 1022
rect 2639 1026 2643 1027
rect 2639 1021 2643 1022
rect 2743 1026 2747 1027
rect 2743 1021 2747 1022
rect 2791 1026 2795 1027
rect 2791 1021 2795 1022
rect 2506 1019 2512 1020
rect 2506 1015 2507 1019
rect 2511 1015 2512 1019
rect 2506 1014 2512 1015
rect 2640 1010 2642 1021
rect 2682 1019 2688 1020
rect 2682 1015 2683 1019
rect 2687 1015 2688 1019
rect 2682 1014 2688 1015
rect 2494 1009 2500 1010
rect 2494 1005 2495 1009
rect 2499 1005 2500 1009
rect 2494 1004 2500 1005
rect 2638 1009 2644 1010
rect 2638 1005 2639 1009
rect 2643 1005 2644 1009
rect 2638 1004 2644 1005
rect 1862 992 1863 996
rect 1867 992 1868 996
rect 1862 991 1868 992
rect 2066 995 2072 996
rect 2066 991 2067 995
rect 2071 991 2072 995
rect 2066 990 2072 991
rect 2418 995 2424 996
rect 2418 991 2419 995
rect 2423 991 2424 995
rect 2418 990 2424 991
rect 1822 979 1828 980
rect 1822 975 1823 979
rect 1827 975 1828 979
rect 1822 974 1828 975
rect 1862 979 1868 980
rect 1862 975 1863 979
rect 1867 975 1868 979
rect 1862 974 1868 975
rect 1824 955 1826 974
rect 1864 955 1866 974
rect 1966 969 1972 970
rect 1966 965 1967 969
rect 1971 965 1972 969
rect 1966 964 1972 965
rect 2086 969 2092 970
rect 2086 965 2087 969
rect 2091 965 2092 969
rect 2086 964 2092 965
rect 2214 969 2220 970
rect 2214 965 2215 969
rect 2219 965 2220 969
rect 2214 964 2220 965
rect 2350 969 2356 970
rect 2350 965 2351 969
rect 2355 965 2356 969
rect 2350 964 2356 965
rect 2486 969 2492 970
rect 2486 965 2487 969
rect 2491 965 2492 969
rect 2486 964 2492 965
rect 2630 969 2636 970
rect 2630 965 2631 969
rect 2635 965 2636 969
rect 2630 964 2636 965
rect 1968 955 1970 964
rect 2088 955 2090 964
rect 2216 955 2218 964
rect 2352 955 2354 964
rect 2488 955 2490 964
rect 2522 963 2528 964
rect 2522 959 2523 963
rect 2527 959 2528 963
rect 2522 958 2528 959
rect 1727 954 1731 955
rect 1727 949 1731 950
rect 1823 954 1827 955
rect 1823 949 1827 950
rect 1863 954 1867 955
rect 1863 949 1867 950
rect 1967 954 1971 955
rect 1967 949 1971 950
rect 2087 954 2091 955
rect 2087 949 2091 950
rect 2143 954 2147 955
rect 2143 949 2147 950
rect 2215 954 2219 955
rect 2215 949 2219 950
rect 2231 954 2235 955
rect 2231 949 2235 950
rect 2319 954 2323 955
rect 2319 949 2323 950
rect 2351 954 2355 955
rect 2351 949 2355 950
rect 2407 954 2411 955
rect 2407 949 2411 950
rect 2487 954 2491 955
rect 2487 949 2491 950
rect 2503 954 2507 955
rect 2503 949 2507 950
rect 1728 944 1730 949
rect 1726 943 1732 944
rect 1726 939 1727 943
rect 1731 939 1732 943
rect 1726 938 1732 939
rect 798 935 804 936
rect 110 933 116 934
rect 110 929 111 933
rect 115 929 116 933
rect 798 931 799 935
rect 803 931 804 935
rect 798 930 804 931
rect 1718 935 1724 936
rect 1718 931 1719 935
rect 1723 931 1724 935
rect 1824 934 1826 949
rect 1864 934 1866 949
rect 2144 944 2146 949
rect 2232 944 2234 949
rect 2320 944 2322 949
rect 2408 944 2410 949
rect 2504 944 2506 949
rect 2142 943 2148 944
rect 2142 939 2143 943
rect 2147 939 2148 943
rect 2142 938 2148 939
rect 2230 943 2236 944
rect 2230 939 2231 943
rect 2235 939 2236 943
rect 2230 938 2236 939
rect 2318 943 2324 944
rect 2318 939 2319 943
rect 2323 939 2324 943
rect 2318 938 2324 939
rect 2406 943 2412 944
rect 2406 939 2407 943
rect 2411 939 2412 943
rect 2406 938 2412 939
rect 2502 943 2508 944
rect 2502 939 2503 943
rect 2507 939 2508 943
rect 2502 938 2508 939
rect 1718 930 1724 931
rect 1822 933 1828 934
rect 110 928 116 929
rect 202 919 208 920
rect 110 916 116 917
rect 110 912 111 916
rect 115 912 116 916
rect 202 915 203 919
rect 207 915 208 919
rect 202 914 208 915
rect 110 911 116 912
rect 112 883 114 911
rect 142 903 148 904
rect 142 899 143 903
rect 147 899 148 903
rect 142 898 148 899
rect 144 883 146 898
rect 204 892 206 914
rect 294 903 300 904
rect 294 899 295 903
rect 299 899 300 903
rect 478 903 484 904
rect 294 898 300 899
rect 303 900 307 901
rect 202 891 208 892
rect 202 887 203 891
rect 207 887 208 891
rect 202 886 208 887
rect 296 883 298 898
rect 478 899 479 903
rect 483 899 484 903
rect 478 898 484 899
rect 670 903 676 904
rect 670 899 671 903
rect 675 899 676 903
rect 800 901 802 930
rect 1822 929 1823 933
rect 1827 929 1828 933
rect 1822 928 1828 929
rect 1862 933 1868 934
rect 1862 929 1863 933
rect 1867 929 1868 933
rect 1862 928 1868 929
rect 2210 919 2216 920
rect 1822 916 1828 917
rect 1822 912 1823 916
rect 1827 912 1828 916
rect 1822 911 1828 912
rect 1862 916 1868 917
rect 1862 912 1863 916
rect 1867 912 1868 916
rect 2210 915 2211 919
rect 2215 915 2216 919
rect 2210 914 2216 915
rect 2298 919 2304 920
rect 2298 915 2299 919
rect 2303 915 2304 919
rect 2298 914 2304 915
rect 2386 919 2392 920
rect 2386 915 2387 919
rect 2391 915 2392 919
rect 2386 914 2392 915
rect 2474 919 2480 920
rect 2474 915 2475 919
rect 2479 915 2480 919
rect 2474 914 2480 915
rect 1862 911 1868 912
rect 862 903 868 904
rect 670 898 676 899
rect 799 900 803 901
rect 303 895 307 896
rect 304 892 306 895
rect 302 891 308 892
rect 302 887 303 891
rect 307 887 308 891
rect 302 886 308 887
rect 480 883 482 898
rect 672 883 674 898
rect 862 899 863 903
rect 867 899 868 903
rect 862 898 868 899
rect 1054 903 1060 904
rect 1054 899 1055 903
rect 1059 899 1060 903
rect 1054 898 1060 899
rect 1230 903 1236 904
rect 1230 899 1231 903
rect 1235 899 1236 903
rect 1230 898 1236 899
rect 1406 903 1412 904
rect 1406 899 1407 903
rect 1411 899 1412 903
rect 1406 898 1412 899
rect 1582 903 1588 904
rect 1582 899 1583 903
rect 1587 899 1588 903
rect 1582 898 1588 899
rect 1734 903 1740 904
rect 1734 899 1735 903
rect 1739 899 1740 903
rect 1734 898 1740 899
rect 799 895 803 896
rect 864 883 866 898
rect 1056 883 1058 898
rect 1206 891 1212 892
rect 1206 887 1207 891
rect 1211 887 1212 891
rect 1206 886 1212 887
rect 111 882 115 883
rect 111 877 115 878
rect 143 882 147 883
rect 143 877 147 878
rect 287 882 291 883
rect 287 877 291 878
rect 295 882 299 883
rect 295 877 299 878
rect 471 882 475 883
rect 471 877 475 878
rect 479 882 483 883
rect 479 877 483 878
rect 655 882 659 883
rect 655 877 659 878
rect 671 882 675 883
rect 671 877 675 878
rect 839 882 843 883
rect 839 877 843 878
rect 863 882 867 883
rect 863 877 867 878
rect 1023 882 1027 883
rect 1023 877 1027 878
rect 1055 882 1059 883
rect 1055 877 1059 878
rect 1191 882 1195 883
rect 1191 877 1195 878
rect 112 853 114 877
rect 144 866 146 877
rect 288 866 290 877
rect 472 866 474 877
rect 656 866 658 877
rect 840 866 842 877
rect 1024 866 1026 877
rect 1086 875 1092 876
rect 1086 871 1087 875
rect 1091 871 1092 875
rect 1086 870 1092 871
rect 142 865 148 866
rect 142 861 143 865
rect 147 861 148 865
rect 142 860 148 861
rect 286 865 292 866
rect 286 861 287 865
rect 291 861 292 865
rect 286 860 292 861
rect 470 865 476 866
rect 470 861 471 865
rect 475 861 476 865
rect 470 860 476 861
rect 654 865 660 866
rect 654 861 655 865
rect 659 861 660 865
rect 654 860 660 861
rect 838 865 844 866
rect 838 861 839 865
rect 843 861 844 865
rect 838 860 844 861
rect 1022 865 1028 866
rect 1022 861 1023 865
rect 1027 861 1028 865
rect 1022 860 1028 861
rect 110 852 116 853
rect 110 848 111 852
rect 115 848 116 852
rect 110 847 116 848
rect 110 835 116 836
rect 110 831 111 835
rect 115 831 116 835
rect 110 830 116 831
rect 750 835 756 836
rect 750 831 751 835
rect 755 831 756 835
rect 750 830 756 831
rect 112 815 114 830
rect 134 825 140 826
rect 134 821 135 825
rect 139 821 140 825
rect 134 820 140 821
rect 278 825 284 826
rect 278 821 279 825
rect 283 821 284 825
rect 278 820 284 821
rect 462 825 468 826
rect 462 821 463 825
rect 467 821 468 825
rect 462 820 468 821
rect 646 825 652 826
rect 646 821 647 825
rect 651 821 652 825
rect 646 820 652 821
rect 136 815 138 820
rect 280 815 282 820
rect 464 815 466 820
rect 648 815 650 820
rect 111 814 115 815
rect 111 809 115 810
rect 135 814 139 815
rect 135 809 139 810
rect 271 814 275 815
rect 271 809 275 810
rect 279 814 283 815
rect 279 809 283 810
rect 423 814 427 815
rect 423 809 427 810
rect 463 814 467 815
rect 463 809 467 810
rect 583 814 587 815
rect 583 809 587 810
rect 647 814 651 815
rect 647 809 651 810
rect 743 814 747 815
rect 743 809 747 810
rect 112 794 114 809
rect 136 804 138 809
rect 272 804 274 809
rect 424 804 426 809
rect 584 804 586 809
rect 744 804 746 809
rect 134 803 140 804
rect 134 799 135 803
rect 139 799 140 803
rect 134 798 140 799
rect 270 803 276 804
rect 270 799 271 803
rect 275 799 276 803
rect 270 798 276 799
rect 422 803 428 804
rect 422 799 423 803
rect 427 799 428 803
rect 422 798 428 799
rect 582 803 588 804
rect 582 799 583 803
rect 587 799 588 803
rect 582 798 588 799
rect 742 803 748 804
rect 742 799 743 803
rect 747 799 748 803
rect 742 798 748 799
rect 752 797 754 830
rect 1088 829 1090 870
rect 1192 866 1194 877
rect 1190 865 1196 866
rect 1190 861 1191 865
rect 1195 861 1196 865
rect 1208 861 1210 886
rect 1232 883 1234 898
rect 1408 883 1410 898
rect 1584 883 1586 898
rect 1736 883 1738 898
rect 1824 883 1826 911
rect 1864 883 1866 911
rect 2150 903 2156 904
rect 2150 899 2151 903
rect 2155 899 2156 903
rect 2150 898 2156 899
rect 2152 883 2154 898
rect 2212 892 2214 914
rect 2238 903 2244 904
rect 2238 899 2239 903
rect 2243 899 2244 903
rect 2238 898 2244 899
rect 2210 891 2216 892
rect 2210 887 2211 891
rect 2215 887 2216 891
rect 2210 886 2216 887
rect 2240 883 2242 898
rect 2300 892 2302 914
rect 2326 903 2332 904
rect 2326 899 2327 903
rect 2331 899 2332 903
rect 2326 898 2332 899
rect 2298 891 2304 892
rect 2298 887 2299 891
rect 2303 887 2304 891
rect 2298 886 2304 887
rect 2328 883 2330 898
rect 2388 892 2390 914
rect 2414 903 2420 904
rect 2414 899 2415 903
rect 2419 899 2420 903
rect 2414 898 2420 899
rect 2386 891 2392 892
rect 2386 887 2387 891
rect 2391 887 2392 891
rect 2386 886 2392 887
rect 2416 883 2418 898
rect 2476 892 2478 914
rect 2510 903 2516 904
rect 2510 899 2511 903
rect 2515 899 2516 903
rect 2510 898 2516 899
rect 2474 891 2480 892
rect 2474 887 2475 891
rect 2479 887 2480 891
rect 2474 886 2480 887
rect 2512 883 2514 898
rect 2524 892 2526 958
rect 2632 955 2634 964
rect 2615 954 2619 955
rect 2615 949 2619 950
rect 2631 954 2635 955
rect 2631 949 2635 950
rect 2616 944 2618 949
rect 2614 943 2620 944
rect 2614 939 2615 943
rect 2619 939 2620 943
rect 2614 938 2620 939
rect 2684 936 2686 1014
rect 2792 1010 2794 1021
rect 2804 1020 2806 1058
rect 2902 1047 2908 1048
rect 2902 1043 2903 1047
rect 2907 1043 2908 1047
rect 2902 1042 2908 1043
rect 2904 1027 2906 1042
rect 2964 1036 2966 1058
rect 3054 1047 3060 1048
rect 3054 1043 3055 1047
rect 3059 1043 3060 1047
rect 3054 1042 3060 1043
rect 2962 1035 2968 1036
rect 2962 1031 2963 1035
rect 2967 1031 2968 1035
rect 2962 1030 2968 1031
rect 3056 1027 3058 1042
rect 3116 1036 3118 1058
rect 3206 1047 3212 1048
rect 3206 1043 3207 1047
rect 3211 1043 3212 1047
rect 3206 1042 3212 1043
rect 3114 1035 3120 1036
rect 3114 1031 3115 1035
rect 3119 1031 3120 1035
rect 3114 1030 3120 1031
rect 3208 1027 3210 1042
rect 3268 1036 3270 1058
rect 3358 1047 3364 1048
rect 3358 1043 3359 1047
rect 3363 1043 3364 1047
rect 3358 1042 3364 1043
rect 3266 1035 3272 1036
rect 3266 1031 3267 1035
rect 3271 1031 3272 1035
rect 3266 1030 3272 1031
rect 3360 1027 3362 1042
rect 3368 1036 3370 1106
rect 3420 1080 3422 1318
rect 3487 1313 3491 1314
rect 3575 1313 3579 1314
rect 3488 1302 3490 1313
rect 3486 1301 3492 1302
rect 3486 1297 3487 1301
rect 3491 1297 3492 1301
rect 3486 1296 3492 1297
rect 3576 1289 3578 1313
rect 3574 1288 3580 1289
rect 3574 1284 3575 1288
rect 3579 1284 3580 1288
rect 3574 1283 3580 1284
rect 3574 1271 3580 1272
rect 3574 1267 3575 1271
rect 3579 1267 3580 1271
rect 3574 1266 3580 1267
rect 3478 1261 3484 1262
rect 3478 1257 3479 1261
rect 3483 1257 3484 1261
rect 3478 1256 3484 1257
rect 3480 1243 3482 1256
rect 3498 1255 3504 1256
rect 3498 1251 3499 1255
rect 3503 1251 3504 1255
rect 3498 1250 3504 1251
rect 3479 1242 3483 1243
rect 3479 1237 3483 1238
rect 3480 1232 3482 1237
rect 3478 1231 3484 1232
rect 3478 1227 3479 1231
rect 3483 1227 3484 1231
rect 3478 1226 3484 1227
rect 3486 1191 3492 1192
rect 3486 1187 3487 1191
rect 3491 1187 3492 1191
rect 3486 1186 3492 1187
rect 3488 1175 3490 1186
rect 3500 1180 3502 1250
rect 3576 1243 3578 1266
rect 3575 1242 3579 1243
rect 3575 1237 3579 1238
rect 3576 1222 3578 1237
rect 3574 1221 3580 1222
rect 3574 1217 3575 1221
rect 3579 1217 3580 1221
rect 3574 1216 3580 1217
rect 3574 1204 3580 1205
rect 3574 1200 3575 1204
rect 3579 1200 3580 1204
rect 3574 1199 3580 1200
rect 3498 1179 3504 1180
rect 3498 1175 3499 1179
rect 3503 1175 3504 1179
rect 3576 1175 3578 1199
rect 3487 1174 3491 1175
rect 3498 1174 3504 1175
rect 3575 1174 3579 1175
rect 3487 1169 3491 1170
rect 3575 1169 3579 1170
rect 3488 1158 3490 1169
rect 3486 1157 3492 1158
rect 3486 1153 3487 1157
rect 3491 1153 3492 1157
rect 3486 1152 3492 1153
rect 3576 1145 3578 1169
rect 3574 1144 3580 1145
rect 3574 1140 3575 1144
rect 3579 1140 3580 1144
rect 3574 1139 3580 1140
rect 3574 1127 3580 1128
rect 3574 1123 3575 1127
rect 3579 1123 3580 1127
rect 3574 1122 3580 1123
rect 3478 1117 3484 1118
rect 3478 1113 3479 1117
rect 3483 1113 3484 1117
rect 3478 1112 3484 1113
rect 3480 1099 3482 1112
rect 3498 1111 3504 1112
rect 3498 1107 3499 1111
rect 3503 1107 3504 1111
rect 3498 1106 3504 1107
rect 3479 1098 3483 1099
rect 3479 1093 3483 1094
rect 3480 1088 3482 1093
rect 3478 1087 3484 1088
rect 3478 1083 3479 1087
rect 3483 1083 3484 1087
rect 3478 1082 3484 1083
rect 3418 1079 3424 1080
rect 3418 1075 3419 1079
rect 3423 1075 3424 1079
rect 3418 1074 3424 1075
rect 3486 1047 3492 1048
rect 3486 1043 3487 1047
rect 3491 1043 3492 1047
rect 3486 1042 3492 1043
rect 3366 1035 3372 1036
rect 3366 1031 3367 1035
rect 3371 1031 3372 1035
rect 3366 1030 3372 1031
rect 3488 1027 3490 1042
rect 2903 1026 2907 1027
rect 2903 1021 2907 1022
rect 2959 1026 2963 1027
rect 2959 1021 2963 1022
rect 3055 1026 3059 1027
rect 3055 1021 3059 1022
rect 3135 1026 3139 1027
rect 3135 1021 3139 1022
rect 3207 1026 3211 1027
rect 3207 1021 3211 1022
rect 3311 1026 3315 1027
rect 3311 1021 3315 1022
rect 3359 1026 3363 1027
rect 3359 1021 3363 1022
rect 3487 1026 3491 1027
rect 3487 1021 3491 1022
rect 2802 1019 2808 1020
rect 2802 1015 2803 1019
rect 2807 1015 2808 1019
rect 2802 1014 2808 1015
rect 2960 1010 2962 1021
rect 3136 1010 3138 1021
rect 3312 1010 3314 1021
rect 3488 1010 3490 1021
rect 3500 1020 3502 1106
rect 3576 1099 3578 1122
rect 3575 1098 3579 1099
rect 3575 1093 3579 1094
rect 3576 1078 3578 1093
rect 3574 1077 3580 1078
rect 3574 1073 3575 1077
rect 3579 1073 3580 1077
rect 3574 1072 3580 1073
rect 3574 1060 3580 1061
rect 3574 1056 3575 1060
rect 3579 1056 3580 1060
rect 3574 1055 3580 1056
rect 3522 1035 3528 1036
rect 3522 1031 3523 1035
rect 3527 1031 3528 1035
rect 3522 1030 3528 1031
rect 3498 1019 3504 1020
rect 3498 1015 3499 1019
rect 3503 1015 3504 1019
rect 3498 1014 3504 1015
rect 2790 1009 2796 1010
rect 2790 1005 2791 1009
rect 2795 1005 2796 1009
rect 2790 1004 2796 1005
rect 2958 1009 2964 1010
rect 2958 1005 2959 1009
rect 2963 1005 2964 1009
rect 2958 1004 2964 1005
rect 3134 1009 3140 1010
rect 3134 1005 3135 1009
rect 3139 1005 3140 1009
rect 3134 1004 3140 1005
rect 3310 1009 3316 1010
rect 3310 1005 3311 1009
rect 3315 1005 3316 1009
rect 3310 1004 3316 1005
rect 3486 1009 3492 1010
rect 3486 1005 3487 1009
rect 3491 1005 3492 1009
rect 3486 1004 3492 1005
rect 3282 979 3288 980
rect 3282 975 3283 979
rect 3287 975 3288 979
rect 3282 974 3288 975
rect 3486 979 3492 980
rect 3486 975 3487 979
rect 3491 975 3492 979
rect 3486 974 3492 975
rect 2782 969 2788 970
rect 2782 965 2783 969
rect 2787 965 2788 969
rect 2782 964 2788 965
rect 2950 969 2956 970
rect 2950 965 2951 969
rect 2955 965 2956 969
rect 2950 964 2956 965
rect 3126 969 3132 970
rect 3126 965 3127 969
rect 3131 965 3132 969
rect 3126 964 3132 965
rect 2784 955 2786 964
rect 2952 955 2954 964
rect 3128 955 3130 964
rect 2751 954 2755 955
rect 2751 949 2755 950
rect 2783 954 2787 955
rect 2783 949 2787 950
rect 2903 954 2907 955
rect 2903 949 2907 950
rect 2951 954 2955 955
rect 2951 949 2955 950
rect 3079 954 3083 955
rect 3079 949 3083 950
rect 3127 954 3131 955
rect 3127 949 3131 950
rect 3263 954 3267 955
rect 3263 949 3267 950
rect 2752 944 2754 949
rect 2904 944 2906 949
rect 3080 944 3082 949
rect 3264 944 3266 949
rect 2750 943 2756 944
rect 2750 939 2751 943
rect 2755 939 2756 943
rect 2750 938 2756 939
rect 2902 943 2908 944
rect 2902 939 2903 943
rect 2907 939 2908 943
rect 2902 938 2908 939
rect 3078 943 3084 944
rect 3078 939 3079 943
rect 3083 939 3084 943
rect 3078 938 3084 939
rect 3262 943 3268 944
rect 3262 939 3263 943
rect 3267 939 3268 943
rect 3262 938 3268 939
rect 2682 935 2688 936
rect 2682 931 2683 935
rect 2687 931 2688 935
rect 2682 930 2688 931
rect 2682 919 2688 920
rect 2682 915 2683 919
rect 2687 915 2688 919
rect 2682 914 2688 915
rect 2818 919 2824 920
rect 2818 915 2819 919
rect 2823 915 2824 919
rect 2818 914 2824 915
rect 2970 919 2976 920
rect 2970 915 2971 919
rect 2975 915 2976 919
rect 2970 914 2976 915
rect 3146 919 3152 920
rect 3146 915 3147 919
rect 3151 915 3152 919
rect 3146 914 3152 915
rect 2622 903 2628 904
rect 2622 899 2623 903
rect 2627 899 2628 903
rect 2622 898 2628 899
rect 2522 891 2528 892
rect 2522 887 2523 891
rect 2527 887 2528 891
rect 2522 886 2528 887
rect 2624 883 2626 898
rect 2684 884 2686 914
rect 2758 903 2764 904
rect 2758 899 2759 903
rect 2763 899 2764 903
rect 2758 898 2764 899
rect 2682 883 2688 884
rect 2760 883 2762 898
rect 2820 892 2822 914
rect 2910 903 2916 904
rect 2910 899 2911 903
rect 2915 899 2916 903
rect 2910 898 2916 899
rect 2818 891 2824 892
rect 2818 887 2819 891
rect 2823 887 2824 891
rect 2818 886 2824 887
rect 2912 883 2914 898
rect 2972 892 2974 914
rect 3086 903 3092 904
rect 3086 899 3087 903
rect 3091 899 3092 903
rect 3086 898 3092 899
rect 2970 891 2976 892
rect 2970 887 2971 891
rect 2975 887 2976 891
rect 2970 886 2976 887
rect 3088 883 3090 898
rect 3148 892 3150 914
rect 3270 903 3276 904
rect 3270 899 3271 903
rect 3275 899 3276 903
rect 3270 898 3276 899
rect 3146 891 3152 892
rect 3146 887 3147 891
rect 3151 887 3152 891
rect 3146 886 3152 887
rect 3272 883 3274 898
rect 3284 892 3286 974
rect 3302 969 3308 970
rect 3302 965 3303 969
rect 3307 965 3308 969
rect 3302 964 3308 965
rect 3478 969 3484 970
rect 3478 965 3479 969
rect 3483 965 3484 969
rect 3478 964 3484 965
rect 3304 955 3306 964
rect 3480 955 3482 964
rect 3303 954 3307 955
rect 3303 949 3307 950
rect 3455 954 3459 955
rect 3455 949 3459 950
rect 3479 954 3483 955
rect 3479 949 3483 950
rect 3456 944 3458 949
rect 3454 943 3460 944
rect 3454 939 3455 943
rect 3459 939 3460 943
rect 3454 938 3460 939
rect 3462 903 3468 904
rect 3462 899 3463 903
rect 3467 899 3468 903
rect 3462 898 3468 899
rect 3282 891 3288 892
rect 3282 887 3283 891
rect 3287 887 3288 891
rect 3282 886 3288 887
rect 3464 883 3466 898
rect 3488 892 3490 974
rect 3524 936 3526 1030
rect 3576 1027 3578 1055
rect 3575 1026 3579 1027
rect 3575 1021 3579 1022
rect 3576 997 3578 1021
rect 3574 996 3580 997
rect 3574 992 3575 996
rect 3579 992 3580 996
rect 3574 991 3580 992
rect 3574 979 3580 980
rect 3574 975 3575 979
rect 3579 975 3580 979
rect 3574 974 3580 975
rect 3576 955 3578 974
rect 3575 954 3579 955
rect 3575 949 3579 950
rect 3522 935 3528 936
rect 3522 931 3523 935
rect 3527 931 3528 935
rect 3576 934 3578 949
rect 3522 930 3528 931
rect 3574 933 3580 934
rect 3574 929 3575 933
rect 3579 929 3580 933
rect 3574 928 3580 929
rect 3574 916 3580 917
rect 3574 912 3575 916
rect 3579 912 3580 916
rect 3574 911 3580 912
rect 3486 891 3492 892
rect 3486 887 3487 891
rect 3491 887 3492 891
rect 3486 886 3492 887
rect 3576 883 3578 911
rect 1231 882 1235 883
rect 1231 877 1235 878
rect 1359 882 1363 883
rect 1359 877 1363 878
rect 1407 882 1411 883
rect 1407 877 1411 878
rect 1527 882 1531 883
rect 1527 877 1531 878
rect 1583 882 1587 883
rect 1583 877 1587 878
rect 1695 882 1699 883
rect 1695 877 1699 878
rect 1735 882 1739 883
rect 1735 877 1739 878
rect 1823 882 1827 883
rect 1823 877 1827 878
rect 1863 882 1867 883
rect 1863 877 1867 878
rect 2103 882 2107 883
rect 2103 877 2107 878
rect 2151 882 2155 883
rect 2151 877 2155 878
rect 2191 882 2195 883
rect 2191 877 2195 878
rect 2239 882 2243 883
rect 2239 877 2243 878
rect 2279 882 2283 883
rect 2279 877 2283 878
rect 2327 882 2331 883
rect 2327 877 2331 878
rect 2367 882 2371 883
rect 2367 877 2371 878
rect 2415 882 2419 883
rect 2415 877 2419 878
rect 2455 882 2459 883
rect 2455 877 2459 878
rect 2511 882 2515 883
rect 2511 877 2515 878
rect 2567 882 2571 883
rect 2567 877 2571 878
rect 2623 882 2627 883
rect 2682 879 2683 883
rect 2687 879 2688 883
rect 2682 878 2688 879
rect 2703 882 2707 883
rect 2623 877 2627 878
rect 2703 877 2707 878
rect 2759 882 2763 883
rect 2759 877 2763 878
rect 2871 882 2875 883
rect 2871 877 2875 878
rect 2911 882 2915 883
rect 2911 877 2915 878
rect 3055 882 3059 883
rect 3055 877 3059 878
rect 3087 882 3091 883
rect 3087 877 3091 878
rect 3255 882 3259 883
rect 3255 877 3259 878
rect 3271 882 3275 883
rect 3271 877 3275 878
rect 3463 882 3467 883
rect 3463 877 3467 878
rect 3575 882 3579 883
rect 3575 877 3579 878
rect 1360 866 1362 877
rect 1528 866 1530 877
rect 1696 866 1698 877
rect 1358 865 1364 866
rect 1358 861 1359 865
rect 1363 861 1364 865
rect 1190 860 1196 861
rect 1207 860 1211 861
rect 1358 860 1364 861
rect 1526 865 1532 866
rect 1526 861 1527 865
rect 1531 861 1532 865
rect 1694 865 1700 866
rect 1694 861 1695 865
rect 1699 861 1700 865
rect 1526 860 1532 861
rect 1627 860 1631 861
rect 1694 860 1700 861
rect 1207 855 1211 856
rect 1627 855 1631 856
rect 1628 848 1630 855
rect 1824 853 1826 877
rect 1864 853 1866 877
rect 2104 866 2106 877
rect 2192 866 2194 877
rect 2280 866 2282 877
rect 2368 866 2370 877
rect 2438 867 2444 868
rect 2102 865 2108 866
rect 2102 861 2103 865
rect 2107 861 2108 865
rect 2102 860 2108 861
rect 2190 865 2196 866
rect 2190 861 2191 865
rect 2195 861 2196 865
rect 2190 860 2196 861
rect 2278 865 2284 866
rect 2278 861 2279 865
rect 2283 861 2284 865
rect 2278 860 2284 861
rect 2366 865 2372 866
rect 2366 861 2367 865
rect 2371 861 2372 865
rect 2438 863 2439 867
rect 2443 863 2444 867
rect 2456 866 2458 877
rect 2568 866 2570 877
rect 2704 866 2706 877
rect 2872 866 2874 877
rect 3056 866 3058 877
rect 3256 866 3258 877
rect 3464 866 3466 877
rect 3506 875 3512 876
rect 3506 871 3507 875
rect 3511 871 3512 875
rect 3506 870 3512 871
rect 2438 862 2444 863
rect 2454 865 2460 866
rect 2366 860 2372 861
rect 1822 852 1828 853
rect 1822 848 1823 852
rect 1827 848 1828 852
rect 1626 847 1632 848
rect 1822 847 1828 848
rect 1862 852 1868 853
rect 1862 848 1863 852
rect 1867 848 1868 852
rect 1862 847 1868 848
rect 1626 843 1627 847
rect 1631 843 1632 847
rect 1626 842 1632 843
rect 1822 835 1828 836
rect 1822 831 1823 835
rect 1827 831 1828 835
rect 1822 830 1828 831
rect 1862 835 1868 836
rect 1862 831 1863 835
rect 1867 831 1868 835
rect 1862 830 1868 831
rect 1087 828 1091 829
rect 830 825 836 826
rect 830 821 831 825
rect 835 821 836 825
rect 830 820 836 821
rect 1014 825 1020 826
rect 1014 821 1015 825
rect 1019 821 1020 825
rect 1399 828 1403 829
rect 1087 823 1091 824
rect 1182 825 1188 826
rect 1014 820 1020 821
rect 1182 821 1183 825
rect 1187 821 1188 825
rect 1182 820 1188 821
rect 1350 825 1356 826
rect 1350 821 1351 825
rect 1355 821 1356 825
rect 1399 823 1403 824
rect 1518 825 1524 826
rect 1350 820 1356 821
rect 832 815 834 820
rect 1016 815 1018 820
rect 1184 815 1186 820
rect 1352 815 1354 820
rect 831 814 835 815
rect 831 809 835 810
rect 895 814 899 815
rect 895 809 899 810
rect 1015 814 1019 815
rect 1015 809 1019 810
rect 1039 814 1043 815
rect 1039 809 1043 810
rect 1183 814 1187 815
rect 1183 809 1187 810
rect 1327 814 1331 815
rect 1327 809 1331 810
rect 1351 814 1355 815
rect 1351 809 1355 810
rect 896 804 898 809
rect 1040 804 1042 809
rect 1184 804 1186 809
rect 1328 804 1330 809
rect 894 803 900 804
rect 894 799 895 803
rect 899 799 900 803
rect 894 798 900 799
rect 1038 803 1044 804
rect 1038 799 1039 803
rect 1043 799 1044 803
rect 1038 798 1044 799
rect 1182 803 1188 804
rect 1182 799 1183 803
rect 1187 799 1188 803
rect 1182 798 1188 799
rect 1326 803 1332 804
rect 1326 799 1327 803
rect 1331 799 1332 803
rect 1326 798 1332 799
rect 155 796 159 797
rect 751 796 755 797
rect 1400 796 1402 823
rect 1518 821 1519 825
rect 1523 821 1524 825
rect 1518 820 1524 821
rect 1686 825 1692 826
rect 1686 821 1687 825
rect 1691 821 1692 825
rect 1686 820 1692 821
rect 1520 815 1522 820
rect 1688 815 1690 820
rect 1824 815 1826 830
rect 1864 815 1866 830
rect 2094 825 2100 826
rect 2094 821 2095 825
rect 2099 821 2100 825
rect 2094 820 2100 821
rect 2182 825 2188 826
rect 2182 821 2183 825
rect 2187 821 2188 825
rect 2182 820 2188 821
rect 2270 825 2276 826
rect 2270 821 2271 825
rect 2275 821 2276 825
rect 2270 820 2276 821
rect 2358 825 2364 826
rect 2358 821 2359 825
rect 2363 821 2364 825
rect 2358 820 2364 821
rect 2096 815 2098 820
rect 2184 815 2186 820
rect 2272 815 2274 820
rect 2306 819 2312 820
rect 2306 815 2307 819
rect 2311 815 2312 819
rect 2360 815 2362 820
rect 1479 814 1483 815
rect 1479 809 1483 810
rect 1519 814 1523 815
rect 1519 809 1523 810
rect 1687 814 1691 815
rect 1687 809 1691 810
rect 1823 814 1827 815
rect 1823 809 1827 810
rect 1863 814 1867 815
rect 1863 809 1867 810
rect 2095 814 2099 815
rect 2095 809 2099 810
rect 2183 814 2187 815
rect 2183 809 2187 810
rect 2199 814 2203 815
rect 2199 809 2203 810
rect 2271 814 2275 815
rect 2271 809 2275 810
rect 2287 814 2291 815
rect 2306 814 2312 815
rect 2359 814 2363 815
rect 2287 809 2291 810
rect 1480 804 1482 809
rect 1478 803 1484 804
rect 1478 799 1479 803
rect 1483 799 1484 803
rect 1478 798 1484 799
rect 110 793 116 794
rect 110 789 111 793
rect 115 789 116 793
rect 155 791 159 792
rect 678 795 684 796
rect 678 791 679 795
rect 683 791 684 795
rect 751 791 755 792
rect 1398 795 1404 796
rect 1398 791 1399 795
rect 1403 791 1404 795
rect 1824 794 1826 809
rect 1864 794 1866 809
rect 2200 804 2202 809
rect 2288 804 2290 809
rect 2198 803 2204 804
rect 2198 799 2199 803
rect 2203 799 2204 803
rect 2198 798 2204 799
rect 2286 803 2292 804
rect 2286 799 2287 803
rect 2291 799 2292 803
rect 2286 798 2292 799
rect 110 788 116 789
rect 110 776 116 777
rect 110 772 111 776
rect 115 772 116 776
rect 110 771 116 772
rect 112 743 114 771
rect 142 763 148 764
rect 142 759 143 763
rect 147 759 148 763
rect 142 758 148 759
rect 144 743 146 758
rect 156 752 158 791
rect 678 790 684 791
rect 1398 790 1404 791
rect 1822 793 1828 794
rect 278 763 284 764
rect 278 759 279 763
rect 283 759 284 763
rect 278 758 284 759
rect 430 763 436 764
rect 430 759 431 763
rect 435 759 436 763
rect 430 758 436 759
rect 590 763 596 764
rect 590 759 591 763
rect 595 759 596 763
rect 590 758 596 759
rect 154 751 160 752
rect 154 747 155 751
rect 159 747 160 751
rect 154 746 160 747
rect 280 743 282 758
rect 371 756 375 757
rect 371 751 375 752
rect 111 742 115 743
rect 111 737 115 738
rect 143 742 147 743
rect 143 737 147 738
rect 279 742 283 743
rect 279 737 283 738
rect 359 742 363 743
rect 359 737 363 738
rect 112 713 114 737
rect 360 726 362 737
rect 372 736 374 751
rect 432 743 434 758
rect 592 743 594 758
rect 680 757 682 790
rect 1822 789 1823 793
rect 1827 789 1828 793
rect 1822 788 1828 789
rect 1862 793 1868 794
rect 1862 789 1863 793
rect 1867 789 1868 793
rect 1862 788 1868 789
rect 2266 779 2272 780
rect 1822 776 1828 777
rect 1822 772 1823 776
rect 1827 772 1828 776
rect 1822 771 1828 772
rect 1862 776 1868 777
rect 1862 772 1863 776
rect 1867 772 1868 776
rect 2266 775 2267 779
rect 2271 775 2272 779
rect 2266 774 2272 775
rect 1862 771 1868 772
rect 750 763 756 764
rect 750 759 751 763
rect 755 759 756 763
rect 750 758 756 759
rect 902 763 908 764
rect 902 759 903 763
rect 907 759 908 763
rect 902 758 908 759
rect 1046 763 1052 764
rect 1046 759 1047 763
rect 1051 759 1052 763
rect 1046 758 1052 759
rect 1190 763 1196 764
rect 1190 759 1191 763
rect 1195 759 1196 763
rect 1190 758 1196 759
rect 1334 763 1340 764
rect 1334 759 1335 763
rect 1339 759 1340 763
rect 1334 758 1340 759
rect 1486 763 1492 764
rect 1486 759 1487 763
rect 1491 759 1492 763
rect 1486 758 1492 759
rect 679 756 683 757
rect 679 751 683 752
rect 752 743 754 758
rect 904 743 906 758
rect 1022 751 1028 752
rect 1022 747 1023 751
rect 1027 747 1028 751
rect 1022 746 1028 747
rect 431 742 435 743
rect 431 737 435 738
rect 447 742 451 743
rect 447 737 451 738
rect 543 742 547 743
rect 543 737 547 738
rect 591 742 595 743
rect 591 737 595 738
rect 639 742 643 743
rect 639 737 643 738
rect 735 742 739 743
rect 735 737 739 738
rect 751 742 755 743
rect 751 737 755 738
rect 831 742 835 743
rect 831 737 835 738
rect 903 742 907 743
rect 903 737 907 738
rect 927 742 931 743
rect 927 737 931 738
rect 370 735 376 736
rect 370 731 371 735
rect 375 731 376 735
rect 370 730 376 731
rect 448 726 450 737
rect 544 726 546 737
rect 640 726 642 737
rect 736 726 738 737
rect 832 726 834 737
rect 898 727 904 728
rect 358 725 364 726
rect 358 721 359 725
rect 363 721 364 725
rect 358 720 364 721
rect 446 725 452 726
rect 446 721 447 725
rect 451 721 452 725
rect 446 720 452 721
rect 542 725 548 726
rect 542 721 543 725
rect 547 721 548 725
rect 542 720 548 721
rect 638 725 644 726
rect 638 721 639 725
rect 643 721 644 725
rect 638 720 644 721
rect 734 725 740 726
rect 734 721 735 725
rect 739 721 740 725
rect 734 720 740 721
rect 830 725 836 726
rect 830 721 831 725
rect 835 721 836 725
rect 898 723 899 727
rect 903 723 904 727
rect 928 726 930 737
rect 1024 733 1026 746
rect 1048 743 1050 758
rect 1192 743 1194 758
rect 1336 743 1338 758
rect 1488 743 1490 758
rect 1824 743 1826 771
rect 1864 743 1866 771
rect 2206 763 2212 764
rect 2206 759 2207 763
rect 2211 759 2212 763
rect 2206 758 2212 759
rect 2208 743 2210 758
rect 1031 742 1035 743
rect 1031 737 1035 738
rect 1047 742 1051 743
rect 1047 737 1051 738
rect 1135 742 1139 743
rect 1135 737 1139 738
rect 1191 742 1195 743
rect 1191 737 1195 738
rect 1239 742 1243 743
rect 1239 737 1243 738
rect 1335 742 1339 743
rect 1335 737 1339 738
rect 1487 742 1491 743
rect 1487 737 1491 738
rect 1823 742 1827 743
rect 1823 737 1827 738
rect 1863 742 1867 743
rect 1863 737 1867 738
rect 1943 742 1947 743
rect 1943 737 1947 738
rect 2103 742 2107 743
rect 2103 737 2107 738
rect 2207 742 2211 743
rect 2207 737 2211 738
rect 2255 742 2259 743
rect 2255 737 2259 738
rect 1023 732 1027 733
rect 1023 727 1027 728
rect 1032 726 1034 737
rect 1136 726 1138 737
rect 1203 732 1207 733
rect 1203 727 1207 728
rect 898 722 904 723
rect 926 725 932 726
rect 830 720 836 721
rect 110 712 116 713
rect 110 708 111 712
rect 115 708 116 712
rect 110 707 116 708
rect 110 695 116 696
rect 110 691 111 695
rect 115 691 116 695
rect 110 690 116 691
rect 112 671 114 690
rect 350 685 356 686
rect 350 681 351 685
rect 355 681 356 685
rect 350 680 356 681
rect 438 685 444 686
rect 438 681 439 685
rect 443 681 444 685
rect 438 680 444 681
rect 534 685 540 686
rect 534 681 535 685
rect 539 681 540 685
rect 534 680 540 681
rect 630 685 636 686
rect 630 681 631 685
rect 635 681 636 685
rect 630 680 636 681
rect 726 685 732 686
rect 726 681 727 685
rect 731 681 732 685
rect 726 680 732 681
rect 822 685 828 686
rect 822 681 823 685
rect 827 681 828 685
rect 822 680 828 681
rect 352 671 354 680
rect 440 671 442 680
rect 510 679 516 680
rect 510 675 511 679
rect 515 675 516 679
rect 510 674 516 675
rect 111 670 115 671
rect 111 665 115 666
rect 351 670 355 671
rect 351 665 355 666
rect 439 670 443 671
rect 439 665 443 666
rect 479 670 483 671
rect 479 665 483 666
rect 112 650 114 665
rect 480 660 482 665
rect 478 659 484 660
rect 478 655 479 659
rect 483 655 484 659
rect 478 654 484 655
rect 110 649 116 650
rect 110 645 111 649
rect 115 645 116 649
rect 110 644 116 645
rect 110 632 116 633
rect 110 628 111 632
rect 115 628 116 632
rect 110 627 116 628
rect 112 603 114 627
rect 486 619 492 620
rect 486 615 487 619
rect 491 615 492 619
rect 486 614 492 615
rect 488 603 490 614
rect 512 608 514 674
rect 536 671 538 680
rect 632 671 634 680
rect 728 671 730 680
rect 824 671 826 680
rect 535 670 539 671
rect 535 665 539 666
rect 567 670 571 671
rect 567 665 571 666
rect 631 670 635 671
rect 631 665 635 666
rect 655 670 659 671
rect 655 665 659 666
rect 727 670 731 671
rect 727 665 731 666
rect 743 670 747 671
rect 743 665 747 666
rect 823 670 827 671
rect 823 665 827 666
rect 831 670 835 671
rect 831 665 835 666
rect 568 660 570 665
rect 656 660 658 665
rect 744 660 746 665
rect 832 660 834 665
rect 566 659 572 660
rect 566 655 567 659
rect 571 655 572 659
rect 566 654 572 655
rect 654 659 660 660
rect 654 655 655 659
rect 659 655 660 659
rect 654 654 660 655
rect 742 659 748 660
rect 742 655 743 659
rect 747 655 748 659
rect 742 654 748 655
rect 830 659 836 660
rect 830 655 831 659
rect 835 655 836 659
rect 830 654 836 655
rect 900 652 902 722
rect 926 721 927 725
rect 931 721 932 725
rect 926 720 932 721
rect 1030 725 1036 726
rect 1030 721 1031 725
rect 1035 721 1036 725
rect 1030 720 1036 721
rect 1134 725 1140 726
rect 1134 721 1135 725
rect 1139 721 1140 725
rect 1134 720 1140 721
rect 1204 696 1206 727
rect 1240 726 1242 737
rect 1238 725 1244 726
rect 1238 721 1239 725
rect 1243 721 1244 725
rect 1238 720 1244 721
rect 1824 713 1826 737
rect 1864 713 1866 737
rect 1944 726 1946 737
rect 2046 735 2052 736
rect 2046 731 2047 735
rect 2051 731 2052 735
rect 2046 730 2052 731
rect 1942 725 1948 726
rect 1942 721 1943 725
rect 1947 721 1948 725
rect 1942 720 1948 721
rect 1822 712 1828 713
rect 1822 708 1823 712
rect 1827 708 1828 712
rect 1822 707 1828 708
rect 1862 712 1868 713
rect 1862 708 1863 712
rect 1867 708 1868 712
rect 2048 708 2050 730
rect 2104 726 2106 737
rect 2114 735 2120 736
rect 2114 731 2115 735
rect 2119 731 2120 735
rect 2114 730 2120 731
rect 2102 725 2108 726
rect 2102 721 2103 725
rect 2107 721 2108 725
rect 2102 720 2108 721
rect 1862 707 1868 708
rect 2046 707 2052 708
rect 2046 703 2047 707
rect 2051 703 2052 707
rect 2046 702 2052 703
rect 1202 695 1208 696
rect 1202 691 1203 695
rect 1207 691 1208 695
rect 1202 690 1208 691
rect 1822 695 1828 696
rect 1822 691 1823 695
rect 1827 691 1828 695
rect 1822 690 1828 691
rect 1862 695 1868 696
rect 1862 691 1863 695
rect 1867 691 1868 695
rect 1862 690 1868 691
rect 1906 695 1912 696
rect 1906 691 1907 695
rect 1911 691 1912 695
rect 1906 690 1912 691
rect 918 685 924 686
rect 918 681 919 685
rect 923 681 924 685
rect 918 680 924 681
rect 1022 685 1028 686
rect 1022 681 1023 685
rect 1027 681 1028 685
rect 1022 680 1028 681
rect 1126 685 1132 686
rect 1126 681 1127 685
rect 1131 681 1132 685
rect 1126 680 1132 681
rect 1230 685 1236 686
rect 1230 681 1231 685
rect 1235 681 1236 685
rect 1230 680 1236 681
rect 920 671 922 680
rect 1024 671 1026 680
rect 1128 671 1130 680
rect 1232 671 1234 680
rect 1824 671 1826 690
rect 1864 671 1866 690
rect 919 670 923 671
rect 919 665 923 666
rect 1007 670 1011 671
rect 1007 665 1011 666
rect 1023 670 1027 671
rect 1023 665 1027 666
rect 1095 670 1099 671
rect 1095 665 1099 666
rect 1127 670 1131 671
rect 1127 665 1131 666
rect 1183 670 1187 671
rect 1183 665 1187 666
rect 1231 670 1235 671
rect 1231 665 1235 666
rect 1271 670 1275 671
rect 1271 665 1275 666
rect 1823 670 1827 671
rect 1823 665 1827 666
rect 1863 670 1867 671
rect 1863 665 1867 666
rect 1887 670 1891 671
rect 1887 665 1891 666
rect 920 660 922 665
rect 1008 660 1010 665
rect 1096 660 1098 665
rect 1184 660 1186 665
rect 1272 660 1274 665
rect 918 659 924 660
rect 918 655 919 659
rect 923 655 924 659
rect 918 654 924 655
rect 1006 659 1012 660
rect 1006 655 1007 659
rect 1011 655 1012 659
rect 1006 654 1012 655
rect 1094 659 1100 660
rect 1094 655 1095 659
rect 1099 655 1100 659
rect 1094 654 1100 655
rect 1182 659 1188 660
rect 1182 655 1183 659
rect 1187 655 1188 659
rect 1182 654 1188 655
rect 1270 659 1276 660
rect 1270 655 1271 659
rect 1275 655 1276 659
rect 1270 654 1276 655
rect 898 651 904 652
rect 898 647 899 651
rect 903 647 904 651
rect 1824 650 1826 665
rect 1864 650 1866 665
rect 1888 660 1890 665
rect 1886 659 1892 660
rect 1886 655 1887 659
rect 1891 655 1892 659
rect 1886 654 1892 655
rect 898 646 904 647
rect 1822 649 1828 650
rect 1822 645 1823 649
rect 1827 645 1828 649
rect 1822 644 1828 645
rect 1862 649 1868 650
rect 1862 645 1863 649
rect 1867 645 1868 649
rect 1862 644 1868 645
rect 986 635 992 636
rect 986 631 987 635
rect 991 631 992 635
rect 986 630 992 631
rect 1074 635 1080 636
rect 1074 631 1075 635
rect 1079 631 1080 635
rect 1074 630 1080 631
rect 1250 635 1256 636
rect 1250 631 1251 635
rect 1255 631 1256 635
rect 1250 630 1256 631
rect 1822 632 1828 633
rect 574 619 580 620
rect 574 615 575 619
rect 579 615 580 619
rect 574 614 580 615
rect 662 619 668 620
rect 662 615 663 619
rect 667 615 668 619
rect 662 614 668 615
rect 750 619 756 620
rect 750 615 751 619
rect 755 615 756 619
rect 750 614 756 615
rect 838 619 844 620
rect 838 615 839 619
rect 843 615 844 619
rect 838 614 844 615
rect 926 619 932 620
rect 926 615 927 619
rect 931 615 932 619
rect 926 614 932 615
rect 510 607 516 608
rect 510 603 511 607
rect 515 603 516 607
rect 576 603 578 614
rect 664 603 666 614
rect 752 603 754 614
rect 840 603 842 614
rect 928 603 930 614
rect 988 608 990 630
rect 1014 619 1020 620
rect 1014 615 1015 619
rect 1019 615 1020 619
rect 1014 614 1020 615
rect 986 607 992 608
rect 986 603 987 607
rect 991 603 992 607
rect 1016 603 1018 614
rect 1076 608 1078 630
rect 1102 619 1108 620
rect 1102 615 1103 619
rect 1107 615 1108 619
rect 1102 614 1108 615
rect 1190 619 1196 620
rect 1190 615 1191 619
rect 1195 615 1196 619
rect 1190 614 1196 615
rect 1074 607 1080 608
rect 1074 603 1075 607
rect 1079 603 1080 607
rect 1104 603 1106 614
rect 1192 603 1194 614
rect 1252 608 1254 630
rect 1822 628 1823 632
rect 1827 628 1828 632
rect 1822 627 1828 628
rect 1862 632 1868 633
rect 1862 628 1863 632
rect 1867 628 1868 632
rect 1862 627 1868 628
rect 1278 619 1284 620
rect 1278 615 1279 619
rect 1283 615 1284 619
rect 1278 614 1284 615
rect 1250 607 1256 608
rect 1250 603 1251 607
rect 1255 603 1256 607
rect 1280 603 1282 614
rect 1824 603 1826 627
rect 1864 603 1866 627
rect 1894 619 1900 620
rect 1894 615 1895 619
rect 1899 615 1900 619
rect 1894 614 1900 615
rect 1896 603 1898 614
rect 1908 608 1910 690
rect 1934 685 1940 686
rect 1934 681 1935 685
rect 1939 681 1940 685
rect 1934 680 1940 681
rect 2094 685 2100 686
rect 2094 681 2095 685
rect 2099 681 2100 685
rect 2094 680 2100 681
rect 1936 671 1938 680
rect 2096 671 2098 680
rect 1935 670 1939 671
rect 1935 665 1939 666
rect 2023 670 2027 671
rect 2023 665 2027 666
rect 2095 670 2099 671
rect 2116 668 2118 730
rect 2256 726 2258 737
rect 2268 736 2270 774
rect 2294 763 2300 764
rect 2294 759 2295 763
rect 2299 759 2300 763
rect 2294 758 2300 759
rect 2296 743 2298 758
rect 2308 752 2310 814
rect 2359 809 2363 810
rect 2375 814 2379 815
rect 2375 809 2379 810
rect 2376 804 2378 809
rect 2374 803 2380 804
rect 2374 799 2375 803
rect 2379 799 2380 803
rect 2440 803 2442 862
rect 2454 861 2455 865
rect 2459 861 2460 865
rect 2454 860 2460 861
rect 2566 865 2572 866
rect 2566 861 2567 865
rect 2571 861 2572 865
rect 2566 860 2572 861
rect 2702 865 2708 866
rect 2702 861 2703 865
rect 2707 861 2708 865
rect 2702 860 2708 861
rect 2870 865 2876 866
rect 2870 861 2871 865
rect 2875 861 2876 865
rect 2870 860 2876 861
rect 3054 865 3060 866
rect 3054 861 3055 865
rect 3059 861 3060 865
rect 3054 860 3060 861
rect 3254 865 3260 866
rect 3254 861 3255 865
rect 3259 861 3260 865
rect 3254 860 3260 861
rect 3462 865 3468 866
rect 3462 861 3463 865
rect 3467 861 3468 865
rect 3462 860 3468 861
rect 3138 835 3144 836
rect 3138 831 3139 835
rect 3143 831 3144 835
rect 3138 830 3144 831
rect 2446 825 2452 826
rect 2446 821 2447 825
rect 2451 821 2452 825
rect 2446 820 2452 821
rect 2558 825 2564 826
rect 2558 821 2559 825
rect 2563 821 2564 825
rect 2558 820 2564 821
rect 2694 825 2700 826
rect 2694 821 2695 825
rect 2699 821 2700 825
rect 2694 820 2700 821
rect 2862 825 2868 826
rect 2862 821 2863 825
rect 2867 821 2868 825
rect 2862 820 2868 821
rect 3046 825 3052 826
rect 3046 821 3047 825
rect 3051 821 3052 825
rect 3046 820 3052 821
rect 2448 815 2450 820
rect 2560 815 2562 820
rect 2696 815 2698 820
rect 2864 815 2866 820
rect 3048 815 3050 820
rect 2447 814 2451 815
rect 2447 809 2451 810
rect 2463 814 2467 815
rect 2463 809 2467 810
rect 2551 814 2555 815
rect 2551 809 2555 810
rect 2559 814 2563 815
rect 2559 809 2563 810
rect 2655 814 2659 815
rect 2655 809 2659 810
rect 2695 814 2699 815
rect 2695 809 2699 810
rect 2783 814 2787 815
rect 2783 809 2787 810
rect 2863 814 2867 815
rect 2863 809 2867 810
rect 2935 814 2939 815
rect 2935 809 2939 810
rect 3047 814 3051 815
rect 3047 809 3051 810
rect 3111 814 3115 815
rect 3111 809 3115 810
rect 2464 804 2466 809
rect 2552 804 2554 809
rect 2656 804 2658 809
rect 2784 804 2786 809
rect 2936 804 2938 809
rect 3112 804 3114 809
rect 2462 803 2468 804
rect 2440 801 2446 803
rect 2374 798 2380 799
rect 2444 796 2446 801
rect 2462 799 2463 803
rect 2467 799 2468 803
rect 2462 798 2468 799
rect 2550 803 2556 804
rect 2550 799 2551 803
rect 2555 799 2556 803
rect 2550 798 2556 799
rect 2654 803 2660 804
rect 2654 799 2655 803
rect 2659 799 2660 803
rect 2654 798 2660 799
rect 2782 803 2788 804
rect 2782 799 2783 803
rect 2787 799 2788 803
rect 2782 798 2788 799
rect 2934 803 2940 804
rect 2934 799 2935 803
rect 2939 799 2940 803
rect 2934 798 2940 799
rect 3110 803 3116 804
rect 3110 799 3111 803
rect 3115 799 3116 803
rect 3110 798 3116 799
rect 2354 795 2360 796
rect 2354 791 2355 795
rect 2359 791 2360 795
rect 2354 790 2360 791
rect 2442 795 2448 796
rect 2442 791 2443 795
rect 2447 791 2448 795
rect 2442 790 2448 791
rect 2306 751 2312 752
rect 2306 747 2307 751
rect 2311 747 2312 751
rect 2306 746 2312 747
rect 2356 744 2358 790
rect 2530 779 2536 780
rect 2530 775 2531 779
rect 2535 775 2536 779
rect 2530 774 2536 775
rect 2382 763 2388 764
rect 2382 759 2383 763
rect 2387 759 2388 763
rect 2382 758 2388 759
rect 2470 763 2476 764
rect 2470 759 2471 763
rect 2475 759 2476 763
rect 2470 758 2476 759
rect 2354 743 2360 744
rect 2384 743 2386 758
rect 2472 743 2474 758
rect 2532 752 2534 774
rect 2707 772 2711 773
rect 2707 767 2711 768
rect 2558 763 2564 764
rect 2558 759 2559 763
rect 2563 759 2564 763
rect 2558 758 2564 759
rect 2662 763 2668 764
rect 2662 759 2663 763
rect 2667 759 2668 763
rect 2662 758 2668 759
rect 2530 751 2536 752
rect 2530 747 2531 751
rect 2535 747 2536 751
rect 2530 746 2536 747
rect 2560 743 2562 758
rect 2610 751 2616 752
rect 2610 747 2611 751
rect 2615 747 2616 751
rect 2610 746 2616 747
rect 2295 742 2299 743
rect 2354 739 2355 743
rect 2359 739 2360 743
rect 2354 738 2360 739
rect 2383 742 2387 743
rect 2295 737 2299 738
rect 2383 737 2387 738
rect 2407 742 2411 743
rect 2407 737 2411 738
rect 2471 742 2475 743
rect 2471 737 2475 738
rect 2551 742 2555 743
rect 2551 737 2555 738
rect 2559 742 2563 743
rect 2559 737 2563 738
rect 2266 735 2272 736
rect 2266 731 2267 735
rect 2271 731 2272 735
rect 2266 730 2272 731
rect 2408 726 2410 737
rect 2552 726 2554 737
rect 2254 725 2260 726
rect 2254 721 2255 725
rect 2259 721 2260 725
rect 2254 720 2260 721
rect 2406 725 2412 726
rect 2406 721 2407 725
rect 2411 721 2412 725
rect 2406 720 2412 721
rect 2550 725 2556 726
rect 2550 721 2551 725
rect 2555 721 2556 725
rect 2550 720 2556 721
rect 2612 712 2614 746
rect 2664 743 2666 758
rect 2675 756 2679 757
rect 2674 751 2680 752
rect 2674 747 2675 751
rect 2679 747 2680 751
rect 2674 746 2680 747
rect 2663 742 2667 743
rect 2663 737 2667 738
rect 2695 742 2699 743
rect 2695 737 2699 738
rect 2696 726 2698 737
rect 2708 736 2710 767
rect 2790 763 2796 764
rect 2790 759 2791 763
rect 2795 759 2796 763
rect 2790 758 2796 759
rect 2942 763 2948 764
rect 2942 759 2943 763
rect 2947 759 2948 763
rect 2942 758 2948 759
rect 3118 763 3124 764
rect 3118 759 3119 763
rect 3123 759 3124 763
rect 3118 758 3124 759
rect 2792 743 2794 758
rect 2944 743 2946 758
rect 3120 743 3122 758
rect 3140 757 3142 830
rect 3246 825 3252 826
rect 3246 821 3247 825
rect 3251 821 3252 825
rect 3246 820 3252 821
rect 3454 825 3460 826
rect 3454 821 3455 825
rect 3459 821 3460 825
rect 3454 820 3460 821
rect 3248 815 3250 820
rect 3456 815 3458 820
rect 3498 819 3504 820
rect 3498 815 3499 819
rect 3503 815 3504 819
rect 3247 814 3251 815
rect 3247 809 3251 810
rect 3295 814 3299 815
rect 3295 809 3299 810
rect 3455 814 3459 815
rect 3455 809 3459 810
rect 3479 814 3483 815
rect 3498 814 3504 815
rect 3479 809 3483 810
rect 3296 804 3298 809
rect 3480 804 3482 809
rect 3294 803 3300 804
rect 3294 799 3295 803
rect 3299 799 3300 803
rect 3294 798 3300 799
rect 3478 803 3484 804
rect 3478 799 3479 803
rect 3483 799 3484 803
rect 3478 798 3484 799
rect 3198 795 3204 796
rect 3198 791 3199 795
rect 3203 791 3204 795
rect 3198 790 3204 791
rect 3200 773 3202 790
rect 3470 779 3476 780
rect 3470 775 3471 779
rect 3475 775 3476 779
rect 3470 774 3476 775
rect 3199 772 3203 773
rect 3199 767 3203 768
rect 3302 763 3308 764
rect 3302 759 3303 763
rect 3307 759 3308 763
rect 3302 758 3308 759
rect 3139 756 3143 757
rect 3139 751 3143 752
rect 3304 743 3306 758
rect 2791 742 2795 743
rect 2791 737 2795 738
rect 2839 742 2843 743
rect 2839 737 2843 738
rect 2943 742 2947 743
rect 2943 737 2947 738
rect 2983 742 2987 743
rect 2983 737 2987 738
rect 3119 742 3123 743
rect 3119 737 3123 738
rect 3135 742 3139 743
rect 3135 737 3139 738
rect 3287 742 3291 743
rect 3287 737 3291 738
rect 3303 742 3307 743
rect 3303 737 3307 738
rect 3439 742 3443 743
rect 3439 737 3443 738
rect 2706 735 2712 736
rect 2706 731 2707 735
rect 2711 731 2712 735
rect 2706 730 2712 731
rect 2840 726 2842 737
rect 2984 726 2986 737
rect 3136 726 3138 737
rect 3190 735 3196 736
rect 3190 731 3191 735
rect 3195 731 3196 735
rect 3190 730 3196 731
rect 2694 725 2700 726
rect 2694 721 2695 725
rect 2699 721 2700 725
rect 2694 720 2700 721
rect 2838 725 2844 726
rect 2838 721 2839 725
rect 2843 721 2844 725
rect 2838 720 2844 721
rect 2982 725 2988 726
rect 2982 721 2983 725
rect 2987 721 2988 725
rect 2982 720 2988 721
rect 3134 725 3140 726
rect 3134 721 3135 725
rect 3139 721 3140 725
rect 3134 720 3140 721
rect 2610 711 2616 712
rect 2610 707 2611 711
rect 2615 707 2616 711
rect 2610 706 2616 707
rect 3078 695 3084 696
rect 3078 691 3079 695
rect 3083 691 3084 695
rect 3078 690 3084 691
rect 2246 685 2252 686
rect 2246 681 2247 685
rect 2251 681 2252 685
rect 2246 680 2252 681
rect 2398 685 2404 686
rect 2398 681 2399 685
rect 2403 681 2404 685
rect 2398 680 2404 681
rect 2542 685 2548 686
rect 2542 681 2543 685
rect 2547 681 2548 685
rect 2542 680 2548 681
rect 2686 685 2692 686
rect 2686 681 2687 685
rect 2691 681 2692 685
rect 2686 680 2692 681
rect 2830 685 2836 686
rect 2830 681 2831 685
rect 2835 681 2836 685
rect 2830 680 2836 681
rect 2974 685 2980 686
rect 2974 681 2975 685
rect 2979 681 2980 685
rect 2974 680 2980 681
rect 2248 671 2250 680
rect 2400 671 2402 680
rect 2544 671 2546 680
rect 2688 671 2690 680
rect 2832 671 2834 680
rect 2976 671 2978 680
rect 2199 670 2203 671
rect 2095 665 2099 666
rect 2114 667 2120 668
rect 2024 660 2026 665
rect 2114 663 2115 667
rect 2119 663 2120 667
rect 2199 665 2203 666
rect 2247 670 2251 671
rect 2247 665 2251 666
rect 2383 670 2387 671
rect 2383 665 2387 666
rect 2399 670 2403 671
rect 2399 665 2403 666
rect 2543 670 2547 671
rect 2543 665 2547 666
rect 2567 670 2571 671
rect 2567 665 2571 666
rect 2687 670 2691 671
rect 2687 665 2691 666
rect 2743 670 2747 671
rect 2743 665 2747 666
rect 2831 670 2835 671
rect 2831 665 2835 666
rect 2911 670 2915 671
rect 2911 665 2915 666
rect 2975 670 2979 671
rect 2975 665 2979 666
rect 3063 670 3067 671
rect 3063 665 3067 666
rect 2114 662 2120 663
rect 2200 660 2202 665
rect 2384 660 2386 665
rect 2568 660 2570 665
rect 2744 660 2746 665
rect 2912 660 2914 665
rect 3064 660 3066 665
rect 2022 659 2028 660
rect 2022 655 2023 659
rect 2027 655 2028 659
rect 2022 654 2028 655
rect 2198 659 2204 660
rect 2198 655 2199 659
rect 2203 655 2204 659
rect 2198 654 2204 655
rect 2382 659 2388 660
rect 2382 655 2383 659
rect 2387 655 2388 659
rect 2382 654 2388 655
rect 2566 659 2572 660
rect 2566 655 2567 659
rect 2571 655 2572 659
rect 2566 654 2572 655
rect 2742 659 2748 660
rect 2742 655 2743 659
rect 2747 655 2748 659
rect 2742 654 2748 655
rect 2910 659 2916 660
rect 2910 655 2911 659
rect 2915 655 2916 659
rect 2910 654 2916 655
rect 3062 659 3068 660
rect 3062 655 3063 659
rect 3067 655 3068 659
rect 3062 654 3068 655
rect 2098 651 2104 652
rect 2098 647 2099 651
rect 2103 647 2104 651
rect 2098 646 2104 647
rect 2030 619 2036 620
rect 2030 615 2031 619
rect 2035 615 2036 619
rect 2030 614 2036 615
rect 1906 607 1912 608
rect 1906 603 1907 607
rect 1911 603 1912 607
rect 2032 603 2034 614
rect 111 602 115 603
rect 111 597 115 598
rect 487 602 491 603
rect 487 597 491 598
rect 503 602 507 603
rect 510 602 516 603
rect 575 602 579 603
rect 503 597 507 598
rect 575 597 579 598
rect 599 602 603 603
rect 599 597 603 598
rect 663 602 667 603
rect 663 597 667 598
rect 703 602 707 603
rect 703 597 707 598
rect 751 602 755 603
rect 751 597 755 598
rect 815 602 819 603
rect 815 597 819 598
rect 839 602 843 603
rect 839 597 843 598
rect 927 602 931 603
rect 927 597 931 598
rect 935 602 939 603
rect 986 602 992 603
rect 1015 602 1019 603
rect 935 597 939 598
rect 1015 597 1019 598
rect 1063 602 1067 603
rect 1074 602 1080 603
rect 1103 602 1107 603
rect 1063 597 1067 598
rect 1103 597 1107 598
rect 1191 602 1195 603
rect 1250 602 1256 603
rect 1279 602 1283 603
rect 1191 597 1195 598
rect 1279 597 1283 598
rect 1327 602 1331 603
rect 1327 597 1331 598
rect 1471 602 1475 603
rect 1471 597 1475 598
rect 1615 602 1619 603
rect 1615 597 1619 598
rect 1735 602 1739 603
rect 1735 597 1739 598
rect 1823 602 1827 603
rect 1823 597 1827 598
rect 1863 602 1867 603
rect 1863 597 1867 598
rect 1895 602 1899 603
rect 1906 602 1912 603
rect 2031 602 2035 603
rect 1895 597 1899 598
rect 2031 597 2035 598
rect 2087 602 2091 603
rect 2087 597 2091 598
rect 112 573 114 597
rect 504 586 506 597
rect 558 595 564 596
rect 558 591 559 595
rect 563 591 564 595
rect 558 590 564 591
rect 502 585 508 586
rect 502 581 503 585
rect 507 581 508 585
rect 502 580 508 581
rect 560 573 562 590
rect 600 586 602 597
rect 704 586 706 597
rect 816 586 818 597
rect 886 595 892 596
rect 886 591 887 595
rect 891 591 892 595
rect 886 590 892 591
rect 598 585 604 586
rect 598 581 599 585
rect 603 581 604 585
rect 598 580 604 581
rect 702 585 708 586
rect 702 581 703 585
rect 707 581 708 585
rect 702 580 708 581
rect 814 585 820 586
rect 814 581 815 585
rect 819 581 820 585
rect 814 580 820 581
rect 110 572 116 573
rect 110 568 111 572
rect 115 568 116 572
rect 110 567 116 568
rect 559 572 563 573
rect 771 572 775 573
rect 888 568 890 590
rect 936 586 938 597
rect 1026 595 1032 596
rect 1026 591 1027 595
rect 1031 591 1032 595
rect 1026 590 1032 591
rect 934 585 940 586
rect 934 581 935 585
rect 939 581 940 585
rect 934 580 940 581
rect 559 567 563 568
rect 770 567 776 568
rect 770 563 771 567
rect 775 563 776 567
rect 770 562 776 563
rect 886 567 892 568
rect 886 563 887 567
rect 891 563 892 567
rect 886 562 892 563
rect 110 555 116 556
rect 110 551 111 555
rect 115 551 116 555
rect 110 550 116 551
rect 814 555 820 556
rect 814 551 815 555
rect 819 551 820 555
rect 814 550 820 551
rect 112 535 114 550
rect 494 545 500 546
rect 494 541 495 545
rect 499 541 500 545
rect 494 540 500 541
rect 590 545 596 546
rect 590 541 591 545
rect 595 541 596 545
rect 590 540 596 541
rect 694 545 700 546
rect 694 541 695 545
rect 699 541 700 545
rect 694 540 700 541
rect 806 545 812 546
rect 806 541 807 545
rect 811 541 812 545
rect 806 540 812 541
rect 496 535 498 540
rect 592 535 594 540
rect 696 535 698 540
rect 808 535 810 540
rect 111 534 115 535
rect 111 529 115 530
rect 159 534 163 535
rect 159 529 163 530
rect 303 534 307 535
rect 303 529 307 530
rect 463 534 467 535
rect 463 529 467 530
rect 495 534 499 535
rect 495 529 499 530
rect 591 534 595 535
rect 591 529 595 530
rect 631 534 635 535
rect 631 529 635 530
rect 695 534 699 535
rect 695 529 699 530
rect 799 534 803 535
rect 799 529 803 530
rect 807 534 811 535
rect 807 529 811 530
rect 112 514 114 529
rect 160 524 162 529
rect 304 524 306 529
rect 464 524 466 529
rect 632 524 634 529
rect 800 524 802 529
rect 158 523 164 524
rect 158 519 159 523
rect 163 519 164 523
rect 158 518 164 519
rect 302 523 308 524
rect 302 519 303 523
rect 307 519 308 523
rect 302 518 308 519
rect 462 523 468 524
rect 462 519 463 523
rect 467 519 468 523
rect 462 518 468 519
rect 630 523 636 524
rect 630 519 631 523
rect 635 519 636 523
rect 630 518 636 519
rect 798 523 804 524
rect 798 519 799 523
rect 803 519 804 523
rect 798 518 804 519
rect 110 513 116 514
rect 110 509 111 513
rect 115 509 116 513
rect 110 508 116 509
rect 150 499 156 500
rect 110 496 116 497
rect 110 492 111 496
rect 115 492 116 496
rect 150 495 151 499
rect 155 495 156 499
rect 150 494 156 495
rect 226 499 232 500
rect 226 495 227 499
rect 231 495 232 499
rect 226 494 232 495
rect 370 499 376 500
rect 370 495 371 499
rect 375 495 376 499
rect 370 494 376 495
rect 530 499 536 500
rect 530 495 531 499
rect 535 495 536 499
rect 530 494 536 495
rect 698 499 704 500
rect 698 495 699 499
rect 703 495 704 499
rect 698 494 704 495
rect 110 491 116 492
rect 112 459 114 491
rect 111 458 115 459
rect 111 453 115 454
rect 143 458 147 459
rect 143 453 147 454
rect 112 429 114 453
rect 144 442 146 453
rect 152 452 154 494
rect 166 483 172 484
rect 166 479 167 483
rect 171 479 172 483
rect 166 478 172 479
rect 168 459 170 478
rect 228 472 230 494
rect 310 483 316 484
rect 310 479 311 483
rect 315 479 316 483
rect 310 478 316 479
rect 226 471 232 472
rect 226 467 227 471
rect 231 467 232 471
rect 226 466 232 467
rect 312 459 314 478
rect 372 472 374 494
rect 470 483 476 484
rect 470 479 471 483
rect 475 479 476 483
rect 470 478 476 479
rect 370 471 376 472
rect 370 467 371 471
rect 375 467 376 471
rect 370 466 376 467
rect 472 459 474 478
rect 532 472 534 494
rect 638 483 644 484
rect 638 479 639 483
rect 643 479 644 483
rect 638 478 644 479
rect 530 471 536 472
rect 530 467 531 471
rect 535 467 536 471
rect 530 466 536 467
rect 640 459 642 478
rect 700 472 702 494
rect 806 483 812 484
rect 806 479 807 483
rect 811 479 812 483
rect 806 478 812 479
rect 698 471 704 472
rect 698 467 699 471
rect 703 467 704 471
rect 698 466 704 467
rect 808 459 810 478
rect 816 472 818 550
rect 926 545 932 546
rect 926 541 927 545
rect 931 541 932 545
rect 926 540 932 541
rect 928 535 930 540
rect 927 534 931 535
rect 927 529 931 530
rect 959 534 963 535
rect 959 529 963 530
rect 960 524 962 529
rect 958 523 964 524
rect 958 519 959 523
rect 963 519 964 523
rect 958 518 964 519
rect 1028 516 1030 590
rect 1064 586 1066 597
rect 1192 586 1194 597
rect 1328 586 1330 597
rect 1472 586 1474 597
rect 1616 586 1618 597
rect 1686 595 1692 596
rect 1686 591 1687 595
rect 1691 591 1692 595
rect 1686 590 1692 591
rect 1694 595 1700 596
rect 1694 591 1695 595
rect 1699 591 1700 595
rect 1694 590 1700 591
rect 1062 585 1068 586
rect 1062 581 1063 585
rect 1067 581 1068 585
rect 1062 580 1068 581
rect 1190 585 1196 586
rect 1190 581 1191 585
rect 1195 581 1196 585
rect 1190 580 1196 581
rect 1326 585 1332 586
rect 1326 581 1327 585
rect 1331 581 1332 585
rect 1326 580 1332 581
rect 1470 585 1476 586
rect 1470 581 1471 585
rect 1475 581 1476 585
rect 1470 580 1476 581
rect 1614 585 1620 586
rect 1614 581 1615 585
rect 1619 581 1620 585
rect 1614 580 1620 581
rect 1688 568 1690 590
rect 1686 567 1692 568
rect 1686 563 1687 567
rect 1691 563 1692 567
rect 1686 562 1692 563
rect 1538 555 1544 556
rect 1538 551 1539 555
rect 1543 551 1544 555
rect 1538 550 1544 551
rect 1054 545 1060 546
rect 1054 541 1055 545
rect 1059 541 1060 545
rect 1054 540 1060 541
rect 1182 545 1188 546
rect 1182 541 1183 545
rect 1187 541 1188 545
rect 1182 540 1188 541
rect 1318 545 1324 546
rect 1318 541 1319 545
rect 1323 541 1324 545
rect 1318 540 1324 541
rect 1462 545 1468 546
rect 1462 541 1463 545
rect 1467 541 1468 545
rect 1462 540 1468 541
rect 1056 535 1058 540
rect 1184 535 1186 540
rect 1320 535 1322 540
rect 1464 535 1466 540
rect 1055 534 1059 535
rect 1055 529 1059 530
rect 1103 534 1107 535
rect 1103 529 1107 530
rect 1183 534 1187 535
rect 1183 529 1187 530
rect 1239 534 1243 535
rect 1239 529 1243 530
rect 1319 534 1323 535
rect 1319 529 1323 530
rect 1367 534 1371 535
rect 1367 529 1371 530
rect 1463 534 1467 535
rect 1463 529 1467 530
rect 1495 534 1499 535
rect 1495 529 1499 530
rect 1104 524 1106 529
rect 1240 524 1242 529
rect 1368 524 1370 529
rect 1496 524 1498 529
rect 1102 523 1108 524
rect 1102 519 1103 523
rect 1107 519 1108 523
rect 1102 518 1108 519
rect 1238 523 1244 524
rect 1238 519 1239 523
rect 1243 519 1244 523
rect 1238 518 1244 519
rect 1366 523 1372 524
rect 1366 519 1367 523
rect 1371 519 1372 523
rect 1366 518 1372 519
rect 1494 523 1500 524
rect 1494 519 1495 523
rect 1499 519 1500 523
rect 1494 518 1500 519
rect 1026 515 1032 516
rect 1026 511 1027 515
rect 1031 511 1032 515
rect 1026 510 1032 511
rect 1026 499 1032 500
rect 1026 495 1027 499
rect 1031 495 1032 499
rect 1026 494 1032 495
rect 1454 499 1460 500
rect 1454 495 1455 499
rect 1459 495 1460 499
rect 1454 494 1460 495
rect 1462 499 1468 500
rect 1462 495 1463 499
rect 1467 495 1468 499
rect 1462 494 1468 495
rect 966 483 972 484
rect 966 479 967 483
rect 971 479 972 483
rect 966 478 972 479
rect 814 471 820 472
rect 814 467 815 471
rect 819 467 820 471
rect 814 466 820 467
rect 968 459 970 478
rect 1028 472 1030 494
rect 1110 483 1116 484
rect 1110 479 1111 483
rect 1115 479 1116 483
rect 1110 478 1116 479
rect 1246 483 1252 484
rect 1246 479 1247 483
rect 1251 479 1252 483
rect 1246 478 1252 479
rect 1374 483 1380 484
rect 1374 479 1375 483
rect 1379 479 1380 483
rect 1374 478 1380 479
rect 1026 471 1032 472
rect 1026 467 1027 471
rect 1031 467 1032 471
rect 1026 466 1032 467
rect 1112 459 1114 478
rect 1238 471 1244 472
rect 1238 467 1239 471
rect 1243 467 1244 471
rect 1238 466 1244 467
rect 167 458 171 459
rect 167 453 171 454
rect 271 458 275 459
rect 271 453 275 454
rect 311 458 315 459
rect 311 453 315 454
rect 439 458 443 459
rect 439 453 443 454
rect 471 458 475 459
rect 471 453 475 454
rect 615 458 619 459
rect 615 453 619 454
rect 639 458 643 459
rect 639 453 643 454
rect 791 458 795 459
rect 791 453 795 454
rect 807 458 811 459
rect 807 453 811 454
rect 967 458 971 459
rect 967 453 971 454
rect 1111 458 1115 459
rect 1111 453 1115 454
rect 1127 458 1131 459
rect 1127 453 1131 454
rect 150 451 156 452
rect 150 447 151 451
rect 155 447 156 451
rect 150 446 156 447
rect 272 442 274 453
rect 382 451 388 452
rect 382 447 383 451
rect 387 447 388 451
rect 382 446 388 447
rect 142 441 148 442
rect 142 437 143 441
rect 147 437 148 441
rect 142 436 148 437
rect 270 441 276 442
rect 270 437 271 441
rect 275 437 276 441
rect 270 436 276 437
rect 110 428 116 429
rect 384 428 386 446
rect 440 442 442 453
rect 616 442 618 453
rect 792 442 794 453
rect 968 442 970 453
rect 1128 442 1130 453
rect 438 441 444 442
rect 438 437 439 441
rect 443 437 444 441
rect 438 436 444 437
rect 614 441 620 442
rect 614 437 615 441
rect 619 437 620 441
rect 614 436 620 437
rect 790 441 796 442
rect 790 437 791 441
rect 795 437 796 441
rect 790 436 796 437
rect 966 441 972 442
rect 966 437 967 441
rect 971 437 972 441
rect 966 436 972 437
rect 1126 441 1132 442
rect 1126 437 1127 441
rect 1131 437 1132 441
rect 1240 437 1242 466
rect 1248 459 1250 478
rect 1376 459 1378 478
rect 1247 458 1251 459
rect 1247 453 1251 454
rect 1287 458 1291 459
rect 1287 453 1291 454
rect 1375 458 1379 459
rect 1375 453 1379 454
rect 1447 458 1451 459
rect 1447 453 1451 454
rect 1288 442 1290 453
rect 1448 442 1450 453
rect 1456 452 1458 494
rect 1464 464 1466 494
rect 1502 483 1508 484
rect 1502 479 1503 483
rect 1507 479 1508 483
rect 1502 478 1508 479
rect 1462 463 1468 464
rect 1462 459 1463 463
rect 1467 459 1468 463
rect 1504 459 1506 478
rect 1540 472 1542 550
rect 1606 545 1612 546
rect 1606 541 1607 545
rect 1611 541 1612 545
rect 1606 540 1612 541
rect 1608 535 1610 540
rect 1607 534 1611 535
rect 1607 529 1611 530
rect 1623 534 1627 535
rect 1623 529 1627 530
rect 1624 524 1626 529
rect 1622 523 1628 524
rect 1622 519 1623 523
rect 1627 519 1628 523
rect 1622 518 1628 519
rect 1696 516 1698 590
rect 1736 586 1738 597
rect 1734 585 1740 586
rect 1734 581 1735 585
rect 1739 581 1740 585
rect 1734 580 1740 581
rect 1824 573 1826 597
rect 1864 573 1866 597
rect 1896 586 1898 597
rect 1970 595 1976 596
rect 1970 591 1971 595
rect 1975 591 1976 595
rect 1970 590 1976 591
rect 1894 585 1900 586
rect 1894 581 1895 585
rect 1899 581 1900 585
rect 1894 580 1900 581
rect 1822 572 1828 573
rect 1822 568 1823 572
rect 1827 568 1828 572
rect 1822 567 1828 568
rect 1862 572 1868 573
rect 1862 568 1863 572
rect 1867 568 1868 572
rect 1972 568 1974 590
rect 2088 586 2090 597
rect 2100 596 2102 646
rect 2450 635 2456 636
rect 2450 631 2451 635
rect 2455 631 2456 635
rect 2450 630 2456 631
rect 2714 635 2720 636
rect 2714 631 2715 635
rect 2719 631 2720 635
rect 2714 630 2720 631
rect 2206 619 2212 620
rect 2206 615 2207 619
rect 2211 615 2212 619
rect 2206 614 2212 615
rect 2390 619 2396 620
rect 2390 615 2391 619
rect 2395 615 2396 619
rect 2390 614 2396 615
rect 2208 603 2210 614
rect 2392 603 2394 614
rect 2452 608 2454 630
rect 2574 619 2580 620
rect 2574 615 2575 619
rect 2579 615 2580 619
rect 2574 614 2580 615
rect 2450 607 2456 608
rect 2450 603 2451 607
rect 2455 603 2456 607
rect 2576 603 2578 614
rect 2207 602 2211 603
rect 2207 597 2211 598
rect 2303 602 2307 603
rect 2303 597 2307 598
rect 2391 602 2395 603
rect 2450 602 2456 603
rect 2511 602 2515 603
rect 2391 597 2395 598
rect 2511 597 2515 598
rect 2575 602 2579 603
rect 2575 597 2579 598
rect 2703 602 2707 603
rect 2703 597 2707 598
rect 2098 595 2104 596
rect 2098 591 2099 595
rect 2103 591 2104 595
rect 2098 590 2104 591
rect 2304 586 2306 597
rect 2512 586 2514 597
rect 2704 586 2706 597
rect 2716 596 2718 630
rect 2750 619 2756 620
rect 2750 615 2751 619
rect 2755 615 2756 619
rect 2750 614 2756 615
rect 2918 619 2924 620
rect 2918 615 2919 619
rect 2923 615 2924 619
rect 2918 614 2924 615
rect 3070 619 3076 620
rect 3070 615 3071 619
rect 3075 615 3076 619
rect 3070 614 3076 615
rect 2752 603 2754 614
rect 2763 612 2767 613
rect 2762 607 2768 608
rect 2762 603 2763 607
rect 2767 603 2768 607
rect 2920 603 2922 614
rect 2938 607 2944 608
rect 2938 603 2939 607
rect 2943 603 2944 607
rect 3072 603 3074 614
rect 3080 613 3082 690
rect 3126 685 3132 686
rect 3126 681 3127 685
rect 3131 681 3132 685
rect 3126 680 3132 681
rect 3128 671 3130 680
rect 3127 670 3131 671
rect 3127 665 3131 666
rect 3192 652 3194 730
rect 3288 726 3290 737
rect 3440 726 3442 737
rect 3450 735 3456 736
rect 3450 731 3451 735
rect 3455 731 3456 735
rect 3450 730 3456 731
rect 3286 725 3292 726
rect 3286 721 3287 725
rect 3291 721 3292 725
rect 3286 720 3292 721
rect 3438 725 3444 726
rect 3438 721 3439 725
rect 3443 721 3444 725
rect 3438 720 3444 721
rect 3226 695 3232 696
rect 3226 691 3227 695
rect 3231 691 3232 695
rect 3226 690 3232 691
rect 3207 670 3211 671
rect 3207 665 3211 666
rect 3208 660 3210 665
rect 3206 659 3212 660
rect 3206 655 3207 659
rect 3211 655 3212 659
rect 3206 654 3212 655
rect 3190 651 3196 652
rect 3190 647 3191 651
rect 3195 647 3196 651
rect 3190 646 3196 647
rect 3214 619 3220 620
rect 3214 615 3215 619
rect 3219 615 3220 619
rect 3214 614 3220 615
rect 3079 612 3083 613
rect 3079 607 3083 608
rect 3216 603 3218 614
rect 3228 608 3230 690
rect 3278 685 3284 686
rect 3278 681 3279 685
rect 3283 681 3284 685
rect 3278 680 3284 681
rect 3430 685 3436 686
rect 3430 681 3431 685
rect 3435 681 3436 685
rect 3430 680 3436 681
rect 3280 671 3282 680
rect 3432 671 3434 680
rect 3279 670 3283 671
rect 3279 665 3283 666
rect 3351 670 3355 671
rect 3351 665 3355 666
rect 3431 670 3435 671
rect 3431 665 3435 666
rect 3352 660 3354 665
rect 3350 659 3356 660
rect 3350 655 3351 659
rect 3355 655 3356 659
rect 3350 654 3356 655
rect 3342 651 3348 652
rect 3342 647 3343 651
rect 3347 647 3348 651
rect 3342 646 3348 647
rect 3226 607 3232 608
rect 3226 603 3227 607
rect 3231 603 3232 607
rect 2751 602 2755 603
rect 2762 602 2768 603
rect 2879 602 2883 603
rect 2751 597 2755 598
rect 2879 597 2883 598
rect 2919 602 2923 603
rect 2938 602 2944 603
rect 3039 602 3043 603
rect 2919 597 2923 598
rect 2714 595 2720 596
rect 2714 591 2715 595
rect 2719 591 2720 595
rect 2714 590 2720 591
rect 2880 586 2882 597
rect 2086 585 2092 586
rect 2086 581 2087 585
rect 2091 581 2092 585
rect 2086 580 2092 581
rect 2302 585 2308 586
rect 2302 581 2303 585
rect 2307 581 2308 585
rect 2302 580 2308 581
rect 2510 585 2516 586
rect 2510 581 2511 585
rect 2515 581 2516 585
rect 2510 580 2516 581
rect 2702 585 2708 586
rect 2702 581 2703 585
rect 2707 581 2708 585
rect 2702 580 2708 581
rect 2878 585 2884 586
rect 2878 581 2879 585
rect 2883 581 2884 585
rect 2878 580 2884 581
rect 2940 572 2942 602
rect 3039 597 3043 598
rect 3071 602 3075 603
rect 3071 597 3075 598
rect 3199 602 3203 603
rect 3199 597 3203 598
rect 3215 602 3219 603
rect 3226 602 3232 603
rect 3215 597 3219 598
rect 3266 599 3272 600
rect 3040 586 3042 597
rect 3200 586 3202 597
rect 3266 595 3267 599
rect 3271 595 3272 599
rect 3344 596 3346 646
rect 3358 619 3364 620
rect 3358 615 3359 619
rect 3363 615 3364 619
rect 3358 614 3364 615
rect 3360 603 3362 614
rect 3351 602 3355 603
rect 3351 597 3355 598
rect 3359 602 3363 603
rect 3359 597 3363 598
rect 3266 594 3272 595
rect 3342 595 3348 596
rect 3038 585 3044 586
rect 3038 581 3039 585
rect 3043 581 3044 585
rect 3038 580 3044 581
rect 3198 585 3204 586
rect 3198 581 3199 585
rect 3203 581 3204 585
rect 3198 580 3204 581
rect 2938 571 2944 572
rect 1862 567 1868 568
rect 1970 567 1976 568
rect 1970 563 1971 567
rect 1975 563 1976 567
rect 2938 567 2939 571
rect 2943 567 2944 571
rect 3268 568 3270 594
rect 3342 591 3343 595
rect 3347 591 3348 595
rect 3342 590 3348 591
rect 3352 586 3354 597
rect 3350 585 3356 586
rect 3350 581 3351 585
rect 3355 581 3356 585
rect 3350 580 3356 581
rect 2938 566 2944 567
rect 3266 567 3272 568
rect 1970 562 1976 563
rect 3266 563 3267 567
rect 3271 563 3272 567
rect 3266 562 3272 563
rect 1822 555 1828 556
rect 1822 551 1823 555
rect 1827 551 1828 555
rect 1822 550 1828 551
rect 1862 555 1868 556
rect 1862 551 1863 555
rect 1867 551 1868 555
rect 1862 550 1868 551
rect 1870 555 1876 556
rect 1870 551 1871 555
rect 1875 551 1876 555
rect 1870 550 1876 551
rect 3350 555 3356 556
rect 3350 551 3351 555
rect 3355 551 3356 555
rect 3350 550 3356 551
rect 1726 545 1732 546
rect 1726 541 1727 545
rect 1731 541 1732 545
rect 1726 540 1732 541
rect 1728 535 1730 540
rect 1824 535 1826 550
rect 1727 534 1731 535
rect 1727 529 1731 530
rect 1823 534 1827 535
rect 1823 529 1827 530
rect 1728 524 1730 529
rect 1726 523 1732 524
rect 1726 519 1727 523
rect 1731 519 1732 523
rect 1726 518 1732 519
rect 1694 515 1700 516
rect 1694 511 1695 515
rect 1699 511 1700 515
rect 1824 514 1826 529
rect 1864 527 1866 550
rect 1863 526 1867 527
rect 1863 521 1867 522
rect 1694 510 1700 511
rect 1822 513 1828 514
rect 1822 509 1823 513
rect 1827 509 1828 513
rect 1822 508 1828 509
rect 1864 506 1866 521
rect 1862 505 1868 506
rect 1862 501 1863 505
rect 1867 501 1868 505
rect 1862 500 1868 501
rect 1822 496 1828 497
rect 1822 492 1823 496
rect 1827 492 1828 496
rect 1822 491 1828 492
rect 1630 483 1636 484
rect 1630 479 1631 483
rect 1635 479 1636 483
rect 1630 478 1636 479
rect 1734 483 1740 484
rect 1734 479 1735 483
rect 1739 479 1740 483
rect 1734 478 1740 479
rect 1538 471 1544 472
rect 1538 467 1539 471
rect 1543 467 1544 471
rect 1538 466 1544 467
rect 1632 459 1634 478
rect 1736 459 1738 478
rect 1824 459 1826 491
rect 1862 488 1868 489
rect 1862 484 1863 488
rect 1867 484 1868 488
rect 1862 483 1868 484
rect 1864 459 1866 483
rect 1872 472 1874 550
rect 1886 545 1892 546
rect 1886 541 1887 545
rect 1891 541 1892 545
rect 1886 540 1892 541
rect 2078 545 2084 546
rect 2078 541 2079 545
rect 2083 541 2084 545
rect 2078 540 2084 541
rect 2294 545 2300 546
rect 2294 541 2295 545
rect 2299 541 2300 545
rect 2294 540 2300 541
rect 2502 545 2508 546
rect 2502 541 2503 545
rect 2507 541 2508 545
rect 2502 540 2508 541
rect 2694 545 2700 546
rect 2694 541 2695 545
rect 2699 541 2700 545
rect 2694 540 2700 541
rect 2870 545 2876 546
rect 2870 541 2871 545
rect 2875 541 2876 545
rect 2870 540 2876 541
rect 3030 545 3036 546
rect 3030 541 3031 545
rect 3035 541 3036 545
rect 3030 540 3036 541
rect 3190 545 3196 546
rect 3190 541 3191 545
rect 3195 541 3196 545
rect 3190 540 3196 541
rect 3342 545 3348 546
rect 3342 541 3343 545
rect 3347 541 3348 545
rect 3342 540 3348 541
rect 1888 527 1890 540
rect 2080 527 2082 540
rect 2296 527 2298 540
rect 2504 527 2506 540
rect 2696 527 2698 540
rect 2872 527 2874 540
rect 3032 527 3034 540
rect 3192 527 3194 540
rect 3344 527 3346 540
rect 1887 526 1891 527
rect 1887 521 1891 522
rect 2079 526 2083 527
rect 2079 521 2083 522
rect 2287 526 2291 527
rect 2287 521 2291 522
rect 2295 526 2299 527
rect 2295 521 2299 522
rect 2487 526 2491 527
rect 2487 521 2491 522
rect 2503 526 2507 527
rect 2503 521 2507 522
rect 2671 526 2675 527
rect 2671 521 2675 522
rect 2695 526 2699 527
rect 2695 521 2699 522
rect 2847 526 2851 527
rect 2847 521 2851 522
rect 2871 526 2875 527
rect 2871 521 2875 522
rect 3015 526 3019 527
rect 3015 521 3019 522
rect 3031 526 3035 527
rect 3031 521 3035 522
rect 3175 526 3179 527
rect 3175 521 3179 522
rect 3191 526 3195 527
rect 3191 521 3195 522
rect 3335 526 3339 527
rect 3335 521 3339 522
rect 3343 526 3347 527
rect 3343 521 3347 522
rect 2080 516 2082 521
rect 2288 516 2290 521
rect 2488 516 2490 521
rect 2672 516 2674 521
rect 2848 516 2850 521
rect 3016 516 3018 521
rect 3176 516 3178 521
rect 3336 516 3338 521
rect 2078 515 2084 516
rect 2078 511 2079 515
rect 2083 511 2084 515
rect 2078 510 2084 511
rect 2286 515 2292 516
rect 2286 511 2287 515
rect 2291 511 2292 515
rect 2286 510 2292 511
rect 2486 515 2492 516
rect 2486 511 2487 515
rect 2491 511 2492 515
rect 2486 510 2492 511
rect 2670 515 2676 516
rect 2670 511 2671 515
rect 2675 511 2676 515
rect 2670 510 2676 511
rect 2846 515 2852 516
rect 2846 511 2847 515
rect 2851 511 2852 515
rect 2846 510 2852 511
rect 3014 515 3020 516
rect 3014 511 3015 515
rect 3019 511 3020 515
rect 3014 510 3020 511
rect 3174 515 3180 516
rect 3174 511 3175 515
rect 3179 511 3180 515
rect 3174 510 3180 511
rect 3334 515 3340 516
rect 3334 511 3335 515
rect 3339 511 3340 515
rect 3334 510 3340 511
rect 3082 507 3088 508
rect 3082 503 3083 507
rect 3087 503 3088 507
rect 3082 502 3088 503
rect 2418 491 2424 492
rect 2418 487 2419 491
rect 2423 487 2424 491
rect 2418 486 2424 487
rect 2086 475 2092 476
rect 1870 471 1876 472
rect 1870 467 1871 471
rect 1875 467 1876 471
rect 2086 471 2087 475
rect 2091 471 2092 475
rect 2086 470 2092 471
rect 2294 475 2300 476
rect 2294 471 2295 475
rect 2299 471 2300 475
rect 2294 470 2300 471
rect 1870 466 1876 467
rect 2088 459 2090 470
rect 2095 468 2099 469
rect 2094 463 2100 464
rect 2094 459 2095 463
rect 2099 459 2100 463
rect 2296 459 2298 470
rect 2420 469 2422 486
rect 2494 475 2500 476
rect 2494 471 2495 475
rect 2499 471 2500 475
rect 2494 470 2500 471
rect 2678 475 2684 476
rect 2678 471 2679 475
rect 2683 471 2684 475
rect 2678 470 2684 471
rect 2854 475 2860 476
rect 2854 471 2855 475
rect 2859 471 2860 475
rect 2854 470 2860 471
rect 3022 475 3028 476
rect 3022 471 3023 475
rect 3027 471 3028 475
rect 3022 470 3028 471
rect 2419 468 2423 469
rect 2419 463 2423 464
rect 2496 459 2498 470
rect 2506 463 2512 464
rect 2506 459 2507 463
rect 2511 459 2512 463
rect 2680 459 2682 470
rect 2687 468 2691 469
rect 2686 463 2692 464
rect 2686 459 2687 463
rect 2691 459 2692 463
rect 2856 459 2858 470
rect 3024 459 3026 470
rect 3084 469 3086 502
rect 3242 491 3248 492
rect 3242 487 3243 491
rect 3247 487 3248 491
rect 3242 486 3248 487
rect 3182 475 3188 476
rect 3182 471 3183 475
rect 3187 471 3188 475
rect 3182 470 3188 471
rect 3083 468 3087 469
rect 3083 463 3087 464
rect 3184 459 3186 470
rect 3244 464 3246 486
rect 3342 475 3348 476
rect 3342 471 3343 475
rect 3347 471 3348 475
rect 3342 470 3348 471
rect 3242 463 3248 464
rect 3242 459 3243 463
rect 3247 459 3248 463
rect 3344 459 3346 470
rect 3352 464 3354 550
rect 3452 508 3454 730
rect 3472 608 3474 774
rect 3486 763 3492 764
rect 3486 759 3487 763
rect 3491 759 3492 763
rect 3486 758 3492 759
rect 3488 743 3490 758
rect 3500 752 3502 814
rect 3498 751 3504 752
rect 3498 747 3499 751
rect 3503 747 3504 751
rect 3498 746 3504 747
rect 3487 742 3491 743
rect 3487 737 3491 738
rect 3508 712 3510 870
rect 3576 853 3578 877
rect 3574 852 3580 853
rect 3574 848 3575 852
rect 3579 848 3580 852
rect 3574 847 3580 848
rect 3574 835 3580 836
rect 3574 831 3575 835
rect 3579 831 3580 835
rect 3574 830 3580 831
rect 3576 815 3578 830
rect 3575 814 3579 815
rect 3575 809 3579 810
rect 3576 794 3578 809
rect 3574 793 3580 794
rect 3574 789 3575 793
rect 3579 789 3580 793
rect 3574 788 3580 789
rect 3574 776 3580 777
rect 3574 772 3575 776
rect 3579 772 3580 776
rect 3574 771 3580 772
rect 3576 743 3578 771
rect 3575 742 3579 743
rect 3575 737 3579 738
rect 3576 713 3578 737
rect 3574 712 3580 713
rect 3506 711 3512 712
rect 3506 707 3507 711
rect 3511 707 3512 711
rect 3574 708 3575 712
rect 3579 708 3580 712
rect 3574 707 3580 708
rect 3506 706 3512 707
rect 3574 695 3580 696
rect 3574 691 3575 695
rect 3579 691 3580 695
rect 3574 690 3580 691
rect 3576 671 3578 690
rect 3479 670 3483 671
rect 3479 665 3483 666
rect 3575 670 3579 671
rect 3575 665 3579 666
rect 3480 660 3482 665
rect 3478 659 3484 660
rect 3478 655 3479 659
rect 3483 655 3484 659
rect 3478 654 3484 655
rect 3576 650 3578 665
rect 3574 649 3580 650
rect 3574 645 3575 649
rect 3579 645 3580 649
rect 3574 644 3580 645
rect 3574 632 3580 633
rect 3574 628 3575 632
rect 3579 628 3580 632
rect 3574 627 3580 628
rect 3486 619 3492 620
rect 3486 615 3487 619
rect 3491 615 3492 619
rect 3486 614 3492 615
rect 3470 607 3476 608
rect 3470 603 3471 607
rect 3475 603 3476 607
rect 3488 603 3490 614
rect 3576 603 3578 627
rect 3470 602 3476 603
rect 3487 602 3491 603
rect 3487 597 3491 598
rect 3575 602 3579 603
rect 3575 597 3579 598
rect 3488 586 3490 597
rect 3486 585 3492 586
rect 3486 581 3487 585
rect 3491 581 3492 585
rect 3486 580 3492 581
rect 3576 573 3578 597
rect 3574 572 3580 573
rect 3574 568 3575 572
rect 3579 568 3580 572
rect 3574 567 3580 568
rect 3574 555 3580 556
rect 3574 551 3575 555
rect 3579 551 3580 555
rect 3574 550 3580 551
rect 3478 545 3484 546
rect 3478 541 3479 545
rect 3483 541 3484 545
rect 3478 540 3484 541
rect 3480 527 3482 540
rect 3576 527 3578 550
rect 3479 526 3483 527
rect 3479 521 3483 522
rect 3575 526 3579 527
rect 3575 521 3579 522
rect 3480 516 3482 521
rect 3478 515 3484 516
rect 3478 511 3479 515
rect 3483 511 3484 515
rect 3478 510 3484 511
rect 3450 507 3456 508
rect 3450 503 3451 507
rect 3455 503 3456 507
rect 3576 506 3578 521
rect 3450 502 3456 503
rect 3574 505 3580 506
rect 3574 501 3575 505
rect 3579 501 3580 505
rect 3574 500 3580 501
rect 3574 488 3580 489
rect 3574 484 3575 488
rect 3579 484 3580 488
rect 3574 483 3580 484
rect 3486 475 3492 476
rect 3486 471 3487 475
rect 3491 471 3492 475
rect 3486 470 3492 471
rect 3350 463 3356 464
rect 3350 459 3351 463
rect 3355 459 3356 463
rect 1462 458 1468 459
rect 1503 458 1507 459
rect 1503 453 1507 454
rect 1607 458 1611 459
rect 1607 453 1611 454
rect 1631 458 1635 459
rect 1631 453 1635 454
rect 1735 458 1739 459
rect 1735 453 1739 454
rect 1823 458 1827 459
rect 1823 453 1827 454
rect 1863 458 1867 459
rect 1863 453 1867 454
rect 2087 458 2091 459
rect 2094 458 2100 459
rect 2247 458 2251 459
rect 2087 453 2091 454
rect 2247 453 2251 454
rect 2295 458 2299 459
rect 2295 453 2299 454
rect 2335 458 2339 459
rect 2335 453 2339 454
rect 2431 458 2435 459
rect 2431 453 2435 454
rect 2495 458 2499 459
rect 2506 458 2512 459
rect 2527 458 2531 459
rect 2495 453 2499 454
rect 1454 451 1460 452
rect 1454 447 1455 451
rect 1459 447 1460 451
rect 1454 446 1460 447
rect 1608 442 1610 453
rect 1286 441 1292 442
rect 1286 437 1287 441
rect 1291 437 1292 441
rect 1126 436 1132 437
rect 1239 436 1243 437
rect 1286 436 1292 437
rect 1446 441 1452 442
rect 1446 437 1447 441
rect 1451 437 1452 441
rect 1606 441 1612 442
rect 1606 437 1607 441
rect 1611 437 1612 441
rect 1446 436 1452 437
rect 1547 436 1551 437
rect 1606 436 1612 437
rect 1239 431 1243 432
rect 1547 431 1551 432
rect 110 424 111 428
rect 115 424 116 428
rect 110 423 116 424
rect 382 427 388 428
rect 382 423 383 427
rect 387 423 388 427
rect 1548 424 1550 431
rect 1824 429 1826 453
rect 1864 429 1866 453
rect 2248 442 2250 453
rect 2302 447 2308 448
rect 2302 442 2303 447
rect 2246 441 2252 442
rect 2246 437 2247 441
rect 2251 437 2252 441
rect 2307 442 2308 447
rect 2336 442 2338 453
rect 2432 442 2434 453
rect 2303 439 2307 440
rect 2334 441 2340 442
rect 2246 436 2252 437
rect 2334 437 2335 441
rect 2339 437 2340 441
rect 2334 436 2340 437
rect 2430 441 2436 442
rect 2430 437 2431 441
rect 2435 437 2436 441
rect 2430 436 2436 437
rect 1822 428 1828 429
rect 1822 424 1823 428
rect 1827 424 1828 428
rect 382 422 388 423
rect 1546 423 1552 424
rect 1822 423 1828 424
rect 1862 428 1868 429
rect 1862 424 1863 428
rect 1867 424 1868 428
rect 2508 424 2510 458
rect 2527 453 2531 454
rect 2623 458 2627 459
rect 2623 453 2627 454
rect 2679 458 2683 459
rect 2686 458 2692 459
rect 2735 458 2739 459
rect 2679 453 2683 454
rect 2735 453 2739 454
rect 2855 458 2859 459
rect 2855 453 2859 454
rect 2863 458 2867 459
rect 2863 453 2867 454
rect 3007 458 3011 459
rect 3007 453 3011 454
rect 3023 458 3027 459
rect 3023 453 3027 454
rect 3167 458 3171 459
rect 3167 453 3171 454
rect 3183 458 3187 459
rect 3242 458 3248 459
rect 3335 458 3339 459
rect 3183 453 3187 454
rect 3335 453 3339 454
rect 3343 458 3347 459
rect 3350 458 3356 459
rect 3478 463 3484 464
rect 3478 459 3479 463
rect 3483 459 3484 463
rect 3488 459 3490 470
rect 3576 459 3578 483
rect 3478 458 3484 459
rect 3487 458 3491 459
rect 3343 453 3347 454
rect 2528 442 2530 453
rect 2578 451 2584 452
rect 2578 447 2579 451
rect 2583 447 2584 451
rect 2578 446 2584 447
rect 2526 441 2532 442
rect 2526 437 2527 441
rect 2531 437 2532 441
rect 2526 436 2532 437
rect 1862 423 1868 424
rect 2506 423 2512 424
rect 1546 419 1547 423
rect 1551 419 1552 423
rect 1546 418 1552 419
rect 2506 419 2507 423
rect 2511 419 2512 423
rect 2506 418 2512 419
rect 110 411 116 412
rect 110 407 111 411
rect 115 407 116 411
rect 110 406 116 407
rect 682 411 688 412
rect 682 407 683 411
rect 687 407 688 411
rect 682 406 688 407
rect 1286 411 1292 412
rect 1286 407 1287 411
rect 1291 407 1292 411
rect 1286 406 1292 407
rect 1822 411 1828 412
rect 1822 407 1823 411
rect 1827 407 1828 411
rect 1822 406 1828 407
rect 1862 411 1868 412
rect 1862 407 1863 411
rect 1867 407 1868 411
rect 1862 406 1868 407
rect 112 391 114 406
rect 134 401 140 402
rect 134 397 135 401
rect 139 397 140 401
rect 134 396 140 397
rect 262 401 268 402
rect 262 397 263 401
rect 267 397 268 401
rect 262 396 268 397
rect 430 401 436 402
rect 430 397 431 401
rect 435 397 436 401
rect 430 396 436 397
rect 606 401 612 402
rect 606 397 607 401
rect 611 397 612 401
rect 606 396 612 397
rect 136 391 138 396
rect 264 391 266 396
rect 432 391 434 396
rect 608 391 610 396
rect 111 390 115 391
rect 111 385 115 386
rect 135 390 139 391
rect 135 385 139 386
rect 263 390 267 391
rect 263 385 267 386
rect 431 390 435 391
rect 431 385 435 386
rect 607 390 611 391
rect 607 385 611 386
rect 112 370 114 385
rect 136 380 138 385
rect 264 380 266 385
rect 432 380 434 385
rect 608 380 610 385
rect 134 379 140 380
rect 134 375 135 379
rect 139 375 140 379
rect 134 374 140 375
rect 262 379 268 380
rect 262 375 263 379
rect 267 375 268 379
rect 262 374 268 375
rect 430 379 436 380
rect 430 375 431 379
rect 435 375 436 379
rect 430 374 436 375
rect 606 379 612 380
rect 606 375 607 379
rect 611 375 612 379
rect 606 374 612 375
rect 684 373 686 406
rect 782 401 788 402
rect 782 397 783 401
rect 787 397 788 401
rect 782 396 788 397
rect 958 401 964 402
rect 958 397 959 401
rect 963 397 964 401
rect 958 396 964 397
rect 1118 401 1124 402
rect 1118 397 1119 401
rect 1123 397 1124 401
rect 1118 396 1124 397
rect 1278 401 1284 402
rect 1278 397 1279 401
rect 1283 397 1284 401
rect 1278 396 1284 397
rect 784 391 786 396
rect 960 391 962 396
rect 1120 391 1122 396
rect 1280 391 1282 396
rect 783 390 787 391
rect 783 385 787 386
rect 951 390 955 391
rect 951 385 955 386
rect 959 390 963 391
rect 959 385 963 386
rect 1111 390 1115 391
rect 1111 385 1115 386
rect 1119 390 1123 391
rect 1119 385 1123 386
rect 1271 390 1275 391
rect 1271 385 1275 386
rect 1279 390 1283 391
rect 1279 385 1283 386
rect 784 380 786 385
rect 952 380 954 385
rect 1112 380 1114 385
rect 1272 380 1274 385
rect 782 379 788 380
rect 782 375 783 379
rect 787 375 788 379
rect 782 374 788 375
rect 950 379 956 380
rect 950 375 951 379
rect 955 375 956 379
rect 950 374 956 375
rect 1110 379 1116 380
rect 1110 375 1111 379
rect 1115 375 1116 379
rect 1110 374 1116 375
rect 1270 379 1276 380
rect 1270 375 1271 379
rect 1275 375 1276 379
rect 1270 374 1276 375
rect 155 372 159 373
rect 110 369 116 370
rect 110 365 111 369
rect 115 365 116 369
rect 155 367 159 368
rect 683 372 687 373
rect 683 367 687 368
rect 690 371 696 372
rect 690 367 691 371
rect 695 367 696 371
rect 110 364 116 365
rect 110 352 116 353
rect 110 348 111 352
rect 115 348 116 352
rect 110 347 116 348
rect 112 319 114 347
rect 142 339 148 340
rect 142 335 143 339
rect 147 335 148 339
rect 142 334 148 335
rect 144 319 146 334
rect 156 328 158 367
rect 690 366 696 367
rect 270 339 276 340
rect 270 335 271 339
rect 275 335 276 339
rect 270 334 276 335
rect 438 339 444 340
rect 438 335 439 339
rect 443 335 444 339
rect 438 334 444 335
rect 614 339 620 340
rect 614 335 615 339
rect 619 335 620 339
rect 614 334 620 335
rect 154 327 160 328
rect 154 323 155 327
rect 159 323 160 327
rect 154 322 160 323
rect 272 319 274 334
rect 351 332 355 333
rect 351 327 355 328
rect 111 318 115 319
rect 111 313 115 314
rect 143 318 147 319
rect 143 313 147 314
rect 263 318 267 319
rect 263 313 267 314
rect 271 318 275 319
rect 352 316 354 327
rect 440 319 442 334
rect 616 319 618 334
rect 692 333 694 366
rect 1018 355 1024 356
rect 1018 351 1019 355
rect 1023 351 1024 355
rect 1018 350 1024 351
rect 790 339 796 340
rect 790 335 791 339
rect 795 335 796 339
rect 790 334 796 335
rect 958 339 964 340
rect 958 335 959 339
rect 963 335 964 339
rect 958 334 964 335
rect 691 332 695 333
rect 691 327 695 328
rect 792 319 794 334
rect 960 319 962 334
rect 1020 328 1022 350
rect 1118 339 1124 340
rect 1118 335 1119 339
rect 1123 335 1124 339
rect 1118 334 1124 335
rect 1278 339 1284 340
rect 1278 335 1279 339
rect 1283 335 1284 339
rect 1278 334 1284 335
rect 1018 327 1024 328
rect 1018 323 1019 327
rect 1023 323 1024 327
rect 1018 322 1024 323
rect 1120 319 1122 334
rect 1242 327 1248 328
rect 1242 323 1243 327
rect 1247 323 1248 327
rect 1242 322 1248 323
rect 391 318 395 319
rect 271 313 275 314
rect 350 315 356 316
rect 112 289 114 313
rect 264 302 266 313
rect 350 311 351 315
rect 355 311 356 315
rect 391 313 395 314
rect 439 318 443 319
rect 439 313 443 314
rect 527 318 531 319
rect 527 313 531 314
rect 615 318 619 319
rect 615 313 619 314
rect 679 318 683 319
rect 679 313 683 314
rect 791 318 795 319
rect 791 313 795 314
rect 839 318 843 319
rect 839 313 843 314
rect 959 318 963 319
rect 959 313 963 314
rect 1007 318 1011 319
rect 1007 313 1011 314
rect 1119 318 1123 319
rect 1119 313 1123 314
rect 1175 318 1179 319
rect 1175 313 1179 314
rect 350 310 356 311
rect 358 311 364 312
rect 358 307 359 311
rect 363 307 364 311
rect 358 306 364 307
rect 262 301 268 302
rect 262 297 263 301
rect 267 297 268 301
rect 262 296 268 297
rect 110 288 116 289
rect 360 288 362 306
rect 392 302 394 313
rect 528 302 530 313
rect 680 302 682 313
rect 840 302 842 313
rect 1008 302 1010 313
rect 1176 302 1178 313
rect 1234 311 1240 312
rect 1234 307 1235 311
rect 1239 307 1240 311
rect 1234 306 1240 307
rect 390 301 396 302
rect 390 297 391 301
rect 395 297 396 301
rect 390 296 396 297
rect 526 301 532 302
rect 526 297 527 301
rect 531 297 532 301
rect 526 296 532 297
rect 678 301 684 302
rect 678 297 679 301
rect 683 297 684 301
rect 678 296 684 297
rect 838 301 844 302
rect 838 297 839 301
rect 843 297 844 301
rect 838 296 844 297
rect 1006 301 1012 302
rect 1006 297 1007 301
rect 1011 297 1012 301
rect 1006 296 1012 297
rect 1174 301 1180 302
rect 1174 297 1175 301
rect 1179 297 1180 301
rect 1174 296 1180 297
rect 1236 288 1238 306
rect 110 284 111 288
rect 115 284 116 288
rect 110 283 116 284
rect 358 287 364 288
rect 358 283 359 287
rect 363 283 364 287
rect 358 282 364 283
rect 1234 287 1240 288
rect 1234 283 1235 287
rect 1239 283 1240 287
rect 1244 284 1246 322
rect 1280 319 1282 334
rect 1288 328 1290 406
rect 1438 401 1444 402
rect 1438 397 1439 401
rect 1443 397 1444 401
rect 1438 396 1444 397
rect 1598 401 1604 402
rect 1598 397 1599 401
rect 1603 397 1604 401
rect 1598 396 1604 397
rect 1440 391 1442 396
rect 1600 391 1602 396
rect 1824 391 1826 406
rect 1864 391 1866 406
rect 2238 401 2244 402
rect 2238 397 2239 401
rect 2243 397 2244 401
rect 2238 396 2244 397
rect 2326 401 2332 402
rect 2326 397 2327 401
rect 2331 397 2332 401
rect 2326 396 2332 397
rect 2422 401 2428 402
rect 2422 397 2423 401
rect 2427 397 2428 401
rect 2422 396 2428 397
rect 2518 401 2524 402
rect 2518 397 2519 401
rect 2523 397 2524 401
rect 2518 396 2524 397
rect 2240 391 2242 396
rect 2328 391 2330 396
rect 2424 391 2426 396
rect 2520 391 2522 396
rect 1431 390 1435 391
rect 1431 385 1435 386
rect 1439 390 1443 391
rect 1439 385 1443 386
rect 1591 390 1595 391
rect 1591 385 1595 386
rect 1599 390 1603 391
rect 1599 385 1603 386
rect 1823 390 1827 391
rect 1823 385 1827 386
rect 1863 390 1867 391
rect 1863 385 1867 386
rect 2151 390 2155 391
rect 2151 385 2155 386
rect 2239 390 2243 391
rect 2239 385 2243 386
rect 2327 390 2331 391
rect 2327 385 2331 386
rect 2415 390 2419 391
rect 2415 385 2419 386
rect 2423 390 2427 391
rect 2423 385 2427 386
rect 2503 390 2507 391
rect 2503 385 2507 386
rect 2519 390 2523 391
rect 2519 385 2523 386
rect 1432 380 1434 385
rect 1592 380 1594 385
rect 1430 379 1436 380
rect 1430 375 1431 379
rect 1435 375 1436 379
rect 1430 374 1436 375
rect 1590 379 1596 380
rect 1590 375 1591 379
rect 1595 375 1596 379
rect 1590 374 1596 375
rect 1824 370 1826 385
rect 1864 370 1866 385
rect 2152 380 2154 385
rect 2240 380 2242 385
rect 2328 380 2330 385
rect 2416 380 2418 385
rect 2504 380 2506 385
rect 2150 379 2156 380
rect 2150 375 2151 379
rect 2155 375 2156 379
rect 2150 374 2156 375
rect 2238 379 2244 380
rect 2238 375 2239 379
rect 2243 375 2244 379
rect 2238 374 2244 375
rect 2326 379 2332 380
rect 2326 375 2327 379
rect 2331 375 2332 379
rect 2326 374 2332 375
rect 2414 379 2420 380
rect 2414 375 2415 379
rect 2419 375 2420 379
rect 2414 374 2420 375
rect 2502 379 2508 380
rect 2502 375 2503 379
rect 2507 375 2508 379
rect 2502 374 2508 375
rect 2580 372 2582 446
rect 2595 444 2599 445
rect 2624 442 2626 453
rect 2736 442 2738 453
rect 2790 451 2796 452
rect 2790 447 2791 451
rect 2795 447 2796 451
rect 2790 446 2796 447
rect 2595 439 2599 440
rect 2622 441 2628 442
rect 2596 424 2598 439
rect 2622 437 2623 441
rect 2627 437 2628 441
rect 2622 436 2628 437
rect 2734 441 2740 442
rect 2734 437 2735 441
rect 2739 437 2740 441
rect 2734 436 2740 437
rect 2594 423 2600 424
rect 2594 419 2595 423
rect 2599 419 2600 423
rect 2594 418 2600 419
rect 2614 401 2620 402
rect 2614 397 2615 401
rect 2619 397 2620 401
rect 2614 396 2620 397
rect 2726 401 2732 402
rect 2726 397 2727 401
rect 2731 397 2732 401
rect 2726 396 2732 397
rect 2792 396 2794 446
rect 2864 442 2866 453
rect 3008 442 3010 453
rect 3168 442 3170 453
rect 3336 442 3338 453
rect 2862 441 2868 442
rect 2862 437 2863 441
rect 2867 437 2868 441
rect 2862 436 2868 437
rect 3006 441 3012 442
rect 3006 437 3007 441
rect 3011 437 3012 441
rect 3006 436 3012 437
rect 3166 441 3172 442
rect 3166 437 3167 441
rect 3171 437 3172 441
rect 3166 436 3172 437
rect 3334 441 3340 442
rect 3334 437 3335 441
rect 3339 437 3340 441
rect 3334 436 3340 437
rect 3480 424 3482 458
rect 3487 453 3491 454
rect 3575 458 3579 459
rect 3575 453 3579 454
rect 3488 442 3490 453
rect 3486 441 3492 442
rect 3486 437 3487 441
rect 3491 437 3492 441
rect 3486 436 3492 437
rect 3576 429 3578 453
rect 3574 428 3580 429
rect 3574 424 3575 428
rect 3579 424 3580 428
rect 3478 423 3484 424
rect 3574 423 3580 424
rect 3478 419 3479 423
rect 3483 419 3484 423
rect 3478 418 3484 419
rect 2934 411 2940 412
rect 2934 407 2935 411
rect 2939 407 2940 411
rect 2934 406 2940 407
rect 3574 411 3580 412
rect 3574 407 3575 411
rect 3579 407 3580 411
rect 3574 406 3580 407
rect 2854 401 2860 402
rect 2854 397 2855 401
rect 2859 397 2860 401
rect 2854 396 2860 397
rect 2616 391 2618 396
rect 2728 391 2730 396
rect 2790 395 2796 396
rect 2790 391 2791 395
rect 2795 391 2796 395
rect 2856 391 2858 396
rect 2615 390 2619 391
rect 2615 385 2619 386
rect 2727 390 2731 391
rect 2727 385 2731 386
rect 2751 390 2755 391
rect 2790 390 2796 391
rect 2855 390 2859 391
rect 2751 385 2755 386
rect 2855 385 2859 386
rect 2919 390 2923 391
rect 2919 385 2923 386
rect 2616 380 2618 385
rect 2752 380 2754 385
rect 2920 380 2922 385
rect 2614 379 2620 380
rect 2614 375 2615 379
rect 2619 375 2620 379
rect 2614 374 2620 375
rect 2750 379 2756 380
rect 2750 375 2751 379
rect 2755 375 2756 379
rect 2750 374 2756 375
rect 2918 379 2924 380
rect 2918 375 2919 379
rect 2923 375 2924 379
rect 2918 374 2924 375
rect 2578 371 2584 372
rect 1822 369 1828 370
rect 1822 365 1823 369
rect 1827 365 1828 369
rect 1822 364 1828 365
rect 1862 369 1868 370
rect 1862 365 1863 369
rect 1867 365 1868 369
rect 2578 367 2579 371
rect 2583 367 2584 371
rect 2578 366 2584 367
rect 1862 364 1868 365
rect 1694 355 1700 356
rect 1694 351 1695 355
rect 1699 351 1700 355
rect 2570 355 2576 356
rect 1694 350 1700 351
rect 1822 352 1828 353
rect 1438 339 1444 340
rect 1438 335 1439 339
rect 1443 335 1444 339
rect 1438 334 1444 335
rect 1598 339 1604 340
rect 1598 335 1599 339
rect 1603 335 1604 339
rect 1598 334 1604 335
rect 1286 327 1292 328
rect 1286 323 1287 327
rect 1291 323 1292 327
rect 1286 322 1292 323
rect 1440 319 1442 334
rect 1600 319 1602 334
rect 1279 318 1283 319
rect 1279 313 1283 314
rect 1343 318 1347 319
rect 1343 313 1347 314
rect 1439 318 1443 319
rect 1439 313 1443 314
rect 1511 318 1515 319
rect 1511 313 1515 314
rect 1599 318 1603 319
rect 1599 313 1603 314
rect 1687 318 1691 319
rect 1687 313 1691 314
rect 1344 302 1346 313
rect 1512 302 1514 313
rect 1688 302 1690 313
rect 1696 312 1698 350
rect 1822 348 1823 352
rect 1827 348 1828 352
rect 1822 347 1828 348
rect 1862 352 1868 353
rect 1862 348 1863 352
rect 1867 348 1868 352
rect 2570 351 2571 355
rect 2575 351 2576 355
rect 2570 350 2576 351
rect 2682 355 2688 356
rect 2682 351 2683 355
rect 2687 351 2688 355
rect 2682 350 2688 351
rect 1862 347 1868 348
rect 1824 319 1826 347
rect 1864 323 1866 347
rect 2158 339 2164 340
rect 2158 335 2159 339
rect 2163 335 2164 339
rect 2158 334 2164 335
rect 2246 339 2252 340
rect 2246 335 2247 339
rect 2251 335 2252 339
rect 2246 334 2252 335
rect 2334 339 2340 340
rect 2334 335 2335 339
rect 2339 335 2340 339
rect 2334 334 2340 335
rect 2422 339 2428 340
rect 2422 335 2423 339
rect 2427 335 2428 339
rect 2422 334 2428 335
rect 2510 339 2516 340
rect 2510 335 2511 339
rect 2515 335 2516 339
rect 2510 334 2516 335
rect 2160 323 2162 334
rect 2214 327 2220 328
rect 2214 323 2215 327
rect 2219 323 2220 327
rect 2248 323 2250 334
rect 2336 323 2338 334
rect 2424 323 2426 334
rect 2512 323 2514 334
rect 1863 322 1867 323
rect 1823 318 1827 319
rect 1863 317 1867 318
rect 2023 322 2027 323
rect 2023 317 2027 318
rect 2119 322 2123 323
rect 2119 317 2123 318
rect 2159 322 2163 323
rect 2214 322 2220 323
rect 2223 322 2227 323
rect 2159 317 2163 318
rect 1823 313 1827 314
rect 1694 311 1700 312
rect 1694 307 1695 311
rect 1699 307 1700 311
rect 1694 306 1700 307
rect 1342 301 1348 302
rect 1342 297 1343 301
rect 1347 297 1348 301
rect 1342 296 1348 297
rect 1510 301 1516 302
rect 1510 297 1511 301
rect 1515 297 1516 301
rect 1510 296 1516 297
rect 1686 301 1692 302
rect 1686 297 1687 301
rect 1691 297 1692 301
rect 1686 296 1692 297
rect 1824 289 1826 313
rect 1864 293 1866 317
rect 2024 306 2026 317
rect 2030 315 2036 316
rect 2030 311 2031 315
rect 2035 311 2036 315
rect 2030 310 2036 311
rect 2022 305 2028 306
rect 2022 301 2023 305
rect 2027 301 2028 305
rect 2022 300 2028 301
rect 1862 292 1868 293
rect 1822 288 1828 289
rect 1822 284 1823 288
rect 1827 284 1828 288
rect 1862 288 1863 292
rect 1867 288 1868 292
rect 1862 287 1868 288
rect 1234 282 1240 283
rect 1242 283 1248 284
rect 1822 283 1828 284
rect 1242 279 1243 283
rect 1247 279 1248 283
rect 1242 278 1248 279
rect 1862 275 1868 276
rect 110 271 116 272
rect 110 267 111 271
rect 115 267 116 271
rect 110 266 116 267
rect 810 271 816 272
rect 810 267 811 271
rect 815 267 816 271
rect 810 266 816 267
rect 1410 271 1416 272
rect 1410 267 1411 271
rect 1415 267 1416 271
rect 1410 266 1416 267
rect 1822 271 1828 272
rect 1822 267 1823 271
rect 1827 267 1828 271
rect 1862 271 1863 275
rect 1867 271 1868 275
rect 1862 270 1868 271
rect 1822 266 1828 267
rect 112 247 114 266
rect 254 261 260 262
rect 254 257 255 261
rect 259 257 260 261
rect 254 256 260 257
rect 382 261 388 262
rect 382 257 383 261
rect 387 257 388 261
rect 382 256 388 257
rect 518 261 524 262
rect 518 257 519 261
rect 523 257 524 261
rect 518 256 524 257
rect 670 261 676 262
rect 670 257 671 261
rect 675 257 676 261
rect 670 256 676 257
rect 256 247 258 256
rect 384 247 386 256
rect 520 247 522 256
rect 672 247 674 256
rect 111 246 115 247
rect 111 241 115 242
rect 255 246 259 247
rect 255 241 259 242
rect 383 246 387 247
rect 383 241 387 242
rect 399 246 403 247
rect 399 241 403 242
rect 503 246 507 247
rect 503 241 507 242
rect 519 246 523 247
rect 519 241 523 242
rect 615 246 619 247
rect 615 241 619 242
rect 671 246 675 247
rect 671 241 675 242
rect 735 246 739 247
rect 735 241 739 242
rect 112 226 114 241
rect 400 236 402 241
rect 504 236 506 241
rect 616 236 618 241
rect 736 236 738 241
rect 398 235 404 236
rect 398 231 399 235
rect 403 231 404 235
rect 398 230 404 231
rect 502 235 508 236
rect 502 231 503 235
rect 507 231 508 235
rect 502 230 508 231
rect 614 235 620 236
rect 614 231 615 235
rect 619 231 620 235
rect 614 230 620 231
rect 734 235 740 236
rect 734 231 735 235
rect 739 231 740 235
rect 734 230 740 231
rect 802 227 808 228
rect 110 225 116 226
rect 110 221 111 225
rect 115 221 116 225
rect 802 223 803 227
rect 807 223 808 227
rect 802 222 808 223
rect 110 220 116 221
rect 110 208 116 209
rect 110 204 111 208
rect 115 204 116 208
rect 110 203 116 204
rect 112 159 114 203
rect 406 195 412 196
rect 406 191 407 195
rect 411 191 412 195
rect 406 190 412 191
rect 510 195 516 196
rect 510 191 511 195
rect 515 191 516 195
rect 510 190 516 191
rect 622 195 628 196
rect 622 191 623 195
rect 627 191 628 195
rect 622 190 628 191
rect 742 195 748 196
rect 742 191 743 195
rect 747 191 748 195
rect 742 190 748 191
rect 408 159 410 190
rect 419 188 423 189
rect 418 183 424 184
rect 418 179 419 183
rect 423 179 424 183
rect 418 178 424 179
rect 512 159 514 190
rect 624 159 626 190
rect 744 159 746 190
rect 804 160 806 222
rect 812 189 814 266
rect 830 261 836 262
rect 830 257 831 261
rect 835 257 836 261
rect 830 256 836 257
rect 998 261 1004 262
rect 998 257 999 261
rect 1003 257 1004 261
rect 998 256 1004 257
rect 1166 261 1172 262
rect 1166 257 1167 261
rect 1171 257 1172 261
rect 1166 256 1172 257
rect 1334 261 1340 262
rect 1334 257 1335 261
rect 1339 257 1340 261
rect 1334 256 1340 257
rect 832 247 834 256
rect 1000 247 1002 256
rect 1168 247 1170 256
rect 1336 247 1338 256
rect 831 246 835 247
rect 831 241 835 242
rect 863 246 867 247
rect 863 241 867 242
rect 991 246 995 247
rect 991 241 995 242
rect 999 246 1003 247
rect 999 241 1003 242
rect 1119 246 1123 247
rect 1119 241 1123 242
rect 1167 246 1171 247
rect 1167 241 1171 242
rect 1247 246 1251 247
rect 1247 241 1251 242
rect 1335 246 1339 247
rect 1335 241 1339 242
rect 1375 246 1379 247
rect 1375 241 1379 242
rect 864 236 866 241
rect 992 236 994 241
rect 1120 236 1122 241
rect 1248 236 1250 241
rect 1376 236 1378 241
rect 862 235 868 236
rect 862 231 863 235
rect 867 231 868 235
rect 862 230 868 231
rect 990 235 996 236
rect 990 231 991 235
rect 995 231 996 235
rect 990 230 996 231
rect 1118 235 1124 236
rect 1118 231 1119 235
rect 1123 231 1124 235
rect 1118 230 1124 231
rect 1246 235 1252 236
rect 1246 231 1247 235
rect 1251 231 1252 235
rect 1246 230 1252 231
rect 1374 235 1380 236
rect 1374 231 1375 235
rect 1379 231 1380 235
rect 1374 230 1380 231
rect 1058 211 1064 212
rect 1058 207 1059 211
rect 1063 207 1064 211
rect 1058 206 1064 207
rect 1214 211 1220 212
rect 1214 207 1215 211
rect 1219 207 1220 211
rect 1214 206 1220 207
rect 870 195 876 196
rect 870 191 871 195
rect 875 191 876 195
rect 870 190 876 191
rect 998 195 1004 196
rect 998 191 999 195
rect 1003 191 1004 195
rect 998 190 1004 191
rect 811 188 815 189
rect 811 183 815 184
rect 802 159 808 160
rect 872 159 874 190
rect 1000 159 1002 190
rect 1060 184 1062 206
rect 1126 195 1132 196
rect 1126 191 1127 195
rect 1131 191 1132 195
rect 1126 190 1132 191
rect 1058 183 1064 184
rect 1058 179 1059 183
rect 1063 179 1064 183
rect 1058 178 1064 179
rect 1128 159 1130 190
rect 1216 184 1218 206
rect 1254 195 1260 196
rect 1254 191 1255 195
rect 1259 191 1260 195
rect 1254 190 1260 191
rect 1382 195 1388 196
rect 1382 191 1383 195
rect 1387 191 1388 195
rect 1382 190 1388 191
rect 1214 183 1220 184
rect 1214 179 1215 183
rect 1219 179 1220 183
rect 1214 178 1220 179
rect 1256 159 1258 190
rect 1384 159 1386 190
rect 1412 184 1414 266
rect 1502 261 1508 262
rect 1502 257 1503 261
rect 1507 257 1508 261
rect 1502 256 1508 257
rect 1678 261 1684 262
rect 1678 257 1679 261
rect 1683 257 1684 261
rect 1678 256 1684 257
rect 1504 247 1506 256
rect 1680 247 1682 256
rect 1824 247 1826 266
rect 1864 255 1866 270
rect 2014 265 2020 266
rect 2014 261 2015 265
rect 2019 261 2020 265
rect 2014 260 2020 261
rect 2016 255 2018 260
rect 1863 254 1867 255
rect 1863 249 1867 250
rect 1959 254 1963 255
rect 1959 249 1963 250
rect 2015 254 2019 255
rect 2015 249 2019 250
rect 1495 246 1499 247
rect 1495 241 1499 242
rect 1503 246 1507 247
rect 1503 241 1507 242
rect 1623 246 1627 247
rect 1623 241 1627 242
rect 1679 246 1683 247
rect 1679 241 1683 242
rect 1727 246 1731 247
rect 1727 241 1731 242
rect 1823 246 1827 247
rect 1823 241 1827 242
rect 1496 236 1498 241
rect 1624 236 1626 241
rect 1728 236 1730 241
rect 1494 235 1500 236
rect 1494 231 1495 235
rect 1499 231 1500 235
rect 1494 230 1500 231
rect 1622 235 1628 236
rect 1622 231 1623 235
rect 1627 231 1628 235
rect 1622 230 1628 231
rect 1726 235 1732 236
rect 1726 231 1727 235
rect 1731 231 1732 235
rect 1726 230 1732 231
rect 1824 226 1826 241
rect 1864 234 1866 249
rect 1960 244 1962 249
rect 1958 243 1964 244
rect 1958 239 1959 243
rect 1963 239 1964 243
rect 1958 238 1964 239
rect 2032 236 2034 310
rect 2120 306 2122 317
rect 2118 305 2124 306
rect 2118 301 2119 305
rect 2123 301 2124 305
rect 2118 300 2124 301
rect 2216 293 2218 322
rect 2223 317 2227 318
rect 2247 322 2251 323
rect 2247 317 2251 318
rect 2327 322 2331 323
rect 2327 317 2331 318
rect 2335 322 2339 323
rect 2335 317 2339 318
rect 2423 322 2427 323
rect 2423 317 2427 318
rect 2431 322 2435 323
rect 2431 317 2435 318
rect 2511 322 2515 323
rect 2511 317 2515 318
rect 2535 322 2539 323
rect 2535 317 2539 318
rect 2224 306 2226 317
rect 2328 306 2330 317
rect 2390 315 2396 316
rect 2390 311 2391 315
rect 2395 311 2396 315
rect 2390 310 2396 311
rect 2222 305 2228 306
rect 2222 301 2223 305
rect 2227 301 2228 305
rect 2222 300 2228 301
rect 2326 305 2332 306
rect 2326 301 2327 305
rect 2331 301 2332 305
rect 2326 300 2332 301
rect 2215 292 2219 293
rect 2392 292 2394 310
rect 2432 306 2434 317
rect 2536 306 2538 317
rect 2572 316 2574 350
rect 2622 339 2628 340
rect 2622 335 2623 339
rect 2627 335 2628 339
rect 2622 334 2628 335
rect 2624 323 2626 334
rect 2684 328 2686 350
rect 2758 339 2764 340
rect 2758 335 2759 339
rect 2763 335 2764 339
rect 2758 334 2764 335
rect 2926 339 2932 340
rect 2926 335 2927 339
rect 2931 335 2932 339
rect 2926 334 2932 335
rect 2682 327 2688 328
rect 2682 323 2683 327
rect 2687 323 2688 327
rect 2760 323 2762 334
rect 2771 332 2775 333
rect 2770 327 2776 328
rect 2770 323 2771 327
rect 2775 323 2776 327
rect 2928 323 2930 334
rect 2936 328 2938 406
rect 2998 401 3004 402
rect 2998 397 2999 401
rect 3003 397 3004 401
rect 2998 396 3004 397
rect 3158 401 3164 402
rect 3158 397 3159 401
rect 3163 397 3164 401
rect 3158 396 3164 397
rect 3326 401 3332 402
rect 3326 397 3327 401
rect 3331 397 3332 401
rect 3326 396 3332 397
rect 3478 401 3484 402
rect 3478 397 3479 401
rect 3483 397 3484 401
rect 3478 396 3484 397
rect 3000 391 3002 396
rect 3160 391 3162 396
rect 3328 391 3330 396
rect 3480 391 3482 396
rect 3576 391 3578 406
rect 2999 390 3003 391
rect 2999 385 3003 386
rect 3103 390 3107 391
rect 3103 385 3107 386
rect 3159 390 3163 391
rect 3159 385 3163 386
rect 3303 390 3307 391
rect 3303 385 3307 386
rect 3327 390 3331 391
rect 3327 385 3331 386
rect 3479 390 3483 391
rect 3479 385 3483 386
rect 3575 390 3579 391
rect 3575 385 3579 386
rect 3104 380 3106 385
rect 3304 380 3306 385
rect 3480 380 3482 385
rect 3102 379 3108 380
rect 3102 375 3103 379
rect 3107 375 3108 379
rect 3102 374 3108 375
rect 3302 379 3308 380
rect 3302 375 3303 379
rect 3307 375 3308 379
rect 3302 374 3308 375
rect 3478 379 3484 380
rect 3478 375 3479 379
rect 3483 375 3484 379
rect 3478 374 3484 375
rect 3198 371 3204 372
rect 3198 367 3199 371
rect 3203 367 3204 371
rect 3576 370 3578 385
rect 3198 366 3204 367
rect 3574 369 3580 370
rect 3110 339 3116 340
rect 3110 335 3111 339
rect 3115 335 3116 339
rect 3110 334 3116 335
rect 2934 327 2940 328
rect 2934 323 2935 327
rect 2939 323 2940 327
rect 3112 323 3114 334
rect 3200 333 3202 366
rect 3574 365 3575 369
rect 3579 365 3580 369
rect 3574 364 3580 365
rect 3574 352 3580 353
rect 3574 348 3575 352
rect 3579 348 3580 352
rect 3574 347 3580 348
rect 3310 339 3316 340
rect 3310 335 3311 339
rect 3315 335 3316 339
rect 3310 334 3316 335
rect 3486 339 3492 340
rect 3486 335 3487 339
rect 3491 335 3492 339
rect 3486 334 3492 335
rect 3199 332 3203 333
rect 3199 327 3203 328
rect 3312 323 3314 334
rect 3488 323 3490 334
rect 3576 323 3578 347
rect 2623 322 2627 323
rect 2623 317 2627 318
rect 2639 322 2643 323
rect 2682 322 2688 323
rect 2743 322 2747 323
rect 2639 317 2643 318
rect 2743 317 2747 318
rect 2759 322 2763 323
rect 2770 322 2776 323
rect 2855 322 2859 323
rect 2759 317 2763 318
rect 2855 317 2859 318
rect 2927 322 2931 323
rect 2934 322 2940 323
rect 2967 322 2971 323
rect 2927 317 2931 318
rect 2967 317 2971 318
rect 3111 322 3115 323
rect 3111 317 3115 318
rect 3311 322 3315 323
rect 3311 317 3315 318
rect 3487 322 3491 323
rect 3487 317 3491 318
rect 3575 322 3579 323
rect 3575 317 3579 318
rect 2570 315 2576 316
rect 2570 311 2571 315
rect 2575 311 2576 315
rect 2570 310 2576 311
rect 2640 306 2642 317
rect 2744 306 2746 317
rect 2856 306 2858 317
rect 2968 306 2970 317
rect 2430 305 2436 306
rect 2430 301 2431 305
rect 2435 301 2436 305
rect 2430 300 2436 301
rect 2534 305 2540 306
rect 2534 301 2535 305
rect 2539 301 2540 305
rect 2534 300 2540 301
rect 2638 305 2644 306
rect 2638 301 2639 305
rect 2643 301 2644 305
rect 2638 300 2644 301
rect 2742 305 2748 306
rect 2742 301 2743 305
rect 2747 301 2748 305
rect 2742 300 2748 301
rect 2854 305 2860 306
rect 2854 301 2855 305
rect 2859 301 2860 305
rect 2854 300 2860 301
rect 2966 305 2972 306
rect 2966 301 2967 305
rect 2971 301 2972 305
rect 2966 300 2972 301
rect 3576 293 3578 317
rect 2399 292 2403 293
rect 2215 287 2219 288
rect 2390 291 2396 292
rect 2390 287 2391 291
rect 2395 287 2396 291
rect 3574 292 3580 293
rect 3574 288 3575 292
rect 3579 288 3580 292
rect 2390 286 2396 287
rect 2398 287 2404 288
rect 3574 287 3580 288
rect 2398 283 2399 287
rect 2403 283 2404 287
rect 2398 282 2404 283
rect 2922 275 2928 276
rect 2922 271 2923 275
rect 2927 271 2928 275
rect 2922 270 2928 271
rect 3574 275 3580 276
rect 3574 271 3575 275
rect 3579 271 3580 275
rect 3574 270 3580 271
rect 2110 265 2116 266
rect 2110 261 2111 265
rect 2115 261 2116 265
rect 2110 260 2116 261
rect 2214 265 2220 266
rect 2214 261 2215 265
rect 2219 261 2220 265
rect 2214 260 2220 261
rect 2318 265 2324 266
rect 2318 261 2319 265
rect 2323 261 2324 265
rect 2318 260 2324 261
rect 2422 265 2428 266
rect 2422 261 2423 265
rect 2427 261 2428 265
rect 2422 260 2428 261
rect 2526 265 2532 266
rect 2526 261 2527 265
rect 2531 261 2532 265
rect 2526 260 2532 261
rect 2630 265 2636 266
rect 2630 261 2631 265
rect 2635 261 2636 265
rect 2630 260 2636 261
rect 2734 265 2740 266
rect 2734 261 2735 265
rect 2739 261 2740 265
rect 2734 260 2740 261
rect 2846 265 2852 266
rect 2846 261 2847 265
rect 2851 261 2852 265
rect 2846 260 2852 261
rect 2112 255 2114 260
rect 2216 255 2218 260
rect 2320 255 2322 260
rect 2424 255 2426 260
rect 2528 255 2530 260
rect 2632 255 2634 260
rect 2736 255 2738 260
rect 2848 255 2850 260
rect 2111 254 2115 255
rect 2111 249 2115 250
rect 2175 254 2179 255
rect 2175 249 2179 250
rect 2215 254 2219 255
rect 2215 249 2219 250
rect 2319 254 2323 255
rect 2319 249 2323 250
rect 2383 254 2387 255
rect 2383 249 2387 250
rect 2423 254 2427 255
rect 2423 249 2427 250
rect 2527 254 2531 255
rect 2527 249 2531 250
rect 2583 254 2587 255
rect 2583 249 2587 250
rect 2631 254 2635 255
rect 2631 249 2635 250
rect 2735 254 2739 255
rect 2735 249 2739 250
rect 2767 254 2771 255
rect 2767 249 2771 250
rect 2847 254 2851 255
rect 2847 249 2851 250
rect 2176 244 2178 249
rect 2384 244 2386 249
rect 2584 244 2586 249
rect 2768 244 2770 249
rect 2174 243 2180 244
rect 2174 239 2175 243
rect 2179 239 2180 243
rect 2174 238 2180 239
rect 2382 243 2388 244
rect 2382 239 2383 243
rect 2387 239 2388 243
rect 2382 238 2388 239
rect 2582 243 2588 244
rect 2582 239 2583 243
rect 2587 239 2588 243
rect 2582 238 2588 239
rect 2766 243 2772 244
rect 2766 239 2767 243
rect 2771 239 2772 243
rect 2766 238 2772 239
rect 2030 235 2036 236
rect 1862 233 1868 234
rect 1862 229 1863 233
rect 1867 229 1868 233
rect 2030 231 2031 235
rect 2035 231 2036 235
rect 2030 230 2036 231
rect 1862 228 1868 229
rect 1822 225 1828 226
rect 1726 223 1732 224
rect 1726 219 1727 223
rect 1731 219 1732 223
rect 1822 221 1823 225
rect 1827 221 1828 225
rect 1822 220 1828 221
rect 1726 218 1732 219
rect 2094 219 2100 220
rect 1502 195 1508 196
rect 1502 191 1503 195
rect 1507 191 1508 195
rect 1502 190 1508 191
rect 1630 195 1636 196
rect 1630 191 1631 195
rect 1635 191 1636 195
rect 1630 190 1636 191
rect 1410 183 1416 184
rect 1410 179 1411 183
rect 1415 179 1416 183
rect 1410 178 1416 179
rect 1504 159 1506 190
rect 1632 159 1634 190
rect 111 158 115 159
rect 111 153 115 154
rect 223 158 227 159
rect 223 153 227 154
rect 311 158 315 159
rect 311 153 315 154
rect 399 158 403 159
rect 399 153 403 154
rect 407 158 411 159
rect 407 153 411 154
rect 487 158 491 159
rect 487 153 491 154
rect 511 158 515 159
rect 511 153 515 154
rect 575 158 579 159
rect 575 153 579 154
rect 623 158 627 159
rect 623 153 627 154
rect 663 158 667 159
rect 663 153 667 154
rect 743 158 747 159
rect 743 153 747 154
rect 751 158 755 159
rect 802 155 803 159
rect 807 155 808 159
rect 802 154 808 155
rect 839 158 843 159
rect 751 153 755 154
rect 839 153 843 154
rect 871 158 875 159
rect 871 153 875 154
rect 927 158 931 159
rect 927 153 931 154
rect 999 158 1003 159
rect 999 153 1003 154
rect 1015 158 1019 159
rect 1015 153 1019 154
rect 1103 158 1107 159
rect 1103 153 1107 154
rect 1127 158 1131 159
rect 1127 153 1131 154
rect 1191 158 1195 159
rect 1191 153 1195 154
rect 1255 158 1259 159
rect 1255 153 1259 154
rect 1295 158 1299 159
rect 1295 153 1299 154
rect 1383 158 1387 159
rect 1383 153 1387 154
rect 1399 158 1403 159
rect 1399 153 1403 154
rect 1503 158 1507 159
rect 1503 153 1507 154
rect 1511 158 1515 159
rect 1511 153 1515 154
rect 1631 158 1635 159
rect 1631 153 1635 154
rect 112 129 114 153
rect 224 142 226 153
rect 312 142 314 153
rect 400 142 402 153
rect 488 142 490 153
rect 576 142 578 153
rect 664 142 666 153
rect 752 142 754 153
rect 840 142 842 153
rect 928 142 930 153
rect 1016 142 1018 153
rect 1104 142 1106 153
rect 1162 151 1168 152
rect 1162 147 1163 151
rect 1167 147 1168 151
rect 1162 146 1168 147
rect 222 141 228 142
rect 222 137 223 141
rect 227 137 228 141
rect 222 136 228 137
rect 310 141 316 142
rect 310 137 311 141
rect 315 137 316 141
rect 310 136 316 137
rect 398 141 404 142
rect 398 137 399 141
rect 403 137 404 141
rect 398 136 404 137
rect 486 141 492 142
rect 486 137 487 141
rect 491 137 492 141
rect 486 136 492 137
rect 574 141 580 142
rect 574 137 575 141
rect 579 137 580 141
rect 574 136 580 137
rect 662 141 668 142
rect 662 137 663 141
rect 667 137 668 141
rect 662 136 668 137
rect 750 141 756 142
rect 750 137 751 141
rect 755 137 756 141
rect 750 136 756 137
rect 838 141 844 142
rect 838 137 839 141
rect 843 137 844 141
rect 838 136 844 137
rect 926 141 932 142
rect 926 137 927 141
rect 931 137 932 141
rect 926 136 932 137
rect 1014 141 1020 142
rect 1014 137 1015 141
rect 1019 137 1020 141
rect 1014 136 1020 137
rect 1102 141 1108 142
rect 1102 137 1103 141
rect 1107 137 1108 141
rect 1102 136 1108 137
rect 110 128 116 129
rect 1164 128 1166 146
rect 1192 142 1194 153
rect 1296 142 1298 153
rect 1400 142 1402 153
rect 1512 142 1514 153
rect 1632 142 1634 153
rect 1728 152 1730 218
rect 1862 216 1868 217
rect 1862 212 1863 216
rect 1867 212 1868 216
rect 2094 215 2095 219
rect 2099 215 2100 219
rect 2094 214 2100 215
rect 2242 219 2248 220
rect 2242 215 2243 219
rect 2247 215 2248 219
rect 2242 214 2248 215
rect 1862 211 1868 212
rect 1822 208 1828 209
rect 1822 204 1823 208
rect 1827 204 1828 208
rect 1822 203 1828 204
rect 1734 195 1740 196
rect 1734 191 1735 195
rect 1739 191 1740 195
rect 1734 190 1740 191
rect 1736 159 1738 190
rect 1824 159 1826 203
rect 1735 158 1739 159
rect 1735 153 1739 154
rect 1823 158 1827 159
rect 1864 155 1866 211
rect 1966 203 1972 204
rect 1966 199 1967 203
rect 1971 199 1972 203
rect 1966 198 1972 199
rect 1968 155 1970 198
rect 2096 192 2098 214
rect 2182 203 2188 204
rect 2182 199 2183 203
rect 2187 199 2188 203
rect 2182 198 2188 199
rect 2094 191 2100 192
rect 2094 187 2095 191
rect 2099 187 2100 191
rect 2094 186 2100 187
rect 2184 155 2186 198
rect 2244 192 2246 214
rect 2390 203 2396 204
rect 2390 199 2391 203
rect 2395 199 2396 203
rect 2390 198 2396 199
rect 2590 203 2596 204
rect 2590 199 2591 203
rect 2595 199 2596 203
rect 2590 198 2596 199
rect 2774 203 2780 204
rect 2774 199 2775 203
rect 2779 199 2780 203
rect 2774 198 2780 199
rect 2242 191 2248 192
rect 2242 187 2243 191
rect 2247 187 2248 191
rect 2242 186 2248 187
rect 2392 155 2394 198
rect 2450 191 2456 192
rect 2450 187 2451 191
rect 2455 187 2456 191
rect 2450 186 2456 187
rect 1823 153 1827 154
rect 1863 154 1867 155
rect 1726 151 1732 152
rect 1726 147 1727 151
rect 1731 147 1732 151
rect 1726 146 1732 147
rect 1736 142 1738 153
rect 1190 141 1196 142
rect 1190 137 1191 141
rect 1195 137 1196 141
rect 1190 136 1196 137
rect 1294 141 1300 142
rect 1294 137 1295 141
rect 1299 137 1300 141
rect 1294 136 1300 137
rect 1398 141 1404 142
rect 1398 137 1399 141
rect 1403 137 1404 141
rect 1398 136 1404 137
rect 1510 141 1516 142
rect 1510 137 1511 141
rect 1515 137 1516 141
rect 1510 136 1516 137
rect 1630 141 1636 142
rect 1630 137 1631 141
rect 1635 137 1636 141
rect 1630 136 1636 137
rect 1734 141 1740 142
rect 1734 137 1735 141
rect 1739 137 1740 141
rect 1734 136 1740 137
rect 1824 129 1826 153
rect 1863 149 1867 150
rect 1895 154 1899 155
rect 1895 149 1899 150
rect 1967 154 1971 155
rect 1967 149 1971 150
rect 1983 154 1987 155
rect 1983 149 1987 150
rect 2071 154 2075 155
rect 2071 149 2075 150
rect 2159 154 2163 155
rect 2159 149 2163 150
rect 2183 154 2187 155
rect 2183 149 2187 150
rect 2271 154 2275 155
rect 2271 149 2275 150
rect 2383 154 2387 155
rect 2383 149 2387 150
rect 2391 154 2395 155
rect 2391 149 2395 150
rect 1822 128 1828 129
rect 110 124 111 128
rect 115 124 116 128
rect 110 123 116 124
rect 1162 127 1168 128
rect 1162 123 1163 127
rect 1167 123 1168 127
rect 1822 124 1823 128
rect 1827 124 1828 128
rect 1864 125 1866 149
rect 1896 138 1898 149
rect 1984 138 1986 149
rect 2072 138 2074 149
rect 2160 138 2162 149
rect 2272 138 2274 149
rect 2384 138 2386 149
rect 2442 147 2448 148
rect 2442 143 2443 147
rect 2447 143 2448 147
rect 2442 142 2448 143
rect 1894 137 1900 138
rect 1894 133 1895 137
rect 1899 133 1900 137
rect 1894 132 1900 133
rect 1982 137 1988 138
rect 1982 133 1983 137
rect 1987 133 1988 137
rect 1982 132 1988 133
rect 2070 137 2076 138
rect 2070 133 2071 137
rect 2075 133 2076 137
rect 2070 132 2076 133
rect 2158 137 2164 138
rect 2158 133 2159 137
rect 2163 133 2164 137
rect 2158 132 2164 133
rect 2270 137 2276 138
rect 2270 133 2271 137
rect 2275 133 2276 137
rect 2270 132 2276 133
rect 2382 137 2388 138
rect 2382 133 2383 137
rect 2387 133 2388 137
rect 2382 132 2388 133
rect 1822 123 1828 124
rect 1862 124 1868 125
rect 2444 124 2446 142
rect 1162 122 1168 123
rect 1862 120 1863 124
rect 1867 120 1868 124
rect 1862 119 1868 120
rect 2442 123 2448 124
rect 2442 119 2443 123
rect 2447 119 2448 123
rect 2452 120 2454 186
rect 2592 155 2594 198
rect 2603 196 2607 197
rect 2602 191 2608 192
rect 2602 187 2603 191
rect 2607 187 2608 191
rect 2602 186 2608 187
rect 2619 164 2623 165
rect 2619 159 2623 160
rect 2495 154 2499 155
rect 2495 149 2499 150
rect 2591 154 2595 155
rect 2591 149 2595 150
rect 2607 154 2611 155
rect 2607 149 2611 150
rect 2496 138 2498 149
rect 2608 138 2610 149
rect 2620 148 2622 159
rect 2776 155 2778 198
rect 2924 197 2926 270
rect 2958 265 2964 266
rect 2958 261 2959 265
rect 2963 261 2964 265
rect 2958 260 2964 261
rect 2960 255 2962 260
rect 3576 255 3578 270
rect 2951 254 2955 255
rect 2951 249 2955 250
rect 2959 254 2963 255
rect 2959 249 2963 250
rect 3127 254 3131 255
rect 3127 249 3131 250
rect 3311 254 3315 255
rect 3311 249 3315 250
rect 3479 254 3483 255
rect 3479 249 3483 250
rect 3575 254 3579 255
rect 3575 249 3579 250
rect 2952 244 2954 249
rect 3128 244 3130 249
rect 3312 244 3314 249
rect 3480 244 3482 249
rect 2950 243 2956 244
rect 2950 239 2951 243
rect 2955 239 2956 243
rect 2950 238 2956 239
rect 3126 243 3132 244
rect 3126 239 3127 243
rect 3131 239 3132 243
rect 3126 238 3132 239
rect 3310 243 3316 244
rect 3310 239 3311 243
rect 3315 239 3316 243
rect 3310 238 3316 239
rect 3478 243 3484 244
rect 3478 239 3479 243
rect 3483 239 3484 243
rect 3478 238 3484 239
rect 3198 235 3204 236
rect 3198 231 3199 235
rect 3203 231 3204 235
rect 3576 234 3578 249
rect 3198 230 3204 231
rect 3574 233 3580 234
rect 2958 203 2964 204
rect 2958 199 2959 203
rect 2963 199 2964 203
rect 2958 198 2964 199
rect 3134 203 3140 204
rect 3134 199 3135 203
rect 3139 199 3140 203
rect 3134 198 3140 199
rect 2923 196 2927 197
rect 2923 191 2927 192
rect 2960 155 2962 198
rect 3136 155 3138 198
rect 3200 165 3202 230
rect 3574 229 3575 233
rect 3579 229 3580 233
rect 3574 228 3580 229
rect 3574 216 3580 217
rect 3574 212 3575 216
rect 3579 212 3580 216
rect 3574 211 3580 212
rect 3318 203 3324 204
rect 3318 199 3319 203
rect 3323 199 3324 203
rect 3318 198 3324 199
rect 3486 203 3492 204
rect 3486 199 3487 203
rect 3491 199 3492 203
rect 3486 198 3492 199
rect 3199 164 3203 165
rect 3199 159 3203 160
rect 3320 155 3322 198
rect 3478 191 3484 192
rect 3478 187 3479 191
rect 3483 187 3484 191
rect 3478 186 3484 187
rect 2719 154 2723 155
rect 2719 149 2723 150
rect 2775 154 2779 155
rect 2775 149 2779 150
rect 2823 154 2827 155
rect 2823 149 2827 150
rect 2927 154 2931 155
rect 2927 149 2931 150
rect 2959 154 2963 155
rect 2959 149 2963 150
rect 3023 154 3027 155
rect 3023 149 3027 150
rect 3119 154 3123 155
rect 3119 149 3123 150
rect 3135 154 3139 155
rect 3135 149 3139 150
rect 3215 154 3219 155
rect 3215 149 3219 150
rect 3311 154 3315 155
rect 3311 149 3315 150
rect 3319 154 3323 155
rect 3319 149 3323 150
rect 3399 154 3403 155
rect 3399 149 3403 150
rect 2618 147 2624 148
rect 2618 143 2619 147
rect 2623 143 2624 147
rect 2618 142 2624 143
rect 2720 138 2722 149
rect 2824 138 2826 149
rect 2928 138 2930 149
rect 3024 138 3026 149
rect 3120 138 3122 149
rect 3216 138 3218 149
rect 3312 138 3314 149
rect 3400 138 3402 149
rect 2494 137 2500 138
rect 2494 133 2495 137
rect 2499 133 2500 137
rect 2494 132 2500 133
rect 2606 137 2612 138
rect 2606 133 2607 137
rect 2611 133 2612 137
rect 2606 132 2612 133
rect 2718 137 2724 138
rect 2718 133 2719 137
rect 2723 133 2724 137
rect 2718 132 2724 133
rect 2822 137 2828 138
rect 2822 133 2823 137
rect 2827 133 2828 137
rect 2822 132 2828 133
rect 2926 137 2932 138
rect 2926 133 2927 137
rect 2931 133 2932 137
rect 2926 132 2932 133
rect 3022 137 3028 138
rect 3022 133 3023 137
rect 3027 133 3028 137
rect 3022 132 3028 133
rect 3118 137 3124 138
rect 3118 133 3119 137
rect 3123 133 3124 137
rect 3118 132 3124 133
rect 3214 137 3220 138
rect 3214 133 3215 137
rect 3219 133 3220 137
rect 3214 132 3220 133
rect 3310 137 3316 138
rect 3310 133 3311 137
rect 3315 133 3316 137
rect 3310 132 3316 133
rect 3398 137 3404 138
rect 3398 133 3399 137
rect 3403 133 3404 137
rect 3398 132 3404 133
rect 3480 120 3482 186
rect 3488 155 3490 198
rect 3576 155 3578 211
rect 3487 154 3491 155
rect 3487 149 3491 150
rect 3575 154 3579 155
rect 3575 149 3579 150
rect 3488 138 3490 149
rect 3486 137 3492 138
rect 3486 133 3487 137
rect 3491 133 3492 137
rect 3486 132 3492 133
rect 3576 125 3578 149
rect 3574 124 3580 125
rect 3574 120 3575 124
rect 3579 120 3580 124
rect 2442 118 2448 119
rect 2450 119 2456 120
rect 2450 115 2451 119
rect 2455 115 2456 119
rect 2450 114 2456 115
rect 3478 119 3484 120
rect 3574 119 3580 120
rect 3478 115 3479 119
rect 3483 115 3484 119
rect 3478 114 3484 115
rect 110 111 116 112
rect 110 107 111 111
rect 115 107 116 111
rect 110 106 116 107
rect 1822 111 1828 112
rect 1822 107 1823 111
rect 1827 107 1828 111
rect 1822 106 1828 107
rect 1862 107 1868 108
rect 112 91 114 106
rect 214 101 220 102
rect 214 97 215 101
rect 219 97 220 101
rect 214 96 220 97
rect 302 101 308 102
rect 302 97 303 101
rect 307 97 308 101
rect 302 96 308 97
rect 390 101 396 102
rect 390 97 391 101
rect 395 97 396 101
rect 390 96 396 97
rect 478 101 484 102
rect 478 97 479 101
rect 483 97 484 101
rect 478 96 484 97
rect 566 101 572 102
rect 566 97 567 101
rect 571 97 572 101
rect 566 96 572 97
rect 654 101 660 102
rect 654 97 655 101
rect 659 97 660 101
rect 654 96 660 97
rect 742 101 748 102
rect 742 97 743 101
rect 747 97 748 101
rect 742 96 748 97
rect 830 101 836 102
rect 830 97 831 101
rect 835 97 836 101
rect 830 96 836 97
rect 918 101 924 102
rect 918 97 919 101
rect 923 97 924 101
rect 918 96 924 97
rect 1006 101 1012 102
rect 1006 97 1007 101
rect 1011 97 1012 101
rect 1006 96 1012 97
rect 1094 101 1100 102
rect 1094 97 1095 101
rect 1099 97 1100 101
rect 1094 96 1100 97
rect 1182 101 1188 102
rect 1182 97 1183 101
rect 1187 97 1188 101
rect 1182 96 1188 97
rect 1286 101 1292 102
rect 1286 97 1287 101
rect 1291 97 1292 101
rect 1286 96 1292 97
rect 1390 101 1396 102
rect 1390 97 1391 101
rect 1395 97 1396 101
rect 1390 96 1396 97
rect 1502 101 1508 102
rect 1502 97 1503 101
rect 1507 97 1508 101
rect 1502 96 1508 97
rect 1622 101 1628 102
rect 1622 97 1623 101
rect 1627 97 1628 101
rect 1622 96 1628 97
rect 1726 101 1732 102
rect 1726 97 1727 101
rect 1731 97 1732 101
rect 1726 96 1732 97
rect 216 91 218 96
rect 304 91 306 96
rect 392 91 394 96
rect 480 91 482 96
rect 568 91 570 96
rect 656 91 658 96
rect 744 91 746 96
rect 832 91 834 96
rect 920 91 922 96
rect 1008 91 1010 96
rect 1096 91 1098 96
rect 1184 91 1186 96
rect 1288 91 1290 96
rect 1392 91 1394 96
rect 1504 91 1506 96
rect 1624 91 1626 96
rect 1728 91 1730 96
rect 1824 91 1826 106
rect 1862 103 1863 107
rect 1867 103 1868 107
rect 1862 102 1868 103
rect 3574 107 3580 108
rect 3574 103 3575 107
rect 3579 103 3580 107
rect 3574 102 3580 103
rect 111 90 115 91
rect 111 85 115 86
rect 215 90 219 91
rect 215 85 219 86
rect 303 90 307 91
rect 303 85 307 86
rect 391 90 395 91
rect 391 85 395 86
rect 479 90 483 91
rect 479 85 483 86
rect 567 90 571 91
rect 567 85 571 86
rect 655 90 659 91
rect 655 85 659 86
rect 743 90 747 91
rect 743 85 747 86
rect 831 90 835 91
rect 831 85 835 86
rect 919 90 923 91
rect 919 85 923 86
rect 1007 90 1011 91
rect 1007 85 1011 86
rect 1095 90 1099 91
rect 1095 85 1099 86
rect 1183 90 1187 91
rect 1183 85 1187 86
rect 1287 90 1291 91
rect 1287 85 1291 86
rect 1391 90 1395 91
rect 1391 85 1395 86
rect 1503 90 1507 91
rect 1503 85 1507 86
rect 1623 90 1627 91
rect 1623 85 1627 86
rect 1727 90 1731 91
rect 1727 85 1731 86
rect 1823 90 1827 91
rect 1864 87 1866 102
rect 1886 97 1892 98
rect 1886 93 1887 97
rect 1891 93 1892 97
rect 1886 92 1892 93
rect 1974 97 1980 98
rect 1974 93 1975 97
rect 1979 93 1980 97
rect 1974 92 1980 93
rect 2062 97 2068 98
rect 2062 93 2063 97
rect 2067 93 2068 97
rect 2062 92 2068 93
rect 2150 97 2156 98
rect 2150 93 2151 97
rect 2155 93 2156 97
rect 2150 92 2156 93
rect 2262 97 2268 98
rect 2262 93 2263 97
rect 2267 93 2268 97
rect 2262 92 2268 93
rect 2374 97 2380 98
rect 2374 93 2375 97
rect 2379 93 2380 97
rect 2374 92 2380 93
rect 2486 97 2492 98
rect 2486 93 2487 97
rect 2491 93 2492 97
rect 2486 92 2492 93
rect 2598 97 2604 98
rect 2598 93 2599 97
rect 2603 93 2604 97
rect 2598 92 2604 93
rect 2710 97 2716 98
rect 2710 93 2711 97
rect 2715 93 2716 97
rect 2710 92 2716 93
rect 2814 97 2820 98
rect 2814 93 2815 97
rect 2819 93 2820 97
rect 2814 92 2820 93
rect 2918 97 2924 98
rect 2918 93 2919 97
rect 2923 93 2924 97
rect 2918 92 2924 93
rect 3014 97 3020 98
rect 3014 93 3015 97
rect 3019 93 3020 97
rect 3014 92 3020 93
rect 3110 97 3116 98
rect 3110 93 3111 97
rect 3115 93 3116 97
rect 3110 92 3116 93
rect 3206 97 3212 98
rect 3206 93 3207 97
rect 3211 93 3212 97
rect 3206 92 3212 93
rect 3302 97 3308 98
rect 3302 93 3303 97
rect 3307 93 3308 97
rect 3302 92 3308 93
rect 3390 97 3396 98
rect 3390 93 3391 97
rect 3395 93 3396 97
rect 3390 92 3396 93
rect 3478 97 3484 98
rect 3478 93 3479 97
rect 3483 93 3484 97
rect 3478 92 3484 93
rect 1888 87 1890 92
rect 1976 87 1978 92
rect 2064 87 2066 92
rect 2152 87 2154 92
rect 2264 87 2266 92
rect 2376 87 2378 92
rect 2488 87 2490 92
rect 2600 87 2602 92
rect 2712 87 2714 92
rect 2816 87 2818 92
rect 2920 87 2922 92
rect 3016 87 3018 92
rect 3112 87 3114 92
rect 3208 87 3210 92
rect 3304 87 3306 92
rect 3392 87 3394 92
rect 3480 87 3482 92
rect 3576 87 3578 102
rect 1823 85 1827 86
rect 1863 86 1867 87
rect 1863 81 1867 82
rect 1887 86 1891 87
rect 1887 81 1891 82
rect 1975 86 1979 87
rect 1975 81 1979 82
rect 2063 86 2067 87
rect 2063 81 2067 82
rect 2151 86 2155 87
rect 2151 81 2155 82
rect 2263 86 2267 87
rect 2263 81 2267 82
rect 2375 86 2379 87
rect 2375 81 2379 82
rect 2487 86 2491 87
rect 2487 81 2491 82
rect 2599 86 2603 87
rect 2599 81 2603 82
rect 2711 86 2715 87
rect 2711 81 2715 82
rect 2815 86 2819 87
rect 2815 81 2819 82
rect 2919 86 2923 87
rect 2919 81 2923 82
rect 3015 86 3019 87
rect 3015 81 3019 82
rect 3111 86 3115 87
rect 3111 81 3115 82
rect 3207 86 3211 87
rect 3207 81 3211 82
rect 3303 86 3307 87
rect 3303 81 3307 82
rect 3391 86 3395 87
rect 3391 81 3395 82
rect 3479 86 3483 87
rect 3479 81 3483 82
rect 3575 86 3579 87
rect 3575 81 3579 82
<< m4c >>
rect 111 3646 115 3650
rect 143 3646 147 3650
rect 231 3646 235 3650
rect 319 3646 323 3650
rect 407 3646 411 3650
rect 495 3646 499 3650
rect 583 3646 587 3650
rect 671 3646 675 3650
rect 1823 3646 1827 3650
rect 111 3570 115 3574
rect 135 3570 139 3574
rect 223 3570 227 3574
rect 287 3570 291 3574
rect 311 3570 315 3574
rect 399 3570 403 3574
rect 463 3570 467 3574
rect 487 3570 491 3574
rect 575 3570 579 3574
rect 631 3570 635 3574
rect 663 3570 667 3574
rect 791 3570 795 3574
rect 935 3570 939 3574
rect 1071 3570 1075 3574
rect 1191 3570 1195 3574
rect 1311 3570 1315 3574
rect 1423 3570 1427 3574
rect 1527 3570 1531 3574
rect 1639 3570 1643 3574
rect 1727 3570 1731 3574
rect 1823 3570 1827 3574
rect 167 3552 171 3556
rect 651 3552 655 3556
rect 159 3512 163 3516
rect 111 3502 115 3506
rect 143 3502 147 3506
rect 151 3502 155 3506
rect 559 3512 563 3516
rect 807 3515 811 3516
rect 807 3512 811 3515
rect 1395 3512 1399 3516
rect 295 3502 299 3506
rect 327 3502 331 3506
rect 471 3502 475 3506
rect 495 3502 499 3506
rect 639 3502 643 3506
rect 655 3502 659 3506
rect 799 3502 803 3506
rect 807 3502 811 3506
rect 943 3502 947 3506
rect 951 3502 955 3506
rect 1079 3502 1083 3506
rect 1087 3502 1091 3506
rect 1199 3502 1203 3506
rect 1207 3502 1211 3506
rect 1319 3502 1323 3506
rect 1431 3502 1435 3506
rect 1535 3502 1539 3506
rect 1647 3502 1651 3506
rect 1735 3502 1739 3506
rect 1823 3502 1827 3506
rect 1863 3498 1867 3502
rect 1895 3498 1899 3502
rect 1983 3498 1987 3502
rect 2071 3498 2075 3502
rect 2159 3498 2163 3502
rect 3575 3498 3579 3502
rect 879 3456 883 3460
rect 1647 3456 1651 3460
rect 111 3434 115 3438
rect 143 3434 147 3438
rect 215 3434 219 3438
rect 319 3434 323 3438
rect 431 3434 435 3438
rect 487 3434 491 3438
rect 235 3376 239 3380
rect 639 3434 643 3438
rect 647 3434 651 3438
rect 799 3434 803 3438
rect 847 3434 851 3438
rect 943 3434 947 3438
rect 1039 3434 1043 3438
rect 1079 3434 1083 3438
rect 1199 3434 1203 3438
rect 1223 3434 1227 3438
rect 1311 3434 1315 3438
rect 1399 3434 1403 3438
rect 1423 3434 1427 3438
rect 1527 3434 1531 3438
rect 1567 3434 1571 3438
rect 1639 3434 1643 3438
rect 1727 3434 1731 3438
rect 1823 3434 1827 3438
rect 1863 3430 1867 3434
rect 1887 3430 1891 3434
rect 563 3376 567 3380
rect 1207 3371 1211 3372
rect 1207 3368 1211 3371
rect 1583 3368 1587 3372
rect 111 3358 115 3362
rect 223 3358 227 3362
rect 239 3358 243 3362
rect 383 3358 387 3362
rect 439 3358 443 3362
rect 543 3358 547 3362
rect 647 3358 651 3362
rect 711 3358 715 3362
rect 855 3358 859 3362
rect 871 3358 875 3362
rect 1031 3358 1035 3362
rect 1047 3358 1051 3362
rect 1183 3358 1187 3362
rect 1231 3358 1235 3362
rect 1335 3358 1339 3362
rect 1407 3358 1411 3362
rect 1487 3358 1491 3362
rect 1575 3358 1579 3362
rect 111 3286 115 3290
rect 231 3286 235 3290
rect 239 3286 243 3290
rect 375 3286 379 3290
rect 407 3286 411 3290
rect 535 3286 539 3290
rect 575 3286 579 3290
rect 703 3286 707 3290
rect 743 3286 747 3290
rect 259 3232 263 3236
rect 499 3232 503 3236
rect 111 3206 115 3210
rect 175 3206 179 3210
rect 247 3206 251 3210
rect 375 3206 379 3210
rect 415 3206 419 3210
rect 559 3206 563 3210
rect 863 3286 867 3290
rect 895 3286 899 3290
rect 1023 3286 1027 3290
rect 1047 3286 1051 3290
rect 1907 3376 1911 3380
rect 1639 3358 1643 3362
rect 1735 3358 1739 3362
rect 1823 3358 1827 3362
rect 1863 3362 1867 3366
rect 1895 3362 1899 3366
rect 1975 3430 1979 3434
rect 1991 3430 1995 3434
rect 2063 3430 2067 3434
rect 2119 3430 2123 3434
rect 2151 3430 2155 3434
rect 2255 3430 2259 3434
rect 2391 3430 2395 3434
rect 2527 3430 2531 3434
rect 2655 3430 2659 3434
rect 2783 3430 2787 3434
rect 2919 3430 2923 3434
rect 3055 3430 3059 3434
rect 3575 3430 3579 3434
rect 2323 3376 2327 3380
rect 1999 3362 2003 3366
rect 2127 3362 2131 3366
rect 2135 3362 2139 3366
rect 2263 3362 2267 3366
rect 2279 3362 2283 3366
rect 2399 3362 2403 3366
rect 2423 3362 2427 3366
rect 2535 3362 2539 3366
rect 2559 3362 2563 3366
rect 2663 3362 2667 3366
rect 2695 3362 2699 3366
rect 2791 3362 2795 3366
rect 2831 3362 2835 3366
rect 2927 3362 2931 3366
rect 2967 3362 2971 3366
rect 3063 3362 3067 3366
rect 3103 3362 3107 3366
rect 1863 3294 1867 3298
rect 1887 3294 1891 3298
rect 1927 3294 1931 3298
rect 1991 3294 1995 3298
rect 2047 3294 2051 3298
rect 2127 3294 2131 3298
rect 2175 3294 2179 3298
rect 2271 3294 2275 3298
rect 2311 3294 2315 3298
rect 1175 3286 1179 3290
rect 1191 3286 1195 3290
rect 1327 3286 1331 3290
rect 1335 3286 1339 3290
rect 1479 3286 1483 3290
rect 1487 3286 1491 3290
rect 1631 3286 1635 3290
rect 1823 3286 1827 3290
rect 583 3206 587 3210
rect 727 3206 731 3210
rect 751 3206 755 3210
rect 887 3206 891 3210
rect 903 3206 907 3210
rect 111 3126 115 3130
rect 135 3126 139 3130
rect 1947 3240 1951 3244
rect 2415 3294 2419 3298
rect 2455 3294 2459 3298
rect 2551 3294 2555 3298
rect 2599 3294 2603 3298
rect 2687 3294 2691 3298
rect 3575 3362 3579 3366
rect 2743 3294 2747 3298
rect 2823 3294 2827 3298
rect 2887 3294 2891 3298
rect 2359 3240 2363 3244
rect 1863 3218 1867 3222
rect 1935 3218 1939 3222
rect 2007 3218 2011 3222
rect 2055 3218 2059 3222
rect 2119 3218 2123 3222
rect 2183 3218 2187 3222
rect 2239 3218 2243 3222
rect 2319 3218 2323 3222
rect 2375 3218 2379 3222
rect 2463 3218 2467 3222
rect 2519 3218 2523 3222
rect 2607 3218 2611 3222
rect 1039 3206 1043 3210
rect 1055 3206 1059 3210
rect 1191 3206 1195 3210
rect 1199 3206 1203 3210
rect 1343 3206 1347 3210
rect 1351 3206 1355 3210
rect 1495 3206 1499 3210
rect 1823 3206 1827 3210
rect 1031 3192 1035 3196
rect 1279 3192 1283 3196
rect 2959 3294 2963 3298
rect 3031 3294 3035 3298
rect 3095 3294 3099 3298
rect 3183 3294 3187 3298
rect 3575 3294 3579 3298
rect 2663 3218 2667 3222
rect 2751 3218 2755 3222
rect 2815 3218 2819 3222
rect 2895 3218 2899 3222
rect 2967 3218 2971 3222
rect 3039 3218 3043 3222
rect 3119 3218 3123 3222
rect 3191 3218 3195 3222
rect 3279 3218 3283 3222
rect 3575 3218 3579 3222
rect 807 3144 811 3148
rect 1243 3144 1247 3148
rect 167 3126 171 3130
rect 263 3126 267 3130
rect 367 3126 371 3130
rect 399 3126 403 3130
rect 527 3126 531 3130
rect 551 3126 555 3130
rect 647 3126 651 3130
rect 719 3126 723 3130
rect 759 3126 763 3130
rect 863 3126 867 3130
rect 879 3126 883 3130
rect 967 3126 971 3130
rect 1031 3126 1035 3130
rect 1071 3126 1075 3130
rect 1175 3126 1179 3130
rect 1183 3126 1187 3130
rect 111 3058 115 3062
rect 143 3058 147 3062
rect 247 3058 251 3062
rect 271 3058 275 3062
rect 367 3058 371 3062
rect 407 3058 411 3062
rect 487 3058 491 3062
rect 535 3058 539 3062
rect 599 3058 603 3062
rect 111 2978 115 2982
rect 135 2978 139 2982
rect 239 2978 243 2982
rect 287 2978 291 2982
rect 359 2978 363 2982
rect 455 2978 459 2982
rect 479 2978 483 2982
rect 1863 3146 1867 3150
rect 1999 3146 2003 3150
rect 2055 3146 2059 3150
rect 2111 3146 2115 3150
rect 2207 3146 2211 3150
rect 2231 3146 2235 3150
rect 2359 3146 2363 3150
rect 2367 3146 2371 3150
rect 2511 3146 2515 3150
rect 1279 3126 1283 3130
rect 1343 3126 1347 3130
rect 1823 3126 1827 3130
rect 1863 3074 1867 3078
rect 1951 3074 1955 3078
rect 655 3058 659 3062
rect 703 3058 707 3062
rect 767 3058 771 3062
rect 799 3058 803 3062
rect 871 3058 875 3062
rect 895 3058 899 3062
rect 975 3058 979 3062
rect 991 3058 995 3062
rect 1079 3058 1083 3062
rect 1087 3058 1091 3062
rect 1183 3058 1187 3062
rect 1287 3058 1291 3062
rect 1823 3058 1827 3062
rect 951 3048 955 3052
rect 591 2978 595 2982
rect 623 2978 627 2982
rect 695 2978 699 2982
rect 783 2978 787 2982
rect 791 2978 795 2982
rect 887 2978 891 2982
rect 927 2978 931 2982
rect 111 2910 115 2914
rect 143 2910 147 2914
rect 295 2910 299 2914
rect 319 2910 323 2914
rect 475 2920 479 2924
rect 691 2920 695 2924
rect 983 2978 987 2982
rect 1251 3048 1255 3052
rect 2655 3146 2659 3150
rect 2791 3146 2795 3150
rect 2807 3146 2811 3150
rect 2919 3146 2923 3150
rect 2959 3146 2963 3150
rect 3039 3146 3043 3150
rect 3111 3146 3115 3150
rect 3159 3146 3163 3150
rect 3271 3146 3275 3150
rect 3383 3146 3387 3150
rect 3479 3146 3483 3150
rect 3575 3146 3579 3150
rect 2063 3074 2067 3078
rect 2079 3074 2083 3078
rect 2215 3074 2219 3078
rect 2367 3074 2371 3078
rect 2519 3074 2523 3078
rect 2527 3074 2531 3078
rect 2663 3074 2667 3078
rect 2679 3074 2683 3078
rect 2799 3074 2803 3078
rect 2831 3074 2835 3078
rect 2927 3074 2931 3078
rect 2975 3074 2979 3078
rect 3047 3074 3051 3078
rect 3111 3074 3115 3078
rect 1863 2994 1867 2998
rect 1887 2994 1891 2998
rect 1943 2994 1947 2998
rect 1975 2994 1979 2998
rect 2063 2994 2067 2998
rect 2071 2994 2075 2998
rect 2151 2994 2155 2998
rect 2207 2994 2211 2998
rect 2239 2994 2243 2998
rect 2351 2994 2355 2998
rect 2359 2994 2363 2998
rect 2463 2994 2467 2998
rect 2519 2994 2523 2998
rect 2575 2994 2579 2998
rect 1063 2978 1067 2982
rect 1079 2978 1083 2982
rect 1175 2978 1179 2982
rect 1191 2978 1195 2982
rect 1279 2978 1283 2982
rect 1311 2978 1315 2982
rect 1423 2978 1427 2982
rect 1527 2978 1531 2982
rect 1639 2978 1643 2982
rect 1727 2978 1731 2982
rect 1823 2978 1827 2982
rect 1119 2920 1123 2924
rect 463 2910 467 2914
rect 519 2910 523 2914
rect 631 2910 635 2914
rect 711 2910 715 2914
rect 791 2910 795 2914
rect 895 2910 899 2914
rect 935 2910 939 2914
rect 1071 2910 1075 2914
rect 1199 2910 1203 2914
rect 1239 2910 1243 2914
rect 1319 2910 1323 2914
rect 1399 2910 1403 2914
rect 111 2838 115 2842
rect 135 2838 139 2842
rect 159 2838 163 2842
rect 311 2838 315 2842
rect 319 2838 323 2842
rect 487 2838 491 2842
rect 511 2838 515 2842
rect 655 2838 659 2842
rect 703 2838 707 2842
rect 823 2838 827 2842
rect 887 2838 891 2842
rect 1119 2888 1123 2892
rect 1415 2920 1419 2924
rect 1863 2918 1867 2922
rect 2671 2994 2675 2998
rect 2687 2994 2691 2998
rect 2799 2994 2803 2998
rect 2823 2994 2827 2998
rect 3167 3074 3171 3078
rect 3239 3074 3243 3078
rect 3279 3074 3283 3078
rect 3375 3074 3379 3078
rect 3391 3074 3395 3078
rect 3487 3074 3491 3078
rect 3575 3074 3579 3078
rect 2903 2994 2907 2998
rect 2967 2994 2971 2998
rect 3007 2994 3011 2998
rect 3103 2994 3107 2998
rect 3199 2994 3203 2998
rect 3231 2994 3235 2998
rect 3295 2994 3299 2998
rect 3367 2994 3371 2998
rect 3391 2994 3395 2998
rect 3479 2994 3483 2998
rect 1431 2910 1435 2914
rect 1535 2910 1539 2914
rect 1551 2910 1555 2914
rect 1647 2910 1651 2914
rect 1711 2910 1715 2914
rect 1735 2910 1739 2914
rect 1823 2910 1827 2914
rect 1651 2896 1655 2900
rect 1895 2918 1899 2922
rect 1983 2918 1987 2922
rect 2071 2918 2075 2922
rect 2159 2918 2163 2922
rect 2247 2918 2251 2922
rect 2359 2918 2363 2922
rect 2471 2918 2475 2922
rect 2583 2918 2587 2922
rect 2695 2918 2699 2922
rect 2807 2918 2811 2922
rect 2895 2918 2899 2922
rect 2911 2918 2915 2922
rect 3575 2994 3579 2998
rect 3015 2918 3019 2922
rect 3111 2918 3115 2922
rect 3199 2918 3203 2922
rect 3207 2918 3211 2922
rect 3303 2918 3307 2922
rect 3399 2918 3403 2922
rect 3487 2918 3491 2922
rect 3575 2918 3579 2922
rect 975 2838 979 2842
rect 1063 2838 1067 2842
rect 1127 2838 1131 2842
rect 1231 2838 1235 2842
rect 1271 2838 1275 2842
rect 111 2762 115 2766
rect 167 2762 171 2766
rect 207 2762 211 2766
rect 327 2762 331 2766
rect 335 2762 339 2766
rect 471 2762 475 2766
rect 495 2762 499 2766
rect 995 2784 999 2788
rect 1863 2850 1867 2854
rect 2831 2850 2835 2854
rect 2887 2850 2891 2854
rect 2919 2850 2923 2854
rect 3007 2850 3011 2854
rect 3095 2850 3099 2854
rect 1391 2838 1395 2842
rect 1415 2838 1419 2842
rect 1543 2838 1547 2842
rect 1559 2838 1563 2842
rect 1703 2838 1707 2842
rect 1823 2838 1827 2842
rect 3191 2850 3195 2854
rect 3479 2850 3483 2854
rect 1483 2784 1487 2788
rect 1863 2782 1867 2786
rect 2671 2782 2675 2786
rect 2807 2782 2811 2786
rect 2839 2782 2843 2786
rect 607 2762 611 2766
rect 663 2762 667 2766
rect 751 2762 755 2766
rect 831 2762 835 2766
rect 887 2762 891 2766
rect 983 2762 987 2766
rect 1023 2762 1027 2766
rect 1135 2762 1139 2766
rect 1151 2762 1155 2766
rect 1279 2762 1283 2766
rect 1287 2762 1291 2766
rect 1423 2762 1427 2766
rect 1567 2762 1571 2766
rect 1823 2762 1827 2766
rect 111 2690 115 2694
rect 199 2690 203 2694
rect 215 2690 219 2694
rect 327 2690 331 2694
rect 335 2690 339 2694
rect 463 2690 467 2694
rect 583 2690 587 2694
rect 599 2690 603 2694
rect 2927 2782 2931 2786
rect 2967 2782 2971 2786
rect 3015 2782 3019 2786
rect 3103 2782 3107 2786
rect 3143 2782 3147 2786
rect 3327 2782 3331 2786
rect 3487 2782 3491 2786
rect 3575 2850 3579 2854
rect 3575 2782 3579 2786
rect 2851 2760 2855 2764
rect 3259 2760 3263 2764
rect 2735 2728 2739 2732
rect 3363 2728 3367 2732
rect 1863 2714 1867 2718
rect 703 2690 707 2694
rect 743 2690 747 2694
rect 823 2690 827 2694
rect 879 2690 883 2694
rect 935 2690 939 2694
rect 1015 2690 1019 2694
rect 1047 2690 1051 2694
rect 1143 2690 1147 2694
rect 1159 2690 1163 2694
rect 111 2618 115 2622
rect 223 2618 227 2622
rect 343 2618 347 2622
rect 471 2618 475 2622
rect 559 2618 563 2622
rect 591 2618 595 2622
rect 647 2618 651 2622
rect 711 2618 715 2622
rect 735 2618 739 2622
rect 111 2542 115 2546
rect 463 2542 467 2546
rect 843 2632 847 2636
rect 823 2618 827 2622
rect 831 2618 835 2622
rect 911 2618 915 2622
rect 943 2618 947 2622
rect 999 2618 1003 2622
rect 1055 2618 1059 2622
rect 1087 2618 1091 2622
rect 1887 2714 1891 2718
rect 1975 2714 1979 2718
rect 2063 2714 2067 2718
rect 2151 2714 2155 2718
rect 2239 2714 2243 2718
rect 2327 2714 2331 2718
rect 2415 2714 2419 2718
rect 2503 2714 2507 2718
rect 2591 2714 2595 2718
rect 2663 2714 2667 2718
rect 2679 2714 2683 2718
rect 2767 2714 2771 2718
rect 2799 2714 2803 2718
rect 2855 2714 2859 2718
rect 2943 2714 2947 2718
rect 2959 2714 2963 2718
rect 3031 2714 3035 2718
rect 3119 2714 3123 2718
rect 3135 2714 3139 2718
rect 3207 2714 3211 2718
rect 3295 2714 3299 2718
rect 3319 2714 3323 2718
rect 3391 2714 3395 2718
rect 3479 2714 3483 2718
rect 1271 2690 1275 2694
rect 1279 2690 1283 2694
rect 1415 2690 1419 2694
rect 1823 2690 1827 2694
rect 1227 2632 1231 2636
rect 1863 2626 1867 2630
rect 1895 2626 1899 2630
rect 1167 2618 1171 2622
rect 1175 2618 1179 2622
rect 1263 2618 1267 2622
rect 1279 2618 1283 2622
rect 1823 2618 1827 2622
rect 1983 2626 1987 2630
rect 2071 2626 2075 2630
rect 2159 2626 2163 2630
rect 2247 2626 2251 2630
rect 2279 2626 2283 2630
rect 2335 2626 2339 2630
rect 2415 2626 2419 2630
rect 2423 2626 2427 2630
rect 2511 2626 2515 2630
rect 1951 2592 1955 2596
rect 495 2542 499 2546
rect 551 2542 555 2546
rect 583 2542 587 2546
rect 639 2542 643 2546
rect 671 2542 675 2546
rect 111 2470 115 2474
rect 359 2470 363 2474
rect 471 2470 475 2474
rect 503 2470 507 2474
rect 415 2459 419 2460
rect 415 2456 419 2459
rect 727 2542 731 2546
rect 759 2542 763 2546
rect 815 2542 819 2546
rect 847 2542 851 2546
rect 903 2542 907 2546
rect 935 2542 939 2546
rect 591 2470 595 2474
rect 679 2470 683 2474
rect 719 2470 723 2474
rect 767 2470 771 2474
rect 1863 2558 1867 2562
rect 2103 2558 2107 2562
rect 2151 2558 2155 2562
rect 2199 2558 2203 2562
rect 2271 2558 2275 2562
rect 2311 2558 2315 2562
rect 2407 2558 2411 2562
rect 2431 2558 2435 2562
rect 991 2542 995 2546
rect 1023 2542 1027 2546
rect 1079 2542 1083 2546
rect 1111 2542 1115 2546
rect 1167 2542 1171 2546
rect 1199 2542 1203 2546
rect 1255 2542 1259 2546
rect 1287 2542 1291 2546
rect 1823 2542 1827 2546
rect 2551 2626 2555 2630
rect 2599 2626 2603 2630
rect 2687 2626 2691 2630
rect 2695 2626 2699 2630
rect 2775 2626 2779 2630
rect 2847 2626 2851 2630
rect 2863 2626 2867 2630
rect 2951 2626 2955 2630
rect 2999 2626 3003 2630
rect 3039 2626 3043 2630
rect 3127 2626 3131 2630
rect 3159 2626 3163 2630
rect 3215 2626 3219 2630
rect 3303 2626 3307 2630
rect 3399 2626 3403 2630
rect 2643 2595 2647 2596
rect 2643 2592 2647 2595
rect 2543 2558 2547 2562
rect 2559 2558 2563 2562
rect 2687 2558 2691 2562
rect 2695 2558 2699 2562
rect 2839 2558 2843 2562
rect 2847 2558 2851 2562
rect 2991 2558 2995 2562
rect 2999 2558 3003 2562
rect 979 2488 983 2492
rect 847 2470 851 2474
rect 855 2470 859 2474
rect 943 2470 947 2474
rect 967 2470 971 2474
rect 111 2398 115 2402
rect 135 2398 139 2402
rect 287 2398 291 2402
rect 351 2398 355 2402
rect 463 2398 467 2402
rect 471 2398 475 2402
rect 583 2398 587 2402
rect 663 2398 667 2402
rect 711 2398 715 2402
rect 787 2456 791 2460
rect 1267 2488 1271 2492
rect 1863 2486 1867 2490
rect 2087 2486 2091 2490
rect 2111 2486 2115 2490
rect 2183 2486 2187 2490
rect 2207 2486 2211 2490
rect 2287 2486 2291 2490
rect 2319 2486 2323 2490
rect 2407 2486 2411 2490
rect 2439 2486 2443 2490
rect 2543 2486 2547 2490
rect 2567 2486 2571 2490
rect 1031 2470 1035 2474
rect 1087 2470 1091 2474
rect 1119 2470 1123 2474
rect 1207 2470 1211 2474
rect 1295 2470 1299 2474
rect 1335 2470 1339 2474
rect 1463 2470 1467 2474
rect 1823 2470 1827 2474
rect 3151 2558 3155 2562
rect 3159 2558 3163 2562
rect 3327 2558 3331 2562
rect 3575 2714 3579 2718
rect 3487 2626 3491 2630
rect 3575 2626 3579 2630
rect 3479 2558 3483 2562
rect 3575 2558 3579 2562
rect 2703 2486 2707 2490
rect 2855 2486 2859 2490
rect 2887 2486 2891 2490
rect 3007 2486 3011 2490
rect 3087 2486 3091 2490
rect 3167 2486 3171 2490
rect 3295 2486 3299 2490
rect 3335 2486 3339 2490
rect 2099 2464 2103 2468
rect 2379 2464 2383 2468
rect 839 2398 843 2402
rect 847 2398 851 2402
rect 959 2398 963 2402
rect 1031 2398 1035 2402
rect 1079 2398 1083 2402
rect 1199 2398 1203 2402
rect 1207 2398 1211 2402
rect 1327 2398 1331 2402
rect 1375 2398 1379 2402
rect 111 2326 115 2330
rect 143 2326 147 2330
rect 295 2326 299 2330
rect 479 2326 483 2330
rect 671 2326 675 2330
rect 111 2250 115 2254
rect 135 2250 139 2254
rect 255 2250 259 2254
rect 287 2250 291 2254
rect 407 2250 411 2254
rect 471 2250 475 2254
rect 1095 2344 1099 2348
rect 1863 2414 1867 2418
rect 1951 2414 1955 2418
rect 2063 2414 2067 2418
rect 2079 2414 2083 2418
rect 2175 2414 2179 2418
rect 2183 2414 2187 2418
rect 2279 2414 2283 2418
rect 2311 2414 2315 2418
rect 1455 2398 1459 2402
rect 1543 2398 1547 2402
rect 1711 2398 1715 2402
rect 1823 2398 1827 2402
rect 3487 2486 3491 2490
rect 3575 2486 3579 2490
rect 2399 2414 2403 2418
rect 2447 2414 2451 2418
rect 2535 2414 2539 2418
rect 2591 2414 2595 2418
rect 2695 2414 2699 2418
rect 1403 2344 1407 2348
rect 855 2326 859 2330
rect 863 2326 867 2330
rect 1039 2326 1043 2330
rect 1055 2326 1059 2330
rect 1215 2326 1219 2330
rect 1231 2326 1235 2330
rect 1383 2326 1387 2330
rect 1407 2326 1411 2330
rect 1551 2326 1555 2330
rect 1583 2326 1587 2330
rect 1719 2326 1723 2330
rect 1735 2326 1739 2330
rect 1151 2296 1155 2300
rect 1339 2296 1343 2300
rect 1863 2338 1867 2342
rect 1895 2338 1899 2342
rect 1959 2338 1963 2342
rect 2007 2338 2011 2342
rect 1823 2326 1827 2330
rect 559 2250 563 2254
rect 663 2250 667 2254
rect 719 2250 723 2254
rect 855 2250 859 2254
rect 871 2250 875 2254
rect 1015 2250 1019 2254
rect 1047 2250 1051 2254
rect 1159 2250 1163 2254
rect 1223 2250 1227 2254
rect 1303 2250 1307 2254
rect 891 2192 895 2196
rect 111 2178 115 2182
rect 143 2178 147 2182
rect 215 2178 219 2182
rect 263 2178 267 2182
rect 311 2178 315 2182
rect 415 2178 419 2182
rect 519 2178 523 2182
rect 567 2178 571 2182
rect 623 2178 627 2182
rect 727 2178 731 2182
rect 831 2178 835 2182
rect 879 2178 883 2182
rect 943 2178 947 2182
rect 111 2102 115 2106
rect 207 2102 211 2106
rect 303 2102 307 2106
rect 319 2102 323 2106
rect 407 2102 411 2106
rect 423 2102 427 2106
rect 1023 2178 1027 2182
rect 1055 2178 1059 2182
rect 1099 2192 1103 2196
rect 1191 2192 1195 2196
rect 1863 2266 1867 2270
rect 1887 2266 1891 2270
rect 1399 2250 1403 2254
rect 1455 2250 1459 2254
rect 1575 2250 1579 2254
rect 1727 2250 1731 2254
rect 1823 2250 1827 2254
rect 2751 2414 2755 2418
rect 2879 2414 2883 2418
rect 2927 2414 2931 2418
rect 3079 2414 3083 2418
rect 3111 2414 3115 2418
rect 3287 2414 3291 2418
rect 3303 2414 3307 2418
rect 3479 2414 3483 2418
rect 3575 2414 3579 2418
rect 2071 2338 2075 2342
rect 2159 2338 2163 2342
rect 2191 2338 2195 2342
rect 2311 2338 2315 2342
rect 2319 2338 2323 2342
rect 2455 2338 2459 2342
rect 2463 2338 2467 2342
rect 2599 2338 2603 2342
rect 2615 2338 2619 2342
rect 2759 2338 2763 2342
rect 2775 2338 2779 2342
rect 2935 2338 2939 2342
rect 2943 2338 2947 2342
rect 3111 2338 3115 2342
rect 3119 2338 3123 2342
rect 3287 2338 3291 2342
rect 3311 2338 3315 2342
rect 3471 2338 3475 2342
rect 3487 2338 3491 2342
rect 3575 2338 3579 2342
rect 2047 2320 2051 2324
rect 2403 2320 2407 2324
rect 1999 2266 2003 2270
rect 2023 2266 2027 2270
rect 2151 2266 2155 2270
rect 2199 2266 2203 2270
rect 2303 2266 2307 2270
rect 2383 2266 2387 2270
rect 2455 2266 2459 2270
rect 2567 2266 2571 2270
rect 2607 2266 2611 2270
rect 2743 2266 2747 2270
rect 2767 2266 2771 2270
rect 1951 2248 1955 2252
rect 2479 2251 2483 2252
rect 2479 2248 2483 2251
rect 1399 2192 1403 2196
rect 1863 2194 1867 2198
rect 1895 2194 1899 2198
rect 1167 2178 1171 2182
rect 1311 2178 1315 2182
rect 1463 2178 1467 2182
rect 1823 2178 1827 2182
rect 2771 2208 2775 2212
rect 2911 2266 2915 2270
rect 2935 2266 2939 2270
rect 3079 2266 3083 2270
rect 3103 2266 3107 2270
rect 3239 2266 3243 2270
rect 3279 2266 3283 2270
rect 3407 2266 3411 2270
rect 3463 2266 3467 2270
rect 2031 2194 2035 2198
rect 2039 2194 2043 2198
rect 2207 2194 2211 2198
rect 2215 2194 2219 2198
rect 2391 2194 2395 2198
rect 2399 2194 2403 2198
rect 2575 2194 2579 2198
rect 2583 2194 2587 2198
rect 2751 2194 2755 2198
rect 2759 2194 2763 2198
rect 3147 2208 3151 2212
rect 2919 2194 2923 2198
rect 3071 2194 3075 2198
rect 3087 2194 3091 2198
rect 3215 2194 3219 2198
rect 3247 2194 3251 2198
rect 3359 2194 3363 2198
rect 3415 2194 3419 2198
rect 2007 2176 2011 2180
rect 2507 2176 2511 2180
rect 511 2102 515 2106
rect 527 2102 531 2106
rect 615 2102 619 2106
rect 631 2102 635 2106
rect 719 2102 723 2106
rect 735 2102 739 2106
rect 823 2102 827 2106
rect 831 2102 835 2106
rect 111 2026 115 2030
rect 215 2026 219 2030
rect 327 2026 331 2030
rect 391 2026 395 2030
rect 431 2026 435 2030
rect 535 2026 539 2030
rect 559 2026 563 2030
rect 639 2026 643 2030
rect 719 2026 723 2030
rect 743 2026 747 2030
rect 111 1950 115 1954
rect 135 1950 139 1954
rect 207 1950 211 1954
rect 311 1950 315 1954
rect 383 1950 387 1954
rect 519 1950 523 1954
rect 551 1950 555 1954
rect 1863 2122 1867 2126
rect 1887 2122 1891 2126
rect 2023 2122 2027 2126
rect 2031 2122 2035 2126
rect 2199 2122 2203 2126
rect 2207 2122 2211 2126
rect 2375 2122 2379 2126
rect 2391 2122 2395 2126
rect 2551 2122 2555 2126
rect 2575 2122 2579 2126
rect 2719 2122 2723 2126
rect 2751 2122 2755 2126
rect 2879 2122 2883 2126
rect 2911 2122 2915 2126
rect 3031 2122 3035 2126
rect 3063 2122 3067 2126
rect 3175 2122 3179 2126
rect 3207 2122 3211 2126
rect 3319 2122 3323 2126
rect 927 2102 931 2106
rect 935 2102 939 2106
rect 1031 2102 1035 2106
rect 1047 2102 1051 2106
rect 1135 2102 1139 2106
rect 1159 2102 1163 2106
rect 1239 2102 1243 2106
rect 1823 2102 1827 2106
rect 2039 2064 2043 2068
rect 1863 2046 1867 2050
rect 1895 2046 1899 2050
rect 2015 2046 2019 2050
rect 2031 2046 2035 2050
rect 2151 2046 2155 2050
rect 2207 2046 2211 2050
rect 839 2026 843 2030
rect 863 2026 867 2030
rect 935 2026 939 2030
rect 999 2026 1003 2030
rect 1039 2026 1043 2030
rect 1127 2026 1131 2030
rect 1143 2026 1147 2030
rect 1247 2026 1251 2030
rect 1367 2026 1371 2030
rect 1495 2026 1499 2030
rect 1823 2026 1827 2030
rect 2007 2027 2011 2028
rect 2007 2024 2011 2027
rect 2479 2064 2483 2068
rect 2295 2046 2299 2050
rect 2383 2046 2387 2050
rect 2439 2046 2443 2050
rect 2559 2046 2563 2050
rect 2591 2046 2595 2050
rect 2223 2024 2227 2028
rect 711 1950 715 1954
rect 719 1950 723 1954
rect 855 1950 859 1954
rect 911 1950 915 1954
rect 991 1950 995 1954
rect 1095 1950 1099 1954
rect 1119 1950 1123 1954
rect 111 1874 115 1878
rect 143 1874 147 1878
rect 311 1874 315 1878
rect 319 1874 323 1878
rect 511 1874 515 1878
rect 527 1874 531 1878
rect 703 1874 707 1878
rect 727 1874 731 1878
rect 887 1874 891 1878
rect 919 1874 923 1878
rect 111 1798 115 1802
rect 135 1798 139 1802
rect 263 1798 267 1802
rect 303 1798 307 1802
rect 415 1798 419 1802
rect 503 1798 507 1802
rect 567 1798 571 1802
rect 1863 1974 1867 1978
rect 1887 1974 1891 1978
rect 2007 1974 2011 1978
rect 2023 1974 2027 1978
rect 2111 1974 2115 1978
rect 2143 1974 2147 1978
rect 2199 1974 2203 1978
rect 2287 1974 2291 1978
rect 2383 1974 2387 1978
rect 2431 1974 2435 1978
rect 3351 2122 3355 2126
rect 3487 2194 3491 2198
rect 3575 2266 3579 2270
rect 3575 2194 3579 2198
rect 3471 2122 3475 2126
rect 3479 2122 3483 2126
rect 2727 2046 2731 2050
rect 2759 2046 2763 2050
rect 2887 2046 2891 2050
rect 2935 2046 2939 2050
rect 3039 2046 3043 2050
rect 3119 2046 3123 2050
rect 3183 2046 3187 2050
rect 3311 2046 3315 2050
rect 3327 2046 3331 2050
rect 2503 1974 2507 1978
rect 2583 1974 2587 1978
rect 2655 1974 2659 1978
rect 2751 1974 2755 1978
rect 2839 1974 2843 1978
rect 2927 1974 2931 1978
rect 3047 1974 3051 1978
rect 3111 1974 3115 1978
rect 3271 1974 3275 1978
rect 3303 1974 3307 1978
rect 1239 1950 1243 1954
rect 1263 1950 1267 1954
rect 1359 1950 1363 1954
rect 1423 1950 1427 1954
rect 1487 1950 1491 1954
rect 1583 1950 1587 1954
rect 1727 1950 1731 1954
rect 1823 1950 1827 1954
rect 1063 1874 1067 1878
rect 1103 1874 1107 1878
rect 1231 1874 1235 1878
rect 1271 1874 1275 1878
rect 1391 1874 1395 1878
rect 1431 1874 1435 1878
rect 1551 1874 1555 1878
rect 1591 1874 1595 1878
rect 1711 1874 1715 1878
rect 1135 1867 1139 1868
rect 1135 1864 1139 1867
rect 1299 1864 1303 1868
rect 1863 1898 1867 1902
rect 2031 1898 2035 1902
rect 1735 1874 1739 1878
rect 1823 1874 1827 1878
rect 2119 1898 2123 1902
rect 2175 1898 2179 1902
rect 2207 1898 2211 1902
rect 2263 1898 2267 1902
rect 2295 1898 2299 1902
rect 2351 1898 2355 1902
rect 2391 1898 2395 1902
rect 2439 1898 2443 1902
rect 2511 1898 2515 1902
rect 2527 1898 2531 1902
rect 2639 1898 2643 1902
rect 1863 1826 1867 1830
rect 695 1798 699 1802
rect 719 1798 723 1802
rect 863 1798 867 1802
rect 879 1798 883 1802
rect 1007 1798 1011 1802
rect 1055 1798 1059 1802
rect 1143 1798 1147 1802
rect 1223 1798 1227 1802
rect 1279 1798 1283 1802
rect 111 1730 115 1734
rect 143 1730 147 1734
rect 271 1730 275 1734
rect 279 1730 283 1734
rect 423 1730 427 1734
rect 431 1730 435 1734
rect 575 1730 579 1734
rect 583 1730 587 1734
rect 727 1730 731 1734
rect 2167 1826 2171 1830
rect 2255 1826 2259 1830
rect 2319 1826 2323 1830
rect 2343 1826 2347 1830
rect 2431 1826 2435 1830
rect 2439 1826 2443 1830
rect 2519 1826 2523 1830
rect 2663 1898 2667 1902
rect 2775 1898 2779 1902
rect 2847 1898 2851 1902
rect 2935 1898 2939 1902
rect 3055 1898 3059 1902
rect 3119 1898 3123 1902
rect 3279 1898 3283 1902
rect 3311 1898 3315 1902
rect 2559 1826 2563 1830
rect 2631 1826 2635 1830
rect 2679 1826 2683 1830
rect 2767 1826 2771 1830
rect 2799 1826 2803 1830
rect 2919 1826 2923 1830
rect 2927 1826 2931 1830
rect 3047 1826 3051 1830
rect 3111 1826 3115 1830
rect 3183 1826 3187 1830
rect 1383 1798 1387 1802
rect 1423 1798 1427 1802
rect 1543 1798 1547 1802
rect 1703 1798 1707 1802
rect 1823 1798 1827 1802
rect 863 1730 867 1734
rect 871 1730 875 1734
rect 991 1730 995 1734
rect 1015 1730 1019 1734
rect 1127 1730 1131 1734
rect 1151 1730 1155 1734
rect 1263 1730 1267 1734
rect 1287 1730 1291 1734
rect 1863 1750 1867 1754
rect 2295 1750 2299 1754
rect 2327 1750 2331 1754
rect 2407 1750 2411 1754
rect 2447 1750 2451 1754
rect 2527 1750 2531 1754
rect 2567 1750 2571 1754
rect 2655 1750 2659 1754
rect 2687 1750 2691 1754
rect 1431 1730 1435 1734
rect 1823 1730 1827 1734
rect 111 1662 115 1666
rect 135 1662 139 1666
rect 263 1662 267 1666
rect 271 1662 275 1666
rect 423 1662 427 1666
rect 575 1662 579 1666
rect 719 1662 723 1666
rect 727 1662 731 1666
rect 855 1662 859 1666
rect 871 1662 875 1666
rect 983 1662 987 1666
rect 1007 1662 1011 1666
rect 1119 1662 1123 1666
rect 1143 1662 1147 1666
rect 111 1590 115 1594
rect 143 1590 147 1594
rect 167 1590 171 1594
rect 443 1608 447 1612
rect 1023 1624 1027 1628
rect 643 1608 647 1612
rect 271 1590 275 1594
rect 335 1590 339 1594
rect 431 1590 435 1594
rect 511 1590 515 1594
rect 583 1590 587 1594
rect 679 1590 683 1594
rect 735 1590 739 1594
rect 891 1608 895 1612
rect 847 1590 851 1594
rect 879 1590 883 1594
rect 999 1590 1003 1594
rect 1015 1590 1019 1594
rect 111 1518 115 1522
rect 159 1518 163 1522
rect 215 1518 219 1522
rect 327 1518 331 1522
rect 391 1518 395 1522
rect 111 1446 115 1450
rect 223 1446 227 1450
rect 255 1446 259 1450
rect 503 1518 507 1522
rect 575 1518 579 1522
rect 671 1518 675 1522
rect 759 1518 763 1522
rect 839 1518 843 1522
rect 1863 1678 1867 1682
rect 2143 1678 2147 1682
rect 2247 1678 2251 1682
rect 2287 1678 2291 1682
rect 2819 1768 2823 1772
rect 3303 1826 3307 1830
rect 3319 1826 3323 1830
rect 3463 1826 3467 1830
rect 3479 2046 3483 2050
rect 3487 2046 3491 2050
rect 3575 2122 3579 2126
rect 3575 2046 3579 2050
rect 3479 1974 3483 1978
rect 3575 1974 3579 1978
rect 3487 1898 3491 1902
rect 3575 1898 3579 1902
rect 3479 1826 3483 1830
rect 3199 1768 3203 1772
rect 2775 1750 2779 1754
rect 2807 1750 2811 1754
rect 2895 1750 2899 1754
rect 2927 1750 2931 1754
rect 3015 1750 3019 1754
rect 3055 1750 3059 1754
rect 3135 1750 3139 1754
rect 3191 1750 3195 1754
rect 3255 1750 3259 1754
rect 3327 1750 3331 1754
rect 3383 1750 3387 1754
rect 1255 1662 1259 1666
rect 1279 1662 1283 1666
rect 1415 1662 1419 1666
rect 1823 1662 1827 1666
rect 2367 1678 2371 1682
rect 2399 1678 2403 1682
rect 2503 1678 2507 1682
rect 2519 1678 2523 1682
rect 2647 1678 2651 1682
rect 2767 1678 2771 1682
rect 2807 1678 2811 1682
rect 1347 1624 1351 1628
rect 1211 1608 1215 1612
rect 2887 1678 2891 1682
rect 2975 1678 2979 1682
rect 3007 1678 3011 1682
rect 3127 1678 3131 1682
rect 3143 1678 3147 1682
rect 3247 1678 3251 1682
rect 3319 1678 3323 1682
rect 1863 1610 1867 1614
rect 2007 1610 2011 1614
rect 2103 1610 2107 1614
rect 2151 1610 2155 1614
rect 2207 1610 2211 1614
rect 1151 1590 1155 1594
rect 1287 1590 1291 1594
rect 1295 1590 1299 1594
rect 1423 1590 1427 1594
rect 1439 1590 1443 1594
rect 1583 1590 1587 1594
rect 1823 1590 1827 1594
rect 2019 1603 2023 1604
rect 2019 1600 2023 1603
rect 935 1518 939 1522
rect 991 1518 995 1522
rect 1095 1518 1099 1522
rect 1143 1518 1147 1522
rect 1255 1518 1259 1522
rect 1287 1518 1291 1522
rect 1407 1518 1411 1522
rect 1431 1518 1435 1522
rect 383 1446 387 1450
rect 399 1446 403 1450
rect 519 1446 523 1450
rect 583 1446 587 1450
rect 671 1446 675 1450
rect 111 1378 115 1382
rect 247 1378 251 1382
rect 351 1378 355 1382
rect 375 1378 379 1382
rect 439 1378 443 1382
rect 511 1378 515 1382
rect 527 1378 531 1382
rect 367 1344 371 1348
rect 515 1347 519 1348
rect 515 1344 519 1347
rect 111 1310 115 1314
rect 359 1310 363 1314
rect 447 1310 451 1314
rect 455 1310 459 1314
rect 623 1378 627 1382
rect 663 1378 667 1382
rect 1115 1464 1119 1468
rect 2255 1610 2259 1614
rect 2327 1610 2331 1614
rect 2375 1610 2379 1614
rect 2463 1610 2467 1614
rect 2511 1610 2515 1614
rect 2607 1610 2611 1614
rect 2655 1610 2659 1614
rect 2767 1610 2771 1614
rect 2815 1610 2819 1614
rect 2943 1610 2947 1614
rect 2307 1600 2311 1604
rect 1863 1534 1867 1538
rect 1887 1534 1891 1538
rect 1975 1534 1979 1538
rect 1999 1534 2003 1538
rect 2095 1534 2099 1538
rect 2103 1534 2107 1538
rect 2199 1534 2203 1538
rect 2239 1534 2243 1538
rect 1559 1518 1563 1522
rect 1575 1518 1579 1522
rect 1711 1518 1715 1522
rect 1823 1518 1827 1522
rect 3375 1678 3379 1682
rect 2983 1610 2987 1614
rect 3127 1610 3131 1614
rect 3151 1610 3155 1614
rect 3319 1610 3323 1614
rect 3327 1610 3331 1614
rect 2319 1534 2323 1538
rect 2383 1534 2387 1538
rect 2455 1534 2459 1538
rect 2543 1534 2547 1538
rect 2599 1534 2603 1538
rect 2711 1534 2715 1538
rect 1519 1464 1523 1468
rect 1863 1462 1867 1466
rect 1895 1462 1899 1466
rect 767 1446 771 1450
rect 831 1446 835 1450
rect 943 1446 947 1450
rect 991 1446 995 1450
rect 1103 1446 1107 1450
rect 1143 1446 1147 1450
rect 1263 1446 1267 1450
rect 1295 1446 1299 1450
rect 1415 1446 1419 1450
rect 1447 1446 1451 1450
rect 1567 1446 1571 1450
rect 1599 1446 1603 1450
rect 1719 1446 1723 1450
rect 1735 1446 1739 1450
rect 1823 1446 1827 1450
rect 727 1378 731 1382
rect 823 1378 827 1382
rect 847 1378 851 1382
rect 983 1378 987 1382
rect 1127 1378 1131 1382
rect 1135 1378 1139 1382
rect 1279 1378 1283 1382
rect 1287 1378 1291 1382
rect 1431 1378 1435 1382
rect 1439 1378 1443 1382
rect 1591 1378 1595 1382
rect 2759 1534 2763 1538
rect 2879 1534 2883 1538
rect 2935 1534 2939 1538
rect 3055 1534 3059 1538
rect 3119 1534 3123 1538
rect 3239 1534 3243 1538
rect 3311 1534 3315 1538
rect 3431 1534 3435 1538
rect 1983 1462 1987 1466
rect 2023 1462 2027 1466
rect 2111 1462 2115 1466
rect 2175 1462 2179 1466
rect 2247 1462 2251 1466
rect 2319 1462 2323 1466
rect 2391 1462 2395 1466
rect 2463 1462 2467 1466
rect 2551 1462 2555 1466
rect 2615 1462 2619 1466
rect 2719 1462 2723 1466
rect 2767 1462 2771 1466
rect 1951 1432 1955 1436
rect 2243 1432 2247 1436
rect 1451 1328 1455 1332
rect 1727 1378 1731 1382
rect 1823 1378 1827 1382
rect 1863 1382 1867 1386
rect 1887 1382 1891 1386
rect 2015 1382 2019 1386
rect 2143 1382 2147 1386
rect 2167 1382 2171 1386
rect 2311 1382 2315 1386
rect 1871 1328 1875 1332
rect 2391 1382 2395 1386
rect 2455 1382 2459 1386
rect 2887 1462 2891 1466
rect 2935 1462 2939 1466
rect 3063 1462 3067 1466
rect 3103 1462 3107 1466
rect 3471 1750 3475 1754
rect 3487 1750 3491 1754
rect 3575 1826 3579 1830
rect 3575 1750 3579 1754
rect 3479 1678 3483 1682
rect 3575 1678 3579 1682
rect 3487 1610 3491 1614
rect 3575 1610 3579 1614
rect 3479 1534 3483 1538
rect 3575 1534 3579 1538
rect 3247 1462 3251 1466
rect 3279 1462 3283 1466
rect 3439 1462 3443 1466
rect 3463 1462 3467 1466
rect 3575 1462 3579 1466
rect 2607 1382 2611 1386
rect 2623 1382 2627 1386
rect 2759 1382 2763 1386
rect 2847 1382 2851 1386
rect 2927 1382 2931 1386
rect 3063 1382 3067 1386
rect 3095 1382 3099 1386
rect 3271 1382 3275 1386
rect 3455 1382 3459 1386
rect 3479 1382 3483 1386
rect 535 1310 539 1314
rect 543 1310 547 1314
rect 631 1310 635 1314
rect 719 1310 723 1314
rect 735 1310 739 1314
rect 831 1310 835 1314
rect 855 1310 859 1314
rect 967 1310 971 1314
rect 991 1310 995 1314
rect 1135 1310 1139 1314
rect 1287 1310 1291 1314
rect 1327 1310 1331 1314
rect 1439 1310 1443 1314
rect 1535 1310 1539 1314
rect 1599 1310 1603 1314
rect 1735 1310 1739 1314
rect 1823 1310 1827 1314
rect 1863 1314 1867 1318
rect 1895 1314 1899 1318
rect 111 1242 115 1246
rect 447 1242 451 1246
rect 535 1242 539 1246
rect 543 1242 547 1246
rect 623 1242 627 1246
rect 631 1242 635 1246
rect 711 1242 715 1246
rect 719 1242 723 1246
rect 807 1242 811 1246
rect 823 1242 827 1246
rect 895 1242 899 1246
rect 959 1242 963 1246
rect 991 1242 995 1246
rect 1095 1242 1099 1246
rect 1127 1242 1131 1246
rect 1207 1242 1211 1246
rect 1319 1242 1323 1246
rect 1335 1242 1339 1246
rect 1471 1242 1475 1246
rect 1527 1242 1531 1246
rect 1927 1314 1931 1318
rect 2111 1314 2115 1318
rect 2151 1314 2155 1318
rect 2287 1314 2291 1318
rect 2399 1314 2403 1318
rect 2455 1314 2459 1318
rect 2623 1314 2627 1318
rect 2631 1314 2635 1318
rect 1607 1242 1611 1246
rect 111 1166 115 1170
rect 359 1166 363 1170
rect 471 1166 475 1170
rect 551 1166 555 1170
rect 591 1166 595 1170
rect 639 1166 643 1170
rect 711 1166 715 1170
rect 727 1166 731 1170
rect 815 1166 819 1170
rect 831 1166 835 1170
rect 903 1166 907 1170
rect 951 1166 955 1170
rect 999 1166 1003 1170
rect 1727 1242 1731 1246
rect 1823 1242 1827 1246
rect 1863 1238 1867 1242
rect 1919 1238 1923 1242
rect 2103 1238 2107 1242
rect 2143 1238 2147 1242
rect 2791 1314 2795 1318
rect 2855 1314 2859 1318
rect 2959 1314 2963 1318
rect 2279 1238 2283 1242
rect 2319 1238 2323 1242
rect 2447 1238 2451 1242
rect 2487 1238 2491 1242
rect 1063 1166 1067 1170
rect 1103 1166 1107 1170
rect 1183 1166 1187 1170
rect 1215 1166 1219 1170
rect 1303 1166 1307 1170
rect 1343 1166 1347 1170
rect 1423 1166 1427 1170
rect 1479 1166 1483 1170
rect 1615 1166 1619 1170
rect 1735 1166 1739 1170
rect 2615 1238 2619 1242
rect 2655 1238 2659 1242
rect 2783 1238 2787 1242
rect 3575 1382 3579 1386
rect 3071 1314 3075 1318
rect 3135 1314 3139 1318
rect 3279 1314 3283 1318
rect 3319 1314 3323 1318
rect 2823 1238 2827 1242
rect 2951 1238 2955 1242
rect 2991 1238 2995 1242
rect 3127 1238 3131 1242
rect 3159 1238 3163 1242
rect 3311 1238 3315 1242
rect 3327 1238 3331 1242
rect 415 1136 419 1140
rect 779 1136 783 1140
rect 111 1094 115 1098
rect 143 1094 147 1098
rect 287 1094 291 1098
rect 351 1094 355 1098
rect 447 1094 451 1098
rect 463 1094 467 1098
rect 583 1094 587 1098
rect 615 1094 619 1098
rect 163 1040 167 1044
rect 111 1022 115 1026
rect 143 1022 147 1026
rect 151 1022 155 1026
rect 287 1022 291 1026
rect 295 1022 299 1026
rect 455 1022 459 1026
rect 471 1022 475 1026
rect 703 1094 707 1098
rect 783 1094 787 1098
rect 823 1094 827 1098
rect 943 1094 947 1098
rect 1055 1094 1059 1098
rect 1103 1094 1107 1098
rect 1175 1094 1179 1098
rect 1255 1094 1259 1098
rect 1295 1094 1299 1098
rect 1823 1166 1827 1170
rect 1863 1170 1867 1174
rect 1895 1170 1899 1174
rect 2007 1170 2011 1174
rect 2143 1170 2147 1174
rect 2151 1170 2155 1174
rect 2295 1170 2299 1174
rect 2327 1170 2331 1174
rect 1407 1094 1411 1098
rect 1415 1094 1419 1098
rect 1559 1094 1563 1098
rect 1823 1094 1827 1098
rect 1863 1094 1867 1098
rect 1887 1094 1891 1098
rect 1895 1094 1899 1098
rect 1999 1094 2003 1098
rect 2047 1094 2051 1098
rect 683 1040 687 1044
rect 959 1040 963 1044
rect 1475 1040 1479 1044
rect 623 1022 627 1026
rect 663 1022 667 1026
rect 791 1022 795 1026
rect 847 1022 851 1026
rect 951 1022 955 1026
rect 1031 1022 1035 1026
rect 1111 1022 1115 1026
rect 1207 1022 1211 1026
rect 1263 1022 1267 1026
rect 1375 1022 1379 1026
rect 1415 1022 1419 1026
rect 247 992 251 996
rect 771 992 775 996
rect 1543 1022 1547 1026
rect 1567 1022 1571 1026
rect 1711 1022 1715 1026
rect 1823 1022 1827 1026
rect 1863 1022 1867 1026
rect 1903 1022 1907 1026
rect 1975 1022 1979 1026
rect 1119 992 1123 996
rect 1459 992 1463 996
rect 111 950 115 954
rect 135 950 139 954
rect 279 950 283 954
rect 287 950 291 954
rect 463 950 467 954
rect 471 950 475 954
rect 655 950 659 954
rect 663 950 667 954
rect 839 950 843 954
rect 855 950 859 954
rect 1023 950 1027 954
rect 1047 950 1051 954
rect 1199 950 1203 954
rect 1223 950 1227 954
rect 1367 950 1371 954
rect 1399 950 1403 954
rect 1535 950 1539 954
rect 1575 950 1579 954
rect 1703 950 1707 954
rect 2135 1094 2139 1098
rect 2215 1094 2219 1098
rect 2287 1094 2291 1098
rect 2455 1170 2459 1174
rect 2495 1170 2499 1174
rect 2623 1170 2627 1174
rect 2663 1170 2667 1174
rect 2391 1094 2395 1098
rect 2447 1094 2451 1098
rect 2567 1094 2571 1098
rect 2055 1022 2059 1026
rect 2095 1022 2099 1026
rect 2223 1022 2227 1026
rect 2359 1022 2363 1026
rect 2399 1022 2403 1026
rect 2495 1022 2499 1026
rect 2791 1170 2795 1174
rect 2831 1170 2835 1174
rect 2967 1170 2971 1174
rect 2999 1170 3003 1174
rect 3143 1170 3147 1174
rect 2615 1094 2619 1098
rect 2735 1094 2739 1098
rect 2783 1094 2787 1098
rect 3167 1170 3171 1174
rect 3327 1170 3331 1174
rect 3335 1170 3339 1174
rect 2895 1094 2899 1098
rect 2959 1094 2963 1098
rect 3047 1094 3051 1098
rect 3135 1094 3139 1098
rect 3199 1094 3203 1098
rect 3319 1094 3323 1098
rect 3351 1094 3355 1098
rect 2575 1022 2579 1026
rect 2639 1022 2643 1026
rect 2743 1022 2747 1026
rect 2791 1022 2795 1026
rect 1727 950 1731 954
rect 1823 950 1827 954
rect 1863 950 1867 954
rect 1967 950 1971 954
rect 2087 950 2091 954
rect 2143 950 2147 954
rect 2215 950 2219 954
rect 2231 950 2235 954
rect 2319 950 2323 954
rect 2351 950 2355 954
rect 2407 950 2411 954
rect 2487 950 2491 954
rect 2503 950 2507 954
rect 303 896 307 900
rect 799 896 803 900
rect 111 878 115 882
rect 143 878 147 882
rect 287 878 291 882
rect 295 878 299 882
rect 471 878 475 882
rect 479 878 483 882
rect 655 878 659 882
rect 671 878 675 882
rect 839 878 843 882
rect 863 878 867 882
rect 1023 878 1027 882
rect 1055 878 1059 882
rect 1191 878 1195 882
rect 111 810 115 814
rect 135 810 139 814
rect 271 810 275 814
rect 279 810 283 814
rect 423 810 427 814
rect 463 810 467 814
rect 583 810 587 814
rect 647 810 651 814
rect 743 810 747 814
rect 2615 950 2619 954
rect 2631 950 2635 954
rect 3487 1314 3491 1318
rect 3575 1314 3579 1318
rect 3479 1238 3483 1242
rect 3575 1238 3579 1242
rect 3487 1170 3491 1174
rect 3575 1170 3579 1174
rect 3479 1094 3483 1098
rect 2903 1022 2907 1026
rect 2959 1022 2963 1026
rect 3055 1022 3059 1026
rect 3135 1022 3139 1026
rect 3207 1022 3211 1026
rect 3311 1022 3315 1026
rect 3359 1022 3363 1026
rect 3487 1022 3491 1026
rect 3575 1094 3579 1098
rect 2751 950 2755 954
rect 2783 950 2787 954
rect 2903 950 2907 954
rect 2951 950 2955 954
rect 3079 950 3083 954
rect 3127 950 3131 954
rect 3263 950 3267 954
rect 3303 950 3307 954
rect 3455 950 3459 954
rect 3479 950 3483 954
rect 3575 1022 3579 1026
rect 3575 950 3579 954
rect 1231 878 1235 882
rect 1359 878 1363 882
rect 1407 878 1411 882
rect 1527 878 1531 882
rect 1583 878 1587 882
rect 1695 878 1699 882
rect 1735 878 1739 882
rect 1823 878 1827 882
rect 1863 878 1867 882
rect 2103 878 2107 882
rect 2151 878 2155 882
rect 2191 878 2195 882
rect 2239 878 2243 882
rect 2279 878 2283 882
rect 2327 878 2331 882
rect 2367 878 2371 882
rect 2415 878 2419 882
rect 2455 878 2459 882
rect 2511 878 2515 882
rect 2567 878 2571 882
rect 2623 878 2627 882
rect 2703 878 2707 882
rect 2759 878 2763 882
rect 2871 878 2875 882
rect 2911 878 2915 882
rect 3055 878 3059 882
rect 3087 878 3091 882
rect 3255 878 3259 882
rect 3271 878 3275 882
rect 3463 878 3467 882
rect 3575 878 3579 882
rect 1207 856 1211 860
rect 1627 856 1631 860
rect 1087 824 1091 828
rect 1399 824 1403 828
rect 831 810 835 814
rect 895 810 899 814
rect 1015 810 1019 814
rect 1039 810 1043 814
rect 1183 810 1187 814
rect 1327 810 1331 814
rect 1351 810 1355 814
rect 1479 810 1483 814
rect 1519 810 1523 814
rect 1687 810 1691 814
rect 1823 810 1827 814
rect 1863 810 1867 814
rect 2095 810 2099 814
rect 2183 810 2187 814
rect 2199 810 2203 814
rect 2271 810 2275 814
rect 2287 810 2291 814
rect 155 792 159 796
rect 751 792 755 796
rect 371 752 375 756
rect 111 738 115 742
rect 143 738 147 742
rect 279 738 283 742
rect 359 738 363 742
rect 679 752 683 756
rect 431 738 435 742
rect 447 738 451 742
rect 543 738 547 742
rect 591 738 595 742
rect 639 738 643 742
rect 735 738 739 742
rect 751 738 755 742
rect 831 738 835 742
rect 903 738 907 742
rect 927 738 931 742
rect 1031 738 1035 742
rect 1047 738 1051 742
rect 1135 738 1139 742
rect 1191 738 1195 742
rect 1239 738 1243 742
rect 1335 738 1339 742
rect 1487 738 1491 742
rect 1823 738 1827 742
rect 1863 738 1867 742
rect 1943 738 1947 742
rect 2103 738 2107 742
rect 2207 738 2211 742
rect 2255 738 2259 742
rect 1023 728 1027 732
rect 1203 728 1207 732
rect 111 666 115 670
rect 351 666 355 670
rect 439 666 443 670
rect 479 666 483 670
rect 535 666 539 670
rect 567 666 571 670
rect 631 666 635 670
rect 655 666 659 670
rect 727 666 731 670
rect 743 666 747 670
rect 823 666 827 670
rect 831 666 835 670
rect 919 666 923 670
rect 1007 666 1011 670
rect 1023 666 1027 670
rect 1095 666 1099 670
rect 1127 666 1131 670
rect 1183 666 1187 670
rect 1231 666 1235 670
rect 1271 666 1275 670
rect 1823 666 1827 670
rect 1863 666 1867 670
rect 1887 666 1891 670
rect 1935 666 1939 670
rect 2023 666 2027 670
rect 2095 666 2099 670
rect 2359 810 2363 814
rect 2375 810 2379 814
rect 2447 810 2451 814
rect 2463 810 2467 814
rect 2551 810 2555 814
rect 2559 810 2563 814
rect 2655 810 2659 814
rect 2695 810 2699 814
rect 2783 810 2787 814
rect 2863 810 2867 814
rect 2935 810 2939 814
rect 3047 810 3051 814
rect 3111 810 3115 814
rect 2707 768 2711 772
rect 2295 738 2299 742
rect 2383 738 2387 742
rect 2407 738 2411 742
rect 2471 738 2475 742
rect 2551 738 2555 742
rect 2559 738 2563 742
rect 2675 752 2679 756
rect 2663 738 2667 742
rect 2695 738 2699 742
rect 3247 810 3251 814
rect 3295 810 3299 814
rect 3455 810 3459 814
rect 3479 810 3483 814
rect 3199 768 3203 772
rect 3139 752 3143 756
rect 2791 738 2795 742
rect 2839 738 2843 742
rect 2943 738 2947 742
rect 2983 738 2987 742
rect 3119 738 3123 742
rect 3135 738 3139 742
rect 3287 738 3291 742
rect 3303 738 3307 742
rect 3439 738 3443 742
rect 2199 666 2203 670
rect 2247 666 2251 670
rect 2383 666 2387 670
rect 2399 666 2403 670
rect 2543 666 2547 670
rect 2567 666 2571 670
rect 2687 666 2691 670
rect 2743 666 2747 670
rect 2831 666 2835 670
rect 2911 666 2915 670
rect 2975 666 2979 670
rect 3063 666 3067 670
rect 111 598 115 602
rect 487 598 491 602
rect 503 598 507 602
rect 575 598 579 602
rect 599 598 603 602
rect 663 598 667 602
rect 703 598 707 602
rect 751 598 755 602
rect 815 598 819 602
rect 839 598 843 602
rect 927 598 931 602
rect 935 598 939 602
rect 1015 598 1019 602
rect 1063 598 1067 602
rect 1103 598 1107 602
rect 1191 598 1195 602
rect 1279 598 1283 602
rect 1327 598 1331 602
rect 1471 598 1475 602
rect 1615 598 1619 602
rect 1735 598 1739 602
rect 1823 598 1827 602
rect 1863 598 1867 602
rect 1895 598 1899 602
rect 2031 598 2035 602
rect 2087 598 2091 602
rect 559 568 563 572
rect 771 568 775 572
rect 111 530 115 534
rect 159 530 163 534
rect 303 530 307 534
rect 463 530 467 534
rect 495 530 499 534
rect 591 530 595 534
rect 631 530 635 534
rect 695 530 699 534
rect 799 530 803 534
rect 807 530 811 534
rect 111 454 115 458
rect 143 454 147 458
rect 927 530 931 534
rect 959 530 963 534
rect 1055 530 1059 534
rect 1103 530 1107 534
rect 1183 530 1187 534
rect 1239 530 1243 534
rect 1319 530 1323 534
rect 1367 530 1371 534
rect 1463 530 1467 534
rect 1495 530 1499 534
rect 167 454 171 458
rect 271 454 275 458
rect 311 454 315 458
rect 439 454 443 458
rect 471 454 475 458
rect 615 454 619 458
rect 639 454 643 458
rect 791 454 795 458
rect 807 454 811 458
rect 967 454 971 458
rect 1111 454 1115 458
rect 1127 454 1131 458
rect 1247 454 1251 458
rect 1287 454 1291 458
rect 1375 454 1379 458
rect 1447 454 1451 458
rect 1607 530 1611 534
rect 1623 530 1627 534
rect 2207 598 2211 602
rect 2303 598 2307 602
rect 2391 598 2395 602
rect 2511 598 2515 602
rect 2575 598 2579 602
rect 2703 598 2707 602
rect 2763 608 2767 612
rect 3127 666 3131 670
rect 3207 666 3211 670
rect 3079 608 3083 612
rect 3279 666 3283 670
rect 3351 666 3355 670
rect 3431 666 3435 670
rect 2751 598 2755 602
rect 2879 598 2883 602
rect 2919 598 2923 602
rect 3039 598 3043 602
rect 3071 598 3075 602
rect 3199 598 3203 602
rect 3215 598 3219 602
rect 3351 598 3355 602
rect 3359 598 3363 602
rect 1727 530 1731 534
rect 1823 530 1827 534
rect 1863 522 1867 526
rect 1887 522 1891 526
rect 2079 522 2083 526
rect 2287 522 2291 526
rect 2295 522 2299 526
rect 2487 522 2491 526
rect 2503 522 2507 526
rect 2671 522 2675 526
rect 2695 522 2699 526
rect 2847 522 2851 526
rect 2871 522 2875 526
rect 3015 522 3019 526
rect 3031 522 3035 526
rect 3175 522 3179 526
rect 3191 522 3195 526
rect 3335 522 3339 526
rect 3343 522 3347 526
rect 2095 464 2099 468
rect 2419 464 2423 468
rect 2687 464 2691 468
rect 3083 464 3087 468
rect 3487 738 3491 742
rect 3575 810 3579 814
rect 3575 738 3579 742
rect 3479 666 3483 670
rect 3575 666 3579 670
rect 3487 598 3491 602
rect 3575 598 3579 602
rect 3479 522 3483 526
rect 3575 522 3579 526
rect 1503 454 1507 458
rect 1607 454 1611 458
rect 1631 454 1635 458
rect 1735 454 1739 458
rect 1823 454 1827 458
rect 1863 454 1867 458
rect 2087 454 2091 458
rect 2247 454 2251 458
rect 2295 454 2299 458
rect 2335 454 2339 458
rect 2431 454 2435 458
rect 2495 454 2499 458
rect 1239 432 1243 436
rect 1547 432 1551 436
rect 2303 443 2307 444
rect 2303 440 2307 443
rect 2527 454 2531 458
rect 2623 454 2627 458
rect 2679 454 2683 458
rect 2735 454 2739 458
rect 2855 454 2859 458
rect 2863 454 2867 458
rect 3007 454 3011 458
rect 3023 454 3027 458
rect 3167 454 3171 458
rect 3183 454 3187 458
rect 3335 454 3339 458
rect 3343 454 3347 458
rect 111 386 115 390
rect 135 386 139 390
rect 263 386 267 390
rect 431 386 435 390
rect 607 386 611 390
rect 783 386 787 390
rect 951 386 955 390
rect 959 386 963 390
rect 1111 386 1115 390
rect 1119 386 1123 390
rect 1271 386 1275 390
rect 1279 386 1283 390
rect 155 368 159 372
rect 683 368 687 372
rect 351 328 355 332
rect 111 314 115 318
rect 143 314 147 318
rect 263 314 267 318
rect 271 314 275 318
rect 691 328 695 332
rect 391 314 395 318
rect 439 314 443 318
rect 527 314 531 318
rect 615 314 619 318
rect 679 314 683 318
rect 791 314 795 318
rect 839 314 843 318
rect 959 314 963 318
rect 1007 314 1011 318
rect 1119 314 1123 318
rect 1175 314 1179 318
rect 1431 386 1435 390
rect 1439 386 1443 390
rect 1591 386 1595 390
rect 1599 386 1603 390
rect 1823 386 1827 390
rect 1863 386 1867 390
rect 2151 386 2155 390
rect 2239 386 2243 390
rect 2327 386 2331 390
rect 2415 386 2419 390
rect 2423 386 2427 390
rect 2503 386 2507 390
rect 2519 386 2523 390
rect 2595 440 2599 444
rect 3487 454 3491 458
rect 3575 454 3579 458
rect 2615 386 2619 390
rect 2727 386 2731 390
rect 2751 386 2755 390
rect 2855 386 2859 390
rect 2919 386 2923 390
rect 1279 314 1283 318
rect 1343 314 1347 318
rect 1439 314 1443 318
rect 1511 314 1515 318
rect 1599 314 1603 318
rect 1687 314 1691 318
rect 1823 314 1827 318
rect 1863 318 1867 322
rect 2023 318 2027 322
rect 2119 318 2123 322
rect 2159 318 2163 322
rect 111 242 115 246
rect 255 242 259 246
rect 383 242 387 246
rect 399 242 403 246
rect 503 242 507 246
rect 519 242 523 246
rect 615 242 619 246
rect 671 242 675 246
rect 735 242 739 246
rect 419 184 423 188
rect 831 242 835 246
rect 863 242 867 246
rect 991 242 995 246
rect 999 242 1003 246
rect 1119 242 1123 246
rect 1167 242 1171 246
rect 1247 242 1251 246
rect 1335 242 1339 246
rect 1375 242 1379 246
rect 811 184 815 188
rect 1863 250 1867 254
rect 1959 250 1963 254
rect 2015 250 2019 254
rect 1495 242 1499 246
rect 1503 242 1507 246
rect 1623 242 1627 246
rect 1679 242 1683 246
rect 1727 242 1731 246
rect 1823 242 1827 246
rect 2223 318 2227 322
rect 2247 318 2251 322
rect 2327 318 2331 322
rect 2335 318 2339 322
rect 2423 318 2427 322
rect 2431 318 2435 322
rect 2511 318 2515 322
rect 2535 318 2539 322
rect 2771 328 2775 332
rect 2999 386 3003 390
rect 3103 386 3107 390
rect 3159 386 3163 390
rect 3303 386 3307 390
rect 3327 386 3331 390
rect 3479 386 3483 390
rect 3575 386 3579 390
rect 3199 328 3203 332
rect 2623 318 2627 322
rect 2639 318 2643 322
rect 2743 318 2747 322
rect 2759 318 2763 322
rect 2855 318 2859 322
rect 2927 318 2931 322
rect 2967 318 2971 322
rect 3111 318 3115 322
rect 3311 318 3315 322
rect 3487 318 3491 322
rect 3575 318 3579 322
rect 2215 288 2219 292
rect 2399 288 2403 292
rect 2111 250 2115 254
rect 2175 250 2179 254
rect 2215 250 2219 254
rect 2319 250 2323 254
rect 2383 250 2387 254
rect 2423 250 2427 254
rect 2527 250 2531 254
rect 2583 250 2587 254
rect 2631 250 2635 254
rect 2735 250 2739 254
rect 2767 250 2771 254
rect 2847 250 2851 254
rect 111 154 115 158
rect 223 154 227 158
rect 311 154 315 158
rect 399 154 403 158
rect 407 154 411 158
rect 487 154 491 158
rect 511 154 515 158
rect 575 154 579 158
rect 623 154 627 158
rect 663 154 667 158
rect 743 154 747 158
rect 751 154 755 158
rect 839 154 843 158
rect 871 154 875 158
rect 927 154 931 158
rect 999 154 1003 158
rect 1015 154 1019 158
rect 1103 154 1107 158
rect 1127 154 1131 158
rect 1191 154 1195 158
rect 1255 154 1259 158
rect 1295 154 1299 158
rect 1383 154 1387 158
rect 1399 154 1403 158
rect 1503 154 1507 158
rect 1511 154 1515 158
rect 1631 154 1635 158
rect 1735 154 1739 158
rect 1823 154 1827 158
rect 1863 150 1867 154
rect 1895 150 1899 154
rect 1967 150 1971 154
rect 1983 150 1987 154
rect 2071 150 2075 154
rect 2159 150 2163 154
rect 2183 150 2187 154
rect 2271 150 2275 154
rect 2383 150 2387 154
rect 2391 150 2395 154
rect 2603 192 2607 196
rect 2619 160 2623 164
rect 2495 150 2499 154
rect 2591 150 2595 154
rect 2607 150 2611 154
rect 2951 250 2955 254
rect 2959 250 2963 254
rect 3127 250 3131 254
rect 3311 250 3315 254
rect 3479 250 3483 254
rect 3575 250 3579 254
rect 2923 192 2927 196
rect 3199 160 3203 164
rect 2719 150 2723 154
rect 2775 150 2779 154
rect 2823 150 2827 154
rect 2927 150 2931 154
rect 2959 150 2963 154
rect 3023 150 3027 154
rect 3119 150 3123 154
rect 3135 150 3139 154
rect 3215 150 3219 154
rect 3311 150 3315 154
rect 3319 150 3323 154
rect 3399 150 3403 154
rect 3487 150 3491 154
rect 3575 150 3579 154
rect 111 86 115 90
rect 215 86 219 90
rect 303 86 307 90
rect 391 86 395 90
rect 479 86 483 90
rect 567 86 571 90
rect 655 86 659 90
rect 743 86 747 90
rect 831 86 835 90
rect 919 86 923 90
rect 1007 86 1011 90
rect 1095 86 1099 90
rect 1183 86 1187 90
rect 1287 86 1291 90
rect 1391 86 1395 90
rect 1503 86 1507 90
rect 1623 86 1627 90
rect 1727 86 1731 90
rect 1823 86 1827 90
rect 1863 82 1867 86
rect 1887 82 1891 86
rect 1975 82 1979 86
rect 2063 82 2067 86
rect 2151 82 2155 86
rect 2263 82 2267 86
rect 2375 82 2379 86
rect 2487 82 2491 86
rect 2599 82 2603 86
rect 2711 82 2715 86
rect 2815 82 2819 86
rect 2919 82 2923 86
rect 3015 82 3019 86
rect 3111 82 3115 86
rect 3207 82 3211 86
rect 3303 82 3307 86
rect 3391 82 3395 86
rect 3479 82 3483 86
rect 3575 82 3579 86
<< m4 >>
rect 96 3645 97 3651
rect 103 3650 1847 3651
rect 103 3646 111 3650
rect 115 3646 143 3650
rect 147 3646 231 3650
rect 235 3646 319 3650
rect 323 3646 407 3650
rect 411 3646 495 3650
rect 499 3646 583 3650
rect 587 3646 671 3650
rect 675 3646 1823 3650
rect 1827 3646 1847 3650
rect 103 3645 1847 3646
rect 1853 3645 1854 3651
rect 84 3569 85 3575
rect 91 3574 1835 3575
rect 91 3570 111 3574
rect 115 3570 135 3574
rect 139 3570 223 3574
rect 227 3570 287 3574
rect 291 3570 311 3574
rect 315 3570 399 3574
rect 403 3570 463 3574
rect 467 3570 487 3574
rect 491 3570 575 3574
rect 579 3570 631 3574
rect 635 3570 663 3574
rect 667 3570 791 3574
rect 795 3570 935 3574
rect 939 3570 1071 3574
rect 1075 3570 1191 3574
rect 1195 3570 1311 3574
rect 1315 3570 1423 3574
rect 1427 3570 1527 3574
rect 1531 3570 1639 3574
rect 1643 3570 1727 3574
rect 1731 3570 1823 3574
rect 1827 3570 1835 3574
rect 91 3569 1835 3570
rect 1841 3569 1842 3575
rect 166 3556 172 3557
rect 650 3556 656 3557
rect 166 3552 167 3556
rect 171 3552 651 3556
rect 655 3552 656 3556
rect 166 3551 172 3552
rect 650 3551 656 3552
rect 158 3516 164 3517
rect 558 3516 564 3517
rect 158 3512 159 3516
rect 163 3512 559 3516
rect 563 3512 564 3516
rect 158 3511 164 3512
rect 558 3511 564 3512
rect 806 3516 812 3517
rect 1394 3516 1400 3517
rect 806 3512 807 3516
rect 811 3512 1395 3516
rect 1399 3512 1400 3516
rect 806 3511 812 3512
rect 1394 3511 1400 3512
rect 96 3501 97 3507
rect 103 3506 1847 3507
rect 103 3502 111 3506
rect 115 3502 143 3506
rect 147 3502 151 3506
rect 155 3502 295 3506
rect 299 3502 327 3506
rect 331 3502 471 3506
rect 475 3502 495 3506
rect 499 3502 639 3506
rect 643 3502 655 3506
rect 659 3502 799 3506
rect 803 3502 807 3506
rect 811 3502 943 3506
rect 947 3502 951 3506
rect 955 3502 1079 3506
rect 1083 3502 1087 3506
rect 1091 3502 1199 3506
rect 1203 3502 1207 3506
rect 1211 3502 1319 3506
rect 1323 3502 1431 3506
rect 1435 3502 1535 3506
rect 1539 3502 1647 3506
rect 1651 3502 1735 3506
rect 1739 3502 1823 3506
rect 1827 3502 1847 3506
rect 103 3501 1847 3502
rect 1853 3503 1854 3507
rect 1853 3502 3618 3503
rect 1853 3501 1863 3502
rect 1846 3498 1863 3501
rect 1867 3498 1895 3502
rect 1899 3498 1983 3502
rect 1987 3498 2071 3502
rect 2075 3498 2159 3502
rect 2163 3498 3575 3502
rect 3579 3498 3618 3502
rect 1846 3497 3618 3498
rect 878 3460 884 3461
rect 1646 3460 1652 3461
rect 878 3456 879 3460
rect 883 3456 1647 3460
rect 1651 3456 1652 3460
rect 878 3455 884 3456
rect 1646 3455 1652 3456
rect 84 3433 85 3439
rect 91 3438 1835 3439
rect 91 3434 111 3438
rect 115 3434 143 3438
rect 147 3434 215 3438
rect 219 3434 319 3438
rect 323 3434 431 3438
rect 435 3434 487 3438
rect 491 3434 639 3438
rect 643 3434 647 3438
rect 651 3434 799 3438
rect 803 3434 847 3438
rect 851 3434 943 3438
rect 947 3434 1039 3438
rect 1043 3434 1079 3438
rect 1083 3434 1199 3438
rect 1203 3434 1223 3438
rect 1227 3434 1311 3438
rect 1315 3434 1399 3438
rect 1403 3434 1423 3438
rect 1427 3434 1527 3438
rect 1531 3434 1567 3438
rect 1571 3434 1639 3438
rect 1643 3434 1727 3438
rect 1731 3434 1823 3438
rect 1827 3434 1835 3438
rect 91 3433 1835 3434
rect 1841 3435 1842 3439
rect 1841 3434 3606 3435
rect 1841 3433 1863 3434
rect 1834 3430 1863 3433
rect 1867 3430 1887 3434
rect 1891 3430 1975 3434
rect 1979 3430 1991 3434
rect 1995 3430 2063 3434
rect 2067 3430 2119 3434
rect 2123 3430 2151 3434
rect 2155 3430 2255 3434
rect 2259 3430 2391 3434
rect 2395 3430 2527 3434
rect 2531 3430 2655 3434
rect 2659 3430 2783 3434
rect 2787 3430 2919 3434
rect 2923 3430 3055 3434
rect 3059 3430 3575 3434
rect 3579 3430 3606 3434
rect 1834 3429 3606 3430
rect 234 3380 240 3381
rect 562 3380 568 3381
rect 234 3376 235 3380
rect 239 3376 563 3380
rect 567 3376 568 3380
rect 234 3375 240 3376
rect 562 3375 568 3376
rect 1906 3380 1912 3381
rect 2322 3380 2328 3381
rect 1906 3376 1907 3380
rect 1911 3376 2323 3380
rect 2327 3376 2328 3380
rect 1906 3375 1912 3376
rect 2322 3375 2328 3376
rect 1206 3372 1212 3373
rect 1582 3372 1588 3373
rect 1206 3368 1207 3372
rect 1211 3368 1583 3372
rect 1587 3368 1588 3372
rect 1206 3367 1212 3368
rect 1582 3367 1588 3368
rect 1846 3366 3618 3367
rect 1846 3363 1863 3366
rect 96 3357 97 3363
rect 103 3362 1847 3363
rect 103 3358 111 3362
rect 115 3358 223 3362
rect 227 3358 239 3362
rect 243 3358 383 3362
rect 387 3358 439 3362
rect 443 3358 543 3362
rect 547 3358 647 3362
rect 651 3358 711 3362
rect 715 3358 855 3362
rect 859 3358 871 3362
rect 875 3358 1031 3362
rect 1035 3358 1047 3362
rect 1051 3358 1183 3362
rect 1187 3358 1231 3362
rect 1235 3358 1335 3362
rect 1339 3358 1407 3362
rect 1411 3358 1487 3362
rect 1491 3358 1575 3362
rect 1579 3358 1639 3362
rect 1643 3358 1735 3362
rect 1739 3358 1823 3362
rect 1827 3358 1847 3362
rect 103 3357 1847 3358
rect 1853 3362 1863 3363
rect 1867 3362 1895 3366
rect 1899 3362 1999 3366
rect 2003 3362 2127 3366
rect 2131 3362 2135 3366
rect 2139 3362 2263 3366
rect 2267 3362 2279 3366
rect 2283 3362 2399 3366
rect 2403 3362 2423 3366
rect 2427 3362 2535 3366
rect 2539 3362 2559 3366
rect 2563 3362 2663 3366
rect 2667 3362 2695 3366
rect 2699 3362 2791 3366
rect 2795 3362 2831 3366
rect 2835 3362 2927 3366
rect 2931 3362 2967 3366
rect 2971 3362 3063 3366
rect 3067 3362 3103 3366
rect 3107 3362 3575 3366
rect 3579 3362 3618 3366
rect 1853 3361 3618 3362
rect 1853 3357 1854 3361
rect 1834 3293 1835 3299
rect 1841 3298 3599 3299
rect 1841 3294 1863 3298
rect 1867 3294 1887 3298
rect 1891 3294 1927 3298
rect 1931 3294 1991 3298
rect 1995 3294 2047 3298
rect 2051 3294 2127 3298
rect 2131 3294 2175 3298
rect 2179 3294 2271 3298
rect 2275 3294 2311 3298
rect 2315 3294 2415 3298
rect 2419 3294 2455 3298
rect 2459 3294 2551 3298
rect 2555 3294 2599 3298
rect 2603 3294 2687 3298
rect 2691 3294 2743 3298
rect 2747 3294 2823 3298
rect 2827 3294 2887 3298
rect 2891 3294 2959 3298
rect 2963 3294 3031 3298
rect 3035 3294 3095 3298
rect 3099 3294 3183 3298
rect 3187 3294 3575 3298
rect 3579 3294 3599 3298
rect 1841 3293 3599 3294
rect 3605 3293 3606 3299
rect 1834 3291 1842 3293
rect 84 3285 85 3291
rect 91 3290 1835 3291
rect 91 3286 111 3290
rect 115 3286 231 3290
rect 235 3286 239 3290
rect 243 3286 375 3290
rect 379 3286 407 3290
rect 411 3286 535 3290
rect 539 3286 575 3290
rect 579 3286 703 3290
rect 707 3286 743 3290
rect 747 3286 863 3290
rect 867 3286 895 3290
rect 899 3286 1023 3290
rect 1027 3286 1047 3290
rect 1051 3286 1175 3290
rect 1179 3286 1191 3290
rect 1195 3286 1327 3290
rect 1331 3286 1335 3290
rect 1339 3286 1479 3290
rect 1483 3286 1487 3290
rect 1491 3286 1631 3290
rect 1635 3286 1823 3290
rect 1827 3286 1835 3290
rect 91 3285 1835 3286
rect 1841 3285 1842 3291
rect 1946 3244 1952 3245
rect 2358 3244 2364 3245
rect 1946 3240 1947 3244
rect 1951 3240 2359 3244
rect 2363 3240 2364 3244
rect 1946 3239 1952 3240
rect 2358 3239 2364 3240
rect 258 3236 264 3237
rect 498 3236 504 3237
rect 258 3232 259 3236
rect 263 3232 499 3236
rect 503 3232 504 3236
rect 258 3231 264 3232
rect 498 3231 504 3232
rect 1846 3217 1847 3223
rect 1853 3222 3611 3223
rect 1853 3218 1863 3222
rect 1867 3218 1935 3222
rect 1939 3218 2007 3222
rect 2011 3218 2055 3222
rect 2059 3218 2119 3222
rect 2123 3218 2183 3222
rect 2187 3218 2239 3222
rect 2243 3218 2319 3222
rect 2323 3218 2375 3222
rect 2379 3218 2463 3222
rect 2467 3218 2519 3222
rect 2523 3218 2607 3222
rect 2611 3218 2663 3222
rect 2667 3218 2751 3222
rect 2755 3218 2815 3222
rect 2819 3218 2895 3222
rect 2899 3218 2967 3222
rect 2971 3218 3039 3222
rect 3043 3218 3119 3222
rect 3123 3218 3191 3222
rect 3195 3218 3279 3222
rect 3283 3218 3575 3222
rect 3579 3218 3611 3222
rect 1853 3217 3611 3218
rect 3617 3217 3618 3223
rect 96 3205 97 3211
rect 103 3210 1847 3211
rect 103 3206 111 3210
rect 115 3206 175 3210
rect 179 3206 247 3210
rect 251 3206 375 3210
rect 379 3206 415 3210
rect 419 3206 559 3210
rect 563 3206 583 3210
rect 587 3206 727 3210
rect 731 3206 751 3210
rect 755 3206 887 3210
rect 891 3206 903 3210
rect 907 3206 1039 3210
rect 1043 3206 1055 3210
rect 1059 3206 1191 3210
rect 1195 3206 1199 3210
rect 1203 3206 1343 3210
rect 1347 3206 1351 3210
rect 1355 3206 1495 3210
rect 1499 3206 1823 3210
rect 1827 3206 1847 3210
rect 103 3205 1847 3206
rect 1853 3205 1854 3211
rect 1030 3196 1036 3197
rect 1278 3196 1284 3197
rect 1030 3192 1031 3196
rect 1035 3192 1279 3196
rect 1283 3192 1284 3196
rect 1030 3191 1036 3192
rect 1278 3191 1284 3192
rect 806 3148 812 3149
rect 1242 3148 1248 3149
rect 806 3144 807 3148
rect 811 3144 1243 3148
rect 1247 3144 1248 3148
rect 1834 3145 1835 3151
rect 1841 3150 3599 3151
rect 1841 3146 1863 3150
rect 1867 3146 1999 3150
rect 2003 3146 2055 3150
rect 2059 3146 2111 3150
rect 2115 3146 2207 3150
rect 2211 3146 2231 3150
rect 2235 3146 2359 3150
rect 2363 3146 2367 3150
rect 2371 3146 2511 3150
rect 2515 3146 2655 3150
rect 2659 3146 2791 3150
rect 2795 3146 2807 3150
rect 2811 3146 2919 3150
rect 2923 3146 2959 3150
rect 2963 3146 3039 3150
rect 3043 3146 3111 3150
rect 3115 3146 3159 3150
rect 3163 3146 3271 3150
rect 3275 3146 3383 3150
rect 3387 3146 3479 3150
rect 3483 3146 3575 3150
rect 3579 3146 3599 3150
rect 1841 3145 3599 3146
rect 3605 3145 3606 3151
rect 806 3143 812 3144
rect 1242 3143 1248 3144
rect 84 3125 85 3131
rect 91 3130 1835 3131
rect 91 3126 111 3130
rect 115 3126 135 3130
rect 139 3126 167 3130
rect 171 3126 263 3130
rect 267 3126 367 3130
rect 371 3126 399 3130
rect 403 3126 527 3130
rect 531 3126 551 3130
rect 555 3126 647 3130
rect 651 3126 719 3130
rect 723 3126 759 3130
rect 763 3126 863 3130
rect 867 3126 879 3130
rect 883 3126 967 3130
rect 971 3126 1031 3130
rect 1035 3126 1071 3130
rect 1075 3126 1175 3130
rect 1179 3126 1183 3130
rect 1187 3126 1279 3130
rect 1283 3126 1343 3130
rect 1347 3126 1823 3130
rect 1827 3126 1835 3130
rect 91 3125 1835 3126
rect 1841 3125 1842 3131
rect 1846 3073 1847 3079
rect 1853 3078 3611 3079
rect 1853 3074 1863 3078
rect 1867 3074 1951 3078
rect 1955 3074 2063 3078
rect 2067 3074 2079 3078
rect 2083 3074 2215 3078
rect 2219 3074 2367 3078
rect 2371 3074 2519 3078
rect 2523 3074 2527 3078
rect 2531 3074 2663 3078
rect 2667 3074 2679 3078
rect 2683 3074 2799 3078
rect 2803 3074 2831 3078
rect 2835 3074 2927 3078
rect 2931 3074 2975 3078
rect 2979 3074 3047 3078
rect 3051 3074 3111 3078
rect 3115 3074 3167 3078
rect 3171 3074 3239 3078
rect 3243 3074 3279 3078
rect 3283 3074 3375 3078
rect 3379 3074 3391 3078
rect 3395 3074 3487 3078
rect 3491 3074 3575 3078
rect 3579 3074 3611 3078
rect 1853 3073 3611 3074
rect 3617 3073 3618 3079
rect 96 3057 97 3063
rect 103 3062 1847 3063
rect 103 3058 111 3062
rect 115 3058 143 3062
rect 147 3058 247 3062
rect 251 3058 271 3062
rect 275 3058 367 3062
rect 371 3058 407 3062
rect 411 3058 487 3062
rect 491 3058 535 3062
rect 539 3058 599 3062
rect 603 3058 655 3062
rect 659 3058 703 3062
rect 707 3058 767 3062
rect 771 3058 799 3062
rect 803 3058 871 3062
rect 875 3058 895 3062
rect 899 3058 975 3062
rect 979 3058 991 3062
rect 995 3058 1079 3062
rect 1083 3058 1087 3062
rect 1091 3058 1183 3062
rect 1187 3058 1287 3062
rect 1291 3058 1823 3062
rect 1827 3058 1847 3062
rect 103 3057 1847 3058
rect 1853 3057 1854 3063
rect 950 3052 956 3053
rect 1250 3052 1256 3053
rect 950 3048 951 3052
rect 955 3048 1251 3052
rect 1255 3048 1256 3052
rect 950 3047 956 3048
rect 1250 3047 1256 3048
rect 1834 2993 1835 2999
rect 1841 2998 3599 2999
rect 1841 2994 1863 2998
rect 1867 2994 1887 2998
rect 1891 2994 1943 2998
rect 1947 2994 1975 2998
rect 1979 2994 2063 2998
rect 2067 2994 2071 2998
rect 2075 2994 2151 2998
rect 2155 2994 2207 2998
rect 2211 2994 2239 2998
rect 2243 2994 2351 2998
rect 2355 2994 2359 2998
rect 2363 2994 2463 2998
rect 2467 2994 2519 2998
rect 2523 2994 2575 2998
rect 2579 2994 2671 2998
rect 2675 2994 2687 2998
rect 2691 2994 2799 2998
rect 2803 2994 2823 2998
rect 2827 2994 2903 2998
rect 2907 2994 2967 2998
rect 2971 2994 3007 2998
rect 3011 2994 3103 2998
rect 3107 2994 3199 2998
rect 3203 2994 3231 2998
rect 3235 2994 3295 2998
rect 3299 2994 3367 2998
rect 3371 2994 3391 2998
rect 3395 2994 3479 2998
rect 3483 2994 3575 2998
rect 3579 2994 3599 2998
rect 1841 2993 3599 2994
rect 3605 2993 3606 2999
rect 84 2977 85 2983
rect 91 2982 1835 2983
rect 91 2978 111 2982
rect 115 2978 135 2982
rect 139 2978 239 2982
rect 243 2978 287 2982
rect 291 2978 359 2982
rect 363 2978 455 2982
rect 459 2978 479 2982
rect 483 2978 591 2982
rect 595 2978 623 2982
rect 627 2978 695 2982
rect 699 2978 783 2982
rect 787 2978 791 2982
rect 795 2978 887 2982
rect 891 2978 927 2982
rect 931 2978 983 2982
rect 987 2978 1063 2982
rect 1067 2978 1079 2982
rect 1083 2978 1175 2982
rect 1179 2978 1191 2982
rect 1195 2978 1279 2982
rect 1283 2978 1311 2982
rect 1315 2978 1423 2982
rect 1427 2978 1527 2982
rect 1531 2978 1639 2982
rect 1643 2978 1727 2982
rect 1731 2978 1823 2982
rect 1827 2978 1835 2982
rect 91 2977 1835 2978
rect 1841 2977 1842 2983
rect 474 2924 480 2925
rect 690 2924 696 2925
rect 474 2920 475 2924
rect 479 2920 691 2924
rect 695 2920 696 2924
rect 474 2919 480 2920
rect 690 2919 696 2920
rect 1118 2924 1124 2925
rect 1414 2924 1420 2925
rect 1118 2920 1119 2924
rect 1123 2920 1415 2924
rect 1419 2920 1420 2924
rect 1118 2919 1124 2920
rect 1414 2919 1420 2920
rect 1846 2917 1847 2923
rect 1853 2922 3611 2923
rect 1853 2918 1863 2922
rect 1867 2918 1895 2922
rect 1899 2918 1983 2922
rect 1987 2918 2071 2922
rect 2075 2918 2159 2922
rect 2163 2918 2247 2922
rect 2251 2918 2359 2922
rect 2363 2918 2471 2922
rect 2475 2918 2583 2922
rect 2587 2918 2695 2922
rect 2699 2918 2807 2922
rect 2811 2918 2895 2922
rect 2899 2918 2911 2922
rect 2915 2918 3015 2922
rect 3019 2918 3111 2922
rect 3115 2918 3199 2922
rect 3203 2918 3207 2922
rect 3211 2918 3303 2922
rect 3307 2918 3399 2922
rect 3403 2918 3487 2922
rect 3491 2918 3575 2922
rect 3579 2918 3611 2922
rect 1853 2917 3611 2918
rect 3617 2917 3618 2923
rect 1846 2915 1854 2917
rect 96 2909 97 2915
rect 103 2914 1847 2915
rect 103 2910 111 2914
rect 115 2910 143 2914
rect 147 2910 295 2914
rect 299 2910 319 2914
rect 323 2910 463 2914
rect 467 2910 519 2914
rect 523 2910 631 2914
rect 635 2910 711 2914
rect 715 2910 791 2914
rect 795 2910 895 2914
rect 899 2910 935 2914
rect 939 2910 1071 2914
rect 1075 2910 1199 2914
rect 1203 2910 1239 2914
rect 1243 2910 1319 2914
rect 1323 2910 1399 2914
rect 1403 2910 1431 2914
rect 1435 2910 1535 2914
rect 1539 2910 1551 2914
rect 1555 2910 1647 2914
rect 1651 2910 1711 2914
rect 1715 2910 1735 2914
rect 1739 2910 1823 2914
rect 1827 2910 1847 2914
rect 103 2909 1847 2910
rect 1853 2909 1854 2915
rect 1650 2900 1656 2901
rect 1158 2896 1651 2900
rect 1655 2896 1656 2900
rect 1118 2892 1124 2893
rect 1158 2892 1162 2896
rect 1650 2895 1656 2896
rect 1118 2888 1119 2892
rect 1123 2888 1162 2892
rect 1118 2887 1124 2888
rect 1834 2849 1835 2855
rect 1841 2854 3599 2855
rect 1841 2850 1863 2854
rect 1867 2850 2831 2854
rect 2835 2850 2887 2854
rect 2891 2850 2919 2854
rect 2923 2850 3007 2854
rect 3011 2850 3095 2854
rect 3099 2850 3191 2854
rect 3195 2850 3479 2854
rect 3483 2850 3575 2854
rect 3579 2850 3599 2854
rect 1841 2849 3599 2850
rect 3605 2849 3606 2855
rect 84 2837 85 2843
rect 91 2842 1835 2843
rect 91 2838 111 2842
rect 115 2838 135 2842
rect 139 2838 159 2842
rect 163 2838 311 2842
rect 315 2838 319 2842
rect 323 2838 487 2842
rect 491 2838 511 2842
rect 515 2838 655 2842
rect 659 2838 703 2842
rect 707 2838 823 2842
rect 827 2838 887 2842
rect 891 2838 975 2842
rect 979 2838 1063 2842
rect 1067 2838 1127 2842
rect 1131 2838 1231 2842
rect 1235 2838 1271 2842
rect 1275 2838 1391 2842
rect 1395 2838 1415 2842
rect 1419 2838 1543 2842
rect 1547 2838 1559 2842
rect 1563 2838 1703 2842
rect 1707 2838 1823 2842
rect 1827 2838 1835 2842
rect 91 2837 1835 2838
rect 1841 2837 1842 2843
rect 994 2788 1000 2789
rect 1482 2788 1488 2789
rect 994 2784 995 2788
rect 999 2784 1483 2788
rect 1487 2784 1488 2788
rect 994 2783 1000 2784
rect 1482 2783 1488 2784
rect 1846 2781 1847 2787
rect 1853 2786 3611 2787
rect 1853 2782 1863 2786
rect 1867 2782 2671 2786
rect 2675 2782 2807 2786
rect 2811 2782 2839 2786
rect 2843 2782 2927 2786
rect 2931 2782 2967 2786
rect 2971 2782 3015 2786
rect 3019 2782 3103 2786
rect 3107 2782 3143 2786
rect 3147 2782 3327 2786
rect 3331 2782 3487 2786
rect 3491 2782 3575 2786
rect 3579 2782 3611 2786
rect 1853 2781 3611 2782
rect 3617 2781 3618 2787
rect 96 2761 97 2767
rect 103 2766 1847 2767
rect 103 2762 111 2766
rect 115 2762 167 2766
rect 171 2762 207 2766
rect 211 2762 327 2766
rect 331 2762 335 2766
rect 339 2762 471 2766
rect 475 2762 495 2766
rect 499 2762 607 2766
rect 611 2762 663 2766
rect 667 2762 751 2766
rect 755 2762 831 2766
rect 835 2762 887 2766
rect 891 2762 983 2766
rect 987 2762 1023 2766
rect 1027 2762 1135 2766
rect 1139 2762 1151 2766
rect 1155 2762 1279 2766
rect 1283 2762 1287 2766
rect 1291 2762 1423 2766
rect 1427 2762 1567 2766
rect 1571 2762 1823 2766
rect 1827 2762 1847 2766
rect 103 2761 1847 2762
rect 1853 2761 1854 2767
rect 2850 2764 2856 2765
rect 3258 2764 3264 2765
rect 2850 2760 2851 2764
rect 2855 2760 3259 2764
rect 3263 2760 3264 2764
rect 2850 2759 2856 2760
rect 3258 2759 3264 2760
rect 2734 2732 2740 2733
rect 3362 2732 3368 2733
rect 2734 2728 2735 2732
rect 2739 2728 3363 2732
rect 3367 2728 3368 2732
rect 2734 2727 2740 2728
rect 3362 2727 3368 2728
rect 1834 2713 1835 2719
rect 1841 2718 3599 2719
rect 1841 2714 1863 2718
rect 1867 2714 1887 2718
rect 1891 2714 1975 2718
rect 1979 2714 2063 2718
rect 2067 2714 2151 2718
rect 2155 2714 2239 2718
rect 2243 2714 2327 2718
rect 2331 2714 2415 2718
rect 2419 2714 2503 2718
rect 2507 2714 2591 2718
rect 2595 2714 2663 2718
rect 2667 2714 2679 2718
rect 2683 2714 2767 2718
rect 2771 2714 2799 2718
rect 2803 2714 2855 2718
rect 2859 2714 2943 2718
rect 2947 2714 2959 2718
rect 2963 2714 3031 2718
rect 3035 2714 3119 2718
rect 3123 2714 3135 2718
rect 3139 2714 3207 2718
rect 3211 2714 3295 2718
rect 3299 2714 3319 2718
rect 3323 2714 3391 2718
rect 3395 2714 3479 2718
rect 3483 2714 3575 2718
rect 3579 2714 3599 2718
rect 1841 2713 3599 2714
rect 3605 2713 3606 2719
rect 84 2689 85 2695
rect 91 2694 1835 2695
rect 91 2690 111 2694
rect 115 2690 199 2694
rect 203 2690 215 2694
rect 219 2690 327 2694
rect 331 2690 335 2694
rect 339 2690 463 2694
rect 467 2690 583 2694
rect 587 2690 599 2694
rect 603 2690 703 2694
rect 707 2690 743 2694
rect 747 2690 823 2694
rect 827 2690 879 2694
rect 883 2690 935 2694
rect 939 2690 1015 2694
rect 1019 2690 1047 2694
rect 1051 2690 1143 2694
rect 1147 2690 1159 2694
rect 1163 2690 1271 2694
rect 1275 2690 1279 2694
rect 1283 2690 1415 2694
rect 1419 2690 1823 2694
rect 1827 2690 1835 2694
rect 91 2689 1835 2690
rect 1841 2689 1842 2695
rect 842 2636 848 2637
rect 1226 2636 1232 2637
rect 842 2632 843 2636
rect 847 2632 1227 2636
rect 1231 2632 1232 2636
rect 842 2631 848 2632
rect 1226 2631 1232 2632
rect 1846 2625 1847 2631
rect 1853 2630 3611 2631
rect 1853 2626 1863 2630
rect 1867 2626 1895 2630
rect 1899 2626 1983 2630
rect 1987 2626 2071 2630
rect 2075 2626 2159 2630
rect 2163 2626 2247 2630
rect 2251 2626 2279 2630
rect 2283 2626 2335 2630
rect 2339 2626 2415 2630
rect 2419 2626 2423 2630
rect 2427 2626 2511 2630
rect 2515 2626 2551 2630
rect 2555 2626 2599 2630
rect 2603 2626 2687 2630
rect 2691 2626 2695 2630
rect 2699 2626 2775 2630
rect 2779 2626 2847 2630
rect 2851 2626 2863 2630
rect 2867 2626 2951 2630
rect 2955 2626 2999 2630
rect 3003 2626 3039 2630
rect 3043 2626 3127 2630
rect 3131 2626 3159 2630
rect 3163 2626 3215 2630
rect 3219 2626 3303 2630
rect 3307 2626 3399 2630
rect 3403 2626 3487 2630
rect 3491 2626 3575 2630
rect 3579 2626 3611 2630
rect 1853 2625 3611 2626
rect 3617 2625 3618 2631
rect 1846 2623 1854 2625
rect 96 2617 97 2623
rect 103 2622 1847 2623
rect 103 2618 111 2622
rect 115 2618 223 2622
rect 227 2618 343 2622
rect 347 2618 471 2622
rect 475 2618 559 2622
rect 563 2618 591 2622
rect 595 2618 647 2622
rect 651 2618 711 2622
rect 715 2618 735 2622
rect 739 2618 823 2622
rect 827 2618 831 2622
rect 835 2618 911 2622
rect 915 2618 943 2622
rect 947 2618 999 2622
rect 1003 2618 1055 2622
rect 1059 2618 1087 2622
rect 1091 2618 1167 2622
rect 1171 2618 1175 2622
rect 1179 2618 1263 2622
rect 1267 2618 1279 2622
rect 1283 2618 1823 2622
rect 1827 2618 1847 2622
rect 103 2617 1847 2618
rect 1853 2617 1854 2623
rect 1950 2596 1956 2597
rect 2642 2596 2648 2597
rect 1950 2592 1951 2596
rect 1955 2592 2643 2596
rect 2647 2592 2648 2596
rect 1950 2591 1956 2592
rect 2642 2591 2648 2592
rect 1834 2557 1835 2563
rect 1841 2562 3599 2563
rect 1841 2558 1863 2562
rect 1867 2558 2103 2562
rect 2107 2558 2151 2562
rect 2155 2558 2199 2562
rect 2203 2558 2271 2562
rect 2275 2558 2311 2562
rect 2315 2558 2407 2562
rect 2411 2558 2431 2562
rect 2435 2558 2543 2562
rect 2547 2558 2559 2562
rect 2563 2558 2687 2562
rect 2691 2558 2695 2562
rect 2699 2558 2839 2562
rect 2843 2558 2847 2562
rect 2851 2558 2991 2562
rect 2995 2558 2999 2562
rect 3003 2558 3151 2562
rect 3155 2558 3159 2562
rect 3163 2558 3327 2562
rect 3331 2558 3479 2562
rect 3483 2558 3575 2562
rect 3579 2558 3599 2562
rect 1841 2557 3599 2558
rect 3605 2557 3606 2563
rect 84 2541 85 2547
rect 91 2546 1835 2547
rect 91 2542 111 2546
rect 115 2542 463 2546
rect 467 2542 495 2546
rect 499 2542 551 2546
rect 555 2542 583 2546
rect 587 2542 639 2546
rect 643 2542 671 2546
rect 675 2542 727 2546
rect 731 2542 759 2546
rect 763 2542 815 2546
rect 819 2542 847 2546
rect 851 2542 903 2546
rect 907 2542 935 2546
rect 939 2542 991 2546
rect 995 2542 1023 2546
rect 1027 2542 1079 2546
rect 1083 2542 1111 2546
rect 1115 2542 1167 2546
rect 1171 2542 1199 2546
rect 1203 2542 1255 2546
rect 1259 2542 1287 2546
rect 1291 2542 1823 2546
rect 1827 2542 1835 2546
rect 91 2541 1835 2542
rect 1841 2541 1842 2547
rect 978 2492 984 2493
rect 1266 2492 1272 2493
rect 978 2488 979 2492
rect 983 2488 1267 2492
rect 1271 2488 1272 2492
rect 978 2487 984 2488
rect 1266 2487 1272 2488
rect 1846 2485 1847 2491
rect 1853 2490 3611 2491
rect 1853 2486 1863 2490
rect 1867 2486 2087 2490
rect 2091 2486 2111 2490
rect 2115 2486 2183 2490
rect 2187 2486 2207 2490
rect 2211 2486 2287 2490
rect 2291 2486 2319 2490
rect 2323 2486 2407 2490
rect 2411 2486 2439 2490
rect 2443 2486 2543 2490
rect 2547 2486 2567 2490
rect 2571 2486 2703 2490
rect 2707 2486 2855 2490
rect 2859 2486 2887 2490
rect 2891 2486 3007 2490
rect 3011 2486 3087 2490
rect 3091 2486 3167 2490
rect 3171 2486 3295 2490
rect 3299 2486 3335 2490
rect 3339 2486 3487 2490
rect 3491 2486 3575 2490
rect 3579 2486 3611 2490
rect 1853 2485 3611 2486
rect 3617 2485 3618 2491
rect 96 2469 97 2475
rect 103 2474 1847 2475
rect 103 2470 111 2474
rect 115 2470 359 2474
rect 363 2470 471 2474
rect 475 2470 503 2474
rect 507 2470 591 2474
rect 595 2470 679 2474
rect 683 2470 719 2474
rect 723 2470 767 2474
rect 771 2470 847 2474
rect 851 2470 855 2474
rect 859 2470 943 2474
rect 947 2470 967 2474
rect 971 2470 1031 2474
rect 1035 2470 1087 2474
rect 1091 2470 1119 2474
rect 1123 2470 1207 2474
rect 1211 2470 1295 2474
rect 1299 2470 1335 2474
rect 1339 2470 1463 2474
rect 1467 2470 1823 2474
rect 1827 2470 1847 2474
rect 103 2469 1847 2470
rect 1853 2469 1854 2475
rect 2098 2468 2104 2469
rect 2378 2468 2384 2469
rect 2098 2464 2099 2468
rect 2103 2464 2379 2468
rect 2383 2464 2384 2468
rect 2098 2463 2104 2464
rect 2378 2463 2384 2464
rect 414 2460 420 2461
rect 786 2460 792 2461
rect 414 2456 415 2460
rect 419 2456 787 2460
rect 791 2456 792 2460
rect 414 2455 420 2456
rect 786 2455 792 2456
rect 1834 2413 1835 2419
rect 1841 2418 3599 2419
rect 1841 2414 1863 2418
rect 1867 2414 1951 2418
rect 1955 2414 2063 2418
rect 2067 2414 2079 2418
rect 2083 2414 2175 2418
rect 2179 2414 2183 2418
rect 2187 2414 2279 2418
rect 2283 2414 2311 2418
rect 2315 2414 2399 2418
rect 2403 2414 2447 2418
rect 2451 2414 2535 2418
rect 2539 2414 2591 2418
rect 2595 2414 2695 2418
rect 2699 2414 2751 2418
rect 2755 2414 2879 2418
rect 2883 2414 2927 2418
rect 2931 2414 3079 2418
rect 3083 2414 3111 2418
rect 3115 2414 3287 2418
rect 3291 2414 3303 2418
rect 3307 2414 3479 2418
rect 3483 2414 3575 2418
rect 3579 2414 3599 2418
rect 1841 2413 3599 2414
rect 3605 2413 3606 2419
rect 84 2397 85 2403
rect 91 2402 1835 2403
rect 91 2398 111 2402
rect 115 2398 135 2402
rect 139 2398 287 2402
rect 291 2398 351 2402
rect 355 2398 463 2402
rect 467 2398 471 2402
rect 475 2398 583 2402
rect 587 2398 663 2402
rect 667 2398 711 2402
rect 715 2398 839 2402
rect 843 2398 847 2402
rect 851 2398 959 2402
rect 963 2398 1031 2402
rect 1035 2398 1079 2402
rect 1083 2398 1199 2402
rect 1203 2398 1207 2402
rect 1211 2398 1327 2402
rect 1331 2398 1375 2402
rect 1379 2398 1455 2402
rect 1459 2398 1543 2402
rect 1547 2398 1711 2402
rect 1715 2398 1823 2402
rect 1827 2398 1835 2402
rect 91 2397 1835 2398
rect 1841 2397 1842 2403
rect 1094 2348 1100 2349
rect 1402 2348 1408 2349
rect 1094 2344 1095 2348
rect 1099 2344 1403 2348
rect 1407 2344 1408 2348
rect 1094 2343 1100 2344
rect 1402 2343 1408 2344
rect 1846 2337 1847 2343
rect 1853 2342 3611 2343
rect 1853 2338 1863 2342
rect 1867 2338 1895 2342
rect 1899 2338 1959 2342
rect 1963 2338 2007 2342
rect 2011 2338 2071 2342
rect 2075 2338 2159 2342
rect 2163 2338 2191 2342
rect 2195 2338 2311 2342
rect 2315 2338 2319 2342
rect 2323 2338 2455 2342
rect 2459 2338 2463 2342
rect 2467 2338 2599 2342
rect 2603 2338 2615 2342
rect 2619 2338 2759 2342
rect 2763 2338 2775 2342
rect 2779 2338 2935 2342
rect 2939 2338 2943 2342
rect 2947 2338 3111 2342
rect 3115 2338 3119 2342
rect 3123 2338 3287 2342
rect 3291 2338 3311 2342
rect 3315 2338 3471 2342
rect 3475 2338 3487 2342
rect 3491 2338 3575 2342
rect 3579 2338 3611 2342
rect 1853 2337 3611 2338
rect 3617 2337 3618 2343
rect 96 2325 97 2331
rect 103 2330 1847 2331
rect 103 2326 111 2330
rect 115 2326 143 2330
rect 147 2326 295 2330
rect 299 2326 479 2330
rect 483 2326 671 2330
rect 675 2326 855 2330
rect 859 2326 863 2330
rect 867 2326 1039 2330
rect 1043 2326 1055 2330
rect 1059 2326 1215 2330
rect 1219 2326 1231 2330
rect 1235 2326 1383 2330
rect 1387 2326 1407 2330
rect 1411 2326 1551 2330
rect 1555 2326 1583 2330
rect 1587 2326 1719 2330
rect 1723 2326 1735 2330
rect 1739 2326 1823 2330
rect 1827 2326 1847 2330
rect 103 2325 1847 2326
rect 1853 2325 1854 2331
rect 2046 2324 2052 2325
rect 2402 2324 2408 2325
rect 2046 2320 2047 2324
rect 2051 2320 2403 2324
rect 2407 2320 2408 2324
rect 2046 2319 2052 2320
rect 2402 2319 2408 2320
rect 1150 2300 1156 2301
rect 1338 2300 1344 2301
rect 1150 2296 1151 2300
rect 1155 2296 1339 2300
rect 1343 2296 1344 2300
rect 1150 2295 1156 2296
rect 1338 2295 1344 2296
rect 1834 2265 1835 2271
rect 1841 2270 3599 2271
rect 1841 2266 1863 2270
rect 1867 2266 1887 2270
rect 1891 2266 1999 2270
rect 2003 2266 2023 2270
rect 2027 2266 2151 2270
rect 2155 2266 2199 2270
rect 2203 2266 2303 2270
rect 2307 2266 2383 2270
rect 2387 2266 2455 2270
rect 2459 2266 2567 2270
rect 2571 2266 2607 2270
rect 2611 2266 2743 2270
rect 2747 2266 2767 2270
rect 2771 2266 2911 2270
rect 2915 2266 2935 2270
rect 2939 2266 3079 2270
rect 3083 2266 3103 2270
rect 3107 2266 3239 2270
rect 3243 2266 3279 2270
rect 3283 2266 3407 2270
rect 3411 2266 3463 2270
rect 3467 2266 3575 2270
rect 3579 2266 3599 2270
rect 1841 2265 3599 2266
rect 3605 2265 3606 2271
rect 84 2249 85 2255
rect 91 2254 1835 2255
rect 91 2250 111 2254
rect 115 2250 135 2254
rect 139 2250 255 2254
rect 259 2250 287 2254
rect 291 2250 407 2254
rect 411 2250 471 2254
rect 475 2250 559 2254
rect 563 2250 663 2254
rect 667 2250 719 2254
rect 723 2250 855 2254
rect 859 2250 871 2254
rect 875 2250 1015 2254
rect 1019 2250 1047 2254
rect 1051 2250 1159 2254
rect 1163 2250 1223 2254
rect 1227 2250 1303 2254
rect 1307 2250 1399 2254
rect 1403 2250 1455 2254
rect 1459 2250 1575 2254
rect 1579 2250 1727 2254
rect 1731 2250 1823 2254
rect 1827 2250 1835 2254
rect 91 2249 1835 2250
rect 1841 2249 1842 2255
rect 1950 2252 1956 2253
rect 2478 2252 2484 2253
rect 1950 2248 1951 2252
rect 1955 2248 2479 2252
rect 2483 2248 2484 2252
rect 1950 2247 1956 2248
rect 2478 2247 2484 2248
rect 2770 2212 2776 2213
rect 3146 2212 3152 2213
rect 2770 2208 2771 2212
rect 2775 2208 3147 2212
rect 3151 2208 3152 2212
rect 2770 2207 2776 2208
rect 3146 2207 3152 2208
rect 890 2196 896 2197
rect 1098 2196 1104 2197
rect 890 2192 891 2196
rect 895 2192 1099 2196
rect 1103 2192 1104 2196
rect 890 2191 896 2192
rect 1098 2191 1104 2192
rect 1190 2196 1196 2197
rect 1398 2196 1404 2197
rect 1190 2192 1191 2196
rect 1195 2192 1399 2196
rect 1403 2192 1404 2196
rect 1846 2193 1847 2199
rect 1853 2198 3611 2199
rect 1853 2194 1863 2198
rect 1867 2194 1895 2198
rect 1899 2194 2031 2198
rect 2035 2194 2039 2198
rect 2043 2194 2207 2198
rect 2211 2194 2215 2198
rect 2219 2194 2391 2198
rect 2395 2194 2399 2198
rect 2403 2194 2575 2198
rect 2579 2194 2583 2198
rect 2587 2194 2751 2198
rect 2755 2194 2759 2198
rect 2763 2194 2919 2198
rect 2923 2194 3071 2198
rect 3075 2194 3087 2198
rect 3091 2194 3215 2198
rect 3219 2194 3247 2198
rect 3251 2194 3359 2198
rect 3363 2194 3415 2198
rect 3419 2194 3487 2198
rect 3491 2194 3575 2198
rect 3579 2194 3611 2198
rect 1853 2193 3611 2194
rect 3617 2193 3618 2199
rect 1190 2191 1196 2192
rect 1398 2191 1404 2192
rect 96 2177 97 2183
rect 103 2182 1847 2183
rect 103 2178 111 2182
rect 115 2178 143 2182
rect 147 2178 215 2182
rect 219 2178 263 2182
rect 267 2178 311 2182
rect 315 2178 415 2182
rect 419 2178 519 2182
rect 523 2178 567 2182
rect 571 2178 623 2182
rect 627 2178 727 2182
rect 731 2178 831 2182
rect 835 2178 879 2182
rect 883 2178 943 2182
rect 947 2178 1023 2182
rect 1027 2178 1055 2182
rect 1059 2178 1167 2182
rect 1171 2178 1311 2182
rect 1315 2178 1463 2182
rect 1467 2178 1823 2182
rect 1827 2178 1847 2182
rect 103 2177 1847 2178
rect 1853 2177 1854 2183
rect 2006 2180 2012 2181
rect 2506 2180 2512 2181
rect 2006 2176 2007 2180
rect 2011 2176 2507 2180
rect 2511 2176 2512 2180
rect 2006 2175 2012 2176
rect 2506 2175 2512 2176
rect 1834 2121 1835 2127
rect 1841 2126 3599 2127
rect 1841 2122 1863 2126
rect 1867 2122 1887 2126
rect 1891 2122 2023 2126
rect 2027 2122 2031 2126
rect 2035 2122 2199 2126
rect 2203 2122 2207 2126
rect 2211 2122 2375 2126
rect 2379 2122 2391 2126
rect 2395 2122 2551 2126
rect 2555 2122 2575 2126
rect 2579 2122 2719 2126
rect 2723 2122 2751 2126
rect 2755 2122 2879 2126
rect 2883 2122 2911 2126
rect 2915 2122 3031 2126
rect 3035 2122 3063 2126
rect 3067 2122 3175 2126
rect 3179 2122 3207 2126
rect 3211 2122 3319 2126
rect 3323 2122 3351 2126
rect 3355 2122 3471 2126
rect 3475 2122 3479 2126
rect 3483 2122 3575 2126
rect 3579 2122 3599 2126
rect 1841 2121 3599 2122
rect 3605 2121 3606 2127
rect 84 2101 85 2107
rect 91 2106 1835 2107
rect 91 2102 111 2106
rect 115 2102 207 2106
rect 211 2102 303 2106
rect 307 2102 319 2106
rect 323 2102 407 2106
rect 411 2102 423 2106
rect 427 2102 511 2106
rect 515 2102 527 2106
rect 531 2102 615 2106
rect 619 2102 631 2106
rect 635 2102 719 2106
rect 723 2102 735 2106
rect 739 2102 823 2106
rect 827 2102 831 2106
rect 835 2102 927 2106
rect 931 2102 935 2106
rect 939 2102 1031 2106
rect 1035 2102 1047 2106
rect 1051 2102 1135 2106
rect 1139 2102 1159 2106
rect 1163 2102 1239 2106
rect 1243 2102 1823 2106
rect 1827 2102 1835 2106
rect 91 2101 1835 2102
rect 1841 2101 1842 2107
rect 2038 2068 2044 2069
rect 2478 2068 2484 2069
rect 2038 2064 2039 2068
rect 2043 2064 2479 2068
rect 2483 2064 2484 2068
rect 2038 2063 2044 2064
rect 2478 2063 2484 2064
rect 1846 2045 1847 2051
rect 1853 2050 3611 2051
rect 1853 2046 1863 2050
rect 1867 2046 1895 2050
rect 1899 2046 2015 2050
rect 2019 2046 2031 2050
rect 2035 2046 2151 2050
rect 2155 2046 2207 2050
rect 2211 2046 2295 2050
rect 2299 2046 2383 2050
rect 2387 2046 2439 2050
rect 2443 2046 2559 2050
rect 2563 2046 2591 2050
rect 2595 2046 2727 2050
rect 2731 2046 2759 2050
rect 2763 2046 2887 2050
rect 2891 2046 2935 2050
rect 2939 2046 3039 2050
rect 3043 2046 3119 2050
rect 3123 2046 3183 2050
rect 3187 2046 3311 2050
rect 3315 2046 3327 2050
rect 3331 2046 3479 2050
rect 3483 2046 3487 2050
rect 3491 2046 3575 2050
rect 3579 2046 3611 2050
rect 1853 2045 3611 2046
rect 3617 2045 3618 2051
rect 96 2025 97 2031
rect 103 2030 1847 2031
rect 103 2026 111 2030
rect 115 2026 215 2030
rect 219 2026 327 2030
rect 331 2026 391 2030
rect 395 2026 431 2030
rect 435 2026 535 2030
rect 539 2026 559 2030
rect 563 2026 639 2030
rect 643 2026 719 2030
rect 723 2026 743 2030
rect 747 2026 839 2030
rect 843 2026 863 2030
rect 867 2026 935 2030
rect 939 2026 999 2030
rect 1003 2026 1039 2030
rect 1043 2026 1127 2030
rect 1131 2026 1143 2030
rect 1147 2026 1247 2030
rect 1251 2026 1367 2030
rect 1371 2026 1495 2030
rect 1499 2026 1823 2030
rect 1827 2026 1847 2030
rect 103 2025 1847 2026
rect 1853 2025 1854 2031
rect 2006 2028 2012 2029
rect 2222 2028 2228 2029
rect 2006 2024 2007 2028
rect 2011 2024 2223 2028
rect 2227 2024 2228 2028
rect 2006 2023 2012 2024
rect 2222 2023 2228 2024
rect 1834 1973 1835 1979
rect 1841 1978 3599 1979
rect 1841 1974 1863 1978
rect 1867 1974 1887 1978
rect 1891 1974 2007 1978
rect 2011 1974 2023 1978
rect 2027 1974 2111 1978
rect 2115 1974 2143 1978
rect 2147 1974 2199 1978
rect 2203 1974 2287 1978
rect 2291 1974 2383 1978
rect 2387 1974 2431 1978
rect 2435 1974 2503 1978
rect 2507 1974 2583 1978
rect 2587 1974 2655 1978
rect 2659 1974 2751 1978
rect 2755 1974 2839 1978
rect 2843 1974 2927 1978
rect 2931 1974 3047 1978
rect 3051 1974 3111 1978
rect 3115 1974 3271 1978
rect 3275 1974 3303 1978
rect 3307 1974 3479 1978
rect 3483 1974 3575 1978
rect 3579 1974 3599 1978
rect 1841 1973 3599 1974
rect 3605 1973 3606 1979
rect 84 1949 85 1955
rect 91 1954 1835 1955
rect 91 1950 111 1954
rect 115 1950 135 1954
rect 139 1950 207 1954
rect 211 1950 311 1954
rect 315 1950 383 1954
rect 387 1950 519 1954
rect 523 1950 551 1954
rect 555 1950 711 1954
rect 715 1950 719 1954
rect 723 1950 855 1954
rect 859 1950 911 1954
rect 915 1950 991 1954
rect 995 1950 1095 1954
rect 1099 1950 1119 1954
rect 1123 1950 1239 1954
rect 1243 1950 1263 1954
rect 1267 1950 1359 1954
rect 1363 1950 1423 1954
rect 1427 1950 1487 1954
rect 1491 1950 1583 1954
rect 1587 1950 1727 1954
rect 1731 1950 1823 1954
rect 1827 1950 1835 1954
rect 91 1949 1835 1950
rect 1841 1949 1842 1955
rect 1846 1897 1847 1903
rect 1853 1902 3611 1903
rect 1853 1898 1863 1902
rect 1867 1898 2031 1902
rect 2035 1898 2119 1902
rect 2123 1898 2175 1902
rect 2179 1898 2207 1902
rect 2211 1898 2263 1902
rect 2267 1898 2295 1902
rect 2299 1898 2351 1902
rect 2355 1898 2391 1902
rect 2395 1898 2439 1902
rect 2443 1898 2511 1902
rect 2515 1898 2527 1902
rect 2531 1898 2639 1902
rect 2643 1898 2663 1902
rect 2667 1898 2775 1902
rect 2779 1898 2847 1902
rect 2851 1898 2935 1902
rect 2939 1898 3055 1902
rect 3059 1898 3119 1902
rect 3123 1898 3279 1902
rect 3283 1898 3311 1902
rect 3315 1898 3487 1902
rect 3491 1898 3575 1902
rect 3579 1898 3611 1902
rect 1853 1897 3611 1898
rect 3617 1897 3618 1903
rect 96 1873 97 1879
rect 103 1878 1847 1879
rect 103 1874 111 1878
rect 115 1874 143 1878
rect 147 1874 311 1878
rect 315 1874 319 1878
rect 323 1874 511 1878
rect 515 1874 527 1878
rect 531 1874 703 1878
rect 707 1874 727 1878
rect 731 1874 887 1878
rect 891 1874 919 1878
rect 923 1874 1063 1878
rect 1067 1874 1103 1878
rect 1107 1874 1231 1878
rect 1235 1874 1271 1878
rect 1275 1874 1391 1878
rect 1395 1874 1431 1878
rect 1435 1874 1551 1878
rect 1555 1874 1591 1878
rect 1595 1874 1711 1878
rect 1715 1874 1735 1878
rect 1739 1874 1823 1878
rect 1827 1874 1847 1878
rect 103 1873 1847 1874
rect 1853 1873 1854 1879
rect 1134 1868 1140 1869
rect 1298 1868 1304 1869
rect 1134 1864 1135 1868
rect 1139 1864 1299 1868
rect 1303 1864 1304 1868
rect 1134 1863 1140 1864
rect 1298 1863 1304 1864
rect 1834 1825 1835 1831
rect 1841 1830 3599 1831
rect 1841 1826 1863 1830
rect 1867 1826 2167 1830
rect 2171 1826 2255 1830
rect 2259 1826 2319 1830
rect 2323 1826 2343 1830
rect 2347 1826 2431 1830
rect 2435 1826 2439 1830
rect 2443 1826 2519 1830
rect 2523 1826 2559 1830
rect 2563 1826 2631 1830
rect 2635 1826 2679 1830
rect 2683 1826 2767 1830
rect 2771 1826 2799 1830
rect 2803 1826 2919 1830
rect 2923 1826 2927 1830
rect 2931 1826 3047 1830
rect 3051 1826 3111 1830
rect 3115 1826 3183 1830
rect 3187 1826 3303 1830
rect 3307 1826 3319 1830
rect 3323 1826 3463 1830
rect 3467 1826 3479 1830
rect 3483 1826 3575 1830
rect 3579 1826 3599 1830
rect 1841 1825 3599 1826
rect 3605 1825 3606 1831
rect 84 1797 85 1803
rect 91 1802 1835 1803
rect 91 1798 111 1802
rect 115 1798 135 1802
rect 139 1798 263 1802
rect 267 1798 303 1802
rect 307 1798 415 1802
rect 419 1798 503 1802
rect 507 1798 567 1802
rect 571 1798 695 1802
rect 699 1798 719 1802
rect 723 1798 863 1802
rect 867 1798 879 1802
rect 883 1798 1007 1802
rect 1011 1798 1055 1802
rect 1059 1798 1143 1802
rect 1147 1798 1223 1802
rect 1227 1798 1279 1802
rect 1283 1798 1383 1802
rect 1387 1798 1423 1802
rect 1427 1798 1543 1802
rect 1547 1798 1703 1802
rect 1707 1798 1823 1802
rect 1827 1798 1835 1802
rect 91 1797 1835 1798
rect 1841 1797 1842 1803
rect 2818 1772 2824 1773
rect 3198 1772 3204 1773
rect 2818 1768 2819 1772
rect 2823 1768 3199 1772
rect 3203 1768 3204 1772
rect 2818 1767 2824 1768
rect 3198 1767 3204 1768
rect 1846 1749 1847 1755
rect 1853 1754 3611 1755
rect 1853 1750 1863 1754
rect 1867 1750 2295 1754
rect 2299 1750 2327 1754
rect 2331 1750 2407 1754
rect 2411 1750 2447 1754
rect 2451 1750 2527 1754
rect 2531 1750 2567 1754
rect 2571 1750 2655 1754
rect 2659 1750 2687 1754
rect 2691 1750 2775 1754
rect 2779 1750 2807 1754
rect 2811 1750 2895 1754
rect 2899 1750 2927 1754
rect 2931 1750 3015 1754
rect 3019 1750 3055 1754
rect 3059 1750 3135 1754
rect 3139 1750 3191 1754
rect 3195 1750 3255 1754
rect 3259 1750 3327 1754
rect 3331 1750 3383 1754
rect 3387 1750 3471 1754
rect 3475 1750 3487 1754
rect 3491 1750 3575 1754
rect 3579 1750 3611 1754
rect 1853 1749 3611 1750
rect 3617 1749 3618 1755
rect 96 1729 97 1735
rect 103 1734 1847 1735
rect 103 1730 111 1734
rect 115 1730 143 1734
rect 147 1730 271 1734
rect 275 1730 279 1734
rect 283 1730 423 1734
rect 427 1730 431 1734
rect 435 1730 575 1734
rect 579 1730 583 1734
rect 587 1730 727 1734
rect 731 1730 863 1734
rect 867 1730 871 1734
rect 875 1730 991 1734
rect 995 1730 1015 1734
rect 1019 1730 1127 1734
rect 1131 1730 1151 1734
rect 1155 1730 1263 1734
rect 1267 1730 1287 1734
rect 1291 1730 1431 1734
rect 1435 1730 1823 1734
rect 1827 1730 1847 1734
rect 103 1729 1847 1730
rect 1853 1729 1854 1735
rect 1834 1677 1835 1683
rect 1841 1682 3599 1683
rect 1841 1678 1863 1682
rect 1867 1678 2143 1682
rect 2147 1678 2247 1682
rect 2251 1678 2287 1682
rect 2291 1678 2367 1682
rect 2371 1678 2399 1682
rect 2403 1678 2503 1682
rect 2507 1678 2519 1682
rect 2523 1678 2647 1682
rect 2651 1678 2767 1682
rect 2771 1678 2807 1682
rect 2811 1678 2887 1682
rect 2891 1678 2975 1682
rect 2979 1678 3007 1682
rect 3011 1678 3127 1682
rect 3131 1678 3143 1682
rect 3147 1678 3247 1682
rect 3251 1678 3319 1682
rect 3323 1678 3375 1682
rect 3379 1678 3479 1682
rect 3483 1678 3575 1682
rect 3579 1678 3599 1682
rect 1841 1677 3599 1678
rect 3605 1677 3606 1683
rect 84 1661 85 1667
rect 91 1666 1835 1667
rect 91 1662 111 1666
rect 115 1662 135 1666
rect 139 1662 263 1666
rect 267 1662 271 1666
rect 275 1662 423 1666
rect 427 1662 575 1666
rect 579 1662 719 1666
rect 723 1662 727 1666
rect 731 1662 855 1666
rect 859 1662 871 1666
rect 875 1662 983 1666
rect 987 1662 1007 1666
rect 1011 1662 1119 1666
rect 1123 1662 1143 1666
rect 1147 1662 1255 1666
rect 1259 1662 1279 1666
rect 1283 1662 1415 1666
rect 1419 1662 1823 1666
rect 1827 1662 1835 1666
rect 91 1661 1835 1662
rect 1841 1661 1842 1667
rect 1022 1628 1028 1629
rect 1346 1628 1352 1629
rect 1022 1624 1023 1628
rect 1027 1624 1347 1628
rect 1351 1624 1352 1628
rect 1022 1623 1028 1624
rect 1346 1623 1352 1624
rect 442 1612 448 1613
rect 642 1612 648 1613
rect 442 1608 443 1612
rect 447 1608 643 1612
rect 647 1608 648 1612
rect 442 1607 448 1608
rect 642 1607 648 1608
rect 890 1612 896 1613
rect 1210 1612 1216 1613
rect 890 1608 891 1612
rect 895 1608 1211 1612
rect 1215 1608 1216 1612
rect 1846 1609 1847 1615
rect 1853 1614 3611 1615
rect 1853 1610 1863 1614
rect 1867 1610 2007 1614
rect 2011 1610 2103 1614
rect 2107 1610 2151 1614
rect 2155 1610 2207 1614
rect 2211 1610 2255 1614
rect 2259 1610 2327 1614
rect 2331 1610 2375 1614
rect 2379 1610 2463 1614
rect 2467 1610 2511 1614
rect 2515 1610 2607 1614
rect 2611 1610 2655 1614
rect 2659 1610 2767 1614
rect 2771 1610 2815 1614
rect 2819 1610 2943 1614
rect 2947 1610 2983 1614
rect 2987 1610 3127 1614
rect 3131 1610 3151 1614
rect 3155 1610 3319 1614
rect 3323 1610 3327 1614
rect 3331 1610 3487 1614
rect 3491 1610 3575 1614
rect 3579 1610 3611 1614
rect 1853 1609 3611 1610
rect 3617 1609 3618 1615
rect 890 1607 896 1608
rect 1210 1607 1216 1608
rect 2018 1604 2024 1605
rect 2306 1604 2312 1605
rect 2018 1600 2019 1604
rect 2023 1600 2307 1604
rect 2311 1600 2312 1604
rect 2018 1599 2024 1600
rect 2306 1599 2312 1600
rect 96 1589 97 1595
rect 103 1594 1847 1595
rect 103 1590 111 1594
rect 115 1590 143 1594
rect 147 1590 167 1594
rect 171 1590 271 1594
rect 275 1590 335 1594
rect 339 1590 431 1594
rect 435 1590 511 1594
rect 515 1590 583 1594
rect 587 1590 679 1594
rect 683 1590 735 1594
rect 739 1590 847 1594
rect 851 1590 879 1594
rect 883 1590 999 1594
rect 1003 1590 1015 1594
rect 1019 1590 1151 1594
rect 1155 1590 1287 1594
rect 1291 1590 1295 1594
rect 1299 1590 1423 1594
rect 1427 1590 1439 1594
rect 1443 1590 1583 1594
rect 1587 1590 1823 1594
rect 1827 1590 1847 1594
rect 103 1589 1847 1590
rect 1853 1589 1854 1595
rect 1834 1533 1835 1539
rect 1841 1538 3599 1539
rect 1841 1534 1863 1538
rect 1867 1534 1887 1538
rect 1891 1534 1975 1538
rect 1979 1534 1999 1538
rect 2003 1534 2095 1538
rect 2099 1534 2103 1538
rect 2107 1534 2199 1538
rect 2203 1534 2239 1538
rect 2243 1534 2319 1538
rect 2323 1534 2383 1538
rect 2387 1534 2455 1538
rect 2459 1534 2543 1538
rect 2547 1534 2599 1538
rect 2603 1534 2711 1538
rect 2715 1534 2759 1538
rect 2763 1534 2879 1538
rect 2883 1534 2935 1538
rect 2939 1534 3055 1538
rect 3059 1534 3119 1538
rect 3123 1534 3239 1538
rect 3243 1534 3311 1538
rect 3315 1534 3431 1538
rect 3435 1534 3479 1538
rect 3483 1534 3575 1538
rect 3579 1534 3599 1538
rect 1841 1533 3599 1534
rect 3605 1533 3606 1539
rect 84 1517 85 1523
rect 91 1522 1835 1523
rect 91 1518 111 1522
rect 115 1518 159 1522
rect 163 1518 215 1522
rect 219 1518 327 1522
rect 331 1518 391 1522
rect 395 1518 503 1522
rect 507 1518 575 1522
rect 579 1518 671 1522
rect 675 1518 759 1522
rect 763 1518 839 1522
rect 843 1518 935 1522
rect 939 1518 991 1522
rect 995 1518 1095 1522
rect 1099 1518 1143 1522
rect 1147 1518 1255 1522
rect 1259 1518 1287 1522
rect 1291 1518 1407 1522
rect 1411 1518 1431 1522
rect 1435 1518 1559 1522
rect 1563 1518 1575 1522
rect 1579 1518 1711 1522
rect 1715 1518 1823 1522
rect 1827 1518 1835 1522
rect 91 1517 1835 1518
rect 1841 1517 1842 1523
rect 1114 1468 1120 1469
rect 1518 1468 1524 1469
rect 1114 1464 1115 1468
rect 1119 1464 1519 1468
rect 1523 1464 1524 1468
rect 1114 1463 1120 1464
rect 1518 1463 1524 1464
rect 1846 1461 1847 1467
rect 1853 1466 3611 1467
rect 1853 1462 1863 1466
rect 1867 1462 1895 1466
rect 1899 1462 1983 1466
rect 1987 1462 2023 1466
rect 2027 1462 2111 1466
rect 2115 1462 2175 1466
rect 2179 1462 2247 1466
rect 2251 1462 2319 1466
rect 2323 1462 2391 1466
rect 2395 1462 2463 1466
rect 2467 1462 2551 1466
rect 2555 1462 2615 1466
rect 2619 1462 2719 1466
rect 2723 1462 2767 1466
rect 2771 1462 2887 1466
rect 2891 1462 2935 1466
rect 2939 1462 3063 1466
rect 3067 1462 3103 1466
rect 3107 1462 3247 1466
rect 3251 1462 3279 1466
rect 3283 1462 3439 1466
rect 3443 1462 3463 1466
rect 3467 1462 3575 1466
rect 3579 1462 3611 1466
rect 1853 1461 3611 1462
rect 3617 1461 3618 1467
rect 96 1445 97 1451
rect 103 1450 1847 1451
rect 103 1446 111 1450
rect 115 1446 223 1450
rect 227 1446 255 1450
rect 259 1446 383 1450
rect 387 1446 399 1450
rect 403 1446 519 1450
rect 523 1446 583 1450
rect 587 1446 671 1450
rect 675 1446 767 1450
rect 771 1446 831 1450
rect 835 1446 943 1450
rect 947 1446 991 1450
rect 995 1446 1103 1450
rect 1107 1446 1143 1450
rect 1147 1446 1263 1450
rect 1267 1446 1295 1450
rect 1299 1446 1415 1450
rect 1419 1446 1447 1450
rect 1451 1446 1567 1450
rect 1571 1446 1599 1450
rect 1603 1446 1719 1450
rect 1723 1446 1735 1450
rect 1739 1446 1823 1450
rect 1827 1446 1847 1450
rect 103 1445 1847 1446
rect 1853 1445 1854 1451
rect 1950 1436 1956 1437
rect 2242 1436 2248 1437
rect 1950 1432 1951 1436
rect 1955 1432 2243 1436
rect 2247 1432 2248 1436
rect 1950 1431 1956 1432
rect 2242 1431 2248 1432
rect 1834 1386 3606 1387
rect 1834 1383 1863 1386
rect 84 1377 85 1383
rect 91 1382 1835 1383
rect 91 1378 111 1382
rect 115 1378 247 1382
rect 251 1378 351 1382
rect 355 1378 375 1382
rect 379 1378 439 1382
rect 443 1378 511 1382
rect 515 1378 527 1382
rect 531 1378 623 1382
rect 627 1378 663 1382
rect 667 1378 727 1382
rect 731 1378 823 1382
rect 827 1378 847 1382
rect 851 1378 983 1382
rect 987 1378 1127 1382
rect 1131 1378 1135 1382
rect 1139 1378 1279 1382
rect 1283 1378 1287 1382
rect 1291 1378 1431 1382
rect 1435 1378 1439 1382
rect 1443 1378 1591 1382
rect 1595 1378 1727 1382
rect 1731 1378 1823 1382
rect 1827 1378 1835 1382
rect 91 1377 1835 1378
rect 1841 1382 1863 1383
rect 1867 1382 1887 1386
rect 1891 1382 2015 1386
rect 2019 1382 2143 1386
rect 2147 1382 2167 1386
rect 2171 1382 2311 1386
rect 2315 1382 2391 1386
rect 2395 1382 2455 1386
rect 2459 1382 2607 1386
rect 2611 1382 2623 1386
rect 2627 1382 2759 1386
rect 2763 1382 2847 1386
rect 2851 1382 2927 1386
rect 2931 1382 3063 1386
rect 3067 1382 3095 1386
rect 3099 1382 3271 1386
rect 3275 1382 3455 1386
rect 3459 1382 3479 1386
rect 3483 1382 3575 1386
rect 3579 1382 3606 1386
rect 1841 1381 3606 1382
rect 1841 1377 1842 1381
rect 366 1348 372 1349
rect 514 1348 520 1349
rect 366 1344 367 1348
rect 371 1344 515 1348
rect 519 1344 520 1348
rect 366 1343 372 1344
rect 514 1343 520 1344
rect 1450 1332 1456 1333
rect 1870 1332 1876 1333
rect 1450 1328 1451 1332
rect 1455 1328 1871 1332
rect 1875 1328 1876 1332
rect 1450 1327 1456 1328
rect 1870 1327 1876 1328
rect 1846 1318 3618 1319
rect 1846 1315 1863 1318
rect 96 1309 97 1315
rect 103 1314 1847 1315
rect 103 1310 111 1314
rect 115 1310 359 1314
rect 363 1310 447 1314
rect 451 1310 455 1314
rect 459 1310 535 1314
rect 539 1310 543 1314
rect 547 1310 631 1314
rect 635 1310 719 1314
rect 723 1310 735 1314
rect 739 1310 831 1314
rect 835 1310 855 1314
rect 859 1310 967 1314
rect 971 1310 991 1314
rect 995 1310 1135 1314
rect 1139 1310 1287 1314
rect 1291 1310 1327 1314
rect 1331 1310 1439 1314
rect 1443 1310 1535 1314
rect 1539 1310 1599 1314
rect 1603 1310 1735 1314
rect 1739 1310 1823 1314
rect 1827 1310 1847 1314
rect 103 1309 1847 1310
rect 1853 1314 1863 1315
rect 1867 1314 1895 1318
rect 1899 1314 1927 1318
rect 1931 1314 2111 1318
rect 2115 1314 2151 1318
rect 2155 1314 2287 1318
rect 2291 1314 2399 1318
rect 2403 1314 2455 1318
rect 2459 1314 2623 1318
rect 2627 1314 2631 1318
rect 2635 1314 2791 1318
rect 2795 1314 2855 1318
rect 2859 1314 2959 1318
rect 2963 1314 3071 1318
rect 3075 1314 3135 1318
rect 3139 1314 3279 1318
rect 3283 1314 3319 1318
rect 3323 1314 3487 1318
rect 3491 1314 3575 1318
rect 3579 1314 3618 1318
rect 1853 1313 3618 1314
rect 1853 1309 1854 1313
rect 84 1241 85 1247
rect 91 1246 1835 1247
rect 91 1242 111 1246
rect 115 1242 447 1246
rect 451 1242 535 1246
rect 539 1242 543 1246
rect 547 1242 623 1246
rect 627 1242 631 1246
rect 635 1242 711 1246
rect 715 1242 719 1246
rect 723 1242 807 1246
rect 811 1242 823 1246
rect 827 1242 895 1246
rect 899 1242 959 1246
rect 963 1242 991 1246
rect 995 1242 1095 1246
rect 1099 1242 1127 1246
rect 1131 1242 1207 1246
rect 1211 1242 1319 1246
rect 1323 1242 1335 1246
rect 1339 1242 1471 1246
rect 1475 1242 1527 1246
rect 1531 1242 1607 1246
rect 1611 1242 1727 1246
rect 1731 1242 1823 1246
rect 1827 1242 1835 1246
rect 91 1241 1835 1242
rect 1841 1243 1842 1247
rect 1841 1242 3606 1243
rect 1841 1241 1863 1242
rect 1834 1238 1863 1241
rect 1867 1238 1919 1242
rect 1923 1238 2103 1242
rect 2107 1238 2143 1242
rect 2147 1238 2279 1242
rect 2283 1238 2319 1242
rect 2323 1238 2447 1242
rect 2451 1238 2487 1242
rect 2491 1238 2615 1242
rect 2619 1238 2655 1242
rect 2659 1238 2783 1242
rect 2787 1238 2823 1242
rect 2827 1238 2951 1242
rect 2955 1238 2991 1242
rect 2995 1238 3127 1242
rect 3131 1238 3159 1242
rect 3163 1238 3311 1242
rect 3315 1238 3327 1242
rect 3331 1238 3479 1242
rect 3483 1238 3575 1242
rect 3579 1238 3606 1242
rect 1834 1237 3606 1238
rect 1846 1174 3618 1175
rect 1846 1171 1863 1174
rect 96 1165 97 1171
rect 103 1170 1847 1171
rect 103 1166 111 1170
rect 115 1166 359 1170
rect 363 1166 471 1170
rect 475 1166 551 1170
rect 555 1166 591 1170
rect 595 1166 639 1170
rect 643 1166 711 1170
rect 715 1166 727 1170
rect 731 1166 815 1170
rect 819 1166 831 1170
rect 835 1166 903 1170
rect 907 1166 951 1170
rect 955 1166 999 1170
rect 1003 1166 1063 1170
rect 1067 1166 1103 1170
rect 1107 1166 1183 1170
rect 1187 1166 1215 1170
rect 1219 1166 1303 1170
rect 1307 1166 1343 1170
rect 1347 1166 1423 1170
rect 1427 1166 1479 1170
rect 1483 1166 1615 1170
rect 1619 1166 1735 1170
rect 1739 1166 1823 1170
rect 1827 1166 1847 1170
rect 103 1165 1847 1166
rect 1853 1170 1863 1171
rect 1867 1170 1895 1174
rect 1899 1170 2007 1174
rect 2011 1170 2143 1174
rect 2147 1170 2151 1174
rect 2155 1170 2295 1174
rect 2299 1170 2327 1174
rect 2331 1170 2455 1174
rect 2459 1170 2495 1174
rect 2499 1170 2623 1174
rect 2627 1170 2663 1174
rect 2667 1170 2791 1174
rect 2795 1170 2831 1174
rect 2835 1170 2967 1174
rect 2971 1170 2999 1174
rect 3003 1170 3143 1174
rect 3147 1170 3167 1174
rect 3171 1170 3327 1174
rect 3331 1170 3335 1174
rect 3339 1170 3487 1174
rect 3491 1170 3575 1174
rect 3579 1170 3618 1174
rect 1853 1169 3618 1170
rect 1853 1165 1854 1169
rect 414 1140 420 1141
rect 778 1140 784 1141
rect 414 1136 415 1140
rect 419 1136 779 1140
rect 783 1136 784 1140
rect 414 1135 420 1136
rect 778 1135 784 1136
rect 84 1093 85 1099
rect 91 1098 1835 1099
rect 91 1094 111 1098
rect 115 1094 143 1098
rect 147 1094 287 1098
rect 291 1094 351 1098
rect 355 1094 447 1098
rect 451 1094 463 1098
rect 467 1094 583 1098
rect 587 1094 615 1098
rect 619 1094 703 1098
rect 707 1094 783 1098
rect 787 1094 823 1098
rect 827 1094 943 1098
rect 947 1094 1055 1098
rect 1059 1094 1103 1098
rect 1107 1094 1175 1098
rect 1179 1094 1255 1098
rect 1259 1094 1295 1098
rect 1299 1094 1407 1098
rect 1411 1094 1415 1098
rect 1419 1094 1559 1098
rect 1563 1094 1823 1098
rect 1827 1094 1835 1098
rect 91 1093 1835 1094
rect 1841 1098 3606 1099
rect 1841 1094 1863 1098
rect 1867 1094 1887 1098
rect 1891 1094 1895 1098
rect 1899 1094 1999 1098
rect 2003 1094 2047 1098
rect 2051 1094 2135 1098
rect 2139 1094 2215 1098
rect 2219 1094 2287 1098
rect 2291 1094 2391 1098
rect 2395 1094 2447 1098
rect 2451 1094 2567 1098
rect 2571 1094 2615 1098
rect 2619 1094 2735 1098
rect 2739 1094 2783 1098
rect 2787 1094 2895 1098
rect 2899 1094 2959 1098
rect 2963 1094 3047 1098
rect 3051 1094 3135 1098
rect 3139 1094 3199 1098
rect 3203 1094 3319 1098
rect 3323 1094 3351 1098
rect 3355 1094 3479 1098
rect 3483 1094 3575 1098
rect 3579 1094 3606 1098
rect 1841 1093 3606 1094
rect 162 1044 168 1045
rect 682 1044 688 1045
rect 162 1040 163 1044
rect 167 1040 683 1044
rect 687 1040 688 1044
rect 162 1039 168 1040
rect 682 1039 688 1040
rect 958 1044 964 1045
rect 1474 1044 1480 1045
rect 958 1040 959 1044
rect 963 1040 1475 1044
rect 1479 1040 1480 1044
rect 958 1039 964 1040
rect 1474 1039 1480 1040
rect 96 1021 97 1027
rect 103 1026 1847 1027
rect 103 1022 111 1026
rect 115 1022 143 1026
rect 147 1022 151 1026
rect 155 1022 287 1026
rect 291 1022 295 1026
rect 299 1022 455 1026
rect 459 1022 471 1026
rect 475 1022 623 1026
rect 627 1022 663 1026
rect 667 1022 791 1026
rect 795 1022 847 1026
rect 851 1022 951 1026
rect 955 1022 1031 1026
rect 1035 1022 1111 1026
rect 1115 1022 1207 1026
rect 1211 1022 1263 1026
rect 1267 1022 1375 1026
rect 1379 1022 1415 1026
rect 1419 1022 1543 1026
rect 1547 1022 1567 1026
rect 1571 1022 1711 1026
rect 1715 1022 1823 1026
rect 1827 1022 1847 1026
rect 103 1021 1847 1022
rect 1853 1026 3618 1027
rect 1853 1022 1863 1026
rect 1867 1022 1903 1026
rect 1907 1022 1975 1026
rect 1979 1022 2055 1026
rect 2059 1022 2095 1026
rect 2099 1022 2223 1026
rect 2227 1022 2359 1026
rect 2363 1022 2399 1026
rect 2403 1022 2495 1026
rect 2499 1022 2575 1026
rect 2579 1022 2639 1026
rect 2643 1022 2743 1026
rect 2747 1022 2791 1026
rect 2795 1022 2903 1026
rect 2907 1022 2959 1026
rect 2963 1022 3055 1026
rect 3059 1022 3135 1026
rect 3139 1022 3207 1026
rect 3211 1022 3311 1026
rect 3315 1022 3359 1026
rect 3363 1022 3487 1026
rect 3491 1022 3575 1026
rect 3579 1022 3618 1026
rect 1853 1021 3618 1022
rect 246 996 252 997
rect 770 996 776 997
rect 246 992 247 996
rect 251 992 771 996
rect 775 992 776 996
rect 246 991 252 992
rect 770 991 776 992
rect 1118 996 1124 997
rect 1458 996 1464 997
rect 1118 992 1119 996
rect 1123 992 1459 996
rect 1463 992 1464 996
rect 1118 991 1124 992
rect 1458 991 1464 992
rect 84 949 85 955
rect 91 954 1835 955
rect 91 950 111 954
rect 115 950 135 954
rect 139 950 279 954
rect 283 950 287 954
rect 291 950 463 954
rect 467 950 471 954
rect 475 950 655 954
rect 659 950 663 954
rect 667 950 839 954
rect 843 950 855 954
rect 859 950 1023 954
rect 1027 950 1047 954
rect 1051 950 1199 954
rect 1203 950 1223 954
rect 1227 950 1367 954
rect 1371 950 1399 954
rect 1403 950 1535 954
rect 1539 950 1575 954
rect 1579 950 1703 954
rect 1707 950 1727 954
rect 1731 950 1823 954
rect 1827 950 1835 954
rect 91 949 1835 950
rect 1841 954 3606 955
rect 1841 950 1863 954
rect 1867 950 1967 954
rect 1971 950 2087 954
rect 2091 950 2143 954
rect 2147 950 2215 954
rect 2219 950 2231 954
rect 2235 950 2319 954
rect 2323 950 2351 954
rect 2355 950 2407 954
rect 2411 950 2487 954
rect 2491 950 2503 954
rect 2507 950 2615 954
rect 2619 950 2631 954
rect 2635 950 2751 954
rect 2755 950 2783 954
rect 2787 950 2903 954
rect 2907 950 2951 954
rect 2955 950 3079 954
rect 3083 950 3127 954
rect 3131 950 3263 954
rect 3267 950 3303 954
rect 3307 950 3455 954
rect 3459 950 3479 954
rect 3483 950 3575 954
rect 3579 950 3606 954
rect 1841 949 3606 950
rect 302 900 308 901
rect 798 900 804 901
rect 302 896 303 900
rect 307 896 799 900
rect 803 896 804 900
rect 302 895 308 896
rect 798 895 804 896
rect 96 877 97 883
rect 103 882 1847 883
rect 103 878 111 882
rect 115 878 143 882
rect 147 878 287 882
rect 291 878 295 882
rect 299 878 471 882
rect 475 878 479 882
rect 483 878 655 882
rect 659 878 671 882
rect 675 878 839 882
rect 843 878 863 882
rect 867 878 1023 882
rect 1027 878 1055 882
rect 1059 878 1191 882
rect 1195 878 1231 882
rect 1235 878 1359 882
rect 1363 878 1407 882
rect 1411 878 1527 882
rect 1531 878 1583 882
rect 1587 878 1695 882
rect 1699 878 1735 882
rect 1739 878 1823 882
rect 1827 878 1847 882
rect 103 877 1847 878
rect 1853 882 3618 883
rect 1853 878 1863 882
rect 1867 878 2103 882
rect 2107 878 2151 882
rect 2155 878 2191 882
rect 2195 878 2239 882
rect 2243 878 2279 882
rect 2283 878 2327 882
rect 2331 878 2367 882
rect 2371 878 2415 882
rect 2419 878 2455 882
rect 2459 878 2511 882
rect 2515 878 2567 882
rect 2571 878 2623 882
rect 2627 878 2703 882
rect 2707 878 2759 882
rect 2763 878 2871 882
rect 2875 878 2911 882
rect 2915 878 3055 882
rect 3059 878 3087 882
rect 3091 878 3255 882
rect 3259 878 3271 882
rect 3275 878 3463 882
rect 3467 878 3575 882
rect 3579 878 3618 882
rect 1853 877 3618 878
rect 1206 860 1212 861
rect 1626 860 1632 861
rect 1206 856 1207 860
rect 1211 856 1627 860
rect 1631 856 1632 860
rect 1206 855 1212 856
rect 1626 855 1632 856
rect 1086 828 1092 829
rect 1398 828 1404 829
rect 1086 824 1087 828
rect 1091 824 1399 828
rect 1403 824 1404 828
rect 1086 823 1092 824
rect 1398 823 1404 824
rect 84 809 85 815
rect 91 814 1835 815
rect 91 810 111 814
rect 115 810 135 814
rect 139 810 271 814
rect 275 810 279 814
rect 283 810 423 814
rect 427 810 463 814
rect 467 810 583 814
rect 587 810 647 814
rect 651 810 743 814
rect 747 810 831 814
rect 835 810 895 814
rect 899 810 1015 814
rect 1019 810 1039 814
rect 1043 810 1183 814
rect 1187 810 1327 814
rect 1331 810 1351 814
rect 1355 810 1479 814
rect 1483 810 1519 814
rect 1523 810 1687 814
rect 1691 810 1823 814
rect 1827 810 1835 814
rect 91 809 1835 810
rect 1841 814 3606 815
rect 1841 810 1863 814
rect 1867 810 2095 814
rect 2099 810 2183 814
rect 2187 810 2199 814
rect 2203 810 2271 814
rect 2275 810 2287 814
rect 2291 810 2359 814
rect 2363 810 2375 814
rect 2379 810 2447 814
rect 2451 810 2463 814
rect 2467 810 2551 814
rect 2555 810 2559 814
rect 2563 810 2655 814
rect 2659 810 2695 814
rect 2699 810 2783 814
rect 2787 810 2863 814
rect 2867 810 2935 814
rect 2939 810 3047 814
rect 3051 810 3111 814
rect 3115 810 3247 814
rect 3251 810 3295 814
rect 3299 810 3455 814
rect 3459 810 3479 814
rect 3483 810 3575 814
rect 3579 810 3606 814
rect 1841 809 3606 810
rect 154 796 160 797
rect 750 796 756 797
rect 154 792 155 796
rect 159 792 751 796
rect 755 792 756 796
rect 154 791 160 792
rect 750 791 756 792
rect 2706 772 2712 773
rect 3198 772 3204 773
rect 2706 768 2707 772
rect 2711 768 3199 772
rect 3203 768 3204 772
rect 2706 767 2712 768
rect 3198 767 3204 768
rect 370 756 376 757
rect 678 756 684 757
rect 370 752 371 756
rect 375 752 679 756
rect 683 752 684 756
rect 370 751 376 752
rect 678 751 684 752
rect 2674 756 2680 757
rect 3138 756 3144 757
rect 2674 752 2675 756
rect 2679 752 3139 756
rect 3143 752 3144 756
rect 2674 751 2680 752
rect 3138 751 3144 752
rect 96 737 97 743
rect 103 742 1847 743
rect 103 738 111 742
rect 115 738 143 742
rect 147 738 279 742
rect 283 738 359 742
rect 363 738 431 742
rect 435 738 447 742
rect 451 738 543 742
rect 547 738 591 742
rect 595 738 639 742
rect 643 738 735 742
rect 739 738 751 742
rect 755 738 831 742
rect 835 738 903 742
rect 907 738 927 742
rect 931 738 1031 742
rect 1035 738 1047 742
rect 1051 738 1135 742
rect 1139 738 1191 742
rect 1195 738 1239 742
rect 1243 738 1335 742
rect 1339 738 1487 742
rect 1491 738 1823 742
rect 1827 738 1847 742
rect 103 737 1847 738
rect 1853 742 3618 743
rect 1853 738 1863 742
rect 1867 738 1943 742
rect 1947 738 2103 742
rect 2107 738 2207 742
rect 2211 738 2255 742
rect 2259 738 2295 742
rect 2299 738 2383 742
rect 2387 738 2407 742
rect 2411 738 2471 742
rect 2475 738 2551 742
rect 2555 738 2559 742
rect 2563 738 2663 742
rect 2667 738 2695 742
rect 2699 738 2791 742
rect 2795 738 2839 742
rect 2843 738 2943 742
rect 2947 738 2983 742
rect 2987 738 3119 742
rect 3123 738 3135 742
rect 3139 738 3287 742
rect 3291 738 3303 742
rect 3307 738 3439 742
rect 3443 738 3487 742
rect 3491 738 3575 742
rect 3579 738 3618 742
rect 1853 737 3618 738
rect 1022 732 1028 733
rect 1202 732 1208 733
rect 1022 728 1023 732
rect 1027 728 1203 732
rect 1207 728 1208 732
rect 1022 727 1028 728
rect 1202 727 1208 728
rect 84 665 85 671
rect 91 670 1835 671
rect 91 666 111 670
rect 115 666 351 670
rect 355 666 439 670
rect 443 666 479 670
rect 483 666 535 670
rect 539 666 567 670
rect 571 666 631 670
rect 635 666 655 670
rect 659 666 727 670
rect 731 666 743 670
rect 747 666 823 670
rect 827 666 831 670
rect 835 666 919 670
rect 923 666 1007 670
rect 1011 666 1023 670
rect 1027 666 1095 670
rect 1099 666 1127 670
rect 1131 666 1183 670
rect 1187 666 1231 670
rect 1235 666 1271 670
rect 1275 666 1823 670
rect 1827 666 1835 670
rect 91 665 1835 666
rect 1841 670 3606 671
rect 1841 666 1863 670
rect 1867 666 1887 670
rect 1891 666 1935 670
rect 1939 666 2023 670
rect 2027 666 2095 670
rect 2099 666 2199 670
rect 2203 666 2247 670
rect 2251 666 2383 670
rect 2387 666 2399 670
rect 2403 666 2543 670
rect 2547 666 2567 670
rect 2571 666 2687 670
rect 2691 666 2743 670
rect 2747 666 2831 670
rect 2835 666 2911 670
rect 2915 666 2975 670
rect 2979 666 3063 670
rect 3067 666 3127 670
rect 3131 666 3207 670
rect 3211 666 3279 670
rect 3283 666 3351 670
rect 3355 666 3431 670
rect 3435 666 3479 670
rect 3483 666 3575 670
rect 3579 666 3606 670
rect 1841 665 3606 666
rect 2762 612 2768 613
rect 3078 612 3084 613
rect 2762 608 2763 612
rect 2767 608 3079 612
rect 3083 608 3084 612
rect 2762 607 2768 608
rect 3078 607 3084 608
rect 96 597 97 603
rect 103 602 1847 603
rect 103 598 111 602
rect 115 598 487 602
rect 491 598 503 602
rect 507 598 575 602
rect 579 598 599 602
rect 603 598 663 602
rect 667 598 703 602
rect 707 598 751 602
rect 755 598 815 602
rect 819 598 839 602
rect 843 598 927 602
rect 931 598 935 602
rect 939 598 1015 602
rect 1019 598 1063 602
rect 1067 598 1103 602
rect 1107 598 1191 602
rect 1195 598 1279 602
rect 1283 598 1327 602
rect 1331 598 1471 602
rect 1475 598 1615 602
rect 1619 598 1735 602
rect 1739 598 1823 602
rect 1827 598 1847 602
rect 103 597 1847 598
rect 1853 602 3618 603
rect 1853 598 1863 602
rect 1867 598 1895 602
rect 1899 598 2031 602
rect 2035 598 2087 602
rect 2091 598 2207 602
rect 2211 598 2303 602
rect 2307 598 2391 602
rect 2395 598 2511 602
rect 2515 598 2575 602
rect 2579 598 2703 602
rect 2707 598 2751 602
rect 2755 598 2879 602
rect 2883 598 2919 602
rect 2923 598 3039 602
rect 3043 598 3071 602
rect 3075 598 3199 602
rect 3203 598 3215 602
rect 3219 598 3351 602
rect 3355 598 3359 602
rect 3363 598 3487 602
rect 3491 598 3575 602
rect 3579 598 3618 602
rect 1853 597 3618 598
rect 558 572 564 573
rect 770 572 776 573
rect 558 568 559 572
rect 563 568 771 572
rect 775 568 776 572
rect 558 567 564 568
rect 770 567 776 568
rect 84 529 85 535
rect 91 534 1835 535
rect 91 530 111 534
rect 115 530 159 534
rect 163 530 303 534
rect 307 530 463 534
rect 467 530 495 534
rect 499 530 591 534
rect 595 530 631 534
rect 635 530 695 534
rect 699 530 799 534
rect 803 530 807 534
rect 811 530 927 534
rect 931 530 959 534
rect 963 530 1055 534
rect 1059 530 1103 534
rect 1107 530 1183 534
rect 1187 530 1239 534
rect 1243 530 1319 534
rect 1323 530 1367 534
rect 1371 530 1463 534
rect 1467 530 1495 534
rect 1499 530 1607 534
rect 1611 530 1623 534
rect 1627 530 1727 534
rect 1731 530 1823 534
rect 1827 530 1835 534
rect 91 529 1835 530
rect 1841 529 1842 535
rect 1834 527 1842 529
rect 1834 521 1835 527
rect 1841 526 3599 527
rect 1841 522 1863 526
rect 1867 522 1887 526
rect 1891 522 2079 526
rect 2083 522 2287 526
rect 2291 522 2295 526
rect 2299 522 2487 526
rect 2491 522 2503 526
rect 2507 522 2671 526
rect 2675 522 2695 526
rect 2699 522 2847 526
rect 2851 522 2871 526
rect 2875 522 3015 526
rect 3019 522 3031 526
rect 3035 522 3175 526
rect 3179 522 3191 526
rect 3195 522 3335 526
rect 3339 522 3343 526
rect 3347 522 3479 526
rect 3483 522 3575 526
rect 3579 522 3599 526
rect 1841 521 3599 522
rect 3605 521 3606 527
rect 2094 468 2100 469
rect 2418 468 2424 469
rect 2094 464 2095 468
rect 2099 464 2419 468
rect 2423 464 2424 468
rect 2094 463 2100 464
rect 2418 463 2424 464
rect 2686 468 2692 469
rect 3082 468 3088 469
rect 2686 464 2687 468
rect 2691 464 3083 468
rect 3087 464 3088 468
rect 2686 463 2692 464
rect 3082 463 3088 464
rect 96 453 97 459
rect 103 458 1847 459
rect 103 454 111 458
rect 115 454 143 458
rect 147 454 167 458
rect 171 454 271 458
rect 275 454 311 458
rect 315 454 439 458
rect 443 454 471 458
rect 475 454 615 458
rect 619 454 639 458
rect 643 454 791 458
rect 795 454 807 458
rect 811 454 967 458
rect 971 454 1111 458
rect 1115 454 1127 458
rect 1131 454 1247 458
rect 1251 454 1287 458
rect 1291 454 1375 458
rect 1379 454 1447 458
rect 1451 454 1503 458
rect 1507 454 1607 458
rect 1611 454 1631 458
rect 1635 454 1735 458
rect 1739 454 1823 458
rect 1827 454 1847 458
rect 103 453 1847 454
rect 1853 458 3618 459
rect 1853 454 1863 458
rect 1867 454 2087 458
rect 2091 454 2247 458
rect 2251 454 2295 458
rect 2299 454 2335 458
rect 2339 454 2431 458
rect 2435 454 2495 458
rect 2499 454 2527 458
rect 2531 454 2623 458
rect 2627 454 2679 458
rect 2683 454 2735 458
rect 2739 454 2855 458
rect 2859 454 2863 458
rect 2867 454 3007 458
rect 3011 454 3023 458
rect 3027 454 3167 458
rect 3171 454 3183 458
rect 3187 454 3335 458
rect 3339 454 3343 458
rect 3347 454 3487 458
rect 3491 454 3575 458
rect 3579 454 3618 458
rect 1853 453 3618 454
rect 2302 444 2308 445
rect 2594 444 2600 445
rect 2302 440 2303 444
rect 2307 440 2595 444
rect 2599 440 2600 444
rect 2302 439 2308 440
rect 2594 439 2600 440
rect 1238 436 1244 437
rect 1546 436 1552 437
rect 1238 432 1239 436
rect 1243 432 1547 436
rect 1551 432 1552 436
rect 1238 431 1244 432
rect 1546 431 1552 432
rect 84 385 85 391
rect 91 390 1835 391
rect 91 386 111 390
rect 115 386 135 390
rect 139 386 263 390
rect 267 386 431 390
rect 435 386 607 390
rect 611 386 783 390
rect 787 386 951 390
rect 955 386 959 390
rect 963 386 1111 390
rect 1115 386 1119 390
rect 1123 386 1271 390
rect 1275 386 1279 390
rect 1283 386 1431 390
rect 1435 386 1439 390
rect 1443 386 1591 390
rect 1595 386 1599 390
rect 1603 386 1823 390
rect 1827 386 1835 390
rect 91 385 1835 386
rect 1841 390 3606 391
rect 1841 386 1863 390
rect 1867 386 2151 390
rect 2155 386 2239 390
rect 2243 386 2327 390
rect 2331 386 2415 390
rect 2419 386 2423 390
rect 2427 386 2503 390
rect 2507 386 2519 390
rect 2523 386 2615 390
rect 2619 386 2727 390
rect 2731 386 2751 390
rect 2755 386 2855 390
rect 2859 386 2919 390
rect 2923 386 2999 390
rect 3003 386 3103 390
rect 3107 386 3159 390
rect 3163 386 3303 390
rect 3307 386 3327 390
rect 3331 386 3479 390
rect 3483 386 3575 390
rect 3579 386 3606 390
rect 1841 385 3606 386
rect 154 372 160 373
rect 682 372 688 373
rect 154 368 155 372
rect 159 368 683 372
rect 687 368 688 372
rect 154 367 160 368
rect 682 367 688 368
rect 350 332 356 333
rect 690 332 696 333
rect 350 328 351 332
rect 355 328 691 332
rect 695 328 696 332
rect 350 327 356 328
rect 690 327 696 328
rect 2770 332 2776 333
rect 3198 332 3204 333
rect 2770 328 2771 332
rect 2775 328 3199 332
rect 3203 328 3204 332
rect 2770 327 2776 328
rect 3198 327 3204 328
rect 1846 322 3618 323
rect 1846 319 1863 322
rect 96 313 97 319
rect 103 318 1847 319
rect 103 314 111 318
rect 115 314 143 318
rect 147 314 263 318
rect 267 314 271 318
rect 275 314 391 318
rect 395 314 439 318
rect 443 314 527 318
rect 531 314 615 318
rect 619 314 679 318
rect 683 314 791 318
rect 795 314 839 318
rect 843 314 959 318
rect 963 314 1007 318
rect 1011 314 1119 318
rect 1123 314 1175 318
rect 1179 314 1279 318
rect 1283 314 1343 318
rect 1347 314 1439 318
rect 1443 314 1511 318
rect 1515 314 1599 318
rect 1603 314 1687 318
rect 1691 314 1823 318
rect 1827 314 1847 318
rect 103 313 1847 314
rect 1853 318 1863 319
rect 1867 318 2023 322
rect 2027 318 2119 322
rect 2123 318 2159 322
rect 2163 318 2223 322
rect 2227 318 2247 322
rect 2251 318 2327 322
rect 2331 318 2335 322
rect 2339 318 2423 322
rect 2427 318 2431 322
rect 2435 318 2511 322
rect 2515 318 2535 322
rect 2539 318 2623 322
rect 2627 318 2639 322
rect 2643 318 2743 322
rect 2747 318 2759 322
rect 2763 318 2855 322
rect 2859 318 2927 322
rect 2931 318 2967 322
rect 2971 318 3111 322
rect 3115 318 3311 322
rect 3315 318 3487 322
rect 3491 318 3575 322
rect 3579 318 3618 322
rect 1853 317 3618 318
rect 1853 313 1854 317
rect 2214 292 2220 293
rect 2398 292 2404 293
rect 2214 288 2215 292
rect 2219 288 2399 292
rect 2403 288 2404 292
rect 2214 287 2220 288
rect 2398 287 2404 288
rect 1834 249 1835 255
rect 1841 254 3599 255
rect 1841 250 1863 254
rect 1867 250 1959 254
rect 1963 250 2015 254
rect 2019 250 2111 254
rect 2115 250 2175 254
rect 2179 250 2215 254
rect 2219 250 2319 254
rect 2323 250 2383 254
rect 2387 250 2423 254
rect 2427 250 2527 254
rect 2531 250 2583 254
rect 2587 250 2631 254
rect 2635 250 2735 254
rect 2739 250 2767 254
rect 2771 250 2847 254
rect 2851 250 2951 254
rect 2955 250 2959 254
rect 2963 250 3127 254
rect 3131 250 3311 254
rect 3315 250 3479 254
rect 3483 250 3575 254
rect 3579 250 3599 254
rect 1841 249 3599 250
rect 3605 249 3606 255
rect 1834 247 1842 249
rect 84 241 85 247
rect 91 246 1835 247
rect 91 242 111 246
rect 115 242 255 246
rect 259 242 383 246
rect 387 242 399 246
rect 403 242 503 246
rect 507 242 519 246
rect 523 242 615 246
rect 619 242 671 246
rect 675 242 735 246
rect 739 242 831 246
rect 835 242 863 246
rect 867 242 991 246
rect 995 242 999 246
rect 1003 242 1119 246
rect 1123 242 1167 246
rect 1171 242 1247 246
rect 1251 242 1335 246
rect 1339 242 1375 246
rect 1379 242 1495 246
rect 1499 242 1503 246
rect 1507 242 1623 246
rect 1627 242 1679 246
rect 1683 242 1727 246
rect 1731 242 1823 246
rect 1827 242 1835 246
rect 91 241 1835 242
rect 1841 241 1842 247
rect 2602 196 2608 197
rect 2922 196 2928 197
rect 2602 192 2603 196
rect 2607 192 2923 196
rect 2927 192 2928 196
rect 2602 191 2608 192
rect 2922 191 2928 192
rect 418 188 424 189
rect 810 188 816 189
rect 418 184 419 188
rect 423 184 811 188
rect 815 184 816 188
rect 418 183 424 184
rect 810 183 816 184
rect 2618 164 2624 165
rect 3198 164 3204 165
rect 2618 160 2619 164
rect 2623 160 3199 164
rect 3203 160 3204 164
rect 2618 159 2624 160
rect 3198 159 3204 160
rect 96 153 97 159
rect 103 158 1847 159
rect 103 154 111 158
rect 115 154 223 158
rect 227 154 311 158
rect 315 154 399 158
rect 403 154 407 158
rect 411 154 487 158
rect 491 154 511 158
rect 515 154 575 158
rect 579 154 623 158
rect 627 154 663 158
rect 667 154 743 158
rect 747 154 751 158
rect 755 154 839 158
rect 843 154 871 158
rect 875 154 927 158
rect 931 154 999 158
rect 1003 154 1015 158
rect 1019 154 1103 158
rect 1107 154 1127 158
rect 1131 154 1191 158
rect 1195 154 1255 158
rect 1259 154 1295 158
rect 1299 154 1383 158
rect 1387 154 1399 158
rect 1403 154 1503 158
rect 1507 154 1511 158
rect 1515 154 1631 158
rect 1635 154 1735 158
rect 1739 154 1823 158
rect 1827 154 1847 158
rect 103 153 1847 154
rect 1853 155 1854 159
rect 1853 154 3618 155
rect 1853 153 1863 154
rect 1846 150 1863 153
rect 1867 150 1895 154
rect 1899 150 1967 154
rect 1971 150 1983 154
rect 1987 150 2071 154
rect 2075 150 2159 154
rect 2163 150 2183 154
rect 2187 150 2271 154
rect 2275 150 2383 154
rect 2387 150 2391 154
rect 2395 150 2495 154
rect 2499 150 2591 154
rect 2595 150 2607 154
rect 2611 150 2719 154
rect 2723 150 2775 154
rect 2779 150 2823 154
rect 2827 150 2927 154
rect 2931 150 2959 154
rect 2963 150 3023 154
rect 3027 150 3119 154
rect 3123 150 3135 154
rect 3139 150 3215 154
rect 3219 150 3311 154
rect 3315 150 3319 154
rect 3323 150 3399 154
rect 3403 150 3487 154
rect 3491 150 3575 154
rect 3579 150 3618 154
rect 1846 149 3618 150
rect 84 85 85 91
rect 91 90 1835 91
rect 91 86 111 90
rect 115 86 215 90
rect 219 86 303 90
rect 307 86 391 90
rect 395 86 479 90
rect 483 86 567 90
rect 571 86 655 90
rect 659 86 743 90
rect 747 86 831 90
rect 835 86 919 90
rect 923 86 1007 90
rect 1011 86 1095 90
rect 1099 86 1183 90
rect 1187 86 1287 90
rect 1291 86 1391 90
rect 1395 86 1503 90
rect 1507 86 1623 90
rect 1627 86 1727 90
rect 1731 86 1823 90
rect 1827 86 1835 90
rect 91 85 1835 86
rect 1841 87 1842 91
rect 1841 86 3606 87
rect 1841 85 1863 86
rect 1834 82 1863 85
rect 1867 82 1887 86
rect 1891 82 1975 86
rect 1979 82 2063 86
rect 2067 82 2151 86
rect 2155 82 2263 86
rect 2267 82 2375 86
rect 2379 82 2487 86
rect 2491 82 2599 86
rect 2603 82 2711 86
rect 2715 82 2815 86
rect 2819 82 2919 86
rect 2923 82 3015 86
rect 3019 82 3111 86
rect 3115 82 3207 86
rect 3211 82 3303 86
rect 3307 82 3391 86
rect 3395 82 3479 86
rect 3483 82 3575 86
rect 3579 82 3606 86
rect 1834 81 3606 82
<< m5c >>
rect 97 3645 103 3651
rect 1847 3645 1853 3651
rect 85 3569 91 3575
rect 1835 3569 1841 3575
rect 97 3501 103 3507
rect 1847 3501 1853 3507
rect 85 3433 91 3439
rect 1835 3433 1841 3439
rect 97 3357 103 3363
rect 1847 3357 1853 3363
rect 1835 3293 1841 3299
rect 3599 3293 3605 3299
rect 85 3285 91 3291
rect 1835 3285 1841 3291
rect 1847 3217 1853 3223
rect 3611 3217 3617 3223
rect 97 3205 103 3211
rect 1847 3205 1853 3211
rect 1835 3145 1841 3151
rect 3599 3145 3605 3151
rect 85 3125 91 3131
rect 1835 3125 1841 3131
rect 1847 3073 1853 3079
rect 3611 3073 3617 3079
rect 97 3057 103 3063
rect 1847 3057 1853 3063
rect 1835 2993 1841 2999
rect 3599 2993 3605 2999
rect 85 2977 91 2983
rect 1835 2977 1841 2983
rect 1847 2917 1853 2923
rect 3611 2917 3617 2923
rect 97 2909 103 2915
rect 1847 2909 1853 2915
rect 1835 2849 1841 2855
rect 3599 2849 3605 2855
rect 85 2837 91 2843
rect 1835 2837 1841 2843
rect 1847 2781 1853 2787
rect 3611 2781 3617 2787
rect 97 2761 103 2767
rect 1847 2761 1853 2767
rect 1835 2713 1841 2719
rect 3599 2713 3605 2719
rect 85 2689 91 2695
rect 1835 2689 1841 2695
rect 1847 2625 1853 2631
rect 3611 2625 3617 2631
rect 97 2617 103 2623
rect 1847 2617 1853 2623
rect 1835 2557 1841 2563
rect 3599 2557 3605 2563
rect 85 2541 91 2547
rect 1835 2541 1841 2547
rect 1847 2485 1853 2491
rect 3611 2485 3617 2491
rect 97 2469 103 2475
rect 1847 2469 1853 2475
rect 1835 2413 1841 2419
rect 3599 2413 3605 2419
rect 85 2397 91 2403
rect 1835 2397 1841 2403
rect 1847 2337 1853 2343
rect 3611 2337 3617 2343
rect 97 2325 103 2331
rect 1847 2325 1853 2331
rect 1835 2265 1841 2271
rect 3599 2265 3605 2271
rect 85 2249 91 2255
rect 1835 2249 1841 2255
rect 1847 2193 1853 2199
rect 3611 2193 3617 2199
rect 97 2177 103 2183
rect 1847 2177 1853 2183
rect 1835 2121 1841 2127
rect 3599 2121 3605 2127
rect 85 2101 91 2107
rect 1835 2101 1841 2107
rect 1847 2045 1853 2051
rect 3611 2045 3617 2051
rect 97 2025 103 2031
rect 1847 2025 1853 2031
rect 1835 1973 1841 1979
rect 3599 1973 3605 1979
rect 85 1949 91 1955
rect 1835 1949 1841 1955
rect 1847 1897 1853 1903
rect 3611 1897 3617 1903
rect 97 1873 103 1879
rect 1847 1873 1853 1879
rect 1835 1825 1841 1831
rect 3599 1825 3605 1831
rect 85 1797 91 1803
rect 1835 1797 1841 1803
rect 1847 1749 1853 1755
rect 3611 1749 3617 1755
rect 97 1729 103 1735
rect 1847 1729 1853 1735
rect 1835 1677 1841 1683
rect 3599 1677 3605 1683
rect 85 1661 91 1667
rect 1835 1661 1841 1667
rect 1847 1609 1853 1615
rect 3611 1609 3617 1615
rect 97 1589 103 1595
rect 1847 1589 1853 1595
rect 1835 1533 1841 1539
rect 3599 1533 3605 1539
rect 85 1517 91 1523
rect 1835 1517 1841 1523
rect 1847 1461 1853 1467
rect 3611 1461 3617 1467
rect 97 1445 103 1451
rect 1847 1445 1853 1451
rect 85 1377 91 1383
rect 1835 1377 1841 1383
rect 97 1309 103 1315
rect 1847 1309 1853 1315
rect 85 1241 91 1247
rect 1835 1241 1841 1247
rect 97 1165 103 1171
rect 1847 1165 1853 1171
rect 85 1093 91 1099
rect 1835 1093 1841 1099
rect 97 1021 103 1027
rect 1847 1021 1853 1027
rect 85 949 91 955
rect 1835 949 1841 955
rect 97 877 103 883
rect 1847 877 1853 883
rect 85 809 91 815
rect 1835 809 1841 815
rect 97 737 103 743
rect 1847 737 1853 743
rect 85 665 91 671
rect 1835 665 1841 671
rect 97 597 103 603
rect 1847 597 1853 603
rect 85 529 91 535
rect 1835 529 1841 535
rect 1835 521 1841 527
rect 3599 521 3605 527
rect 97 453 103 459
rect 1847 453 1853 459
rect 85 385 91 391
rect 1835 385 1841 391
rect 97 313 103 319
rect 1847 313 1853 319
rect 1835 249 1841 255
rect 3599 249 3605 255
rect 85 241 91 247
rect 1835 241 1841 247
rect 97 153 103 159
rect 1847 153 1853 159
rect 85 85 91 91
rect 1835 85 1841 91
<< m5 >>
rect 84 3575 92 3672
rect 84 3569 85 3575
rect 91 3569 92 3575
rect 84 3439 92 3569
rect 84 3433 85 3439
rect 91 3433 92 3439
rect 84 3291 92 3433
rect 84 3285 85 3291
rect 91 3285 92 3291
rect 84 3131 92 3285
rect 84 3125 85 3131
rect 91 3125 92 3131
rect 84 2983 92 3125
rect 84 2977 85 2983
rect 91 2977 92 2983
rect 84 2843 92 2977
rect 84 2837 85 2843
rect 91 2837 92 2843
rect 84 2695 92 2837
rect 84 2689 85 2695
rect 91 2689 92 2695
rect 84 2547 92 2689
rect 84 2541 85 2547
rect 91 2541 92 2547
rect 84 2403 92 2541
rect 84 2397 85 2403
rect 91 2397 92 2403
rect 84 2255 92 2397
rect 84 2249 85 2255
rect 91 2249 92 2255
rect 84 2107 92 2249
rect 84 2101 85 2107
rect 91 2101 92 2107
rect 84 1955 92 2101
rect 84 1949 85 1955
rect 91 1949 92 1955
rect 84 1803 92 1949
rect 84 1797 85 1803
rect 91 1797 92 1803
rect 84 1667 92 1797
rect 84 1661 85 1667
rect 91 1661 92 1667
rect 84 1523 92 1661
rect 84 1517 85 1523
rect 91 1517 92 1523
rect 84 1383 92 1517
rect 84 1377 85 1383
rect 91 1377 92 1383
rect 84 1247 92 1377
rect 84 1241 85 1247
rect 91 1241 92 1247
rect 84 1099 92 1241
rect 84 1093 85 1099
rect 91 1093 92 1099
rect 84 955 92 1093
rect 84 949 85 955
rect 91 949 92 955
rect 84 815 92 949
rect 84 809 85 815
rect 91 809 92 815
rect 84 671 92 809
rect 84 665 85 671
rect 91 665 92 671
rect 84 535 92 665
rect 84 529 85 535
rect 91 529 92 535
rect 84 391 92 529
rect 84 385 85 391
rect 91 385 92 391
rect 84 247 92 385
rect 84 241 85 247
rect 91 241 92 247
rect 84 91 92 241
rect 84 85 85 91
rect 91 85 92 91
rect 84 72 92 85
rect 96 3651 104 3672
rect 96 3645 97 3651
rect 103 3645 104 3651
rect 96 3507 104 3645
rect 96 3501 97 3507
rect 103 3501 104 3507
rect 96 3363 104 3501
rect 96 3357 97 3363
rect 103 3357 104 3363
rect 96 3211 104 3357
rect 96 3205 97 3211
rect 103 3205 104 3211
rect 96 3063 104 3205
rect 96 3057 97 3063
rect 103 3057 104 3063
rect 96 2915 104 3057
rect 96 2909 97 2915
rect 103 2909 104 2915
rect 96 2767 104 2909
rect 96 2761 97 2767
rect 103 2761 104 2767
rect 96 2623 104 2761
rect 96 2617 97 2623
rect 103 2617 104 2623
rect 96 2475 104 2617
rect 96 2469 97 2475
rect 103 2469 104 2475
rect 96 2331 104 2469
rect 96 2325 97 2331
rect 103 2325 104 2331
rect 96 2183 104 2325
rect 96 2177 97 2183
rect 103 2177 104 2183
rect 96 2031 104 2177
rect 96 2025 97 2031
rect 103 2025 104 2031
rect 96 1879 104 2025
rect 96 1873 97 1879
rect 103 1873 104 1879
rect 96 1735 104 1873
rect 96 1729 97 1735
rect 103 1729 104 1735
rect 96 1595 104 1729
rect 96 1589 97 1595
rect 103 1589 104 1595
rect 96 1451 104 1589
rect 96 1445 97 1451
rect 103 1445 104 1451
rect 96 1315 104 1445
rect 96 1309 97 1315
rect 103 1309 104 1315
rect 96 1171 104 1309
rect 96 1165 97 1171
rect 103 1165 104 1171
rect 96 1027 104 1165
rect 96 1021 97 1027
rect 103 1021 104 1027
rect 96 883 104 1021
rect 96 877 97 883
rect 103 877 104 883
rect 96 743 104 877
rect 96 737 97 743
rect 103 737 104 743
rect 96 603 104 737
rect 96 597 97 603
rect 103 597 104 603
rect 96 459 104 597
rect 96 453 97 459
rect 103 453 104 459
rect 96 319 104 453
rect 96 313 97 319
rect 103 313 104 319
rect 96 159 104 313
rect 96 153 97 159
rect 103 153 104 159
rect 96 72 104 153
rect 1834 3575 1842 3672
rect 1834 3569 1835 3575
rect 1841 3569 1842 3575
rect 1834 3439 1842 3569
rect 1834 3433 1835 3439
rect 1841 3433 1842 3439
rect 1834 3299 1842 3433
rect 1834 3293 1835 3299
rect 1841 3293 1842 3299
rect 1834 3291 1842 3293
rect 1834 3285 1835 3291
rect 1841 3285 1842 3291
rect 1834 3151 1842 3285
rect 1834 3145 1835 3151
rect 1841 3145 1842 3151
rect 1834 3131 1842 3145
rect 1834 3125 1835 3131
rect 1841 3125 1842 3131
rect 1834 2999 1842 3125
rect 1834 2993 1835 2999
rect 1841 2993 1842 2999
rect 1834 2983 1842 2993
rect 1834 2977 1835 2983
rect 1841 2977 1842 2983
rect 1834 2855 1842 2977
rect 1834 2849 1835 2855
rect 1841 2849 1842 2855
rect 1834 2843 1842 2849
rect 1834 2837 1835 2843
rect 1841 2837 1842 2843
rect 1834 2719 1842 2837
rect 1834 2713 1835 2719
rect 1841 2713 1842 2719
rect 1834 2695 1842 2713
rect 1834 2689 1835 2695
rect 1841 2689 1842 2695
rect 1834 2563 1842 2689
rect 1834 2557 1835 2563
rect 1841 2557 1842 2563
rect 1834 2547 1842 2557
rect 1834 2541 1835 2547
rect 1841 2541 1842 2547
rect 1834 2419 1842 2541
rect 1834 2413 1835 2419
rect 1841 2413 1842 2419
rect 1834 2403 1842 2413
rect 1834 2397 1835 2403
rect 1841 2397 1842 2403
rect 1834 2271 1842 2397
rect 1834 2265 1835 2271
rect 1841 2265 1842 2271
rect 1834 2255 1842 2265
rect 1834 2249 1835 2255
rect 1841 2249 1842 2255
rect 1834 2127 1842 2249
rect 1834 2121 1835 2127
rect 1841 2121 1842 2127
rect 1834 2107 1842 2121
rect 1834 2101 1835 2107
rect 1841 2101 1842 2107
rect 1834 1979 1842 2101
rect 1834 1973 1835 1979
rect 1841 1973 1842 1979
rect 1834 1955 1842 1973
rect 1834 1949 1835 1955
rect 1841 1949 1842 1955
rect 1834 1831 1842 1949
rect 1834 1825 1835 1831
rect 1841 1825 1842 1831
rect 1834 1803 1842 1825
rect 1834 1797 1835 1803
rect 1841 1797 1842 1803
rect 1834 1683 1842 1797
rect 1834 1677 1835 1683
rect 1841 1677 1842 1683
rect 1834 1667 1842 1677
rect 1834 1661 1835 1667
rect 1841 1661 1842 1667
rect 1834 1539 1842 1661
rect 1834 1533 1835 1539
rect 1841 1533 1842 1539
rect 1834 1523 1842 1533
rect 1834 1517 1835 1523
rect 1841 1517 1842 1523
rect 1834 1383 1842 1517
rect 1834 1377 1835 1383
rect 1841 1377 1842 1383
rect 1834 1247 1842 1377
rect 1834 1241 1835 1247
rect 1841 1241 1842 1247
rect 1834 1099 1842 1241
rect 1834 1093 1835 1099
rect 1841 1093 1842 1099
rect 1834 955 1842 1093
rect 1834 949 1835 955
rect 1841 949 1842 955
rect 1834 815 1842 949
rect 1834 809 1835 815
rect 1841 809 1842 815
rect 1834 671 1842 809
rect 1834 665 1835 671
rect 1841 665 1842 671
rect 1834 535 1842 665
rect 1834 529 1835 535
rect 1841 529 1842 535
rect 1834 527 1842 529
rect 1834 521 1835 527
rect 1841 521 1842 527
rect 1834 391 1842 521
rect 1834 385 1835 391
rect 1841 385 1842 391
rect 1834 255 1842 385
rect 1834 249 1835 255
rect 1841 249 1842 255
rect 1834 247 1842 249
rect 1834 241 1835 247
rect 1841 241 1842 247
rect 1834 91 1842 241
rect 1834 85 1835 91
rect 1841 85 1842 91
rect 1834 72 1842 85
rect 1846 3651 1854 3672
rect 1846 3645 1847 3651
rect 1853 3645 1854 3651
rect 1846 3507 1854 3645
rect 1846 3501 1847 3507
rect 1853 3501 1854 3507
rect 1846 3363 1854 3501
rect 1846 3357 1847 3363
rect 1853 3357 1854 3363
rect 1846 3223 1854 3357
rect 1846 3217 1847 3223
rect 1853 3217 1854 3223
rect 1846 3211 1854 3217
rect 1846 3205 1847 3211
rect 1853 3205 1854 3211
rect 1846 3079 1854 3205
rect 1846 3073 1847 3079
rect 1853 3073 1854 3079
rect 1846 3063 1854 3073
rect 1846 3057 1847 3063
rect 1853 3057 1854 3063
rect 1846 2923 1854 3057
rect 1846 2917 1847 2923
rect 1853 2917 1854 2923
rect 1846 2915 1854 2917
rect 1846 2909 1847 2915
rect 1853 2909 1854 2915
rect 1846 2787 1854 2909
rect 1846 2781 1847 2787
rect 1853 2781 1854 2787
rect 1846 2767 1854 2781
rect 1846 2761 1847 2767
rect 1853 2761 1854 2767
rect 1846 2631 1854 2761
rect 1846 2625 1847 2631
rect 1853 2625 1854 2631
rect 1846 2623 1854 2625
rect 1846 2617 1847 2623
rect 1853 2617 1854 2623
rect 1846 2491 1854 2617
rect 1846 2485 1847 2491
rect 1853 2485 1854 2491
rect 1846 2475 1854 2485
rect 1846 2469 1847 2475
rect 1853 2469 1854 2475
rect 1846 2343 1854 2469
rect 1846 2337 1847 2343
rect 1853 2337 1854 2343
rect 1846 2331 1854 2337
rect 1846 2325 1847 2331
rect 1853 2325 1854 2331
rect 1846 2199 1854 2325
rect 1846 2193 1847 2199
rect 1853 2193 1854 2199
rect 1846 2183 1854 2193
rect 1846 2177 1847 2183
rect 1853 2177 1854 2183
rect 1846 2051 1854 2177
rect 1846 2045 1847 2051
rect 1853 2045 1854 2051
rect 1846 2031 1854 2045
rect 1846 2025 1847 2031
rect 1853 2025 1854 2031
rect 1846 1903 1854 2025
rect 1846 1897 1847 1903
rect 1853 1897 1854 1903
rect 1846 1879 1854 1897
rect 1846 1873 1847 1879
rect 1853 1873 1854 1879
rect 1846 1755 1854 1873
rect 1846 1749 1847 1755
rect 1853 1749 1854 1755
rect 1846 1735 1854 1749
rect 1846 1729 1847 1735
rect 1853 1729 1854 1735
rect 1846 1615 1854 1729
rect 1846 1609 1847 1615
rect 1853 1609 1854 1615
rect 1846 1595 1854 1609
rect 1846 1589 1847 1595
rect 1853 1589 1854 1595
rect 1846 1467 1854 1589
rect 1846 1461 1847 1467
rect 1853 1461 1854 1467
rect 1846 1451 1854 1461
rect 1846 1445 1847 1451
rect 1853 1445 1854 1451
rect 1846 1315 1854 1445
rect 1846 1309 1847 1315
rect 1853 1309 1854 1315
rect 1846 1171 1854 1309
rect 1846 1165 1847 1171
rect 1853 1165 1854 1171
rect 1846 1027 1854 1165
rect 1846 1021 1847 1027
rect 1853 1021 1854 1027
rect 1846 883 1854 1021
rect 1846 877 1847 883
rect 1853 877 1854 883
rect 1846 743 1854 877
rect 1846 737 1847 743
rect 1853 737 1854 743
rect 1846 603 1854 737
rect 1846 597 1847 603
rect 1853 597 1854 603
rect 1846 459 1854 597
rect 1846 453 1847 459
rect 1853 453 1854 459
rect 1846 319 1854 453
rect 1846 313 1847 319
rect 1853 313 1854 319
rect 1846 159 1854 313
rect 1846 153 1847 159
rect 1853 153 1854 159
rect 1846 72 1854 153
rect 3598 3299 3606 3672
rect 3598 3293 3599 3299
rect 3605 3293 3606 3299
rect 3598 3151 3606 3293
rect 3598 3145 3599 3151
rect 3605 3145 3606 3151
rect 3598 2999 3606 3145
rect 3598 2993 3599 2999
rect 3605 2993 3606 2999
rect 3598 2855 3606 2993
rect 3598 2849 3599 2855
rect 3605 2849 3606 2855
rect 3598 2719 3606 2849
rect 3598 2713 3599 2719
rect 3605 2713 3606 2719
rect 3598 2563 3606 2713
rect 3598 2557 3599 2563
rect 3605 2557 3606 2563
rect 3598 2419 3606 2557
rect 3598 2413 3599 2419
rect 3605 2413 3606 2419
rect 3598 2271 3606 2413
rect 3598 2265 3599 2271
rect 3605 2265 3606 2271
rect 3598 2127 3606 2265
rect 3598 2121 3599 2127
rect 3605 2121 3606 2127
rect 3598 1979 3606 2121
rect 3598 1973 3599 1979
rect 3605 1973 3606 1979
rect 3598 1831 3606 1973
rect 3598 1825 3599 1831
rect 3605 1825 3606 1831
rect 3598 1683 3606 1825
rect 3598 1677 3599 1683
rect 3605 1677 3606 1683
rect 3598 1539 3606 1677
rect 3598 1533 3599 1539
rect 3605 1533 3606 1539
rect 3598 527 3606 1533
rect 3598 521 3599 527
rect 3605 521 3606 527
rect 3598 255 3606 521
rect 3598 249 3599 255
rect 3605 249 3606 255
rect 3598 72 3606 249
rect 3610 3223 3618 3672
rect 3610 3217 3611 3223
rect 3617 3217 3618 3223
rect 3610 3079 3618 3217
rect 3610 3073 3611 3079
rect 3617 3073 3618 3079
rect 3610 2923 3618 3073
rect 3610 2917 3611 2923
rect 3617 2917 3618 2923
rect 3610 2787 3618 2917
rect 3610 2781 3611 2787
rect 3617 2781 3618 2787
rect 3610 2631 3618 2781
rect 3610 2625 3611 2631
rect 3617 2625 3618 2631
rect 3610 2491 3618 2625
rect 3610 2485 3611 2491
rect 3617 2485 3618 2491
rect 3610 2343 3618 2485
rect 3610 2337 3611 2343
rect 3617 2337 3618 2343
rect 3610 2199 3618 2337
rect 3610 2193 3611 2199
rect 3617 2193 3618 2199
rect 3610 2051 3618 2193
rect 3610 2045 3611 2051
rect 3617 2045 3618 2051
rect 3610 1903 3618 2045
rect 3610 1897 3611 1903
rect 3617 1897 3618 1903
rect 3610 1755 3618 1897
rect 3610 1749 3611 1755
rect 3617 1749 3618 1755
rect 3610 1615 3618 1749
rect 3610 1609 3611 1615
rect 3617 1609 3618 1615
rect 3610 1467 3618 1609
rect 3610 1461 3611 1467
rect 3617 1461 3618 1467
rect 3610 72 3618 1461
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__191
timestamp 1731220617
transform 1 0 3568 0 1 3448
box 7 3 12 24
use welltap_svt  __well_tap__190
timestamp 1731220617
transform 1 0 1856 0 1 3448
box 7 3 12 24
use welltap_svt  __well_tap__189
timestamp 1731220617
transform 1 0 3568 0 -1 3416
box 7 3 12 24
use welltap_svt  __well_tap__188
timestamp 1731220617
transform 1 0 1856 0 -1 3416
box 7 3 12 24
use welltap_svt  __well_tap__187
timestamp 1731220617
transform 1 0 3568 0 1 3312
box 7 3 12 24
use welltap_svt  __well_tap__186
timestamp 1731220617
transform 1 0 1856 0 1 3312
box 7 3 12 24
use welltap_svt  __well_tap__185
timestamp 1731220617
transform 1 0 3568 0 -1 3280
box 7 3 12 24
use welltap_svt  __well_tap__184
timestamp 1731220617
transform 1 0 1856 0 -1 3280
box 7 3 12 24
use welltap_svt  __well_tap__183
timestamp 1731220617
transform 1 0 3568 0 1 3168
box 7 3 12 24
use welltap_svt  __well_tap__182
timestamp 1731220617
transform 1 0 1856 0 1 3168
box 7 3 12 24
use welltap_svt  __well_tap__181
timestamp 1731220617
transform 1 0 3568 0 -1 3132
box 7 3 12 24
use welltap_svt  __well_tap__180
timestamp 1731220617
transform 1 0 1856 0 -1 3132
box 7 3 12 24
use welltap_svt  __well_tap__179
timestamp 1731220617
transform 1 0 3568 0 1 3024
box 7 3 12 24
use welltap_svt  __well_tap__178
timestamp 1731220617
transform 1 0 1856 0 1 3024
box 7 3 12 24
use welltap_svt  __well_tap__177
timestamp 1731220617
transform 1 0 3568 0 -1 2980
box 7 3 12 24
use welltap_svt  __well_tap__176
timestamp 1731220617
transform 1 0 1856 0 -1 2980
box 7 3 12 24
use welltap_svt  __well_tap__175
timestamp 1731220617
transform 1 0 3568 0 1 2868
box 7 3 12 24
use welltap_svt  __well_tap__174
timestamp 1731220617
transform 1 0 1856 0 1 2868
box 7 3 12 24
use welltap_svt  __well_tap__173
timestamp 1731220617
transform 1 0 3568 0 -1 2836
box 7 3 12 24
use welltap_svt  __well_tap__172
timestamp 1731220617
transform 1 0 1856 0 -1 2836
box 7 3 12 24
use welltap_svt  __well_tap__171
timestamp 1731220617
transform 1 0 3568 0 1 2732
box 7 3 12 24
use welltap_svt  __well_tap__170
timestamp 1731220617
transform 1 0 1856 0 1 2732
box 7 3 12 24
use welltap_svt  __well_tap__169
timestamp 1731220617
transform 1 0 3568 0 -1 2700
box 7 3 12 24
use welltap_svt  __well_tap__168
timestamp 1731220617
transform 1 0 1856 0 -1 2700
box 7 3 12 24
use welltap_svt  __well_tap__167
timestamp 1731220617
transform 1 0 3568 0 1 2576
box 7 3 12 24
use welltap_svt  __well_tap__166
timestamp 1731220617
transform 1 0 1856 0 1 2576
box 7 3 12 24
use welltap_svt  __well_tap__165
timestamp 1731220617
transform 1 0 3568 0 -1 2544
box 7 3 12 24
use welltap_svt  __well_tap__164
timestamp 1731220617
transform 1 0 1856 0 -1 2544
box 7 3 12 24
use welltap_svt  __well_tap__163
timestamp 1731220617
transform 1 0 3568 0 1 2436
box 7 3 12 24
use welltap_svt  __well_tap__162
timestamp 1731220617
transform 1 0 1856 0 1 2436
box 7 3 12 24
use welltap_svt  __well_tap__161
timestamp 1731220617
transform 1 0 3568 0 -1 2400
box 7 3 12 24
use welltap_svt  __well_tap__160
timestamp 1731220617
transform 1 0 1856 0 -1 2400
box 7 3 12 24
use welltap_svt  __well_tap__159
timestamp 1731220617
transform 1 0 3568 0 1 2288
box 7 3 12 24
use welltap_svt  __well_tap__158
timestamp 1731220617
transform 1 0 1856 0 1 2288
box 7 3 12 24
use welltap_svt  __well_tap__157
timestamp 1731220617
transform 1 0 3568 0 -1 2252
box 7 3 12 24
use welltap_svt  __well_tap__156
timestamp 1731220617
transform 1 0 1856 0 -1 2252
box 7 3 12 24
use welltap_svt  __well_tap__155
timestamp 1731220617
transform 1 0 3568 0 1 2144
box 7 3 12 24
use welltap_svt  __well_tap__154
timestamp 1731220617
transform 1 0 1856 0 1 2144
box 7 3 12 24
use welltap_svt  __well_tap__153
timestamp 1731220617
transform 1 0 3568 0 -1 2108
box 7 3 12 24
use welltap_svt  __well_tap__152
timestamp 1731220617
transform 1 0 1856 0 -1 2108
box 7 3 12 24
use welltap_svt  __well_tap__151
timestamp 1731220617
transform 1 0 3568 0 1 1996
box 7 3 12 24
use welltap_svt  __well_tap__150
timestamp 1731220617
transform 1 0 1856 0 1 1996
box 7 3 12 24
use welltap_svt  __well_tap__149
timestamp 1731220617
transform 1 0 3568 0 -1 1960
box 7 3 12 24
use welltap_svt  __well_tap__148
timestamp 1731220617
transform 1 0 1856 0 -1 1960
box 7 3 12 24
use welltap_svt  __well_tap__147
timestamp 1731220617
transform 1 0 3568 0 1 1848
box 7 3 12 24
use welltap_svt  __well_tap__146
timestamp 1731220617
transform 1 0 1856 0 1 1848
box 7 3 12 24
use welltap_svt  __well_tap__145
timestamp 1731220617
transform 1 0 3568 0 -1 1812
box 7 3 12 24
use welltap_svt  __well_tap__144
timestamp 1731220617
transform 1 0 1856 0 -1 1812
box 7 3 12 24
use welltap_svt  __well_tap__143
timestamp 1731220617
transform 1 0 3568 0 1 1700
box 7 3 12 24
use welltap_svt  __well_tap__142
timestamp 1731220617
transform 1 0 1856 0 1 1700
box 7 3 12 24
use welltap_svt  __well_tap__141
timestamp 1731220617
transform 1 0 3568 0 -1 1664
box 7 3 12 24
use welltap_svt  __well_tap__140
timestamp 1731220617
transform 1 0 1856 0 -1 1664
box 7 3 12 24
use welltap_svt  __well_tap__139
timestamp 1731220617
transform 1 0 3568 0 1 1560
box 7 3 12 24
use welltap_svt  __well_tap__138
timestamp 1731220617
transform 1 0 1856 0 1 1560
box 7 3 12 24
use welltap_svt  __well_tap__137
timestamp 1731220617
transform 1 0 3568 0 -1 1520
box 7 3 12 24
use welltap_svt  __well_tap__136
timestamp 1731220617
transform 1 0 1856 0 -1 1520
box 7 3 12 24
use welltap_svt  __well_tap__135
timestamp 1731220617
transform 1 0 3568 0 1 1412
box 7 3 12 24
use welltap_svt  __well_tap__134
timestamp 1731220617
transform 1 0 1856 0 1 1412
box 7 3 12 24
use welltap_svt  __well_tap__133
timestamp 1731220617
transform 1 0 3568 0 -1 1368
box 7 3 12 24
use welltap_svt  __well_tap__132
timestamp 1731220617
transform 1 0 1856 0 -1 1368
box 7 3 12 24
use welltap_svt  __well_tap__131
timestamp 1731220617
transform 1 0 3568 0 1 1264
box 7 3 12 24
use welltap_svt  __well_tap__130
timestamp 1731220617
transform 1 0 1856 0 1 1264
box 7 3 12 24
use welltap_svt  __well_tap__129
timestamp 1731220617
transform 1 0 3568 0 -1 1224
box 7 3 12 24
use welltap_svt  __well_tap__128
timestamp 1731220617
transform 1 0 1856 0 -1 1224
box 7 3 12 24
use welltap_svt  __well_tap__127
timestamp 1731220617
transform 1 0 3568 0 1 1120
box 7 3 12 24
use welltap_svt  __well_tap__126
timestamp 1731220617
transform 1 0 1856 0 1 1120
box 7 3 12 24
use welltap_svt  __well_tap__125
timestamp 1731220617
transform 1 0 3568 0 -1 1080
box 7 3 12 24
use welltap_svt  __well_tap__124
timestamp 1731220617
transform 1 0 1856 0 -1 1080
box 7 3 12 24
use welltap_svt  __well_tap__123
timestamp 1731220617
transform 1 0 3568 0 1 972
box 7 3 12 24
use welltap_svt  __well_tap__122
timestamp 1731220617
transform 1 0 1856 0 1 972
box 7 3 12 24
use welltap_svt  __well_tap__121
timestamp 1731220617
transform 1 0 3568 0 -1 936
box 7 3 12 24
use welltap_svt  __well_tap__120
timestamp 1731220617
transform 1 0 1856 0 -1 936
box 7 3 12 24
use welltap_svt  __well_tap__119
timestamp 1731220617
transform 1 0 3568 0 1 828
box 7 3 12 24
use welltap_svt  __well_tap__118
timestamp 1731220617
transform 1 0 1856 0 1 828
box 7 3 12 24
use welltap_svt  __well_tap__117
timestamp 1731220617
transform 1 0 3568 0 -1 796
box 7 3 12 24
use welltap_svt  __well_tap__116
timestamp 1731220617
transform 1 0 1856 0 -1 796
box 7 3 12 24
use welltap_svt  __well_tap__115
timestamp 1731220617
transform 1 0 3568 0 1 688
box 7 3 12 24
use welltap_svt  __well_tap__114
timestamp 1731220617
transform 1 0 1856 0 1 688
box 7 3 12 24
use welltap_svt  __well_tap__113
timestamp 1731220617
transform 1 0 3568 0 -1 652
box 7 3 12 24
use welltap_svt  __well_tap__112
timestamp 1731220617
transform 1 0 1856 0 -1 652
box 7 3 12 24
use welltap_svt  __well_tap__111
timestamp 1731220617
transform 1 0 3568 0 1 548
box 7 3 12 24
use welltap_svt  __well_tap__110
timestamp 1731220617
transform 1 0 1856 0 1 548
box 7 3 12 24
use welltap_svt  __well_tap__109
timestamp 1731220617
transform 1 0 3568 0 -1 508
box 7 3 12 24
use welltap_svt  __well_tap__108
timestamp 1731220617
transform 1 0 1856 0 -1 508
box 7 3 12 24
use welltap_svt  __well_tap__107
timestamp 1731220617
transform 1 0 3568 0 1 404
box 7 3 12 24
use welltap_svt  __well_tap__106
timestamp 1731220617
transform 1 0 1856 0 1 404
box 7 3 12 24
use welltap_svt  __well_tap__105
timestamp 1731220617
transform 1 0 3568 0 -1 372
box 7 3 12 24
use welltap_svt  __well_tap__104
timestamp 1731220617
transform 1 0 1856 0 -1 372
box 7 3 12 24
use welltap_svt  __well_tap__103
timestamp 1731220617
transform 1 0 3568 0 1 268
box 7 3 12 24
use welltap_svt  __well_tap__102
timestamp 1731220617
transform 1 0 1856 0 1 268
box 7 3 12 24
use welltap_svt  __well_tap__101
timestamp 1731220617
transform 1 0 3568 0 -1 236
box 7 3 12 24
use welltap_svt  __well_tap__100
timestamp 1731220617
transform 1 0 1856 0 -1 236
box 7 3 12 24
use welltap_svt  __well_tap__99
timestamp 1731220617
transform 1 0 3568 0 1 100
box 7 3 12 24
use welltap_svt  __well_tap__98
timestamp 1731220617
transform 1 0 1856 0 1 100
box 7 3 12 24
use welltap_svt  __well_tap__97
timestamp 1731220617
transform 1 0 1816 0 1 3596
box 7 3 12 24
use welltap_svt  __well_tap__96
timestamp 1731220617
transform 1 0 104 0 1 3596
box 7 3 12 24
use welltap_svt  __well_tap__95
timestamp 1731220617
transform 1 0 1816 0 -1 3556
box 7 3 12 24
use welltap_svt  __well_tap__94
timestamp 1731220617
transform 1 0 104 0 -1 3556
box 7 3 12 24
use welltap_svt  __well_tap__93
timestamp 1731220617
transform 1 0 1816 0 1 3452
box 7 3 12 24
use welltap_svt  __well_tap__92
timestamp 1731220617
transform 1 0 104 0 1 3452
box 7 3 12 24
use welltap_svt  __well_tap__91
timestamp 1731220617
transform 1 0 1816 0 -1 3420
box 7 3 12 24
use welltap_svt  __well_tap__90
timestamp 1731220617
transform 1 0 104 0 -1 3420
box 7 3 12 24
use welltap_svt  __well_tap__89
timestamp 1731220617
transform 1 0 1816 0 1 3308
box 7 3 12 24
use welltap_svt  __well_tap__88
timestamp 1731220617
transform 1 0 104 0 1 3308
box 7 3 12 24
use welltap_svt  __well_tap__87
timestamp 1731220617
transform 1 0 1816 0 -1 3272
box 7 3 12 24
use welltap_svt  __well_tap__86
timestamp 1731220617
transform 1 0 104 0 -1 3272
box 7 3 12 24
use welltap_svt  __well_tap__85
timestamp 1731220617
transform 1 0 1816 0 1 3156
box 7 3 12 24
use welltap_svt  __well_tap__84
timestamp 1731220617
transform 1 0 104 0 1 3156
box 7 3 12 24
use welltap_svt  __well_tap__83
timestamp 1731220617
transform 1 0 1816 0 -1 3112
box 7 3 12 24
use welltap_svt  __well_tap__82
timestamp 1731220617
transform 1 0 104 0 -1 3112
box 7 3 12 24
use welltap_svt  __well_tap__81
timestamp 1731220617
transform 1 0 1816 0 1 3008
box 7 3 12 24
use welltap_svt  __well_tap__80
timestamp 1731220617
transform 1 0 104 0 1 3008
box 7 3 12 24
use welltap_svt  __well_tap__79
timestamp 1731220617
transform 1 0 1816 0 -1 2964
box 7 3 12 24
use welltap_svt  __well_tap__78
timestamp 1731220617
transform 1 0 104 0 -1 2964
box 7 3 12 24
use welltap_svt  __well_tap__77
timestamp 1731220617
transform 1 0 1816 0 1 2860
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220617
transform 1 0 104 0 1 2860
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220617
transform 1 0 1816 0 -1 2824
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220617
transform 1 0 104 0 -1 2824
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220617
transform 1 0 1816 0 1 2712
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220617
transform 1 0 104 0 1 2712
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220617
transform 1 0 1816 0 -1 2676
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220617
transform 1 0 104 0 -1 2676
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220617
transform 1 0 1816 0 1 2568
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220617
transform 1 0 104 0 1 2568
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220617
transform 1 0 1816 0 -1 2528
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220617
transform 1 0 104 0 -1 2528
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220617
transform 1 0 1816 0 1 2420
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220617
transform 1 0 104 0 1 2420
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220617
transform 1 0 1816 0 -1 2384
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220617
transform 1 0 104 0 -1 2384
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220617
transform 1 0 1816 0 1 2276
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220617
transform 1 0 104 0 1 2276
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220617
transform 1 0 1816 0 -1 2236
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220617
transform 1 0 104 0 -1 2236
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220617
transform 1 0 1816 0 1 2128
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220617
transform 1 0 104 0 1 2128
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220617
transform 1 0 1816 0 -1 2088
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220617
transform 1 0 104 0 -1 2088
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220617
transform 1 0 1816 0 1 1976
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220617
transform 1 0 104 0 1 1976
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220617
transform 1 0 1816 0 -1 1936
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220617
transform 1 0 104 0 -1 1936
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220617
transform 1 0 1816 0 1 1824
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220617
transform 1 0 104 0 1 1824
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220617
transform 1 0 1816 0 -1 1784
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220617
transform 1 0 104 0 -1 1784
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220617
transform 1 0 1816 0 1 1680
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220617
transform 1 0 104 0 1 1680
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220617
transform 1 0 1816 0 -1 1648
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220617
transform 1 0 104 0 -1 1648
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220617
transform 1 0 1816 0 1 1540
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220617
transform 1 0 104 0 1 1540
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220617
transform 1 0 1816 0 -1 1504
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220617
transform 1 0 104 0 -1 1504
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220617
transform 1 0 1816 0 1 1396
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220617
transform 1 0 104 0 1 1396
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220617
transform 1 0 1816 0 -1 1364
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220617
transform 1 0 104 0 -1 1364
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220617
transform 1 0 1816 0 1 1260
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220617
transform 1 0 104 0 1 1260
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220617
transform 1 0 1816 0 -1 1228
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220617
transform 1 0 104 0 -1 1228
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220617
transform 1 0 1816 0 1 1116
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220617
transform 1 0 104 0 1 1116
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220617
transform 1 0 1816 0 -1 1080
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220617
transform 1 0 104 0 -1 1080
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220617
transform 1 0 1816 0 1 972
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220617
transform 1 0 104 0 1 972
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220617
transform 1 0 1816 0 -1 936
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220617
transform 1 0 104 0 -1 936
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220617
transform 1 0 1816 0 1 828
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220617
transform 1 0 104 0 1 828
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220617
transform 1 0 1816 0 -1 796
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220617
transform 1 0 104 0 -1 796
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220617
transform 1 0 1816 0 1 688
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220617
transform 1 0 104 0 1 688
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220617
transform 1 0 1816 0 -1 652
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220617
transform 1 0 104 0 -1 652
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220617
transform 1 0 1816 0 1 548
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220617
transform 1 0 104 0 1 548
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220617
transform 1 0 1816 0 -1 516
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220617
transform 1 0 104 0 -1 516
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220617
transform 1 0 1816 0 1 404
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220617
transform 1 0 104 0 1 404
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220617
transform 1 0 1816 0 -1 372
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220617
transform 1 0 104 0 -1 372
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220617
transform 1 0 1816 0 1 264
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220617
transform 1 0 104 0 1 264
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220617
transform 1 0 1816 0 -1 228
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220617
transform 1 0 104 0 -1 228
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220617
transform 1 0 1816 0 1 104
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220617
transform 1 0 104 0 1 104
box 7 3 12 24
use _0_0std_0_0cells_0_0MUX2X1  tst_5999_6
timestamp 1731220617
transform 1 0 3472 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5998_6
timestamp 1731220617
transform 1 0 3472 0 -1 668
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5997_6
timestamp 1731220617
transform 1 0 3472 0 -1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5996_6
timestamp 1731220617
transform 1 0 3448 0 1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5995_6
timestamp 1731220617
transform 1 0 3424 0 1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5994_6
timestamp 1731220617
transform 1 0 3472 0 -1 524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5993_6
timestamp 1731220617
transform 1 0 3472 0 1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5992_6
timestamp 1731220617
transform 1 0 3472 0 -1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5991_6
timestamp 1731220617
transform 1 0 3472 0 -1 252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5990_6
timestamp 1731220617
transform 1 0 3472 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5989_6
timestamp 1731220617
transform 1 0 3384 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5988_6
timestamp 1731220617
transform 1 0 3296 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5987_6
timestamp 1731220617
transform 1 0 3200 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5986_6
timestamp 1731220617
transform 1 0 3104 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5985_6
timestamp 1731220617
transform 1 0 3008 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5984_6
timestamp 1731220617
transform 1 0 2912 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5983_6
timestamp 1731220617
transform 1 0 2808 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5982_6
timestamp 1731220617
transform 1 0 2704 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5981_6
timestamp 1731220617
transform 1 0 2592 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5980_6
timestamp 1731220617
transform 1 0 3304 0 -1 252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5979_6
timestamp 1731220617
transform 1 0 3120 0 -1 252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5978_6
timestamp 1731220617
transform 1 0 2944 0 -1 252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5977_6
timestamp 1731220617
transform 1 0 2760 0 -1 252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5976_6
timestamp 1731220617
transform 1 0 2576 0 -1 252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5975_6
timestamp 1731220617
transform 1 0 2952 0 1 252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5974_6
timestamp 1731220617
transform 1 0 2840 0 1 252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5973_6
timestamp 1731220617
transform 1 0 2728 0 1 252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5972_6
timestamp 1731220617
transform 1 0 2624 0 1 252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5971_6
timestamp 1731220617
transform 1 0 2520 0 1 252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5970_6
timestamp 1731220617
transform 1 0 2608 0 -1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5969_6
timestamp 1731220617
transform 1 0 2744 0 -1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5968_6
timestamp 1731220617
transform 1 0 3296 0 -1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5967_6
timestamp 1731220617
transform 1 0 3096 0 -1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5966_6
timestamp 1731220617
transform 1 0 2912 0 -1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5965_6
timestamp 1731220617
transform 1 0 2848 0 1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5964_6
timestamp 1731220617
transform 1 0 2720 0 1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5963_6
timestamp 1731220617
transform 1 0 2992 0 1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5962_6
timestamp 1731220617
transform 1 0 3320 0 1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5961_6
timestamp 1731220617
transform 1 0 3152 0 1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5960_6
timestamp 1731220617
transform 1 0 3008 0 -1 524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5959_6
timestamp 1731220617
transform 1 0 2840 0 -1 524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5958_6
timestamp 1731220617
transform 1 0 2664 0 -1 524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5957_6
timestamp 1731220617
transform 1 0 3168 0 -1 524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5956_6
timestamp 1731220617
transform 1 0 3328 0 -1 524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5955_6
timestamp 1731220617
transform 1 0 3184 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5954_6
timestamp 1731220617
transform 1 0 3024 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5953_6
timestamp 1731220617
transform 1 0 3336 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5952_6
timestamp 1731220617
transform 1 0 3344 0 -1 668
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5951_6
timestamp 1731220617
transform 1 0 3200 0 -1 668
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5950_6
timestamp 1731220617
transform 1 0 3272 0 1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5949_6
timestamp 1731220617
transform 1 0 3056 0 -1 668
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5948_6
timestamp 1731220617
transform 1 0 2904 0 -1 668
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5947_6
timestamp 1731220617
transform 1 0 2864 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5946_6
timestamp 1731220617
transform 1 0 2688 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5945_6
timestamp 1731220617
transform 1 0 2736 0 -1 668
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5944_6
timestamp 1731220617
transform 1 0 3120 0 1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5943_6
timestamp 1731220617
transform 1 0 2968 0 1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5942_6
timestamp 1731220617
transform 1 0 2824 0 1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5941_6
timestamp 1731220617
transform 1 0 2680 0 1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5940_6
timestamp 1731220617
transform 1 0 3288 0 -1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5939_6
timestamp 1731220617
transform 1 0 3104 0 -1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5938_6
timestamp 1731220617
transform 1 0 2928 0 -1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5937_6
timestamp 1731220617
transform 1 0 2776 0 -1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5936_6
timestamp 1731220617
transform 1 0 2648 0 -1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5935_6
timestamp 1731220617
transform 1 0 3240 0 1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5934_6
timestamp 1731220617
transform 1 0 3040 0 1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5933_6
timestamp 1731220617
transform 1 0 2856 0 1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5932_6
timestamp 1731220617
transform 1 0 2688 0 1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5931_6
timestamp 1731220617
transform 1 0 2552 0 1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5930_6
timestamp 1731220617
transform 1 0 2744 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5929_6
timestamp 1731220617
transform 1 0 2896 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5928_6
timestamp 1731220617
transform 1 0 3072 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5927_6
timestamp 1731220617
transform 1 0 3256 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5926_6
timestamp 1731220617
transform 1 0 3296 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5925_6
timestamp 1731220617
transform 1 0 3120 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5924_6
timestamp 1731220617
transform 1 0 2944 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5923_6
timestamp 1731220617
transform 1 0 2776 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5922_6
timestamp 1731220617
transform 1 0 2888 0 -1 1096
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5921_6
timestamp 1731220617
transform 1 0 3040 0 -1 1096
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5920_6
timestamp 1731220617
transform 1 0 3192 0 -1 1096
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5919_6
timestamp 1731220617
transform 1 0 3344 0 -1 1096
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5918_6
timestamp 1731220617
transform 1 0 3312 0 1 1104
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5917_6
timestamp 1731220617
transform 1 0 3128 0 1 1104
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5916_6
timestamp 1731220617
transform 1 0 2984 0 -1 1240
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5915_6
timestamp 1731220617
transform 1 0 3152 0 -1 1240
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5914_6
timestamp 1731220617
transform 1 0 3320 0 -1 1240
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5913_6
timestamp 1731220617
transform 1 0 3304 0 1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5912_6
timestamp 1731220617
transform 1 0 3120 0 1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5911_6
timestamp 1731220617
transform 1 0 2944 0 1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5910_6
timestamp 1731220617
transform 1 0 3056 0 -1 1384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5909_6
timestamp 1731220617
transform 1 0 2840 0 -1 1384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5908_6
timestamp 1731220617
transform 1 0 2920 0 1 1396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5907_6
timestamp 1731220617
transform 1 0 3264 0 1 1396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5906_6
timestamp 1731220617
transform 1 0 3088 0 1 1396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5905_6
timestamp 1731220617
transform 1 0 3048 0 -1 1536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5904_6
timestamp 1731220617
transform 1 0 2872 0 -1 1536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5903_6
timestamp 1731220617
transform 1 0 2752 0 1 1396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5902_6
timestamp 1731220617
transform 1 0 2600 0 1 1396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5901_6
timestamp 1731220617
transform 1 0 2384 0 -1 1384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5900_6
timestamp 1731220617
transform 1 0 2616 0 -1 1384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5899_6
timestamp 1731220617
transform 1 0 2608 0 1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5898_6
timestamp 1731220617
transform 1 0 2776 0 1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5897_6
timestamp 1731220617
transform 1 0 2816 0 -1 1240
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5896_6
timestamp 1731220617
transform 1 0 2648 0 -1 1240
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5895_6
timestamp 1731220617
transform 1 0 2608 0 1 1104
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5894_6
timestamp 1731220617
transform 1 0 2952 0 1 1104
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5893_6
timestamp 1731220617
transform 1 0 2776 0 1 1104
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5892_6
timestamp 1731220617
transform 1 0 2728 0 -1 1096
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5891_6
timestamp 1731220617
transform 1 0 2624 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5890_6
timestamp 1731220617
transform 1 0 2608 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5889_6
timestamp 1731220617
transform 1 0 2440 0 1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5888_6
timestamp 1731220617
transform 1 0 2352 0 1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5887_6
timestamp 1731220617
transform 1 0 2456 0 -1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5886_6
timestamp 1731220617
transform 1 0 2544 0 -1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5885_6
timestamp 1731220617
transform 1 0 2536 0 1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5884_6
timestamp 1731220617
transform 1 0 2392 0 1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5883_6
timestamp 1731220617
transform 1 0 2240 0 1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5882_6
timestamp 1731220617
transform 1 0 2192 0 -1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5881_6
timestamp 1731220617
transform 1 0 2368 0 -1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5880_6
timestamp 1731220617
transform 1 0 2280 0 -1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5879_6
timestamp 1731220617
transform 1 0 2264 0 1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5878_6
timestamp 1731220617
transform 1 0 2176 0 1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5877_6
timestamp 1731220617
transform 1 0 2088 0 1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5876_6
timestamp 1731220617
transform 1 0 2136 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5875_6
timestamp 1731220617
transform 1 0 2224 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5874_6
timestamp 1731220617
transform 1 0 2312 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5873_6
timestamp 1731220617
transform 1 0 2400 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5872_6
timestamp 1731220617
transform 1 0 2496 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5871_6
timestamp 1731220617
transform 1 0 2480 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5870_6
timestamp 1731220617
transform 1 0 2560 0 -1 1096
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5869_6
timestamp 1731220617
transform 1 0 2440 0 1 1104
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5868_6
timestamp 1731220617
transform 1 0 2480 0 -1 1240
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5867_6
timestamp 1731220617
transform 1 0 2440 0 1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5866_6
timestamp 1731220617
transform 1 0 2136 0 -1 1384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5865_6
timestamp 1731220617
transform 1 0 2448 0 1 1396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5864_6
timestamp 1731220617
transform 1 0 2536 0 -1 1536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5863_6
timestamp 1731220617
transform 1 0 2704 0 -1 1536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5862_6
timestamp 1731220617
transform 1 0 2592 0 1 1544
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5861_6
timestamp 1731220617
transform 1 0 2752 0 1 1544
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5860_6
timestamp 1731220617
transform 1 0 2928 0 1 1544
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5859_6
timestamp 1731220617
transform 1 0 2968 0 -1 1680
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5858_6
timestamp 1731220617
transform 1 0 2800 0 -1 1680
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5857_6
timestamp 1731220617
transform 1 0 2880 0 1 1684
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5856_6
timestamp 1731220617
transform 1 0 3000 0 1 1684
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5855_6
timestamp 1731220617
transform 1 0 3136 0 -1 1680
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5854_6
timestamp 1731220617
transform 1 0 3112 0 1 1544
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5853_6
timestamp 1731220617
transform 1 0 3304 0 1 1544
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5852_6
timestamp 1731220617
transform 1 0 3232 0 -1 1536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5851_6
timestamp 1731220617
transform 1 0 3264 0 -1 1384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5850_6
timestamp 1731220617
transform 1 0 3472 0 -1 1096
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5849_6
timestamp 1731220617
transform 1 0 3448 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5848_6
timestamp 1731220617
transform 1 0 3472 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5847_6
timestamp 1731220617
transform 1 0 3472 0 1 1104
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5846_6
timestamp 1731220617
transform 1 0 3472 0 -1 1240
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5845_6
timestamp 1731220617
transform 1 0 3472 0 1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5844_6
timestamp 1731220617
transform 1 0 3472 0 -1 1384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5843_6
timestamp 1731220617
transform 1 0 3448 0 1 1396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5842_6
timestamp 1731220617
transform 1 0 3424 0 -1 1536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5841_6
timestamp 1731220617
transform 1 0 3312 0 -1 1680
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5840_6
timestamp 1731220617
transform 1 0 3240 0 1 1684
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5839_6
timestamp 1731220617
transform 1 0 3120 0 1 1684
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5838_6
timestamp 1731220617
transform 1 0 3368 0 1 1684
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5837_6
timestamp 1731220617
transform 1 0 3312 0 -1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5836_6
timestamp 1731220617
transform 1 0 3176 0 -1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5835_6
timestamp 1731220617
transform 1 0 3040 0 -1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5834_6
timestamp 1731220617
transform 1 0 2912 0 -1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5833_6
timestamp 1731220617
transform 1 0 2792 0 -1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5832_6
timestamp 1731220617
transform 1 0 3296 0 1 1832
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5831_6
timestamp 1731220617
transform 1 0 3104 0 1 1832
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5830_6
timestamp 1731220617
transform 1 0 2920 0 1 1832
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5829_6
timestamp 1731220617
transform 1 0 2760 0 1 1832
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5828_6
timestamp 1731220617
transform 1 0 2624 0 1 1832
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5827_6
timestamp 1731220617
transform 1 0 2496 0 -1 1976
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5826_6
timestamp 1731220617
transform 1 0 2648 0 -1 1976
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5825_6
timestamp 1731220617
transform 1 0 2832 0 -1 1976
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5824_6
timestamp 1731220617
transform 1 0 3040 0 -1 1976
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5823_6
timestamp 1731220617
transform 1 0 3264 0 -1 1976
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5822_6
timestamp 1731220617
transform 1 0 3296 0 1 1980
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5821_6
timestamp 1731220617
transform 1 0 3104 0 1 1980
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5820_6
timestamp 1731220617
transform 1 0 2920 0 1 1980
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5819_6
timestamp 1731220617
transform 1 0 2744 0 1 1980
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5818_6
timestamp 1731220617
transform 1 0 2576 0 1 1980
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5817_6
timestamp 1731220617
transform 1 0 2712 0 -1 2124
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5816_6
timestamp 1731220617
transform 1 0 2872 0 -1 2124
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5815_6
timestamp 1731220617
transform 1 0 3024 0 -1 2124
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5814_6
timestamp 1731220617
transform 1 0 3168 0 -1 2124
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5813_6
timestamp 1731220617
transform 1 0 3312 0 -1 2124
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5812_6
timestamp 1731220617
transform 1 0 3344 0 1 2128
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5811_6
timestamp 1731220617
transform 1 0 3200 0 1 2128
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5810_6
timestamp 1731220617
transform 1 0 3056 0 1 2128
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5809_6
timestamp 1731220617
transform 1 0 2904 0 1 2128
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5808_6
timestamp 1731220617
transform 1 0 2744 0 1 2128
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5807_6
timestamp 1731220617
transform 1 0 3232 0 -1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5806_6
timestamp 1731220617
transform 1 0 3072 0 -1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5805_6
timestamp 1731220617
transform 1 0 2904 0 -1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5804_6
timestamp 1731220617
transform 1 0 2736 0 -1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5803_6
timestamp 1731220617
transform 1 0 3272 0 1 2272
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5802_6
timestamp 1731220617
transform 1 0 3096 0 1 2272
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5801_6
timestamp 1731220617
transform 1 0 2928 0 1 2272
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5800_6
timestamp 1731220617
transform 1 0 2760 0 1 2272
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5799_6
timestamp 1731220617
transform 1 0 2600 0 1 2272
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5798_6
timestamp 1731220617
transform 1 0 3104 0 -1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5797_6
timestamp 1731220617
transform 1 0 2920 0 -1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5796_6
timestamp 1731220617
transform 1 0 2744 0 -1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5795_6
timestamp 1731220617
transform 1 0 2584 0 -1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5794_6
timestamp 1731220617
transform 1 0 3072 0 1 2420
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5793_6
timestamp 1731220617
transform 1 0 2872 0 1 2420
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5792_6
timestamp 1731220617
transform 1 0 2688 0 1 2420
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5791_6
timestamp 1731220617
transform 1 0 2528 0 1 2420
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5790_6
timestamp 1731220617
transform 1 0 2688 0 -1 2560
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5789_6
timestamp 1731220617
transform 1 0 2840 0 -1 2560
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5788_6
timestamp 1731220617
transform 1 0 2992 0 -1 2560
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5787_6
timestamp 1731220617
transform 1 0 2984 0 1 2560
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5786_6
timestamp 1731220617
transform 1 0 2832 0 1 2560
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5785_6
timestamp 1731220617
transform 1 0 3144 0 1 2560
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5784_6
timestamp 1731220617
transform 1 0 3152 0 -1 2560
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5783_6
timestamp 1731220617
transform 1 0 3320 0 -1 2560
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5782_6
timestamp 1731220617
transform 1 0 3280 0 1 2420
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5781_6
timestamp 1731220617
transform 1 0 3296 0 -1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5780_6
timestamp 1731220617
transform 1 0 3400 0 -1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5779_6
timestamp 1731220617
transform 1 0 3464 0 -1 2124
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5778_6
timestamp 1731220617
transform 1 0 3456 0 -1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5777_6
timestamp 1731220617
transform 1 0 3472 0 1 1544
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5776_6
timestamp 1731220617
transform 1 0 3472 0 -1 1680
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5775_6
timestamp 1731220617
transform 1 0 3472 0 1 1684
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5774_6
timestamp 1731220617
transform 1 0 3472 0 1 1832
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5773_6
timestamp 1731220617
transform 1 0 3472 0 -1 1976
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5772_6
timestamp 1731220617
transform 1 0 3472 0 1 1980
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5771_6
timestamp 1731220617
transform 1 0 3472 0 1 2128
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5770_6
timestamp 1731220617
transform 1 0 3456 0 1 2272
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5769_6
timestamp 1731220617
transform 1 0 3472 0 -1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5768_6
timestamp 1731220617
transform 1 0 3472 0 1 2420
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5767_6
timestamp 1731220617
transform 1 0 3472 0 -1 2560
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5766_6
timestamp 1731220617
transform 1 0 3472 0 -1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5765_6
timestamp 1731220617
transform 1 0 3472 0 1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5764_6
timestamp 1731220617
transform 1 0 3472 0 1 2852
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5763_6
timestamp 1731220617
transform 1 0 3472 0 -1 2996
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5762_6
timestamp 1731220617
transform 1 0 3472 0 1 3008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5761_6
timestamp 1731220617
transform 1 0 3360 0 1 3008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5760_6
timestamp 1731220617
transform 1 0 3472 0 -1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5759_6
timestamp 1731220617
transform 1 0 3376 0 -1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5758_6
timestamp 1731220617
transform 1 0 3264 0 -1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5757_6
timestamp 1731220617
transform 1 0 3152 0 -1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5756_6
timestamp 1731220617
transform 1 0 3224 0 1 3008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5755_6
timestamp 1731220617
transform 1 0 3384 0 -1 2996
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5754_6
timestamp 1731220617
transform 1 0 3288 0 -1 2996
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5753_6
timestamp 1731220617
transform 1 0 3192 0 -1 2996
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5752_6
timestamp 1731220617
transform 1 0 3096 0 -1 2996
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5751_6
timestamp 1731220617
transform 1 0 3000 0 -1 2996
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5750_6
timestamp 1731220617
transform 1 0 2792 0 -1 2996
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5749_6
timestamp 1731220617
transform 1 0 2680 0 -1 2996
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5748_6
timestamp 1731220617
transform 1 0 2960 0 1 3008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5747_6
timestamp 1731220617
transform 1 0 3096 0 1 3008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5746_6
timestamp 1731220617
transform 1 0 3032 0 -1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5745_6
timestamp 1731220617
transform 1 0 2912 0 -1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5744_6
timestamp 1731220617
transform 1 0 2784 0 -1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5743_6
timestamp 1731220617
transform 1 0 2952 0 1 3152
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5742_6
timestamp 1731220617
transform 1 0 3104 0 1 3152
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5741_6
timestamp 1731220617
transform 1 0 3264 0 1 3152
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5740_6
timestamp 1731220617
transform 1 0 3176 0 -1 3296
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5739_6
timestamp 1731220617
transform 1 0 3024 0 -1 3296
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5738_6
timestamp 1731220617
transform 1 0 2880 0 -1 3296
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5737_6
timestamp 1731220617
transform 1 0 2816 0 1 3296
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5736_6
timestamp 1731220617
transform 1 0 2952 0 1 3296
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5735_6
timestamp 1731220617
transform 1 0 3088 0 1 3296
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5734_6
timestamp 1731220617
transform 1 0 3048 0 -1 3432
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5733_6
timestamp 1731220617
transform 1 0 2912 0 -1 3432
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5732_6
timestamp 1731220617
transform 1 0 2776 0 -1 3432
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5731_6
timestamp 1731220617
transform 1 0 2648 0 -1 3432
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5730_6
timestamp 1731220617
transform 1 0 2520 0 -1 3432
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5729_6
timestamp 1731220617
transform 1 0 2544 0 1 3296
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5728_6
timestamp 1731220617
transform 1 0 2680 0 1 3296
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5727_6
timestamp 1731220617
transform 1 0 2736 0 -1 3296
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5726_6
timestamp 1731220617
transform 1 0 2592 0 -1 3296
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5725_6
timestamp 1731220617
transform 1 0 2648 0 1 3152
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5724_6
timestamp 1731220617
transform 1 0 2800 0 1 3152
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5723_6
timestamp 1731220617
transform 1 0 2648 0 -1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5722_6
timestamp 1731220617
transform 1 0 2664 0 1 3008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5721_6
timestamp 1731220617
transform 1 0 2816 0 1 3008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5720_6
timestamp 1731220617
transform 1 0 2896 0 -1 2996
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5719_6
timestamp 1731220617
transform 1 0 2880 0 1 2852
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5718_6
timestamp 1731220617
transform 1 0 3184 0 1 2852
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5717_6
timestamp 1731220617
transform 1 0 3088 0 -1 2852
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5716_6
timestamp 1731220617
transform 1 0 3000 0 -1 2852
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5715_6
timestamp 1731220617
transform 1 0 2912 0 -1 2852
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5714_6
timestamp 1731220617
transform 1 0 2824 0 -1 2852
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5713_6
timestamp 1731220617
transform 1 0 3312 0 1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5712_6
timestamp 1731220617
transform 1 0 3128 0 1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5711_6
timestamp 1731220617
transform 1 0 2952 0 1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5710_6
timestamp 1731220617
transform 1 0 2792 0 1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5709_6
timestamp 1731220617
transform 1 0 2656 0 1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5708_6
timestamp 1731220617
transform 1 0 3384 0 -1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5707_6
timestamp 1731220617
transform 1 0 3288 0 -1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5706_6
timestamp 1731220617
transform 1 0 3200 0 -1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5705_6
timestamp 1731220617
transform 1 0 3112 0 -1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5704_6
timestamp 1731220617
transform 1 0 3024 0 -1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5703_6
timestamp 1731220617
transform 1 0 2936 0 -1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5702_6
timestamp 1731220617
transform 1 0 2848 0 -1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5701_6
timestamp 1731220617
transform 1 0 2760 0 -1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5700_6
timestamp 1731220617
transform 1 0 2672 0 -1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5699_6
timestamp 1731220617
transform 1 0 2584 0 -1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5698_6
timestamp 1731220617
transform 1 0 2496 0 -1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5697_6
timestamp 1731220617
transform 1 0 2408 0 -1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5696_6
timestamp 1731220617
transform 1 0 2320 0 -1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5695_6
timestamp 1731220617
transform 1 0 2232 0 -1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5694_6
timestamp 1731220617
transform 1 0 2144 0 -1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5693_6
timestamp 1731220617
transform 1 0 2056 0 -1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5692_6
timestamp 1731220617
transform 1 0 1968 0 -1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5691_6
timestamp 1731220617
transform 1 0 1880 0 -1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5690_6
timestamp 1731220617
transform 1 0 2680 0 1 2560
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5689_6
timestamp 1731220617
transform 1 0 2536 0 1 2560
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5688_6
timestamp 1731220617
transform 1 0 2400 0 1 2560
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5687_6
timestamp 1731220617
transform 1 0 2264 0 1 2560
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5686_6
timestamp 1731220617
transform 1 0 2144 0 1 2560
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5685_6
timestamp 1731220617
transform 1 0 2552 0 -1 2560
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5684_6
timestamp 1731220617
transform 1 0 2424 0 -1 2560
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5683_6
timestamp 1731220617
transform 1 0 2304 0 -1 2560
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5682_6
timestamp 1731220617
transform 1 0 2192 0 -1 2560
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5681_6
timestamp 1731220617
transform 1 0 2096 0 -1 2560
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5680_6
timestamp 1731220617
transform 1 0 2392 0 1 2420
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5679_6
timestamp 1731220617
transform 1 0 2272 0 1 2420
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5678_6
timestamp 1731220617
transform 1 0 2168 0 1 2420
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5677_6
timestamp 1731220617
transform 1 0 2072 0 1 2420
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5676_6
timestamp 1731220617
transform 1 0 2440 0 -1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5675_6
timestamp 1731220617
transform 1 0 2304 0 -1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5674_6
timestamp 1731220617
transform 1 0 2176 0 -1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5673_6
timestamp 1731220617
transform 1 0 2056 0 -1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5672_6
timestamp 1731220617
transform 1 0 1944 0 -1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5671_6
timestamp 1731220617
transform 1 0 2448 0 1 2272
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5670_6
timestamp 1731220617
transform 1 0 2296 0 1 2272
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5669_6
timestamp 1731220617
transform 1 0 2144 0 1 2272
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5668_6
timestamp 1731220617
transform 1 0 1992 0 1 2272
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5667_6
timestamp 1731220617
transform 1 0 1880 0 1 2272
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5666_6
timestamp 1731220617
transform 1 0 2560 0 -1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5665_6
timestamp 1731220617
transform 1 0 2376 0 -1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5664_6
timestamp 1731220617
transform 1 0 2192 0 -1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5663_6
timestamp 1731220617
transform 1 0 2016 0 -1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5662_6
timestamp 1731220617
transform 1 0 1880 0 -1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5661_6
timestamp 1731220617
transform 1 0 2568 0 1 2128
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5660_6
timestamp 1731220617
transform 1 0 2384 0 1 2128
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5659_6
timestamp 1731220617
transform 1 0 2200 0 1 2128
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5658_6
timestamp 1731220617
transform 1 0 2024 0 1 2128
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5657_6
timestamp 1731220617
transform 1 0 1880 0 1 2128
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5656_6
timestamp 1731220617
transform 1 0 1880 0 -1 2124
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5655_6
timestamp 1731220617
transform 1 0 2016 0 -1 2124
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5654_6
timestamp 1731220617
transform 1 0 2544 0 -1 2124
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5653_6
timestamp 1731220617
transform 1 0 2368 0 -1 2124
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5652_6
timestamp 1731220617
transform 1 0 2192 0 -1 2124
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5651_6
timestamp 1731220617
transform 1 0 2136 0 1 1980
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5650_6
timestamp 1731220617
transform 1 0 2000 0 1 1980
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5649_6
timestamp 1731220617
transform 1 0 1880 0 1 1980
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5648_6
timestamp 1731220617
transform 1 0 2280 0 1 1980
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5647_6
timestamp 1731220617
transform 1 0 2424 0 1 1980
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5646_6
timestamp 1731220617
transform 1 0 2376 0 -1 1976
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5645_6
timestamp 1731220617
transform 1 0 2280 0 -1 1976
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5644_6
timestamp 1731220617
transform 1 0 2192 0 -1 1976
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5643_6
timestamp 1731220617
transform 1 0 2104 0 -1 1976
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5642_6
timestamp 1731220617
transform 1 0 2016 0 -1 1976
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5641_6
timestamp 1731220617
transform 1 0 2160 0 1 1832
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5640_6
timestamp 1731220617
transform 1 0 2248 0 1 1832
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5639_6
timestamp 1731220617
transform 1 0 2336 0 1 1832
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5638_6
timestamp 1731220617
transform 1 0 2424 0 1 1832
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5637_6
timestamp 1731220617
transform 1 0 2512 0 1 1832
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5636_6
timestamp 1731220617
transform 1 0 2432 0 -1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5635_6
timestamp 1731220617
transform 1 0 2312 0 -1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5634_6
timestamp 1731220617
transform 1 0 2552 0 -1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5633_6
timestamp 1731220617
transform 1 0 2672 0 -1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5632_6
timestamp 1731220617
transform 1 0 2760 0 1 1684
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5631_6
timestamp 1731220617
transform 1 0 2640 0 1 1684
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5630_6
timestamp 1731220617
transform 1 0 2512 0 1 1684
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5629_6
timestamp 1731220617
transform 1 0 2392 0 1 1684
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5628_6
timestamp 1731220617
transform 1 0 2280 0 1 1684
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5627_6
timestamp 1731220617
transform 1 0 2640 0 -1 1680
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5626_6
timestamp 1731220617
transform 1 0 2496 0 -1 1680
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5625_6
timestamp 1731220617
transform 1 0 2360 0 -1 1680
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5624_6
timestamp 1731220617
transform 1 0 2240 0 -1 1680
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5623_6
timestamp 1731220617
transform 1 0 2136 0 -1 1680
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5622_6
timestamp 1731220617
transform 1 0 2448 0 1 1544
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5621_6
timestamp 1731220617
transform 1 0 2312 0 1 1544
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5620_6
timestamp 1731220617
transform 1 0 2192 0 1 1544
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5619_6
timestamp 1731220617
transform 1 0 2088 0 1 1544
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5618_6
timestamp 1731220617
transform 1 0 1992 0 1 1544
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5617_6
timestamp 1731220617
transform 1 0 2376 0 -1 1536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5616_6
timestamp 1731220617
transform 1 0 2232 0 -1 1536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5615_6
timestamp 1731220617
transform 1 0 2096 0 -1 1536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5614_6
timestamp 1731220617
transform 1 0 1968 0 -1 1536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5613_6
timestamp 1731220617
transform 1 0 1880 0 -1 1536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5612_6
timestamp 1731220617
transform 1 0 2304 0 1 1396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5611_6
timestamp 1731220617
transform 1 0 2160 0 1 1396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5610_6
timestamp 1731220617
transform 1 0 2008 0 1 1396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5609_6
timestamp 1731220617
transform 1 0 1880 0 1 1396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5608_6
timestamp 1731220617
transform 1 0 1720 0 1 1380
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5607_6
timestamp 1731220617
transform 1 0 1584 0 -1 1380
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5606_6
timestamp 1731220617
transform 1 0 1424 0 -1 1380
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5605_6
timestamp 1731220617
transform 1 0 1880 0 -1 1384
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5604_6
timestamp 1731220617
transform 1 0 1912 0 1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5603_6
timestamp 1731220617
transform 1 0 2096 0 1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5602_6
timestamp 1731220617
transform 1 0 2272 0 1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5601_6
timestamp 1731220617
transform 1 0 2136 0 -1 1240
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5600_6
timestamp 1731220617
transform 1 0 2312 0 -1 1240
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5599_6
timestamp 1731220617
transform 1 0 2280 0 1 1104
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5598_6
timestamp 1731220617
transform 1 0 2208 0 -1 1096
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5597_6
timestamp 1731220617
transform 1 0 2384 0 -1 1096
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5596_6
timestamp 1731220617
transform 1 0 2344 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5595_6
timestamp 1731220617
transform 1 0 2208 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5594_6
timestamp 1731220617
transform 1 0 2080 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5593_6
timestamp 1731220617
transform 1 0 1960 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5592_6
timestamp 1731220617
transform 1 0 1888 0 -1 1096
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5591_6
timestamp 1731220617
transform 1 0 2040 0 -1 1096
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5590_6
timestamp 1731220617
transform 1 0 2128 0 1 1104
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5589_6
timestamp 1731220617
transform 1 0 1992 0 1 1104
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5588_6
timestamp 1731220617
transform 1 0 1880 0 1 1104
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5587_6
timestamp 1731220617
transform 1 0 1720 0 -1 1244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5586_6
timestamp 1731220617
transform 1 0 1600 0 -1 1244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5585_6
timestamp 1731220617
transform 1 0 1720 0 1 1244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5584_6
timestamp 1731220617
transform 1 0 1720 0 -1 1380
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5583_6
timestamp 1731220617
transform 1 0 1584 0 1 1380
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5582_6
timestamp 1731220617
transform 1 0 1432 0 1 1380
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5581_6
timestamp 1731220617
transform 1 0 1280 0 1 1380
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5580_6
timestamp 1731220617
transform 1 0 1704 0 -1 1520
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5579_6
timestamp 1731220617
transform 1 0 1552 0 -1 1520
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5578_6
timestamp 1731220617
transform 1 0 1400 0 -1 1520
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5577_6
timestamp 1731220617
transform 1 0 1248 0 -1 1520
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5576_6
timestamp 1731220617
transform 1 0 1088 0 -1 1520
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5575_6
timestamp 1731220617
transform 1 0 1568 0 1 1524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5574_6
timestamp 1731220617
transform 1 0 1424 0 1 1524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5573_6
timestamp 1731220617
transform 1 0 1280 0 1 1524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5572_6
timestamp 1731220617
transform 1 0 1136 0 1 1524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5571_6
timestamp 1731220617
transform 1 0 984 0 1 1524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5570_6
timestamp 1731220617
transform 1 0 1408 0 -1 1664
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5569_6
timestamp 1731220617
transform 1 0 1272 0 -1 1664
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5568_6
timestamp 1731220617
transform 1 0 1136 0 -1 1664
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5567_6
timestamp 1731220617
transform 1 0 1000 0 -1 1664
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5566_6
timestamp 1731220617
transform 1 0 864 0 -1 1664
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5565_6
timestamp 1731220617
transform 1 0 1248 0 1 1664
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5564_6
timestamp 1731220617
transform 1 0 1112 0 1 1664
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5563_6
timestamp 1731220617
transform 1 0 976 0 1 1664
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5562_6
timestamp 1731220617
transform 1 0 848 0 1 1664
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5561_6
timestamp 1731220617
transform 1 0 712 0 1 1664
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5560_6
timestamp 1731220617
transform 1 0 856 0 -1 1800
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5559_6
timestamp 1731220617
transform 1 0 1000 0 -1 1800
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5558_6
timestamp 1731220617
transform 1 0 1136 0 -1 1800
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5557_6
timestamp 1731220617
transform 1 0 1416 0 -1 1800
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5556_6
timestamp 1731220617
transform 1 0 1272 0 -1 1800
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5555_6
timestamp 1731220617
transform 1 0 1216 0 1 1808
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5554_6
timestamp 1731220617
transform 1 0 1048 0 1 1808
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5553_6
timestamp 1731220617
transform 1 0 1376 0 1 1808
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5552_6
timestamp 1731220617
transform 1 0 1536 0 1 1808
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5551_6
timestamp 1731220617
transform 1 0 1696 0 1 1808
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5550_6
timestamp 1731220617
transform 1 0 1720 0 -1 1952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5549_6
timestamp 1731220617
transform 1 0 1576 0 -1 1952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5548_6
timestamp 1731220617
transform 1 0 1416 0 -1 1952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5547_6
timestamp 1731220617
transform 1 0 1256 0 -1 1952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5546_6
timestamp 1731220617
transform 1 0 1088 0 -1 1952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5545_6
timestamp 1731220617
transform 1 0 1480 0 1 1960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5544_6
timestamp 1731220617
transform 1 0 1352 0 1 1960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5543_6
timestamp 1731220617
transform 1 0 1232 0 1 1960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5542_6
timestamp 1731220617
transform 1 0 1112 0 1 1960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5541_6
timestamp 1731220617
transform 1 0 984 0 1 1960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5540_6
timestamp 1731220617
transform 1 0 1232 0 -1 2104
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5539_6
timestamp 1731220617
transform 1 0 1128 0 -1 2104
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5538_6
timestamp 1731220617
transform 1 0 1024 0 -1 2104
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5537_6
timestamp 1731220617
transform 1 0 920 0 -1 2104
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5536_6
timestamp 1731220617
transform 1 0 824 0 -1 2104
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5535_6
timestamp 1731220617
transform 1 0 816 0 1 2112
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5534_6
timestamp 1731220617
transform 1 0 712 0 1 2112
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5533_6
timestamp 1731220617
transform 1 0 928 0 1 2112
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5532_6
timestamp 1731220617
transform 1 0 1152 0 1 2112
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5531_6
timestamp 1731220617
transform 1 0 1040 0 1 2112
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5530_6
timestamp 1731220617
transform 1 0 1008 0 -1 2252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5529_6
timestamp 1731220617
transform 1 0 864 0 -1 2252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5528_6
timestamp 1731220617
transform 1 0 1152 0 -1 2252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5527_6
timestamp 1731220617
transform 1 0 1448 0 -1 2252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5526_6
timestamp 1731220617
transform 1 0 1296 0 -1 2252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5525_6
timestamp 1731220617
transform 1 0 1216 0 1 2260
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5524_6
timestamp 1731220617
transform 1 0 1040 0 1 2260
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5523_6
timestamp 1731220617
transform 1 0 1392 0 1 2260
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5522_6
timestamp 1731220617
transform 1 0 1568 0 1 2260
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5521_6
timestamp 1731220617
transform 1 0 1720 0 1 2260
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5520_6
timestamp 1731220617
transform 1 0 1704 0 -1 2400
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5519_6
timestamp 1731220617
transform 1 0 1536 0 -1 2400
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5518_6
timestamp 1731220617
transform 1 0 1368 0 -1 2400
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5517_6
timestamp 1731220617
transform 1 0 1200 0 -1 2400
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5516_6
timestamp 1731220617
transform 1 0 1024 0 -1 2400
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5515_6
timestamp 1731220617
transform 1 0 1448 0 1 2404
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5514_6
timestamp 1731220617
transform 1 0 1320 0 1 2404
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5513_6
timestamp 1731220617
transform 1 0 1192 0 1 2404
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5512_6
timestamp 1731220617
transform 1 0 1072 0 1 2404
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5511_6
timestamp 1731220617
transform 1 0 952 0 1 2404
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5510_6
timestamp 1731220617
transform 1 0 1280 0 -1 2544
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5509_6
timestamp 1731220617
transform 1 0 1192 0 -1 2544
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5508_6
timestamp 1731220617
transform 1 0 1104 0 -1 2544
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5507_6
timestamp 1731220617
transform 1 0 1016 0 -1 2544
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5506_6
timestamp 1731220617
transform 1 0 928 0 -1 2544
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5505_6
timestamp 1731220617
transform 1 0 1072 0 1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5504_6
timestamp 1731220617
transform 1 0 984 0 1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5503_6
timestamp 1731220617
transform 1 0 896 0 1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5502_6
timestamp 1731220617
transform 1 0 808 0 1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5501_6
timestamp 1731220617
transform 1 0 696 0 -1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5500_6
timestamp 1731220617
transform 1 0 632 0 1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5499_6
timestamp 1731220617
transform 1 0 544 0 1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5498_6
timestamp 1731220617
transform 1 0 456 0 1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5497_6
timestamp 1731220617
transform 1 0 488 0 -1 2544
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5496_6
timestamp 1731220617
transform 1 0 576 0 -1 2544
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5495_6
timestamp 1731220617
transform 1 0 576 0 1 2404
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5494_6
timestamp 1731220617
transform 1 0 704 0 1 2404
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5493_6
timestamp 1731220617
transform 1 0 656 0 -1 2400
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5492_6
timestamp 1731220617
transform 1 0 840 0 -1 2400
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5491_6
timestamp 1731220617
transform 1 0 848 0 1 2260
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5490_6
timestamp 1731220617
transform 1 0 656 0 1 2260
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5489_6
timestamp 1731220617
transform 1 0 464 0 1 2260
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5488_6
timestamp 1731220617
transform 1 0 552 0 -1 2252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5487_6
timestamp 1731220617
transform 1 0 712 0 -1 2252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5486_6
timestamp 1731220617
transform 1 0 608 0 1 2112
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5485_6
timestamp 1731220617
transform 1 0 504 0 1 2112
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5484_6
timestamp 1731220617
transform 1 0 400 0 1 2112
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5483_6
timestamp 1731220617
transform 1 0 520 0 -1 2104
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5482_6
timestamp 1731220617
transform 1 0 624 0 -1 2104
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5481_6
timestamp 1731220617
transform 1 0 728 0 -1 2104
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5480_6
timestamp 1731220617
transform 1 0 848 0 1 1960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5479_6
timestamp 1731220617
transform 1 0 704 0 1 1960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5478_6
timestamp 1731220617
transform 1 0 544 0 1 1960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5477_6
timestamp 1731220617
transform 1 0 712 0 -1 1952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5476_6
timestamp 1731220617
transform 1 0 904 0 -1 1952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5475_6
timestamp 1731220617
transform 1 0 872 0 1 1808
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5474_6
timestamp 1731220617
transform 1 0 688 0 1 1808
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5473_6
timestamp 1731220617
transform 1 0 496 0 1 1808
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5472_6
timestamp 1731220617
transform 1 0 712 0 -1 1800
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5471_6
timestamp 1731220617
transform 1 0 560 0 -1 1800
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5470_6
timestamp 1731220617
transform 1 0 408 0 -1 1800
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5469_6
timestamp 1731220617
transform 1 0 416 0 1 1664
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5468_6
timestamp 1731220617
transform 1 0 568 0 1 1664
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5467_6
timestamp 1731220617
transform 1 0 568 0 -1 1664
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5466_6
timestamp 1731220617
transform 1 0 416 0 -1 1664
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5465_6
timestamp 1731220617
transform 1 0 720 0 -1 1664
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5464_6
timestamp 1731220617
transform 1 0 664 0 1 1524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5463_6
timestamp 1731220617
transform 1 0 496 0 1 1524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5462_6
timestamp 1731220617
transform 1 0 832 0 1 1524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5461_6
timestamp 1731220617
transform 1 0 928 0 -1 1520
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5460_6
timestamp 1731220617
transform 1 0 752 0 -1 1520
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5459_6
timestamp 1731220617
transform 1 0 568 0 -1 1520
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5458_6
timestamp 1731220617
transform 1 0 816 0 1 1380
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5457_6
timestamp 1731220617
transform 1 0 656 0 1 1380
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5456_6
timestamp 1731220617
transform 1 0 616 0 -1 1380
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5455_6
timestamp 1731220617
transform 1 0 720 0 -1 1380
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5454_6
timestamp 1731220617
transform 1 0 840 0 -1 1380
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5453_6
timestamp 1731220617
transform 1 0 976 0 1 1380
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5452_6
timestamp 1731220617
transform 1 0 1128 0 1 1380
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5451_6
timestamp 1731220617
transform 1 0 1272 0 -1 1380
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5450_6
timestamp 1731220617
transform 1 0 1120 0 -1 1380
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5449_6
timestamp 1731220617
transform 1 0 976 0 -1 1380
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5448_6
timestamp 1731220617
transform 1 0 952 0 1 1244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5447_6
timestamp 1731220617
transform 1 0 1120 0 1 1244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5446_6
timestamp 1731220617
transform 1 0 1312 0 1 1244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5445_6
timestamp 1731220617
transform 1 0 1520 0 1 1244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5444_6
timestamp 1731220617
transform 1 0 1464 0 -1 1244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5443_6
timestamp 1731220617
transform 1 0 1328 0 -1 1244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5442_6
timestamp 1731220617
transform 1 0 1200 0 -1 1244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5441_6
timestamp 1731220617
transform 1 0 1088 0 -1 1244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5440_6
timestamp 1731220617
transform 1 0 984 0 -1 1244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5439_6
timestamp 1731220617
transform 1 0 936 0 1 1100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5438_6
timestamp 1731220617
transform 1 0 1048 0 1 1100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5437_6
timestamp 1731220617
transform 1 0 1168 0 1 1100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5436_6
timestamp 1731220617
transform 1 0 1408 0 1 1100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5435_6
timestamp 1731220617
transform 1 0 1288 0 1 1100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5434_6
timestamp 1731220617
transform 1 0 1248 0 -1 1096
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5433_6
timestamp 1731220617
transform 1 0 1096 0 -1 1096
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5432_6
timestamp 1731220617
transform 1 0 936 0 -1 1096
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5431_6
timestamp 1731220617
transform 1 0 1552 0 -1 1096
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5430_6
timestamp 1731220617
transform 1 0 1400 0 -1 1096
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5429_6
timestamp 1731220617
transform 1 0 1360 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5428_6
timestamp 1731220617
transform 1 0 1192 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5427_6
timestamp 1731220617
transform 1 0 1016 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5426_6
timestamp 1731220617
transform 1 0 1528 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5425_6
timestamp 1731220617
transform 1 0 1696 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5424_6
timestamp 1731220617
transform 1 0 1720 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5423_6
timestamp 1731220617
transform 1 0 1568 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5422_6
timestamp 1731220617
transform 1 0 1392 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5421_6
timestamp 1731220617
transform 1 0 1216 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5420_6
timestamp 1731220617
transform 1 0 1040 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5419_6
timestamp 1731220617
transform 1 0 1680 0 1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5418_6
timestamp 1731220617
transform 1 0 1512 0 1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5417_6
timestamp 1731220617
transform 1 0 1344 0 1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5416_6
timestamp 1731220617
transform 1 0 1176 0 1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5415_6
timestamp 1731220617
transform 1 0 1008 0 1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5414_6
timestamp 1731220617
transform 1 0 1472 0 -1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5413_6
timestamp 1731220617
transform 1 0 1320 0 -1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5412_6
timestamp 1731220617
transform 1 0 1176 0 -1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5411_6
timestamp 1731220617
transform 1 0 1032 0 -1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5410_6
timestamp 1731220617
transform 1 0 888 0 -1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5409_6
timestamp 1731220617
transform 1 0 1224 0 1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5408_6
timestamp 1731220617
transform 1 0 1120 0 1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5407_6
timestamp 1731220617
transform 1 0 1016 0 1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5406_6
timestamp 1731220617
transform 1 0 912 0 1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5405_6
timestamp 1731220617
transform 1 0 816 0 1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5404_6
timestamp 1731220617
transform 1 0 912 0 -1 668
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5403_6
timestamp 1731220617
transform 1 0 1000 0 -1 668
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5402_6
timestamp 1731220617
transform 1 0 1088 0 -1 668
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5401_6
timestamp 1731220617
transform 1 0 1176 0 -1 668
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5400_6
timestamp 1731220617
transform 1 0 1264 0 -1 668
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5399_6
timestamp 1731220617
transform 1 0 1456 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5398_6
timestamp 1731220617
transform 1 0 1312 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5397_6
timestamp 1731220617
transform 1 0 1176 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5396_6
timestamp 1731220617
transform 1 0 1048 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5395_6
timestamp 1731220617
transform 1 0 952 0 -1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5394_6
timestamp 1731220617
transform 1 0 1096 0 -1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5393_6
timestamp 1731220617
transform 1 0 1592 0 1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5392_6
timestamp 1731220617
transform 1 0 1432 0 1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5391_6
timestamp 1731220617
transform 1 0 1360 0 -1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5390_6
timestamp 1731220617
transform 1 0 1232 0 -1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5389_6
timestamp 1731220617
transform 1 0 1488 0 -1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5388_6
timestamp 1731220617
transform 1 0 1600 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5387_6
timestamp 1731220617
transform 1 0 1720 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5386_6
timestamp 1731220617
transform 1 0 1616 0 -1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5385_6
timestamp 1731220617
transform 1 0 1720 0 -1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5384_6
timestamp 1731220617
transform 1 0 1880 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5383_6
timestamp 1731220617
transform 1 0 2072 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5382_6
timestamp 1731220617
transform 1 0 2192 0 -1 668
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5381_6
timestamp 1731220617
transform 1 0 2016 0 -1 668
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5380_6
timestamp 1731220617
transform 1 0 1880 0 -1 668
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5379_6
timestamp 1731220617
transform 1 0 1928 0 1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5378_6
timestamp 1731220617
transform 1 0 2088 0 1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5377_6
timestamp 1731220617
transform 1 0 2376 0 -1 668
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5376_6
timestamp 1731220617
transform 1 0 2560 0 -1 668
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5375_6
timestamp 1731220617
transform 1 0 2496 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5374_6
timestamp 1731220617
transform 1 0 2288 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5373_6
timestamp 1731220617
transform 1 0 2280 0 -1 524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5372_6
timestamp 1731220617
transform 1 0 2072 0 -1 524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5371_6
timestamp 1731220617
transform 1 0 2480 0 -1 524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5370_6
timestamp 1731220617
transform 1 0 2512 0 1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5369_6
timestamp 1731220617
transform 1 0 2416 0 1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5368_6
timestamp 1731220617
transform 1 0 2320 0 1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5367_6
timestamp 1731220617
transform 1 0 2232 0 1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5366_6
timestamp 1731220617
transform 1 0 2608 0 1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5365_6
timestamp 1731220617
transform 1 0 2496 0 -1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5364_6
timestamp 1731220617
transform 1 0 2408 0 -1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5363_6
timestamp 1731220617
transform 1 0 2320 0 -1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5362_6
timestamp 1731220617
transform 1 0 2232 0 -1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5361_6
timestamp 1731220617
transform 1 0 2144 0 -1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5360_6
timestamp 1731220617
transform 1 0 2416 0 1 252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5359_6
timestamp 1731220617
transform 1 0 2312 0 1 252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5358_6
timestamp 1731220617
transform 1 0 2208 0 1 252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5357_6
timestamp 1731220617
transform 1 0 2104 0 1 252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5356_6
timestamp 1731220617
transform 1 0 2008 0 1 252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5355_6
timestamp 1731220617
transform 1 0 1952 0 -1 252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5354_6
timestamp 1731220617
transform 1 0 2168 0 -1 252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5353_6
timestamp 1731220617
transform 1 0 2376 0 -1 252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5352_6
timestamp 1731220617
transform 1 0 2480 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5351_6
timestamp 1731220617
transform 1 0 2368 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5350_6
timestamp 1731220617
transform 1 0 2256 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5349_6
timestamp 1731220617
transform 1 0 2144 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5348_6
timestamp 1731220617
transform 1 0 2056 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5347_6
timestamp 1731220617
transform 1 0 1968 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5346_6
timestamp 1731220617
transform 1 0 1880 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5345_6
timestamp 1731220617
transform 1 0 1720 0 1 88
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5344_6
timestamp 1731220617
transform 1 0 1720 0 -1 244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5343_6
timestamp 1731220617
transform 1 0 1616 0 -1 244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5342_6
timestamp 1731220617
transform 1 0 1488 0 -1 244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5341_6
timestamp 1731220617
transform 1 0 1368 0 -1 244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5340_6
timestamp 1731220617
transform 1 0 1496 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5339_6
timestamp 1731220617
transform 1 0 1672 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5338_6
timestamp 1731220617
transform 1 0 1584 0 -1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5337_6
timestamp 1731220617
transform 1 0 1424 0 -1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5336_6
timestamp 1731220617
transform 1 0 1264 0 -1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5335_6
timestamp 1731220617
transform 1 0 1272 0 1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5334_6
timestamp 1731220617
transform 1 0 1112 0 1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5333_6
timestamp 1731220617
transform 1 0 952 0 1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5332_6
timestamp 1731220617
transform 1 0 944 0 -1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5331_6
timestamp 1731220617
transform 1 0 1104 0 -1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5330_6
timestamp 1731220617
transform 1 0 1328 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5329_6
timestamp 1731220617
transform 1 0 1160 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5328_6
timestamp 1731220617
transform 1 0 992 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5327_6
timestamp 1731220617
transform 1 0 984 0 -1 244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5326_6
timestamp 1731220617
transform 1 0 1112 0 -1 244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5325_6
timestamp 1731220617
transform 1 0 1240 0 -1 244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5324_6
timestamp 1731220617
transform 1 0 1616 0 1 88
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5323_6
timestamp 1731220617
transform 1 0 1496 0 1 88
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5322_6
timestamp 1731220617
transform 1 0 1384 0 1 88
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5321_6
timestamp 1731220617
transform 1 0 1280 0 1 88
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5320_6
timestamp 1731220617
transform 1 0 1176 0 1 88
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5319_6
timestamp 1731220617
transform 1 0 1088 0 1 88
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5318_6
timestamp 1731220617
transform 1 0 1000 0 1 88
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5317_6
timestamp 1731220617
transform 1 0 912 0 1 88
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5316_6
timestamp 1731220617
transform 1 0 824 0 1 88
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5315_6
timestamp 1731220617
transform 1 0 736 0 1 88
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5314_6
timestamp 1731220617
transform 1 0 648 0 1 88
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5313_6
timestamp 1731220617
transform 1 0 560 0 1 88
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5312_6
timestamp 1731220617
transform 1 0 472 0 1 88
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5311_6
timestamp 1731220617
transform 1 0 384 0 1 88
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5310_6
timestamp 1731220617
transform 1 0 296 0 1 88
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5309_6
timestamp 1731220617
transform 1 0 208 0 1 88
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5308_6
timestamp 1731220617
transform 1 0 856 0 -1 244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5307_6
timestamp 1731220617
transform 1 0 728 0 -1 244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5306_6
timestamp 1731220617
transform 1 0 608 0 -1 244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5305_6
timestamp 1731220617
transform 1 0 496 0 -1 244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5304_6
timestamp 1731220617
transform 1 0 392 0 -1 244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5303_6
timestamp 1731220617
transform 1 0 824 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5302_6
timestamp 1731220617
transform 1 0 664 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5301_6
timestamp 1731220617
transform 1 0 512 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5300_6
timestamp 1731220617
transform 1 0 376 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5299_6
timestamp 1731220617
transform 1 0 248 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5298_6
timestamp 1731220617
transform 1 0 776 0 -1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5297_6
timestamp 1731220617
transform 1 0 600 0 -1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5296_6
timestamp 1731220617
transform 1 0 424 0 -1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5295_6
timestamp 1731220617
transform 1 0 256 0 -1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5294_6
timestamp 1731220617
transform 1 0 128 0 -1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5293_6
timestamp 1731220617
transform 1 0 776 0 1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5292_6
timestamp 1731220617
transform 1 0 600 0 1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5291_6
timestamp 1731220617
transform 1 0 424 0 1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5290_6
timestamp 1731220617
transform 1 0 256 0 1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5289_6
timestamp 1731220617
transform 1 0 128 0 1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5288_6
timestamp 1731220617
transform 1 0 152 0 -1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5287_6
timestamp 1731220617
transform 1 0 296 0 -1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5286_6
timestamp 1731220617
transform 1 0 456 0 -1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5285_6
timestamp 1731220617
transform 1 0 624 0 -1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5284_6
timestamp 1731220617
transform 1 0 792 0 -1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5283_6
timestamp 1731220617
transform 1 0 688 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5282_6
timestamp 1731220617
transform 1 0 584 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5281_6
timestamp 1731220617
transform 1 0 488 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5280_6
timestamp 1731220617
transform 1 0 800 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5279_6
timestamp 1731220617
transform 1 0 920 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5278_6
timestamp 1731220617
transform 1 0 824 0 -1 668
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5277_6
timestamp 1731220617
transform 1 0 736 0 -1 668
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5276_6
timestamp 1731220617
transform 1 0 648 0 -1 668
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5275_6
timestamp 1731220617
transform 1 0 560 0 -1 668
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5274_6
timestamp 1731220617
transform 1 0 472 0 -1 668
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5273_6
timestamp 1731220617
transform 1 0 720 0 1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5272_6
timestamp 1731220617
transform 1 0 624 0 1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5271_6
timestamp 1731220617
transform 1 0 528 0 1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5270_6
timestamp 1731220617
transform 1 0 432 0 1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5269_6
timestamp 1731220617
transform 1 0 344 0 1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5268_6
timestamp 1731220617
transform 1 0 736 0 -1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5267_6
timestamp 1731220617
transform 1 0 576 0 -1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5266_6
timestamp 1731220617
transform 1 0 416 0 -1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5265_6
timestamp 1731220617
transform 1 0 264 0 -1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5264_6
timestamp 1731220617
transform 1 0 128 0 -1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5263_6
timestamp 1731220617
transform 1 0 824 0 1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5262_6
timestamp 1731220617
transform 1 0 640 0 1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5261_6
timestamp 1731220617
transform 1 0 456 0 1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5260_6
timestamp 1731220617
transform 1 0 272 0 1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5259_6
timestamp 1731220617
transform 1 0 128 0 1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5258_6
timestamp 1731220617
transform 1 0 128 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5257_6
timestamp 1731220617
transform 1 0 280 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5256_6
timestamp 1731220617
transform 1 0 848 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5255_6
timestamp 1731220617
transform 1 0 656 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5254_6
timestamp 1731220617
transform 1 0 464 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5253_6
timestamp 1731220617
transform 1 0 272 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5252_6
timestamp 1731220617
transform 1 0 128 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5251_6
timestamp 1731220617
transform 1 0 832 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5250_6
timestamp 1731220617
transform 1 0 648 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5249_6
timestamp 1731220617
transform 1 0 456 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5248_6
timestamp 1731220617
transform 1 0 440 0 -1 1096
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5247_6
timestamp 1731220617
transform 1 0 280 0 -1 1096
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5246_6
timestamp 1731220617
transform 1 0 136 0 -1 1096
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5245_6
timestamp 1731220617
transform 1 0 776 0 -1 1096
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5244_6
timestamp 1731220617
transform 1 0 608 0 -1 1096
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5243_6
timestamp 1731220617
transform 1 0 576 0 1 1100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5242_6
timestamp 1731220617
transform 1 0 456 0 1 1100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5241_6
timestamp 1731220617
transform 1 0 344 0 1 1100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5240_6
timestamp 1731220617
transform 1 0 816 0 1 1100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5239_6
timestamp 1731220617
transform 1 0 696 0 1 1100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5238_6
timestamp 1731220617
transform 1 0 624 0 -1 1244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5237_6
timestamp 1731220617
transform 1 0 536 0 -1 1244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5236_6
timestamp 1731220617
transform 1 0 712 0 -1 1244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5235_6
timestamp 1731220617
transform 1 0 888 0 -1 1244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5234_6
timestamp 1731220617
transform 1 0 800 0 -1 1244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5233_6
timestamp 1731220617
transform 1 0 816 0 1 1244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5232_6
timestamp 1731220617
transform 1 0 704 0 1 1244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5231_6
timestamp 1731220617
transform 1 0 616 0 1 1244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5230_6
timestamp 1731220617
transform 1 0 528 0 1 1244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5229_6
timestamp 1731220617
transform 1 0 440 0 1 1244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5228_6
timestamp 1731220617
transform 1 0 432 0 -1 1380
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5227_6
timestamp 1731220617
transform 1 0 344 0 -1 1380
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5226_6
timestamp 1731220617
transform 1 0 520 0 -1 1380
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5225_6
timestamp 1731220617
transform 1 0 504 0 1 1380
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5224_6
timestamp 1731220617
transform 1 0 368 0 1 1380
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5223_6
timestamp 1731220617
transform 1 0 240 0 1 1380
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5222_6
timestamp 1731220617
transform 1 0 208 0 -1 1520
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5221_6
timestamp 1731220617
transform 1 0 384 0 -1 1520
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5220_6
timestamp 1731220617
transform 1 0 320 0 1 1524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5219_6
timestamp 1731220617
transform 1 0 152 0 1 1524
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5218_6
timestamp 1731220617
transform 1 0 256 0 -1 1664
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5217_6
timestamp 1731220617
transform 1 0 128 0 -1 1664
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5216_6
timestamp 1731220617
transform 1 0 128 0 1 1664
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5215_6
timestamp 1731220617
transform 1 0 264 0 1 1664
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5214_6
timestamp 1731220617
transform 1 0 256 0 -1 1800
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5213_6
timestamp 1731220617
transform 1 0 128 0 -1 1800
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5212_6
timestamp 1731220617
transform 1 0 128 0 1 1808
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5211_6
timestamp 1731220617
transform 1 0 296 0 1 1808
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5210_6
timestamp 1731220617
transform 1 0 512 0 -1 1952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5209_6
timestamp 1731220617
transform 1 0 304 0 -1 1952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5208_6
timestamp 1731220617
transform 1 0 128 0 -1 1952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5207_6
timestamp 1731220617
transform 1 0 200 0 1 1960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5206_6
timestamp 1731220617
transform 1 0 376 0 1 1960
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5205_6
timestamp 1731220617
transform 1 0 416 0 -1 2104
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5204_6
timestamp 1731220617
transform 1 0 312 0 -1 2104
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5203_6
timestamp 1731220617
transform 1 0 296 0 1 2112
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5202_6
timestamp 1731220617
transform 1 0 200 0 1 2112
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5201_6
timestamp 1731220617
transform 1 0 400 0 -1 2252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5200_6
timestamp 1731220617
transform 1 0 248 0 -1 2252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5199_6
timestamp 1731220617
transform 1 0 128 0 -1 2252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5198_6
timestamp 1731220617
transform 1 0 128 0 1 2260
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5197_6
timestamp 1731220617
transform 1 0 280 0 1 2260
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5196_6
timestamp 1731220617
transform 1 0 128 0 -1 2400
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5195_6
timestamp 1731220617
transform 1 0 280 0 -1 2400
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5194_6
timestamp 1731220617
transform 1 0 464 0 -1 2400
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5193_6
timestamp 1731220617
transform 1 0 456 0 1 2404
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5192_6
timestamp 1731220617
transform 1 0 344 0 1 2404
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5191_6
timestamp 1731220617
transform 1 0 832 0 1 2404
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5190_6
timestamp 1731220617
transform 1 0 840 0 -1 2544
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5189_6
timestamp 1731220617
transform 1 0 752 0 -1 2544
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5188_6
timestamp 1731220617
transform 1 0 664 0 -1 2544
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5187_6
timestamp 1731220617
transform 1 0 720 0 1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5186_6
timestamp 1731220617
transform 1 0 1248 0 1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5185_6
timestamp 1731220617
transform 1 0 1160 0 1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5184_6
timestamp 1731220617
transform 1 0 1040 0 -1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5183_6
timestamp 1731220617
transform 1 0 928 0 -1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5182_6
timestamp 1731220617
transform 1 0 816 0 -1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5181_6
timestamp 1731220617
transform 1 0 1264 0 -1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5180_6
timestamp 1731220617
transform 1 0 1152 0 -1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5179_6
timestamp 1731220617
transform 1 0 1136 0 1 2696
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5178_6
timestamp 1731220617
transform 1 0 1008 0 1 2696
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5177_6
timestamp 1731220617
transform 1 0 872 0 1 2696
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5176_6
timestamp 1731220617
transform 1 0 1408 0 1 2696
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5175_6
timestamp 1731220617
transform 1 0 1272 0 1 2696
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5174_6
timestamp 1731220617
transform 1 0 1120 0 -1 2840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5173_6
timestamp 1731220617
transform 1 0 968 0 -1 2840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5172_6
timestamp 1731220617
transform 1 0 1552 0 -1 2840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5171_6
timestamp 1731220617
transform 1 0 1408 0 -1 2840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5170_6
timestamp 1731220617
transform 1 0 1264 0 -1 2840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5169_6
timestamp 1731220617
transform 1 0 1224 0 1 2844
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5168_6
timestamp 1731220617
transform 1 0 1056 0 1 2844
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5167_6
timestamp 1731220617
transform 1 0 1696 0 1 2844
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5166_6
timestamp 1731220617
transform 1 0 1536 0 1 2844
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5165_6
timestamp 1731220617
transform 1 0 1384 0 1 2844
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5164_6
timestamp 1731220617
transform 1 0 1304 0 -1 2980
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5163_6
timestamp 1731220617
transform 1 0 1184 0 -1 2980
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5162_6
timestamp 1731220617
transform 1 0 1056 0 -1 2980
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5161_6
timestamp 1731220617
transform 1 0 1416 0 -1 2980
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5160_6
timestamp 1731220617
transform 1 0 1520 0 -1 2980
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5159_6
timestamp 1731220617
transform 1 0 1632 0 -1 2980
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5158_6
timestamp 1731220617
transform 1 0 1720 0 -1 2980
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5157_6
timestamp 1731220617
transform 1 0 1880 0 -1 2996
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5156_6
timestamp 1731220617
transform 1 0 1968 0 -1 2996
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5155_6
timestamp 1731220617
transform 1 0 2056 0 -1 2996
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5154_6
timestamp 1731220617
transform 1 0 2144 0 -1 2996
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5153_6
timestamp 1731220617
transform 1 0 2232 0 -1 2996
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5152_6
timestamp 1731220617
transform 1 0 2344 0 -1 2996
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5151_6
timestamp 1731220617
transform 1 0 2456 0 -1 2996
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5150_6
timestamp 1731220617
transform 1 0 2568 0 -1 2996
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5149_6
timestamp 1731220617
transform 1 0 2512 0 1 3008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5148_6
timestamp 1731220617
transform 1 0 2352 0 1 3008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5147_6
timestamp 1731220617
transform 1 0 2200 0 1 3008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5146_6
timestamp 1731220617
transform 1 0 2064 0 1 3008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5145_6
timestamp 1731220617
transform 1 0 1936 0 1 3008
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5144_6
timestamp 1731220617
transform 1 0 2048 0 -1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5143_6
timestamp 1731220617
transform 1 0 2200 0 -1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5142_6
timestamp 1731220617
transform 1 0 2352 0 -1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5141_6
timestamp 1731220617
transform 1 0 2504 0 -1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5140_6
timestamp 1731220617
transform 1 0 2504 0 1 3152
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5139_6
timestamp 1731220617
transform 1 0 2360 0 1 3152
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5138_6
timestamp 1731220617
transform 1 0 2224 0 1 3152
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5137_6
timestamp 1731220617
transform 1 0 2104 0 1 3152
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5136_6
timestamp 1731220617
transform 1 0 1992 0 1 3152
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5135_6
timestamp 1731220617
transform 1 0 2448 0 -1 3296
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5134_6
timestamp 1731220617
transform 1 0 2304 0 -1 3296
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5133_6
timestamp 1731220617
transform 1 0 2168 0 -1 3296
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5132_6
timestamp 1731220617
transform 1 0 2040 0 -1 3296
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5131_6
timestamp 1731220617
transform 1 0 1920 0 -1 3296
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5130_6
timestamp 1731220617
transform 1 0 2408 0 1 3296
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5129_6
timestamp 1731220617
transform 1 0 2264 0 1 3296
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5128_6
timestamp 1731220617
transform 1 0 2120 0 1 3296
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5127_6
timestamp 1731220617
transform 1 0 1984 0 1 3296
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5126_6
timestamp 1731220617
transform 1 0 1880 0 1 3296
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5125_6
timestamp 1731220617
transform 1 0 2384 0 -1 3432
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5124_6
timestamp 1731220617
transform 1 0 2248 0 -1 3432
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5123_6
timestamp 1731220617
transform 1 0 2112 0 -1 3432
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5122_6
timestamp 1731220617
transform 1 0 1984 0 -1 3432
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5121_6
timestamp 1731220617
transform 1 0 1880 0 -1 3432
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5120_6
timestamp 1731220617
transform 1 0 2144 0 1 3432
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5119_6
timestamp 1731220617
transform 1 0 2056 0 1 3432
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5118_6
timestamp 1731220617
transform 1 0 1968 0 1 3432
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5117_6
timestamp 1731220617
transform 1 0 1880 0 1 3432
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5116_6
timestamp 1731220617
transform 1 0 1720 0 1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5115_6
timestamp 1731220617
transform 1 0 1632 0 1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5114_6
timestamp 1731220617
transform 1 0 1520 0 1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5113_6
timestamp 1731220617
transform 1 0 1720 0 -1 3572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5112_6
timestamp 1731220617
transform 1 0 1632 0 -1 3572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5111_6
timestamp 1731220617
transform 1 0 1520 0 -1 3572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5110_6
timestamp 1731220617
transform 1 0 1416 0 -1 3572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5109_6
timestamp 1731220617
transform 1 0 1304 0 -1 3572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5108_6
timestamp 1731220617
transform 1 0 1184 0 -1 3572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5107_6
timestamp 1731220617
transform 1 0 1064 0 -1 3572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5106_6
timestamp 1731220617
transform 1 0 928 0 -1 3572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5105_6
timestamp 1731220617
transform 1 0 784 0 -1 3572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5104_6
timestamp 1731220617
transform 1 0 1416 0 1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5103_6
timestamp 1731220617
transform 1 0 1304 0 1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5102_6
timestamp 1731220617
transform 1 0 1192 0 1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5101_6
timestamp 1731220617
transform 1 0 1072 0 1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5100_6
timestamp 1731220617
transform 1 0 936 0 1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_599_6
timestamp 1731220617
transform 1 0 792 0 1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_598_6
timestamp 1731220617
transform 1 0 1720 0 -1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_597_6
timestamp 1731220617
transform 1 0 1560 0 -1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_596_6
timestamp 1731220617
transform 1 0 1392 0 -1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_595_6
timestamp 1731220617
transform 1 0 1216 0 -1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_594_6
timestamp 1731220617
transform 1 0 1032 0 -1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_593_6
timestamp 1731220617
transform 1 0 1624 0 1 3292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_592_6
timestamp 1731220617
transform 1 0 1472 0 1 3292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_591_6
timestamp 1731220617
transform 1 0 1320 0 1 3292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_590_6
timestamp 1731220617
transform 1 0 1168 0 1 3292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_589_6
timestamp 1731220617
transform 1 0 1016 0 1 3292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_588_6
timestamp 1731220617
transform 1 0 1480 0 -1 3288
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_587_6
timestamp 1731220617
transform 1 0 1328 0 -1 3288
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_586_6
timestamp 1731220617
transform 1 0 1184 0 -1 3288
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_585_6
timestamp 1731220617
transform 1 0 1040 0 -1 3288
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_584_6
timestamp 1731220617
transform 1 0 888 0 -1 3288
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_583_6
timestamp 1731220617
transform 1 0 1336 0 1 3140
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_582_6
timestamp 1731220617
transform 1 0 1176 0 1 3140
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_581_6
timestamp 1731220617
transform 1 0 1024 0 1 3140
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_580_6
timestamp 1731220617
transform 1 0 872 0 1 3140
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_579_6
timestamp 1731220617
transform 1 0 712 0 1 3140
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_578_6
timestamp 1731220617
transform 1 0 1272 0 -1 3128
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_577_6
timestamp 1731220617
transform 1 0 1168 0 -1 3128
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_576_6
timestamp 1731220617
transform 1 0 1064 0 -1 3128
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_575_6
timestamp 1731220617
transform 1 0 960 0 -1 3128
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_574_6
timestamp 1731220617
transform 1 0 856 0 -1 3128
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_573_6
timestamp 1731220617
transform 1 0 1272 0 1 2992
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_572_6
timestamp 1731220617
transform 1 0 1168 0 1 2992
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_571_6
timestamp 1731220617
transform 1 0 1072 0 1 2992
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_570_6
timestamp 1731220617
transform 1 0 976 0 1 2992
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_569_6
timestamp 1731220617
transform 1 0 920 0 -1 2980
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_568_6
timestamp 1731220617
transform 1 0 880 0 1 2992
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_567_6
timestamp 1731220617
transform 1 0 784 0 1 2992
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_566_6
timestamp 1731220617
transform 1 0 688 0 1 2992
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_565_6
timestamp 1731220617
transform 1 0 584 0 1 2992
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_564_6
timestamp 1731220617
transform 1 0 752 0 -1 3128
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_563_6
timestamp 1731220617
transform 1 0 640 0 -1 3128
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_562_6
timestamp 1731220617
transform 1 0 520 0 -1 3128
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_561_6
timestamp 1731220617
transform 1 0 392 0 -1 3128
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_560_6
timestamp 1731220617
transform 1 0 352 0 1 2992
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_559_6
timestamp 1731220617
transform 1 0 472 0 1 2992
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_558_6
timestamp 1731220617
transform 1 0 448 0 -1 2980
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_557_6
timestamp 1731220617
transform 1 0 776 0 -1 2980
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_556_6
timestamp 1731220617
transform 1 0 616 0 -1 2980
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_555_6
timestamp 1731220617
transform 1 0 504 0 1 2844
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_554_6
timestamp 1731220617
transform 1 0 696 0 1 2844
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_553_6
timestamp 1731220617
transform 1 0 880 0 1 2844
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_552_6
timestamp 1731220617
transform 1 0 816 0 -1 2840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_551_6
timestamp 1731220617
transform 1 0 648 0 -1 2840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_550_6
timestamp 1731220617
transform 1 0 480 0 -1 2840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_549_6
timestamp 1731220617
transform 1 0 456 0 1 2696
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_548_6
timestamp 1731220617
transform 1 0 736 0 1 2696
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_547_6
timestamp 1731220617
transform 1 0 592 0 1 2696
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_546_6
timestamp 1731220617
transform 1 0 576 0 -1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_545_6
timestamp 1731220617
transform 1 0 456 0 -1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_544_6
timestamp 1731220617
transform 1 0 328 0 -1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_543_6
timestamp 1731220617
transform 1 0 208 0 -1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_542_6
timestamp 1731220617
transform 1 0 192 0 1 2696
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_541_6
timestamp 1731220617
transform 1 0 320 0 1 2696
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_540_6
timestamp 1731220617
transform 1 0 312 0 -1 2840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_539_6
timestamp 1731220617
transform 1 0 152 0 -1 2840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_538_6
timestamp 1731220617
transform 1 0 128 0 1 2844
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_537_6
timestamp 1731220617
transform 1 0 304 0 1 2844
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_536_6
timestamp 1731220617
transform 1 0 280 0 -1 2980
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_535_6
timestamp 1731220617
transform 1 0 128 0 -1 2980
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_534_6
timestamp 1731220617
transform 1 0 128 0 1 2992
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_533_6
timestamp 1731220617
transform 1 0 232 0 1 2992
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_532_6
timestamp 1731220617
transform 1 0 256 0 -1 3128
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_531_6
timestamp 1731220617
transform 1 0 128 0 -1 3128
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_530_6
timestamp 1731220617
transform 1 0 160 0 1 3140
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_529_6
timestamp 1731220617
transform 1 0 360 0 1 3140
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_528_6
timestamp 1731220617
transform 1 0 544 0 1 3140
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_527_6
timestamp 1731220617
transform 1 0 400 0 -1 3288
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_526_6
timestamp 1731220617
transform 1 0 232 0 -1 3288
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_525_6
timestamp 1731220617
transform 1 0 568 0 -1 3288
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_524_6
timestamp 1731220617
transform 1 0 736 0 -1 3288
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_523_6
timestamp 1731220617
transform 1 0 856 0 1 3292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_522_6
timestamp 1731220617
transform 1 0 696 0 1 3292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_521_6
timestamp 1731220617
transform 1 0 528 0 1 3292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_520_6
timestamp 1731220617
transform 1 0 368 0 1 3292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_519_6
timestamp 1731220617
transform 1 0 224 0 1 3292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_518_6
timestamp 1731220617
transform 1 0 840 0 -1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_517_6
timestamp 1731220617
transform 1 0 632 0 -1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_516_6
timestamp 1731220617
transform 1 0 424 0 -1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_515_6
timestamp 1731220617
transform 1 0 208 0 -1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_514_6
timestamp 1731220617
transform 1 0 640 0 1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_513_6
timestamp 1731220617
transform 1 0 480 0 1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_512_6
timestamp 1731220617
transform 1 0 312 0 1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_511_6
timestamp 1731220617
transform 1 0 136 0 1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_510_6
timestamp 1731220617
transform 1 0 624 0 -1 3572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_59_6
timestamp 1731220617
transform 1 0 456 0 -1 3572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_58_6
timestamp 1731220617
transform 1 0 280 0 -1 3572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_57_6
timestamp 1731220617
transform 1 0 128 0 -1 3572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_56_6
timestamp 1731220617
transform 1 0 656 0 1 3580
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_55_6
timestamp 1731220617
transform 1 0 568 0 1 3580
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_54_6
timestamp 1731220617
transform 1 0 480 0 1 3580
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_53_6
timestamp 1731220617
transform 1 0 392 0 1 3580
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_52_6
timestamp 1731220617
transform 1 0 304 0 1 3580
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_51_6
timestamp 1731220617
transform 1 0 216 0 1 3580
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_50_6
timestamp 1731220617
transform 1 0 128 0 1 3580
box 8 4 80 64
<< end >>
