magic
tech TSMC180
timestamp 1734111263
<< ndiffusion >>
rect 6 21 12 22
rect 6 19 8 21
rect 10 19 12 21
rect 6 12 12 19
rect 14 12 20 22
rect 22 17 28 22
rect 30 21 36 22
rect 30 19 33 21
rect 35 19 36 21
rect 30 17 36 19
rect 22 15 26 17
rect 22 13 23 15
rect 25 13 26 15
rect 22 12 26 13
<< ndcontact >>
rect 8 19 10 21
rect 33 19 35 21
rect 23 13 25 15
<< ntransistor >>
rect 12 12 14 22
rect 20 12 22 22
rect 28 17 30 22
<< pdiffusion >>
rect 6 45 12 46
rect 6 43 7 45
rect 9 43 12 45
rect 6 38 12 43
rect 14 41 20 46
rect 14 39 15 41
rect 17 39 20 41
rect 14 38 20 39
rect 22 45 28 46
rect 22 43 23 45
rect 25 43 28 45
rect 22 38 28 43
rect 30 41 36 46
rect 30 39 33 41
rect 35 39 36 41
rect 30 38 36 39
<< pdcontact >>
rect 7 43 9 45
rect 15 39 17 41
rect 23 43 25 45
rect 33 39 35 41
<< ptransistor >>
rect 12 38 14 46
rect 20 38 22 46
rect 28 38 30 46
<< polysilicon >>
rect 18 53 22 54
rect 18 51 19 53
rect 21 51 22 53
rect 18 50 22 51
rect 12 46 14 49
rect 20 46 22 50
rect 28 46 30 49
rect 12 22 14 38
rect 20 22 22 38
rect 28 31 30 38
rect 28 30 43 31
rect 28 29 40 30
rect 28 22 30 29
rect 39 28 40 29
rect 42 28 43 30
rect 39 27 43 28
rect 28 14 30 17
rect 12 10 14 12
rect 6 9 14 10
rect 20 9 22 12
rect 6 7 7 9
rect 9 8 14 9
rect 9 7 10 8
rect 6 6 10 7
<< polycontact >>
rect 19 51 21 53
rect 40 28 42 30
rect 7 7 9 9
<< m1 >>
rect 6 57 21 60
rect 18 54 21 57
rect 33 57 45 60
rect 18 53 22 54
rect 18 51 19 53
rect 21 51 22 53
rect 18 50 22 51
rect 6 46 11 47
rect 6 43 7 46
rect 10 43 11 46
rect 6 42 11 43
rect 21 46 26 47
rect 21 43 22 46
rect 25 43 26 46
rect 21 42 26 43
rect 33 42 36 57
rect 14 41 18 42
rect 14 39 15 41
rect 17 39 18 41
rect 14 38 18 39
rect 32 41 36 42
rect 32 39 33 41
rect 35 39 36 41
rect 32 38 36 39
rect 14 32 17 38
rect 6 31 11 32
rect 6 28 7 31
rect 10 28 11 31
rect 6 27 11 28
rect 14 31 19 32
rect 14 28 15 31
rect 18 28 19 31
rect 14 27 19 28
rect 8 22 11 27
rect 33 22 36 38
rect 39 31 44 32
rect 39 28 40 31
rect 43 28 44 31
rect 39 27 44 28
rect 7 21 11 22
rect 7 19 8 21
rect 10 19 11 21
rect 7 18 11 19
rect 32 21 36 22
rect 32 19 33 21
rect 35 19 36 21
rect 32 18 36 19
rect 21 15 26 16
rect 21 12 22 15
rect 25 12 26 15
rect 21 11 26 12
rect 6 9 10 10
rect 6 7 7 9
rect 9 7 10 9
rect 6 6 10 7
rect 6 1 9 6
<< m2c >>
rect 7 45 10 46
rect 7 43 9 45
rect 9 43 10 45
rect 22 45 25 46
rect 22 43 23 45
rect 23 43 25 45
rect 7 28 10 31
rect 15 28 18 31
rect 40 30 43 31
rect 40 28 42 30
rect 42 28 43 30
rect 22 13 23 15
rect 23 13 25 15
rect 22 12 25 13
<< m2 >>
rect -5 46 26 47
rect -5 43 7 46
rect 10 43 22 46
rect 25 43 26 46
rect -5 42 26 43
rect 6 31 44 32
rect 6 28 7 31
rect 10 28 15 31
rect 18 28 40 31
rect 43 28 44 31
rect 6 27 44 28
rect 21 15 26 16
rect 21 12 22 15
rect 25 12 26 15
rect 21 0 26 12
<< labels >>
rlabel ndiffusion 31 18 31 18 3 Y
rlabel polysilicon 29 23 29 23 3 _Y
rlabel polysilicon 29 36 29 36 3 _Y
rlabel pdiffusion 31 39 31 39 3 Y
rlabel ndiffusion 23 13 23 13 3 GND
rlabel pdiffusion 23 39 23 39 3 Vdd
rlabel polysilicon 21 23 21 23 3 A
rlabel polysilicon 21 36 21 36 3 A
rlabel pdiffusion 15 39 15 39 3 _Y
rlabel polysilicon 13 23 13 23 3 B
rlabel polysilicon 13 36 13 36 3 B
rlabel ndiffusion 7 13 7 13 3 _Y
rlabel pdiffusion 7 39 7 39 3 Vdd
rlabel m1 7 58 7 58 3 A
port 5 e
rlabel m2 -4 43 -4 43 3 Vdd
rlabel m2 22 1 22 1 1 GND
rlabel m1 43 58 43 58 3 Y
rlabel m1 7 2 7 2 3 B
<< end >>
