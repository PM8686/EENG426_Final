magic
tech sky130l
timestamp 1731220637
<< m2 >>
rect 230 2479 236 2480
rect 230 2475 231 2479
rect 235 2475 236 2479
rect 230 2474 236 2475
rect 270 2479 276 2480
rect 270 2475 271 2479
rect 275 2475 276 2479
rect 270 2474 276 2475
rect 310 2479 316 2480
rect 310 2475 311 2479
rect 315 2475 316 2479
rect 310 2474 316 2475
rect 350 2479 356 2480
rect 350 2475 351 2479
rect 355 2475 356 2479
rect 350 2474 356 2475
rect 398 2479 404 2480
rect 398 2475 399 2479
rect 403 2475 404 2479
rect 398 2474 404 2475
rect 454 2479 460 2480
rect 454 2475 455 2479
rect 459 2475 460 2479
rect 454 2474 460 2475
rect 510 2479 516 2480
rect 510 2475 511 2479
rect 515 2475 516 2479
rect 510 2474 516 2475
rect 574 2479 580 2480
rect 574 2475 575 2479
rect 579 2475 580 2479
rect 574 2474 580 2475
rect 638 2479 644 2480
rect 638 2475 639 2479
rect 643 2475 644 2479
rect 638 2474 644 2475
rect 702 2479 708 2480
rect 702 2475 703 2479
rect 707 2475 708 2479
rect 702 2474 708 2475
rect 766 2479 772 2480
rect 766 2475 767 2479
rect 771 2475 772 2479
rect 766 2474 772 2475
rect 822 2479 828 2480
rect 822 2475 823 2479
rect 827 2475 828 2479
rect 822 2474 828 2475
rect 878 2479 884 2480
rect 878 2475 879 2479
rect 883 2475 884 2479
rect 878 2474 884 2475
rect 926 2479 932 2480
rect 926 2475 927 2479
rect 931 2475 932 2479
rect 926 2474 932 2475
rect 974 2479 980 2480
rect 974 2475 975 2479
rect 979 2475 980 2479
rect 974 2474 980 2475
rect 1022 2479 1028 2480
rect 1022 2475 1023 2479
rect 1027 2475 1028 2479
rect 1022 2474 1028 2475
rect 1070 2479 1076 2480
rect 1070 2475 1071 2479
rect 1075 2475 1076 2479
rect 1070 2474 1076 2475
rect 1110 2479 1116 2480
rect 1110 2475 1111 2479
rect 1115 2475 1116 2479
rect 1110 2474 1116 2475
rect 1150 2479 1156 2480
rect 1150 2475 1151 2479
rect 1155 2475 1156 2479
rect 1150 2474 1156 2475
rect 1190 2479 1196 2480
rect 1190 2475 1191 2479
rect 1195 2475 1196 2479
rect 1190 2474 1196 2475
rect 1302 2475 1308 2476
rect 1302 2471 1303 2475
rect 1307 2471 1308 2475
rect 1302 2470 1308 2471
rect 1342 2475 1348 2476
rect 1342 2471 1343 2475
rect 1347 2471 1348 2475
rect 1342 2470 1348 2471
rect 1382 2475 1388 2476
rect 1382 2471 1383 2475
rect 1387 2471 1388 2475
rect 1382 2470 1388 2471
rect 1438 2475 1444 2476
rect 1438 2471 1439 2475
rect 1443 2471 1444 2475
rect 1438 2470 1444 2471
rect 1510 2475 1516 2476
rect 1510 2471 1511 2475
rect 1515 2471 1516 2475
rect 1510 2470 1516 2471
rect 1582 2475 1588 2476
rect 1582 2471 1583 2475
rect 1587 2471 1588 2475
rect 1582 2470 1588 2471
rect 1662 2475 1668 2476
rect 1662 2471 1663 2475
rect 1667 2471 1668 2475
rect 1662 2470 1668 2471
rect 1734 2475 1740 2476
rect 1734 2471 1735 2475
rect 1739 2471 1740 2475
rect 1734 2470 1740 2471
rect 1806 2475 1812 2476
rect 1806 2471 1807 2475
rect 1811 2471 1812 2475
rect 1806 2470 1812 2471
rect 1886 2475 1892 2476
rect 1886 2471 1887 2475
rect 1891 2471 1892 2475
rect 1886 2470 1892 2471
rect 1966 2475 1972 2476
rect 1966 2471 1967 2475
rect 1971 2471 1972 2475
rect 1966 2470 1972 2471
rect 2062 2475 2068 2476
rect 2062 2471 2063 2475
rect 2067 2471 2068 2475
rect 2062 2470 2068 2471
rect 2166 2475 2172 2476
rect 2166 2471 2167 2475
rect 2171 2471 2172 2475
rect 2166 2470 2172 2471
rect 2270 2475 2276 2476
rect 2270 2471 2271 2475
rect 2275 2471 2276 2475
rect 2270 2470 2276 2471
rect 2358 2475 2364 2476
rect 2358 2471 2359 2475
rect 2363 2471 2364 2475
rect 2358 2470 2364 2471
rect 110 2456 116 2457
rect 110 2452 111 2456
rect 115 2452 116 2456
rect 110 2451 116 2452
rect 1238 2456 1244 2457
rect 1238 2452 1239 2456
rect 1243 2452 1244 2456
rect 1238 2451 1244 2452
rect 1278 2452 1284 2453
rect 1278 2448 1279 2452
rect 1283 2448 1284 2452
rect 1278 2447 1284 2448
rect 2406 2452 2412 2453
rect 2406 2448 2407 2452
rect 2411 2448 2412 2452
rect 2406 2447 2412 2448
rect 110 2439 116 2440
rect 110 2435 111 2439
rect 115 2435 116 2439
rect 110 2434 116 2435
rect 1238 2439 1244 2440
rect 1238 2435 1239 2439
rect 1243 2435 1244 2439
rect 1238 2434 1244 2435
rect 1278 2435 1284 2436
rect 230 2432 236 2433
rect 230 2428 231 2432
rect 235 2428 236 2432
rect 230 2427 236 2428
rect 270 2432 276 2433
rect 270 2428 271 2432
rect 275 2428 276 2432
rect 270 2427 276 2428
rect 310 2432 316 2433
rect 310 2428 311 2432
rect 315 2428 316 2432
rect 310 2427 316 2428
rect 350 2432 356 2433
rect 350 2428 351 2432
rect 355 2428 356 2432
rect 350 2427 356 2428
rect 398 2432 404 2433
rect 398 2428 399 2432
rect 403 2428 404 2432
rect 398 2427 404 2428
rect 454 2432 460 2433
rect 454 2428 455 2432
rect 459 2428 460 2432
rect 454 2427 460 2428
rect 510 2432 516 2433
rect 510 2428 511 2432
rect 515 2428 516 2432
rect 510 2427 516 2428
rect 574 2432 580 2433
rect 574 2428 575 2432
rect 579 2428 580 2432
rect 574 2427 580 2428
rect 638 2432 644 2433
rect 638 2428 639 2432
rect 643 2428 644 2432
rect 638 2427 644 2428
rect 702 2432 708 2433
rect 702 2428 703 2432
rect 707 2428 708 2432
rect 702 2427 708 2428
rect 766 2432 772 2433
rect 766 2428 767 2432
rect 771 2428 772 2432
rect 766 2427 772 2428
rect 822 2432 828 2433
rect 822 2428 823 2432
rect 827 2428 828 2432
rect 822 2427 828 2428
rect 878 2432 884 2433
rect 878 2428 879 2432
rect 883 2428 884 2432
rect 878 2427 884 2428
rect 926 2432 932 2433
rect 926 2428 927 2432
rect 931 2428 932 2432
rect 926 2427 932 2428
rect 974 2432 980 2433
rect 974 2428 975 2432
rect 979 2428 980 2432
rect 974 2427 980 2428
rect 1022 2432 1028 2433
rect 1022 2428 1023 2432
rect 1027 2428 1028 2432
rect 1022 2427 1028 2428
rect 1070 2432 1076 2433
rect 1070 2428 1071 2432
rect 1075 2428 1076 2432
rect 1070 2427 1076 2428
rect 1110 2432 1116 2433
rect 1110 2428 1111 2432
rect 1115 2428 1116 2432
rect 1110 2427 1116 2428
rect 1150 2432 1156 2433
rect 1150 2428 1151 2432
rect 1155 2428 1156 2432
rect 1150 2427 1156 2428
rect 1190 2432 1196 2433
rect 1190 2428 1191 2432
rect 1195 2428 1196 2432
rect 1278 2431 1279 2435
rect 1283 2431 1284 2435
rect 1278 2430 1284 2431
rect 2406 2435 2412 2436
rect 2406 2431 2407 2435
rect 2411 2431 2412 2435
rect 2406 2430 2412 2431
rect 1190 2427 1196 2428
rect 1302 2428 1308 2429
rect 1302 2424 1303 2428
rect 1307 2424 1308 2428
rect 1302 2423 1308 2424
rect 1342 2428 1348 2429
rect 1342 2424 1343 2428
rect 1347 2424 1348 2428
rect 1342 2423 1348 2424
rect 1382 2428 1388 2429
rect 1382 2424 1383 2428
rect 1387 2424 1388 2428
rect 1382 2423 1388 2424
rect 1438 2428 1444 2429
rect 1438 2424 1439 2428
rect 1443 2424 1444 2428
rect 1438 2423 1444 2424
rect 1510 2428 1516 2429
rect 1510 2424 1511 2428
rect 1515 2424 1516 2428
rect 1510 2423 1516 2424
rect 1582 2428 1588 2429
rect 1582 2424 1583 2428
rect 1587 2424 1588 2428
rect 1582 2423 1588 2424
rect 1662 2428 1668 2429
rect 1662 2424 1663 2428
rect 1667 2424 1668 2428
rect 1662 2423 1668 2424
rect 1734 2428 1740 2429
rect 1734 2424 1735 2428
rect 1739 2424 1740 2428
rect 1734 2423 1740 2424
rect 1806 2428 1812 2429
rect 1806 2424 1807 2428
rect 1811 2424 1812 2428
rect 1806 2423 1812 2424
rect 1886 2428 1892 2429
rect 1886 2424 1887 2428
rect 1891 2424 1892 2428
rect 1886 2423 1892 2424
rect 1966 2428 1972 2429
rect 1966 2424 1967 2428
rect 1971 2424 1972 2428
rect 1966 2423 1972 2424
rect 2062 2428 2068 2429
rect 2062 2424 2063 2428
rect 2067 2424 2068 2428
rect 2062 2423 2068 2424
rect 2166 2428 2172 2429
rect 2166 2424 2167 2428
rect 2171 2424 2172 2428
rect 2166 2423 2172 2424
rect 2270 2428 2276 2429
rect 2270 2424 2271 2428
rect 2275 2424 2276 2428
rect 2270 2423 2276 2424
rect 2358 2428 2364 2429
rect 2358 2424 2359 2428
rect 2363 2424 2364 2428
rect 2358 2423 2364 2424
rect 1374 2416 1380 2417
rect 198 2412 204 2413
rect 198 2408 199 2412
rect 203 2408 204 2412
rect 198 2407 204 2408
rect 262 2412 268 2413
rect 262 2408 263 2412
rect 267 2408 268 2412
rect 262 2407 268 2408
rect 326 2412 332 2413
rect 326 2408 327 2412
rect 331 2408 332 2412
rect 326 2407 332 2408
rect 398 2412 404 2413
rect 398 2408 399 2412
rect 403 2408 404 2412
rect 398 2407 404 2408
rect 470 2412 476 2413
rect 470 2408 471 2412
rect 475 2408 476 2412
rect 470 2407 476 2408
rect 542 2412 548 2413
rect 542 2408 543 2412
rect 547 2408 548 2412
rect 542 2407 548 2408
rect 614 2412 620 2413
rect 614 2408 615 2412
rect 619 2408 620 2412
rect 614 2407 620 2408
rect 686 2412 692 2413
rect 686 2408 687 2412
rect 691 2408 692 2412
rect 686 2407 692 2408
rect 750 2412 756 2413
rect 750 2408 751 2412
rect 755 2408 756 2412
rect 750 2407 756 2408
rect 822 2412 828 2413
rect 822 2408 823 2412
rect 827 2408 828 2412
rect 822 2407 828 2408
rect 894 2412 900 2413
rect 894 2408 895 2412
rect 899 2408 900 2412
rect 894 2407 900 2408
rect 966 2412 972 2413
rect 966 2408 967 2412
rect 971 2408 972 2412
rect 1374 2412 1375 2416
rect 1379 2412 1380 2416
rect 1374 2411 1380 2412
rect 1414 2416 1420 2417
rect 1414 2412 1415 2416
rect 1419 2412 1420 2416
rect 1414 2411 1420 2412
rect 1454 2416 1460 2417
rect 1454 2412 1455 2416
rect 1459 2412 1460 2416
rect 1454 2411 1460 2412
rect 1502 2416 1508 2417
rect 1502 2412 1503 2416
rect 1507 2412 1508 2416
rect 1502 2411 1508 2412
rect 1558 2416 1564 2417
rect 1558 2412 1559 2416
rect 1563 2412 1564 2416
rect 1558 2411 1564 2412
rect 1614 2416 1620 2417
rect 1614 2412 1615 2416
rect 1619 2412 1620 2416
rect 1614 2411 1620 2412
rect 1678 2416 1684 2417
rect 1678 2412 1679 2416
rect 1683 2412 1684 2416
rect 1678 2411 1684 2412
rect 1734 2416 1740 2417
rect 1734 2412 1735 2416
rect 1739 2412 1740 2416
rect 1734 2411 1740 2412
rect 1798 2416 1804 2417
rect 1798 2412 1799 2416
rect 1803 2412 1804 2416
rect 1798 2411 1804 2412
rect 1870 2416 1876 2417
rect 1870 2412 1871 2416
rect 1875 2412 1876 2416
rect 1870 2411 1876 2412
rect 1950 2416 1956 2417
rect 1950 2412 1951 2416
rect 1955 2412 1956 2416
rect 1950 2411 1956 2412
rect 2046 2416 2052 2417
rect 2046 2412 2047 2416
rect 2051 2412 2052 2416
rect 2046 2411 2052 2412
rect 2150 2416 2156 2417
rect 2150 2412 2151 2416
rect 2155 2412 2156 2416
rect 2150 2411 2156 2412
rect 2262 2416 2268 2417
rect 2262 2412 2263 2416
rect 2267 2412 2268 2416
rect 2262 2411 2268 2412
rect 2358 2416 2364 2417
rect 2358 2412 2359 2416
rect 2363 2412 2364 2416
rect 2358 2411 2364 2412
rect 966 2407 972 2408
rect 1278 2409 1284 2410
rect 110 2405 116 2406
rect 110 2401 111 2405
rect 115 2401 116 2405
rect 110 2400 116 2401
rect 1238 2405 1244 2406
rect 1238 2401 1239 2405
rect 1243 2401 1244 2405
rect 1278 2405 1279 2409
rect 1283 2405 1284 2409
rect 1278 2404 1284 2405
rect 2406 2409 2412 2410
rect 2406 2405 2407 2409
rect 2411 2405 2412 2409
rect 2406 2404 2412 2405
rect 1238 2400 1244 2401
rect 1278 2392 1284 2393
rect 110 2388 116 2389
rect 110 2384 111 2388
rect 115 2384 116 2388
rect 110 2383 116 2384
rect 1238 2388 1244 2389
rect 1238 2384 1239 2388
rect 1243 2384 1244 2388
rect 1278 2388 1279 2392
rect 1283 2388 1284 2392
rect 1278 2387 1284 2388
rect 2406 2392 2412 2393
rect 2406 2388 2407 2392
rect 2411 2388 2412 2392
rect 2406 2387 2412 2388
rect 1238 2383 1244 2384
rect 1374 2369 1380 2370
rect 198 2365 204 2366
rect 198 2361 199 2365
rect 203 2361 204 2365
rect 198 2360 204 2361
rect 262 2365 268 2366
rect 262 2361 263 2365
rect 267 2361 268 2365
rect 262 2360 268 2361
rect 326 2365 332 2366
rect 326 2361 327 2365
rect 331 2361 332 2365
rect 326 2360 332 2361
rect 398 2365 404 2366
rect 398 2361 399 2365
rect 403 2361 404 2365
rect 398 2360 404 2361
rect 470 2365 476 2366
rect 470 2361 471 2365
rect 475 2361 476 2365
rect 470 2360 476 2361
rect 542 2365 548 2366
rect 542 2361 543 2365
rect 547 2361 548 2365
rect 542 2360 548 2361
rect 614 2365 620 2366
rect 614 2361 615 2365
rect 619 2361 620 2365
rect 614 2360 620 2361
rect 686 2365 692 2366
rect 686 2361 687 2365
rect 691 2361 692 2365
rect 686 2360 692 2361
rect 750 2365 756 2366
rect 750 2361 751 2365
rect 755 2361 756 2365
rect 750 2360 756 2361
rect 822 2365 828 2366
rect 822 2361 823 2365
rect 827 2361 828 2365
rect 822 2360 828 2361
rect 894 2365 900 2366
rect 894 2361 895 2365
rect 899 2361 900 2365
rect 894 2360 900 2361
rect 966 2365 972 2366
rect 966 2361 967 2365
rect 971 2361 972 2365
rect 1374 2365 1375 2369
rect 1379 2365 1380 2369
rect 1374 2364 1380 2365
rect 1414 2369 1420 2370
rect 1414 2365 1415 2369
rect 1419 2365 1420 2369
rect 1414 2364 1420 2365
rect 1454 2369 1460 2370
rect 1454 2365 1455 2369
rect 1459 2365 1460 2369
rect 1454 2364 1460 2365
rect 1502 2369 1508 2370
rect 1502 2365 1503 2369
rect 1507 2365 1508 2369
rect 1502 2364 1508 2365
rect 1558 2369 1564 2370
rect 1558 2365 1559 2369
rect 1563 2365 1564 2369
rect 1558 2364 1564 2365
rect 1614 2369 1620 2370
rect 1614 2365 1615 2369
rect 1619 2365 1620 2369
rect 1614 2364 1620 2365
rect 1678 2369 1684 2370
rect 1678 2365 1679 2369
rect 1683 2365 1684 2369
rect 1678 2364 1684 2365
rect 1734 2369 1740 2370
rect 1734 2365 1735 2369
rect 1739 2365 1740 2369
rect 1734 2364 1740 2365
rect 1798 2369 1804 2370
rect 1798 2365 1799 2369
rect 1803 2365 1804 2369
rect 1798 2364 1804 2365
rect 1870 2369 1876 2370
rect 1870 2365 1871 2369
rect 1875 2365 1876 2369
rect 1870 2364 1876 2365
rect 1950 2369 1956 2370
rect 1950 2365 1951 2369
rect 1955 2365 1956 2369
rect 1950 2364 1956 2365
rect 2046 2369 2052 2370
rect 2046 2365 2047 2369
rect 2051 2365 2052 2369
rect 2046 2364 2052 2365
rect 2150 2369 2156 2370
rect 2150 2365 2151 2369
rect 2155 2365 2156 2369
rect 2150 2364 2156 2365
rect 2262 2369 2268 2370
rect 2262 2365 2263 2369
rect 2267 2365 2268 2369
rect 2262 2364 2268 2365
rect 2358 2369 2364 2370
rect 2358 2365 2359 2369
rect 2363 2365 2364 2369
rect 2358 2364 2364 2365
rect 966 2360 972 2361
rect 1326 2335 1332 2336
rect 270 2331 276 2332
rect 270 2327 271 2331
rect 275 2327 276 2331
rect 270 2326 276 2327
rect 326 2331 332 2332
rect 326 2327 327 2331
rect 331 2327 332 2331
rect 326 2326 332 2327
rect 398 2331 404 2332
rect 398 2327 399 2331
rect 403 2327 404 2331
rect 398 2326 404 2327
rect 470 2331 476 2332
rect 470 2327 471 2331
rect 475 2327 476 2331
rect 470 2326 476 2327
rect 550 2331 556 2332
rect 550 2327 551 2331
rect 555 2327 556 2331
rect 550 2326 556 2327
rect 630 2331 636 2332
rect 630 2327 631 2331
rect 635 2327 636 2331
rect 630 2326 636 2327
rect 710 2331 716 2332
rect 710 2327 711 2331
rect 715 2327 716 2331
rect 710 2326 716 2327
rect 782 2331 788 2332
rect 782 2327 783 2331
rect 787 2327 788 2331
rect 782 2326 788 2327
rect 854 2331 860 2332
rect 854 2327 855 2331
rect 859 2327 860 2331
rect 854 2326 860 2327
rect 918 2331 924 2332
rect 918 2327 919 2331
rect 923 2327 924 2331
rect 918 2326 924 2327
rect 990 2331 996 2332
rect 990 2327 991 2331
rect 995 2327 996 2331
rect 990 2326 996 2327
rect 1062 2331 1068 2332
rect 1062 2327 1063 2331
rect 1067 2327 1068 2331
rect 1326 2331 1327 2335
rect 1331 2331 1332 2335
rect 1326 2330 1332 2331
rect 1382 2335 1388 2336
rect 1382 2331 1383 2335
rect 1387 2331 1388 2335
rect 1382 2330 1388 2331
rect 1438 2335 1444 2336
rect 1438 2331 1439 2335
rect 1443 2331 1444 2335
rect 1438 2330 1444 2331
rect 1502 2335 1508 2336
rect 1502 2331 1503 2335
rect 1507 2331 1508 2335
rect 1502 2330 1508 2331
rect 1574 2335 1580 2336
rect 1574 2331 1575 2335
rect 1579 2331 1580 2335
rect 1574 2330 1580 2331
rect 1646 2335 1652 2336
rect 1646 2331 1647 2335
rect 1651 2331 1652 2335
rect 1646 2330 1652 2331
rect 1718 2335 1724 2336
rect 1718 2331 1719 2335
rect 1723 2331 1724 2335
rect 1718 2330 1724 2331
rect 1798 2335 1804 2336
rect 1798 2331 1799 2335
rect 1803 2331 1804 2335
rect 1798 2330 1804 2331
rect 1878 2335 1884 2336
rect 1878 2331 1879 2335
rect 1883 2331 1884 2335
rect 1878 2330 1884 2331
rect 1966 2335 1972 2336
rect 1966 2331 1967 2335
rect 1971 2331 1972 2335
rect 1966 2330 1972 2331
rect 2062 2335 2068 2336
rect 2062 2331 2063 2335
rect 2067 2331 2068 2335
rect 2062 2330 2068 2331
rect 2166 2335 2172 2336
rect 2166 2331 2167 2335
rect 2171 2331 2172 2335
rect 2166 2330 2172 2331
rect 2270 2335 2276 2336
rect 2270 2331 2271 2335
rect 2275 2331 2276 2335
rect 2270 2330 2276 2331
rect 2358 2335 2364 2336
rect 2358 2331 2359 2335
rect 2363 2331 2364 2335
rect 2358 2330 2364 2331
rect 1062 2326 1068 2327
rect 1278 2312 1284 2313
rect 110 2308 116 2309
rect 110 2304 111 2308
rect 115 2304 116 2308
rect 110 2303 116 2304
rect 1238 2308 1244 2309
rect 1238 2304 1239 2308
rect 1243 2304 1244 2308
rect 1278 2308 1279 2312
rect 1283 2308 1284 2312
rect 1278 2307 1284 2308
rect 2406 2312 2412 2313
rect 2406 2308 2407 2312
rect 2411 2308 2412 2312
rect 2406 2307 2412 2308
rect 1238 2303 1244 2304
rect 1278 2295 1284 2296
rect 110 2291 116 2292
rect 110 2287 111 2291
rect 115 2287 116 2291
rect 110 2286 116 2287
rect 1238 2291 1244 2292
rect 1238 2287 1239 2291
rect 1243 2287 1244 2291
rect 1278 2291 1279 2295
rect 1283 2291 1284 2295
rect 1278 2290 1284 2291
rect 2406 2295 2412 2296
rect 2406 2291 2407 2295
rect 2411 2291 2412 2295
rect 2406 2290 2412 2291
rect 1238 2286 1244 2287
rect 1326 2288 1332 2289
rect 270 2284 276 2285
rect 270 2280 271 2284
rect 275 2280 276 2284
rect 270 2279 276 2280
rect 326 2284 332 2285
rect 326 2280 327 2284
rect 331 2280 332 2284
rect 326 2279 332 2280
rect 398 2284 404 2285
rect 398 2280 399 2284
rect 403 2280 404 2284
rect 398 2279 404 2280
rect 470 2284 476 2285
rect 470 2280 471 2284
rect 475 2280 476 2284
rect 470 2279 476 2280
rect 550 2284 556 2285
rect 550 2280 551 2284
rect 555 2280 556 2284
rect 550 2279 556 2280
rect 630 2284 636 2285
rect 630 2280 631 2284
rect 635 2280 636 2284
rect 630 2279 636 2280
rect 710 2284 716 2285
rect 710 2280 711 2284
rect 715 2280 716 2284
rect 710 2279 716 2280
rect 782 2284 788 2285
rect 782 2280 783 2284
rect 787 2280 788 2284
rect 782 2279 788 2280
rect 854 2284 860 2285
rect 854 2280 855 2284
rect 859 2280 860 2284
rect 854 2279 860 2280
rect 918 2284 924 2285
rect 918 2280 919 2284
rect 923 2280 924 2284
rect 918 2279 924 2280
rect 990 2284 996 2285
rect 990 2280 991 2284
rect 995 2280 996 2284
rect 990 2279 996 2280
rect 1062 2284 1068 2285
rect 1062 2280 1063 2284
rect 1067 2280 1068 2284
rect 1326 2284 1327 2288
rect 1331 2284 1332 2288
rect 1326 2283 1332 2284
rect 1382 2288 1388 2289
rect 1382 2284 1383 2288
rect 1387 2284 1388 2288
rect 1382 2283 1388 2284
rect 1438 2288 1444 2289
rect 1438 2284 1439 2288
rect 1443 2284 1444 2288
rect 1438 2283 1444 2284
rect 1502 2288 1508 2289
rect 1502 2284 1503 2288
rect 1507 2284 1508 2288
rect 1502 2283 1508 2284
rect 1574 2288 1580 2289
rect 1574 2284 1575 2288
rect 1579 2284 1580 2288
rect 1574 2283 1580 2284
rect 1646 2288 1652 2289
rect 1646 2284 1647 2288
rect 1651 2284 1652 2288
rect 1646 2283 1652 2284
rect 1718 2288 1724 2289
rect 1718 2284 1719 2288
rect 1723 2284 1724 2288
rect 1718 2283 1724 2284
rect 1798 2288 1804 2289
rect 1798 2284 1799 2288
rect 1803 2284 1804 2288
rect 1798 2283 1804 2284
rect 1878 2288 1884 2289
rect 1878 2284 1879 2288
rect 1883 2284 1884 2288
rect 1878 2283 1884 2284
rect 1966 2288 1972 2289
rect 1966 2284 1967 2288
rect 1971 2284 1972 2288
rect 1966 2283 1972 2284
rect 2062 2288 2068 2289
rect 2062 2284 2063 2288
rect 2067 2284 2068 2288
rect 2062 2283 2068 2284
rect 2166 2288 2172 2289
rect 2166 2284 2167 2288
rect 2171 2284 2172 2288
rect 2166 2283 2172 2284
rect 2270 2288 2276 2289
rect 2270 2284 2271 2288
rect 2275 2284 2276 2288
rect 2270 2283 2276 2284
rect 2358 2288 2364 2289
rect 2358 2284 2359 2288
rect 2363 2284 2364 2288
rect 2358 2283 2364 2284
rect 1062 2279 1068 2280
rect 1334 2276 1340 2277
rect 1334 2272 1335 2276
rect 1339 2272 1340 2276
rect 1334 2271 1340 2272
rect 1406 2276 1412 2277
rect 1406 2272 1407 2276
rect 1411 2272 1412 2276
rect 1406 2271 1412 2272
rect 1486 2276 1492 2277
rect 1486 2272 1487 2276
rect 1491 2272 1492 2276
rect 1486 2271 1492 2272
rect 1558 2276 1564 2277
rect 1558 2272 1559 2276
rect 1563 2272 1564 2276
rect 1558 2271 1564 2272
rect 1630 2276 1636 2277
rect 1630 2272 1631 2276
rect 1635 2272 1636 2276
rect 1630 2271 1636 2272
rect 1702 2276 1708 2277
rect 1702 2272 1703 2276
rect 1707 2272 1708 2276
rect 1702 2271 1708 2272
rect 1774 2276 1780 2277
rect 1774 2272 1775 2276
rect 1779 2272 1780 2276
rect 1774 2271 1780 2272
rect 1838 2276 1844 2277
rect 1838 2272 1839 2276
rect 1843 2272 1844 2276
rect 1838 2271 1844 2272
rect 1910 2276 1916 2277
rect 1910 2272 1911 2276
rect 1915 2272 1916 2276
rect 1910 2271 1916 2272
rect 1990 2276 1996 2277
rect 1990 2272 1991 2276
rect 1995 2272 1996 2276
rect 1990 2271 1996 2272
rect 2078 2276 2084 2277
rect 2078 2272 2079 2276
rect 2083 2272 2084 2276
rect 2078 2271 2084 2272
rect 2174 2276 2180 2277
rect 2174 2272 2175 2276
rect 2179 2272 2180 2276
rect 2174 2271 2180 2272
rect 2278 2276 2284 2277
rect 2278 2272 2279 2276
rect 2283 2272 2284 2276
rect 2278 2271 2284 2272
rect 2358 2276 2364 2277
rect 2358 2272 2359 2276
rect 2363 2272 2364 2276
rect 2358 2271 2364 2272
rect 1278 2269 1284 2270
rect 1278 2265 1279 2269
rect 1283 2265 1284 2269
rect 142 2264 148 2265
rect 142 2260 143 2264
rect 147 2260 148 2264
rect 142 2259 148 2260
rect 182 2264 188 2265
rect 182 2260 183 2264
rect 187 2260 188 2264
rect 182 2259 188 2260
rect 222 2264 228 2265
rect 222 2260 223 2264
rect 227 2260 228 2264
rect 222 2259 228 2260
rect 278 2264 284 2265
rect 278 2260 279 2264
rect 283 2260 284 2264
rect 278 2259 284 2260
rect 334 2264 340 2265
rect 334 2260 335 2264
rect 339 2260 340 2264
rect 334 2259 340 2260
rect 406 2264 412 2265
rect 406 2260 407 2264
rect 411 2260 412 2264
rect 406 2259 412 2260
rect 478 2264 484 2265
rect 478 2260 479 2264
rect 483 2260 484 2264
rect 478 2259 484 2260
rect 558 2264 564 2265
rect 558 2260 559 2264
rect 563 2260 564 2264
rect 558 2259 564 2260
rect 646 2264 652 2265
rect 646 2260 647 2264
rect 651 2260 652 2264
rect 646 2259 652 2260
rect 726 2264 732 2265
rect 726 2260 727 2264
rect 731 2260 732 2264
rect 726 2259 732 2260
rect 806 2264 812 2265
rect 806 2260 807 2264
rect 811 2260 812 2264
rect 806 2259 812 2260
rect 886 2264 892 2265
rect 886 2260 887 2264
rect 891 2260 892 2264
rect 886 2259 892 2260
rect 966 2264 972 2265
rect 966 2260 967 2264
rect 971 2260 972 2264
rect 966 2259 972 2260
rect 1046 2264 1052 2265
rect 1046 2260 1047 2264
rect 1051 2260 1052 2264
rect 1046 2259 1052 2260
rect 1126 2264 1132 2265
rect 1278 2264 1284 2265
rect 2406 2269 2412 2270
rect 2406 2265 2407 2269
rect 2411 2265 2412 2269
rect 2406 2264 2412 2265
rect 1126 2260 1127 2264
rect 1131 2260 1132 2264
rect 1126 2259 1132 2260
rect 110 2257 116 2258
rect 110 2253 111 2257
rect 115 2253 116 2257
rect 110 2252 116 2253
rect 1238 2257 1244 2258
rect 1238 2253 1239 2257
rect 1243 2253 1244 2257
rect 1238 2252 1244 2253
rect 1278 2252 1284 2253
rect 1278 2248 1279 2252
rect 1283 2248 1284 2252
rect 1278 2247 1284 2248
rect 2406 2252 2412 2253
rect 2406 2248 2407 2252
rect 2411 2248 2412 2252
rect 2406 2247 2412 2248
rect 110 2240 116 2241
rect 110 2236 111 2240
rect 115 2236 116 2240
rect 110 2235 116 2236
rect 1238 2240 1244 2241
rect 1238 2236 1239 2240
rect 1243 2236 1244 2240
rect 1238 2235 1244 2236
rect 1334 2229 1340 2230
rect 1334 2225 1335 2229
rect 1339 2225 1340 2229
rect 1334 2224 1340 2225
rect 1406 2229 1412 2230
rect 1406 2225 1407 2229
rect 1411 2225 1412 2229
rect 1406 2224 1412 2225
rect 1486 2229 1492 2230
rect 1486 2225 1487 2229
rect 1491 2225 1492 2229
rect 1486 2224 1492 2225
rect 1558 2229 1564 2230
rect 1558 2225 1559 2229
rect 1563 2225 1564 2229
rect 1558 2224 1564 2225
rect 1630 2229 1636 2230
rect 1630 2225 1631 2229
rect 1635 2225 1636 2229
rect 1630 2224 1636 2225
rect 1702 2229 1708 2230
rect 1702 2225 1703 2229
rect 1707 2225 1708 2229
rect 1702 2224 1708 2225
rect 1774 2229 1780 2230
rect 1774 2225 1775 2229
rect 1779 2225 1780 2229
rect 1774 2224 1780 2225
rect 1838 2229 1844 2230
rect 1838 2225 1839 2229
rect 1843 2225 1844 2229
rect 1838 2224 1844 2225
rect 1910 2229 1916 2230
rect 1910 2225 1911 2229
rect 1915 2225 1916 2229
rect 1910 2224 1916 2225
rect 1990 2229 1996 2230
rect 1990 2225 1991 2229
rect 1995 2225 1996 2229
rect 1990 2224 1996 2225
rect 2078 2229 2084 2230
rect 2078 2225 2079 2229
rect 2083 2225 2084 2229
rect 2078 2224 2084 2225
rect 2174 2229 2180 2230
rect 2174 2225 2175 2229
rect 2179 2225 2180 2229
rect 2174 2224 2180 2225
rect 2278 2229 2284 2230
rect 2278 2225 2279 2229
rect 2283 2225 2284 2229
rect 2278 2224 2284 2225
rect 2358 2229 2364 2230
rect 2358 2225 2359 2229
rect 2363 2225 2364 2229
rect 2358 2224 2364 2225
rect 142 2217 148 2218
rect 142 2213 143 2217
rect 147 2213 148 2217
rect 142 2212 148 2213
rect 182 2217 188 2218
rect 182 2213 183 2217
rect 187 2213 188 2217
rect 182 2212 188 2213
rect 222 2217 228 2218
rect 222 2213 223 2217
rect 227 2213 228 2217
rect 222 2212 228 2213
rect 278 2217 284 2218
rect 278 2213 279 2217
rect 283 2213 284 2217
rect 278 2212 284 2213
rect 334 2217 340 2218
rect 334 2213 335 2217
rect 339 2213 340 2217
rect 334 2212 340 2213
rect 406 2217 412 2218
rect 406 2213 407 2217
rect 411 2213 412 2217
rect 406 2212 412 2213
rect 478 2217 484 2218
rect 478 2213 479 2217
rect 483 2213 484 2217
rect 478 2212 484 2213
rect 558 2217 564 2218
rect 558 2213 559 2217
rect 563 2213 564 2217
rect 558 2212 564 2213
rect 646 2217 652 2218
rect 646 2213 647 2217
rect 651 2213 652 2217
rect 646 2212 652 2213
rect 726 2217 732 2218
rect 726 2213 727 2217
rect 731 2213 732 2217
rect 726 2212 732 2213
rect 806 2217 812 2218
rect 806 2213 807 2217
rect 811 2213 812 2217
rect 806 2212 812 2213
rect 886 2217 892 2218
rect 886 2213 887 2217
rect 891 2213 892 2217
rect 886 2212 892 2213
rect 966 2217 972 2218
rect 966 2213 967 2217
rect 971 2213 972 2217
rect 966 2212 972 2213
rect 1046 2217 1052 2218
rect 1046 2213 1047 2217
rect 1051 2213 1052 2217
rect 1046 2212 1052 2213
rect 1126 2217 1132 2218
rect 1126 2213 1127 2217
rect 1131 2213 1132 2217
rect 1126 2212 1132 2213
rect 1374 2191 1380 2192
rect 134 2187 140 2188
rect 134 2183 135 2187
rect 139 2183 140 2187
rect 134 2182 140 2183
rect 206 2187 212 2188
rect 206 2183 207 2187
rect 211 2183 212 2187
rect 206 2182 212 2183
rect 278 2187 284 2188
rect 278 2183 279 2187
rect 283 2183 284 2187
rect 278 2182 284 2183
rect 358 2187 364 2188
rect 358 2183 359 2187
rect 363 2183 364 2187
rect 358 2182 364 2183
rect 438 2187 444 2188
rect 438 2183 439 2187
rect 443 2183 444 2187
rect 438 2182 444 2183
rect 518 2187 524 2188
rect 518 2183 519 2187
rect 523 2183 524 2187
rect 518 2182 524 2183
rect 598 2187 604 2188
rect 598 2183 599 2187
rect 603 2183 604 2187
rect 598 2182 604 2183
rect 678 2187 684 2188
rect 678 2183 679 2187
rect 683 2183 684 2187
rect 678 2182 684 2183
rect 758 2187 764 2188
rect 758 2183 759 2187
rect 763 2183 764 2187
rect 758 2182 764 2183
rect 830 2187 836 2188
rect 830 2183 831 2187
rect 835 2183 836 2187
rect 830 2182 836 2183
rect 902 2187 908 2188
rect 902 2183 903 2187
rect 907 2183 908 2187
rect 902 2182 908 2183
rect 974 2187 980 2188
rect 974 2183 975 2187
rect 979 2183 980 2187
rect 974 2182 980 2183
rect 1046 2187 1052 2188
rect 1046 2183 1047 2187
rect 1051 2183 1052 2187
rect 1046 2182 1052 2183
rect 1118 2187 1124 2188
rect 1118 2183 1119 2187
rect 1123 2183 1124 2187
rect 1374 2187 1375 2191
rect 1379 2187 1380 2191
rect 1374 2186 1380 2187
rect 1438 2191 1444 2192
rect 1438 2187 1439 2191
rect 1443 2187 1444 2191
rect 1438 2186 1444 2187
rect 1510 2191 1516 2192
rect 1510 2187 1511 2191
rect 1515 2187 1516 2191
rect 1510 2186 1516 2187
rect 1590 2191 1596 2192
rect 1590 2187 1591 2191
rect 1595 2187 1596 2191
rect 1590 2186 1596 2187
rect 1670 2191 1676 2192
rect 1670 2187 1671 2191
rect 1675 2187 1676 2191
rect 1670 2186 1676 2187
rect 1750 2191 1756 2192
rect 1750 2187 1751 2191
rect 1755 2187 1756 2191
rect 1750 2186 1756 2187
rect 1830 2191 1836 2192
rect 1830 2187 1831 2191
rect 1835 2187 1836 2191
rect 1830 2186 1836 2187
rect 1902 2191 1908 2192
rect 1902 2187 1903 2191
rect 1907 2187 1908 2191
rect 1902 2186 1908 2187
rect 1966 2191 1972 2192
rect 1966 2187 1967 2191
rect 1971 2187 1972 2191
rect 1966 2186 1972 2187
rect 2030 2191 2036 2192
rect 2030 2187 2031 2191
rect 2035 2187 2036 2191
rect 2030 2186 2036 2187
rect 2094 2191 2100 2192
rect 2094 2187 2095 2191
rect 2099 2187 2100 2191
rect 2094 2186 2100 2187
rect 2166 2191 2172 2192
rect 2166 2187 2167 2191
rect 2171 2187 2172 2191
rect 2166 2186 2172 2187
rect 2238 2191 2244 2192
rect 2238 2187 2239 2191
rect 2243 2187 2244 2191
rect 2238 2186 2244 2187
rect 2310 2191 2316 2192
rect 2310 2187 2311 2191
rect 2315 2187 2316 2191
rect 2310 2186 2316 2187
rect 2358 2191 2364 2192
rect 2358 2187 2359 2191
rect 2363 2187 2364 2191
rect 2358 2186 2364 2187
rect 1118 2182 1124 2183
rect 1278 2168 1284 2169
rect 110 2164 116 2165
rect 110 2160 111 2164
rect 115 2160 116 2164
rect 110 2159 116 2160
rect 1238 2164 1244 2165
rect 1238 2160 1239 2164
rect 1243 2160 1244 2164
rect 1278 2164 1279 2168
rect 1283 2164 1284 2168
rect 1278 2163 1284 2164
rect 2406 2168 2412 2169
rect 2406 2164 2407 2168
rect 2411 2164 2412 2168
rect 2406 2163 2412 2164
rect 1238 2159 1244 2160
rect 1278 2151 1284 2152
rect 110 2147 116 2148
rect 110 2143 111 2147
rect 115 2143 116 2147
rect 110 2142 116 2143
rect 1238 2147 1244 2148
rect 1238 2143 1239 2147
rect 1243 2143 1244 2147
rect 1278 2147 1279 2151
rect 1283 2147 1284 2151
rect 1278 2146 1284 2147
rect 2406 2151 2412 2152
rect 2406 2147 2407 2151
rect 2411 2147 2412 2151
rect 2406 2146 2412 2147
rect 1238 2142 1244 2143
rect 1374 2144 1380 2145
rect 134 2140 140 2141
rect 134 2136 135 2140
rect 139 2136 140 2140
rect 134 2135 140 2136
rect 206 2140 212 2141
rect 206 2136 207 2140
rect 211 2136 212 2140
rect 206 2135 212 2136
rect 278 2140 284 2141
rect 278 2136 279 2140
rect 283 2136 284 2140
rect 278 2135 284 2136
rect 358 2140 364 2141
rect 358 2136 359 2140
rect 363 2136 364 2140
rect 358 2135 364 2136
rect 438 2140 444 2141
rect 438 2136 439 2140
rect 443 2136 444 2140
rect 438 2135 444 2136
rect 518 2140 524 2141
rect 518 2136 519 2140
rect 523 2136 524 2140
rect 518 2135 524 2136
rect 598 2140 604 2141
rect 598 2136 599 2140
rect 603 2136 604 2140
rect 598 2135 604 2136
rect 678 2140 684 2141
rect 678 2136 679 2140
rect 683 2136 684 2140
rect 678 2135 684 2136
rect 758 2140 764 2141
rect 758 2136 759 2140
rect 763 2136 764 2140
rect 758 2135 764 2136
rect 830 2140 836 2141
rect 830 2136 831 2140
rect 835 2136 836 2140
rect 830 2135 836 2136
rect 902 2140 908 2141
rect 902 2136 903 2140
rect 907 2136 908 2140
rect 902 2135 908 2136
rect 974 2140 980 2141
rect 974 2136 975 2140
rect 979 2136 980 2140
rect 974 2135 980 2136
rect 1046 2140 1052 2141
rect 1046 2136 1047 2140
rect 1051 2136 1052 2140
rect 1046 2135 1052 2136
rect 1118 2140 1124 2141
rect 1118 2136 1119 2140
rect 1123 2136 1124 2140
rect 1374 2140 1375 2144
rect 1379 2140 1380 2144
rect 1374 2139 1380 2140
rect 1438 2144 1444 2145
rect 1438 2140 1439 2144
rect 1443 2140 1444 2144
rect 1438 2139 1444 2140
rect 1510 2144 1516 2145
rect 1510 2140 1511 2144
rect 1515 2140 1516 2144
rect 1510 2139 1516 2140
rect 1590 2144 1596 2145
rect 1590 2140 1591 2144
rect 1595 2140 1596 2144
rect 1590 2139 1596 2140
rect 1670 2144 1676 2145
rect 1670 2140 1671 2144
rect 1675 2140 1676 2144
rect 1670 2139 1676 2140
rect 1750 2144 1756 2145
rect 1750 2140 1751 2144
rect 1755 2140 1756 2144
rect 1750 2139 1756 2140
rect 1830 2144 1836 2145
rect 1830 2140 1831 2144
rect 1835 2140 1836 2144
rect 1830 2139 1836 2140
rect 1902 2144 1908 2145
rect 1902 2140 1903 2144
rect 1907 2140 1908 2144
rect 1902 2139 1908 2140
rect 1966 2144 1972 2145
rect 1966 2140 1967 2144
rect 1971 2140 1972 2144
rect 1966 2139 1972 2140
rect 2030 2144 2036 2145
rect 2030 2140 2031 2144
rect 2035 2140 2036 2144
rect 2030 2139 2036 2140
rect 2094 2144 2100 2145
rect 2094 2140 2095 2144
rect 2099 2140 2100 2144
rect 2094 2139 2100 2140
rect 2166 2144 2172 2145
rect 2166 2140 2167 2144
rect 2171 2140 2172 2144
rect 2166 2139 2172 2140
rect 2238 2144 2244 2145
rect 2238 2140 2239 2144
rect 2243 2140 2244 2144
rect 2238 2139 2244 2140
rect 2310 2144 2316 2145
rect 2310 2140 2311 2144
rect 2315 2140 2316 2144
rect 2310 2139 2316 2140
rect 2358 2144 2364 2145
rect 2358 2140 2359 2144
rect 2363 2140 2364 2144
rect 2358 2139 2364 2140
rect 1118 2135 1124 2136
rect 1398 2132 1404 2133
rect 1398 2128 1399 2132
rect 1403 2128 1404 2132
rect 1398 2127 1404 2128
rect 1438 2132 1444 2133
rect 1438 2128 1439 2132
rect 1443 2128 1444 2132
rect 1438 2127 1444 2128
rect 1494 2132 1500 2133
rect 1494 2128 1495 2132
rect 1499 2128 1500 2132
rect 1494 2127 1500 2128
rect 1566 2132 1572 2133
rect 1566 2128 1567 2132
rect 1571 2128 1572 2132
rect 1566 2127 1572 2128
rect 1646 2132 1652 2133
rect 1646 2128 1647 2132
rect 1651 2128 1652 2132
rect 1646 2127 1652 2128
rect 1734 2132 1740 2133
rect 1734 2128 1735 2132
rect 1739 2128 1740 2132
rect 1734 2127 1740 2128
rect 1822 2132 1828 2133
rect 1822 2128 1823 2132
rect 1827 2128 1828 2132
rect 1822 2127 1828 2128
rect 1910 2132 1916 2133
rect 1910 2128 1911 2132
rect 1915 2128 1916 2132
rect 1910 2127 1916 2128
rect 1998 2132 2004 2133
rect 1998 2128 1999 2132
rect 2003 2128 2004 2132
rect 1998 2127 2004 2128
rect 2086 2132 2092 2133
rect 2086 2128 2087 2132
rect 2091 2128 2092 2132
rect 2086 2127 2092 2128
rect 2174 2132 2180 2133
rect 2174 2128 2175 2132
rect 2179 2128 2180 2132
rect 2174 2127 2180 2128
rect 2270 2132 2276 2133
rect 2270 2128 2271 2132
rect 2275 2128 2276 2132
rect 2270 2127 2276 2128
rect 2358 2132 2364 2133
rect 2358 2128 2359 2132
rect 2363 2128 2364 2132
rect 2358 2127 2364 2128
rect 1278 2125 1284 2126
rect 1278 2121 1279 2125
rect 1283 2121 1284 2125
rect 134 2120 140 2121
rect 134 2116 135 2120
rect 139 2116 140 2120
rect 134 2115 140 2116
rect 190 2120 196 2121
rect 190 2116 191 2120
rect 195 2116 196 2120
rect 190 2115 196 2116
rect 270 2120 276 2121
rect 270 2116 271 2120
rect 275 2116 276 2120
rect 270 2115 276 2116
rect 342 2120 348 2121
rect 342 2116 343 2120
rect 347 2116 348 2120
rect 342 2115 348 2116
rect 414 2120 420 2121
rect 414 2116 415 2120
rect 419 2116 420 2120
rect 414 2115 420 2116
rect 478 2120 484 2121
rect 478 2116 479 2120
rect 483 2116 484 2120
rect 478 2115 484 2116
rect 542 2120 548 2121
rect 542 2116 543 2120
rect 547 2116 548 2120
rect 542 2115 548 2116
rect 606 2120 612 2121
rect 606 2116 607 2120
rect 611 2116 612 2120
rect 606 2115 612 2116
rect 670 2120 676 2121
rect 670 2116 671 2120
rect 675 2116 676 2120
rect 670 2115 676 2116
rect 734 2120 740 2121
rect 734 2116 735 2120
rect 739 2116 740 2120
rect 734 2115 740 2116
rect 790 2120 796 2121
rect 790 2116 791 2120
rect 795 2116 796 2120
rect 790 2115 796 2116
rect 838 2120 844 2121
rect 838 2116 839 2120
rect 843 2116 844 2120
rect 838 2115 844 2116
rect 886 2120 892 2121
rect 886 2116 887 2120
rect 891 2116 892 2120
rect 886 2115 892 2116
rect 934 2120 940 2121
rect 934 2116 935 2120
rect 939 2116 940 2120
rect 934 2115 940 2116
rect 990 2120 996 2121
rect 990 2116 991 2120
rect 995 2116 996 2120
rect 990 2115 996 2116
rect 1046 2120 1052 2121
rect 1278 2120 1284 2121
rect 2406 2125 2412 2126
rect 2406 2121 2407 2125
rect 2411 2121 2412 2125
rect 2406 2120 2412 2121
rect 1046 2116 1047 2120
rect 1051 2116 1052 2120
rect 1046 2115 1052 2116
rect 110 2113 116 2114
rect 110 2109 111 2113
rect 115 2109 116 2113
rect 110 2108 116 2109
rect 1238 2113 1244 2114
rect 1238 2109 1239 2113
rect 1243 2109 1244 2113
rect 1238 2108 1244 2109
rect 1278 2108 1284 2109
rect 1278 2104 1279 2108
rect 1283 2104 1284 2108
rect 1278 2103 1284 2104
rect 2406 2108 2412 2109
rect 2406 2104 2407 2108
rect 2411 2104 2412 2108
rect 2406 2103 2412 2104
rect 110 2096 116 2097
rect 110 2092 111 2096
rect 115 2092 116 2096
rect 110 2091 116 2092
rect 1238 2096 1244 2097
rect 1238 2092 1239 2096
rect 1243 2092 1244 2096
rect 1238 2091 1244 2092
rect 1398 2085 1404 2086
rect 1398 2081 1399 2085
rect 1403 2081 1404 2085
rect 1398 2080 1404 2081
rect 1438 2085 1444 2086
rect 1438 2081 1439 2085
rect 1443 2081 1444 2085
rect 1438 2080 1444 2081
rect 1494 2085 1500 2086
rect 1494 2081 1495 2085
rect 1499 2081 1500 2085
rect 1494 2080 1500 2081
rect 1566 2085 1572 2086
rect 1566 2081 1567 2085
rect 1571 2081 1572 2085
rect 1566 2080 1572 2081
rect 1646 2085 1652 2086
rect 1646 2081 1647 2085
rect 1651 2081 1652 2085
rect 1646 2080 1652 2081
rect 1734 2085 1740 2086
rect 1734 2081 1735 2085
rect 1739 2081 1740 2085
rect 1734 2080 1740 2081
rect 1822 2085 1828 2086
rect 1822 2081 1823 2085
rect 1827 2081 1828 2085
rect 1822 2080 1828 2081
rect 1910 2085 1916 2086
rect 1910 2081 1911 2085
rect 1915 2081 1916 2085
rect 1910 2080 1916 2081
rect 1998 2085 2004 2086
rect 1998 2081 1999 2085
rect 2003 2081 2004 2085
rect 1998 2080 2004 2081
rect 2086 2085 2092 2086
rect 2086 2081 2087 2085
rect 2091 2081 2092 2085
rect 2086 2080 2092 2081
rect 2174 2085 2180 2086
rect 2174 2081 2175 2085
rect 2179 2081 2180 2085
rect 2174 2080 2180 2081
rect 2270 2085 2276 2086
rect 2270 2081 2271 2085
rect 2275 2081 2276 2085
rect 2270 2080 2276 2081
rect 2358 2085 2364 2086
rect 2358 2081 2359 2085
rect 2363 2081 2364 2085
rect 2358 2080 2364 2081
rect 134 2073 140 2074
rect 134 2069 135 2073
rect 139 2069 140 2073
rect 134 2068 140 2069
rect 190 2073 196 2074
rect 190 2069 191 2073
rect 195 2069 196 2073
rect 190 2068 196 2069
rect 270 2073 276 2074
rect 270 2069 271 2073
rect 275 2069 276 2073
rect 270 2068 276 2069
rect 342 2073 348 2074
rect 342 2069 343 2073
rect 347 2069 348 2073
rect 342 2068 348 2069
rect 414 2073 420 2074
rect 414 2069 415 2073
rect 419 2069 420 2073
rect 414 2068 420 2069
rect 478 2073 484 2074
rect 478 2069 479 2073
rect 483 2069 484 2073
rect 478 2068 484 2069
rect 542 2073 548 2074
rect 542 2069 543 2073
rect 547 2069 548 2073
rect 542 2068 548 2069
rect 606 2073 612 2074
rect 606 2069 607 2073
rect 611 2069 612 2073
rect 606 2068 612 2069
rect 670 2073 676 2074
rect 670 2069 671 2073
rect 675 2069 676 2073
rect 670 2068 676 2069
rect 734 2073 740 2074
rect 734 2069 735 2073
rect 739 2069 740 2073
rect 734 2068 740 2069
rect 790 2073 796 2074
rect 790 2069 791 2073
rect 795 2069 796 2073
rect 790 2068 796 2069
rect 838 2073 844 2074
rect 838 2069 839 2073
rect 843 2069 844 2073
rect 838 2068 844 2069
rect 886 2073 892 2074
rect 886 2069 887 2073
rect 891 2069 892 2073
rect 886 2068 892 2069
rect 934 2073 940 2074
rect 934 2069 935 2073
rect 939 2069 940 2073
rect 934 2068 940 2069
rect 990 2073 996 2074
rect 990 2069 991 2073
rect 995 2069 996 2073
rect 990 2068 996 2069
rect 1046 2073 1052 2074
rect 1046 2069 1047 2073
rect 1051 2069 1052 2073
rect 1046 2068 1052 2069
rect 2038 2055 2044 2056
rect 2038 2051 2039 2055
rect 2043 2051 2044 2055
rect 2038 2050 2044 2051
rect 2078 2055 2084 2056
rect 2078 2051 2079 2055
rect 2083 2051 2084 2055
rect 2078 2050 2084 2051
rect 2118 2055 2124 2056
rect 2118 2051 2119 2055
rect 2123 2051 2124 2055
rect 2118 2050 2124 2051
rect 2158 2055 2164 2056
rect 2158 2051 2159 2055
rect 2163 2051 2164 2055
rect 2158 2050 2164 2051
rect 2198 2055 2204 2056
rect 2198 2051 2199 2055
rect 2203 2051 2204 2055
rect 2198 2050 2204 2051
rect 2238 2055 2244 2056
rect 2238 2051 2239 2055
rect 2243 2051 2244 2055
rect 2238 2050 2244 2051
rect 2278 2055 2284 2056
rect 2278 2051 2279 2055
rect 2283 2051 2284 2055
rect 2278 2050 2284 2051
rect 2318 2055 2324 2056
rect 2318 2051 2319 2055
rect 2323 2051 2324 2055
rect 2318 2050 2324 2051
rect 2358 2055 2364 2056
rect 2358 2051 2359 2055
rect 2363 2051 2364 2055
rect 2358 2050 2364 2051
rect 134 2039 140 2040
rect 134 2035 135 2039
rect 139 2035 140 2039
rect 134 2034 140 2035
rect 174 2039 180 2040
rect 174 2035 175 2039
rect 179 2035 180 2039
rect 174 2034 180 2035
rect 214 2039 220 2040
rect 214 2035 215 2039
rect 219 2035 220 2039
rect 214 2034 220 2035
rect 278 2039 284 2040
rect 278 2035 279 2039
rect 283 2035 284 2039
rect 278 2034 284 2035
rect 350 2039 356 2040
rect 350 2035 351 2039
rect 355 2035 356 2039
rect 350 2034 356 2035
rect 422 2039 428 2040
rect 422 2035 423 2039
rect 427 2035 428 2039
rect 422 2034 428 2035
rect 486 2039 492 2040
rect 486 2035 487 2039
rect 491 2035 492 2039
rect 486 2034 492 2035
rect 550 2039 556 2040
rect 550 2035 551 2039
rect 555 2035 556 2039
rect 550 2034 556 2035
rect 614 2039 620 2040
rect 614 2035 615 2039
rect 619 2035 620 2039
rect 614 2034 620 2035
rect 678 2039 684 2040
rect 678 2035 679 2039
rect 683 2035 684 2039
rect 678 2034 684 2035
rect 742 2039 748 2040
rect 742 2035 743 2039
rect 747 2035 748 2039
rect 742 2034 748 2035
rect 814 2039 820 2040
rect 814 2035 815 2039
rect 819 2035 820 2039
rect 814 2034 820 2035
rect 1278 2032 1284 2033
rect 1278 2028 1279 2032
rect 1283 2028 1284 2032
rect 1278 2027 1284 2028
rect 2406 2032 2412 2033
rect 2406 2028 2407 2032
rect 2411 2028 2412 2032
rect 2406 2027 2412 2028
rect 110 2016 116 2017
rect 110 2012 111 2016
rect 115 2012 116 2016
rect 110 2011 116 2012
rect 1238 2016 1244 2017
rect 1238 2012 1239 2016
rect 1243 2012 1244 2016
rect 1238 2011 1244 2012
rect 1278 2015 1284 2016
rect 1278 2011 1279 2015
rect 1283 2011 1284 2015
rect 1278 2010 1284 2011
rect 2406 2015 2412 2016
rect 2406 2011 2407 2015
rect 2411 2011 2412 2015
rect 2406 2010 2412 2011
rect 2038 2008 2044 2009
rect 2038 2004 2039 2008
rect 2043 2004 2044 2008
rect 2038 2003 2044 2004
rect 2078 2008 2084 2009
rect 2078 2004 2079 2008
rect 2083 2004 2084 2008
rect 2078 2003 2084 2004
rect 2118 2008 2124 2009
rect 2118 2004 2119 2008
rect 2123 2004 2124 2008
rect 2118 2003 2124 2004
rect 2158 2008 2164 2009
rect 2158 2004 2159 2008
rect 2163 2004 2164 2008
rect 2158 2003 2164 2004
rect 2198 2008 2204 2009
rect 2198 2004 2199 2008
rect 2203 2004 2204 2008
rect 2198 2003 2204 2004
rect 2238 2008 2244 2009
rect 2238 2004 2239 2008
rect 2243 2004 2244 2008
rect 2238 2003 2244 2004
rect 2278 2008 2284 2009
rect 2278 2004 2279 2008
rect 2283 2004 2284 2008
rect 2278 2003 2284 2004
rect 2318 2008 2324 2009
rect 2318 2004 2319 2008
rect 2323 2004 2324 2008
rect 2318 2003 2324 2004
rect 2358 2008 2364 2009
rect 2358 2004 2359 2008
rect 2363 2004 2364 2008
rect 2358 2003 2364 2004
rect 110 1999 116 2000
rect 110 1995 111 1999
rect 115 1995 116 1999
rect 110 1994 116 1995
rect 1238 1999 1244 2000
rect 1238 1995 1239 1999
rect 1243 1995 1244 1999
rect 1238 1994 1244 1995
rect 1398 1996 1404 1997
rect 134 1992 140 1993
rect 134 1988 135 1992
rect 139 1988 140 1992
rect 134 1987 140 1988
rect 174 1992 180 1993
rect 174 1988 175 1992
rect 179 1988 180 1992
rect 174 1987 180 1988
rect 214 1992 220 1993
rect 214 1988 215 1992
rect 219 1988 220 1992
rect 214 1987 220 1988
rect 278 1992 284 1993
rect 278 1988 279 1992
rect 283 1988 284 1992
rect 278 1987 284 1988
rect 350 1992 356 1993
rect 350 1988 351 1992
rect 355 1988 356 1992
rect 350 1987 356 1988
rect 422 1992 428 1993
rect 422 1988 423 1992
rect 427 1988 428 1992
rect 422 1987 428 1988
rect 486 1992 492 1993
rect 486 1988 487 1992
rect 491 1988 492 1992
rect 486 1987 492 1988
rect 550 1992 556 1993
rect 550 1988 551 1992
rect 555 1988 556 1992
rect 550 1987 556 1988
rect 614 1992 620 1993
rect 614 1988 615 1992
rect 619 1988 620 1992
rect 614 1987 620 1988
rect 678 1992 684 1993
rect 678 1988 679 1992
rect 683 1988 684 1992
rect 678 1987 684 1988
rect 742 1992 748 1993
rect 742 1988 743 1992
rect 747 1988 748 1992
rect 742 1987 748 1988
rect 814 1992 820 1993
rect 814 1988 815 1992
rect 819 1988 820 1992
rect 1398 1992 1399 1996
rect 1403 1992 1404 1996
rect 1398 1991 1404 1992
rect 1438 1996 1444 1997
rect 1438 1992 1439 1996
rect 1443 1992 1444 1996
rect 1438 1991 1444 1992
rect 1478 1996 1484 1997
rect 1478 1992 1479 1996
rect 1483 1992 1484 1996
rect 1478 1991 1484 1992
rect 1518 1996 1524 1997
rect 1518 1992 1519 1996
rect 1523 1992 1524 1996
rect 1518 1991 1524 1992
rect 1558 1996 1564 1997
rect 1558 1992 1559 1996
rect 1563 1992 1564 1996
rect 1558 1991 1564 1992
rect 1598 1996 1604 1997
rect 1598 1992 1599 1996
rect 1603 1992 1604 1996
rect 1598 1991 1604 1992
rect 1638 1996 1644 1997
rect 1638 1992 1639 1996
rect 1643 1992 1644 1996
rect 1638 1991 1644 1992
rect 1678 1996 1684 1997
rect 1678 1992 1679 1996
rect 1683 1992 1684 1996
rect 1678 1991 1684 1992
rect 1718 1996 1724 1997
rect 1718 1992 1719 1996
rect 1723 1992 1724 1996
rect 1718 1991 1724 1992
rect 1766 1996 1772 1997
rect 1766 1992 1767 1996
rect 1771 1992 1772 1996
rect 1766 1991 1772 1992
rect 1822 1996 1828 1997
rect 1822 1992 1823 1996
rect 1827 1992 1828 1996
rect 1822 1991 1828 1992
rect 1870 1996 1876 1997
rect 1870 1992 1871 1996
rect 1875 1992 1876 1996
rect 1870 1991 1876 1992
rect 1918 1996 1924 1997
rect 1918 1992 1919 1996
rect 1923 1992 1924 1996
rect 1918 1991 1924 1992
rect 1966 1996 1972 1997
rect 1966 1992 1967 1996
rect 1971 1992 1972 1996
rect 1966 1991 1972 1992
rect 2014 1996 2020 1997
rect 2014 1992 2015 1996
rect 2019 1992 2020 1996
rect 2014 1991 2020 1992
rect 2054 1996 2060 1997
rect 2054 1992 2055 1996
rect 2059 1992 2060 1996
rect 2054 1991 2060 1992
rect 2094 1996 2100 1997
rect 2094 1992 2095 1996
rect 2099 1992 2100 1996
rect 2094 1991 2100 1992
rect 2142 1996 2148 1997
rect 2142 1992 2143 1996
rect 2147 1992 2148 1996
rect 2142 1991 2148 1992
rect 2190 1996 2196 1997
rect 2190 1992 2191 1996
rect 2195 1992 2196 1996
rect 2190 1991 2196 1992
rect 2238 1996 2244 1997
rect 2238 1992 2239 1996
rect 2243 1992 2244 1996
rect 2238 1991 2244 1992
rect 2278 1996 2284 1997
rect 2278 1992 2279 1996
rect 2283 1992 2284 1996
rect 2278 1991 2284 1992
rect 2318 1996 2324 1997
rect 2318 1992 2319 1996
rect 2323 1992 2324 1996
rect 2318 1991 2324 1992
rect 2358 1996 2364 1997
rect 2358 1992 2359 1996
rect 2363 1992 2364 1996
rect 2358 1991 2364 1992
rect 814 1987 820 1988
rect 1278 1989 1284 1990
rect 1278 1985 1279 1989
rect 1283 1985 1284 1989
rect 1278 1984 1284 1985
rect 2406 1989 2412 1990
rect 2406 1985 2407 1989
rect 2411 1985 2412 1989
rect 2406 1984 2412 1985
rect 134 1980 140 1981
rect 134 1976 135 1980
rect 139 1976 140 1980
rect 134 1975 140 1976
rect 174 1980 180 1981
rect 174 1976 175 1980
rect 179 1976 180 1980
rect 174 1975 180 1976
rect 214 1980 220 1981
rect 214 1976 215 1980
rect 219 1976 220 1980
rect 214 1975 220 1976
rect 270 1980 276 1981
rect 270 1976 271 1980
rect 275 1976 276 1980
rect 270 1975 276 1976
rect 342 1980 348 1981
rect 342 1976 343 1980
rect 347 1976 348 1980
rect 342 1975 348 1976
rect 414 1980 420 1981
rect 414 1976 415 1980
rect 419 1976 420 1980
rect 414 1975 420 1976
rect 494 1980 500 1981
rect 494 1976 495 1980
rect 499 1976 500 1980
rect 494 1975 500 1976
rect 574 1980 580 1981
rect 574 1976 575 1980
rect 579 1976 580 1980
rect 574 1975 580 1976
rect 646 1980 652 1981
rect 646 1976 647 1980
rect 651 1976 652 1980
rect 646 1975 652 1976
rect 718 1980 724 1981
rect 718 1976 719 1980
rect 723 1976 724 1980
rect 718 1975 724 1976
rect 790 1980 796 1981
rect 790 1976 791 1980
rect 795 1976 796 1980
rect 790 1975 796 1976
rect 862 1980 868 1981
rect 862 1976 863 1980
rect 867 1976 868 1980
rect 862 1975 868 1976
rect 934 1980 940 1981
rect 934 1976 935 1980
rect 939 1976 940 1980
rect 934 1975 940 1976
rect 1006 1980 1012 1981
rect 1006 1976 1007 1980
rect 1011 1976 1012 1980
rect 1006 1975 1012 1976
rect 110 1973 116 1974
rect 110 1969 111 1973
rect 115 1969 116 1973
rect 110 1968 116 1969
rect 1238 1973 1244 1974
rect 1238 1969 1239 1973
rect 1243 1969 1244 1973
rect 1238 1968 1244 1969
rect 1278 1972 1284 1973
rect 1278 1968 1279 1972
rect 1283 1968 1284 1972
rect 1278 1967 1284 1968
rect 2406 1972 2412 1973
rect 2406 1968 2407 1972
rect 2411 1968 2412 1972
rect 2406 1967 2412 1968
rect 110 1956 116 1957
rect 110 1952 111 1956
rect 115 1952 116 1956
rect 110 1951 116 1952
rect 1238 1956 1244 1957
rect 1238 1952 1239 1956
rect 1243 1952 1244 1956
rect 1238 1951 1244 1952
rect 1398 1949 1404 1950
rect 1398 1945 1399 1949
rect 1403 1945 1404 1949
rect 1398 1944 1404 1945
rect 1438 1949 1444 1950
rect 1438 1945 1439 1949
rect 1443 1945 1444 1949
rect 1438 1944 1444 1945
rect 1478 1949 1484 1950
rect 1478 1945 1479 1949
rect 1483 1945 1484 1949
rect 1478 1944 1484 1945
rect 1518 1949 1524 1950
rect 1518 1945 1519 1949
rect 1523 1945 1524 1949
rect 1518 1944 1524 1945
rect 1558 1949 1564 1950
rect 1558 1945 1559 1949
rect 1563 1945 1564 1949
rect 1558 1944 1564 1945
rect 1598 1949 1604 1950
rect 1598 1945 1599 1949
rect 1603 1945 1604 1949
rect 1598 1944 1604 1945
rect 1638 1949 1644 1950
rect 1638 1945 1639 1949
rect 1643 1945 1644 1949
rect 1638 1944 1644 1945
rect 1678 1949 1684 1950
rect 1678 1945 1679 1949
rect 1683 1945 1684 1949
rect 1678 1944 1684 1945
rect 1718 1949 1724 1950
rect 1718 1945 1719 1949
rect 1723 1945 1724 1949
rect 1718 1944 1724 1945
rect 1766 1949 1772 1950
rect 1766 1945 1767 1949
rect 1771 1945 1772 1949
rect 1766 1944 1772 1945
rect 1822 1949 1828 1950
rect 1822 1945 1823 1949
rect 1827 1945 1828 1949
rect 1822 1944 1828 1945
rect 1870 1949 1876 1950
rect 1870 1945 1871 1949
rect 1875 1945 1876 1949
rect 1870 1944 1876 1945
rect 1918 1949 1924 1950
rect 1918 1945 1919 1949
rect 1923 1945 1924 1949
rect 1918 1944 1924 1945
rect 1966 1949 1972 1950
rect 1966 1945 1967 1949
rect 1971 1945 1972 1949
rect 1966 1944 1972 1945
rect 2014 1949 2020 1950
rect 2014 1945 2015 1949
rect 2019 1945 2020 1949
rect 2014 1944 2020 1945
rect 2054 1949 2060 1950
rect 2054 1945 2055 1949
rect 2059 1945 2060 1949
rect 2054 1944 2060 1945
rect 2094 1949 2100 1950
rect 2094 1945 2095 1949
rect 2099 1945 2100 1949
rect 2094 1944 2100 1945
rect 2142 1949 2148 1950
rect 2142 1945 2143 1949
rect 2147 1945 2148 1949
rect 2142 1944 2148 1945
rect 2190 1949 2196 1950
rect 2190 1945 2191 1949
rect 2195 1945 2196 1949
rect 2190 1944 2196 1945
rect 2238 1949 2244 1950
rect 2238 1945 2239 1949
rect 2243 1945 2244 1949
rect 2238 1944 2244 1945
rect 2278 1949 2284 1950
rect 2278 1945 2279 1949
rect 2283 1945 2284 1949
rect 2278 1944 2284 1945
rect 2318 1949 2324 1950
rect 2318 1945 2319 1949
rect 2323 1945 2324 1949
rect 2318 1944 2324 1945
rect 2358 1949 2364 1950
rect 2358 1945 2359 1949
rect 2363 1945 2364 1949
rect 2358 1944 2364 1945
rect 134 1933 140 1934
rect 134 1929 135 1933
rect 139 1929 140 1933
rect 134 1928 140 1929
rect 174 1933 180 1934
rect 174 1929 175 1933
rect 179 1929 180 1933
rect 174 1928 180 1929
rect 214 1933 220 1934
rect 214 1929 215 1933
rect 219 1929 220 1933
rect 214 1928 220 1929
rect 270 1933 276 1934
rect 270 1929 271 1933
rect 275 1929 276 1933
rect 270 1928 276 1929
rect 342 1933 348 1934
rect 342 1929 343 1933
rect 347 1929 348 1933
rect 342 1928 348 1929
rect 414 1933 420 1934
rect 414 1929 415 1933
rect 419 1929 420 1933
rect 414 1928 420 1929
rect 494 1933 500 1934
rect 494 1929 495 1933
rect 499 1929 500 1933
rect 494 1928 500 1929
rect 574 1933 580 1934
rect 574 1929 575 1933
rect 579 1929 580 1933
rect 574 1928 580 1929
rect 646 1933 652 1934
rect 646 1929 647 1933
rect 651 1929 652 1933
rect 646 1928 652 1929
rect 718 1933 724 1934
rect 718 1929 719 1933
rect 723 1929 724 1933
rect 718 1928 724 1929
rect 790 1933 796 1934
rect 790 1929 791 1933
rect 795 1929 796 1933
rect 790 1928 796 1929
rect 862 1933 868 1934
rect 862 1929 863 1933
rect 867 1929 868 1933
rect 862 1928 868 1929
rect 934 1933 940 1934
rect 934 1929 935 1933
rect 939 1929 940 1933
rect 934 1928 940 1929
rect 1006 1933 1012 1934
rect 1006 1929 1007 1933
rect 1011 1929 1012 1933
rect 1006 1928 1012 1929
rect 1342 1915 1348 1916
rect 1342 1911 1343 1915
rect 1347 1911 1348 1915
rect 1342 1910 1348 1911
rect 1382 1915 1388 1916
rect 1382 1911 1383 1915
rect 1387 1911 1388 1915
rect 1382 1910 1388 1911
rect 1422 1915 1428 1916
rect 1422 1911 1423 1915
rect 1427 1911 1428 1915
rect 1422 1910 1428 1911
rect 1462 1915 1468 1916
rect 1462 1911 1463 1915
rect 1467 1911 1468 1915
rect 1462 1910 1468 1911
rect 1510 1915 1516 1916
rect 1510 1911 1511 1915
rect 1515 1911 1516 1915
rect 1510 1910 1516 1911
rect 1566 1915 1572 1916
rect 1566 1911 1567 1915
rect 1571 1911 1572 1915
rect 1566 1910 1572 1911
rect 1630 1915 1636 1916
rect 1630 1911 1631 1915
rect 1635 1911 1636 1915
rect 1630 1910 1636 1911
rect 1710 1915 1716 1916
rect 1710 1911 1711 1915
rect 1715 1911 1716 1915
rect 1710 1910 1716 1911
rect 1806 1915 1812 1916
rect 1806 1911 1807 1915
rect 1811 1911 1812 1915
rect 1806 1910 1812 1911
rect 1918 1915 1924 1916
rect 1918 1911 1919 1915
rect 1923 1911 1924 1915
rect 1918 1910 1924 1911
rect 2030 1915 2036 1916
rect 2030 1911 2031 1915
rect 2035 1911 2036 1915
rect 2030 1910 2036 1911
rect 2150 1915 2156 1916
rect 2150 1911 2151 1915
rect 2155 1911 2156 1915
rect 2150 1910 2156 1911
rect 246 1899 252 1900
rect 246 1895 247 1899
rect 251 1895 252 1899
rect 246 1894 252 1895
rect 286 1899 292 1900
rect 286 1895 287 1899
rect 291 1895 292 1899
rect 286 1894 292 1895
rect 326 1899 332 1900
rect 326 1895 327 1899
rect 331 1895 332 1899
rect 326 1894 332 1895
rect 366 1899 372 1900
rect 366 1895 367 1899
rect 371 1895 372 1899
rect 366 1894 372 1895
rect 414 1899 420 1900
rect 414 1895 415 1899
rect 419 1895 420 1899
rect 414 1894 420 1895
rect 470 1899 476 1900
rect 470 1895 471 1899
rect 475 1895 476 1899
rect 470 1894 476 1895
rect 534 1899 540 1900
rect 534 1895 535 1899
rect 539 1895 540 1899
rect 534 1894 540 1895
rect 598 1899 604 1900
rect 598 1895 599 1899
rect 603 1895 604 1899
rect 598 1894 604 1895
rect 662 1899 668 1900
rect 662 1895 663 1899
rect 667 1895 668 1899
rect 662 1894 668 1895
rect 726 1899 732 1900
rect 726 1895 727 1899
rect 731 1895 732 1899
rect 726 1894 732 1895
rect 790 1899 796 1900
rect 790 1895 791 1899
rect 795 1895 796 1899
rect 790 1894 796 1895
rect 854 1899 860 1900
rect 854 1895 855 1899
rect 859 1895 860 1899
rect 854 1894 860 1895
rect 918 1899 924 1900
rect 918 1895 919 1899
rect 923 1895 924 1899
rect 918 1894 924 1895
rect 982 1899 988 1900
rect 982 1895 983 1899
rect 987 1895 988 1899
rect 982 1894 988 1895
rect 1054 1899 1060 1900
rect 1054 1895 1055 1899
rect 1059 1895 1060 1899
rect 1054 1894 1060 1895
rect 1126 1899 1132 1900
rect 1126 1895 1127 1899
rect 1131 1895 1132 1899
rect 1126 1894 1132 1895
rect 1278 1892 1284 1893
rect 1278 1888 1279 1892
rect 1283 1888 1284 1892
rect 1278 1887 1284 1888
rect 2406 1892 2412 1893
rect 2406 1888 2407 1892
rect 2411 1888 2412 1892
rect 2406 1887 2412 1888
rect 110 1876 116 1877
rect 110 1872 111 1876
rect 115 1872 116 1876
rect 110 1871 116 1872
rect 1238 1876 1244 1877
rect 1238 1872 1239 1876
rect 1243 1872 1244 1876
rect 1238 1871 1244 1872
rect 1278 1875 1284 1876
rect 1278 1871 1279 1875
rect 1283 1871 1284 1875
rect 1278 1870 1284 1871
rect 2406 1875 2412 1876
rect 2406 1871 2407 1875
rect 2411 1871 2412 1875
rect 2406 1870 2412 1871
rect 1342 1868 1348 1869
rect 1342 1864 1343 1868
rect 1347 1864 1348 1868
rect 1342 1863 1348 1864
rect 1382 1868 1388 1869
rect 1382 1864 1383 1868
rect 1387 1864 1388 1868
rect 1382 1863 1388 1864
rect 1422 1868 1428 1869
rect 1422 1864 1423 1868
rect 1427 1864 1428 1868
rect 1422 1863 1428 1864
rect 1462 1868 1468 1869
rect 1462 1864 1463 1868
rect 1467 1864 1468 1868
rect 1462 1863 1468 1864
rect 1510 1868 1516 1869
rect 1510 1864 1511 1868
rect 1515 1864 1516 1868
rect 1510 1863 1516 1864
rect 1566 1868 1572 1869
rect 1566 1864 1567 1868
rect 1571 1864 1572 1868
rect 1566 1863 1572 1864
rect 1630 1868 1636 1869
rect 1630 1864 1631 1868
rect 1635 1864 1636 1868
rect 1630 1863 1636 1864
rect 1710 1868 1716 1869
rect 1710 1864 1711 1868
rect 1715 1864 1716 1868
rect 1710 1863 1716 1864
rect 1806 1868 1812 1869
rect 1806 1864 1807 1868
rect 1811 1864 1812 1868
rect 1806 1863 1812 1864
rect 1918 1868 1924 1869
rect 1918 1864 1919 1868
rect 1923 1864 1924 1868
rect 1918 1863 1924 1864
rect 2030 1868 2036 1869
rect 2030 1864 2031 1868
rect 2035 1864 2036 1868
rect 2030 1863 2036 1864
rect 2150 1868 2156 1869
rect 2150 1864 2151 1868
rect 2155 1864 2156 1868
rect 2150 1863 2156 1864
rect 110 1859 116 1860
rect 110 1855 111 1859
rect 115 1855 116 1859
rect 110 1854 116 1855
rect 1238 1859 1244 1860
rect 1238 1855 1239 1859
rect 1243 1855 1244 1859
rect 1238 1854 1244 1855
rect 246 1852 252 1853
rect 246 1848 247 1852
rect 251 1848 252 1852
rect 246 1847 252 1848
rect 286 1852 292 1853
rect 286 1848 287 1852
rect 291 1848 292 1852
rect 286 1847 292 1848
rect 326 1852 332 1853
rect 326 1848 327 1852
rect 331 1848 332 1852
rect 326 1847 332 1848
rect 366 1852 372 1853
rect 366 1848 367 1852
rect 371 1848 372 1852
rect 366 1847 372 1848
rect 414 1852 420 1853
rect 414 1848 415 1852
rect 419 1848 420 1852
rect 414 1847 420 1848
rect 470 1852 476 1853
rect 470 1848 471 1852
rect 475 1848 476 1852
rect 470 1847 476 1848
rect 534 1852 540 1853
rect 534 1848 535 1852
rect 539 1848 540 1852
rect 534 1847 540 1848
rect 598 1852 604 1853
rect 598 1848 599 1852
rect 603 1848 604 1852
rect 598 1847 604 1848
rect 662 1852 668 1853
rect 662 1848 663 1852
rect 667 1848 668 1852
rect 662 1847 668 1848
rect 726 1852 732 1853
rect 726 1848 727 1852
rect 731 1848 732 1852
rect 726 1847 732 1848
rect 790 1852 796 1853
rect 790 1848 791 1852
rect 795 1848 796 1852
rect 790 1847 796 1848
rect 854 1852 860 1853
rect 854 1848 855 1852
rect 859 1848 860 1852
rect 854 1847 860 1848
rect 918 1852 924 1853
rect 918 1848 919 1852
rect 923 1848 924 1852
rect 918 1847 924 1848
rect 982 1852 988 1853
rect 982 1848 983 1852
rect 987 1848 988 1852
rect 982 1847 988 1848
rect 1054 1852 1060 1853
rect 1054 1848 1055 1852
rect 1059 1848 1060 1852
rect 1054 1847 1060 1848
rect 1126 1852 1132 1853
rect 1126 1848 1127 1852
rect 1131 1848 1132 1852
rect 1126 1847 1132 1848
rect 1358 1848 1364 1849
rect 1358 1844 1359 1848
rect 1363 1844 1364 1848
rect 1358 1843 1364 1844
rect 1398 1848 1404 1849
rect 1398 1844 1399 1848
rect 1403 1844 1404 1848
rect 1398 1843 1404 1844
rect 1446 1848 1452 1849
rect 1446 1844 1447 1848
rect 1451 1844 1452 1848
rect 1446 1843 1452 1844
rect 1502 1848 1508 1849
rect 1502 1844 1503 1848
rect 1507 1844 1508 1848
rect 1502 1843 1508 1844
rect 1558 1848 1564 1849
rect 1558 1844 1559 1848
rect 1563 1844 1564 1848
rect 1558 1843 1564 1844
rect 1614 1848 1620 1849
rect 1614 1844 1615 1848
rect 1619 1844 1620 1848
rect 1614 1843 1620 1844
rect 1670 1848 1676 1849
rect 1670 1844 1671 1848
rect 1675 1844 1676 1848
rect 1670 1843 1676 1844
rect 1726 1848 1732 1849
rect 1726 1844 1727 1848
rect 1731 1844 1732 1848
rect 1726 1843 1732 1844
rect 1782 1848 1788 1849
rect 1782 1844 1783 1848
rect 1787 1844 1788 1848
rect 1782 1843 1788 1844
rect 1838 1848 1844 1849
rect 1838 1844 1839 1848
rect 1843 1844 1844 1848
rect 1838 1843 1844 1844
rect 1894 1848 1900 1849
rect 1894 1844 1895 1848
rect 1899 1844 1900 1848
rect 1894 1843 1900 1844
rect 1950 1848 1956 1849
rect 1950 1844 1951 1848
rect 1955 1844 1956 1848
rect 1950 1843 1956 1844
rect 1278 1841 1284 1842
rect 1278 1837 1279 1841
rect 1283 1837 1284 1841
rect 398 1836 404 1837
rect 398 1832 399 1836
rect 403 1832 404 1836
rect 398 1831 404 1832
rect 438 1836 444 1837
rect 438 1832 439 1836
rect 443 1832 444 1836
rect 438 1831 444 1832
rect 478 1836 484 1837
rect 478 1832 479 1836
rect 483 1832 484 1836
rect 478 1831 484 1832
rect 518 1836 524 1837
rect 518 1832 519 1836
rect 523 1832 524 1836
rect 518 1831 524 1832
rect 566 1836 572 1837
rect 566 1832 567 1836
rect 571 1832 572 1836
rect 566 1831 572 1832
rect 622 1836 628 1837
rect 622 1832 623 1836
rect 627 1832 628 1836
rect 622 1831 628 1832
rect 686 1836 692 1837
rect 686 1832 687 1836
rect 691 1832 692 1836
rect 686 1831 692 1832
rect 758 1836 764 1837
rect 758 1832 759 1836
rect 763 1832 764 1836
rect 758 1831 764 1832
rect 830 1836 836 1837
rect 830 1832 831 1836
rect 835 1832 836 1836
rect 830 1831 836 1832
rect 902 1836 908 1837
rect 902 1832 903 1836
rect 907 1832 908 1836
rect 902 1831 908 1832
rect 974 1836 980 1837
rect 974 1832 975 1836
rect 979 1832 980 1836
rect 974 1831 980 1832
rect 1046 1836 1052 1837
rect 1046 1832 1047 1836
rect 1051 1832 1052 1836
rect 1046 1831 1052 1832
rect 1126 1836 1132 1837
rect 1126 1832 1127 1836
rect 1131 1832 1132 1836
rect 1126 1831 1132 1832
rect 1190 1836 1196 1837
rect 1278 1836 1284 1837
rect 2406 1841 2412 1842
rect 2406 1837 2407 1841
rect 2411 1837 2412 1841
rect 2406 1836 2412 1837
rect 1190 1832 1191 1836
rect 1195 1832 1196 1836
rect 1190 1831 1196 1832
rect 110 1829 116 1830
rect 110 1825 111 1829
rect 115 1825 116 1829
rect 110 1824 116 1825
rect 1238 1829 1244 1830
rect 1238 1825 1239 1829
rect 1243 1825 1244 1829
rect 1238 1824 1244 1825
rect 1278 1824 1284 1825
rect 1278 1820 1279 1824
rect 1283 1820 1284 1824
rect 1278 1819 1284 1820
rect 2406 1824 2412 1825
rect 2406 1820 2407 1824
rect 2411 1820 2412 1824
rect 2406 1819 2412 1820
rect 110 1812 116 1813
rect 110 1808 111 1812
rect 115 1808 116 1812
rect 110 1807 116 1808
rect 1238 1812 1244 1813
rect 1238 1808 1239 1812
rect 1243 1808 1244 1812
rect 1238 1807 1244 1808
rect 1358 1801 1364 1802
rect 1358 1797 1359 1801
rect 1363 1797 1364 1801
rect 1358 1796 1364 1797
rect 1398 1801 1404 1802
rect 1398 1797 1399 1801
rect 1403 1797 1404 1801
rect 1398 1796 1404 1797
rect 1446 1801 1452 1802
rect 1446 1797 1447 1801
rect 1451 1797 1452 1801
rect 1446 1796 1452 1797
rect 1502 1801 1508 1802
rect 1502 1797 1503 1801
rect 1507 1797 1508 1801
rect 1502 1796 1508 1797
rect 1558 1801 1564 1802
rect 1558 1797 1559 1801
rect 1563 1797 1564 1801
rect 1558 1796 1564 1797
rect 1614 1801 1620 1802
rect 1614 1797 1615 1801
rect 1619 1797 1620 1801
rect 1614 1796 1620 1797
rect 1670 1801 1676 1802
rect 1670 1797 1671 1801
rect 1675 1797 1676 1801
rect 1670 1796 1676 1797
rect 1726 1801 1732 1802
rect 1726 1797 1727 1801
rect 1731 1797 1732 1801
rect 1726 1796 1732 1797
rect 1782 1801 1788 1802
rect 1782 1797 1783 1801
rect 1787 1797 1788 1801
rect 1782 1796 1788 1797
rect 1838 1801 1844 1802
rect 1838 1797 1839 1801
rect 1843 1797 1844 1801
rect 1838 1796 1844 1797
rect 1894 1801 1900 1802
rect 1894 1797 1895 1801
rect 1899 1797 1900 1801
rect 1894 1796 1900 1797
rect 1950 1801 1956 1802
rect 1950 1797 1951 1801
rect 1955 1797 1956 1801
rect 1950 1796 1956 1797
rect 398 1789 404 1790
rect 398 1785 399 1789
rect 403 1785 404 1789
rect 398 1784 404 1785
rect 438 1789 444 1790
rect 438 1785 439 1789
rect 443 1785 444 1789
rect 438 1784 444 1785
rect 478 1789 484 1790
rect 478 1785 479 1789
rect 483 1785 484 1789
rect 478 1784 484 1785
rect 518 1789 524 1790
rect 518 1785 519 1789
rect 523 1785 524 1789
rect 518 1784 524 1785
rect 566 1789 572 1790
rect 566 1785 567 1789
rect 571 1785 572 1789
rect 566 1784 572 1785
rect 622 1789 628 1790
rect 622 1785 623 1789
rect 627 1785 628 1789
rect 622 1784 628 1785
rect 686 1789 692 1790
rect 686 1785 687 1789
rect 691 1785 692 1789
rect 686 1784 692 1785
rect 758 1789 764 1790
rect 758 1785 759 1789
rect 763 1785 764 1789
rect 758 1784 764 1785
rect 830 1789 836 1790
rect 830 1785 831 1789
rect 835 1785 836 1789
rect 830 1784 836 1785
rect 902 1789 908 1790
rect 902 1785 903 1789
rect 907 1785 908 1789
rect 902 1784 908 1785
rect 974 1789 980 1790
rect 974 1785 975 1789
rect 979 1785 980 1789
rect 974 1784 980 1785
rect 1046 1789 1052 1790
rect 1046 1785 1047 1789
rect 1051 1785 1052 1789
rect 1046 1784 1052 1785
rect 1126 1789 1132 1790
rect 1126 1785 1127 1789
rect 1131 1785 1132 1789
rect 1126 1784 1132 1785
rect 1190 1789 1196 1790
rect 1190 1785 1191 1789
rect 1195 1785 1196 1789
rect 1190 1784 1196 1785
rect 406 1759 412 1760
rect 406 1755 407 1759
rect 411 1755 412 1759
rect 406 1754 412 1755
rect 446 1759 452 1760
rect 446 1755 447 1759
rect 451 1755 452 1759
rect 446 1754 452 1755
rect 486 1759 492 1760
rect 486 1755 487 1759
rect 491 1755 492 1759
rect 486 1754 492 1755
rect 526 1759 532 1760
rect 526 1755 527 1759
rect 531 1755 532 1759
rect 526 1754 532 1755
rect 566 1759 572 1760
rect 566 1755 567 1759
rect 571 1755 572 1759
rect 566 1754 572 1755
rect 606 1759 612 1760
rect 606 1755 607 1759
rect 611 1755 612 1759
rect 606 1754 612 1755
rect 646 1759 652 1760
rect 646 1755 647 1759
rect 651 1755 652 1759
rect 646 1754 652 1755
rect 694 1759 700 1760
rect 694 1755 695 1759
rect 699 1755 700 1759
rect 694 1754 700 1755
rect 750 1759 756 1760
rect 750 1755 751 1759
rect 755 1755 756 1759
rect 750 1754 756 1755
rect 806 1759 812 1760
rect 806 1755 807 1759
rect 811 1755 812 1759
rect 806 1754 812 1755
rect 870 1759 876 1760
rect 870 1755 871 1759
rect 875 1755 876 1759
rect 870 1754 876 1755
rect 934 1759 940 1760
rect 934 1755 935 1759
rect 939 1755 940 1759
rect 934 1754 940 1755
rect 998 1759 1004 1760
rect 998 1755 999 1759
rect 1003 1755 1004 1759
rect 998 1754 1004 1755
rect 1070 1759 1076 1760
rect 1070 1755 1071 1759
rect 1075 1755 1076 1759
rect 1070 1754 1076 1755
rect 1142 1759 1148 1760
rect 1142 1755 1143 1759
rect 1147 1755 1148 1759
rect 1142 1754 1148 1755
rect 1190 1759 1196 1760
rect 1190 1755 1191 1759
rect 1195 1755 1196 1759
rect 1190 1754 1196 1755
rect 1302 1759 1308 1760
rect 1302 1755 1303 1759
rect 1307 1755 1308 1759
rect 1302 1754 1308 1755
rect 1342 1759 1348 1760
rect 1342 1755 1343 1759
rect 1347 1755 1348 1759
rect 1342 1754 1348 1755
rect 1390 1759 1396 1760
rect 1390 1755 1391 1759
rect 1395 1755 1396 1759
rect 1390 1754 1396 1755
rect 1454 1759 1460 1760
rect 1454 1755 1455 1759
rect 1459 1755 1460 1759
rect 1454 1754 1460 1755
rect 1518 1759 1524 1760
rect 1518 1755 1519 1759
rect 1523 1755 1524 1759
rect 1518 1754 1524 1755
rect 1582 1759 1588 1760
rect 1582 1755 1583 1759
rect 1587 1755 1588 1759
rect 1582 1754 1588 1755
rect 1646 1759 1652 1760
rect 1646 1755 1647 1759
rect 1651 1755 1652 1759
rect 1646 1754 1652 1755
rect 1702 1759 1708 1760
rect 1702 1755 1703 1759
rect 1707 1755 1708 1759
rect 1702 1754 1708 1755
rect 1758 1759 1764 1760
rect 1758 1755 1759 1759
rect 1763 1755 1764 1759
rect 1758 1754 1764 1755
rect 1806 1759 1812 1760
rect 1806 1755 1807 1759
rect 1811 1755 1812 1759
rect 1806 1754 1812 1755
rect 1862 1759 1868 1760
rect 1862 1755 1863 1759
rect 1867 1755 1868 1759
rect 1862 1754 1868 1755
rect 1918 1759 1924 1760
rect 1918 1755 1919 1759
rect 1923 1755 1924 1759
rect 1918 1754 1924 1755
rect 1974 1759 1980 1760
rect 1974 1755 1975 1759
rect 1979 1755 1980 1759
rect 1974 1754 1980 1755
rect 110 1736 116 1737
rect 110 1732 111 1736
rect 115 1732 116 1736
rect 110 1731 116 1732
rect 1238 1736 1244 1737
rect 1238 1732 1239 1736
rect 1243 1732 1244 1736
rect 1238 1731 1244 1732
rect 1278 1736 1284 1737
rect 1278 1732 1279 1736
rect 1283 1732 1284 1736
rect 1278 1731 1284 1732
rect 2406 1736 2412 1737
rect 2406 1732 2407 1736
rect 2411 1732 2412 1736
rect 2406 1731 2412 1732
rect 110 1719 116 1720
rect 110 1715 111 1719
rect 115 1715 116 1719
rect 110 1714 116 1715
rect 1238 1719 1244 1720
rect 1238 1715 1239 1719
rect 1243 1715 1244 1719
rect 1238 1714 1244 1715
rect 1278 1719 1284 1720
rect 1278 1715 1279 1719
rect 1283 1715 1284 1719
rect 1278 1714 1284 1715
rect 2406 1719 2412 1720
rect 2406 1715 2407 1719
rect 2411 1715 2412 1719
rect 2406 1714 2412 1715
rect 406 1712 412 1713
rect 406 1708 407 1712
rect 411 1708 412 1712
rect 406 1707 412 1708
rect 446 1712 452 1713
rect 446 1708 447 1712
rect 451 1708 452 1712
rect 446 1707 452 1708
rect 486 1712 492 1713
rect 486 1708 487 1712
rect 491 1708 492 1712
rect 486 1707 492 1708
rect 526 1712 532 1713
rect 526 1708 527 1712
rect 531 1708 532 1712
rect 526 1707 532 1708
rect 566 1712 572 1713
rect 566 1708 567 1712
rect 571 1708 572 1712
rect 566 1707 572 1708
rect 606 1712 612 1713
rect 606 1708 607 1712
rect 611 1708 612 1712
rect 606 1707 612 1708
rect 646 1712 652 1713
rect 646 1708 647 1712
rect 651 1708 652 1712
rect 646 1707 652 1708
rect 694 1712 700 1713
rect 694 1708 695 1712
rect 699 1708 700 1712
rect 694 1707 700 1708
rect 750 1712 756 1713
rect 750 1708 751 1712
rect 755 1708 756 1712
rect 750 1707 756 1708
rect 806 1712 812 1713
rect 806 1708 807 1712
rect 811 1708 812 1712
rect 806 1707 812 1708
rect 870 1712 876 1713
rect 870 1708 871 1712
rect 875 1708 876 1712
rect 870 1707 876 1708
rect 934 1712 940 1713
rect 934 1708 935 1712
rect 939 1708 940 1712
rect 934 1707 940 1708
rect 998 1712 1004 1713
rect 998 1708 999 1712
rect 1003 1708 1004 1712
rect 998 1707 1004 1708
rect 1070 1712 1076 1713
rect 1070 1708 1071 1712
rect 1075 1708 1076 1712
rect 1070 1707 1076 1708
rect 1142 1712 1148 1713
rect 1142 1708 1143 1712
rect 1147 1708 1148 1712
rect 1142 1707 1148 1708
rect 1190 1712 1196 1713
rect 1190 1708 1191 1712
rect 1195 1708 1196 1712
rect 1190 1707 1196 1708
rect 1302 1712 1308 1713
rect 1302 1708 1303 1712
rect 1307 1708 1308 1712
rect 1302 1707 1308 1708
rect 1342 1712 1348 1713
rect 1342 1708 1343 1712
rect 1347 1708 1348 1712
rect 1342 1707 1348 1708
rect 1390 1712 1396 1713
rect 1390 1708 1391 1712
rect 1395 1708 1396 1712
rect 1390 1707 1396 1708
rect 1454 1712 1460 1713
rect 1454 1708 1455 1712
rect 1459 1708 1460 1712
rect 1454 1707 1460 1708
rect 1518 1712 1524 1713
rect 1518 1708 1519 1712
rect 1523 1708 1524 1712
rect 1518 1707 1524 1708
rect 1582 1712 1588 1713
rect 1582 1708 1583 1712
rect 1587 1708 1588 1712
rect 1582 1707 1588 1708
rect 1646 1712 1652 1713
rect 1646 1708 1647 1712
rect 1651 1708 1652 1712
rect 1646 1707 1652 1708
rect 1702 1712 1708 1713
rect 1702 1708 1703 1712
rect 1707 1708 1708 1712
rect 1702 1707 1708 1708
rect 1758 1712 1764 1713
rect 1758 1708 1759 1712
rect 1763 1708 1764 1712
rect 1758 1707 1764 1708
rect 1806 1712 1812 1713
rect 1806 1708 1807 1712
rect 1811 1708 1812 1712
rect 1806 1707 1812 1708
rect 1862 1712 1868 1713
rect 1862 1708 1863 1712
rect 1867 1708 1868 1712
rect 1862 1707 1868 1708
rect 1918 1712 1924 1713
rect 1918 1708 1919 1712
rect 1923 1708 1924 1712
rect 1918 1707 1924 1708
rect 1974 1712 1980 1713
rect 1974 1708 1975 1712
rect 1979 1708 1980 1712
rect 1974 1707 1980 1708
rect 278 1696 284 1697
rect 278 1692 279 1696
rect 283 1692 284 1696
rect 278 1691 284 1692
rect 318 1696 324 1697
rect 318 1692 319 1696
rect 323 1692 324 1696
rect 318 1691 324 1692
rect 358 1696 364 1697
rect 358 1692 359 1696
rect 363 1692 364 1696
rect 358 1691 364 1692
rect 398 1696 404 1697
rect 398 1692 399 1696
rect 403 1692 404 1696
rect 398 1691 404 1692
rect 446 1696 452 1697
rect 446 1692 447 1696
rect 451 1692 452 1696
rect 446 1691 452 1692
rect 494 1696 500 1697
rect 494 1692 495 1696
rect 499 1692 500 1696
rect 494 1691 500 1692
rect 542 1696 548 1697
rect 542 1692 543 1696
rect 547 1692 548 1696
rect 542 1691 548 1692
rect 590 1696 596 1697
rect 590 1692 591 1696
rect 595 1692 596 1696
rect 590 1691 596 1692
rect 638 1696 644 1697
rect 638 1692 639 1696
rect 643 1692 644 1696
rect 638 1691 644 1692
rect 686 1696 692 1697
rect 686 1692 687 1696
rect 691 1692 692 1696
rect 686 1691 692 1692
rect 734 1696 740 1697
rect 734 1692 735 1696
rect 739 1692 740 1696
rect 734 1691 740 1692
rect 782 1696 788 1697
rect 782 1692 783 1696
rect 787 1692 788 1696
rect 782 1691 788 1692
rect 838 1696 844 1697
rect 838 1692 839 1696
rect 843 1692 844 1696
rect 838 1691 844 1692
rect 894 1696 900 1697
rect 894 1692 895 1696
rect 899 1692 900 1696
rect 894 1691 900 1692
rect 1302 1696 1308 1697
rect 1302 1692 1303 1696
rect 1307 1692 1308 1696
rect 1302 1691 1308 1692
rect 1342 1696 1348 1697
rect 1342 1692 1343 1696
rect 1347 1692 1348 1696
rect 1342 1691 1348 1692
rect 1382 1696 1388 1697
rect 1382 1692 1383 1696
rect 1387 1692 1388 1696
rect 1382 1691 1388 1692
rect 1422 1696 1428 1697
rect 1422 1692 1423 1696
rect 1427 1692 1428 1696
rect 1422 1691 1428 1692
rect 1462 1696 1468 1697
rect 1462 1692 1463 1696
rect 1467 1692 1468 1696
rect 1462 1691 1468 1692
rect 1502 1696 1508 1697
rect 1502 1692 1503 1696
rect 1507 1692 1508 1696
rect 1502 1691 1508 1692
rect 1558 1696 1564 1697
rect 1558 1692 1559 1696
rect 1563 1692 1564 1696
rect 1558 1691 1564 1692
rect 1622 1696 1628 1697
rect 1622 1692 1623 1696
rect 1627 1692 1628 1696
rect 1622 1691 1628 1692
rect 1686 1696 1692 1697
rect 1686 1692 1687 1696
rect 1691 1692 1692 1696
rect 1686 1691 1692 1692
rect 1750 1696 1756 1697
rect 1750 1692 1751 1696
rect 1755 1692 1756 1696
rect 1750 1691 1756 1692
rect 1806 1696 1812 1697
rect 1806 1692 1807 1696
rect 1811 1692 1812 1696
rect 1806 1691 1812 1692
rect 1862 1696 1868 1697
rect 1862 1692 1863 1696
rect 1867 1692 1868 1696
rect 1862 1691 1868 1692
rect 1918 1696 1924 1697
rect 1918 1692 1919 1696
rect 1923 1692 1924 1696
rect 1918 1691 1924 1692
rect 1974 1696 1980 1697
rect 1974 1692 1975 1696
rect 1979 1692 1980 1696
rect 1974 1691 1980 1692
rect 2030 1696 2036 1697
rect 2030 1692 2031 1696
rect 2035 1692 2036 1696
rect 2030 1691 2036 1692
rect 2086 1696 2092 1697
rect 2086 1692 2087 1696
rect 2091 1692 2092 1696
rect 2086 1691 2092 1692
rect 110 1689 116 1690
rect 110 1685 111 1689
rect 115 1685 116 1689
rect 110 1684 116 1685
rect 1238 1689 1244 1690
rect 1238 1685 1239 1689
rect 1243 1685 1244 1689
rect 1238 1684 1244 1685
rect 1278 1689 1284 1690
rect 1278 1685 1279 1689
rect 1283 1685 1284 1689
rect 1278 1684 1284 1685
rect 2406 1689 2412 1690
rect 2406 1685 2407 1689
rect 2411 1685 2412 1689
rect 2406 1684 2412 1685
rect 110 1672 116 1673
rect 110 1668 111 1672
rect 115 1668 116 1672
rect 110 1667 116 1668
rect 1238 1672 1244 1673
rect 1238 1668 1239 1672
rect 1243 1668 1244 1672
rect 1238 1667 1244 1668
rect 1278 1672 1284 1673
rect 1278 1668 1279 1672
rect 1283 1668 1284 1672
rect 1278 1667 1284 1668
rect 2406 1672 2412 1673
rect 2406 1668 2407 1672
rect 2411 1668 2412 1672
rect 2406 1667 2412 1668
rect 278 1649 284 1650
rect 278 1645 279 1649
rect 283 1645 284 1649
rect 278 1644 284 1645
rect 318 1649 324 1650
rect 318 1645 319 1649
rect 323 1645 324 1649
rect 318 1644 324 1645
rect 358 1649 364 1650
rect 358 1645 359 1649
rect 363 1645 364 1649
rect 358 1644 364 1645
rect 398 1649 404 1650
rect 398 1645 399 1649
rect 403 1645 404 1649
rect 398 1644 404 1645
rect 446 1649 452 1650
rect 446 1645 447 1649
rect 451 1645 452 1649
rect 446 1644 452 1645
rect 494 1649 500 1650
rect 494 1645 495 1649
rect 499 1645 500 1649
rect 494 1644 500 1645
rect 542 1649 548 1650
rect 542 1645 543 1649
rect 547 1645 548 1649
rect 542 1644 548 1645
rect 590 1649 596 1650
rect 590 1645 591 1649
rect 595 1645 596 1649
rect 590 1644 596 1645
rect 638 1649 644 1650
rect 638 1645 639 1649
rect 643 1645 644 1649
rect 638 1644 644 1645
rect 686 1649 692 1650
rect 686 1645 687 1649
rect 691 1645 692 1649
rect 686 1644 692 1645
rect 734 1649 740 1650
rect 734 1645 735 1649
rect 739 1645 740 1649
rect 734 1644 740 1645
rect 782 1649 788 1650
rect 782 1645 783 1649
rect 787 1645 788 1649
rect 782 1644 788 1645
rect 838 1649 844 1650
rect 838 1645 839 1649
rect 843 1645 844 1649
rect 838 1644 844 1645
rect 894 1649 900 1650
rect 894 1645 895 1649
rect 899 1645 900 1649
rect 894 1644 900 1645
rect 1302 1649 1308 1650
rect 1302 1645 1303 1649
rect 1307 1645 1308 1649
rect 1302 1644 1308 1645
rect 1342 1649 1348 1650
rect 1342 1645 1343 1649
rect 1347 1645 1348 1649
rect 1342 1644 1348 1645
rect 1382 1649 1388 1650
rect 1382 1645 1383 1649
rect 1387 1645 1388 1649
rect 1382 1644 1388 1645
rect 1422 1649 1428 1650
rect 1422 1645 1423 1649
rect 1427 1645 1428 1649
rect 1422 1644 1428 1645
rect 1462 1649 1468 1650
rect 1462 1645 1463 1649
rect 1467 1645 1468 1649
rect 1462 1644 1468 1645
rect 1502 1649 1508 1650
rect 1502 1645 1503 1649
rect 1507 1645 1508 1649
rect 1502 1644 1508 1645
rect 1558 1649 1564 1650
rect 1558 1645 1559 1649
rect 1563 1645 1564 1649
rect 1558 1644 1564 1645
rect 1622 1649 1628 1650
rect 1622 1645 1623 1649
rect 1627 1645 1628 1649
rect 1622 1644 1628 1645
rect 1686 1649 1692 1650
rect 1686 1645 1687 1649
rect 1691 1645 1692 1649
rect 1686 1644 1692 1645
rect 1750 1649 1756 1650
rect 1750 1645 1751 1649
rect 1755 1645 1756 1649
rect 1750 1644 1756 1645
rect 1806 1649 1812 1650
rect 1806 1645 1807 1649
rect 1811 1645 1812 1649
rect 1806 1644 1812 1645
rect 1862 1649 1868 1650
rect 1862 1645 1863 1649
rect 1867 1645 1868 1649
rect 1862 1644 1868 1645
rect 1918 1649 1924 1650
rect 1918 1645 1919 1649
rect 1923 1645 1924 1649
rect 1918 1644 1924 1645
rect 1974 1649 1980 1650
rect 1974 1645 1975 1649
rect 1979 1645 1980 1649
rect 1974 1644 1980 1645
rect 2030 1649 2036 1650
rect 2030 1645 2031 1649
rect 2035 1645 2036 1649
rect 2030 1644 2036 1645
rect 2086 1649 2092 1650
rect 2086 1645 2087 1649
rect 2091 1645 2092 1649
rect 2086 1644 2092 1645
rect 134 1615 140 1616
rect 134 1611 135 1615
rect 139 1611 140 1615
rect 134 1610 140 1611
rect 174 1615 180 1616
rect 174 1611 175 1615
rect 179 1611 180 1615
rect 174 1610 180 1611
rect 214 1615 220 1616
rect 214 1611 215 1615
rect 219 1611 220 1615
rect 214 1610 220 1611
rect 254 1615 260 1616
rect 254 1611 255 1615
rect 259 1611 260 1615
rect 254 1610 260 1611
rect 310 1615 316 1616
rect 310 1611 311 1615
rect 315 1611 316 1615
rect 310 1610 316 1611
rect 390 1615 396 1616
rect 390 1611 391 1615
rect 395 1611 396 1615
rect 390 1610 396 1611
rect 470 1615 476 1616
rect 470 1611 471 1615
rect 475 1611 476 1615
rect 470 1610 476 1611
rect 558 1615 564 1616
rect 558 1611 559 1615
rect 563 1611 564 1615
rect 558 1610 564 1611
rect 638 1615 644 1616
rect 638 1611 639 1615
rect 643 1611 644 1615
rect 638 1610 644 1611
rect 718 1615 724 1616
rect 718 1611 719 1615
rect 723 1611 724 1615
rect 718 1610 724 1611
rect 790 1615 796 1616
rect 790 1611 791 1615
rect 795 1611 796 1615
rect 790 1610 796 1611
rect 854 1615 860 1616
rect 854 1611 855 1615
rect 859 1611 860 1615
rect 854 1610 860 1611
rect 918 1615 924 1616
rect 918 1611 919 1615
rect 923 1611 924 1615
rect 918 1610 924 1611
rect 982 1615 988 1616
rect 982 1611 983 1615
rect 987 1611 988 1615
rect 982 1610 988 1611
rect 1046 1615 1052 1616
rect 1046 1611 1047 1615
rect 1051 1611 1052 1615
rect 1046 1610 1052 1611
rect 1302 1615 1308 1616
rect 1302 1611 1303 1615
rect 1307 1611 1308 1615
rect 1302 1610 1308 1611
rect 1342 1615 1348 1616
rect 1342 1611 1343 1615
rect 1347 1611 1348 1615
rect 1342 1610 1348 1611
rect 1382 1615 1388 1616
rect 1382 1611 1383 1615
rect 1387 1611 1388 1615
rect 1382 1610 1388 1611
rect 1422 1615 1428 1616
rect 1422 1611 1423 1615
rect 1427 1611 1428 1615
rect 1422 1610 1428 1611
rect 1462 1615 1468 1616
rect 1462 1611 1463 1615
rect 1467 1611 1468 1615
rect 1462 1610 1468 1611
rect 1502 1615 1508 1616
rect 1502 1611 1503 1615
rect 1507 1611 1508 1615
rect 1502 1610 1508 1611
rect 1558 1615 1564 1616
rect 1558 1611 1559 1615
rect 1563 1611 1564 1615
rect 1558 1610 1564 1611
rect 1630 1615 1636 1616
rect 1630 1611 1631 1615
rect 1635 1611 1636 1615
rect 1630 1610 1636 1611
rect 1702 1615 1708 1616
rect 1702 1611 1703 1615
rect 1707 1611 1708 1615
rect 1702 1610 1708 1611
rect 1782 1615 1788 1616
rect 1782 1611 1783 1615
rect 1787 1611 1788 1615
rect 1782 1610 1788 1611
rect 1854 1615 1860 1616
rect 1854 1611 1855 1615
rect 1859 1611 1860 1615
rect 1854 1610 1860 1611
rect 1926 1615 1932 1616
rect 1926 1611 1927 1615
rect 1931 1611 1932 1615
rect 1926 1610 1932 1611
rect 1998 1615 2004 1616
rect 1998 1611 1999 1615
rect 2003 1611 2004 1615
rect 1998 1610 2004 1611
rect 2062 1615 2068 1616
rect 2062 1611 2063 1615
rect 2067 1611 2068 1615
rect 2062 1610 2068 1611
rect 2126 1615 2132 1616
rect 2126 1611 2127 1615
rect 2131 1611 2132 1615
rect 2126 1610 2132 1611
rect 2190 1615 2196 1616
rect 2190 1611 2191 1615
rect 2195 1611 2196 1615
rect 2190 1610 2196 1611
rect 2254 1615 2260 1616
rect 2254 1611 2255 1615
rect 2259 1611 2260 1615
rect 2254 1610 2260 1611
rect 2318 1615 2324 1616
rect 2318 1611 2319 1615
rect 2323 1611 2324 1615
rect 2318 1610 2324 1611
rect 2358 1615 2364 1616
rect 2358 1611 2359 1615
rect 2363 1611 2364 1615
rect 2358 1610 2364 1611
rect 110 1592 116 1593
rect 110 1588 111 1592
rect 115 1588 116 1592
rect 110 1587 116 1588
rect 1238 1592 1244 1593
rect 1238 1588 1239 1592
rect 1243 1588 1244 1592
rect 1238 1587 1244 1588
rect 1278 1592 1284 1593
rect 1278 1588 1279 1592
rect 1283 1588 1284 1592
rect 1278 1587 1284 1588
rect 2406 1592 2412 1593
rect 2406 1588 2407 1592
rect 2411 1588 2412 1592
rect 2406 1587 2412 1588
rect 110 1575 116 1576
rect 110 1571 111 1575
rect 115 1571 116 1575
rect 110 1570 116 1571
rect 1238 1575 1244 1576
rect 1238 1571 1239 1575
rect 1243 1571 1244 1575
rect 1238 1570 1244 1571
rect 1278 1575 1284 1576
rect 1278 1571 1279 1575
rect 1283 1571 1284 1575
rect 1278 1570 1284 1571
rect 2406 1575 2412 1576
rect 2406 1571 2407 1575
rect 2411 1571 2412 1575
rect 2406 1570 2412 1571
rect 134 1568 140 1569
rect 134 1564 135 1568
rect 139 1564 140 1568
rect 134 1563 140 1564
rect 174 1568 180 1569
rect 174 1564 175 1568
rect 179 1564 180 1568
rect 174 1563 180 1564
rect 214 1568 220 1569
rect 214 1564 215 1568
rect 219 1564 220 1568
rect 214 1563 220 1564
rect 254 1568 260 1569
rect 254 1564 255 1568
rect 259 1564 260 1568
rect 254 1563 260 1564
rect 310 1568 316 1569
rect 310 1564 311 1568
rect 315 1564 316 1568
rect 310 1563 316 1564
rect 390 1568 396 1569
rect 390 1564 391 1568
rect 395 1564 396 1568
rect 390 1563 396 1564
rect 470 1568 476 1569
rect 470 1564 471 1568
rect 475 1564 476 1568
rect 470 1563 476 1564
rect 558 1568 564 1569
rect 558 1564 559 1568
rect 563 1564 564 1568
rect 558 1563 564 1564
rect 638 1568 644 1569
rect 638 1564 639 1568
rect 643 1564 644 1568
rect 638 1563 644 1564
rect 718 1568 724 1569
rect 718 1564 719 1568
rect 723 1564 724 1568
rect 718 1563 724 1564
rect 790 1568 796 1569
rect 790 1564 791 1568
rect 795 1564 796 1568
rect 790 1563 796 1564
rect 854 1568 860 1569
rect 854 1564 855 1568
rect 859 1564 860 1568
rect 854 1563 860 1564
rect 918 1568 924 1569
rect 918 1564 919 1568
rect 923 1564 924 1568
rect 918 1563 924 1564
rect 982 1568 988 1569
rect 982 1564 983 1568
rect 987 1564 988 1568
rect 982 1563 988 1564
rect 1046 1568 1052 1569
rect 1046 1564 1047 1568
rect 1051 1564 1052 1568
rect 1046 1563 1052 1564
rect 1302 1568 1308 1569
rect 1302 1564 1303 1568
rect 1307 1564 1308 1568
rect 1302 1563 1308 1564
rect 1342 1568 1348 1569
rect 1342 1564 1343 1568
rect 1347 1564 1348 1568
rect 1342 1563 1348 1564
rect 1382 1568 1388 1569
rect 1382 1564 1383 1568
rect 1387 1564 1388 1568
rect 1382 1563 1388 1564
rect 1422 1568 1428 1569
rect 1422 1564 1423 1568
rect 1427 1564 1428 1568
rect 1422 1563 1428 1564
rect 1462 1568 1468 1569
rect 1462 1564 1463 1568
rect 1467 1564 1468 1568
rect 1462 1563 1468 1564
rect 1502 1568 1508 1569
rect 1502 1564 1503 1568
rect 1507 1564 1508 1568
rect 1502 1563 1508 1564
rect 1558 1568 1564 1569
rect 1558 1564 1559 1568
rect 1563 1564 1564 1568
rect 1558 1563 1564 1564
rect 1630 1568 1636 1569
rect 1630 1564 1631 1568
rect 1635 1564 1636 1568
rect 1630 1563 1636 1564
rect 1702 1568 1708 1569
rect 1702 1564 1703 1568
rect 1707 1564 1708 1568
rect 1702 1563 1708 1564
rect 1782 1568 1788 1569
rect 1782 1564 1783 1568
rect 1787 1564 1788 1568
rect 1782 1563 1788 1564
rect 1854 1568 1860 1569
rect 1854 1564 1855 1568
rect 1859 1564 1860 1568
rect 1854 1563 1860 1564
rect 1926 1568 1932 1569
rect 1926 1564 1927 1568
rect 1931 1564 1932 1568
rect 1926 1563 1932 1564
rect 1998 1568 2004 1569
rect 1998 1564 1999 1568
rect 2003 1564 2004 1568
rect 1998 1563 2004 1564
rect 2062 1568 2068 1569
rect 2062 1564 2063 1568
rect 2067 1564 2068 1568
rect 2062 1563 2068 1564
rect 2126 1568 2132 1569
rect 2126 1564 2127 1568
rect 2131 1564 2132 1568
rect 2126 1563 2132 1564
rect 2190 1568 2196 1569
rect 2190 1564 2191 1568
rect 2195 1564 2196 1568
rect 2190 1563 2196 1564
rect 2254 1568 2260 1569
rect 2254 1564 2255 1568
rect 2259 1564 2260 1568
rect 2254 1563 2260 1564
rect 2318 1568 2324 1569
rect 2318 1564 2319 1568
rect 2323 1564 2324 1568
rect 2318 1563 2324 1564
rect 2358 1568 2364 1569
rect 2358 1564 2359 1568
rect 2363 1564 2364 1568
rect 2358 1563 2364 1564
rect 1470 1556 1476 1557
rect 150 1552 156 1553
rect 150 1548 151 1552
rect 155 1548 156 1552
rect 150 1547 156 1548
rect 198 1552 204 1553
rect 198 1548 199 1552
rect 203 1548 204 1552
rect 198 1547 204 1548
rect 262 1552 268 1553
rect 262 1548 263 1552
rect 267 1548 268 1552
rect 262 1547 268 1548
rect 342 1552 348 1553
rect 342 1548 343 1552
rect 347 1548 348 1552
rect 342 1547 348 1548
rect 438 1552 444 1553
rect 438 1548 439 1552
rect 443 1548 444 1552
rect 438 1547 444 1548
rect 534 1552 540 1553
rect 534 1548 535 1552
rect 539 1548 540 1552
rect 534 1547 540 1548
rect 638 1552 644 1553
rect 638 1548 639 1552
rect 643 1548 644 1552
rect 638 1547 644 1548
rect 734 1552 740 1553
rect 734 1548 735 1552
rect 739 1548 740 1552
rect 734 1547 740 1548
rect 822 1552 828 1553
rect 822 1548 823 1552
rect 827 1548 828 1552
rect 822 1547 828 1548
rect 902 1552 908 1553
rect 902 1548 903 1552
rect 907 1548 908 1552
rect 902 1547 908 1548
rect 974 1552 980 1553
rect 974 1548 975 1552
rect 979 1548 980 1552
rect 974 1547 980 1548
rect 1046 1552 1052 1553
rect 1046 1548 1047 1552
rect 1051 1548 1052 1552
rect 1046 1547 1052 1548
rect 1118 1552 1124 1553
rect 1118 1548 1119 1552
rect 1123 1548 1124 1552
rect 1118 1547 1124 1548
rect 1190 1552 1196 1553
rect 1190 1548 1191 1552
rect 1195 1548 1196 1552
rect 1470 1552 1471 1556
rect 1475 1552 1476 1556
rect 1470 1551 1476 1552
rect 1622 1556 1628 1557
rect 1622 1552 1623 1556
rect 1627 1552 1628 1556
rect 1622 1551 1628 1552
rect 1758 1556 1764 1557
rect 1758 1552 1759 1556
rect 1763 1552 1764 1556
rect 1758 1551 1764 1552
rect 1870 1556 1876 1557
rect 1870 1552 1871 1556
rect 1875 1552 1876 1556
rect 1870 1551 1876 1552
rect 1966 1556 1972 1557
rect 1966 1552 1967 1556
rect 1971 1552 1972 1556
rect 1966 1551 1972 1552
rect 2054 1556 2060 1557
rect 2054 1552 2055 1556
rect 2059 1552 2060 1556
rect 2054 1551 2060 1552
rect 2126 1556 2132 1557
rect 2126 1552 2127 1556
rect 2131 1552 2132 1556
rect 2126 1551 2132 1552
rect 2190 1556 2196 1557
rect 2190 1552 2191 1556
rect 2195 1552 2196 1556
rect 2190 1551 2196 1552
rect 2254 1556 2260 1557
rect 2254 1552 2255 1556
rect 2259 1552 2260 1556
rect 2254 1551 2260 1552
rect 2318 1556 2324 1557
rect 2318 1552 2319 1556
rect 2323 1552 2324 1556
rect 2318 1551 2324 1552
rect 2358 1556 2364 1557
rect 2358 1552 2359 1556
rect 2363 1552 2364 1556
rect 2358 1551 2364 1552
rect 1190 1547 1196 1548
rect 1278 1549 1284 1550
rect 110 1545 116 1546
rect 110 1541 111 1545
rect 115 1541 116 1545
rect 110 1540 116 1541
rect 1238 1545 1244 1546
rect 1238 1541 1239 1545
rect 1243 1541 1244 1545
rect 1278 1545 1279 1549
rect 1283 1545 1284 1549
rect 1278 1544 1284 1545
rect 2406 1549 2412 1550
rect 2406 1545 2407 1549
rect 2411 1545 2412 1549
rect 2406 1544 2412 1545
rect 1238 1540 1244 1541
rect 1278 1532 1284 1533
rect 110 1528 116 1529
rect 110 1524 111 1528
rect 115 1524 116 1528
rect 110 1523 116 1524
rect 1238 1528 1244 1529
rect 1238 1524 1239 1528
rect 1243 1524 1244 1528
rect 1278 1528 1279 1532
rect 1283 1528 1284 1532
rect 1278 1527 1284 1528
rect 2406 1532 2412 1533
rect 2406 1528 2407 1532
rect 2411 1528 2412 1532
rect 2406 1527 2412 1528
rect 1238 1523 1244 1524
rect 1470 1509 1476 1510
rect 150 1505 156 1506
rect 150 1501 151 1505
rect 155 1501 156 1505
rect 150 1500 156 1501
rect 198 1505 204 1506
rect 198 1501 199 1505
rect 203 1501 204 1505
rect 198 1500 204 1501
rect 262 1505 268 1506
rect 262 1501 263 1505
rect 267 1501 268 1505
rect 262 1500 268 1501
rect 342 1505 348 1506
rect 342 1501 343 1505
rect 347 1501 348 1505
rect 342 1500 348 1501
rect 438 1505 444 1506
rect 438 1501 439 1505
rect 443 1501 444 1505
rect 438 1500 444 1501
rect 534 1505 540 1506
rect 534 1501 535 1505
rect 539 1501 540 1505
rect 534 1500 540 1501
rect 638 1505 644 1506
rect 638 1501 639 1505
rect 643 1501 644 1505
rect 638 1500 644 1501
rect 734 1505 740 1506
rect 734 1501 735 1505
rect 739 1501 740 1505
rect 734 1500 740 1501
rect 822 1505 828 1506
rect 822 1501 823 1505
rect 827 1501 828 1505
rect 822 1500 828 1501
rect 902 1505 908 1506
rect 902 1501 903 1505
rect 907 1501 908 1505
rect 902 1500 908 1501
rect 974 1505 980 1506
rect 974 1501 975 1505
rect 979 1501 980 1505
rect 974 1500 980 1501
rect 1046 1505 1052 1506
rect 1046 1501 1047 1505
rect 1051 1501 1052 1505
rect 1046 1500 1052 1501
rect 1118 1505 1124 1506
rect 1118 1501 1119 1505
rect 1123 1501 1124 1505
rect 1118 1500 1124 1501
rect 1190 1505 1196 1506
rect 1190 1501 1191 1505
rect 1195 1501 1196 1505
rect 1470 1505 1471 1509
rect 1475 1505 1476 1509
rect 1470 1504 1476 1505
rect 1622 1509 1628 1510
rect 1622 1505 1623 1509
rect 1627 1505 1628 1509
rect 1622 1504 1628 1505
rect 1758 1509 1764 1510
rect 1758 1505 1759 1509
rect 1763 1505 1764 1509
rect 1758 1504 1764 1505
rect 1870 1509 1876 1510
rect 1870 1505 1871 1509
rect 1875 1505 1876 1509
rect 1870 1504 1876 1505
rect 1966 1509 1972 1510
rect 1966 1505 1967 1509
rect 1971 1505 1972 1509
rect 1966 1504 1972 1505
rect 2054 1509 2060 1510
rect 2054 1505 2055 1509
rect 2059 1505 2060 1509
rect 2054 1504 2060 1505
rect 2126 1509 2132 1510
rect 2126 1505 2127 1509
rect 2131 1505 2132 1509
rect 2126 1504 2132 1505
rect 2190 1509 2196 1510
rect 2190 1505 2191 1509
rect 2195 1505 2196 1509
rect 2190 1504 2196 1505
rect 2254 1509 2260 1510
rect 2254 1505 2255 1509
rect 2259 1505 2260 1509
rect 2254 1504 2260 1505
rect 2318 1509 2324 1510
rect 2318 1505 2319 1509
rect 2323 1505 2324 1509
rect 2318 1504 2324 1505
rect 2358 1509 2364 1510
rect 2358 1505 2359 1509
rect 2363 1505 2364 1509
rect 2358 1504 2364 1505
rect 1190 1500 1196 1501
rect 318 1471 324 1472
rect 318 1467 319 1471
rect 323 1467 324 1471
rect 318 1466 324 1467
rect 358 1471 364 1472
rect 358 1467 359 1471
rect 363 1467 364 1471
rect 358 1466 364 1467
rect 398 1471 404 1472
rect 398 1467 399 1471
rect 403 1467 404 1471
rect 398 1466 404 1467
rect 446 1471 452 1472
rect 446 1467 447 1471
rect 451 1467 452 1471
rect 446 1466 452 1467
rect 502 1471 508 1472
rect 502 1467 503 1471
rect 507 1467 508 1471
rect 502 1466 508 1467
rect 558 1471 564 1472
rect 558 1467 559 1471
rect 563 1467 564 1471
rect 558 1466 564 1467
rect 614 1471 620 1472
rect 614 1467 615 1471
rect 619 1467 620 1471
rect 614 1466 620 1467
rect 670 1471 676 1472
rect 670 1467 671 1471
rect 675 1467 676 1471
rect 670 1466 676 1467
rect 734 1471 740 1472
rect 734 1467 735 1471
rect 739 1467 740 1471
rect 734 1466 740 1467
rect 798 1471 804 1472
rect 798 1467 799 1471
rect 803 1467 804 1471
rect 798 1466 804 1467
rect 854 1471 860 1472
rect 854 1467 855 1471
rect 859 1467 860 1471
rect 854 1466 860 1467
rect 910 1471 916 1472
rect 910 1467 911 1471
rect 915 1467 916 1471
rect 910 1466 916 1467
rect 966 1471 972 1472
rect 966 1467 967 1471
rect 971 1467 972 1471
rect 966 1466 972 1467
rect 1022 1471 1028 1472
rect 1022 1467 1023 1471
rect 1027 1467 1028 1471
rect 1022 1466 1028 1467
rect 1086 1471 1092 1472
rect 1086 1467 1087 1471
rect 1091 1467 1092 1471
rect 1086 1466 1092 1467
rect 1150 1471 1156 1472
rect 1150 1467 1151 1471
rect 1155 1467 1156 1471
rect 1150 1466 1156 1467
rect 1190 1471 1196 1472
rect 1190 1467 1191 1471
rect 1195 1467 1196 1471
rect 1190 1466 1196 1467
rect 1302 1459 1308 1460
rect 1302 1455 1303 1459
rect 1307 1455 1308 1459
rect 1302 1454 1308 1455
rect 1374 1459 1380 1460
rect 1374 1455 1375 1459
rect 1379 1455 1380 1459
rect 1374 1454 1380 1455
rect 1478 1459 1484 1460
rect 1478 1455 1479 1459
rect 1483 1455 1484 1459
rect 1478 1454 1484 1455
rect 1582 1459 1588 1460
rect 1582 1455 1583 1459
rect 1587 1455 1588 1459
rect 1582 1454 1588 1455
rect 1686 1459 1692 1460
rect 1686 1455 1687 1459
rect 1691 1455 1692 1459
rect 1686 1454 1692 1455
rect 1782 1459 1788 1460
rect 1782 1455 1783 1459
rect 1787 1455 1788 1459
rect 1782 1454 1788 1455
rect 1870 1459 1876 1460
rect 1870 1455 1871 1459
rect 1875 1455 1876 1459
rect 1870 1454 1876 1455
rect 1950 1459 1956 1460
rect 1950 1455 1951 1459
rect 1955 1455 1956 1459
rect 1950 1454 1956 1455
rect 2030 1459 2036 1460
rect 2030 1455 2031 1459
rect 2035 1455 2036 1459
rect 2030 1454 2036 1455
rect 2102 1459 2108 1460
rect 2102 1455 2103 1459
rect 2107 1455 2108 1459
rect 2102 1454 2108 1455
rect 2166 1459 2172 1460
rect 2166 1455 2167 1459
rect 2171 1455 2172 1459
rect 2166 1454 2172 1455
rect 2238 1459 2244 1460
rect 2238 1455 2239 1459
rect 2243 1455 2244 1459
rect 2238 1454 2244 1455
rect 2310 1459 2316 1460
rect 2310 1455 2311 1459
rect 2315 1455 2316 1459
rect 2310 1454 2316 1455
rect 2358 1459 2364 1460
rect 2358 1455 2359 1459
rect 2363 1455 2364 1459
rect 2358 1454 2364 1455
rect 110 1448 116 1449
rect 110 1444 111 1448
rect 115 1444 116 1448
rect 110 1443 116 1444
rect 1238 1448 1244 1449
rect 1238 1444 1239 1448
rect 1243 1444 1244 1448
rect 1238 1443 1244 1444
rect 1278 1436 1284 1437
rect 1278 1432 1279 1436
rect 1283 1432 1284 1436
rect 110 1431 116 1432
rect 110 1427 111 1431
rect 115 1427 116 1431
rect 110 1426 116 1427
rect 1238 1431 1244 1432
rect 1278 1431 1284 1432
rect 2406 1436 2412 1437
rect 2406 1432 2407 1436
rect 2411 1432 2412 1436
rect 2406 1431 2412 1432
rect 1238 1427 1239 1431
rect 1243 1427 1244 1431
rect 1238 1426 1244 1427
rect 318 1424 324 1425
rect 318 1420 319 1424
rect 323 1420 324 1424
rect 318 1419 324 1420
rect 358 1424 364 1425
rect 358 1420 359 1424
rect 363 1420 364 1424
rect 358 1419 364 1420
rect 398 1424 404 1425
rect 398 1420 399 1424
rect 403 1420 404 1424
rect 398 1419 404 1420
rect 446 1424 452 1425
rect 446 1420 447 1424
rect 451 1420 452 1424
rect 446 1419 452 1420
rect 502 1424 508 1425
rect 502 1420 503 1424
rect 507 1420 508 1424
rect 502 1419 508 1420
rect 558 1424 564 1425
rect 558 1420 559 1424
rect 563 1420 564 1424
rect 558 1419 564 1420
rect 614 1424 620 1425
rect 614 1420 615 1424
rect 619 1420 620 1424
rect 614 1419 620 1420
rect 670 1424 676 1425
rect 670 1420 671 1424
rect 675 1420 676 1424
rect 670 1419 676 1420
rect 734 1424 740 1425
rect 734 1420 735 1424
rect 739 1420 740 1424
rect 734 1419 740 1420
rect 798 1424 804 1425
rect 798 1420 799 1424
rect 803 1420 804 1424
rect 798 1419 804 1420
rect 854 1424 860 1425
rect 854 1420 855 1424
rect 859 1420 860 1424
rect 854 1419 860 1420
rect 910 1424 916 1425
rect 910 1420 911 1424
rect 915 1420 916 1424
rect 910 1419 916 1420
rect 966 1424 972 1425
rect 966 1420 967 1424
rect 971 1420 972 1424
rect 966 1419 972 1420
rect 1022 1424 1028 1425
rect 1022 1420 1023 1424
rect 1027 1420 1028 1424
rect 1022 1419 1028 1420
rect 1086 1424 1092 1425
rect 1086 1420 1087 1424
rect 1091 1420 1092 1424
rect 1086 1419 1092 1420
rect 1150 1424 1156 1425
rect 1150 1420 1151 1424
rect 1155 1420 1156 1424
rect 1150 1419 1156 1420
rect 1190 1424 1196 1425
rect 1190 1420 1191 1424
rect 1195 1420 1196 1424
rect 1190 1419 1196 1420
rect 1278 1419 1284 1420
rect 1278 1415 1279 1419
rect 1283 1415 1284 1419
rect 1278 1414 1284 1415
rect 2406 1419 2412 1420
rect 2406 1415 2407 1419
rect 2411 1415 2412 1419
rect 2406 1414 2412 1415
rect 1302 1412 1308 1413
rect 262 1408 268 1409
rect 262 1404 263 1408
rect 267 1404 268 1408
rect 262 1403 268 1404
rect 302 1408 308 1409
rect 302 1404 303 1408
rect 307 1404 308 1408
rect 302 1403 308 1404
rect 342 1408 348 1409
rect 342 1404 343 1408
rect 347 1404 348 1408
rect 342 1403 348 1404
rect 390 1408 396 1409
rect 390 1404 391 1408
rect 395 1404 396 1408
rect 390 1403 396 1404
rect 446 1408 452 1409
rect 446 1404 447 1408
rect 451 1404 452 1408
rect 446 1403 452 1404
rect 502 1408 508 1409
rect 502 1404 503 1408
rect 507 1404 508 1408
rect 502 1403 508 1404
rect 558 1408 564 1409
rect 558 1404 559 1408
rect 563 1404 564 1408
rect 558 1403 564 1404
rect 622 1408 628 1409
rect 622 1404 623 1408
rect 627 1404 628 1408
rect 622 1403 628 1404
rect 686 1408 692 1409
rect 686 1404 687 1408
rect 691 1404 692 1408
rect 686 1403 692 1404
rect 750 1408 756 1409
rect 750 1404 751 1408
rect 755 1404 756 1408
rect 750 1403 756 1404
rect 814 1408 820 1409
rect 814 1404 815 1408
rect 819 1404 820 1408
rect 814 1403 820 1404
rect 878 1408 884 1409
rect 878 1404 879 1408
rect 883 1404 884 1408
rect 878 1403 884 1404
rect 950 1408 956 1409
rect 950 1404 951 1408
rect 955 1404 956 1408
rect 950 1403 956 1404
rect 1022 1408 1028 1409
rect 1022 1404 1023 1408
rect 1027 1404 1028 1408
rect 1302 1408 1303 1412
rect 1307 1408 1308 1412
rect 1302 1407 1308 1408
rect 1374 1412 1380 1413
rect 1374 1408 1375 1412
rect 1379 1408 1380 1412
rect 1374 1407 1380 1408
rect 1478 1412 1484 1413
rect 1478 1408 1479 1412
rect 1483 1408 1484 1412
rect 1478 1407 1484 1408
rect 1582 1412 1588 1413
rect 1582 1408 1583 1412
rect 1587 1408 1588 1412
rect 1582 1407 1588 1408
rect 1686 1412 1692 1413
rect 1686 1408 1687 1412
rect 1691 1408 1692 1412
rect 1686 1407 1692 1408
rect 1782 1412 1788 1413
rect 1782 1408 1783 1412
rect 1787 1408 1788 1412
rect 1782 1407 1788 1408
rect 1870 1412 1876 1413
rect 1870 1408 1871 1412
rect 1875 1408 1876 1412
rect 1870 1407 1876 1408
rect 1950 1412 1956 1413
rect 1950 1408 1951 1412
rect 1955 1408 1956 1412
rect 1950 1407 1956 1408
rect 2030 1412 2036 1413
rect 2030 1408 2031 1412
rect 2035 1408 2036 1412
rect 2030 1407 2036 1408
rect 2102 1412 2108 1413
rect 2102 1408 2103 1412
rect 2107 1408 2108 1412
rect 2102 1407 2108 1408
rect 2166 1412 2172 1413
rect 2166 1408 2167 1412
rect 2171 1408 2172 1412
rect 2166 1407 2172 1408
rect 2238 1412 2244 1413
rect 2238 1408 2239 1412
rect 2243 1408 2244 1412
rect 2238 1407 2244 1408
rect 2310 1412 2316 1413
rect 2310 1408 2311 1412
rect 2315 1408 2316 1412
rect 2310 1407 2316 1408
rect 2358 1412 2364 1413
rect 2358 1408 2359 1412
rect 2363 1408 2364 1412
rect 2358 1407 2364 1408
rect 1022 1403 1028 1404
rect 110 1401 116 1402
rect 110 1397 111 1401
rect 115 1397 116 1401
rect 110 1396 116 1397
rect 1238 1401 1244 1402
rect 1238 1397 1239 1401
rect 1243 1397 1244 1401
rect 1238 1396 1244 1397
rect 1302 1400 1308 1401
rect 1302 1396 1303 1400
rect 1307 1396 1308 1400
rect 1302 1395 1308 1396
rect 1342 1400 1348 1401
rect 1342 1396 1343 1400
rect 1347 1396 1348 1400
rect 1342 1395 1348 1396
rect 1398 1400 1404 1401
rect 1398 1396 1399 1400
rect 1403 1396 1404 1400
rect 1398 1395 1404 1396
rect 1470 1400 1476 1401
rect 1470 1396 1471 1400
rect 1475 1396 1476 1400
rect 1470 1395 1476 1396
rect 1550 1400 1556 1401
rect 1550 1396 1551 1400
rect 1555 1396 1556 1400
rect 1550 1395 1556 1396
rect 1638 1400 1644 1401
rect 1638 1396 1639 1400
rect 1643 1396 1644 1400
rect 1638 1395 1644 1396
rect 1726 1400 1732 1401
rect 1726 1396 1727 1400
rect 1731 1396 1732 1400
rect 1726 1395 1732 1396
rect 1814 1400 1820 1401
rect 1814 1396 1815 1400
rect 1819 1396 1820 1400
rect 1814 1395 1820 1396
rect 1902 1400 1908 1401
rect 1902 1396 1903 1400
rect 1907 1396 1908 1400
rect 1902 1395 1908 1396
rect 1990 1400 1996 1401
rect 1990 1396 1991 1400
rect 1995 1396 1996 1400
rect 1990 1395 1996 1396
rect 2070 1400 2076 1401
rect 2070 1396 2071 1400
rect 2075 1396 2076 1400
rect 2070 1395 2076 1396
rect 2150 1400 2156 1401
rect 2150 1396 2151 1400
rect 2155 1396 2156 1400
rect 2150 1395 2156 1396
rect 2222 1400 2228 1401
rect 2222 1396 2223 1400
rect 2227 1396 2228 1400
rect 2222 1395 2228 1396
rect 2302 1400 2308 1401
rect 2302 1396 2303 1400
rect 2307 1396 2308 1400
rect 2302 1395 2308 1396
rect 2358 1400 2364 1401
rect 2358 1396 2359 1400
rect 2363 1396 2364 1400
rect 2358 1395 2364 1396
rect 1278 1393 1284 1394
rect 1278 1389 1279 1393
rect 1283 1389 1284 1393
rect 1278 1388 1284 1389
rect 2406 1393 2412 1394
rect 2406 1389 2407 1393
rect 2411 1389 2412 1393
rect 2406 1388 2412 1389
rect 110 1384 116 1385
rect 110 1380 111 1384
rect 115 1380 116 1384
rect 110 1379 116 1380
rect 1238 1384 1244 1385
rect 1238 1380 1239 1384
rect 1243 1380 1244 1384
rect 1238 1379 1244 1380
rect 1278 1376 1284 1377
rect 1278 1372 1279 1376
rect 1283 1372 1284 1376
rect 1278 1371 1284 1372
rect 2406 1376 2412 1377
rect 2406 1372 2407 1376
rect 2411 1372 2412 1376
rect 2406 1371 2412 1372
rect 262 1361 268 1362
rect 262 1357 263 1361
rect 267 1357 268 1361
rect 262 1356 268 1357
rect 302 1361 308 1362
rect 302 1357 303 1361
rect 307 1357 308 1361
rect 302 1356 308 1357
rect 342 1361 348 1362
rect 342 1357 343 1361
rect 347 1357 348 1361
rect 342 1356 348 1357
rect 390 1361 396 1362
rect 390 1357 391 1361
rect 395 1357 396 1361
rect 390 1356 396 1357
rect 446 1361 452 1362
rect 446 1357 447 1361
rect 451 1357 452 1361
rect 446 1356 452 1357
rect 502 1361 508 1362
rect 502 1357 503 1361
rect 507 1357 508 1361
rect 502 1356 508 1357
rect 558 1361 564 1362
rect 558 1357 559 1361
rect 563 1357 564 1361
rect 558 1356 564 1357
rect 622 1361 628 1362
rect 622 1357 623 1361
rect 627 1357 628 1361
rect 622 1356 628 1357
rect 686 1361 692 1362
rect 686 1357 687 1361
rect 691 1357 692 1361
rect 686 1356 692 1357
rect 750 1361 756 1362
rect 750 1357 751 1361
rect 755 1357 756 1361
rect 750 1356 756 1357
rect 814 1361 820 1362
rect 814 1357 815 1361
rect 819 1357 820 1361
rect 814 1356 820 1357
rect 878 1361 884 1362
rect 878 1357 879 1361
rect 883 1357 884 1361
rect 878 1356 884 1357
rect 950 1361 956 1362
rect 950 1357 951 1361
rect 955 1357 956 1361
rect 950 1356 956 1357
rect 1022 1361 1028 1362
rect 1022 1357 1023 1361
rect 1027 1357 1028 1361
rect 1022 1356 1028 1357
rect 1302 1353 1308 1354
rect 1302 1349 1303 1353
rect 1307 1349 1308 1353
rect 1302 1348 1308 1349
rect 1342 1353 1348 1354
rect 1342 1349 1343 1353
rect 1347 1349 1348 1353
rect 1342 1348 1348 1349
rect 1398 1353 1404 1354
rect 1398 1349 1399 1353
rect 1403 1349 1404 1353
rect 1398 1348 1404 1349
rect 1470 1353 1476 1354
rect 1470 1349 1471 1353
rect 1475 1349 1476 1353
rect 1470 1348 1476 1349
rect 1550 1353 1556 1354
rect 1550 1349 1551 1353
rect 1555 1349 1556 1353
rect 1550 1348 1556 1349
rect 1638 1353 1644 1354
rect 1638 1349 1639 1353
rect 1643 1349 1644 1353
rect 1638 1348 1644 1349
rect 1726 1353 1732 1354
rect 1726 1349 1727 1353
rect 1731 1349 1732 1353
rect 1726 1348 1732 1349
rect 1814 1353 1820 1354
rect 1814 1349 1815 1353
rect 1819 1349 1820 1353
rect 1814 1348 1820 1349
rect 1902 1353 1908 1354
rect 1902 1349 1903 1353
rect 1907 1349 1908 1353
rect 1902 1348 1908 1349
rect 1990 1353 1996 1354
rect 1990 1349 1991 1353
rect 1995 1349 1996 1353
rect 1990 1348 1996 1349
rect 2070 1353 2076 1354
rect 2070 1349 2071 1353
rect 2075 1349 2076 1353
rect 2070 1348 2076 1349
rect 2150 1353 2156 1354
rect 2150 1349 2151 1353
rect 2155 1349 2156 1353
rect 2150 1348 2156 1349
rect 2222 1353 2228 1354
rect 2222 1349 2223 1353
rect 2227 1349 2228 1353
rect 2222 1348 2228 1349
rect 2302 1353 2308 1354
rect 2302 1349 2303 1353
rect 2307 1349 2308 1353
rect 2302 1348 2308 1349
rect 2358 1353 2364 1354
rect 2358 1349 2359 1353
rect 2363 1349 2364 1353
rect 2358 1348 2364 1349
rect 134 1327 140 1328
rect 134 1323 135 1327
rect 139 1323 140 1327
rect 134 1322 140 1323
rect 174 1327 180 1328
rect 174 1323 175 1327
rect 179 1323 180 1327
rect 174 1322 180 1323
rect 214 1327 220 1328
rect 214 1323 215 1327
rect 219 1323 220 1327
rect 214 1322 220 1323
rect 254 1327 260 1328
rect 254 1323 255 1327
rect 259 1323 260 1327
rect 254 1322 260 1323
rect 326 1327 332 1328
rect 326 1323 327 1327
rect 331 1323 332 1327
rect 326 1322 332 1323
rect 406 1327 412 1328
rect 406 1323 407 1327
rect 411 1323 412 1327
rect 406 1322 412 1323
rect 494 1327 500 1328
rect 494 1323 495 1327
rect 499 1323 500 1327
rect 494 1322 500 1323
rect 582 1327 588 1328
rect 582 1323 583 1327
rect 587 1323 588 1327
rect 582 1322 588 1323
rect 670 1327 676 1328
rect 670 1323 671 1327
rect 675 1323 676 1327
rect 670 1322 676 1323
rect 758 1327 764 1328
rect 758 1323 759 1327
rect 763 1323 764 1327
rect 758 1322 764 1323
rect 838 1327 844 1328
rect 838 1323 839 1327
rect 843 1323 844 1327
rect 838 1322 844 1323
rect 918 1327 924 1328
rect 918 1323 919 1327
rect 923 1323 924 1327
rect 918 1322 924 1323
rect 1006 1327 1012 1328
rect 1006 1323 1007 1327
rect 1011 1323 1012 1327
rect 1006 1322 1012 1323
rect 1094 1327 1100 1328
rect 1094 1323 1095 1327
rect 1099 1323 1100 1327
rect 1094 1322 1100 1323
rect 1446 1319 1452 1320
rect 1446 1315 1447 1319
rect 1451 1315 1452 1319
rect 1446 1314 1452 1315
rect 1486 1319 1492 1320
rect 1486 1315 1487 1319
rect 1491 1315 1492 1319
rect 1486 1314 1492 1315
rect 1526 1319 1532 1320
rect 1526 1315 1527 1319
rect 1531 1315 1532 1319
rect 1526 1314 1532 1315
rect 1566 1319 1572 1320
rect 1566 1315 1567 1319
rect 1571 1315 1572 1319
rect 1566 1314 1572 1315
rect 1614 1319 1620 1320
rect 1614 1315 1615 1319
rect 1619 1315 1620 1319
rect 1614 1314 1620 1315
rect 1670 1319 1676 1320
rect 1670 1315 1671 1319
rect 1675 1315 1676 1319
rect 1670 1314 1676 1315
rect 1718 1319 1724 1320
rect 1718 1315 1719 1319
rect 1723 1315 1724 1319
rect 1718 1314 1724 1315
rect 1774 1319 1780 1320
rect 1774 1315 1775 1319
rect 1779 1315 1780 1319
rect 1774 1314 1780 1315
rect 1830 1319 1836 1320
rect 1830 1315 1831 1319
rect 1835 1315 1836 1319
rect 1830 1314 1836 1315
rect 1902 1319 1908 1320
rect 1902 1315 1903 1319
rect 1907 1315 1908 1319
rect 1902 1314 1908 1315
rect 1982 1319 1988 1320
rect 1982 1315 1983 1319
rect 1987 1315 1988 1319
rect 1982 1314 1988 1315
rect 2070 1319 2076 1320
rect 2070 1315 2071 1319
rect 2075 1315 2076 1319
rect 2070 1314 2076 1315
rect 2166 1319 2172 1320
rect 2166 1315 2167 1319
rect 2171 1315 2172 1319
rect 2166 1314 2172 1315
rect 2270 1319 2276 1320
rect 2270 1315 2271 1319
rect 2275 1315 2276 1319
rect 2270 1314 2276 1315
rect 2358 1319 2364 1320
rect 2358 1315 2359 1319
rect 2363 1315 2364 1319
rect 2358 1314 2364 1315
rect 110 1304 116 1305
rect 110 1300 111 1304
rect 115 1300 116 1304
rect 110 1299 116 1300
rect 1238 1304 1244 1305
rect 1238 1300 1239 1304
rect 1243 1300 1244 1304
rect 1238 1299 1244 1300
rect 1278 1296 1284 1297
rect 1278 1292 1279 1296
rect 1283 1292 1284 1296
rect 1278 1291 1284 1292
rect 2406 1296 2412 1297
rect 2406 1292 2407 1296
rect 2411 1292 2412 1296
rect 2406 1291 2412 1292
rect 110 1287 116 1288
rect 110 1283 111 1287
rect 115 1283 116 1287
rect 110 1282 116 1283
rect 1238 1287 1244 1288
rect 1238 1283 1239 1287
rect 1243 1283 1244 1287
rect 1238 1282 1244 1283
rect 134 1280 140 1281
rect 134 1276 135 1280
rect 139 1276 140 1280
rect 134 1275 140 1276
rect 174 1280 180 1281
rect 174 1276 175 1280
rect 179 1276 180 1280
rect 174 1275 180 1276
rect 214 1280 220 1281
rect 214 1276 215 1280
rect 219 1276 220 1280
rect 214 1275 220 1276
rect 254 1280 260 1281
rect 254 1276 255 1280
rect 259 1276 260 1280
rect 254 1275 260 1276
rect 326 1280 332 1281
rect 326 1276 327 1280
rect 331 1276 332 1280
rect 326 1275 332 1276
rect 406 1280 412 1281
rect 406 1276 407 1280
rect 411 1276 412 1280
rect 406 1275 412 1276
rect 494 1280 500 1281
rect 494 1276 495 1280
rect 499 1276 500 1280
rect 494 1275 500 1276
rect 582 1280 588 1281
rect 582 1276 583 1280
rect 587 1276 588 1280
rect 582 1275 588 1276
rect 670 1280 676 1281
rect 670 1276 671 1280
rect 675 1276 676 1280
rect 670 1275 676 1276
rect 758 1280 764 1281
rect 758 1276 759 1280
rect 763 1276 764 1280
rect 758 1275 764 1276
rect 838 1280 844 1281
rect 838 1276 839 1280
rect 843 1276 844 1280
rect 838 1275 844 1276
rect 918 1280 924 1281
rect 918 1276 919 1280
rect 923 1276 924 1280
rect 918 1275 924 1276
rect 1006 1280 1012 1281
rect 1006 1276 1007 1280
rect 1011 1276 1012 1280
rect 1006 1275 1012 1276
rect 1094 1280 1100 1281
rect 1094 1276 1095 1280
rect 1099 1276 1100 1280
rect 1094 1275 1100 1276
rect 1278 1279 1284 1280
rect 1278 1275 1279 1279
rect 1283 1275 1284 1279
rect 1278 1274 1284 1275
rect 2406 1279 2412 1280
rect 2406 1275 2407 1279
rect 2411 1275 2412 1279
rect 2406 1274 2412 1275
rect 1446 1272 1452 1273
rect 1446 1268 1447 1272
rect 1451 1268 1452 1272
rect 1446 1267 1452 1268
rect 1486 1272 1492 1273
rect 1486 1268 1487 1272
rect 1491 1268 1492 1272
rect 1486 1267 1492 1268
rect 1526 1272 1532 1273
rect 1526 1268 1527 1272
rect 1531 1268 1532 1272
rect 1526 1267 1532 1268
rect 1566 1272 1572 1273
rect 1566 1268 1567 1272
rect 1571 1268 1572 1272
rect 1566 1267 1572 1268
rect 1614 1272 1620 1273
rect 1614 1268 1615 1272
rect 1619 1268 1620 1272
rect 1614 1267 1620 1268
rect 1670 1272 1676 1273
rect 1670 1268 1671 1272
rect 1675 1268 1676 1272
rect 1670 1267 1676 1268
rect 1718 1272 1724 1273
rect 1718 1268 1719 1272
rect 1723 1268 1724 1272
rect 1718 1267 1724 1268
rect 1774 1272 1780 1273
rect 1774 1268 1775 1272
rect 1779 1268 1780 1272
rect 1774 1267 1780 1268
rect 1830 1272 1836 1273
rect 1830 1268 1831 1272
rect 1835 1268 1836 1272
rect 1830 1267 1836 1268
rect 1902 1272 1908 1273
rect 1902 1268 1903 1272
rect 1907 1268 1908 1272
rect 1902 1267 1908 1268
rect 1982 1272 1988 1273
rect 1982 1268 1983 1272
rect 1987 1268 1988 1272
rect 1982 1267 1988 1268
rect 2070 1272 2076 1273
rect 2070 1268 2071 1272
rect 2075 1268 2076 1272
rect 2070 1267 2076 1268
rect 2166 1272 2172 1273
rect 2166 1268 2167 1272
rect 2171 1268 2172 1272
rect 2166 1267 2172 1268
rect 2270 1272 2276 1273
rect 2270 1268 2271 1272
rect 2275 1268 2276 1272
rect 2270 1267 2276 1268
rect 2358 1272 2364 1273
rect 2358 1268 2359 1272
rect 2363 1268 2364 1272
rect 2358 1267 2364 1268
rect 134 1264 140 1265
rect 134 1260 135 1264
rect 139 1260 140 1264
rect 134 1259 140 1260
rect 174 1264 180 1265
rect 174 1260 175 1264
rect 179 1260 180 1264
rect 174 1259 180 1260
rect 246 1264 252 1265
rect 246 1260 247 1264
rect 251 1260 252 1264
rect 246 1259 252 1260
rect 326 1264 332 1265
rect 326 1260 327 1264
rect 331 1260 332 1264
rect 326 1259 332 1260
rect 414 1264 420 1265
rect 414 1260 415 1264
rect 419 1260 420 1264
rect 414 1259 420 1260
rect 502 1264 508 1265
rect 502 1260 503 1264
rect 507 1260 508 1264
rect 502 1259 508 1260
rect 590 1264 596 1265
rect 590 1260 591 1264
rect 595 1260 596 1264
rect 590 1259 596 1260
rect 670 1264 676 1265
rect 670 1260 671 1264
rect 675 1260 676 1264
rect 670 1259 676 1260
rect 742 1264 748 1265
rect 742 1260 743 1264
rect 747 1260 748 1264
rect 742 1259 748 1260
rect 814 1264 820 1265
rect 814 1260 815 1264
rect 819 1260 820 1264
rect 814 1259 820 1260
rect 878 1264 884 1265
rect 878 1260 879 1264
rect 883 1260 884 1264
rect 878 1259 884 1260
rect 942 1264 948 1265
rect 942 1260 943 1264
rect 947 1260 948 1264
rect 942 1259 948 1260
rect 1006 1264 1012 1265
rect 1006 1260 1007 1264
rect 1011 1260 1012 1264
rect 1006 1259 1012 1260
rect 1070 1264 1076 1265
rect 1070 1260 1071 1264
rect 1075 1260 1076 1264
rect 1070 1259 1076 1260
rect 110 1257 116 1258
rect 110 1253 111 1257
rect 115 1253 116 1257
rect 110 1252 116 1253
rect 1238 1257 1244 1258
rect 1238 1253 1239 1257
rect 1243 1253 1244 1257
rect 1238 1252 1244 1253
rect 1510 1256 1516 1257
rect 1510 1252 1511 1256
rect 1515 1252 1516 1256
rect 1510 1251 1516 1252
rect 1550 1256 1556 1257
rect 1550 1252 1551 1256
rect 1555 1252 1556 1256
rect 1550 1251 1556 1252
rect 1590 1256 1596 1257
rect 1590 1252 1591 1256
rect 1595 1252 1596 1256
rect 1590 1251 1596 1252
rect 1630 1256 1636 1257
rect 1630 1252 1631 1256
rect 1635 1252 1636 1256
rect 1630 1251 1636 1252
rect 1670 1256 1676 1257
rect 1670 1252 1671 1256
rect 1675 1252 1676 1256
rect 1670 1251 1676 1252
rect 1710 1256 1716 1257
rect 1710 1252 1711 1256
rect 1715 1252 1716 1256
rect 1710 1251 1716 1252
rect 1750 1256 1756 1257
rect 1750 1252 1751 1256
rect 1755 1252 1756 1256
rect 1750 1251 1756 1252
rect 1790 1256 1796 1257
rect 1790 1252 1791 1256
rect 1795 1252 1796 1256
rect 1790 1251 1796 1252
rect 1838 1256 1844 1257
rect 1838 1252 1839 1256
rect 1843 1252 1844 1256
rect 1838 1251 1844 1252
rect 1902 1256 1908 1257
rect 1902 1252 1903 1256
rect 1907 1252 1908 1256
rect 1902 1251 1908 1252
rect 1966 1256 1972 1257
rect 1966 1252 1967 1256
rect 1971 1252 1972 1256
rect 1966 1251 1972 1252
rect 2038 1256 2044 1257
rect 2038 1252 2039 1256
rect 2043 1252 2044 1256
rect 2038 1251 2044 1252
rect 2118 1256 2124 1257
rect 2118 1252 2119 1256
rect 2123 1252 2124 1256
rect 2118 1251 2124 1252
rect 2206 1256 2212 1257
rect 2206 1252 2207 1256
rect 2211 1252 2212 1256
rect 2206 1251 2212 1252
rect 2294 1256 2300 1257
rect 2294 1252 2295 1256
rect 2299 1252 2300 1256
rect 2294 1251 2300 1252
rect 2358 1256 2364 1257
rect 2358 1252 2359 1256
rect 2363 1252 2364 1256
rect 2358 1251 2364 1252
rect 1278 1249 1284 1250
rect 1278 1245 1279 1249
rect 1283 1245 1284 1249
rect 1278 1244 1284 1245
rect 2406 1249 2412 1250
rect 2406 1245 2407 1249
rect 2411 1245 2412 1249
rect 2406 1244 2412 1245
rect 110 1240 116 1241
rect 110 1236 111 1240
rect 115 1236 116 1240
rect 110 1235 116 1236
rect 1238 1240 1244 1241
rect 1238 1236 1239 1240
rect 1243 1236 1244 1240
rect 1238 1235 1244 1236
rect 1278 1232 1284 1233
rect 1278 1228 1279 1232
rect 1283 1228 1284 1232
rect 1278 1227 1284 1228
rect 2406 1232 2412 1233
rect 2406 1228 2407 1232
rect 2411 1228 2412 1232
rect 2406 1227 2412 1228
rect 134 1217 140 1218
rect 134 1213 135 1217
rect 139 1213 140 1217
rect 134 1212 140 1213
rect 174 1217 180 1218
rect 174 1213 175 1217
rect 179 1213 180 1217
rect 174 1212 180 1213
rect 246 1217 252 1218
rect 246 1213 247 1217
rect 251 1213 252 1217
rect 246 1212 252 1213
rect 326 1217 332 1218
rect 326 1213 327 1217
rect 331 1213 332 1217
rect 326 1212 332 1213
rect 414 1217 420 1218
rect 414 1213 415 1217
rect 419 1213 420 1217
rect 414 1212 420 1213
rect 502 1217 508 1218
rect 502 1213 503 1217
rect 507 1213 508 1217
rect 502 1212 508 1213
rect 590 1217 596 1218
rect 590 1213 591 1217
rect 595 1213 596 1217
rect 590 1212 596 1213
rect 670 1217 676 1218
rect 670 1213 671 1217
rect 675 1213 676 1217
rect 670 1212 676 1213
rect 742 1217 748 1218
rect 742 1213 743 1217
rect 747 1213 748 1217
rect 742 1212 748 1213
rect 814 1217 820 1218
rect 814 1213 815 1217
rect 819 1213 820 1217
rect 814 1212 820 1213
rect 878 1217 884 1218
rect 878 1213 879 1217
rect 883 1213 884 1217
rect 878 1212 884 1213
rect 942 1217 948 1218
rect 942 1213 943 1217
rect 947 1213 948 1217
rect 942 1212 948 1213
rect 1006 1217 1012 1218
rect 1006 1213 1007 1217
rect 1011 1213 1012 1217
rect 1006 1212 1012 1213
rect 1070 1217 1076 1218
rect 1070 1213 1071 1217
rect 1075 1213 1076 1217
rect 1070 1212 1076 1213
rect 1510 1209 1516 1210
rect 1510 1205 1511 1209
rect 1515 1205 1516 1209
rect 1510 1204 1516 1205
rect 1550 1209 1556 1210
rect 1550 1205 1551 1209
rect 1555 1205 1556 1209
rect 1550 1204 1556 1205
rect 1590 1209 1596 1210
rect 1590 1205 1591 1209
rect 1595 1205 1596 1209
rect 1590 1204 1596 1205
rect 1630 1209 1636 1210
rect 1630 1205 1631 1209
rect 1635 1205 1636 1209
rect 1630 1204 1636 1205
rect 1670 1209 1676 1210
rect 1670 1205 1671 1209
rect 1675 1205 1676 1209
rect 1670 1204 1676 1205
rect 1710 1209 1716 1210
rect 1710 1205 1711 1209
rect 1715 1205 1716 1209
rect 1710 1204 1716 1205
rect 1750 1209 1756 1210
rect 1750 1205 1751 1209
rect 1755 1205 1756 1209
rect 1750 1204 1756 1205
rect 1790 1209 1796 1210
rect 1790 1205 1791 1209
rect 1795 1205 1796 1209
rect 1790 1204 1796 1205
rect 1838 1209 1844 1210
rect 1838 1205 1839 1209
rect 1843 1205 1844 1209
rect 1838 1204 1844 1205
rect 1902 1209 1908 1210
rect 1902 1205 1903 1209
rect 1907 1205 1908 1209
rect 1902 1204 1908 1205
rect 1966 1209 1972 1210
rect 1966 1205 1967 1209
rect 1971 1205 1972 1209
rect 1966 1204 1972 1205
rect 2038 1209 2044 1210
rect 2038 1205 2039 1209
rect 2043 1205 2044 1209
rect 2038 1204 2044 1205
rect 2118 1209 2124 1210
rect 2118 1205 2119 1209
rect 2123 1205 2124 1209
rect 2118 1204 2124 1205
rect 2206 1209 2212 1210
rect 2206 1205 2207 1209
rect 2211 1205 2212 1209
rect 2206 1204 2212 1205
rect 2294 1209 2300 1210
rect 2294 1205 2295 1209
rect 2299 1205 2300 1209
rect 2294 1204 2300 1205
rect 2358 1209 2364 1210
rect 2358 1205 2359 1209
rect 2363 1205 2364 1209
rect 2358 1204 2364 1205
rect 134 1179 140 1180
rect 134 1175 135 1179
rect 139 1175 140 1179
rect 134 1174 140 1175
rect 174 1179 180 1180
rect 174 1175 175 1179
rect 179 1175 180 1179
rect 174 1174 180 1175
rect 230 1179 236 1180
rect 230 1175 231 1179
rect 235 1175 236 1179
rect 230 1174 236 1175
rect 302 1179 308 1180
rect 302 1175 303 1179
rect 307 1175 308 1179
rect 302 1174 308 1175
rect 382 1179 388 1180
rect 382 1175 383 1179
rect 387 1175 388 1179
rect 382 1174 388 1175
rect 470 1179 476 1180
rect 470 1175 471 1179
rect 475 1175 476 1179
rect 470 1174 476 1175
rect 558 1179 564 1180
rect 558 1175 559 1179
rect 563 1175 564 1179
rect 558 1174 564 1175
rect 638 1179 644 1180
rect 638 1175 639 1179
rect 643 1175 644 1179
rect 638 1174 644 1175
rect 718 1179 724 1180
rect 718 1175 719 1179
rect 723 1175 724 1179
rect 718 1174 724 1175
rect 798 1179 804 1180
rect 798 1175 799 1179
rect 803 1175 804 1179
rect 798 1174 804 1175
rect 870 1179 876 1180
rect 870 1175 871 1179
rect 875 1175 876 1179
rect 870 1174 876 1175
rect 934 1179 940 1180
rect 934 1175 935 1179
rect 939 1175 940 1179
rect 934 1174 940 1175
rect 990 1179 996 1180
rect 990 1175 991 1179
rect 995 1175 996 1179
rect 990 1174 996 1175
rect 1046 1179 1052 1180
rect 1046 1175 1047 1179
rect 1051 1175 1052 1179
rect 1046 1174 1052 1175
rect 1102 1179 1108 1180
rect 1102 1175 1103 1179
rect 1107 1175 1108 1179
rect 1102 1174 1108 1175
rect 1150 1179 1156 1180
rect 1150 1175 1151 1179
rect 1155 1175 1156 1179
rect 1150 1174 1156 1175
rect 1190 1179 1196 1180
rect 1190 1175 1191 1179
rect 1195 1175 1196 1179
rect 1190 1174 1196 1175
rect 1558 1175 1564 1176
rect 1558 1171 1559 1175
rect 1563 1171 1564 1175
rect 1558 1170 1564 1171
rect 1598 1175 1604 1176
rect 1598 1171 1599 1175
rect 1603 1171 1604 1175
rect 1598 1170 1604 1171
rect 1638 1175 1644 1176
rect 1638 1171 1639 1175
rect 1643 1171 1644 1175
rect 1638 1170 1644 1171
rect 1678 1175 1684 1176
rect 1678 1171 1679 1175
rect 1683 1171 1684 1175
rect 1678 1170 1684 1171
rect 1718 1175 1724 1176
rect 1718 1171 1719 1175
rect 1723 1171 1724 1175
rect 1718 1170 1724 1171
rect 1758 1175 1764 1176
rect 1758 1171 1759 1175
rect 1763 1171 1764 1175
rect 1758 1170 1764 1171
rect 1798 1175 1804 1176
rect 1798 1171 1799 1175
rect 1803 1171 1804 1175
rect 1798 1170 1804 1171
rect 1854 1175 1860 1176
rect 1854 1171 1855 1175
rect 1859 1171 1860 1175
rect 1854 1170 1860 1171
rect 1926 1175 1932 1176
rect 1926 1171 1927 1175
rect 1931 1171 1932 1175
rect 1926 1170 1932 1171
rect 2022 1175 2028 1176
rect 2022 1171 2023 1175
rect 2027 1171 2028 1175
rect 2022 1170 2028 1171
rect 2134 1175 2140 1176
rect 2134 1171 2135 1175
rect 2139 1171 2140 1175
rect 2134 1170 2140 1171
rect 2254 1175 2260 1176
rect 2254 1171 2255 1175
rect 2259 1171 2260 1175
rect 2254 1170 2260 1171
rect 2358 1175 2364 1176
rect 2358 1171 2359 1175
rect 2363 1171 2364 1175
rect 2358 1170 2364 1171
rect 110 1156 116 1157
rect 110 1152 111 1156
rect 115 1152 116 1156
rect 110 1151 116 1152
rect 1238 1156 1244 1157
rect 1238 1152 1239 1156
rect 1243 1152 1244 1156
rect 1238 1151 1244 1152
rect 1278 1152 1284 1153
rect 1278 1148 1279 1152
rect 1283 1148 1284 1152
rect 1278 1147 1284 1148
rect 2406 1152 2412 1153
rect 2406 1148 2407 1152
rect 2411 1148 2412 1152
rect 2406 1147 2412 1148
rect 110 1139 116 1140
rect 110 1135 111 1139
rect 115 1135 116 1139
rect 110 1134 116 1135
rect 1238 1139 1244 1140
rect 1238 1135 1239 1139
rect 1243 1135 1244 1139
rect 1238 1134 1244 1135
rect 1278 1135 1284 1136
rect 134 1132 140 1133
rect 134 1128 135 1132
rect 139 1128 140 1132
rect 134 1127 140 1128
rect 174 1132 180 1133
rect 174 1128 175 1132
rect 179 1128 180 1132
rect 174 1127 180 1128
rect 230 1132 236 1133
rect 230 1128 231 1132
rect 235 1128 236 1132
rect 230 1127 236 1128
rect 302 1132 308 1133
rect 302 1128 303 1132
rect 307 1128 308 1132
rect 302 1127 308 1128
rect 382 1132 388 1133
rect 382 1128 383 1132
rect 387 1128 388 1132
rect 382 1127 388 1128
rect 470 1132 476 1133
rect 470 1128 471 1132
rect 475 1128 476 1132
rect 470 1127 476 1128
rect 558 1132 564 1133
rect 558 1128 559 1132
rect 563 1128 564 1132
rect 558 1127 564 1128
rect 638 1132 644 1133
rect 638 1128 639 1132
rect 643 1128 644 1132
rect 638 1127 644 1128
rect 718 1132 724 1133
rect 718 1128 719 1132
rect 723 1128 724 1132
rect 718 1127 724 1128
rect 798 1132 804 1133
rect 798 1128 799 1132
rect 803 1128 804 1132
rect 798 1127 804 1128
rect 870 1132 876 1133
rect 870 1128 871 1132
rect 875 1128 876 1132
rect 870 1127 876 1128
rect 934 1132 940 1133
rect 934 1128 935 1132
rect 939 1128 940 1132
rect 934 1127 940 1128
rect 990 1132 996 1133
rect 990 1128 991 1132
rect 995 1128 996 1132
rect 990 1127 996 1128
rect 1046 1132 1052 1133
rect 1046 1128 1047 1132
rect 1051 1128 1052 1132
rect 1046 1127 1052 1128
rect 1102 1132 1108 1133
rect 1102 1128 1103 1132
rect 1107 1128 1108 1132
rect 1102 1127 1108 1128
rect 1150 1132 1156 1133
rect 1150 1128 1151 1132
rect 1155 1128 1156 1132
rect 1150 1127 1156 1128
rect 1190 1132 1196 1133
rect 1190 1128 1191 1132
rect 1195 1128 1196 1132
rect 1278 1131 1279 1135
rect 1283 1131 1284 1135
rect 1278 1130 1284 1131
rect 2406 1135 2412 1136
rect 2406 1131 2407 1135
rect 2411 1131 2412 1135
rect 2406 1130 2412 1131
rect 1190 1127 1196 1128
rect 1558 1128 1564 1129
rect 1558 1124 1559 1128
rect 1563 1124 1564 1128
rect 1558 1123 1564 1124
rect 1598 1128 1604 1129
rect 1598 1124 1599 1128
rect 1603 1124 1604 1128
rect 1598 1123 1604 1124
rect 1638 1128 1644 1129
rect 1638 1124 1639 1128
rect 1643 1124 1644 1128
rect 1638 1123 1644 1124
rect 1678 1128 1684 1129
rect 1678 1124 1679 1128
rect 1683 1124 1684 1128
rect 1678 1123 1684 1124
rect 1718 1128 1724 1129
rect 1718 1124 1719 1128
rect 1723 1124 1724 1128
rect 1718 1123 1724 1124
rect 1758 1128 1764 1129
rect 1758 1124 1759 1128
rect 1763 1124 1764 1128
rect 1758 1123 1764 1124
rect 1798 1128 1804 1129
rect 1798 1124 1799 1128
rect 1803 1124 1804 1128
rect 1798 1123 1804 1124
rect 1854 1128 1860 1129
rect 1854 1124 1855 1128
rect 1859 1124 1860 1128
rect 1854 1123 1860 1124
rect 1926 1128 1932 1129
rect 1926 1124 1927 1128
rect 1931 1124 1932 1128
rect 1926 1123 1932 1124
rect 2022 1128 2028 1129
rect 2022 1124 2023 1128
rect 2027 1124 2028 1128
rect 2022 1123 2028 1124
rect 2134 1128 2140 1129
rect 2134 1124 2135 1128
rect 2139 1124 2140 1128
rect 2134 1123 2140 1124
rect 2254 1128 2260 1129
rect 2254 1124 2255 1128
rect 2259 1124 2260 1128
rect 2254 1123 2260 1124
rect 2358 1128 2364 1129
rect 2358 1124 2359 1128
rect 2363 1124 2364 1128
rect 2358 1123 2364 1124
rect 134 1120 140 1121
rect 134 1116 135 1120
rect 139 1116 140 1120
rect 134 1115 140 1116
rect 214 1120 220 1121
rect 214 1116 215 1120
rect 219 1116 220 1120
rect 214 1115 220 1116
rect 302 1120 308 1121
rect 302 1116 303 1120
rect 307 1116 308 1120
rect 302 1115 308 1116
rect 390 1120 396 1121
rect 390 1116 391 1120
rect 395 1116 396 1120
rect 390 1115 396 1116
rect 478 1120 484 1121
rect 478 1116 479 1120
rect 483 1116 484 1120
rect 478 1115 484 1116
rect 558 1120 564 1121
rect 558 1116 559 1120
rect 563 1116 564 1120
rect 558 1115 564 1116
rect 638 1120 644 1121
rect 638 1116 639 1120
rect 643 1116 644 1120
rect 638 1115 644 1116
rect 710 1120 716 1121
rect 710 1116 711 1120
rect 715 1116 716 1120
rect 710 1115 716 1116
rect 774 1120 780 1121
rect 774 1116 775 1120
rect 779 1116 780 1120
rect 774 1115 780 1116
rect 838 1120 844 1121
rect 838 1116 839 1120
rect 843 1116 844 1120
rect 838 1115 844 1116
rect 902 1120 908 1121
rect 902 1116 903 1120
rect 907 1116 908 1120
rect 902 1115 908 1116
rect 958 1120 964 1121
rect 958 1116 959 1120
rect 963 1116 964 1120
rect 958 1115 964 1116
rect 1022 1120 1028 1121
rect 1022 1116 1023 1120
rect 1027 1116 1028 1120
rect 1022 1115 1028 1116
rect 1086 1120 1092 1121
rect 1086 1116 1087 1120
rect 1091 1116 1092 1120
rect 1086 1115 1092 1116
rect 1150 1120 1156 1121
rect 1150 1116 1151 1120
rect 1155 1116 1156 1120
rect 1150 1115 1156 1116
rect 1190 1120 1196 1121
rect 1190 1116 1191 1120
rect 1195 1116 1196 1120
rect 1190 1115 1196 1116
rect 110 1113 116 1114
rect 110 1109 111 1113
rect 115 1109 116 1113
rect 110 1108 116 1109
rect 1238 1113 1244 1114
rect 1238 1109 1239 1113
rect 1243 1109 1244 1113
rect 1238 1108 1244 1109
rect 1534 1108 1540 1109
rect 1534 1104 1535 1108
rect 1539 1104 1540 1108
rect 1534 1103 1540 1104
rect 1598 1108 1604 1109
rect 1598 1104 1599 1108
rect 1603 1104 1604 1108
rect 1598 1103 1604 1104
rect 1662 1108 1668 1109
rect 1662 1104 1663 1108
rect 1667 1104 1668 1108
rect 1662 1103 1668 1104
rect 1726 1108 1732 1109
rect 1726 1104 1727 1108
rect 1731 1104 1732 1108
rect 1726 1103 1732 1104
rect 1790 1108 1796 1109
rect 1790 1104 1791 1108
rect 1795 1104 1796 1108
rect 1790 1103 1796 1104
rect 1854 1108 1860 1109
rect 1854 1104 1855 1108
rect 1859 1104 1860 1108
rect 1854 1103 1860 1104
rect 1910 1108 1916 1109
rect 1910 1104 1911 1108
rect 1915 1104 1916 1108
rect 1910 1103 1916 1104
rect 1966 1108 1972 1109
rect 1966 1104 1967 1108
rect 1971 1104 1972 1108
rect 1966 1103 1972 1104
rect 2022 1108 2028 1109
rect 2022 1104 2023 1108
rect 2027 1104 2028 1108
rect 2022 1103 2028 1104
rect 2078 1108 2084 1109
rect 2078 1104 2079 1108
rect 2083 1104 2084 1108
rect 2078 1103 2084 1104
rect 2134 1108 2140 1109
rect 2134 1104 2135 1108
rect 2139 1104 2140 1108
rect 2134 1103 2140 1104
rect 2190 1108 2196 1109
rect 2190 1104 2191 1108
rect 2195 1104 2196 1108
rect 2190 1103 2196 1104
rect 2254 1108 2260 1109
rect 2254 1104 2255 1108
rect 2259 1104 2260 1108
rect 2254 1103 2260 1104
rect 2318 1108 2324 1109
rect 2318 1104 2319 1108
rect 2323 1104 2324 1108
rect 2318 1103 2324 1104
rect 2358 1108 2364 1109
rect 2358 1104 2359 1108
rect 2363 1104 2364 1108
rect 2358 1103 2364 1104
rect 1278 1101 1284 1102
rect 1278 1097 1279 1101
rect 1283 1097 1284 1101
rect 110 1096 116 1097
rect 110 1092 111 1096
rect 115 1092 116 1096
rect 110 1091 116 1092
rect 1238 1096 1244 1097
rect 1278 1096 1284 1097
rect 2406 1101 2412 1102
rect 2406 1097 2407 1101
rect 2411 1097 2412 1101
rect 2406 1096 2412 1097
rect 1238 1092 1239 1096
rect 1243 1092 1244 1096
rect 1238 1091 1244 1092
rect 1278 1084 1284 1085
rect 1278 1080 1279 1084
rect 1283 1080 1284 1084
rect 1278 1079 1284 1080
rect 2406 1084 2412 1085
rect 2406 1080 2407 1084
rect 2411 1080 2412 1084
rect 2406 1079 2412 1080
rect 134 1073 140 1074
rect 134 1069 135 1073
rect 139 1069 140 1073
rect 134 1068 140 1069
rect 214 1073 220 1074
rect 214 1069 215 1073
rect 219 1069 220 1073
rect 214 1068 220 1069
rect 302 1073 308 1074
rect 302 1069 303 1073
rect 307 1069 308 1073
rect 302 1068 308 1069
rect 390 1073 396 1074
rect 390 1069 391 1073
rect 395 1069 396 1073
rect 390 1068 396 1069
rect 478 1073 484 1074
rect 478 1069 479 1073
rect 483 1069 484 1073
rect 478 1068 484 1069
rect 558 1073 564 1074
rect 558 1069 559 1073
rect 563 1069 564 1073
rect 558 1068 564 1069
rect 638 1073 644 1074
rect 638 1069 639 1073
rect 643 1069 644 1073
rect 638 1068 644 1069
rect 710 1073 716 1074
rect 710 1069 711 1073
rect 715 1069 716 1073
rect 710 1068 716 1069
rect 774 1073 780 1074
rect 774 1069 775 1073
rect 779 1069 780 1073
rect 774 1068 780 1069
rect 838 1073 844 1074
rect 838 1069 839 1073
rect 843 1069 844 1073
rect 838 1068 844 1069
rect 902 1073 908 1074
rect 902 1069 903 1073
rect 907 1069 908 1073
rect 902 1068 908 1069
rect 958 1073 964 1074
rect 958 1069 959 1073
rect 963 1069 964 1073
rect 958 1068 964 1069
rect 1022 1073 1028 1074
rect 1022 1069 1023 1073
rect 1027 1069 1028 1073
rect 1022 1068 1028 1069
rect 1086 1073 1092 1074
rect 1086 1069 1087 1073
rect 1091 1069 1092 1073
rect 1086 1068 1092 1069
rect 1150 1073 1156 1074
rect 1150 1069 1151 1073
rect 1155 1069 1156 1073
rect 1150 1068 1156 1069
rect 1190 1073 1196 1074
rect 1190 1069 1191 1073
rect 1195 1069 1196 1073
rect 1190 1068 1196 1069
rect 1534 1061 1540 1062
rect 1534 1057 1535 1061
rect 1539 1057 1540 1061
rect 1534 1056 1540 1057
rect 1598 1061 1604 1062
rect 1598 1057 1599 1061
rect 1603 1057 1604 1061
rect 1598 1056 1604 1057
rect 1662 1061 1668 1062
rect 1662 1057 1663 1061
rect 1667 1057 1668 1061
rect 1662 1056 1668 1057
rect 1726 1061 1732 1062
rect 1726 1057 1727 1061
rect 1731 1057 1732 1061
rect 1726 1056 1732 1057
rect 1790 1061 1796 1062
rect 1790 1057 1791 1061
rect 1795 1057 1796 1061
rect 1790 1056 1796 1057
rect 1854 1061 1860 1062
rect 1854 1057 1855 1061
rect 1859 1057 1860 1061
rect 1854 1056 1860 1057
rect 1910 1061 1916 1062
rect 1910 1057 1911 1061
rect 1915 1057 1916 1061
rect 1910 1056 1916 1057
rect 1966 1061 1972 1062
rect 1966 1057 1967 1061
rect 1971 1057 1972 1061
rect 1966 1056 1972 1057
rect 2022 1061 2028 1062
rect 2022 1057 2023 1061
rect 2027 1057 2028 1061
rect 2022 1056 2028 1057
rect 2078 1061 2084 1062
rect 2078 1057 2079 1061
rect 2083 1057 2084 1061
rect 2078 1056 2084 1057
rect 2134 1061 2140 1062
rect 2134 1057 2135 1061
rect 2139 1057 2140 1061
rect 2134 1056 2140 1057
rect 2190 1061 2196 1062
rect 2190 1057 2191 1061
rect 2195 1057 2196 1061
rect 2190 1056 2196 1057
rect 2254 1061 2260 1062
rect 2254 1057 2255 1061
rect 2259 1057 2260 1061
rect 2254 1056 2260 1057
rect 2318 1061 2324 1062
rect 2318 1057 2319 1061
rect 2323 1057 2324 1061
rect 2318 1056 2324 1057
rect 2358 1061 2364 1062
rect 2358 1057 2359 1061
rect 2363 1057 2364 1061
rect 2358 1056 2364 1057
rect 198 1039 204 1040
rect 198 1035 199 1039
rect 203 1035 204 1039
rect 198 1034 204 1035
rect 238 1039 244 1040
rect 238 1035 239 1039
rect 243 1035 244 1039
rect 238 1034 244 1035
rect 286 1039 292 1040
rect 286 1035 287 1039
rect 291 1035 292 1039
rect 286 1034 292 1035
rect 342 1039 348 1040
rect 342 1035 343 1039
rect 347 1035 348 1039
rect 342 1034 348 1035
rect 390 1039 396 1040
rect 390 1035 391 1039
rect 395 1035 396 1039
rect 390 1034 396 1035
rect 438 1039 444 1040
rect 438 1035 439 1039
rect 443 1035 444 1039
rect 438 1034 444 1035
rect 486 1039 492 1040
rect 486 1035 487 1039
rect 491 1035 492 1039
rect 486 1034 492 1035
rect 534 1039 540 1040
rect 534 1035 535 1039
rect 539 1035 540 1039
rect 534 1034 540 1035
rect 582 1039 588 1040
rect 582 1035 583 1039
rect 587 1035 588 1039
rect 582 1034 588 1035
rect 630 1039 636 1040
rect 630 1035 631 1039
rect 635 1035 636 1039
rect 630 1034 636 1035
rect 678 1039 684 1040
rect 678 1035 679 1039
rect 683 1035 684 1039
rect 678 1034 684 1035
rect 726 1039 732 1040
rect 726 1035 727 1039
rect 731 1035 732 1039
rect 726 1034 732 1035
rect 782 1039 788 1040
rect 782 1035 783 1039
rect 787 1035 788 1039
rect 782 1034 788 1035
rect 838 1039 844 1040
rect 838 1035 839 1039
rect 843 1035 844 1039
rect 838 1034 844 1035
rect 894 1039 900 1040
rect 894 1035 895 1039
rect 899 1035 900 1039
rect 894 1034 900 1035
rect 958 1039 964 1040
rect 958 1035 959 1039
rect 963 1035 964 1039
rect 958 1034 964 1035
rect 1022 1039 1028 1040
rect 1022 1035 1023 1039
rect 1027 1035 1028 1039
rect 1022 1034 1028 1035
rect 1086 1039 1092 1040
rect 1086 1035 1087 1039
rect 1091 1035 1092 1039
rect 1086 1034 1092 1035
rect 1150 1039 1156 1040
rect 1150 1035 1151 1039
rect 1155 1035 1156 1039
rect 1150 1034 1156 1035
rect 1190 1039 1196 1040
rect 1190 1035 1191 1039
rect 1195 1035 1196 1039
rect 1190 1034 1196 1035
rect 1502 1019 1508 1020
rect 110 1016 116 1017
rect 110 1012 111 1016
rect 115 1012 116 1016
rect 110 1011 116 1012
rect 1238 1016 1244 1017
rect 1238 1012 1239 1016
rect 1243 1012 1244 1016
rect 1502 1015 1503 1019
rect 1507 1015 1508 1019
rect 1502 1014 1508 1015
rect 1622 1019 1628 1020
rect 1622 1015 1623 1019
rect 1627 1015 1628 1019
rect 1622 1014 1628 1015
rect 1734 1019 1740 1020
rect 1734 1015 1735 1019
rect 1739 1015 1740 1019
rect 1734 1014 1740 1015
rect 1830 1019 1836 1020
rect 1830 1015 1831 1019
rect 1835 1015 1836 1019
rect 1830 1014 1836 1015
rect 1918 1019 1924 1020
rect 1918 1015 1919 1019
rect 1923 1015 1924 1019
rect 1918 1014 1924 1015
rect 1998 1019 2004 1020
rect 1998 1015 1999 1019
rect 2003 1015 2004 1019
rect 1998 1014 2004 1015
rect 2070 1019 2076 1020
rect 2070 1015 2071 1019
rect 2075 1015 2076 1019
rect 2070 1014 2076 1015
rect 2142 1019 2148 1020
rect 2142 1015 2143 1019
rect 2147 1015 2148 1019
rect 2142 1014 2148 1015
rect 2206 1019 2212 1020
rect 2206 1015 2207 1019
rect 2211 1015 2212 1019
rect 2206 1014 2212 1015
rect 2278 1019 2284 1020
rect 2278 1015 2279 1019
rect 2283 1015 2284 1019
rect 2278 1014 2284 1015
rect 1238 1011 1244 1012
rect 110 999 116 1000
rect 110 995 111 999
rect 115 995 116 999
rect 110 994 116 995
rect 1238 999 1244 1000
rect 1238 995 1239 999
rect 1243 995 1244 999
rect 1238 994 1244 995
rect 1278 996 1284 997
rect 198 992 204 993
rect 198 988 199 992
rect 203 988 204 992
rect 198 987 204 988
rect 238 992 244 993
rect 238 988 239 992
rect 243 988 244 992
rect 238 987 244 988
rect 286 992 292 993
rect 286 988 287 992
rect 291 988 292 992
rect 286 987 292 988
rect 342 992 348 993
rect 342 988 343 992
rect 347 988 348 992
rect 342 987 348 988
rect 390 992 396 993
rect 390 988 391 992
rect 395 988 396 992
rect 390 987 396 988
rect 438 992 444 993
rect 438 988 439 992
rect 443 988 444 992
rect 438 987 444 988
rect 486 992 492 993
rect 486 988 487 992
rect 491 988 492 992
rect 486 987 492 988
rect 534 992 540 993
rect 534 988 535 992
rect 539 988 540 992
rect 534 987 540 988
rect 582 992 588 993
rect 582 988 583 992
rect 587 988 588 992
rect 582 987 588 988
rect 630 992 636 993
rect 630 988 631 992
rect 635 988 636 992
rect 630 987 636 988
rect 678 992 684 993
rect 678 988 679 992
rect 683 988 684 992
rect 678 987 684 988
rect 726 992 732 993
rect 726 988 727 992
rect 731 988 732 992
rect 726 987 732 988
rect 782 992 788 993
rect 782 988 783 992
rect 787 988 788 992
rect 782 987 788 988
rect 838 992 844 993
rect 838 988 839 992
rect 843 988 844 992
rect 838 987 844 988
rect 894 992 900 993
rect 894 988 895 992
rect 899 988 900 992
rect 894 987 900 988
rect 958 992 964 993
rect 958 988 959 992
rect 963 988 964 992
rect 958 987 964 988
rect 1022 992 1028 993
rect 1022 988 1023 992
rect 1027 988 1028 992
rect 1022 987 1028 988
rect 1086 992 1092 993
rect 1086 988 1087 992
rect 1091 988 1092 992
rect 1086 987 1092 988
rect 1150 992 1156 993
rect 1150 988 1151 992
rect 1155 988 1156 992
rect 1150 987 1156 988
rect 1190 992 1196 993
rect 1190 988 1191 992
rect 1195 988 1196 992
rect 1278 992 1279 996
rect 1283 992 1284 996
rect 1278 991 1284 992
rect 2406 996 2412 997
rect 2406 992 2407 996
rect 2411 992 2412 996
rect 2406 991 2412 992
rect 1190 987 1196 988
rect 1278 979 1284 980
rect 1278 975 1279 979
rect 1283 975 1284 979
rect 1278 974 1284 975
rect 2406 979 2412 980
rect 2406 975 2407 979
rect 2411 975 2412 979
rect 2406 974 2412 975
rect 1502 972 1508 973
rect 294 968 300 969
rect 294 964 295 968
rect 299 964 300 968
rect 294 963 300 964
rect 342 968 348 969
rect 342 964 343 968
rect 347 964 348 968
rect 342 963 348 964
rect 398 968 404 969
rect 398 964 399 968
rect 403 964 404 968
rect 398 963 404 964
rect 470 968 476 969
rect 470 964 471 968
rect 475 964 476 968
rect 470 963 476 964
rect 550 968 556 969
rect 550 964 551 968
rect 555 964 556 968
rect 550 963 556 964
rect 638 968 644 969
rect 638 964 639 968
rect 643 964 644 968
rect 638 963 644 964
rect 726 968 732 969
rect 726 964 727 968
rect 731 964 732 968
rect 726 963 732 964
rect 806 968 812 969
rect 806 964 807 968
rect 811 964 812 968
rect 806 963 812 964
rect 886 968 892 969
rect 886 964 887 968
rect 891 964 892 968
rect 886 963 892 964
rect 958 968 964 969
rect 958 964 959 968
rect 963 964 964 968
rect 958 963 964 964
rect 1022 968 1028 969
rect 1022 964 1023 968
rect 1027 964 1028 968
rect 1022 963 1028 964
rect 1086 968 1092 969
rect 1086 964 1087 968
rect 1091 964 1092 968
rect 1086 963 1092 964
rect 1150 968 1156 969
rect 1150 964 1151 968
rect 1155 964 1156 968
rect 1150 963 1156 964
rect 1190 968 1196 969
rect 1190 964 1191 968
rect 1195 964 1196 968
rect 1502 968 1503 972
rect 1507 968 1508 972
rect 1502 967 1508 968
rect 1622 972 1628 973
rect 1622 968 1623 972
rect 1627 968 1628 972
rect 1622 967 1628 968
rect 1734 972 1740 973
rect 1734 968 1735 972
rect 1739 968 1740 972
rect 1734 967 1740 968
rect 1830 972 1836 973
rect 1830 968 1831 972
rect 1835 968 1836 972
rect 1830 967 1836 968
rect 1918 972 1924 973
rect 1918 968 1919 972
rect 1923 968 1924 972
rect 1918 967 1924 968
rect 1998 972 2004 973
rect 1998 968 1999 972
rect 2003 968 2004 972
rect 1998 967 2004 968
rect 2070 972 2076 973
rect 2070 968 2071 972
rect 2075 968 2076 972
rect 2070 967 2076 968
rect 2142 972 2148 973
rect 2142 968 2143 972
rect 2147 968 2148 972
rect 2142 967 2148 968
rect 2206 972 2212 973
rect 2206 968 2207 972
rect 2211 968 2212 972
rect 2206 967 2212 968
rect 2278 972 2284 973
rect 2278 968 2279 972
rect 2283 968 2284 972
rect 2278 967 2284 968
rect 1190 963 1196 964
rect 110 961 116 962
rect 110 957 111 961
rect 115 957 116 961
rect 110 956 116 957
rect 1238 961 1244 962
rect 1238 957 1239 961
rect 1243 957 1244 961
rect 1238 956 1244 957
rect 1318 952 1324 953
rect 1318 948 1319 952
rect 1323 948 1324 952
rect 1318 947 1324 948
rect 1358 952 1364 953
rect 1358 948 1359 952
rect 1363 948 1364 952
rect 1358 947 1364 948
rect 1398 952 1404 953
rect 1398 948 1399 952
rect 1403 948 1404 952
rect 1398 947 1404 948
rect 1462 952 1468 953
rect 1462 948 1463 952
rect 1467 948 1468 952
rect 1462 947 1468 948
rect 1542 952 1548 953
rect 1542 948 1543 952
rect 1547 948 1548 952
rect 1542 947 1548 948
rect 1638 952 1644 953
rect 1638 948 1639 952
rect 1643 948 1644 952
rect 1638 947 1644 948
rect 1734 952 1740 953
rect 1734 948 1735 952
rect 1739 948 1740 952
rect 1734 947 1740 948
rect 1838 952 1844 953
rect 1838 948 1839 952
rect 1843 948 1844 952
rect 1838 947 1844 948
rect 1934 952 1940 953
rect 1934 948 1935 952
rect 1939 948 1940 952
rect 1934 947 1940 948
rect 2022 952 2028 953
rect 2022 948 2023 952
rect 2027 948 2028 952
rect 2022 947 2028 948
rect 2102 952 2108 953
rect 2102 948 2103 952
rect 2107 948 2108 952
rect 2102 947 2108 948
rect 2174 952 2180 953
rect 2174 948 2175 952
rect 2179 948 2180 952
rect 2174 947 2180 948
rect 2238 952 2244 953
rect 2238 948 2239 952
rect 2243 948 2244 952
rect 2238 947 2244 948
rect 2310 952 2316 953
rect 2310 948 2311 952
rect 2315 948 2316 952
rect 2310 947 2316 948
rect 2358 952 2364 953
rect 2358 948 2359 952
rect 2363 948 2364 952
rect 2358 947 2364 948
rect 1278 945 1284 946
rect 110 944 116 945
rect 110 940 111 944
rect 115 940 116 944
rect 110 939 116 940
rect 1238 944 1244 945
rect 1238 940 1239 944
rect 1243 940 1244 944
rect 1278 941 1279 945
rect 1283 941 1284 945
rect 1278 940 1284 941
rect 2406 945 2412 946
rect 2406 941 2407 945
rect 2411 941 2412 945
rect 2406 940 2412 941
rect 1238 939 1244 940
rect 1278 928 1284 929
rect 1278 924 1279 928
rect 1283 924 1284 928
rect 1278 923 1284 924
rect 2406 928 2412 929
rect 2406 924 2407 928
rect 2411 924 2412 928
rect 2406 923 2412 924
rect 294 921 300 922
rect 294 917 295 921
rect 299 917 300 921
rect 294 916 300 917
rect 342 921 348 922
rect 342 917 343 921
rect 347 917 348 921
rect 342 916 348 917
rect 398 921 404 922
rect 398 917 399 921
rect 403 917 404 921
rect 398 916 404 917
rect 470 921 476 922
rect 470 917 471 921
rect 475 917 476 921
rect 470 916 476 917
rect 550 921 556 922
rect 550 917 551 921
rect 555 917 556 921
rect 550 916 556 917
rect 638 921 644 922
rect 638 917 639 921
rect 643 917 644 921
rect 638 916 644 917
rect 726 921 732 922
rect 726 917 727 921
rect 731 917 732 921
rect 726 916 732 917
rect 806 921 812 922
rect 806 917 807 921
rect 811 917 812 921
rect 806 916 812 917
rect 886 921 892 922
rect 886 917 887 921
rect 891 917 892 921
rect 886 916 892 917
rect 958 921 964 922
rect 958 917 959 921
rect 963 917 964 921
rect 958 916 964 917
rect 1022 921 1028 922
rect 1022 917 1023 921
rect 1027 917 1028 921
rect 1022 916 1028 917
rect 1086 921 1092 922
rect 1086 917 1087 921
rect 1091 917 1092 921
rect 1086 916 1092 917
rect 1150 921 1156 922
rect 1150 917 1151 921
rect 1155 917 1156 921
rect 1150 916 1156 917
rect 1190 921 1196 922
rect 1190 917 1191 921
rect 1195 917 1196 921
rect 1190 916 1196 917
rect 1318 905 1324 906
rect 1318 901 1319 905
rect 1323 901 1324 905
rect 1318 900 1324 901
rect 1358 905 1364 906
rect 1358 901 1359 905
rect 1363 901 1364 905
rect 1358 900 1364 901
rect 1398 905 1404 906
rect 1398 901 1399 905
rect 1403 901 1404 905
rect 1398 900 1404 901
rect 1462 905 1468 906
rect 1462 901 1463 905
rect 1467 901 1468 905
rect 1462 900 1468 901
rect 1542 905 1548 906
rect 1542 901 1543 905
rect 1547 901 1548 905
rect 1542 900 1548 901
rect 1638 905 1644 906
rect 1638 901 1639 905
rect 1643 901 1644 905
rect 1638 900 1644 901
rect 1734 905 1740 906
rect 1734 901 1735 905
rect 1739 901 1740 905
rect 1734 900 1740 901
rect 1838 905 1844 906
rect 1838 901 1839 905
rect 1843 901 1844 905
rect 1838 900 1844 901
rect 1934 905 1940 906
rect 1934 901 1935 905
rect 1939 901 1940 905
rect 1934 900 1940 901
rect 2022 905 2028 906
rect 2022 901 2023 905
rect 2027 901 2028 905
rect 2022 900 2028 901
rect 2102 905 2108 906
rect 2102 901 2103 905
rect 2107 901 2108 905
rect 2102 900 2108 901
rect 2174 905 2180 906
rect 2174 901 2175 905
rect 2179 901 2180 905
rect 2174 900 2180 901
rect 2238 905 2244 906
rect 2238 901 2239 905
rect 2243 901 2244 905
rect 2238 900 2244 901
rect 2310 905 2316 906
rect 2310 901 2311 905
rect 2315 901 2316 905
rect 2310 900 2316 901
rect 2358 905 2364 906
rect 2358 901 2359 905
rect 2363 901 2364 905
rect 2358 900 2364 901
rect 254 883 260 884
rect 254 879 255 883
rect 259 879 260 883
rect 254 878 260 879
rect 310 883 316 884
rect 310 879 311 883
rect 315 879 316 883
rect 310 878 316 879
rect 374 883 380 884
rect 374 879 375 883
rect 379 879 380 883
rect 374 878 380 879
rect 454 883 460 884
rect 454 879 455 883
rect 459 879 460 883
rect 454 878 460 879
rect 534 883 540 884
rect 534 879 535 883
rect 539 879 540 883
rect 534 878 540 879
rect 622 883 628 884
rect 622 879 623 883
rect 627 879 628 883
rect 622 878 628 879
rect 710 883 716 884
rect 710 879 711 883
rect 715 879 716 883
rect 710 878 716 879
rect 790 883 796 884
rect 790 879 791 883
rect 795 879 796 883
rect 790 878 796 879
rect 862 883 868 884
rect 862 879 863 883
rect 867 879 868 883
rect 862 878 868 879
rect 934 883 940 884
rect 934 879 935 883
rect 939 879 940 883
rect 934 878 940 879
rect 998 883 1004 884
rect 998 879 999 883
rect 1003 879 1004 883
rect 998 878 1004 879
rect 1054 883 1060 884
rect 1054 879 1055 883
rect 1059 879 1060 883
rect 1054 878 1060 879
rect 1118 883 1124 884
rect 1118 879 1119 883
rect 1123 879 1124 883
rect 1118 878 1124 879
rect 1182 883 1188 884
rect 1182 879 1183 883
rect 1187 879 1188 883
rect 1182 878 1188 879
rect 1334 867 1340 868
rect 1334 863 1335 867
rect 1339 863 1340 867
rect 1334 862 1340 863
rect 1374 867 1380 868
rect 1374 863 1375 867
rect 1379 863 1380 867
rect 1374 862 1380 863
rect 1414 867 1420 868
rect 1414 863 1415 867
rect 1419 863 1420 867
rect 1414 862 1420 863
rect 1470 867 1476 868
rect 1470 863 1471 867
rect 1475 863 1476 867
rect 1470 862 1476 863
rect 1534 867 1540 868
rect 1534 863 1535 867
rect 1539 863 1540 867
rect 1534 862 1540 863
rect 1606 867 1612 868
rect 1606 863 1607 867
rect 1611 863 1612 867
rect 1606 862 1612 863
rect 1678 867 1684 868
rect 1678 863 1679 867
rect 1683 863 1684 867
rect 1678 862 1684 863
rect 1750 867 1756 868
rect 1750 863 1751 867
rect 1755 863 1756 867
rect 1750 862 1756 863
rect 1822 867 1828 868
rect 1822 863 1823 867
rect 1827 863 1828 867
rect 1822 862 1828 863
rect 1894 867 1900 868
rect 1894 863 1895 867
rect 1899 863 1900 867
rect 1894 862 1900 863
rect 1958 867 1964 868
rect 1958 863 1959 867
rect 1963 863 1964 867
rect 1958 862 1964 863
rect 2022 867 2028 868
rect 2022 863 2023 867
rect 2027 863 2028 867
rect 2022 862 2028 863
rect 2086 867 2092 868
rect 2086 863 2087 867
rect 2091 863 2092 867
rect 2086 862 2092 863
rect 2142 867 2148 868
rect 2142 863 2143 867
rect 2147 863 2148 867
rect 2142 862 2148 863
rect 2198 867 2204 868
rect 2198 863 2199 867
rect 2203 863 2204 867
rect 2198 862 2204 863
rect 2254 867 2260 868
rect 2254 863 2255 867
rect 2259 863 2260 867
rect 2254 862 2260 863
rect 2318 867 2324 868
rect 2318 863 2319 867
rect 2323 863 2324 867
rect 2318 862 2324 863
rect 2358 867 2364 868
rect 2358 863 2359 867
rect 2363 863 2364 867
rect 2358 862 2364 863
rect 110 860 116 861
rect 110 856 111 860
rect 115 856 116 860
rect 110 855 116 856
rect 1238 860 1244 861
rect 1238 856 1239 860
rect 1243 856 1244 860
rect 1238 855 1244 856
rect 1278 844 1284 845
rect 110 843 116 844
rect 110 839 111 843
rect 115 839 116 843
rect 110 838 116 839
rect 1238 843 1244 844
rect 1238 839 1239 843
rect 1243 839 1244 843
rect 1278 840 1279 844
rect 1283 840 1284 844
rect 1278 839 1284 840
rect 2406 844 2412 845
rect 2406 840 2407 844
rect 2411 840 2412 844
rect 2406 839 2412 840
rect 1238 838 1244 839
rect 254 836 260 837
rect 254 832 255 836
rect 259 832 260 836
rect 254 831 260 832
rect 310 836 316 837
rect 310 832 311 836
rect 315 832 316 836
rect 310 831 316 832
rect 374 836 380 837
rect 374 832 375 836
rect 379 832 380 836
rect 374 831 380 832
rect 454 836 460 837
rect 454 832 455 836
rect 459 832 460 836
rect 454 831 460 832
rect 534 836 540 837
rect 534 832 535 836
rect 539 832 540 836
rect 534 831 540 832
rect 622 836 628 837
rect 622 832 623 836
rect 627 832 628 836
rect 622 831 628 832
rect 710 836 716 837
rect 710 832 711 836
rect 715 832 716 836
rect 710 831 716 832
rect 790 836 796 837
rect 790 832 791 836
rect 795 832 796 836
rect 790 831 796 832
rect 862 836 868 837
rect 862 832 863 836
rect 867 832 868 836
rect 862 831 868 832
rect 934 836 940 837
rect 934 832 935 836
rect 939 832 940 836
rect 934 831 940 832
rect 998 836 1004 837
rect 998 832 999 836
rect 1003 832 1004 836
rect 998 831 1004 832
rect 1054 836 1060 837
rect 1054 832 1055 836
rect 1059 832 1060 836
rect 1054 831 1060 832
rect 1118 836 1124 837
rect 1118 832 1119 836
rect 1123 832 1124 836
rect 1118 831 1124 832
rect 1182 836 1188 837
rect 1182 832 1183 836
rect 1187 832 1188 836
rect 1182 831 1188 832
rect 1278 827 1284 828
rect 190 824 196 825
rect 190 820 191 824
rect 195 820 196 824
rect 190 819 196 820
rect 246 824 252 825
rect 246 820 247 824
rect 251 820 252 824
rect 246 819 252 820
rect 310 824 316 825
rect 310 820 311 824
rect 315 820 316 824
rect 310 819 316 820
rect 382 824 388 825
rect 382 820 383 824
rect 387 820 388 824
rect 382 819 388 820
rect 462 824 468 825
rect 462 820 463 824
rect 467 820 468 824
rect 462 819 468 820
rect 542 824 548 825
rect 542 820 543 824
rect 547 820 548 824
rect 542 819 548 820
rect 614 824 620 825
rect 614 820 615 824
rect 619 820 620 824
rect 614 819 620 820
rect 686 824 692 825
rect 686 820 687 824
rect 691 820 692 824
rect 686 819 692 820
rect 750 824 756 825
rect 750 820 751 824
rect 755 820 756 824
rect 750 819 756 820
rect 814 824 820 825
rect 814 820 815 824
rect 819 820 820 824
rect 814 819 820 820
rect 870 824 876 825
rect 870 820 871 824
rect 875 820 876 824
rect 870 819 876 820
rect 926 824 932 825
rect 926 820 927 824
rect 931 820 932 824
rect 926 819 932 820
rect 982 824 988 825
rect 982 820 983 824
rect 987 820 988 824
rect 982 819 988 820
rect 1046 824 1052 825
rect 1046 820 1047 824
rect 1051 820 1052 824
rect 1278 823 1279 827
rect 1283 823 1284 827
rect 1278 822 1284 823
rect 2406 827 2412 828
rect 2406 823 2407 827
rect 2411 823 2412 827
rect 2406 822 2412 823
rect 1046 819 1052 820
rect 1334 820 1340 821
rect 110 817 116 818
rect 110 813 111 817
rect 115 813 116 817
rect 110 812 116 813
rect 1238 817 1244 818
rect 1238 813 1239 817
rect 1243 813 1244 817
rect 1334 816 1335 820
rect 1339 816 1340 820
rect 1334 815 1340 816
rect 1374 820 1380 821
rect 1374 816 1375 820
rect 1379 816 1380 820
rect 1374 815 1380 816
rect 1414 820 1420 821
rect 1414 816 1415 820
rect 1419 816 1420 820
rect 1414 815 1420 816
rect 1470 820 1476 821
rect 1470 816 1471 820
rect 1475 816 1476 820
rect 1470 815 1476 816
rect 1534 820 1540 821
rect 1534 816 1535 820
rect 1539 816 1540 820
rect 1534 815 1540 816
rect 1606 820 1612 821
rect 1606 816 1607 820
rect 1611 816 1612 820
rect 1606 815 1612 816
rect 1678 820 1684 821
rect 1678 816 1679 820
rect 1683 816 1684 820
rect 1678 815 1684 816
rect 1750 820 1756 821
rect 1750 816 1751 820
rect 1755 816 1756 820
rect 1750 815 1756 816
rect 1822 820 1828 821
rect 1822 816 1823 820
rect 1827 816 1828 820
rect 1822 815 1828 816
rect 1894 820 1900 821
rect 1894 816 1895 820
rect 1899 816 1900 820
rect 1894 815 1900 816
rect 1958 820 1964 821
rect 1958 816 1959 820
rect 1963 816 1964 820
rect 1958 815 1964 816
rect 2022 820 2028 821
rect 2022 816 2023 820
rect 2027 816 2028 820
rect 2022 815 2028 816
rect 2086 820 2092 821
rect 2086 816 2087 820
rect 2091 816 2092 820
rect 2086 815 2092 816
rect 2142 820 2148 821
rect 2142 816 2143 820
rect 2147 816 2148 820
rect 2142 815 2148 816
rect 2198 820 2204 821
rect 2198 816 2199 820
rect 2203 816 2204 820
rect 2198 815 2204 816
rect 2254 820 2260 821
rect 2254 816 2255 820
rect 2259 816 2260 820
rect 2254 815 2260 816
rect 2318 820 2324 821
rect 2318 816 2319 820
rect 2323 816 2324 820
rect 2318 815 2324 816
rect 2358 820 2364 821
rect 2358 816 2359 820
rect 2363 816 2364 820
rect 2358 815 2364 816
rect 1238 812 1244 813
rect 1302 804 1308 805
rect 110 800 116 801
rect 110 796 111 800
rect 115 796 116 800
rect 110 795 116 796
rect 1238 800 1244 801
rect 1238 796 1239 800
rect 1243 796 1244 800
rect 1302 800 1303 804
rect 1307 800 1308 804
rect 1302 799 1308 800
rect 1342 804 1348 805
rect 1342 800 1343 804
rect 1347 800 1348 804
rect 1342 799 1348 800
rect 1406 804 1412 805
rect 1406 800 1407 804
rect 1411 800 1412 804
rect 1406 799 1412 800
rect 1478 804 1484 805
rect 1478 800 1479 804
rect 1483 800 1484 804
rect 1478 799 1484 800
rect 1550 804 1556 805
rect 1550 800 1551 804
rect 1555 800 1556 804
rect 1550 799 1556 800
rect 1622 804 1628 805
rect 1622 800 1623 804
rect 1627 800 1628 804
rect 1622 799 1628 800
rect 1694 804 1700 805
rect 1694 800 1695 804
rect 1699 800 1700 804
rect 1694 799 1700 800
rect 1758 804 1764 805
rect 1758 800 1759 804
rect 1763 800 1764 804
rect 1758 799 1764 800
rect 1822 804 1828 805
rect 1822 800 1823 804
rect 1827 800 1828 804
rect 1822 799 1828 800
rect 1886 804 1892 805
rect 1886 800 1887 804
rect 1891 800 1892 804
rect 1886 799 1892 800
rect 1950 804 1956 805
rect 1950 800 1951 804
rect 1955 800 1956 804
rect 1950 799 1956 800
rect 2022 804 2028 805
rect 2022 800 2023 804
rect 2027 800 2028 804
rect 2022 799 2028 800
rect 2102 804 2108 805
rect 2102 800 2103 804
rect 2107 800 2108 804
rect 2102 799 2108 800
rect 2190 804 2196 805
rect 2190 800 2191 804
rect 2195 800 2196 804
rect 2190 799 2196 800
rect 2278 804 2284 805
rect 2278 800 2279 804
rect 2283 800 2284 804
rect 2278 799 2284 800
rect 2358 804 2364 805
rect 2358 800 2359 804
rect 2363 800 2364 804
rect 2358 799 2364 800
rect 1238 795 1244 796
rect 1278 797 1284 798
rect 1278 793 1279 797
rect 1283 793 1284 797
rect 1278 792 1284 793
rect 2406 797 2412 798
rect 2406 793 2407 797
rect 2411 793 2412 797
rect 2406 792 2412 793
rect 1278 780 1284 781
rect 190 777 196 778
rect 190 773 191 777
rect 195 773 196 777
rect 190 772 196 773
rect 246 777 252 778
rect 246 773 247 777
rect 251 773 252 777
rect 246 772 252 773
rect 310 777 316 778
rect 310 773 311 777
rect 315 773 316 777
rect 310 772 316 773
rect 382 777 388 778
rect 382 773 383 777
rect 387 773 388 777
rect 382 772 388 773
rect 462 777 468 778
rect 462 773 463 777
rect 467 773 468 777
rect 462 772 468 773
rect 542 777 548 778
rect 542 773 543 777
rect 547 773 548 777
rect 542 772 548 773
rect 614 777 620 778
rect 614 773 615 777
rect 619 773 620 777
rect 614 772 620 773
rect 686 777 692 778
rect 686 773 687 777
rect 691 773 692 777
rect 686 772 692 773
rect 750 777 756 778
rect 750 773 751 777
rect 755 773 756 777
rect 750 772 756 773
rect 814 777 820 778
rect 814 773 815 777
rect 819 773 820 777
rect 814 772 820 773
rect 870 777 876 778
rect 870 773 871 777
rect 875 773 876 777
rect 870 772 876 773
rect 926 777 932 778
rect 926 773 927 777
rect 931 773 932 777
rect 926 772 932 773
rect 982 777 988 778
rect 982 773 983 777
rect 987 773 988 777
rect 982 772 988 773
rect 1046 777 1052 778
rect 1046 773 1047 777
rect 1051 773 1052 777
rect 1278 776 1279 780
rect 1283 776 1284 780
rect 1278 775 1284 776
rect 2406 780 2412 781
rect 2406 776 2407 780
rect 2411 776 2412 780
rect 2406 775 2412 776
rect 1046 772 1052 773
rect 1302 757 1308 758
rect 1302 753 1303 757
rect 1307 753 1308 757
rect 1302 752 1308 753
rect 1342 757 1348 758
rect 1342 753 1343 757
rect 1347 753 1348 757
rect 1342 752 1348 753
rect 1406 757 1412 758
rect 1406 753 1407 757
rect 1411 753 1412 757
rect 1406 752 1412 753
rect 1478 757 1484 758
rect 1478 753 1479 757
rect 1483 753 1484 757
rect 1478 752 1484 753
rect 1550 757 1556 758
rect 1550 753 1551 757
rect 1555 753 1556 757
rect 1550 752 1556 753
rect 1622 757 1628 758
rect 1622 753 1623 757
rect 1627 753 1628 757
rect 1622 752 1628 753
rect 1694 757 1700 758
rect 1694 753 1695 757
rect 1699 753 1700 757
rect 1694 752 1700 753
rect 1758 757 1764 758
rect 1758 753 1759 757
rect 1763 753 1764 757
rect 1758 752 1764 753
rect 1822 757 1828 758
rect 1822 753 1823 757
rect 1827 753 1828 757
rect 1822 752 1828 753
rect 1886 757 1892 758
rect 1886 753 1887 757
rect 1891 753 1892 757
rect 1886 752 1892 753
rect 1950 757 1956 758
rect 1950 753 1951 757
rect 1955 753 1956 757
rect 1950 752 1956 753
rect 2022 757 2028 758
rect 2022 753 2023 757
rect 2027 753 2028 757
rect 2022 752 2028 753
rect 2102 757 2108 758
rect 2102 753 2103 757
rect 2107 753 2108 757
rect 2102 752 2108 753
rect 2190 757 2196 758
rect 2190 753 2191 757
rect 2195 753 2196 757
rect 2190 752 2196 753
rect 2278 757 2284 758
rect 2278 753 2279 757
rect 2283 753 2284 757
rect 2278 752 2284 753
rect 2358 757 2364 758
rect 2358 753 2359 757
rect 2363 753 2364 757
rect 2358 752 2364 753
rect 134 747 140 748
rect 134 743 135 747
rect 139 743 140 747
rect 134 742 140 743
rect 174 747 180 748
rect 174 743 175 747
rect 179 743 180 747
rect 174 742 180 743
rect 214 747 220 748
rect 214 743 215 747
rect 219 743 220 747
rect 214 742 220 743
rect 278 747 284 748
rect 278 743 279 747
rect 283 743 284 747
rect 278 742 284 743
rect 350 747 356 748
rect 350 743 351 747
rect 355 743 356 747
rect 350 742 356 743
rect 422 747 428 748
rect 422 743 423 747
rect 427 743 428 747
rect 422 742 428 743
rect 494 747 500 748
rect 494 743 495 747
rect 499 743 500 747
rect 494 742 500 743
rect 558 747 564 748
rect 558 743 559 747
rect 563 743 564 747
rect 558 742 564 743
rect 622 747 628 748
rect 622 743 623 747
rect 627 743 628 747
rect 622 742 628 743
rect 694 747 700 748
rect 694 743 695 747
rect 699 743 700 747
rect 694 742 700 743
rect 782 747 788 748
rect 782 743 783 747
rect 787 743 788 747
rect 782 742 788 743
rect 878 747 884 748
rect 878 743 879 747
rect 883 743 884 747
rect 878 742 884 743
rect 982 747 988 748
rect 982 743 983 747
rect 987 743 988 747
rect 982 742 988 743
rect 1094 747 1100 748
rect 1094 743 1095 747
rect 1099 743 1100 747
rect 1094 742 1100 743
rect 1190 747 1196 748
rect 1190 743 1191 747
rect 1195 743 1196 747
rect 1190 742 1196 743
rect 1302 727 1308 728
rect 110 724 116 725
rect 110 720 111 724
rect 115 720 116 724
rect 110 719 116 720
rect 1238 724 1244 725
rect 1238 720 1239 724
rect 1243 720 1244 724
rect 1302 723 1303 727
rect 1307 723 1308 727
rect 1302 722 1308 723
rect 1366 727 1372 728
rect 1366 723 1367 727
rect 1371 723 1372 727
rect 1366 722 1372 723
rect 1454 727 1460 728
rect 1454 723 1455 727
rect 1459 723 1460 727
rect 1454 722 1460 723
rect 1534 727 1540 728
rect 1534 723 1535 727
rect 1539 723 1540 727
rect 1534 722 1540 723
rect 1614 727 1620 728
rect 1614 723 1615 727
rect 1619 723 1620 727
rect 1614 722 1620 723
rect 1694 727 1700 728
rect 1694 723 1695 727
rect 1699 723 1700 727
rect 1694 722 1700 723
rect 1774 727 1780 728
rect 1774 723 1775 727
rect 1779 723 1780 727
rect 1774 722 1780 723
rect 1854 727 1860 728
rect 1854 723 1855 727
rect 1859 723 1860 727
rect 1854 722 1860 723
rect 1942 727 1948 728
rect 1942 723 1943 727
rect 1947 723 1948 727
rect 1942 722 1948 723
rect 2030 727 2036 728
rect 2030 723 2031 727
rect 2035 723 2036 727
rect 2030 722 2036 723
rect 2118 727 2124 728
rect 2118 723 2119 727
rect 2123 723 2124 727
rect 2118 722 2124 723
rect 2206 727 2212 728
rect 2206 723 2207 727
rect 2211 723 2212 727
rect 2206 722 2212 723
rect 2294 727 2300 728
rect 2294 723 2295 727
rect 2299 723 2300 727
rect 2294 722 2300 723
rect 2358 727 2364 728
rect 2358 723 2359 727
rect 2363 723 2364 727
rect 2358 722 2364 723
rect 1238 719 1244 720
rect 110 707 116 708
rect 110 703 111 707
rect 115 703 116 707
rect 110 702 116 703
rect 1238 707 1244 708
rect 1238 703 1239 707
rect 1243 703 1244 707
rect 1238 702 1244 703
rect 1278 704 1284 705
rect 134 700 140 701
rect 134 696 135 700
rect 139 696 140 700
rect 134 695 140 696
rect 174 700 180 701
rect 174 696 175 700
rect 179 696 180 700
rect 174 695 180 696
rect 214 700 220 701
rect 214 696 215 700
rect 219 696 220 700
rect 214 695 220 696
rect 278 700 284 701
rect 278 696 279 700
rect 283 696 284 700
rect 278 695 284 696
rect 350 700 356 701
rect 350 696 351 700
rect 355 696 356 700
rect 350 695 356 696
rect 422 700 428 701
rect 422 696 423 700
rect 427 696 428 700
rect 422 695 428 696
rect 494 700 500 701
rect 494 696 495 700
rect 499 696 500 700
rect 494 695 500 696
rect 558 700 564 701
rect 558 696 559 700
rect 563 696 564 700
rect 558 695 564 696
rect 622 700 628 701
rect 622 696 623 700
rect 627 696 628 700
rect 622 695 628 696
rect 694 700 700 701
rect 694 696 695 700
rect 699 696 700 700
rect 694 695 700 696
rect 782 700 788 701
rect 782 696 783 700
rect 787 696 788 700
rect 782 695 788 696
rect 878 700 884 701
rect 878 696 879 700
rect 883 696 884 700
rect 878 695 884 696
rect 982 700 988 701
rect 982 696 983 700
rect 987 696 988 700
rect 982 695 988 696
rect 1094 700 1100 701
rect 1094 696 1095 700
rect 1099 696 1100 700
rect 1094 695 1100 696
rect 1190 700 1196 701
rect 1190 696 1191 700
rect 1195 696 1196 700
rect 1278 700 1279 704
rect 1283 700 1284 704
rect 1278 699 1284 700
rect 2406 704 2412 705
rect 2406 700 2407 704
rect 2411 700 2412 704
rect 2406 699 2412 700
rect 1190 695 1196 696
rect 1278 687 1284 688
rect 1278 683 1279 687
rect 1283 683 1284 687
rect 1278 682 1284 683
rect 2406 687 2412 688
rect 2406 683 2407 687
rect 2411 683 2412 687
rect 2406 682 2412 683
rect 134 680 140 681
rect 134 676 135 680
rect 139 676 140 680
rect 134 675 140 676
rect 174 680 180 681
rect 174 676 175 680
rect 179 676 180 680
rect 174 675 180 676
rect 230 680 236 681
rect 230 676 231 680
rect 235 676 236 680
rect 230 675 236 676
rect 286 680 292 681
rect 286 676 287 680
rect 291 676 292 680
rect 286 675 292 676
rect 342 680 348 681
rect 342 676 343 680
rect 347 676 348 680
rect 342 675 348 676
rect 398 680 404 681
rect 398 676 399 680
rect 403 676 404 680
rect 398 675 404 676
rect 454 680 460 681
rect 454 676 455 680
rect 459 676 460 680
rect 454 675 460 676
rect 502 680 508 681
rect 502 676 503 680
rect 507 676 508 680
rect 502 675 508 676
rect 558 680 564 681
rect 558 676 559 680
rect 563 676 564 680
rect 558 675 564 676
rect 622 680 628 681
rect 622 676 623 680
rect 627 676 628 680
rect 622 675 628 676
rect 694 680 700 681
rect 694 676 695 680
rect 699 676 700 680
rect 694 675 700 676
rect 766 680 772 681
rect 766 676 767 680
rect 771 676 772 680
rect 766 675 772 676
rect 838 680 844 681
rect 838 676 839 680
rect 843 676 844 680
rect 838 675 844 676
rect 902 680 908 681
rect 902 676 903 680
rect 907 676 908 680
rect 902 675 908 676
rect 966 680 972 681
rect 966 676 967 680
rect 971 676 972 680
rect 966 675 972 676
rect 1022 680 1028 681
rect 1022 676 1023 680
rect 1027 676 1028 680
rect 1022 675 1028 676
rect 1086 680 1092 681
rect 1086 676 1087 680
rect 1091 676 1092 680
rect 1086 675 1092 676
rect 1150 680 1156 681
rect 1150 676 1151 680
rect 1155 676 1156 680
rect 1150 675 1156 676
rect 1190 680 1196 681
rect 1190 676 1191 680
rect 1195 676 1196 680
rect 1190 675 1196 676
rect 1302 680 1308 681
rect 1302 676 1303 680
rect 1307 676 1308 680
rect 1302 675 1308 676
rect 1366 680 1372 681
rect 1366 676 1367 680
rect 1371 676 1372 680
rect 1366 675 1372 676
rect 1454 680 1460 681
rect 1454 676 1455 680
rect 1459 676 1460 680
rect 1454 675 1460 676
rect 1534 680 1540 681
rect 1534 676 1535 680
rect 1539 676 1540 680
rect 1534 675 1540 676
rect 1614 680 1620 681
rect 1614 676 1615 680
rect 1619 676 1620 680
rect 1614 675 1620 676
rect 1694 680 1700 681
rect 1694 676 1695 680
rect 1699 676 1700 680
rect 1694 675 1700 676
rect 1774 680 1780 681
rect 1774 676 1775 680
rect 1779 676 1780 680
rect 1774 675 1780 676
rect 1854 680 1860 681
rect 1854 676 1855 680
rect 1859 676 1860 680
rect 1854 675 1860 676
rect 1942 680 1948 681
rect 1942 676 1943 680
rect 1947 676 1948 680
rect 1942 675 1948 676
rect 2030 680 2036 681
rect 2030 676 2031 680
rect 2035 676 2036 680
rect 2030 675 2036 676
rect 2118 680 2124 681
rect 2118 676 2119 680
rect 2123 676 2124 680
rect 2118 675 2124 676
rect 2206 680 2212 681
rect 2206 676 2207 680
rect 2211 676 2212 680
rect 2206 675 2212 676
rect 2294 680 2300 681
rect 2294 676 2295 680
rect 2299 676 2300 680
rect 2294 675 2300 676
rect 2358 680 2364 681
rect 2358 676 2359 680
rect 2363 676 2364 680
rect 2358 675 2364 676
rect 110 673 116 674
rect 110 669 111 673
rect 115 669 116 673
rect 110 668 116 669
rect 1238 673 1244 674
rect 1238 669 1239 673
rect 1243 669 1244 673
rect 1238 668 1244 669
rect 1590 668 1596 669
rect 1590 664 1591 668
rect 1595 664 1596 668
rect 1590 663 1596 664
rect 1638 668 1644 669
rect 1638 664 1639 668
rect 1643 664 1644 668
rect 1638 663 1644 664
rect 1686 668 1692 669
rect 1686 664 1687 668
rect 1691 664 1692 668
rect 1686 663 1692 664
rect 1742 668 1748 669
rect 1742 664 1743 668
rect 1747 664 1748 668
rect 1742 663 1748 664
rect 1798 668 1804 669
rect 1798 664 1799 668
rect 1803 664 1804 668
rect 1798 663 1804 664
rect 1870 668 1876 669
rect 1870 664 1871 668
rect 1875 664 1876 668
rect 1870 663 1876 664
rect 1950 668 1956 669
rect 1950 664 1951 668
rect 1955 664 1956 668
rect 1950 663 1956 664
rect 2046 668 2052 669
rect 2046 664 2047 668
rect 2051 664 2052 668
rect 2046 663 2052 664
rect 2150 668 2156 669
rect 2150 664 2151 668
rect 2155 664 2156 668
rect 2150 663 2156 664
rect 2262 668 2268 669
rect 2262 664 2263 668
rect 2267 664 2268 668
rect 2262 663 2268 664
rect 2358 668 2364 669
rect 2358 664 2359 668
rect 2363 664 2364 668
rect 2358 663 2364 664
rect 1278 661 1284 662
rect 1278 657 1279 661
rect 1283 657 1284 661
rect 110 656 116 657
rect 110 652 111 656
rect 115 652 116 656
rect 110 651 116 652
rect 1238 656 1244 657
rect 1278 656 1284 657
rect 2406 661 2412 662
rect 2406 657 2407 661
rect 2411 657 2412 661
rect 2406 656 2412 657
rect 1238 652 1239 656
rect 1243 652 1244 656
rect 1238 651 1244 652
rect 1278 644 1284 645
rect 1278 640 1279 644
rect 1283 640 1284 644
rect 1278 639 1284 640
rect 2406 644 2412 645
rect 2406 640 2407 644
rect 2411 640 2412 644
rect 2406 639 2412 640
rect 134 633 140 634
rect 134 629 135 633
rect 139 629 140 633
rect 134 628 140 629
rect 174 633 180 634
rect 174 629 175 633
rect 179 629 180 633
rect 174 628 180 629
rect 230 633 236 634
rect 230 629 231 633
rect 235 629 236 633
rect 230 628 236 629
rect 286 633 292 634
rect 286 629 287 633
rect 291 629 292 633
rect 286 628 292 629
rect 342 633 348 634
rect 342 629 343 633
rect 347 629 348 633
rect 342 628 348 629
rect 398 633 404 634
rect 398 629 399 633
rect 403 629 404 633
rect 398 628 404 629
rect 454 633 460 634
rect 454 629 455 633
rect 459 629 460 633
rect 454 628 460 629
rect 502 633 508 634
rect 502 629 503 633
rect 507 629 508 633
rect 502 628 508 629
rect 558 633 564 634
rect 558 629 559 633
rect 563 629 564 633
rect 558 628 564 629
rect 622 633 628 634
rect 622 629 623 633
rect 627 629 628 633
rect 622 628 628 629
rect 694 633 700 634
rect 694 629 695 633
rect 699 629 700 633
rect 694 628 700 629
rect 766 633 772 634
rect 766 629 767 633
rect 771 629 772 633
rect 766 628 772 629
rect 838 633 844 634
rect 838 629 839 633
rect 843 629 844 633
rect 838 628 844 629
rect 902 633 908 634
rect 902 629 903 633
rect 907 629 908 633
rect 902 628 908 629
rect 966 633 972 634
rect 966 629 967 633
rect 971 629 972 633
rect 966 628 972 629
rect 1022 633 1028 634
rect 1022 629 1023 633
rect 1027 629 1028 633
rect 1022 628 1028 629
rect 1086 633 1092 634
rect 1086 629 1087 633
rect 1091 629 1092 633
rect 1086 628 1092 629
rect 1150 633 1156 634
rect 1150 629 1151 633
rect 1155 629 1156 633
rect 1150 628 1156 629
rect 1190 633 1196 634
rect 1190 629 1191 633
rect 1195 629 1196 633
rect 1190 628 1196 629
rect 1590 621 1596 622
rect 1590 617 1591 621
rect 1595 617 1596 621
rect 1590 616 1596 617
rect 1638 621 1644 622
rect 1638 617 1639 621
rect 1643 617 1644 621
rect 1638 616 1644 617
rect 1686 621 1692 622
rect 1686 617 1687 621
rect 1691 617 1692 621
rect 1686 616 1692 617
rect 1742 621 1748 622
rect 1742 617 1743 621
rect 1747 617 1748 621
rect 1742 616 1748 617
rect 1798 621 1804 622
rect 1798 617 1799 621
rect 1803 617 1804 621
rect 1798 616 1804 617
rect 1870 621 1876 622
rect 1870 617 1871 621
rect 1875 617 1876 621
rect 1870 616 1876 617
rect 1950 621 1956 622
rect 1950 617 1951 621
rect 1955 617 1956 621
rect 1950 616 1956 617
rect 2046 621 2052 622
rect 2046 617 2047 621
rect 2051 617 2052 621
rect 2046 616 2052 617
rect 2150 621 2156 622
rect 2150 617 2151 621
rect 2155 617 2156 621
rect 2150 616 2156 617
rect 2262 621 2268 622
rect 2262 617 2263 621
rect 2267 617 2268 621
rect 2262 616 2268 617
rect 2358 621 2364 622
rect 2358 617 2359 621
rect 2363 617 2364 621
rect 2358 616 2364 617
rect 134 603 140 604
rect 134 599 135 603
rect 139 599 140 603
rect 134 598 140 599
rect 182 603 188 604
rect 182 599 183 603
rect 187 599 188 603
rect 182 598 188 599
rect 254 603 260 604
rect 254 599 255 603
rect 259 599 260 603
rect 254 598 260 599
rect 326 603 332 604
rect 326 599 327 603
rect 331 599 332 603
rect 326 598 332 599
rect 398 603 404 604
rect 398 599 399 603
rect 403 599 404 603
rect 398 598 404 599
rect 478 603 484 604
rect 478 599 479 603
rect 483 599 484 603
rect 478 598 484 599
rect 558 603 564 604
rect 558 599 559 603
rect 563 599 564 603
rect 558 598 564 599
rect 638 603 644 604
rect 638 599 639 603
rect 643 599 644 603
rect 638 598 644 599
rect 718 603 724 604
rect 718 599 719 603
rect 723 599 724 603
rect 718 598 724 599
rect 798 603 804 604
rect 798 599 799 603
rect 803 599 804 603
rect 798 598 804 599
rect 878 603 884 604
rect 878 599 879 603
rect 883 599 884 603
rect 878 598 884 599
rect 950 603 956 604
rect 950 599 951 603
rect 955 599 956 603
rect 950 598 956 599
rect 1014 603 1020 604
rect 1014 599 1015 603
rect 1019 599 1020 603
rect 1014 598 1020 599
rect 1078 603 1084 604
rect 1078 599 1079 603
rect 1083 599 1084 603
rect 1078 598 1084 599
rect 1142 603 1148 604
rect 1142 599 1143 603
rect 1147 599 1148 603
rect 1142 598 1148 599
rect 1190 603 1196 604
rect 1190 599 1191 603
rect 1195 599 1196 603
rect 1190 598 1196 599
rect 1558 583 1564 584
rect 110 580 116 581
rect 110 576 111 580
rect 115 576 116 580
rect 110 575 116 576
rect 1238 580 1244 581
rect 1238 576 1239 580
rect 1243 576 1244 580
rect 1558 579 1559 583
rect 1563 579 1564 583
rect 1558 578 1564 579
rect 1598 583 1604 584
rect 1598 579 1599 583
rect 1603 579 1604 583
rect 1598 578 1604 579
rect 1638 583 1644 584
rect 1638 579 1639 583
rect 1643 579 1644 583
rect 1638 578 1644 579
rect 1678 583 1684 584
rect 1678 579 1679 583
rect 1683 579 1684 583
rect 1678 578 1684 579
rect 1718 583 1724 584
rect 1718 579 1719 583
rect 1723 579 1724 583
rect 1718 578 1724 579
rect 1758 583 1764 584
rect 1758 579 1759 583
rect 1763 579 1764 583
rect 1758 578 1764 579
rect 1806 583 1812 584
rect 1806 579 1807 583
rect 1811 579 1812 583
rect 1806 578 1812 579
rect 1854 583 1860 584
rect 1854 579 1855 583
rect 1859 579 1860 583
rect 1854 578 1860 579
rect 1910 583 1916 584
rect 1910 579 1911 583
rect 1915 579 1916 583
rect 1910 578 1916 579
rect 1966 583 1972 584
rect 1966 579 1967 583
rect 1971 579 1972 583
rect 1966 578 1972 579
rect 2030 583 2036 584
rect 2030 579 2031 583
rect 2035 579 2036 583
rect 2030 578 2036 579
rect 2094 583 2100 584
rect 2094 579 2095 583
rect 2099 579 2100 583
rect 2094 578 2100 579
rect 2166 583 2172 584
rect 2166 579 2167 583
rect 2171 579 2172 583
rect 2166 578 2172 579
rect 2238 583 2244 584
rect 2238 579 2239 583
rect 2243 579 2244 583
rect 2238 578 2244 579
rect 2310 583 2316 584
rect 2310 579 2311 583
rect 2315 579 2316 583
rect 2310 578 2316 579
rect 2358 583 2364 584
rect 2358 579 2359 583
rect 2363 579 2364 583
rect 2358 578 2364 579
rect 1238 575 1244 576
rect 110 563 116 564
rect 110 559 111 563
rect 115 559 116 563
rect 110 558 116 559
rect 1238 563 1244 564
rect 1238 559 1239 563
rect 1243 559 1244 563
rect 1238 558 1244 559
rect 1278 560 1284 561
rect 134 556 140 557
rect 134 552 135 556
rect 139 552 140 556
rect 134 551 140 552
rect 182 556 188 557
rect 182 552 183 556
rect 187 552 188 556
rect 182 551 188 552
rect 254 556 260 557
rect 254 552 255 556
rect 259 552 260 556
rect 254 551 260 552
rect 326 556 332 557
rect 326 552 327 556
rect 331 552 332 556
rect 326 551 332 552
rect 398 556 404 557
rect 398 552 399 556
rect 403 552 404 556
rect 398 551 404 552
rect 478 556 484 557
rect 478 552 479 556
rect 483 552 484 556
rect 478 551 484 552
rect 558 556 564 557
rect 558 552 559 556
rect 563 552 564 556
rect 558 551 564 552
rect 638 556 644 557
rect 638 552 639 556
rect 643 552 644 556
rect 638 551 644 552
rect 718 556 724 557
rect 718 552 719 556
rect 723 552 724 556
rect 718 551 724 552
rect 798 556 804 557
rect 798 552 799 556
rect 803 552 804 556
rect 798 551 804 552
rect 878 556 884 557
rect 878 552 879 556
rect 883 552 884 556
rect 878 551 884 552
rect 950 556 956 557
rect 950 552 951 556
rect 955 552 956 556
rect 950 551 956 552
rect 1014 556 1020 557
rect 1014 552 1015 556
rect 1019 552 1020 556
rect 1014 551 1020 552
rect 1078 556 1084 557
rect 1078 552 1079 556
rect 1083 552 1084 556
rect 1078 551 1084 552
rect 1142 556 1148 557
rect 1142 552 1143 556
rect 1147 552 1148 556
rect 1142 551 1148 552
rect 1190 556 1196 557
rect 1190 552 1191 556
rect 1195 552 1196 556
rect 1278 556 1279 560
rect 1283 556 1284 560
rect 1278 555 1284 556
rect 2406 560 2412 561
rect 2406 556 2407 560
rect 2411 556 2412 560
rect 2406 555 2412 556
rect 1190 551 1196 552
rect 1278 543 1284 544
rect 150 540 156 541
rect 150 536 151 540
rect 155 536 156 540
rect 150 535 156 536
rect 222 540 228 541
rect 222 536 223 540
rect 227 536 228 540
rect 222 535 228 536
rect 286 540 292 541
rect 286 536 287 540
rect 291 536 292 540
rect 286 535 292 536
rect 350 540 356 541
rect 350 536 351 540
rect 355 536 356 540
rect 350 535 356 536
rect 414 540 420 541
rect 414 536 415 540
rect 419 536 420 540
rect 414 535 420 536
rect 478 540 484 541
rect 478 536 479 540
rect 483 536 484 540
rect 478 535 484 536
rect 550 540 556 541
rect 550 536 551 540
rect 555 536 556 540
rect 550 535 556 536
rect 622 540 628 541
rect 622 536 623 540
rect 627 536 628 540
rect 622 535 628 536
rect 694 540 700 541
rect 694 536 695 540
rect 699 536 700 540
rect 694 535 700 536
rect 766 540 772 541
rect 766 536 767 540
rect 771 536 772 540
rect 766 535 772 536
rect 838 540 844 541
rect 838 536 839 540
rect 843 536 844 540
rect 838 535 844 536
rect 918 540 924 541
rect 918 536 919 540
rect 923 536 924 540
rect 918 535 924 536
rect 998 540 1004 541
rect 998 536 999 540
rect 1003 536 1004 540
rect 998 535 1004 536
rect 1078 540 1084 541
rect 1078 536 1079 540
rect 1083 536 1084 540
rect 1278 539 1279 543
rect 1283 539 1284 543
rect 1278 538 1284 539
rect 2406 543 2412 544
rect 2406 539 2407 543
rect 2411 539 2412 543
rect 2406 538 2412 539
rect 1078 535 1084 536
rect 1558 536 1564 537
rect 110 533 116 534
rect 110 529 111 533
rect 115 529 116 533
rect 110 528 116 529
rect 1238 533 1244 534
rect 1238 529 1239 533
rect 1243 529 1244 533
rect 1558 532 1559 536
rect 1563 532 1564 536
rect 1558 531 1564 532
rect 1598 536 1604 537
rect 1598 532 1599 536
rect 1603 532 1604 536
rect 1598 531 1604 532
rect 1638 536 1644 537
rect 1638 532 1639 536
rect 1643 532 1644 536
rect 1638 531 1644 532
rect 1678 536 1684 537
rect 1678 532 1679 536
rect 1683 532 1684 536
rect 1678 531 1684 532
rect 1718 536 1724 537
rect 1718 532 1719 536
rect 1723 532 1724 536
rect 1718 531 1724 532
rect 1758 536 1764 537
rect 1758 532 1759 536
rect 1763 532 1764 536
rect 1758 531 1764 532
rect 1806 536 1812 537
rect 1806 532 1807 536
rect 1811 532 1812 536
rect 1806 531 1812 532
rect 1854 536 1860 537
rect 1854 532 1855 536
rect 1859 532 1860 536
rect 1854 531 1860 532
rect 1910 536 1916 537
rect 1910 532 1911 536
rect 1915 532 1916 536
rect 1910 531 1916 532
rect 1966 536 1972 537
rect 1966 532 1967 536
rect 1971 532 1972 536
rect 1966 531 1972 532
rect 2030 536 2036 537
rect 2030 532 2031 536
rect 2035 532 2036 536
rect 2030 531 2036 532
rect 2094 536 2100 537
rect 2094 532 2095 536
rect 2099 532 2100 536
rect 2094 531 2100 532
rect 2166 536 2172 537
rect 2166 532 2167 536
rect 2171 532 2172 536
rect 2166 531 2172 532
rect 2238 536 2244 537
rect 2238 532 2239 536
rect 2243 532 2244 536
rect 2238 531 2244 532
rect 2310 536 2316 537
rect 2310 532 2311 536
rect 2315 532 2316 536
rect 2310 531 2316 532
rect 2358 536 2364 537
rect 2358 532 2359 536
rect 2363 532 2364 536
rect 2358 531 2364 532
rect 1238 528 1244 529
rect 1406 524 1412 525
rect 1406 520 1407 524
rect 1411 520 1412 524
rect 1406 519 1412 520
rect 1446 524 1452 525
rect 1446 520 1447 524
rect 1451 520 1452 524
rect 1446 519 1452 520
rect 1486 524 1492 525
rect 1486 520 1487 524
rect 1491 520 1492 524
rect 1486 519 1492 520
rect 1534 524 1540 525
rect 1534 520 1535 524
rect 1539 520 1540 524
rect 1534 519 1540 520
rect 1590 524 1596 525
rect 1590 520 1591 524
rect 1595 520 1596 524
rect 1590 519 1596 520
rect 1646 524 1652 525
rect 1646 520 1647 524
rect 1651 520 1652 524
rect 1646 519 1652 520
rect 1710 524 1716 525
rect 1710 520 1711 524
rect 1715 520 1716 524
rect 1710 519 1716 520
rect 1782 524 1788 525
rect 1782 520 1783 524
rect 1787 520 1788 524
rect 1782 519 1788 520
rect 1862 524 1868 525
rect 1862 520 1863 524
rect 1867 520 1868 524
rect 1862 519 1868 520
rect 1942 524 1948 525
rect 1942 520 1943 524
rect 1947 520 1948 524
rect 1942 519 1948 520
rect 2022 524 2028 525
rect 2022 520 2023 524
rect 2027 520 2028 524
rect 2022 519 2028 520
rect 2102 524 2108 525
rect 2102 520 2103 524
rect 2107 520 2108 524
rect 2102 519 2108 520
rect 2190 524 2196 525
rect 2190 520 2191 524
rect 2195 520 2196 524
rect 2190 519 2196 520
rect 2286 524 2292 525
rect 2286 520 2287 524
rect 2291 520 2292 524
rect 2286 519 2292 520
rect 2358 524 2364 525
rect 2358 520 2359 524
rect 2363 520 2364 524
rect 2358 519 2364 520
rect 1278 517 1284 518
rect 110 516 116 517
rect 110 512 111 516
rect 115 512 116 516
rect 110 511 116 512
rect 1238 516 1244 517
rect 1238 512 1239 516
rect 1243 512 1244 516
rect 1278 513 1279 517
rect 1283 513 1284 517
rect 1278 512 1284 513
rect 2406 517 2412 518
rect 2406 513 2407 517
rect 2411 513 2412 517
rect 2406 512 2412 513
rect 1238 511 1244 512
rect 1278 500 1284 501
rect 1278 496 1279 500
rect 1283 496 1284 500
rect 1278 495 1284 496
rect 2406 500 2412 501
rect 2406 496 2407 500
rect 2411 496 2412 500
rect 2406 495 2412 496
rect 150 493 156 494
rect 150 489 151 493
rect 155 489 156 493
rect 150 488 156 489
rect 222 493 228 494
rect 222 489 223 493
rect 227 489 228 493
rect 222 488 228 489
rect 286 493 292 494
rect 286 489 287 493
rect 291 489 292 493
rect 286 488 292 489
rect 350 493 356 494
rect 350 489 351 493
rect 355 489 356 493
rect 350 488 356 489
rect 414 493 420 494
rect 414 489 415 493
rect 419 489 420 493
rect 414 488 420 489
rect 478 493 484 494
rect 478 489 479 493
rect 483 489 484 493
rect 478 488 484 489
rect 550 493 556 494
rect 550 489 551 493
rect 555 489 556 493
rect 550 488 556 489
rect 622 493 628 494
rect 622 489 623 493
rect 627 489 628 493
rect 622 488 628 489
rect 694 493 700 494
rect 694 489 695 493
rect 699 489 700 493
rect 694 488 700 489
rect 766 493 772 494
rect 766 489 767 493
rect 771 489 772 493
rect 766 488 772 489
rect 838 493 844 494
rect 838 489 839 493
rect 843 489 844 493
rect 838 488 844 489
rect 918 493 924 494
rect 918 489 919 493
rect 923 489 924 493
rect 918 488 924 489
rect 998 493 1004 494
rect 998 489 999 493
rect 1003 489 1004 493
rect 998 488 1004 489
rect 1078 493 1084 494
rect 1078 489 1079 493
rect 1083 489 1084 493
rect 1078 488 1084 489
rect 1406 477 1412 478
rect 1406 473 1407 477
rect 1411 473 1412 477
rect 1406 472 1412 473
rect 1446 477 1452 478
rect 1446 473 1447 477
rect 1451 473 1452 477
rect 1446 472 1452 473
rect 1486 477 1492 478
rect 1486 473 1487 477
rect 1491 473 1492 477
rect 1486 472 1492 473
rect 1534 477 1540 478
rect 1534 473 1535 477
rect 1539 473 1540 477
rect 1534 472 1540 473
rect 1590 477 1596 478
rect 1590 473 1591 477
rect 1595 473 1596 477
rect 1590 472 1596 473
rect 1646 477 1652 478
rect 1646 473 1647 477
rect 1651 473 1652 477
rect 1646 472 1652 473
rect 1710 477 1716 478
rect 1710 473 1711 477
rect 1715 473 1716 477
rect 1710 472 1716 473
rect 1782 477 1788 478
rect 1782 473 1783 477
rect 1787 473 1788 477
rect 1782 472 1788 473
rect 1862 477 1868 478
rect 1862 473 1863 477
rect 1867 473 1868 477
rect 1862 472 1868 473
rect 1942 477 1948 478
rect 1942 473 1943 477
rect 1947 473 1948 477
rect 1942 472 1948 473
rect 2022 477 2028 478
rect 2022 473 2023 477
rect 2027 473 2028 477
rect 2022 472 2028 473
rect 2102 477 2108 478
rect 2102 473 2103 477
rect 2107 473 2108 477
rect 2102 472 2108 473
rect 2190 477 2196 478
rect 2190 473 2191 477
rect 2195 473 2196 477
rect 2190 472 2196 473
rect 2286 477 2292 478
rect 2286 473 2287 477
rect 2291 473 2292 477
rect 2286 472 2292 473
rect 2358 477 2364 478
rect 2358 473 2359 477
rect 2363 473 2364 477
rect 2358 472 2364 473
rect 238 463 244 464
rect 238 459 239 463
rect 243 459 244 463
rect 238 458 244 459
rect 278 463 284 464
rect 278 459 279 463
rect 283 459 284 463
rect 278 458 284 459
rect 326 463 332 464
rect 326 459 327 463
rect 331 459 332 463
rect 326 458 332 459
rect 382 463 388 464
rect 382 459 383 463
rect 387 459 388 463
rect 382 458 388 459
rect 438 463 444 464
rect 438 459 439 463
rect 443 459 444 463
rect 438 458 444 459
rect 502 463 508 464
rect 502 459 503 463
rect 507 459 508 463
rect 502 458 508 459
rect 566 463 572 464
rect 566 459 567 463
rect 571 459 572 463
rect 566 458 572 459
rect 630 463 636 464
rect 630 459 631 463
rect 635 459 636 463
rect 630 458 636 459
rect 694 463 700 464
rect 694 459 695 463
rect 699 459 700 463
rect 694 458 700 459
rect 758 463 764 464
rect 758 459 759 463
rect 763 459 764 463
rect 758 458 764 459
rect 822 463 828 464
rect 822 459 823 463
rect 827 459 828 463
rect 822 458 828 459
rect 886 463 892 464
rect 886 459 887 463
rect 891 459 892 463
rect 886 458 892 459
rect 950 463 956 464
rect 950 459 951 463
rect 955 459 956 463
rect 950 458 956 459
rect 1014 463 1020 464
rect 1014 459 1015 463
rect 1019 459 1020 463
rect 1014 458 1020 459
rect 1302 447 1308 448
rect 1302 443 1303 447
rect 1307 443 1308 447
rect 1302 442 1308 443
rect 1342 447 1348 448
rect 1342 443 1343 447
rect 1347 443 1348 447
rect 1342 442 1348 443
rect 1382 447 1388 448
rect 1382 443 1383 447
rect 1387 443 1388 447
rect 1382 442 1388 443
rect 1446 447 1452 448
rect 1446 443 1447 447
rect 1451 443 1452 447
rect 1446 442 1452 443
rect 1534 447 1540 448
rect 1534 443 1535 447
rect 1539 443 1540 447
rect 1534 442 1540 443
rect 1630 447 1636 448
rect 1630 443 1631 447
rect 1635 443 1636 447
rect 1630 442 1636 443
rect 1734 447 1740 448
rect 1734 443 1735 447
rect 1739 443 1740 447
rect 1734 442 1740 443
rect 1830 447 1836 448
rect 1830 443 1831 447
rect 1835 443 1836 447
rect 1830 442 1836 443
rect 1918 447 1924 448
rect 1918 443 1919 447
rect 1923 443 1924 447
rect 1918 442 1924 443
rect 1998 447 2004 448
rect 1998 443 1999 447
rect 2003 443 2004 447
rect 1998 442 2004 443
rect 2070 447 2076 448
rect 2070 443 2071 447
rect 2075 443 2076 447
rect 2070 442 2076 443
rect 2134 447 2140 448
rect 2134 443 2135 447
rect 2139 443 2140 447
rect 2134 442 2140 443
rect 2198 447 2204 448
rect 2198 443 2199 447
rect 2203 443 2204 447
rect 2198 442 2204 443
rect 2254 447 2260 448
rect 2254 443 2255 447
rect 2259 443 2260 447
rect 2254 442 2260 443
rect 2318 447 2324 448
rect 2318 443 2319 447
rect 2323 443 2324 447
rect 2318 442 2324 443
rect 2358 447 2364 448
rect 2358 443 2359 447
rect 2363 443 2364 447
rect 2358 442 2364 443
rect 110 440 116 441
rect 110 436 111 440
rect 115 436 116 440
rect 110 435 116 436
rect 1238 440 1244 441
rect 1238 436 1239 440
rect 1243 436 1244 440
rect 1238 435 1244 436
rect 1278 424 1284 425
rect 110 423 116 424
rect 110 419 111 423
rect 115 419 116 423
rect 110 418 116 419
rect 1238 423 1244 424
rect 1238 419 1239 423
rect 1243 419 1244 423
rect 1278 420 1279 424
rect 1283 420 1284 424
rect 1278 419 1284 420
rect 2406 424 2412 425
rect 2406 420 2407 424
rect 2411 420 2412 424
rect 2406 419 2412 420
rect 1238 418 1244 419
rect 238 416 244 417
rect 238 412 239 416
rect 243 412 244 416
rect 238 411 244 412
rect 278 416 284 417
rect 278 412 279 416
rect 283 412 284 416
rect 278 411 284 412
rect 326 416 332 417
rect 326 412 327 416
rect 331 412 332 416
rect 326 411 332 412
rect 382 416 388 417
rect 382 412 383 416
rect 387 412 388 416
rect 382 411 388 412
rect 438 416 444 417
rect 438 412 439 416
rect 443 412 444 416
rect 438 411 444 412
rect 502 416 508 417
rect 502 412 503 416
rect 507 412 508 416
rect 502 411 508 412
rect 566 416 572 417
rect 566 412 567 416
rect 571 412 572 416
rect 566 411 572 412
rect 630 416 636 417
rect 630 412 631 416
rect 635 412 636 416
rect 630 411 636 412
rect 694 416 700 417
rect 694 412 695 416
rect 699 412 700 416
rect 694 411 700 412
rect 758 416 764 417
rect 758 412 759 416
rect 763 412 764 416
rect 758 411 764 412
rect 822 416 828 417
rect 822 412 823 416
rect 827 412 828 416
rect 822 411 828 412
rect 886 416 892 417
rect 886 412 887 416
rect 891 412 892 416
rect 886 411 892 412
rect 950 416 956 417
rect 950 412 951 416
rect 955 412 956 416
rect 950 411 956 412
rect 1014 416 1020 417
rect 1014 412 1015 416
rect 1019 412 1020 416
rect 1014 411 1020 412
rect 1278 407 1284 408
rect 1278 403 1279 407
rect 1283 403 1284 407
rect 1278 402 1284 403
rect 2406 407 2412 408
rect 2406 403 2407 407
rect 2411 403 2412 407
rect 2406 402 2412 403
rect 142 400 148 401
rect 142 396 143 400
rect 147 396 148 400
rect 142 395 148 396
rect 182 400 188 401
rect 182 396 183 400
rect 187 396 188 400
rect 182 395 188 396
rect 222 400 228 401
rect 222 396 223 400
rect 227 396 228 400
rect 222 395 228 396
rect 270 400 276 401
rect 270 396 271 400
rect 275 396 276 400
rect 270 395 276 396
rect 334 400 340 401
rect 334 396 335 400
rect 339 396 340 400
rect 334 395 340 396
rect 398 400 404 401
rect 398 396 399 400
rect 403 396 404 400
rect 398 395 404 396
rect 470 400 476 401
rect 470 396 471 400
rect 475 396 476 400
rect 470 395 476 396
rect 542 400 548 401
rect 542 396 543 400
rect 547 396 548 400
rect 542 395 548 396
rect 614 400 620 401
rect 614 396 615 400
rect 619 396 620 400
rect 614 395 620 396
rect 686 400 692 401
rect 686 396 687 400
rect 691 396 692 400
rect 686 395 692 396
rect 750 400 756 401
rect 750 396 751 400
rect 755 396 756 400
rect 750 395 756 396
rect 806 400 812 401
rect 806 396 807 400
rect 811 396 812 400
rect 806 395 812 396
rect 862 400 868 401
rect 862 396 863 400
rect 867 396 868 400
rect 862 395 868 396
rect 918 400 924 401
rect 918 396 919 400
rect 923 396 924 400
rect 918 395 924 396
rect 974 400 980 401
rect 974 396 975 400
rect 979 396 980 400
rect 974 395 980 396
rect 1030 400 1036 401
rect 1030 396 1031 400
rect 1035 396 1036 400
rect 1030 395 1036 396
rect 1302 400 1308 401
rect 1302 396 1303 400
rect 1307 396 1308 400
rect 1302 395 1308 396
rect 1342 400 1348 401
rect 1342 396 1343 400
rect 1347 396 1348 400
rect 1342 395 1348 396
rect 1382 400 1388 401
rect 1382 396 1383 400
rect 1387 396 1388 400
rect 1382 395 1388 396
rect 1446 400 1452 401
rect 1446 396 1447 400
rect 1451 396 1452 400
rect 1446 395 1452 396
rect 1534 400 1540 401
rect 1534 396 1535 400
rect 1539 396 1540 400
rect 1534 395 1540 396
rect 1630 400 1636 401
rect 1630 396 1631 400
rect 1635 396 1636 400
rect 1630 395 1636 396
rect 1734 400 1740 401
rect 1734 396 1735 400
rect 1739 396 1740 400
rect 1734 395 1740 396
rect 1830 400 1836 401
rect 1830 396 1831 400
rect 1835 396 1836 400
rect 1830 395 1836 396
rect 1918 400 1924 401
rect 1918 396 1919 400
rect 1923 396 1924 400
rect 1918 395 1924 396
rect 1998 400 2004 401
rect 1998 396 1999 400
rect 2003 396 2004 400
rect 1998 395 2004 396
rect 2070 400 2076 401
rect 2070 396 2071 400
rect 2075 396 2076 400
rect 2070 395 2076 396
rect 2134 400 2140 401
rect 2134 396 2135 400
rect 2139 396 2140 400
rect 2134 395 2140 396
rect 2198 400 2204 401
rect 2198 396 2199 400
rect 2203 396 2204 400
rect 2198 395 2204 396
rect 2254 400 2260 401
rect 2254 396 2255 400
rect 2259 396 2260 400
rect 2254 395 2260 396
rect 2318 400 2324 401
rect 2318 396 2319 400
rect 2323 396 2324 400
rect 2318 395 2324 396
rect 2358 400 2364 401
rect 2358 396 2359 400
rect 2363 396 2364 400
rect 2358 395 2364 396
rect 110 393 116 394
rect 110 389 111 393
rect 115 389 116 393
rect 110 388 116 389
rect 1238 393 1244 394
rect 1238 389 1239 393
rect 1243 389 1244 393
rect 1238 388 1244 389
rect 1358 388 1364 389
rect 1358 384 1359 388
rect 1363 384 1364 388
rect 1358 383 1364 384
rect 1398 388 1404 389
rect 1398 384 1399 388
rect 1403 384 1404 388
rect 1398 383 1404 384
rect 1438 388 1444 389
rect 1438 384 1439 388
rect 1443 384 1444 388
rect 1438 383 1444 384
rect 1486 388 1492 389
rect 1486 384 1487 388
rect 1491 384 1492 388
rect 1486 383 1492 384
rect 1542 388 1548 389
rect 1542 384 1543 388
rect 1547 384 1548 388
rect 1542 383 1548 384
rect 1606 388 1612 389
rect 1606 384 1607 388
rect 1611 384 1612 388
rect 1606 383 1612 384
rect 1678 388 1684 389
rect 1678 384 1679 388
rect 1683 384 1684 388
rect 1678 383 1684 384
rect 1758 388 1764 389
rect 1758 384 1759 388
rect 1763 384 1764 388
rect 1758 383 1764 384
rect 1838 388 1844 389
rect 1838 384 1839 388
rect 1843 384 1844 388
rect 1838 383 1844 384
rect 1918 388 1924 389
rect 1918 384 1919 388
rect 1923 384 1924 388
rect 1918 383 1924 384
rect 1998 388 2004 389
rect 1998 384 1999 388
rect 2003 384 2004 388
rect 1998 383 2004 384
rect 2078 388 2084 389
rect 2078 384 2079 388
rect 2083 384 2084 388
rect 2078 383 2084 384
rect 2158 388 2164 389
rect 2158 384 2159 388
rect 2163 384 2164 388
rect 2158 383 2164 384
rect 2246 388 2252 389
rect 2246 384 2247 388
rect 2251 384 2252 388
rect 2246 383 2252 384
rect 2334 388 2340 389
rect 2334 384 2335 388
rect 2339 384 2340 388
rect 2334 383 2340 384
rect 1278 381 1284 382
rect 1278 377 1279 381
rect 1283 377 1284 381
rect 110 376 116 377
rect 110 372 111 376
rect 115 372 116 376
rect 110 371 116 372
rect 1238 376 1244 377
rect 1278 376 1284 377
rect 2406 381 2412 382
rect 2406 377 2407 381
rect 2411 377 2412 381
rect 2406 376 2412 377
rect 1238 372 1239 376
rect 1243 372 1244 376
rect 1238 371 1244 372
rect 1278 364 1284 365
rect 1278 360 1279 364
rect 1283 360 1284 364
rect 1278 359 1284 360
rect 2406 364 2412 365
rect 2406 360 2407 364
rect 2411 360 2412 364
rect 2406 359 2412 360
rect 142 353 148 354
rect 142 349 143 353
rect 147 349 148 353
rect 142 348 148 349
rect 182 353 188 354
rect 182 349 183 353
rect 187 349 188 353
rect 182 348 188 349
rect 222 353 228 354
rect 222 349 223 353
rect 227 349 228 353
rect 222 348 228 349
rect 270 353 276 354
rect 270 349 271 353
rect 275 349 276 353
rect 270 348 276 349
rect 334 353 340 354
rect 334 349 335 353
rect 339 349 340 353
rect 334 348 340 349
rect 398 353 404 354
rect 398 349 399 353
rect 403 349 404 353
rect 398 348 404 349
rect 470 353 476 354
rect 470 349 471 353
rect 475 349 476 353
rect 470 348 476 349
rect 542 353 548 354
rect 542 349 543 353
rect 547 349 548 353
rect 542 348 548 349
rect 614 353 620 354
rect 614 349 615 353
rect 619 349 620 353
rect 614 348 620 349
rect 686 353 692 354
rect 686 349 687 353
rect 691 349 692 353
rect 686 348 692 349
rect 750 353 756 354
rect 750 349 751 353
rect 755 349 756 353
rect 750 348 756 349
rect 806 353 812 354
rect 806 349 807 353
rect 811 349 812 353
rect 806 348 812 349
rect 862 353 868 354
rect 862 349 863 353
rect 867 349 868 353
rect 862 348 868 349
rect 918 353 924 354
rect 918 349 919 353
rect 923 349 924 353
rect 918 348 924 349
rect 974 353 980 354
rect 974 349 975 353
rect 979 349 980 353
rect 974 348 980 349
rect 1030 353 1036 354
rect 1030 349 1031 353
rect 1035 349 1036 353
rect 1030 348 1036 349
rect 1358 341 1364 342
rect 1358 337 1359 341
rect 1363 337 1364 341
rect 1358 336 1364 337
rect 1398 341 1404 342
rect 1398 337 1399 341
rect 1403 337 1404 341
rect 1398 336 1404 337
rect 1438 341 1444 342
rect 1438 337 1439 341
rect 1443 337 1444 341
rect 1438 336 1444 337
rect 1486 341 1492 342
rect 1486 337 1487 341
rect 1491 337 1492 341
rect 1486 336 1492 337
rect 1542 341 1548 342
rect 1542 337 1543 341
rect 1547 337 1548 341
rect 1542 336 1548 337
rect 1606 341 1612 342
rect 1606 337 1607 341
rect 1611 337 1612 341
rect 1606 336 1612 337
rect 1678 341 1684 342
rect 1678 337 1679 341
rect 1683 337 1684 341
rect 1678 336 1684 337
rect 1758 341 1764 342
rect 1758 337 1759 341
rect 1763 337 1764 341
rect 1758 336 1764 337
rect 1838 341 1844 342
rect 1838 337 1839 341
rect 1843 337 1844 341
rect 1838 336 1844 337
rect 1918 341 1924 342
rect 1918 337 1919 341
rect 1923 337 1924 341
rect 1918 336 1924 337
rect 1998 341 2004 342
rect 1998 337 1999 341
rect 2003 337 2004 341
rect 1998 336 2004 337
rect 2078 341 2084 342
rect 2078 337 2079 341
rect 2083 337 2084 341
rect 2078 336 2084 337
rect 2158 341 2164 342
rect 2158 337 2159 341
rect 2163 337 2164 341
rect 2158 336 2164 337
rect 2246 341 2252 342
rect 2246 337 2247 341
rect 2251 337 2252 341
rect 2246 336 2252 337
rect 2334 341 2340 342
rect 2334 337 2335 341
rect 2339 337 2340 341
rect 2334 336 2340 337
rect 134 315 140 316
rect 134 311 135 315
rect 139 311 140 315
rect 134 310 140 311
rect 174 315 180 316
rect 174 311 175 315
rect 179 311 180 315
rect 174 310 180 311
rect 214 315 220 316
rect 214 311 215 315
rect 219 311 220 315
rect 214 310 220 311
rect 254 315 260 316
rect 254 311 255 315
rect 259 311 260 315
rect 254 310 260 311
rect 294 315 300 316
rect 294 311 295 315
rect 299 311 300 315
rect 294 310 300 311
rect 334 315 340 316
rect 334 311 335 315
rect 339 311 340 315
rect 334 310 340 311
rect 390 315 396 316
rect 390 311 391 315
rect 395 311 396 315
rect 390 310 396 311
rect 446 315 452 316
rect 446 311 447 315
rect 451 311 452 315
rect 446 310 452 311
rect 494 315 500 316
rect 494 311 495 315
rect 499 311 500 315
rect 494 310 500 311
rect 542 315 548 316
rect 542 311 543 315
rect 547 311 548 315
rect 542 310 548 311
rect 590 315 596 316
rect 590 311 591 315
rect 595 311 596 315
rect 590 310 596 311
rect 638 315 644 316
rect 638 311 639 315
rect 643 311 644 315
rect 638 310 644 311
rect 686 315 692 316
rect 686 311 687 315
rect 691 311 692 315
rect 686 310 692 311
rect 734 315 740 316
rect 734 311 735 315
rect 739 311 740 315
rect 734 310 740 311
rect 782 315 788 316
rect 782 311 783 315
rect 787 311 788 315
rect 782 310 788 311
rect 838 315 844 316
rect 838 311 839 315
rect 843 311 844 315
rect 838 310 844 311
rect 1510 303 1516 304
rect 1510 299 1511 303
rect 1515 299 1516 303
rect 1510 298 1516 299
rect 1550 303 1556 304
rect 1550 299 1551 303
rect 1555 299 1556 303
rect 1550 298 1556 299
rect 1590 303 1596 304
rect 1590 299 1591 303
rect 1595 299 1596 303
rect 1590 298 1596 299
rect 1630 303 1636 304
rect 1630 299 1631 303
rect 1635 299 1636 303
rect 1630 298 1636 299
rect 1670 303 1676 304
rect 1670 299 1671 303
rect 1675 299 1676 303
rect 1670 298 1676 299
rect 1710 303 1716 304
rect 1710 299 1711 303
rect 1715 299 1716 303
rect 1710 298 1716 299
rect 1750 303 1756 304
rect 1750 299 1751 303
rect 1755 299 1756 303
rect 1750 298 1756 299
rect 1790 303 1796 304
rect 1790 299 1791 303
rect 1795 299 1796 303
rect 1790 298 1796 299
rect 1838 303 1844 304
rect 1838 299 1839 303
rect 1843 299 1844 303
rect 1838 298 1844 299
rect 1902 303 1908 304
rect 1902 299 1903 303
rect 1907 299 1908 303
rect 1902 298 1908 299
rect 1966 303 1972 304
rect 1966 299 1967 303
rect 1971 299 1972 303
rect 1966 298 1972 299
rect 2038 303 2044 304
rect 2038 299 2039 303
rect 2043 299 2044 303
rect 2038 298 2044 299
rect 2118 303 2124 304
rect 2118 299 2119 303
rect 2123 299 2124 303
rect 2118 298 2124 299
rect 2198 303 2204 304
rect 2198 299 2199 303
rect 2203 299 2204 303
rect 2198 298 2204 299
rect 2278 303 2284 304
rect 2278 299 2279 303
rect 2283 299 2284 303
rect 2278 298 2284 299
rect 2358 303 2364 304
rect 2358 299 2359 303
rect 2363 299 2364 303
rect 2358 298 2364 299
rect 110 292 116 293
rect 110 288 111 292
rect 115 288 116 292
rect 110 287 116 288
rect 1238 292 1244 293
rect 1238 288 1239 292
rect 1243 288 1244 292
rect 1238 287 1244 288
rect 1278 280 1284 281
rect 1278 276 1279 280
rect 1283 276 1284 280
rect 110 275 116 276
rect 110 271 111 275
rect 115 271 116 275
rect 110 270 116 271
rect 1238 275 1244 276
rect 1278 275 1284 276
rect 2406 280 2412 281
rect 2406 276 2407 280
rect 2411 276 2412 280
rect 2406 275 2412 276
rect 1238 271 1239 275
rect 1243 271 1244 275
rect 1238 270 1244 271
rect 134 268 140 269
rect 134 264 135 268
rect 139 264 140 268
rect 134 263 140 264
rect 174 268 180 269
rect 174 264 175 268
rect 179 264 180 268
rect 174 263 180 264
rect 214 268 220 269
rect 214 264 215 268
rect 219 264 220 268
rect 214 263 220 264
rect 254 268 260 269
rect 254 264 255 268
rect 259 264 260 268
rect 254 263 260 264
rect 294 268 300 269
rect 294 264 295 268
rect 299 264 300 268
rect 294 263 300 264
rect 334 268 340 269
rect 334 264 335 268
rect 339 264 340 268
rect 334 263 340 264
rect 390 268 396 269
rect 390 264 391 268
rect 395 264 396 268
rect 390 263 396 264
rect 446 268 452 269
rect 446 264 447 268
rect 451 264 452 268
rect 446 263 452 264
rect 494 268 500 269
rect 494 264 495 268
rect 499 264 500 268
rect 494 263 500 264
rect 542 268 548 269
rect 542 264 543 268
rect 547 264 548 268
rect 542 263 548 264
rect 590 268 596 269
rect 590 264 591 268
rect 595 264 596 268
rect 590 263 596 264
rect 638 268 644 269
rect 638 264 639 268
rect 643 264 644 268
rect 638 263 644 264
rect 686 268 692 269
rect 686 264 687 268
rect 691 264 692 268
rect 686 263 692 264
rect 734 268 740 269
rect 734 264 735 268
rect 739 264 740 268
rect 734 263 740 264
rect 782 268 788 269
rect 782 264 783 268
rect 787 264 788 268
rect 782 263 788 264
rect 838 268 844 269
rect 838 264 839 268
rect 843 264 844 268
rect 838 263 844 264
rect 1278 263 1284 264
rect 1278 259 1279 263
rect 1283 259 1284 263
rect 1278 258 1284 259
rect 2406 263 2412 264
rect 2406 259 2407 263
rect 2411 259 2412 263
rect 2406 258 2412 259
rect 1510 256 1516 257
rect 1510 252 1511 256
rect 1515 252 1516 256
rect 1510 251 1516 252
rect 1550 256 1556 257
rect 1550 252 1551 256
rect 1555 252 1556 256
rect 1550 251 1556 252
rect 1590 256 1596 257
rect 1590 252 1591 256
rect 1595 252 1596 256
rect 1590 251 1596 252
rect 1630 256 1636 257
rect 1630 252 1631 256
rect 1635 252 1636 256
rect 1630 251 1636 252
rect 1670 256 1676 257
rect 1670 252 1671 256
rect 1675 252 1676 256
rect 1670 251 1676 252
rect 1710 256 1716 257
rect 1710 252 1711 256
rect 1715 252 1716 256
rect 1710 251 1716 252
rect 1750 256 1756 257
rect 1750 252 1751 256
rect 1755 252 1756 256
rect 1750 251 1756 252
rect 1790 256 1796 257
rect 1790 252 1791 256
rect 1795 252 1796 256
rect 1790 251 1796 252
rect 1838 256 1844 257
rect 1838 252 1839 256
rect 1843 252 1844 256
rect 1838 251 1844 252
rect 1902 256 1908 257
rect 1902 252 1903 256
rect 1907 252 1908 256
rect 1902 251 1908 252
rect 1966 256 1972 257
rect 1966 252 1967 256
rect 1971 252 1972 256
rect 1966 251 1972 252
rect 2038 256 2044 257
rect 2038 252 2039 256
rect 2043 252 2044 256
rect 2038 251 2044 252
rect 2118 256 2124 257
rect 2118 252 2119 256
rect 2123 252 2124 256
rect 2118 251 2124 252
rect 2198 256 2204 257
rect 2198 252 2199 256
rect 2203 252 2204 256
rect 2198 251 2204 252
rect 2278 256 2284 257
rect 2278 252 2279 256
rect 2283 252 2284 256
rect 2278 251 2284 252
rect 2358 256 2364 257
rect 2358 252 2359 256
rect 2363 252 2364 256
rect 2358 251 2364 252
rect 134 248 140 249
rect 134 244 135 248
rect 139 244 140 248
rect 134 243 140 244
rect 222 248 228 249
rect 222 244 223 248
rect 227 244 228 248
rect 222 243 228 244
rect 310 248 316 249
rect 310 244 311 248
rect 315 244 316 248
rect 310 243 316 244
rect 390 248 396 249
rect 390 244 391 248
rect 395 244 396 248
rect 390 243 396 244
rect 462 248 468 249
rect 462 244 463 248
rect 467 244 468 248
rect 462 243 468 244
rect 526 248 532 249
rect 526 244 527 248
rect 531 244 532 248
rect 526 243 532 244
rect 590 248 596 249
rect 590 244 591 248
rect 595 244 596 248
rect 590 243 596 244
rect 646 248 652 249
rect 646 244 647 248
rect 651 244 652 248
rect 646 243 652 244
rect 694 248 700 249
rect 694 244 695 248
rect 699 244 700 248
rect 694 243 700 244
rect 734 248 740 249
rect 734 244 735 248
rect 739 244 740 248
rect 734 243 740 244
rect 782 248 788 249
rect 782 244 783 248
rect 787 244 788 248
rect 782 243 788 244
rect 830 248 836 249
rect 830 244 831 248
rect 835 244 836 248
rect 830 243 836 244
rect 878 248 884 249
rect 878 244 879 248
rect 883 244 884 248
rect 878 243 884 244
rect 926 248 932 249
rect 926 244 927 248
rect 931 244 932 248
rect 926 243 932 244
rect 974 248 980 249
rect 974 244 975 248
rect 979 244 980 248
rect 974 243 980 244
rect 1022 248 1028 249
rect 1022 244 1023 248
rect 1027 244 1028 248
rect 1022 243 1028 244
rect 110 241 116 242
rect 110 237 111 241
rect 115 237 116 241
rect 110 236 116 237
rect 1238 241 1244 242
rect 1238 237 1239 241
rect 1243 237 1244 241
rect 1238 236 1244 237
rect 1366 240 1372 241
rect 1366 236 1367 240
rect 1371 236 1372 240
rect 1366 235 1372 236
rect 1406 240 1412 241
rect 1406 236 1407 240
rect 1411 236 1412 240
rect 1406 235 1412 236
rect 1454 240 1460 241
rect 1454 236 1455 240
rect 1459 236 1460 240
rect 1454 235 1460 236
rect 1510 240 1516 241
rect 1510 236 1511 240
rect 1515 236 1516 240
rect 1510 235 1516 236
rect 1566 240 1572 241
rect 1566 236 1567 240
rect 1571 236 1572 240
rect 1566 235 1572 236
rect 1630 240 1636 241
rect 1630 236 1631 240
rect 1635 236 1636 240
rect 1630 235 1636 236
rect 1702 240 1708 241
rect 1702 236 1703 240
rect 1707 236 1708 240
rect 1702 235 1708 236
rect 1774 240 1780 241
rect 1774 236 1775 240
rect 1779 236 1780 240
rect 1774 235 1780 236
rect 1854 240 1860 241
rect 1854 236 1855 240
rect 1859 236 1860 240
rect 1854 235 1860 236
rect 1942 240 1948 241
rect 1942 236 1943 240
rect 1947 236 1948 240
rect 1942 235 1948 236
rect 2030 240 2036 241
rect 2030 236 2031 240
rect 2035 236 2036 240
rect 2030 235 2036 236
rect 2118 240 2124 241
rect 2118 236 2119 240
rect 2123 236 2124 240
rect 2118 235 2124 236
rect 2206 240 2212 241
rect 2206 236 2207 240
rect 2211 236 2212 240
rect 2206 235 2212 236
rect 2294 240 2300 241
rect 2294 236 2295 240
rect 2299 236 2300 240
rect 2294 235 2300 236
rect 2358 240 2364 241
rect 2358 236 2359 240
rect 2363 236 2364 240
rect 2358 235 2364 236
rect 1278 233 1284 234
rect 1278 229 1279 233
rect 1283 229 1284 233
rect 1278 228 1284 229
rect 2406 233 2412 234
rect 2406 229 2407 233
rect 2411 229 2412 233
rect 2406 228 2412 229
rect 110 224 116 225
rect 110 220 111 224
rect 115 220 116 224
rect 110 219 116 220
rect 1238 224 1244 225
rect 1238 220 1239 224
rect 1243 220 1244 224
rect 1238 219 1244 220
rect 1278 216 1284 217
rect 1278 212 1279 216
rect 1283 212 1284 216
rect 1278 211 1284 212
rect 2406 216 2412 217
rect 2406 212 2407 216
rect 2411 212 2412 216
rect 2406 211 2412 212
rect 134 201 140 202
rect 134 197 135 201
rect 139 197 140 201
rect 134 196 140 197
rect 222 201 228 202
rect 222 197 223 201
rect 227 197 228 201
rect 222 196 228 197
rect 310 201 316 202
rect 310 197 311 201
rect 315 197 316 201
rect 310 196 316 197
rect 390 201 396 202
rect 390 197 391 201
rect 395 197 396 201
rect 390 196 396 197
rect 462 201 468 202
rect 462 197 463 201
rect 467 197 468 201
rect 462 196 468 197
rect 526 201 532 202
rect 526 197 527 201
rect 531 197 532 201
rect 526 196 532 197
rect 590 201 596 202
rect 590 197 591 201
rect 595 197 596 201
rect 590 196 596 197
rect 646 201 652 202
rect 646 197 647 201
rect 651 197 652 201
rect 646 196 652 197
rect 694 201 700 202
rect 694 197 695 201
rect 699 197 700 201
rect 694 196 700 197
rect 734 201 740 202
rect 734 197 735 201
rect 739 197 740 201
rect 734 196 740 197
rect 782 201 788 202
rect 782 197 783 201
rect 787 197 788 201
rect 782 196 788 197
rect 830 201 836 202
rect 830 197 831 201
rect 835 197 836 201
rect 830 196 836 197
rect 878 201 884 202
rect 878 197 879 201
rect 883 197 884 201
rect 878 196 884 197
rect 926 201 932 202
rect 926 197 927 201
rect 931 197 932 201
rect 926 196 932 197
rect 974 201 980 202
rect 974 197 975 201
rect 979 197 980 201
rect 974 196 980 197
rect 1022 201 1028 202
rect 1022 197 1023 201
rect 1027 197 1028 201
rect 1022 196 1028 197
rect 1366 193 1372 194
rect 1366 189 1367 193
rect 1371 189 1372 193
rect 1366 188 1372 189
rect 1406 193 1412 194
rect 1406 189 1407 193
rect 1411 189 1412 193
rect 1406 188 1412 189
rect 1454 193 1460 194
rect 1454 189 1455 193
rect 1459 189 1460 193
rect 1454 188 1460 189
rect 1510 193 1516 194
rect 1510 189 1511 193
rect 1515 189 1516 193
rect 1510 188 1516 189
rect 1566 193 1572 194
rect 1566 189 1567 193
rect 1571 189 1572 193
rect 1566 188 1572 189
rect 1630 193 1636 194
rect 1630 189 1631 193
rect 1635 189 1636 193
rect 1630 188 1636 189
rect 1702 193 1708 194
rect 1702 189 1703 193
rect 1707 189 1708 193
rect 1702 188 1708 189
rect 1774 193 1780 194
rect 1774 189 1775 193
rect 1779 189 1780 193
rect 1774 188 1780 189
rect 1854 193 1860 194
rect 1854 189 1855 193
rect 1859 189 1860 193
rect 1854 188 1860 189
rect 1942 193 1948 194
rect 1942 189 1943 193
rect 1947 189 1948 193
rect 1942 188 1948 189
rect 2030 193 2036 194
rect 2030 189 2031 193
rect 2035 189 2036 193
rect 2030 188 2036 189
rect 2118 193 2124 194
rect 2118 189 2119 193
rect 2123 189 2124 193
rect 2118 188 2124 189
rect 2206 193 2212 194
rect 2206 189 2207 193
rect 2211 189 2212 193
rect 2206 188 2212 189
rect 2294 193 2300 194
rect 2294 189 2295 193
rect 2299 189 2300 193
rect 2294 188 2300 189
rect 2358 193 2364 194
rect 2358 189 2359 193
rect 2363 189 2364 193
rect 2358 188 2364 189
rect 1302 155 1308 156
rect 1302 151 1303 155
rect 1307 151 1308 155
rect 1302 150 1308 151
rect 1342 155 1348 156
rect 1342 151 1343 155
rect 1347 151 1348 155
rect 1342 150 1348 151
rect 1382 155 1388 156
rect 1382 151 1383 155
rect 1387 151 1388 155
rect 1382 150 1388 151
rect 1422 155 1428 156
rect 1422 151 1423 155
rect 1427 151 1428 155
rect 1422 150 1428 151
rect 1462 155 1468 156
rect 1462 151 1463 155
rect 1467 151 1468 155
rect 1462 150 1468 151
rect 1518 155 1524 156
rect 1518 151 1519 155
rect 1523 151 1524 155
rect 1518 150 1524 151
rect 1582 155 1588 156
rect 1582 151 1583 155
rect 1587 151 1588 155
rect 1582 150 1588 151
rect 1646 155 1652 156
rect 1646 151 1647 155
rect 1651 151 1652 155
rect 1646 150 1652 151
rect 1710 155 1716 156
rect 1710 151 1711 155
rect 1715 151 1716 155
rect 1710 150 1716 151
rect 1774 155 1780 156
rect 1774 151 1775 155
rect 1779 151 1780 155
rect 1774 150 1780 151
rect 1830 155 1836 156
rect 1830 151 1831 155
rect 1835 151 1836 155
rect 1830 150 1836 151
rect 1886 155 1892 156
rect 1886 151 1887 155
rect 1891 151 1892 155
rect 1886 150 1892 151
rect 1934 155 1940 156
rect 1934 151 1935 155
rect 1939 151 1940 155
rect 1934 150 1940 151
rect 1974 155 1980 156
rect 1974 151 1975 155
rect 1979 151 1980 155
rect 1974 150 1980 151
rect 2014 155 2020 156
rect 2014 151 2015 155
rect 2019 151 2020 155
rect 2014 150 2020 151
rect 2054 155 2060 156
rect 2054 151 2055 155
rect 2059 151 2060 155
rect 2054 150 2060 151
rect 2094 155 2100 156
rect 2094 151 2095 155
rect 2099 151 2100 155
rect 2094 150 2100 151
rect 2142 155 2148 156
rect 2142 151 2143 155
rect 2147 151 2148 155
rect 2142 150 2148 151
rect 2190 155 2196 156
rect 2190 151 2191 155
rect 2195 151 2196 155
rect 2190 150 2196 151
rect 2238 155 2244 156
rect 2238 151 2239 155
rect 2243 151 2244 155
rect 2238 150 2244 151
rect 2278 155 2284 156
rect 2278 151 2279 155
rect 2283 151 2284 155
rect 2278 150 2284 151
rect 2318 155 2324 156
rect 2318 151 2319 155
rect 2323 151 2324 155
rect 2318 150 2324 151
rect 2358 155 2364 156
rect 2358 151 2359 155
rect 2363 151 2364 155
rect 2358 150 2364 151
rect 150 139 156 140
rect 150 135 151 139
rect 155 135 156 139
rect 150 134 156 135
rect 190 139 196 140
rect 190 135 191 139
rect 195 135 196 139
rect 190 134 196 135
rect 230 139 236 140
rect 230 135 231 139
rect 235 135 236 139
rect 230 134 236 135
rect 270 139 276 140
rect 270 135 271 139
rect 275 135 276 139
rect 270 134 276 135
rect 310 139 316 140
rect 310 135 311 139
rect 315 135 316 139
rect 310 134 316 135
rect 350 139 356 140
rect 350 135 351 139
rect 355 135 356 139
rect 350 134 356 135
rect 390 139 396 140
rect 390 135 391 139
rect 395 135 396 139
rect 390 134 396 135
rect 430 139 436 140
rect 430 135 431 139
rect 435 135 436 139
rect 430 134 436 135
rect 470 139 476 140
rect 470 135 471 139
rect 475 135 476 139
rect 470 134 476 135
rect 510 139 516 140
rect 510 135 511 139
rect 515 135 516 139
rect 510 134 516 135
rect 550 139 556 140
rect 550 135 551 139
rect 555 135 556 139
rect 550 134 556 135
rect 590 139 596 140
rect 590 135 591 139
rect 595 135 596 139
rect 590 134 596 135
rect 630 139 636 140
rect 630 135 631 139
rect 635 135 636 139
rect 630 134 636 135
rect 670 139 676 140
rect 670 135 671 139
rect 675 135 676 139
rect 670 134 676 135
rect 710 139 716 140
rect 710 135 711 139
rect 715 135 716 139
rect 710 134 716 135
rect 750 139 756 140
rect 750 135 751 139
rect 755 135 756 139
rect 750 134 756 135
rect 790 139 796 140
rect 790 135 791 139
rect 795 135 796 139
rect 790 134 796 135
rect 830 139 836 140
rect 830 135 831 139
rect 835 135 836 139
rect 830 134 836 135
rect 870 139 876 140
rect 870 135 871 139
rect 875 135 876 139
rect 870 134 876 135
rect 910 139 916 140
rect 910 135 911 139
rect 915 135 916 139
rect 910 134 916 135
rect 950 139 956 140
rect 950 135 951 139
rect 955 135 956 139
rect 950 134 956 135
rect 990 139 996 140
rect 990 135 991 139
rect 995 135 996 139
rect 990 134 996 135
rect 1030 139 1036 140
rect 1030 135 1031 139
rect 1035 135 1036 139
rect 1030 134 1036 135
rect 1070 139 1076 140
rect 1070 135 1071 139
rect 1075 135 1076 139
rect 1070 134 1076 135
rect 1110 139 1116 140
rect 1110 135 1111 139
rect 1115 135 1116 139
rect 1110 134 1116 135
rect 1150 139 1156 140
rect 1150 135 1151 139
rect 1155 135 1156 139
rect 1150 134 1156 135
rect 1190 139 1196 140
rect 1190 135 1191 139
rect 1195 135 1196 139
rect 1190 134 1196 135
rect 1278 132 1284 133
rect 1278 128 1279 132
rect 1283 128 1284 132
rect 1278 127 1284 128
rect 2406 132 2412 133
rect 2406 128 2407 132
rect 2411 128 2412 132
rect 2406 127 2412 128
rect 110 116 116 117
rect 110 112 111 116
rect 115 112 116 116
rect 110 111 116 112
rect 1238 116 1244 117
rect 1238 112 1239 116
rect 1243 112 1244 116
rect 1238 111 1244 112
rect 1278 115 1284 116
rect 1278 111 1279 115
rect 1283 111 1284 115
rect 1278 110 1284 111
rect 2406 115 2412 116
rect 2406 111 2407 115
rect 2411 111 2412 115
rect 2406 110 2412 111
rect 1302 108 1308 109
rect 1302 104 1303 108
rect 1307 104 1308 108
rect 1302 103 1308 104
rect 1342 108 1348 109
rect 1342 104 1343 108
rect 1347 104 1348 108
rect 1342 103 1348 104
rect 1382 108 1388 109
rect 1382 104 1383 108
rect 1387 104 1388 108
rect 1382 103 1388 104
rect 1422 108 1428 109
rect 1422 104 1423 108
rect 1427 104 1428 108
rect 1422 103 1428 104
rect 1462 108 1468 109
rect 1462 104 1463 108
rect 1467 104 1468 108
rect 1462 103 1468 104
rect 1518 108 1524 109
rect 1518 104 1519 108
rect 1523 104 1524 108
rect 1518 103 1524 104
rect 1582 108 1588 109
rect 1582 104 1583 108
rect 1587 104 1588 108
rect 1582 103 1588 104
rect 1646 108 1652 109
rect 1646 104 1647 108
rect 1651 104 1652 108
rect 1646 103 1652 104
rect 1710 108 1716 109
rect 1710 104 1711 108
rect 1715 104 1716 108
rect 1710 103 1716 104
rect 1774 108 1780 109
rect 1774 104 1775 108
rect 1779 104 1780 108
rect 1774 103 1780 104
rect 1830 108 1836 109
rect 1830 104 1831 108
rect 1835 104 1836 108
rect 1830 103 1836 104
rect 1886 108 1892 109
rect 1886 104 1887 108
rect 1891 104 1892 108
rect 1886 103 1892 104
rect 1934 108 1940 109
rect 1934 104 1935 108
rect 1939 104 1940 108
rect 1934 103 1940 104
rect 1974 108 1980 109
rect 1974 104 1975 108
rect 1979 104 1980 108
rect 1974 103 1980 104
rect 2014 108 2020 109
rect 2014 104 2015 108
rect 2019 104 2020 108
rect 2014 103 2020 104
rect 2054 108 2060 109
rect 2054 104 2055 108
rect 2059 104 2060 108
rect 2054 103 2060 104
rect 2094 108 2100 109
rect 2094 104 2095 108
rect 2099 104 2100 108
rect 2094 103 2100 104
rect 2142 108 2148 109
rect 2142 104 2143 108
rect 2147 104 2148 108
rect 2142 103 2148 104
rect 2190 108 2196 109
rect 2190 104 2191 108
rect 2195 104 2196 108
rect 2190 103 2196 104
rect 2238 108 2244 109
rect 2238 104 2239 108
rect 2243 104 2244 108
rect 2238 103 2244 104
rect 2278 108 2284 109
rect 2278 104 2279 108
rect 2283 104 2284 108
rect 2278 103 2284 104
rect 2318 108 2324 109
rect 2318 104 2319 108
rect 2323 104 2324 108
rect 2318 103 2324 104
rect 2358 108 2364 109
rect 2358 104 2359 108
rect 2363 104 2364 108
rect 2358 103 2364 104
rect 110 99 116 100
rect 110 95 111 99
rect 115 95 116 99
rect 110 94 116 95
rect 1238 99 1244 100
rect 1238 95 1239 99
rect 1243 95 1244 99
rect 1238 94 1244 95
rect 150 92 156 93
rect 150 88 151 92
rect 155 88 156 92
rect 150 87 156 88
rect 190 92 196 93
rect 190 88 191 92
rect 195 88 196 92
rect 190 87 196 88
rect 230 92 236 93
rect 230 88 231 92
rect 235 88 236 92
rect 230 87 236 88
rect 270 92 276 93
rect 270 88 271 92
rect 275 88 276 92
rect 270 87 276 88
rect 310 92 316 93
rect 310 88 311 92
rect 315 88 316 92
rect 310 87 316 88
rect 350 92 356 93
rect 350 88 351 92
rect 355 88 356 92
rect 350 87 356 88
rect 390 92 396 93
rect 390 88 391 92
rect 395 88 396 92
rect 390 87 396 88
rect 430 92 436 93
rect 430 88 431 92
rect 435 88 436 92
rect 430 87 436 88
rect 470 92 476 93
rect 470 88 471 92
rect 475 88 476 92
rect 470 87 476 88
rect 510 92 516 93
rect 510 88 511 92
rect 515 88 516 92
rect 510 87 516 88
rect 550 92 556 93
rect 550 88 551 92
rect 555 88 556 92
rect 550 87 556 88
rect 590 92 596 93
rect 590 88 591 92
rect 595 88 596 92
rect 590 87 596 88
rect 630 92 636 93
rect 630 88 631 92
rect 635 88 636 92
rect 630 87 636 88
rect 670 92 676 93
rect 670 88 671 92
rect 675 88 676 92
rect 670 87 676 88
rect 710 92 716 93
rect 710 88 711 92
rect 715 88 716 92
rect 710 87 716 88
rect 750 92 756 93
rect 750 88 751 92
rect 755 88 756 92
rect 750 87 756 88
rect 790 92 796 93
rect 790 88 791 92
rect 795 88 796 92
rect 790 87 796 88
rect 830 92 836 93
rect 830 88 831 92
rect 835 88 836 92
rect 830 87 836 88
rect 870 92 876 93
rect 870 88 871 92
rect 875 88 876 92
rect 870 87 876 88
rect 910 92 916 93
rect 910 88 911 92
rect 915 88 916 92
rect 910 87 916 88
rect 950 92 956 93
rect 950 88 951 92
rect 955 88 956 92
rect 950 87 956 88
rect 990 92 996 93
rect 990 88 991 92
rect 995 88 996 92
rect 990 87 996 88
rect 1030 92 1036 93
rect 1030 88 1031 92
rect 1035 88 1036 92
rect 1030 87 1036 88
rect 1070 92 1076 93
rect 1070 88 1071 92
rect 1075 88 1076 92
rect 1070 87 1076 88
rect 1110 92 1116 93
rect 1110 88 1111 92
rect 1115 88 1116 92
rect 1110 87 1116 88
rect 1150 92 1156 93
rect 1150 88 1151 92
rect 1155 88 1156 92
rect 1150 87 1156 88
rect 1190 92 1196 93
rect 1190 88 1191 92
rect 1195 88 1196 92
rect 1190 87 1196 88
<< m3c >>
rect 231 2475 235 2479
rect 271 2475 275 2479
rect 311 2475 315 2479
rect 351 2475 355 2479
rect 399 2475 403 2479
rect 455 2475 459 2479
rect 511 2475 515 2479
rect 575 2475 579 2479
rect 639 2475 643 2479
rect 703 2475 707 2479
rect 767 2475 771 2479
rect 823 2475 827 2479
rect 879 2475 883 2479
rect 927 2475 931 2479
rect 975 2475 979 2479
rect 1023 2475 1027 2479
rect 1071 2475 1075 2479
rect 1111 2475 1115 2479
rect 1151 2475 1155 2479
rect 1191 2475 1195 2479
rect 1303 2471 1307 2475
rect 1343 2471 1347 2475
rect 1383 2471 1387 2475
rect 1439 2471 1443 2475
rect 1511 2471 1515 2475
rect 1583 2471 1587 2475
rect 1663 2471 1667 2475
rect 1735 2471 1739 2475
rect 1807 2471 1811 2475
rect 1887 2471 1891 2475
rect 1967 2471 1971 2475
rect 2063 2471 2067 2475
rect 2167 2471 2171 2475
rect 2271 2471 2275 2475
rect 2359 2471 2363 2475
rect 111 2452 115 2456
rect 1239 2452 1243 2456
rect 1279 2448 1283 2452
rect 2407 2448 2411 2452
rect 111 2435 115 2439
rect 1239 2435 1243 2439
rect 231 2428 235 2432
rect 271 2428 275 2432
rect 311 2428 315 2432
rect 351 2428 355 2432
rect 399 2428 403 2432
rect 455 2428 459 2432
rect 511 2428 515 2432
rect 575 2428 579 2432
rect 639 2428 643 2432
rect 703 2428 707 2432
rect 767 2428 771 2432
rect 823 2428 827 2432
rect 879 2428 883 2432
rect 927 2428 931 2432
rect 975 2428 979 2432
rect 1023 2428 1027 2432
rect 1071 2428 1075 2432
rect 1111 2428 1115 2432
rect 1151 2428 1155 2432
rect 1191 2428 1195 2432
rect 1279 2431 1283 2435
rect 2407 2431 2411 2435
rect 1303 2424 1307 2428
rect 1343 2424 1347 2428
rect 1383 2424 1387 2428
rect 1439 2424 1443 2428
rect 1511 2424 1515 2428
rect 1583 2424 1587 2428
rect 1663 2424 1667 2428
rect 1735 2424 1739 2428
rect 1807 2424 1811 2428
rect 1887 2424 1891 2428
rect 1967 2424 1971 2428
rect 2063 2424 2067 2428
rect 2167 2424 2171 2428
rect 2271 2424 2275 2428
rect 2359 2424 2363 2428
rect 199 2408 203 2412
rect 263 2408 267 2412
rect 327 2408 331 2412
rect 399 2408 403 2412
rect 471 2408 475 2412
rect 543 2408 547 2412
rect 615 2408 619 2412
rect 687 2408 691 2412
rect 751 2408 755 2412
rect 823 2408 827 2412
rect 895 2408 899 2412
rect 967 2408 971 2412
rect 1375 2412 1379 2416
rect 1415 2412 1419 2416
rect 1455 2412 1459 2416
rect 1503 2412 1507 2416
rect 1559 2412 1563 2416
rect 1615 2412 1619 2416
rect 1679 2412 1683 2416
rect 1735 2412 1739 2416
rect 1799 2412 1803 2416
rect 1871 2412 1875 2416
rect 1951 2412 1955 2416
rect 2047 2412 2051 2416
rect 2151 2412 2155 2416
rect 2263 2412 2267 2416
rect 2359 2412 2363 2416
rect 111 2401 115 2405
rect 1239 2401 1243 2405
rect 1279 2405 1283 2409
rect 2407 2405 2411 2409
rect 111 2384 115 2388
rect 1239 2384 1243 2388
rect 1279 2388 1283 2392
rect 2407 2388 2411 2392
rect 199 2361 203 2365
rect 263 2361 267 2365
rect 327 2361 331 2365
rect 399 2361 403 2365
rect 471 2361 475 2365
rect 543 2361 547 2365
rect 615 2361 619 2365
rect 687 2361 691 2365
rect 751 2361 755 2365
rect 823 2361 827 2365
rect 895 2361 899 2365
rect 967 2361 971 2365
rect 1375 2365 1379 2369
rect 1415 2365 1419 2369
rect 1455 2365 1459 2369
rect 1503 2365 1507 2369
rect 1559 2365 1563 2369
rect 1615 2365 1619 2369
rect 1679 2365 1683 2369
rect 1735 2365 1739 2369
rect 1799 2365 1803 2369
rect 1871 2365 1875 2369
rect 1951 2365 1955 2369
rect 2047 2365 2051 2369
rect 2151 2365 2155 2369
rect 2263 2365 2267 2369
rect 2359 2365 2363 2369
rect 271 2327 275 2331
rect 327 2327 331 2331
rect 399 2327 403 2331
rect 471 2327 475 2331
rect 551 2327 555 2331
rect 631 2327 635 2331
rect 711 2327 715 2331
rect 783 2327 787 2331
rect 855 2327 859 2331
rect 919 2327 923 2331
rect 991 2327 995 2331
rect 1063 2327 1067 2331
rect 1327 2331 1331 2335
rect 1383 2331 1387 2335
rect 1439 2331 1443 2335
rect 1503 2331 1507 2335
rect 1575 2331 1579 2335
rect 1647 2331 1651 2335
rect 1719 2331 1723 2335
rect 1799 2331 1803 2335
rect 1879 2331 1883 2335
rect 1967 2331 1971 2335
rect 2063 2331 2067 2335
rect 2167 2331 2171 2335
rect 2271 2331 2275 2335
rect 2359 2331 2363 2335
rect 111 2304 115 2308
rect 1239 2304 1243 2308
rect 1279 2308 1283 2312
rect 2407 2308 2411 2312
rect 111 2287 115 2291
rect 1239 2287 1243 2291
rect 1279 2291 1283 2295
rect 2407 2291 2411 2295
rect 271 2280 275 2284
rect 327 2280 331 2284
rect 399 2280 403 2284
rect 471 2280 475 2284
rect 551 2280 555 2284
rect 631 2280 635 2284
rect 711 2280 715 2284
rect 783 2280 787 2284
rect 855 2280 859 2284
rect 919 2280 923 2284
rect 991 2280 995 2284
rect 1063 2280 1067 2284
rect 1327 2284 1331 2288
rect 1383 2284 1387 2288
rect 1439 2284 1443 2288
rect 1503 2284 1507 2288
rect 1575 2284 1579 2288
rect 1647 2284 1651 2288
rect 1719 2284 1723 2288
rect 1799 2284 1803 2288
rect 1879 2284 1883 2288
rect 1967 2284 1971 2288
rect 2063 2284 2067 2288
rect 2167 2284 2171 2288
rect 2271 2284 2275 2288
rect 2359 2284 2363 2288
rect 1335 2272 1339 2276
rect 1407 2272 1411 2276
rect 1487 2272 1491 2276
rect 1559 2272 1563 2276
rect 1631 2272 1635 2276
rect 1703 2272 1707 2276
rect 1775 2272 1779 2276
rect 1839 2272 1843 2276
rect 1911 2272 1915 2276
rect 1991 2272 1995 2276
rect 2079 2272 2083 2276
rect 2175 2272 2179 2276
rect 2279 2272 2283 2276
rect 2359 2272 2363 2276
rect 1279 2265 1283 2269
rect 143 2260 147 2264
rect 183 2260 187 2264
rect 223 2260 227 2264
rect 279 2260 283 2264
rect 335 2260 339 2264
rect 407 2260 411 2264
rect 479 2260 483 2264
rect 559 2260 563 2264
rect 647 2260 651 2264
rect 727 2260 731 2264
rect 807 2260 811 2264
rect 887 2260 891 2264
rect 967 2260 971 2264
rect 1047 2260 1051 2264
rect 2407 2265 2411 2269
rect 1127 2260 1131 2264
rect 111 2253 115 2257
rect 1239 2253 1243 2257
rect 1279 2248 1283 2252
rect 2407 2248 2411 2252
rect 111 2236 115 2240
rect 1239 2236 1243 2240
rect 1335 2225 1339 2229
rect 1407 2225 1411 2229
rect 1487 2225 1491 2229
rect 1559 2225 1563 2229
rect 1631 2225 1635 2229
rect 1703 2225 1707 2229
rect 1775 2225 1779 2229
rect 1839 2225 1843 2229
rect 1911 2225 1915 2229
rect 1991 2225 1995 2229
rect 2079 2225 2083 2229
rect 2175 2225 2179 2229
rect 2279 2225 2283 2229
rect 2359 2225 2363 2229
rect 143 2213 147 2217
rect 183 2213 187 2217
rect 223 2213 227 2217
rect 279 2213 283 2217
rect 335 2213 339 2217
rect 407 2213 411 2217
rect 479 2213 483 2217
rect 559 2213 563 2217
rect 647 2213 651 2217
rect 727 2213 731 2217
rect 807 2213 811 2217
rect 887 2213 891 2217
rect 967 2213 971 2217
rect 1047 2213 1051 2217
rect 1127 2213 1131 2217
rect 135 2183 139 2187
rect 207 2183 211 2187
rect 279 2183 283 2187
rect 359 2183 363 2187
rect 439 2183 443 2187
rect 519 2183 523 2187
rect 599 2183 603 2187
rect 679 2183 683 2187
rect 759 2183 763 2187
rect 831 2183 835 2187
rect 903 2183 907 2187
rect 975 2183 979 2187
rect 1047 2183 1051 2187
rect 1119 2183 1123 2187
rect 1375 2187 1379 2191
rect 1439 2187 1443 2191
rect 1511 2187 1515 2191
rect 1591 2187 1595 2191
rect 1671 2187 1675 2191
rect 1751 2187 1755 2191
rect 1831 2187 1835 2191
rect 1903 2187 1907 2191
rect 1967 2187 1971 2191
rect 2031 2187 2035 2191
rect 2095 2187 2099 2191
rect 2167 2187 2171 2191
rect 2239 2187 2243 2191
rect 2311 2187 2315 2191
rect 2359 2187 2363 2191
rect 111 2160 115 2164
rect 1239 2160 1243 2164
rect 1279 2164 1283 2168
rect 2407 2164 2411 2168
rect 111 2143 115 2147
rect 1239 2143 1243 2147
rect 1279 2147 1283 2151
rect 2407 2147 2411 2151
rect 135 2136 139 2140
rect 207 2136 211 2140
rect 279 2136 283 2140
rect 359 2136 363 2140
rect 439 2136 443 2140
rect 519 2136 523 2140
rect 599 2136 603 2140
rect 679 2136 683 2140
rect 759 2136 763 2140
rect 831 2136 835 2140
rect 903 2136 907 2140
rect 975 2136 979 2140
rect 1047 2136 1051 2140
rect 1119 2136 1123 2140
rect 1375 2140 1379 2144
rect 1439 2140 1443 2144
rect 1511 2140 1515 2144
rect 1591 2140 1595 2144
rect 1671 2140 1675 2144
rect 1751 2140 1755 2144
rect 1831 2140 1835 2144
rect 1903 2140 1907 2144
rect 1967 2140 1971 2144
rect 2031 2140 2035 2144
rect 2095 2140 2099 2144
rect 2167 2140 2171 2144
rect 2239 2140 2243 2144
rect 2311 2140 2315 2144
rect 2359 2140 2363 2144
rect 1399 2128 1403 2132
rect 1439 2128 1443 2132
rect 1495 2128 1499 2132
rect 1567 2128 1571 2132
rect 1647 2128 1651 2132
rect 1735 2128 1739 2132
rect 1823 2128 1827 2132
rect 1911 2128 1915 2132
rect 1999 2128 2003 2132
rect 2087 2128 2091 2132
rect 2175 2128 2179 2132
rect 2271 2128 2275 2132
rect 2359 2128 2363 2132
rect 1279 2121 1283 2125
rect 135 2116 139 2120
rect 191 2116 195 2120
rect 271 2116 275 2120
rect 343 2116 347 2120
rect 415 2116 419 2120
rect 479 2116 483 2120
rect 543 2116 547 2120
rect 607 2116 611 2120
rect 671 2116 675 2120
rect 735 2116 739 2120
rect 791 2116 795 2120
rect 839 2116 843 2120
rect 887 2116 891 2120
rect 935 2116 939 2120
rect 991 2116 995 2120
rect 2407 2121 2411 2125
rect 1047 2116 1051 2120
rect 111 2109 115 2113
rect 1239 2109 1243 2113
rect 1279 2104 1283 2108
rect 2407 2104 2411 2108
rect 111 2092 115 2096
rect 1239 2092 1243 2096
rect 1399 2081 1403 2085
rect 1439 2081 1443 2085
rect 1495 2081 1499 2085
rect 1567 2081 1571 2085
rect 1647 2081 1651 2085
rect 1735 2081 1739 2085
rect 1823 2081 1827 2085
rect 1911 2081 1915 2085
rect 1999 2081 2003 2085
rect 2087 2081 2091 2085
rect 2175 2081 2179 2085
rect 2271 2081 2275 2085
rect 2359 2081 2363 2085
rect 135 2069 139 2073
rect 191 2069 195 2073
rect 271 2069 275 2073
rect 343 2069 347 2073
rect 415 2069 419 2073
rect 479 2069 483 2073
rect 543 2069 547 2073
rect 607 2069 611 2073
rect 671 2069 675 2073
rect 735 2069 739 2073
rect 791 2069 795 2073
rect 839 2069 843 2073
rect 887 2069 891 2073
rect 935 2069 939 2073
rect 991 2069 995 2073
rect 1047 2069 1051 2073
rect 2039 2051 2043 2055
rect 2079 2051 2083 2055
rect 2119 2051 2123 2055
rect 2159 2051 2163 2055
rect 2199 2051 2203 2055
rect 2239 2051 2243 2055
rect 2279 2051 2283 2055
rect 2319 2051 2323 2055
rect 2359 2051 2363 2055
rect 135 2035 139 2039
rect 175 2035 179 2039
rect 215 2035 219 2039
rect 279 2035 283 2039
rect 351 2035 355 2039
rect 423 2035 427 2039
rect 487 2035 491 2039
rect 551 2035 555 2039
rect 615 2035 619 2039
rect 679 2035 683 2039
rect 743 2035 747 2039
rect 815 2035 819 2039
rect 1279 2028 1283 2032
rect 2407 2028 2411 2032
rect 111 2012 115 2016
rect 1239 2012 1243 2016
rect 1279 2011 1283 2015
rect 2407 2011 2411 2015
rect 2039 2004 2043 2008
rect 2079 2004 2083 2008
rect 2119 2004 2123 2008
rect 2159 2004 2163 2008
rect 2199 2004 2203 2008
rect 2239 2004 2243 2008
rect 2279 2004 2283 2008
rect 2319 2004 2323 2008
rect 2359 2004 2363 2008
rect 111 1995 115 1999
rect 1239 1995 1243 1999
rect 135 1988 139 1992
rect 175 1988 179 1992
rect 215 1988 219 1992
rect 279 1988 283 1992
rect 351 1988 355 1992
rect 423 1988 427 1992
rect 487 1988 491 1992
rect 551 1988 555 1992
rect 615 1988 619 1992
rect 679 1988 683 1992
rect 743 1988 747 1992
rect 815 1988 819 1992
rect 1399 1992 1403 1996
rect 1439 1992 1443 1996
rect 1479 1992 1483 1996
rect 1519 1992 1523 1996
rect 1559 1992 1563 1996
rect 1599 1992 1603 1996
rect 1639 1992 1643 1996
rect 1679 1992 1683 1996
rect 1719 1992 1723 1996
rect 1767 1992 1771 1996
rect 1823 1992 1827 1996
rect 1871 1992 1875 1996
rect 1919 1992 1923 1996
rect 1967 1992 1971 1996
rect 2015 1992 2019 1996
rect 2055 1992 2059 1996
rect 2095 1992 2099 1996
rect 2143 1992 2147 1996
rect 2191 1992 2195 1996
rect 2239 1992 2243 1996
rect 2279 1992 2283 1996
rect 2319 1992 2323 1996
rect 2359 1992 2363 1996
rect 1279 1985 1283 1989
rect 2407 1985 2411 1989
rect 135 1976 139 1980
rect 175 1976 179 1980
rect 215 1976 219 1980
rect 271 1976 275 1980
rect 343 1976 347 1980
rect 415 1976 419 1980
rect 495 1976 499 1980
rect 575 1976 579 1980
rect 647 1976 651 1980
rect 719 1976 723 1980
rect 791 1976 795 1980
rect 863 1976 867 1980
rect 935 1976 939 1980
rect 1007 1976 1011 1980
rect 111 1969 115 1973
rect 1239 1969 1243 1973
rect 1279 1968 1283 1972
rect 2407 1968 2411 1972
rect 111 1952 115 1956
rect 1239 1952 1243 1956
rect 1399 1945 1403 1949
rect 1439 1945 1443 1949
rect 1479 1945 1483 1949
rect 1519 1945 1523 1949
rect 1559 1945 1563 1949
rect 1599 1945 1603 1949
rect 1639 1945 1643 1949
rect 1679 1945 1683 1949
rect 1719 1945 1723 1949
rect 1767 1945 1771 1949
rect 1823 1945 1827 1949
rect 1871 1945 1875 1949
rect 1919 1945 1923 1949
rect 1967 1945 1971 1949
rect 2015 1945 2019 1949
rect 2055 1945 2059 1949
rect 2095 1945 2099 1949
rect 2143 1945 2147 1949
rect 2191 1945 2195 1949
rect 2239 1945 2243 1949
rect 2279 1945 2283 1949
rect 2319 1945 2323 1949
rect 2359 1945 2363 1949
rect 135 1929 139 1933
rect 175 1929 179 1933
rect 215 1929 219 1933
rect 271 1929 275 1933
rect 343 1929 347 1933
rect 415 1929 419 1933
rect 495 1929 499 1933
rect 575 1929 579 1933
rect 647 1929 651 1933
rect 719 1929 723 1933
rect 791 1929 795 1933
rect 863 1929 867 1933
rect 935 1929 939 1933
rect 1007 1929 1011 1933
rect 1343 1911 1347 1915
rect 1383 1911 1387 1915
rect 1423 1911 1427 1915
rect 1463 1911 1467 1915
rect 1511 1911 1515 1915
rect 1567 1911 1571 1915
rect 1631 1911 1635 1915
rect 1711 1911 1715 1915
rect 1807 1911 1811 1915
rect 1919 1911 1923 1915
rect 2031 1911 2035 1915
rect 2151 1911 2155 1915
rect 247 1895 251 1899
rect 287 1895 291 1899
rect 327 1895 331 1899
rect 367 1895 371 1899
rect 415 1895 419 1899
rect 471 1895 475 1899
rect 535 1895 539 1899
rect 599 1895 603 1899
rect 663 1895 667 1899
rect 727 1895 731 1899
rect 791 1895 795 1899
rect 855 1895 859 1899
rect 919 1895 923 1899
rect 983 1895 987 1899
rect 1055 1895 1059 1899
rect 1127 1895 1131 1899
rect 1279 1888 1283 1892
rect 2407 1888 2411 1892
rect 111 1872 115 1876
rect 1239 1872 1243 1876
rect 1279 1871 1283 1875
rect 2407 1871 2411 1875
rect 1343 1864 1347 1868
rect 1383 1864 1387 1868
rect 1423 1864 1427 1868
rect 1463 1864 1467 1868
rect 1511 1864 1515 1868
rect 1567 1864 1571 1868
rect 1631 1864 1635 1868
rect 1711 1864 1715 1868
rect 1807 1864 1811 1868
rect 1919 1864 1923 1868
rect 2031 1864 2035 1868
rect 2151 1864 2155 1868
rect 111 1855 115 1859
rect 1239 1855 1243 1859
rect 247 1848 251 1852
rect 287 1848 291 1852
rect 327 1848 331 1852
rect 367 1848 371 1852
rect 415 1848 419 1852
rect 471 1848 475 1852
rect 535 1848 539 1852
rect 599 1848 603 1852
rect 663 1848 667 1852
rect 727 1848 731 1852
rect 791 1848 795 1852
rect 855 1848 859 1852
rect 919 1848 923 1852
rect 983 1848 987 1852
rect 1055 1848 1059 1852
rect 1127 1848 1131 1852
rect 1359 1844 1363 1848
rect 1399 1844 1403 1848
rect 1447 1844 1451 1848
rect 1503 1844 1507 1848
rect 1559 1844 1563 1848
rect 1615 1844 1619 1848
rect 1671 1844 1675 1848
rect 1727 1844 1731 1848
rect 1783 1844 1787 1848
rect 1839 1844 1843 1848
rect 1895 1844 1899 1848
rect 1951 1844 1955 1848
rect 1279 1837 1283 1841
rect 399 1832 403 1836
rect 439 1832 443 1836
rect 479 1832 483 1836
rect 519 1832 523 1836
rect 567 1832 571 1836
rect 623 1832 627 1836
rect 687 1832 691 1836
rect 759 1832 763 1836
rect 831 1832 835 1836
rect 903 1832 907 1836
rect 975 1832 979 1836
rect 1047 1832 1051 1836
rect 1127 1832 1131 1836
rect 2407 1837 2411 1841
rect 1191 1832 1195 1836
rect 111 1825 115 1829
rect 1239 1825 1243 1829
rect 1279 1820 1283 1824
rect 2407 1820 2411 1824
rect 111 1808 115 1812
rect 1239 1808 1243 1812
rect 1359 1797 1363 1801
rect 1399 1797 1403 1801
rect 1447 1797 1451 1801
rect 1503 1797 1507 1801
rect 1559 1797 1563 1801
rect 1615 1797 1619 1801
rect 1671 1797 1675 1801
rect 1727 1797 1731 1801
rect 1783 1797 1787 1801
rect 1839 1797 1843 1801
rect 1895 1797 1899 1801
rect 1951 1797 1955 1801
rect 399 1785 403 1789
rect 439 1785 443 1789
rect 479 1785 483 1789
rect 519 1785 523 1789
rect 567 1785 571 1789
rect 623 1785 627 1789
rect 687 1785 691 1789
rect 759 1785 763 1789
rect 831 1785 835 1789
rect 903 1785 907 1789
rect 975 1785 979 1789
rect 1047 1785 1051 1789
rect 1127 1785 1131 1789
rect 1191 1785 1195 1789
rect 407 1755 411 1759
rect 447 1755 451 1759
rect 487 1755 491 1759
rect 527 1755 531 1759
rect 567 1755 571 1759
rect 607 1755 611 1759
rect 647 1755 651 1759
rect 695 1755 699 1759
rect 751 1755 755 1759
rect 807 1755 811 1759
rect 871 1755 875 1759
rect 935 1755 939 1759
rect 999 1755 1003 1759
rect 1071 1755 1075 1759
rect 1143 1755 1147 1759
rect 1191 1755 1195 1759
rect 1303 1755 1307 1759
rect 1343 1755 1347 1759
rect 1391 1755 1395 1759
rect 1455 1755 1459 1759
rect 1519 1755 1523 1759
rect 1583 1755 1587 1759
rect 1647 1755 1651 1759
rect 1703 1755 1707 1759
rect 1759 1755 1763 1759
rect 1807 1755 1811 1759
rect 1863 1755 1867 1759
rect 1919 1755 1923 1759
rect 1975 1755 1979 1759
rect 111 1732 115 1736
rect 1239 1732 1243 1736
rect 1279 1732 1283 1736
rect 2407 1732 2411 1736
rect 111 1715 115 1719
rect 1239 1715 1243 1719
rect 1279 1715 1283 1719
rect 2407 1715 2411 1719
rect 407 1708 411 1712
rect 447 1708 451 1712
rect 487 1708 491 1712
rect 527 1708 531 1712
rect 567 1708 571 1712
rect 607 1708 611 1712
rect 647 1708 651 1712
rect 695 1708 699 1712
rect 751 1708 755 1712
rect 807 1708 811 1712
rect 871 1708 875 1712
rect 935 1708 939 1712
rect 999 1708 1003 1712
rect 1071 1708 1075 1712
rect 1143 1708 1147 1712
rect 1191 1708 1195 1712
rect 1303 1708 1307 1712
rect 1343 1708 1347 1712
rect 1391 1708 1395 1712
rect 1455 1708 1459 1712
rect 1519 1708 1523 1712
rect 1583 1708 1587 1712
rect 1647 1708 1651 1712
rect 1703 1708 1707 1712
rect 1759 1708 1763 1712
rect 1807 1708 1811 1712
rect 1863 1708 1867 1712
rect 1919 1708 1923 1712
rect 1975 1708 1979 1712
rect 279 1692 283 1696
rect 319 1692 323 1696
rect 359 1692 363 1696
rect 399 1692 403 1696
rect 447 1692 451 1696
rect 495 1692 499 1696
rect 543 1692 547 1696
rect 591 1692 595 1696
rect 639 1692 643 1696
rect 687 1692 691 1696
rect 735 1692 739 1696
rect 783 1692 787 1696
rect 839 1692 843 1696
rect 895 1692 899 1696
rect 1303 1692 1307 1696
rect 1343 1692 1347 1696
rect 1383 1692 1387 1696
rect 1423 1692 1427 1696
rect 1463 1692 1467 1696
rect 1503 1692 1507 1696
rect 1559 1692 1563 1696
rect 1623 1692 1627 1696
rect 1687 1692 1691 1696
rect 1751 1692 1755 1696
rect 1807 1692 1811 1696
rect 1863 1692 1867 1696
rect 1919 1692 1923 1696
rect 1975 1692 1979 1696
rect 2031 1692 2035 1696
rect 2087 1692 2091 1696
rect 111 1685 115 1689
rect 1239 1685 1243 1689
rect 1279 1685 1283 1689
rect 2407 1685 2411 1689
rect 111 1668 115 1672
rect 1239 1668 1243 1672
rect 1279 1668 1283 1672
rect 2407 1668 2411 1672
rect 279 1645 283 1649
rect 319 1645 323 1649
rect 359 1645 363 1649
rect 399 1645 403 1649
rect 447 1645 451 1649
rect 495 1645 499 1649
rect 543 1645 547 1649
rect 591 1645 595 1649
rect 639 1645 643 1649
rect 687 1645 691 1649
rect 735 1645 739 1649
rect 783 1645 787 1649
rect 839 1645 843 1649
rect 895 1645 899 1649
rect 1303 1645 1307 1649
rect 1343 1645 1347 1649
rect 1383 1645 1387 1649
rect 1423 1645 1427 1649
rect 1463 1645 1467 1649
rect 1503 1645 1507 1649
rect 1559 1645 1563 1649
rect 1623 1645 1627 1649
rect 1687 1645 1691 1649
rect 1751 1645 1755 1649
rect 1807 1645 1811 1649
rect 1863 1645 1867 1649
rect 1919 1645 1923 1649
rect 1975 1645 1979 1649
rect 2031 1645 2035 1649
rect 2087 1645 2091 1649
rect 135 1611 139 1615
rect 175 1611 179 1615
rect 215 1611 219 1615
rect 255 1611 259 1615
rect 311 1611 315 1615
rect 391 1611 395 1615
rect 471 1611 475 1615
rect 559 1611 563 1615
rect 639 1611 643 1615
rect 719 1611 723 1615
rect 791 1611 795 1615
rect 855 1611 859 1615
rect 919 1611 923 1615
rect 983 1611 987 1615
rect 1047 1611 1051 1615
rect 1303 1611 1307 1615
rect 1343 1611 1347 1615
rect 1383 1611 1387 1615
rect 1423 1611 1427 1615
rect 1463 1611 1467 1615
rect 1503 1611 1507 1615
rect 1559 1611 1563 1615
rect 1631 1611 1635 1615
rect 1703 1611 1707 1615
rect 1783 1611 1787 1615
rect 1855 1611 1859 1615
rect 1927 1611 1931 1615
rect 1999 1611 2003 1615
rect 2063 1611 2067 1615
rect 2127 1611 2131 1615
rect 2191 1611 2195 1615
rect 2255 1611 2259 1615
rect 2319 1611 2323 1615
rect 2359 1611 2363 1615
rect 111 1588 115 1592
rect 1239 1588 1243 1592
rect 1279 1588 1283 1592
rect 2407 1588 2411 1592
rect 111 1571 115 1575
rect 1239 1571 1243 1575
rect 1279 1571 1283 1575
rect 2407 1571 2411 1575
rect 135 1564 139 1568
rect 175 1564 179 1568
rect 215 1564 219 1568
rect 255 1564 259 1568
rect 311 1564 315 1568
rect 391 1564 395 1568
rect 471 1564 475 1568
rect 559 1564 563 1568
rect 639 1564 643 1568
rect 719 1564 723 1568
rect 791 1564 795 1568
rect 855 1564 859 1568
rect 919 1564 923 1568
rect 983 1564 987 1568
rect 1047 1564 1051 1568
rect 1303 1564 1307 1568
rect 1343 1564 1347 1568
rect 1383 1564 1387 1568
rect 1423 1564 1427 1568
rect 1463 1564 1467 1568
rect 1503 1564 1507 1568
rect 1559 1564 1563 1568
rect 1631 1564 1635 1568
rect 1703 1564 1707 1568
rect 1783 1564 1787 1568
rect 1855 1564 1859 1568
rect 1927 1564 1931 1568
rect 1999 1564 2003 1568
rect 2063 1564 2067 1568
rect 2127 1564 2131 1568
rect 2191 1564 2195 1568
rect 2255 1564 2259 1568
rect 2319 1564 2323 1568
rect 2359 1564 2363 1568
rect 151 1548 155 1552
rect 199 1548 203 1552
rect 263 1548 267 1552
rect 343 1548 347 1552
rect 439 1548 443 1552
rect 535 1548 539 1552
rect 639 1548 643 1552
rect 735 1548 739 1552
rect 823 1548 827 1552
rect 903 1548 907 1552
rect 975 1548 979 1552
rect 1047 1548 1051 1552
rect 1119 1548 1123 1552
rect 1191 1548 1195 1552
rect 1471 1552 1475 1556
rect 1623 1552 1627 1556
rect 1759 1552 1763 1556
rect 1871 1552 1875 1556
rect 1967 1552 1971 1556
rect 2055 1552 2059 1556
rect 2127 1552 2131 1556
rect 2191 1552 2195 1556
rect 2255 1552 2259 1556
rect 2319 1552 2323 1556
rect 2359 1552 2363 1556
rect 111 1541 115 1545
rect 1239 1541 1243 1545
rect 1279 1545 1283 1549
rect 2407 1545 2411 1549
rect 111 1524 115 1528
rect 1239 1524 1243 1528
rect 1279 1528 1283 1532
rect 2407 1528 2411 1532
rect 151 1501 155 1505
rect 199 1501 203 1505
rect 263 1501 267 1505
rect 343 1501 347 1505
rect 439 1501 443 1505
rect 535 1501 539 1505
rect 639 1501 643 1505
rect 735 1501 739 1505
rect 823 1501 827 1505
rect 903 1501 907 1505
rect 975 1501 979 1505
rect 1047 1501 1051 1505
rect 1119 1501 1123 1505
rect 1191 1501 1195 1505
rect 1471 1505 1475 1509
rect 1623 1505 1627 1509
rect 1759 1505 1763 1509
rect 1871 1505 1875 1509
rect 1967 1505 1971 1509
rect 2055 1505 2059 1509
rect 2127 1505 2131 1509
rect 2191 1505 2195 1509
rect 2255 1505 2259 1509
rect 2319 1505 2323 1509
rect 2359 1505 2363 1509
rect 319 1467 323 1471
rect 359 1467 363 1471
rect 399 1467 403 1471
rect 447 1467 451 1471
rect 503 1467 507 1471
rect 559 1467 563 1471
rect 615 1467 619 1471
rect 671 1467 675 1471
rect 735 1467 739 1471
rect 799 1467 803 1471
rect 855 1467 859 1471
rect 911 1467 915 1471
rect 967 1467 971 1471
rect 1023 1467 1027 1471
rect 1087 1467 1091 1471
rect 1151 1467 1155 1471
rect 1191 1467 1195 1471
rect 1303 1455 1307 1459
rect 1375 1455 1379 1459
rect 1479 1455 1483 1459
rect 1583 1455 1587 1459
rect 1687 1455 1691 1459
rect 1783 1455 1787 1459
rect 1871 1455 1875 1459
rect 1951 1455 1955 1459
rect 2031 1455 2035 1459
rect 2103 1455 2107 1459
rect 2167 1455 2171 1459
rect 2239 1455 2243 1459
rect 2311 1455 2315 1459
rect 2359 1455 2363 1459
rect 111 1444 115 1448
rect 1239 1444 1243 1448
rect 1279 1432 1283 1436
rect 111 1427 115 1431
rect 2407 1432 2411 1436
rect 1239 1427 1243 1431
rect 319 1420 323 1424
rect 359 1420 363 1424
rect 399 1420 403 1424
rect 447 1420 451 1424
rect 503 1420 507 1424
rect 559 1420 563 1424
rect 615 1420 619 1424
rect 671 1420 675 1424
rect 735 1420 739 1424
rect 799 1420 803 1424
rect 855 1420 859 1424
rect 911 1420 915 1424
rect 967 1420 971 1424
rect 1023 1420 1027 1424
rect 1087 1420 1091 1424
rect 1151 1420 1155 1424
rect 1191 1420 1195 1424
rect 1279 1415 1283 1419
rect 2407 1415 2411 1419
rect 263 1404 267 1408
rect 303 1404 307 1408
rect 343 1404 347 1408
rect 391 1404 395 1408
rect 447 1404 451 1408
rect 503 1404 507 1408
rect 559 1404 563 1408
rect 623 1404 627 1408
rect 687 1404 691 1408
rect 751 1404 755 1408
rect 815 1404 819 1408
rect 879 1404 883 1408
rect 951 1404 955 1408
rect 1023 1404 1027 1408
rect 1303 1408 1307 1412
rect 1375 1408 1379 1412
rect 1479 1408 1483 1412
rect 1583 1408 1587 1412
rect 1687 1408 1691 1412
rect 1783 1408 1787 1412
rect 1871 1408 1875 1412
rect 1951 1408 1955 1412
rect 2031 1408 2035 1412
rect 2103 1408 2107 1412
rect 2167 1408 2171 1412
rect 2239 1408 2243 1412
rect 2311 1408 2315 1412
rect 2359 1408 2363 1412
rect 111 1397 115 1401
rect 1239 1397 1243 1401
rect 1303 1396 1307 1400
rect 1343 1396 1347 1400
rect 1399 1396 1403 1400
rect 1471 1396 1475 1400
rect 1551 1396 1555 1400
rect 1639 1396 1643 1400
rect 1727 1396 1731 1400
rect 1815 1396 1819 1400
rect 1903 1396 1907 1400
rect 1991 1396 1995 1400
rect 2071 1396 2075 1400
rect 2151 1396 2155 1400
rect 2223 1396 2227 1400
rect 2303 1396 2307 1400
rect 2359 1396 2363 1400
rect 1279 1389 1283 1393
rect 2407 1389 2411 1393
rect 111 1380 115 1384
rect 1239 1380 1243 1384
rect 1279 1372 1283 1376
rect 2407 1372 2411 1376
rect 263 1357 267 1361
rect 303 1357 307 1361
rect 343 1357 347 1361
rect 391 1357 395 1361
rect 447 1357 451 1361
rect 503 1357 507 1361
rect 559 1357 563 1361
rect 623 1357 627 1361
rect 687 1357 691 1361
rect 751 1357 755 1361
rect 815 1357 819 1361
rect 879 1357 883 1361
rect 951 1357 955 1361
rect 1023 1357 1027 1361
rect 1303 1349 1307 1353
rect 1343 1349 1347 1353
rect 1399 1349 1403 1353
rect 1471 1349 1475 1353
rect 1551 1349 1555 1353
rect 1639 1349 1643 1353
rect 1727 1349 1731 1353
rect 1815 1349 1819 1353
rect 1903 1349 1907 1353
rect 1991 1349 1995 1353
rect 2071 1349 2075 1353
rect 2151 1349 2155 1353
rect 2223 1349 2227 1353
rect 2303 1349 2307 1353
rect 2359 1349 2363 1353
rect 135 1323 139 1327
rect 175 1323 179 1327
rect 215 1323 219 1327
rect 255 1323 259 1327
rect 327 1323 331 1327
rect 407 1323 411 1327
rect 495 1323 499 1327
rect 583 1323 587 1327
rect 671 1323 675 1327
rect 759 1323 763 1327
rect 839 1323 843 1327
rect 919 1323 923 1327
rect 1007 1323 1011 1327
rect 1095 1323 1099 1327
rect 1447 1315 1451 1319
rect 1487 1315 1491 1319
rect 1527 1315 1531 1319
rect 1567 1315 1571 1319
rect 1615 1315 1619 1319
rect 1671 1315 1675 1319
rect 1719 1315 1723 1319
rect 1775 1315 1779 1319
rect 1831 1315 1835 1319
rect 1903 1315 1907 1319
rect 1983 1315 1987 1319
rect 2071 1315 2075 1319
rect 2167 1315 2171 1319
rect 2271 1315 2275 1319
rect 2359 1315 2363 1319
rect 111 1300 115 1304
rect 1239 1300 1243 1304
rect 1279 1292 1283 1296
rect 2407 1292 2411 1296
rect 111 1283 115 1287
rect 1239 1283 1243 1287
rect 135 1276 139 1280
rect 175 1276 179 1280
rect 215 1276 219 1280
rect 255 1276 259 1280
rect 327 1276 331 1280
rect 407 1276 411 1280
rect 495 1276 499 1280
rect 583 1276 587 1280
rect 671 1276 675 1280
rect 759 1276 763 1280
rect 839 1276 843 1280
rect 919 1276 923 1280
rect 1007 1276 1011 1280
rect 1095 1276 1099 1280
rect 1279 1275 1283 1279
rect 2407 1275 2411 1279
rect 1447 1268 1451 1272
rect 1487 1268 1491 1272
rect 1527 1268 1531 1272
rect 1567 1268 1571 1272
rect 1615 1268 1619 1272
rect 1671 1268 1675 1272
rect 1719 1268 1723 1272
rect 1775 1268 1779 1272
rect 1831 1268 1835 1272
rect 1903 1268 1907 1272
rect 1983 1268 1987 1272
rect 2071 1268 2075 1272
rect 2167 1268 2171 1272
rect 2271 1268 2275 1272
rect 2359 1268 2363 1272
rect 135 1260 139 1264
rect 175 1260 179 1264
rect 247 1260 251 1264
rect 327 1260 331 1264
rect 415 1260 419 1264
rect 503 1260 507 1264
rect 591 1260 595 1264
rect 671 1260 675 1264
rect 743 1260 747 1264
rect 815 1260 819 1264
rect 879 1260 883 1264
rect 943 1260 947 1264
rect 1007 1260 1011 1264
rect 1071 1260 1075 1264
rect 111 1253 115 1257
rect 1239 1253 1243 1257
rect 1511 1252 1515 1256
rect 1551 1252 1555 1256
rect 1591 1252 1595 1256
rect 1631 1252 1635 1256
rect 1671 1252 1675 1256
rect 1711 1252 1715 1256
rect 1751 1252 1755 1256
rect 1791 1252 1795 1256
rect 1839 1252 1843 1256
rect 1903 1252 1907 1256
rect 1967 1252 1971 1256
rect 2039 1252 2043 1256
rect 2119 1252 2123 1256
rect 2207 1252 2211 1256
rect 2295 1252 2299 1256
rect 2359 1252 2363 1256
rect 1279 1245 1283 1249
rect 2407 1245 2411 1249
rect 111 1236 115 1240
rect 1239 1236 1243 1240
rect 1279 1228 1283 1232
rect 2407 1228 2411 1232
rect 135 1213 139 1217
rect 175 1213 179 1217
rect 247 1213 251 1217
rect 327 1213 331 1217
rect 415 1213 419 1217
rect 503 1213 507 1217
rect 591 1213 595 1217
rect 671 1213 675 1217
rect 743 1213 747 1217
rect 815 1213 819 1217
rect 879 1213 883 1217
rect 943 1213 947 1217
rect 1007 1213 1011 1217
rect 1071 1213 1075 1217
rect 1511 1205 1515 1209
rect 1551 1205 1555 1209
rect 1591 1205 1595 1209
rect 1631 1205 1635 1209
rect 1671 1205 1675 1209
rect 1711 1205 1715 1209
rect 1751 1205 1755 1209
rect 1791 1205 1795 1209
rect 1839 1205 1843 1209
rect 1903 1205 1907 1209
rect 1967 1205 1971 1209
rect 2039 1205 2043 1209
rect 2119 1205 2123 1209
rect 2207 1205 2211 1209
rect 2295 1205 2299 1209
rect 2359 1205 2363 1209
rect 135 1175 139 1179
rect 175 1175 179 1179
rect 231 1175 235 1179
rect 303 1175 307 1179
rect 383 1175 387 1179
rect 471 1175 475 1179
rect 559 1175 563 1179
rect 639 1175 643 1179
rect 719 1175 723 1179
rect 799 1175 803 1179
rect 871 1175 875 1179
rect 935 1175 939 1179
rect 991 1175 995 1179
rect 1047 1175 1051 1179
rect 1103 1175 1107 1179
rect 1151 1175 1155 1179
rect 1191 1175 1195 1179
rect 1559 1171 1563 1175
rect 1599 1171 1603 1175
rect 1639 1171 1643 1175
rect 1679 1171 1683 1175
rect 1719 1171 1723 1175
rect 1759 1171 1763 1175
rect 1799 1171 1803 1175
rect 1855 1171 1859 1175
rect 1927 1171 1931 1175
rect 2023 1171 2027 1175
rect 2135 1171 2139 1175
rect 2255 1171 2259 1175
rect 2359 1171 2363 1175
rect 111 1152 115 1156
rect 1239 1152 1243 1156
rect 1279 1148 1283 1152
rect 2407 1148 2411 1152
rect 111 1135 115 1139
rect 1239 1135 1243 1139
rect 135 1128 139 1132
rect 175 1128 179 1132
rect 231 1128 235 1132
rect 303 1128 307 1132
rect 383 1128 387 1132
rect 471 1128 475 1132
rect 559 1128 563 1132
rect 639 1128 643 1132
rect 719 1128 723 1132
rect 799 1128 803 1132
rect 871 1128 875 1132
rect 935 1128 939 1132
rect 991 1128 995 1132
rect 1047 1128 1051 1132
rect 1103 1128 1107 1132
rect 1151 1128 1155 1132
rect 1191 1128 1195 1132
rect 1279 1131 1283 1135
rect 2407 1131 2411 1135
rect 1559 1124 1563 1128
rect 1599 1124 1603 1128
rect 1639 1124 1643 1128
rect 1679 1124 1683 1128
rect 1719 1124 1723 1128
rect 1759 1124 1763 1128
rect 1799 1124 1803 1128
rect 1855 1124 1859 1128
rect 1927 1124 1931 1128
rect 2023 1124 2027 1128
rect 2135 1124 2139 1128
rect 2255 1124 2259 1128
rect 2359 1124 2363 1128
rect 135 1116 139 1120
rect 215 1116 219 1120
rect 303 1116 307 1120
rect 391 1116 395 1120
rect 479 1116 483 1120
rect 559 1116 563 1120
rect 639 1116 643 1120
rect 711 1116 715 1120
rect 775 1116 779 1120
rect 839 1116 843 1120
rect 903 1116 907 1120
rect 959 1116 963 1120
rect 1023 1116 1027 1120
rect 1087 1116 1091 1120
rect 1151 1116 1155 1120
rect 1191 1116 1195 1120
rect 111 1109 115 1113
rect 1239 1109 1243 1113
rect 1535 1104 1539 1108
rect 1599 1104 1603 1108
rect 1663 1104 1667 1108
rect 1727 1104 1731 1108
rect 1791 1104 1795 1108
rect 1855 1104 1859 1108
rect 1911 1104 1915 1108
rect 1967 1104 1971 1108
rect 2023 1104 2027 1108
rect 2079 1104 2083 1108
rect 2135 1104 2139 1108
rect 2191 1104 2195 1108
rect 2255 1104 2259 1108
rect 2319 1104 2323 1108
rect 2359 1104 2363 1108
rect 1279 1097 1283 1101
rect 111 1092 115 1096
rect 2407 1097 2411 1101
rect 1239 1092 1243 1096
rect 1279 1080 1283 1084
rect 2407 1080 2411 1084
rect 135 1069 139 1073
rect 215 1069 219 1073
rect 303 1069 307 1073
rect 391 1069 395 1073
rect 479 1069 483 1073
rect 559 1069 563 1073
rect 639 1069 643 1073
rect 711 1069 715 1073
rect 775 1069 779 1073
rect 839 1069 843 1073
rect 903 1069 907 1073
rect 959 1069 963 1073
rect 1023 1069 1027 1073
rect 1087 1069 1091 1073
rect 1151 1069 1155 1073
rect 1191 1069 1195 1073
rect 1535 1057 1539 1061
rect 1599 1057 1603 1061
rect 1663 1057 1667 1061
rect 1727 1057 1731 1061
rect 1791 1057 1795 1061
rect 1855 1057 1859 1061
rect 1911 1057 1915 1061
rect 1967 1057 1971 1061
rect 2023 1057 2027 1061
rect 2079 1057 2083 1061
rect 2135 1057 2139 1061
rect 2191 1057 2195 1061
rect 2255 1057 2259 1061
rect 2319 1057 2323 1061
rect 2359 1057 2363 1061
rect 199 1035 203 1039
rect 239 1035 243 1039
rect 287 1035 291 1039
rect 343 1035 347 1039
rect 391 1035 395 1039
rect 439 1035 443 1039
rect 487 1035 491 1039
rect 535 1035 539 1039
rect 583 1035 587 1039
rect 631 1035 635 1039
rect 679 1035 683 1039
rect 727 1035 731 1039
rect 783 1035 787 1039
rect 839 1035 843 1039
rect 895 1035 899 1039
rect 959 1035 963 1039
rect 1023 1035 1027 1039
rect 1087 1035 1091 1039
rect 1151 1035 1155 1039
rect 1191 1035 1195 1039
rect 111 1012 115 1016
rect 1239 1012 1243 1016
rect 1503 1015 1507 1019
rect 1623 1015 1627 1019
rect 1735 1015 1739 1019
rect 1831 1015 1835 1019
rect 1919 1015 1923 1019
rect 1999 1015 2003 1019
rect 2071 1015 2075 1019
rect 2143 1015 2147 1019
rect 2207 1015 2211 1019
rect 2279 1015 2283 1019
rect 111 995 115 999
rect 1239 995 1243 999
rect 199 988 203 992
rect 239 988 243 992
rect 287 988 291 992
rect 343 988 347 992
rect 391 988 395 992
rect 439 988 443 992
rect 487 988 491 992
rect 535 988 539 992
rect 583 988 587 992
rect 631 988 635 992
rect 679 988 683 992
rect 727 988 731 992
rect 783 988 787 992
rect 839 988 843 992
rect 895 988 899 992
rect 959 988 963 992
rect 1023 988 1027 992
rect 1087 988 1091 992
rect 1151 988 1155 992
rect 1191 988 1195 992
rect 1279 992 1283 996
rect 2407 992 2411 996
rect 1279 975 1283 979
rect 2407 975 2411 979
rect 295 964 299 968
rect 343 964 347 968
rect 399 964 403 968
rect 471 964 475 968
rect 551 964 555 968
rect 639 964 643 968
rect 727 964 731 968
rect 807 964 811 968
rect 887 964 891 968
rect 959 964 963 968
rect 1023 964 1027 968
rect 1087 964 1091 968
rect 1151 964 1155 968
rect 1191 964 1195 968
rect 1503 968 1507 972
rect 1623 968 1627 972
rect 1735 968 1739 972
rect 1831 968 1835 972
rect 1919 968 1923 972
rect 1999 968 2003 972
rect 2071 968 2075 972
rect 2143 968 2147 972
rect 2207 968 2211 972
rect 2279 968 2283 972
rect 111 957 115 961
rect 1239 957 1243 961
rect 1319 948 1323 952
rect 1359 948 1363 952
rect 1399 948 1403 952
rect 1463 948 1467 952
rect 1543 948 1547 952
rect 1639 948 1643 952
rect 1735 948 1739 952
rect 1839 948 1843 952
rect 1935 948 1939 952
rect 2023 948 2027 952
rect 2103 948 2107 952
rect 2175 948 2179 952
rect 2239 948 2243 952
rect 2311 948 2315 952
rect 2359 948 2363 952
rect 111 940 115 944
rect 1239 940 1243 944
rect 1279 941 1283 945
rect 2407 941 2411 945
rect 1279 924 1283 928
rect 2407 924 2411 928
rect 295 917 299 921
rect 343 917 347 921
rect 399 917 403 921
rect 471 917 475 921
rect 551 917 555 921
rect 639 917 643 921
rect 727 917 731 921
rect 807 917 811 921
rect 887 917 891 921
rect 959 917 963 921
rect 1023 917 1027 921
rect 1087 917 1091 921
rect 1151 917 1155 921
rect 1191 917 1195 921
rect 1319 901 1323 905
rect 1359 901 1363 905
rect 1399 901 1403 905
rect 1463 901 1467 905
rect 1543 901 1547 905
rect 1639 901 1643 905
rect 1735 901 1739 905
rect 1839 901 1843 905
rect 1935 901 1939 905
rect 2023 901 2027 905
rect 2103 901 2107 905
rect 2175 901 2179 905
rect 2239 901 2243 905
rect 2311 901 2315 905
rect 2359 901 2363 905
rect 255 879 259 883
rect 311 879 315 883
rect 375 879 379 883
rect 455 879 459 883
rect 535 879 539 883
rect 623 879 627 883
rect 711 879 715 883
rect 791 879 795 883
rect 863 879 867 883
rect 935 879 939 883
rect 999 879 1003 883
rect 1055 879 1059 883
rect 1119 879 1123 883
rect 1183 879 1187 883
rect 1335 863 1339 867
rect 1375 863 1379 867
rect 1415 863 1419 867
rect 1471 863 1475 867
rect 1535 863 1539 867
rect 1607 863 1611 867
rect 1679 863 1683 867
rect 1751 863 1755 867
rect 1823 863 1827 867
rect 1895 863 1899 867
rect 1959 863 1963 867
rect 2023 863 2027 867
rect 2087 863 2091 867
rect 2143 863 2147 867
rect 2199 863 2203 867
rect 2255 863 2259 867
rect 2319 863 2323 867
rect 2359 863 2363 867
rect 111 856 115 860
rect 1239 856 1243 860
rect 111 839 115 843
rect 1239 839 1243 843
rect 1279 840 1283 844
rect 2407 840 2411 844
rect 255 832 259 836
rect 311 832 315 836
rect 375 832 379 836
rect 455 832 459 836
rect 535 832 539 836
rect 623 832 627 836
rect 711 832 715 836
rect 791 832 795 836
rect 863 832 867 836
rect 935 832 939 836
rect 999 832 1003 836
rect 1055 832 1059 836
rect 1119 832 1123 836
rect 1183 832 1187 836
rect 191 820 195 824
rect 247 820 251 824
rect 311 820 315 824
rect 383 820 387 824
rect 463 820 467 824
rect 543 820 547 824
rect 615 820 619 824
rect 687 820 691 824
rect 751 820 755 824
rect 815 820 819 824
rect 871 820 875 824
rect 927 820 931 824
rect 983 820 987 824
rect 1047 820 1051 824
rect 1279 823 1283 827
rect 2407 823 2411 827
rect 111 813 115 817
rect 1239 813 1243 817
rect 1335 816 1339 820
rect 1375 816 1379 820
rect 1415 816 1419 820
rect 1471 816 1475 820
rect 1535 816 1539 820
rect 1607 816 1611 820
rect 1679 816 1683 820
rect 1751 816 1755 820
rect 1823 816 1827 820
rect 1895 816 1899 820
rect 1959 816 1963 820
rect 2023 816 2027 820
rect 2087 816 2091 820
rect 2143 816 2147 820
rect 2199 816 2203 820
rect 2255 816 2259 820
rect 2319 816 2323 820
rect 2359 816 2363 820
rect 111 796 115 800
rect 1239 796 1243 800
rect 1303 800 1307 804
rect 1343 800 1347 804
rect 1407 800 1411 804
rect 1479 800 1483 804
rect 1551 800 1555 804
rect 1623 800 1627 804
rect 1695 800 1699 804
rect 1759 800 1763 804
rect 1823 800 1827 804
rect 1887 800 1891 804
rect 1951 800 1955 804
rect 2023 800 2027 804
rect 2103 800 2107 804
rect 2191 800 2195 804
rect 2279 800 2283 804
rect 2359 800 2363 804
rect 1279 793 1283 797
rect 2407 793 2411 797
rect 191 773 195 777
rect 247 773 251 777
rect 311 773 315 777
rect 383 773 387 777
rect 463 773 467 777
rect 543 773 547 777
rect 615 773 619 777
rect 687 773 691 777
rect 751 773 755 777
rect 815 773 819 777
rect 871 773 875 777
rect 927 773 931 777
rect 983 773 987 777
rect 1047 773 1051 777
rect 1279 776 1283 780
rect 2407 776 2411 780
rect 1303 753 1307 757
rect 1343 753 1347 757
rect 1407 753 1411 757
rect 1479 753 1483 757
rect 1551 753 1555 757
rect 1623 753 1627 757
rect 1695 753 1699 757
rect 1759 753 1763 757
rect 1823 753 1827 757
rect 1887 753 1891 757
rect 1951 753 1955 757
rect 2023 753 2027 757
rect 2103 753 2107 757
rect 2191 753 2195 757
rect 2279 753 2283 757
rect 2359 753 2363 757
rect 135 743 139 747
rect 175 743 179 747
rect 215 743 219 747
rect 279 743 283 747
rect 351 743 355 747
rect 423 743 427 747
rect 495 743 499 747
rect 559 743 563 747
rect 623 743 627 747
rect 695 743 699 747
rect 783 743 787 747
rect 879 743 883 747
rect 983 743 987 747
rect 1095 743 1099 747
rect 1191 743 1195 747
rect 111 720 115 724
rect 1239 720 1243 724
rect 1303 723 1307 727
rect 1367 723 1371 727
rect 1455 723 1459 727
rect 1535 723 1539 727
rect 1615 723 1619 727
rect 1695 723 1699 727
rect 1775 723 1779 727
rect 1855 723 1859 727
rect 1943 723 1947 727
rect 2031 723 2035 727
rect 2119 723 2123 727
rect 2207 723 2211 727
rect 2295 723 2299 727
rect 2359 723 2363 727
rect 111 703 115 707
rect 1239 703 1243 707
rect 135 696 139 700
rect 175 696 179 700
rect 215 696 219 700
rect 279 696 283 700
rect 351 696 355 700
rect 423 696 427 700
rect 495 696 499 700
rect 559 696 563 700
rect 623 696 627 700
rect 695 696 699 700
rect 783 696 787 700
rect 879 696 883 700
rect 983 696 987 700
rect 1095 696 1099 700
rect 1191 696 1195 700
rect 1279 700 1283 704
rect 2407 700 2411 704
rect 1279 683 1283 687
rect 2407 683 2411 687
rect 135 676 139 680
rect 175 676 179 680
rect 231 676 235 680
rect 287 676 291 680
rect 343 676 347 680
rect 399 676 403 680
rect 455 676 459 680
rect 503 676 507 680
rect 559 676 563 680
rect 623 676 627 680
rect 695 676 699 680
rect 767 676 771 680
rect 839 676 843 680
rect 903 676 907 680
rect 967 676 971 680
rect 1023 676 1027 680
rect 1087 676 1091 680
rect 1151 676 1155 680
rect 1191 676 1195 680
rect 1303 676 1307 680
rect 1367 676 1371 680
rect 1455 676 1459 680
rect 1535 676 1539 680
rect 1615 676 1619 680
rect 1695 676 1699 680
rect 1775 676 1779 680
rect 1855 676 1859 680
rect 1943 676 1947 680
rect 2031 676 2035 680
rect 2119 676 2123 680
rect 2207 676 2211 680
rect 2295 676 2299 680
rect 2359 676 2363 680
rect 111 669 115 673
rect 1239 669 1243 673
rect 1591 664 1595 668
rect 1639 664 1643 668
rect 1687 664 1691 668
rect 1743 664 1747 668
rect 1799 664 1803 668
rect 1871 664 1875 668
rect 1951 664 1955 668
rect 2047 664 2051 668
rect 2151 664 2155 668
rect 2263 664 2267 668
rect 2359 664 2363 668
rect 1279 657 1283 661
rect 111 652 115 656
rect 2407 657 2411 661
rect 1239 652 1243 656
rect 1279 640 1283 644
rect 2407 640 2411 644
rect 135 629 139 633
rect 175 629 179 633
rect 231 629 235 633
rect 287 629 291 633
rect 343 629 347 633
rect 399 629 403 633
rect 455 629 459 633
rect 503 629 507 633
rect 559 629 563 633
rect 623 629 627 633
rect 695 629 699 633
rect 767 629 771 633
rect 839 629 843 633
rect 903 629 907 633
rect 967 629 971 633
rect 1023 629 1027 633
rect 1087 629 1091 633
rect 1151 629 1155 633
rect 1191 629 1195 633
rect 1591 617 1595 621
rect 1639 617 1643 621
rect 1687 617 1691 621
rect 1743 617 1747 621
rect 1799 617 1803 621
rect 1871 617 1875 621
rect 1951 617 1955 621
rect 2047 617 2051 621
rect 2151 617 2155 621
rect 2263 617 2267 621
rect 2359 617 2363 621
rect 135 599 139 603
rect 183 599 187 603
rect 255 599 259 603
rect 327 599 331 603
rect 399 599 403 603
rect 479 599 483 603
rect 559 599 563 603
rect 639 599 643 603
rect 719 599 723 603
rect 799 599 803 603
rect 879 599 883 603
rect 951 599 955 603
rect 1015 599 1019 603
rect 1079 599 1083 603
rect 1143 599 1147 603
rect 1191 599 1195 603
rect 111 576 115 580
rect 1239 576 1243 580
rect 1559 579 1563 583
rect 1599 579 1603 583
rect 1639 579 1643 583
rect 1679 579 1683 583
rect 1719 579 1723 583
rect 1759 579 1763 583
rect 1807 579 1811 583
rect 1855 579 1859 583
rect 1911 579 1915 583
rect 1967 579 1971 583
rect 2031 579 2035 583
rect 2095 579 2099 583
rect 2167 579 2171 583
rect 2239 579 2243 583
rect 2311 579 2315 583
rect 2359 579 2363 583
rect 111 559 115 563
rect 1239 559 1243 563
rect 135 552 139 556
rect 183 552 187 556
rect 255 552 259 556
rect 327 552 331 556
rect 399 552 403 556
rect 479 552 483 556
rect 559 552 563 556
rect 639 552 643 556
rect 719 552 723 556
rect 799 552 803 556
rect 879 552 883 556
rect 951 552 955 556
rect 1015 552 1019 556
rect 1079 552 1083 556
rect 1143 552 1147 556
rect 1191 552 1195 556
rect 1279 556 1283 560
rect 2407 556 2411 560
rect 151 536 155 540
rect 223 536 227 540
rect 287 536 291 540
rect 351 536 355 540
rect 415 536 419 540
rect 479 536 483 540
rect 551 536 555 540
rect 623 536 627 540
rect 695 536 699 540
rect 767 536 771 540
rect 839 536 843 540
rect 919 536 923 540
rect 999 536 1003 540
rect 1079 536 1083 540
rect 1279 539 1283 543
rect 2407 539 2411 543
rect 111 529 115 533
rect 1239 529 1243 533
rect 1559 532 1563 536
rect 1599 532 1603 536
rect 1639 532 1643 536
rect 1679 532 1683 536
rect 1719 532 1723 536
rect 1759 532 1763 536
rect 1807 532 1811 536
rect 1855 532 1859 536
rect 1911 532 1915 536
rect 1967 532 1971 536
rect 2031 532 2035 536
rect 2095 532 2099 536
rect 2167 532 2171 536
rect 2239 532 2243 536
rect 2311 532 2315 536
rect 2359 532 2363 536
rect 1407 520 1411 524
rect 1447 520 1451 524
rect 1487 520 1491 524
rect 1535 520 1539 524
rect 1591 520 1595 524
rect 1647 520 1651 524
rect 1711 520 1715 524
rect 1783 520 1787 524
rect 1863 520 1867 524
rect 1943 520 1947 524
rect 2023 520 2027 524
rect 2103 520 2107 524
rect 2191 520 2195 524
rect 2287 520 2291 524
rect 2359 520 2363 524
rect 111 512 115 516
rect 1239 512 1243 516
rect 1279 513 1283 517
rect 2407 513 2411 517
rect 1279 496 1283 500
rect 2407 496 2411 500
rect 151 489 155 493
rect 223 489 227 493
rect 287 489 291 493
rect 351 489 355 493
rect 415 489 419 493
rect 479 489 483 493
rect 551 489 555 493
rect 623 489 627 493
rect 695 489 699 493
rect 767 489 771 493
rect 839 489 843 493
rect 919 489 923 493
rect 999 489 1003 493
rect 1079 489 1083 493
rect 1407 473 1411 477
rect 1447 473 1451 477
rect 1487 473 1491 477
rect 1535 473 1539 477
rect 1591 473 1595 477
rect 1647 473 1651 477
rect 1711 473 1715 477
rect 1783 473 1787 477
rect 1863 473 1867 477
rect 1943 473 1947 477
rect 2023 473 2027 477
rect 2103 473 2107 477
rect 2191 473 2195 477
rect 2287 473 2291 477
rect 2359 473 2363 477
rect 239 459 243 463
rect 279 459 283 463
rect 327 459 331 463
rect 383 459 387 463
rect 439 459 443 463
rect 503 459 507 463
rect 567 459 571 463
rect 631 459 635 463
rect 695 459 699 463
rect 759 459 763 463
rect 823 459 827 463
rect 887 459 891 463
rect 951 459 955 463
rect 1015 459 1019 463
rect 1303 443 1307 447
rect 1343 443 1347 447
rect 1383 443 1387 447
rect 1447 443 1451 447
rect 1535 443 1539 447
rect 1631 443 1635 447
rect 1735 443 1739 447
rect 1831 443 1835 447
rect 1919 443 1923 447
rect 1999 443 2003 447
rect 2071 443 2075 447
rect 2135 443 2139 447
rect 2199 443 2203 447
rect 2255 443 2259 447
rect 2319 443 2323 447
rect 2359 443 2363 447
rect 111 436 115 440
rect 1239 436 1243 440
rect 111 419 115 423
rect 1239 419 1243 423
rect 1279 420 1283 424
rect 2407 420 2411 424
rect 239 412 243 416
rect 279 412 283 416
rect 327 412 331 416
rect 383 412 387 416
rect 439 412 443 416
rect 503 412 507 416
rect 567 412 571 416
rect 631 412 635 416
rect 695 412 699 416
rect 759 412 763 416
rect 823 412 827 416
rect 887 412 891 416
rect 951 412 955 416
rect 1015 412 1019 416
rect 1279 403 1283 407
rect 2407 403 2411 407
rect 143 396 147 400
rect 183 396 187 400
rect 223 396 227 400
rect 271 396 275 400
rect 335 396 339 400
rect 399 396 403 400
rect 471 396 475 400
rect 543 396 547 400
rect 615 396 619 400
rect 687 396 691 400
rect 751 396 755 400
rect 807 396 811 400
rect 863 396 867 400
rect 919 396 923 400
rect 975 396 979 400
rect 1031 396 1035 400
rect 1303 396 1307 400
rect 1343 396 1347 400
rect 1383 396 1387 400
rect 1447 396 1451 400
rect 1535 396 1539 400
rect 1631 396 1635 400
rect 1735 396 1739 400
rect 1831 396 1835 400
rect 1919 396 1923 400
rect 1999 396 2003 400
rect 2071 396 2075 400
rect 2135 396 2139 400
rect 2199 396 2203 400
rect 2255 396 2259 400
rect 2319 396 2323 400
rect 2359 396 2363 400
rect 111 389 115 393
rect 1239 389 1243 393
rect 1359 384 1363 388
rect 1399 384 1403 388
rect 1439 384 1443 388
rect 1487 384 1491 388
rect 1543 384 1547 388
rect 1607 384 1611 388
rect 1679 384 1683 388
rect 1759 384 1763 388
rect 1839 384 1843 388
rect 1919 384 1923 388
rect 1999 384 2003 388
rect 2079 384 2083 388
rect 2159 384 2163 388
rect 2247 384 2251 388
rect 2335 384 2339 388
rect 1279 377 1283 381
rect 111 372 115 376
rect 2407 377 2411 381
rect 1239 372 1243 376
rect 1279 360 1283 364
rect 2407 360 2411 364
rect 143 349 147 353
rect 183 349 187 353
rect 223 349 227 353
rect 271 349 275 353
rect 335 349 339 353
rect 399 349 403 353
rect 471 349 475 353
rect 543 349 547 353
rect 615 349 619 353
rect 687 349 691 353
rect 751 349 755 353
rect 807 349 811 353
rect 863 349 867 353
rect 919 349 923 353
rect 975 349 979 353
rect 1031 349 1035 353
rect 1359 337 1363 341
rect 1399 337 1403 341
rect 1439 337 1443 341
rect 1487 337 1491 341
rect 1543 337 1547 341
rect 1607 337 1611 341
rect 1679 337 1683 341
rect 1759 337 1763 341
rect 1839 337 1843 341
rect 1919 337 1923 341
rect 1999 337 2003 341
rect 2079 337 2083 341
rect 2159 337 2163 341
rect 2247 337 2251 341
rect 2335 337 2339 341
rect 135 311 139 315
rect 175 311 179 315
rect 215 311 219 315
rect 255 311 259 315
rect 295 311 299 315
rect 335 311 339 315
rect 391 311 395 315
rect 447 311 451 315
rect 495 311 499 315
rect 543 311 547 315
rect 591 311 595 315
rect 639 311 643 315
rect 687 311 691 315
rect 735 311 739 315
rect 783 311 787 315
rect 839 311 843 315
rect 1511 299 1515 303
rect 1551 299 1555 303
rect 1591 299 1595 303
rect 1631 299 1635 303
rect 1671 299 1675 303
rect 1711 299 1715 303
rect 1751 299 1755 303
rect 1791 299 1795 303
rect 1839 299 1843 303
rect 1903 299 1907 303
rect 1967 299 1971 303
rect 2039 299 2043 303
rect 2119 299 2123 303
rect 2199 299 2203 303
rect 2279 299 2283 303
rect 2359 299 2363 303
rect 111 288 115 292
rect 1239 288 1243 292
rect 1279 276 1283 280
rect 111 271 115 275
rect 2407 276 2411 280
rect 1239 271 1243 275
rect 135 264 139 268
rect 175 264 179 268
rect 215 264 219 268
rect 255 264 259 268
rect 295 264 299 268
rect 335 264 339 268
rect 391 264 395 268
rect 447 264 451 268
rect 495 264 499 268
rect 543 264 547 268
rect 591 264 595 268
rect 639 264 643 268
rect 687 264 691 268
rect 735 264 739 268
rect 783 264 787 268
rect 839 264 843 268
rect 1279 259 1283 263
rect 2407 259 2411 263
rect 1511 252 1515 256
rect 1551 252 1555 256
rect 1591 252 1595 256
rect 1631 252 1635 256
rect 1671 252 1675 256
rect 1711 252 1715 256
rect 1751 252 1755 256
rect 1791 252 1795 256
rect 1839 252 1843 256
rect 1903 252 1907 256
rect 1967 252 1971 256
rect 2039 252 2043 256
rect 2119 252 2123 256
rect 2199 252 2203 256
rect 2279 252 2283 256
rect 2359 252 2363 256
rect 135 244 139 248
rect 223 244 227 248
rect 311 244 315 248
rect 391 244 395 248
rect 463 244 467 248
rect 527 244 531 248
rect 591 244 595 248
rect 647 244 651 248
rect 695 244 699 248
rect 735 244 739 248
rect 783 244 787 248
rect 831 244 835 248
rect 879 244 883 248
rect 927 244 931 248
rect 975 244 979 248
rect 1023 244 1027 248
rect 111 237 115 241
rect 1239 237 1243 241
rect 1367 236 1371 240
rect 1407 236 1411 240
rect 1455 236 1459 240
rect 1511 236 1515 240
rect 1567 236 1571 240
rect 1631 236 1635 240
rect 1703 236 1707 240
rect 1775 236 1779 240
rect 1855 236 1859 240
rect 1943 236 1947 240
rect 2031 236 2035 240
rect 2119 236 2123 240
rect 2207 236 2211 240
rect 2295 236 2299 240
rect 2359 236 2363 240
rect 1279 229 1283 233
rect 2407 229 2411 233
rect 111 220 115 224
rect 1239 220 1243 224
rect 1279 212 1283 216
rect 2407 212 2411 216
rect 135 197 139 201
rect 223 197 227 201
rect 311 197 315 201
rect 391 197 395 201
rect 463 197 467 201
rect 527 197 531 201
rect 591 197 595 201
rect 647 197 651 201
rect 695 197 699 201
rect 735 197 739 201
rect 783 197 787 201
rect 831 197 835 201
rect 879 197 883 201
rect 927 197 931 201
rect 975 197 979 201
rect 1023 197 1027 201
rect 1367 189 1371 193
rect 1407 189 1411 193
rect 1455 189 1459 193
rect 1511 189 1515 193
rect 1567 189 1571 193
rect 1631 189 1635 193
rect 1703 189 1707 193
rect 1775 189 1779 193
rect 1855 189 1859 193
rect 1943 189 1947 193
rect 2031 189 2035 193
rect 2119 189 2123 193
rect 2207 189 2211 193
rect 2295 189 2299 193
rect 2359 189 2363 193
rect 1303 151 1307 155
rect 1343 151 1347 155
rect 1383 151 1387 155
rect 1423 151 1427 155
rect 1463 151 1467 155
rect 1519 151 1523 155
rect 1583 151 1587 155
rect 1647 151 1651 155
rect 1711 151 1715 155
rect 1775 151 1779 155
rect 1831 151 1835 155
rect 1887 151 1891 155
rect 1935 151 1939 155
rect 1975 151 1979 155
rect 2015 151 2019 155
rect 2055 151 2059 155
rect 2095 151 2099 155
rect 2143 151 2147 155
rect 2191 151 2195 155
rect 2239 151 2243 155
rect 2279 151 2283 155
rect 2319 151 2323 155
rect 2359 151 2363 155
rect 151 135 155 139
rect 191 135 195 139
rect 231 135 235 139
rect 271 135 275 139
rect 311 135 315 139
rect 351 135 355 139
rect 391 135 395 139
rect 431 135 435 139
rect 471 135 475 139
rect 511 135 515 139
rect 551 135 555 139
rect 591 135 595 139
rect 631 135 635 139
rect 671 135 675 139
rect 711 135 715 139
rect 751 135 755 139
rect 791 135 795 139
rect 831 135 835 139
rect 871 135 875 139
rect 911 135 915 139
rect 951 135 955 139
rect 991 135 995 139
rect 1031 135 1035 139
rect 1071 135 1075 139
rect 1111 135 1115 139
rect 1151 135 1155 139
rect 1191 135 1195 139
rect 1279 128 1283 132
rect 2407 128 2411 132
rect 111 112 115 116
rect 1239 112 1243 116
rect 1279 111 1283 115
rect 2407 111 2411 115
rect 1303 104 1307 108
rect 1343 104 1347 108
rect 1383 104 1387 108
rect 1423 104 1427 108
rect 1463 104 1467 108
rect 1519 104 1523 108
rect 1583 104 1587 108
rect 1647 104 1651 108
rect 1711 104 1715 108
rect 1775 104 1779 108
rect 1831 104 1835 108
rect 1887 104 1891 108
rect 1935 104 1939 108
rect 1975 104 1979 108
rect 2015 104 2019 108
rect 2055 104 2059 108
rect 2095 104 2099 108
rect 2143 104 2147 108
rect 2191 104 2195 108
rect 2239 104 2243 108
rect 2279 104 2283 108
rect 2319 104 2323 108
rect 2359 104 2363 108
rect 111 95 115 99
rect 1239 95 1243 99
rect 151 88 155 92
rect 191 88 195 92
rect 231 88 235 92
rect 271 88 275 92
rect 311 88 315 92
rect 351 88 355 92
rect 391 88 395 92
rect 431 88 435 92
rect 471 88 475 92
rect 511 88 515 92
rect 551 88 555 92
rect 591 88 595 92
rect 631 88 635 92
rect 671 88 675 92
rect 711 88 715 92
rect 751 88 755 92
rect 791 88 795 92
rect 831 88 835 92
rect 871 88 875 92
rect 911 88 915 92
rect 951 88 955 92
rect 991 88 995 92
rect 1031 88 1035 92
rect 1071 88 1075 92
rect 1111 88 1115 92
rect 1151 88 1155 92
rect 1191 88 1195 92
<< m3 >>
rect 111 2494 115 2495
rect 111 2489 115 2490
rect 231 2494 235 2495
rect 231 2489 235 2490
rect 271 2494 275 2495
rect 271 2489 275 2490
rect 311 2494 315 2495
rect 311 2489 315 2490
rect 351 2494 355 2495
rect 351 2489 355 2490
rect 399 2494 403 2495
rect 399 2489 403 2490
rect 455 2494 459 2495
rect 455 2489 459 2490
rect 511 2494 515 2495
rect 511 2489 515 2490
rect 575 2494 579 2495
rect 575 2489 579 2490
rect 639 2494 643 2495
rect 639 2489 643 2490
rect 703 2494 707 2495
rect 703 2489 707 2490
rect 767 2494 771 2495
rect 767 2489 771 2490
rect 823 2494 827 2495
rect 823 2489 827 2490
rect 879 2494 883 2495
rect 879 2489 883 2490
rect 927 2494 931 2495
rect 927 2489 931 2490
rect 975 2494 979 2495
rect 975 2489 979 2490
rect 1023 2494 1027 2495
rect 1023 2489 1027 2490
rect 1071 2494 1075 2495
rect 1071 2489 1075 2490
rect 1111 2494 1115 2495
rect 1111 2489 1115 2490
rect 1151 2494 1155 2495
rect 1151 2489 1155 2490
rect 1191 2494 1195 2495
rect 1191 2489 1195 2490
rect 1239 2494 1243 2495
rect 1239 2489 1243 2490
rect 1279 2490 1283 2491
rect 112 2457 114 2489
rect 232 2480 234 2489
rect 272 2480 274 2489
rect 312 2480 314 2489
rect 352 2480 354 2489
rect 400 2480 402 2489
rect 456 2480 458 2489
rect 512 2480 514 2489
rect 576 2480 578 2489
rect 640 2480 642 2489
rect 704 2480 706 2489
rect 768 2480 770 2489
rect 824 2480 826 2489
rect 880 2480 882 2489
rect 928 2480 930 2489
rect 976 2480 978 2489
rect 1024 2480 1026 2489
rect 1072 2480 1074 2489
rect 1112 2480 1114 2489
rect 1152 2480 1154 2489
rect 1192 2480 1194 2489
rect 230 2479 236 2480
rect 230 2475 231 2479
rect 235 2475 236 2479
rect 230 2474 236 2475
rect 270 2479 276 2480
rect 270 2475 271 2479
rect 275 2475 276 2479
rect 270 2474 276 2475
rect 310 2479 316 2480
rect 310 2475 311 2479
rect 315 2475 316 2479
rect 310 2474 316 2475
rect 350 2479 356 2480
rect 350 2475 351 2479
rect 355 2475 356 2479
rect 350 2474 356 2475
rect 398 2479 404 2480
rect 398 2475 399 2479
rect 403 2475 404 2479
rect 398 2474 404 2475
rect 454 2479 460 2480
rect 454 2475 455 2479
rect 459 2475 460 2479
rect 454 2474 460 2475
rect 510 2479 516 2480
rect 510 2475 511 2479
rect 515 2475 516 2479
rect 510 2474 516 2475
rect 574 2479 580 2480
rect 574 2475 575 2479
rect 579 2475 580 2479
rect 574 2474 580 2475
rect 638 2479 644 2480
rect 638 2475 639 2479
rect 643 2475 644 2479
rect 638 2474 644 2475
rect 702 2479 708 2480
rect 702 2475 703 2479
rect 707 2475 708 2479
rect 702 2474 708 2475
rect 766 2479 772 2480
rect 766 2475 767 2479
rect 771 2475 772 2479
rect 766 2474 772 2475
rect 822 2479 828 2480
rect 822 2475 823 2479
rect 827 2475 828 2479
rect 822 2474 828 2475
rect 878 2479 884 2480
rect 878 2475 879 2479
rect 883 2475 884 2479
rect 878 2474 884 2475
rect 926 2479 932 2480
rect 926 2475 927 2479
rect 931 2475 932 2479
rect 926 2474 932 2475
rect 974 2479 980 2480
rect 974 2475 975 2479
rect 979 2475 980 2479
rect 974 2474 980 2475
rect 1022 2479 1028 2480
rect 1022 2475 1023 2479
rect 1027 2475 1028 2479
rect 1022 2474 1028 2475
rect 1070 2479 1076 2480
rect 1070 2475 1071 2479
rect 1075 2475 1076 2479
rect 1070 2474 1076 2475
rect 1110 2479 1116 2480
rect 1110 2475 1111 2479
rect 1115 2475 1116 2479
rect 1110 2474 1116 2475
rect 1150 2479 1156 2480
rect 1150 2475 1151 2479
rect 1155 2475 1156 2479
rect 1150 2474 1156 2475
rect 1190 2479 1196 2480
rect 1190 2475 1191 2479
rect 1195 2475 1196 2479
rect 1190 2474 1196 2475
rect 1240 2457 1242 2489
rect 1279 2485 1283 2486
rect 1303 2490 1307 2491
rect 1303 2485 1307 2486
rect 1343 2490 1347 2491
rect 1343 2485 1347 2486
rect 1383 2490 1387 2491
rect 1383 2485 1387 2486
rect 1439 2490 1443 2491
rect 1439 2485 1443 2486
rect 1511 2490 1515 2491
rect 1511 2485 1515 2486
rect 1583 2490 1587 2491
rect 1583 2485 1587 2486
rect 1663 2490 1667 2491
rect 1663 2485 1667 2486
rect 1735 2490 1739 2491
rect 1735 2485 1739 2486
rect 1807 2490 1811 2491
rect 1807 2485 1811 2486
rect 1887 2490 1891 2491
rect 1887 2485 1891 2486
rect 1967 2490 1971 2491
rect 1967 2485 1971 2486
rect 2063 2490 2067 2491
rect 2063 2485 2067 2486
rect 2167 2490 2171 2491
rect 2167 2485 2171 2486
rect 2271 2490 2275 2491
rect 2271 2485 2275 2486
rect 2359 2490 2363 2491
rect 2359 2485 2363 2486
rect 2407 2490 2411 2491
rect 2407 2485 2411 2486
rect 110 2456 116 2457
rect 110 2452 111 2456
rect 115 2452 116 2456
rect 110 2451 116 2452
rect 1238 2456 1244 2457
rect 1238 2452 1239 2456
rect 1243 2452 1244 2456
rect 1280 2453 1282 2485
rect 1304 2476 1306 2485
rect 1344 2476 1346 2485
rect 1384 2476 1386 2485
rect 1440 2476 1442 2485
rect 1512 2476 1514 2485
rect 1584 2476 1586 2485
rect 1664 2476 1666 2485
rect 1736 2476 1738 2485
rect 1808 2476 1810 2485
rect 1888 2476 1890 2485
rect 1968 2476 1970 2485
rect 2064 2476 2066 2485
rect 2168 2476 2170 2485
rect 2272 2476 2274 2485
rect 2360 2476 2362 2485
rect 1302 2475 1308 2476
rect 1302 2471 1303 2475
rect 1307 2471 1308 2475
rect 1302 2470 1308 2471
rect 1342 2475 1348 2476
rect 1342 2471 1343 2475
rect 1347 2471 1348 2475
rect 1342 2470 1348 2471
rect 1382 2475 1388 2476
rect 1382 2471 1383 2475
rect 1387 2471 1388 2475
rect 1382 2470 1388 2471
rect 1438 2475 1444 2476
rect 1438 2471 1439 2475
rect 1443 2471 1444 2475
rect 1438 2470 1444 2471
rect 1510 2475 1516 2476
rect 1510 2471 1511 2475
rect 1515 2471 1516 2475
rect 1510 2470 1516 2471
rect 1582 2475 1588 2476
rect 1582 2471 1583 2475
rect 1587 2471 1588 2475
rect 1582 2470 1588 2471
rect 1662 2475 1668 2476
rect 1662 2471 1663 2475
rect 1667 2471 1668 2475
rect 1662 2470 1668 2471
rect 1734 2475 1740 2476
rect 1734 2471 1735 2475
rect 1739 2471 1740 2475
rect 1734 2470 1740 2471
rect 1806 2475 1812 2476
rect 1806 2471 1807 2475
rect 1811 2471 1812 2475
rect 1806 2470 1812 2471
rect 1886 2475 1892 2476
rect 1886 2471 1887 2475
rect 1891 2471 1892 2475
rect 1886 2470 1892 2471
rect 1966 2475 1972 2476
rect 1966 2471 1967 2475
rect 1971 2471 1972 2475
rect 1966 2470 1972 2471
rect 2062 2475 2068 2476
rect 2062 2471 2063 2475
rect 2067 2471 2068 2475
rect 2062 2470 2068 2471
rect 2166 2475 2172 2476
rect 2166 2471 2167 2475
rect 2171 2471 2172 2475
rect 2166 2470 2172 2471
rect 2270 2475 2276 2476
rect 2270 2471 2271 2475
rect 2275 2471 2276 2475
rect 2270 2470 2276 2471
rect 2358 2475 2364 2476
rect 2358 2471 2359 2475
rect 2363 2471 2364 2475
rect 2358 2470 2364 2471
rect 2408 2453 2410 2485
rect 1238 2451 1244 2452
rect 1278 2452 1284 2453
rect 1278 2448 1279 2452
rect 1283 2448 1284 2452
rect 1278 2447 1284 2448
rect 2406 2452 2412 2453
rect 2406 2448 2407 2452
rect 2411 2448 2412 2452
rect 2406 2447 2412 2448
rect 110 2439 116 2440
rect 110 2435 111 2439
rect 115 2435 116 2439
rect 110 2434 116 2435
rect 1238 2439 1244 2440
rect 1238 2435 1239 2439
rect 1243 2435 1244 2439
rect 1238 2434 1244 2435
rect 1278 2435 1284 2436
rect 112 2419 114 2434
rect 230 2432 236 2433
rect 230 2428 231 2432
rect 235 2428 236 2432
rect 230 2427 236 2428
rect 270 2432 276 2433
rect 270 2428 271 2432
rect 275 2428 276 2432
rect 270 2427 276 2428
rect 310 2432 316 2433
rect 310 2428 311 2432
rect 315 2428 316 2432
rect 310 2427 316 2428
rect 350 2432 356 2433
rect 350 2428 351 2432
rect 355 2428 356 2432
rect 350 2427 356 2428
rect 398 2432 404 2433
rect 398 2428 399 2432
rect 403 2428 404 2432
rect 398 2427 404 2428
rect 454 2432 460 2433
rect 454 2428 455 2432
rect 459 2428 460 2432
rect 454 2427 460 2428
rect 510 2432 516 2433
rect 510 2428 511 2432
rect 515 2428 516 2432
rect 510 2427 516 2428
rect 574 2432 580 2433
rect 574 2428 575 2432
rect 579 2428 580 2432
rect 574 2427 580 2428
rect 638 2432 644 2433
rect 638 2428 639 2432
rect 643 2428 644 2432
rect 638 2427 644 2428
rect 702 2432 708 2433
rect 702 2428 703 2432
rect 707 2428 708 2432
rect 702 2427 708 2428
rect 766 2432 772 2433
rect 766 2428 767 2432
rect 771 2428 772 2432
rect 766 2427 772 2428
rect 822 2432 828 2433
rect 822 2428 823 2432
rect 827 2428 828 2432
rect 822 2427 828 2428
rect 878 2432 884 2433
rect 878 2428 879 2432
rect 883 2428 884 2432
rect 878 2427 884 2428
rect 926 2432 932 2433
rect 926 2428 927 2432
rect 931 2428 932 2432
rect 926 2427 932 2428
rect 974 2432 980 2433
rect 974 2428 975 2432
rect 979 2428 980 2432
rect 974 2427 980 2428
rect 1022 2432 1028 2433
rect 1022 2428 1023 2432
rect 1027 2428 1028 2432
rect 1022 2427 1028 2428
rect 1070 2432 1076 2433
rect 1070 2428 1071 2432
rect 1075 2428 1076 2432
rect 1070 2427 1076 2428
rect 1110 2432 1116 2433
rect 1110 2428 1111 2432
rect 1115 2428 1116 2432
rect 1110 2427 1116 2428
rect 1150 2432 1156 2433
rect 1150 2428 1151 2432
rect 1155 2428 1156 2432
rect 1150 2427 1156 2428
rect 1190 2432 1196 2433
rect 1190 2428 1191 2432
rect 1195 2428 1196 2432
rect 1190 2427 1196 2428
rect 232 2419 234 2427
rect 272 2419 274 2427
rect 312 2419 314 2427
rect 352 2419 354 2427
rect 400 2419 402 2427
rect 456 2419 458 2427
rect 512 2419 514 2427
rect 576 2419 578 2427
rect 640 2419 642 2427
rect 704 2419 706 2427
rect 768 2419 770 2427
rect 824 2419 826 2427
rect 880 2419 882 2427
rect 928 2419 930 2427
rect 976 2419 978 2427
rect 1024 2419 1026 2427
rect 1072 2419 1074 2427
rect 1112 2419 1114 2427
rect 1152 2419 1154 2427
rect 1192 2419 1194 2427
rect 1240 2419 1242 2434
rect 1278 2431 1279 2435
rect 1283 2431 1284 2435
rect 1278 2430 1284 2431
rect 2406 2435 2412 2436
rect 2406 2431 2407 2435
rect 2411 2431 2412 2435
rect 2406 2430 2412 2431
rect 1280 2423 1282 2430
rect 1302 2428 1308 2429
rect 1302 2424 1303 2428
rect 1307 2424 1308 2428
rect 1302 2423 1308 2424
rect 1342 2428 1348 2429
rect 1342 2424 1343 2428
rect 1347 2424 1348 2428
rect 1342 2423 1348 2424
rect 1382 2428 1388 2429
rect 1382 2424 1383 2428
rect 1387 2424 1388 2428
rect 1382 2423 1388 2424
rect 1438 2428 1444 2429
rect 1438 2424 1439 2428
rect 1443 2424 1444 2428
rect 1438 2423 1444 2424
rect 1510 2428 1516 2429
rect 1510 2424 1511 2428
rect 1515 2424 1516 2428
rect 1510 2423 1516 2424
rect 1582 2428 1588 2429
rect 1582 2424 1583 2428
rect 1587 2424 1588 2428
rect 1582 2423 1588 2424
rect 1662 2428 1668 2429
rect 1662 2424 1663 2428
rect 1667 2424 1668 2428
rect 1662 2423 1668 2424
rect 1734 2428 1740 2429
rect 1734 2424 1735 2428
rect 1739 2424 1740 2428
rect 1734 2423 1740 2424
rect 1806 2428 1812 2429
rect 1806 2424 1807 2428
rect 1811 2424 1812 2428
rect 1806 2423 1812 2424
rect 1886 2428 1892 2429
rect 1886 2424 1887 2428
rect 1891 2424 1892 2428
rect 1886 2423 1892 2424
rect 1966 2428 1972 2429
rect 1966 2424 1967 2428
rect 1971 2424 1972 2428
rect 1966 2423 1972 2424
rect 2062 2428 2068 2429
rect 2062 2424 2063 2428
rect 2067 2424 2068 2428
rect 2062 2423 2068 2424
rect 2166 2428 2172 2429
rect 2166 2424 2167 2428
rect 2171 2424 2172 2428
rect 2166 2423 2172 2424
rect 2270 2428 2276 2429
rect 2270 2424 2271 2428
rect 2275 2424 2276 2428
rect 2270 2423 2276 2424
rect 2358 2428 2364 2429
rect 2358 2424 2359 2428
rect 2363 2424 2364 2428
rect 2358 2423 2364 2424
rect 2408 2423 2410 2430
rect 1279 2422 1283 2423
rect 111 2418 115 2419
rect 111 2413 115 2414
rect 199 2418 203 2419
rect 199 2413 203 2414
rect 231 2418 235 2419
rect 231 2413 235 2414
rect 263 2418 267 2419
rect 263 2413 267 2414
rect 271 2418 275 2419
rect 271 2413 275 2414
rect 311 2418 315 2419
rect 311 2413 315 2414
rect 327 2418 331 2419
rect 327 2413 331 2414
rect 351 2418 355 2419
rect 351 2413 355 2414
rect 399 2418 403 2419
rect 399 2413 403 2414
rect 455 2418 459 2419
rect 455 2413 459 2414
rect 471 2418 475 2419
rect 471 2413 475 2414
rect 511 2418 515 2419
rect 511 2413 515 2414
rect 543 2418 547 2419
rect 543 2413 547 2414
rect 575 2418 579 2419
rect 575 2413 579 2414
rect 615 2418 619 2419
rect 615 2413 619 2414
rect 639 2418 643 2419
rect 639 2413 643 2414
rect 687 2418 691 2419
rect 687 2413 691 2414
rect 703 2418 707 2419
rect 703 2413 707 2414
rect 751 2418 755 2419
rect 751 2413 755 2414
rect 767 2418 771 2419
rect 767 2413 771 2414
rect 823 2418 827 2419
rect 823 2413 827 2414
rect 879 2418 883 2419
rect 879 2413 883 2414
rect 895 2418 899 2419
rect 895 2413 899 2414
rect 927 2418 931 2419
rect 927 2413 931 2414
rect 967 2418 971 2419
rect 967 2413 971 2414
rect 975 2418 979 2419
rect 975 2413 979 2414
rect 1023 2418 1027 2419
rect 1023 2413 1027 2414
rect 1071 2418 1075 2419
rect 1071 2413 1075 2414
rect 1111 2418 1115 2419
rect 1111 2413 1115 2414
rect 1151 2418 1155 2419
rect 1151 2413 1155 2414
rect 1191 2418 1195 2419
rect 1191 2413 1195 2414
rect 1239 2418 1243 2419
rect 1279 2417 1283 2418
rect 1303 2422 1307 2423
rect 1303 2417 1307 2418
rect 1343 2422 1347 2423
rect 1343 2417 1347 2418
rect 1375 2422 1379 2423
rect 1375 2417 1379 2418
rect 1383 2422 1387 2423
rect 1383 2417 1387 2418
rect 1415 2422 1419 2423
rect 1415 2417 1419 2418
rect 1439 2422 1443 2423
rect 1439 2417 1443 2418
rect 1455 2422 1459 2423
rect 1455 2417 1459 2418
rect 1503 2422 1507 2423
rect 1503 2417 1507 2418
rect 1511 2422 1515 2423
rect 1511 2417 1515 2418
rect 1559 2422 1563 2423
rect 1559 2417 1563 2418
rect 1583 2422 1587 2423
rect 1583 2417 1587 2418
rect 1615 2422 1619 2423
rect 1615 2417 1619 2418
rect 1663 2422 1667 2423
rect 1663 2417 1667 2418
rect 1679 2422 1683 2423
rect 1679 2417 1683 2418
rect 1735 2422 1739 2423
rect 1735 2417 1739 2418
rect 1799 2422 1803 2423
rect 1799 2417 1803 2418
rect 1807 2422 1811 2423
rect 1807 2417 1811 2418
rect 1871 2422 1875 2423
rect 1871 2417 1875 2418
rect 1887 2422 1891 2423
rect 1887 2417 1891 2418
rect 1951 2422 1955 2423
rect 1951 2417 1955 2418
rect 1967 2422 1971 2423
rect 1967 2417 1971 2418
rect 2047 2422 2051 2423
rect 2047 2417 2051 2418
rect 2063 2422 2067 2423
rect 2063 2417 2067 2418
rect 2151 2422 2155 2423
rect 2151 2417 2155 2418
rect 2167 2422 2171 2423
rect 2167 2417 2171 2418
rect 2263 2422 2267 2423
rect 2263 2417 2267 2418
rect 2271 2422 2275 2423
rect 2271 2417 2275 2418
rect 2359 2422 2363 2423
rect 2359 2417 2363 2418
rect 2407 2422 2411 2423
rect 2407 2417 2411 2418
rect 1239 2413 1243 2414
rect 112 2406 114 2413
rect 198 2412 204 2413
rect 198 2408 199 2412
rect 203 2408 204 2412
rect 198 2407 204 2408
rect 262 2412 268 2413
rect 262 2408 263 2412
rect 267 2408 268 2412
rect 262 2407 268 2408
rect 326 2412 332 2413
rect 326 2408 327 2412
rect 331 2408 332 2412
rect 326 2407 332 2408
rect 398 2412 404 2413
rect 398 2408 399 2412
rect 403 2408 404 2412
rect 398 2407 404 2408
rect 470 2412 476 2413
rect 470 2408 471 2412
rect 475 2408 476 2412
rect 470 2407 476 2408
rect 542 2412 548 2413
rect 542 2408 543 2412
rect 547 2408 548 2412
rect 542 2407 548 2408
rect 614 2412 620 2413
rect 614 2408 615 2412
rect 619 2408 620 2412
rect 614 2407 620 2408
rect 686 2412 692 2413
rect 686 2408 687 2412
rect 691 2408 692 2412
rect 686 2407 692 2408
rect 750 2412 756 2413
rect 750 2408 751 2412
rect 755 2408 756 2412
rect 750 2407 756 2408
rect 822 2412 828 2413
rect 822 2408 823 2412
rect 827 2408 828 2412
rect 822 2407 828 2408
rect 894 2412 900 2413
rect 894 2408 895 2412
rect 899 2408 900 2412
rect 894 2407 900 2408
rect 966 2412 972 2413
rect 966 2408 967 2412
rect 971 2408 972 2412
rect 966 2407 972 2408
rect 1240 2406 1242 2413
rect 1280 2410 1282 2417
rect 1374 2416 1380 2417
rect 1374 2412 1375 2416
rect 1379 2412 1380 2416
rect 1374 2411 1380 2412
rect 1414 2416 1420 2417
rect 1414 2412 1415 2416
rect 1419 2412 1420 2416
rect 1414 2411 1420 2412
rect 1454 2416 1460 2417
rect 1454 2412 1455 2416
rect 1459 2412 1460 2416
rect 1454 2411 1460 2412
rect 1502 2416 1508 2417
rect 1502 2412 1503 2416
rect 1507 2412 1508 2416
rect 1502 2411 1508 2412
rect 1558 2416 1564 2417
rect 1558 2412 1559 2416
rect 1563 2412 1564 2416
rect 1558 2411 1564 2412
rect 1614 2416 1620 2417
rect 1614 2412 1615 2416
rect 1619 2412 1620 2416
rect 1614 2411 1620 2412
rect 1678 2416 1684 2417
rect 1678 2412 1679 2416
rect 1683 2412 1684 2416
rect 1678 2411 1684 2412
rect 1734 2416 1740 2417
rect 1734 2412 1735 2416
rect 1739 2412 1740 2416
rect 1734 2411 1740 2412
rect 1798 2416 1804 2417
rect 1798 2412 1799 2416
rect 1803 2412 1804 2416
rect 1798 2411 1804 2412
rect 1870 2416 1876 2417
rect 1870 2412 1871 2416
rect 1875 2412 1876 2416
rect 1870 2411 1876 2412
rect 1950 2416 1956 2417
rect 1950 2412 1951 2416
rect 1955 2412 1956 2416
rect 1950 2411 1956 2412
rect 2046 2416 2052 2417
rect 2046 2412 2047 2416
rect 2051 2412 2052 2416
rect 2046 2411 2052 2412
rect 2150 2416 2156 2417
rect 2150 2412 2151 2416
rect 2155 2412 2156 2416
rect 2150 2411 2156 2412
rect 2262 2416 2268 2417
rect 2262 2412 2263 2416
rect 2267 2412 2268 2416
rect 2262 2411 2268 2412
rect 2358 2416 2364 2417
rect 2358 2412 2359 2416
rect 2363 2412 2364 2416
rect 2358 2411 2364 2412
rect 2408 2410 2410 2417
rect 1278 2409 1284 2410
rect 110 2405 116 2406
rect 110 2401 111 2405
rect 115 2401 116 2405
rect 110 2400 116 2401
rect 1238 2405 1244 2406
rect 1238 2401 1239 2405
rect 1243 2401 1244 2405
rect 1278 2405 1279 2409
rect 1283 2405 1284 2409
rect 1278 2404 1284 2405
rect 2406 2409 2412 2410
rect 2406 2405 2407 2409
rect 2411 2405 2412 2409
rect 2406 2404 2412 2405
rect 1238 2400 1244 2401
rect 1278 2392 1284 2393
rect 110 2388 116 2389
rect 110 2384 111 2388
rect 115 2384 116 2388
rect 110 2383 116 2384
rect 1238 2388 1244 2389
rect 1238 2384 1239 2388
rect 1243 2384 1244 2388
rect 1278 2388 1279 2392
rect 1283 2388 1284 2392
rect 1278 2387 1284 2388
rect 2406 2392 2412 2393
rect 2406 2388 2407 2392
rect 2411 2388 2412 2392
rect 2406 2387 2412 2388
rect 1238 2383 1244 2384
rect 112 2347 114 2383
rect 198 2365 204 2366
rect 198 2361 199 2365
rect 203 2361 204 2365
rect 198 2360 204 2361
rect 262 2365 268 2366
rect 262 2361 263 2365
rect 267 2361 268 2365
rect 262 2360 268 2361
rect 326 2365 332 2366
rect 326 2361 327 2365
rect 331 2361 332 2365
rect 326 2360 332 2361
rect 398 2365 404 2366
rect 398 2361 399 2365
rect 403 2361 404 2365
rect 398 2360 404 2361
rect 470 2365 476 2366
rect 470 2361 471 2365
rect 475 2361 476 2365
rect 470 2360 476 2361
rect 542 2365 548 2366
rect 542 2361 543 2365
rect 547 2361 548 2365
rect 542 2360 548 2361
rect 614 2365 620 2366
rect 614 2361 615 2365
rect 619 2361 620 2365
rect 614 2360 620 2361
rect 686 2365 692 2366
rect 686 2361 687 2365
rect 691 2361 692 2365
rect 686 2360 692 2361
rect 750 2365 756 2366
rect 750 2361 751 2365
rect 755 2361 756 2365
rect 750 2360 756 2361
rect 822 2365 828 2366
rect 822 2361 823 2365
rect 827 2361 828 2365
rect 822 2360 828 2361
rect 894 2365 900 2366
rect 894 2361 895 2365
rect 899 2361 900 2365
rect 894 2360 900 2361
rect 966 2365 972 2366
rect 966 2361 967 2365
rect 971 2361 972 2365
rect 966 2360 972 2361
rect 200 2347 202 2360
rect 264 2347 266 2360
rect 328 2347 330 2360
rect 400 2347 402 2360
rect 472 2347 474 2360
rect 544 2347 546 2360
rect 616 2347 618 2360
rect 688 2347 690 2360
rect 752 2347 754 2360
rect 824 2347 826 2360
rect 896 2347 898 2360
rect 968 2347 970 2360
rect 1240 2347 1242 2383
rect 1280 2351 1282 2387
rect 1374 2369 1380 2370
rect 1374 2365 1375 2369
rect 1379 2365 1380 2369
rect 1374 2364 1380 2365
rect 1414 2369 1420 2370
rect 1414 2365 1415 2369
rect 1419 2365 1420 2369
rect 1414 2364 1420 2365
rect 1454 2369 1460 2370
rect 1454 2365 1455 2369
rect 1459 2365 1460 2369
rect 1454 2364 1460 2365
rect 1502 2369 1508 2370
rect 1502 2365 1503 2369
rect 1507 2365 1508 2369
rect 1502 2364 1508 2365
rect 1558 2369 1564 2370
rect 1558 2365 1559 2369
rect 1563 2365 1564 2369
rect 1558 2364 1564 2365
rect 1614 2369 1620 2370
rect 1614 2365 1615 2369
rect 1619 2365 1620 2369
rect 1614 2364 1620 2365
rect 1678 2369 1684 2370
rect 1678 2365 1679 2369
rect 1683 2365 1684 2369
rect 1678 2364 1684 2365
rect 1734 2369 1740 2370
rect 1734 2365 1735 2369
rect 1739 2365 1740 2369
rect 1734 2364 1740 2365
rect 1798 2369 1804 2370
rect 1798 2365 1799 2369
rect 1803 2365 1804 2369
rect 1798 2364 1804 2365
rect 1870 2369 1876 2370
rect 1870 2365 1871 2369
rect 1875 2365 1876 2369
rect 1870 2364 1876 2365
rect 1950 2369 1956 2370
rect 1950 2365 1951 2369
rect 1955 2365 1956 2369
rect 1950 2364 1956 2365
rect 2046 2369 2052 2370
rect 2046 2365 2047 2369
rect 2051 2365 2052 2369
rect 2046 2364 2052 2365
rect 2150 2369 2156 2370
rect 2150 2365 2151 2369
rect 2155 2365 2156 2369
rect 2150 2364 2156 2365
rect 2262 2369 2268 2370
rect 2262 2365 2263 2369
rect 2267 2365 2268 2369
rect 2262 2364 2268 2365
rect 2358 2369 2364 2370
rect 2358 2365 2359 2369
rect 2363 2365 2364 2369
rect 2358 2364 2364 2365
rect 1376 2351 1378 2364
rect 1416 2351 1418 2364
rect 1456 2351 1458 2364
rect 1504 2351 1506 2364
rect 1560 2351 1562 2364
rect 1616 2351 1618 2364
rect 1680 2351 1682 2364
rect 1736 2351 1738 2364
rect 1800 2351 1802 2364
rect 1872 2351 1874 2364
rect 1952 2351 1954 2364
rect 2048 2351 2050 2364
rect 2152 2351 2154 2364
rect 2264 2351 2266 2364
rect 2360 2351 2362 2364
rect 2408 2351 2410 2387
rect 1279 2350 1283 2351
rect 111 2346 115 2347
rect 111 2341 115 2342
rect 199 2346 203 2347
rect 199 2341 203 2342
rect 263 2346 267 2347
rect 263 2341 267 2342
rect 271 2346 275 2347
rect 271 2341 275 2342
rect 327 2346 331 2347
rect 327 2341 331 2342
rect 399 2346 403 2347
rect 399 2341 403 2342
rect 471 2346 475 2347
rect 471 2341 475 2342
rect 543 2346 547 2347
rect 543 2341 547 2342
rect 551 2346 555 2347
rect 551 2341 555 2342
rect 615 2346 619 2347
rect 615 2341 619 2342
rect 631 2346 635 2347
rect 631 2341 635 2342
rect 687 2346 691 2347
rect 687 2341 691 2342
rect 711 2346 715 2347
rect 711 2341 715 2342
rect 751 2346 755 2347
rect 751 2341 755 2342
rect 783 2346 787 2347
rect 783 2341 787 2342
rect 823 2346 827 2347
rect 823 2341 827 2342
rect 855 2346 859 2347
rect 855 2341 859 2342
rect 895 2346 899 2347
rect 895 2341 899 2342
rect 919 2346 923 2347
rect 919 2341 923 2342
rect 967 2346 971 2347
rect 967 2341 971 2342
rect 991 2346 995 2347
rect 991 2341 995 2342
rect 1063 2346 1067 2347
rect 1063 2341 1067 2342
rect 1239 2346 1243 2347
rect 1279 2345 1283 2346
rect 1327 2350 1331 2351
rect 1327 2345 1331 2346
rect 1375 2350 1379 2351
rect 1375 2345 1379 2346
rect 1383 2350 1387 2351
rect 1383 2345 1387 2346
rect 1415 2350 1419 2351
rect 1415 2345 1419 2346
rect 1439 2350 1443 2351
rect 1439 2345 1443 2346
rect 1455 2350 1459 2351
rect 1455 2345 1459 2346
rect 1503 2350 1507 2351
rect 1503 2345 1507 2346
rect 1559 2350 1563 2351
rect 1559 2345 1563 2346
rect 1575 2350 1579 2351
rect 1575 2345 1579 2346
rect 1615 2350 1619 2351
rect 1615 2345 1619 2346
rect 1647 2350 1651 2351
rect 1647 2345 1651 2346
rect 1679 2350 1683 2351
rect 1679 2345 1683 2346
rect 1719 2350 1723 2351
rect 1719 2345 1723 2346
rect 1735 2350 1739 2351
rect 1735 2345 1739 2346
rect 1799 2350 1803 2351
rect 1799 2345 1803 2346
rect 1871 2350 1875 2351
rect 1871 2345 1875 2346
rect 1879 2350 1883 2351
rect 1879 2345 1883 2346
rect 1951 2350 1955 2351
rect 1951 2345 1955 2346
rect 1967 2350 1971 2351
rect 1967 2345 1971 2346
rect 2047 2350 2051 2351
rect 2047 2345 2051 2346
rect 2063 2350 2067 2351
rect 2063 2345 2067 2346
rect 2151 2350 2155 2351
rect 2151 2345 2155 2346
rect 2167 2350 2171 2351
rect 2167 2345 2171 2346
rect 2263 2350 2267 2351
rect 2263 2345 2267 2346
rect 2271 2350 2275 2351
rect 2271 2345 2275 2346
rect 2359 2350 2363 2351
rect 2359 2345 2363 2346
rect 2407 2350 2411 2351
rect 2407 2345 2411 2346
rect 1239 2341 1243 2342
rect 112 2309 114 2341
rect 272 2332 274 2341
rect 328 2332 330 2341
rect 400 2332 402 2341
rect 472 2332 474 2341
rect 552 2332 554 2341
rect 632 2332 634 2341
rect 712 2332 714 2341
rect 784 2332 786 2341
rect 856 2332 858 2341
rect 920 2332 922 2341
rect 992 2332 994 2341
rect 1064 2332 1066 2341
rect 270 2331 276 2332
rect 270 2327 271 2331
rect 275 2327 276 2331
rect 270 2326 276 2327
rect 326 2331 332 2332
rect 326 2327 327 2331
rect 331 2327 332 2331
rect 326 2326 332 2327
rect 398 2331 404 2332
rect 398 2327 399 2331
rect 403 2327 404 2331
rect 398 2326 404 2327
rect 470 2331 476 2332
rect 470 2327 471 2331
rect 475 2327 476 2331
rect 470 2326 476 2327
rect 550 2331 556 2332
rect 550 2327 551 2331
rect 555 2327 556 2331
rect 550 2326 556 2327
rect 630 2331 636 2332
rect 630 2327 631 2331
rect 635 2327 636 2331
rect 630 2326 636 2327
rect 710 2331 716 2332
rect 710 2327 711 2331
rect 715 2327 716 2331
rect 710 2326 716 2327
rect 782 2331 788 2332
rect 782 2327 783 2331
rect 787 2327 788 2331
rect 782 2326 788 2327
rect 854 2331 860 2332
rect 854 2327 855 2331
rect 859 2327 860 2331
rect 854 2326 860 2327
rect 918 2331 924 2332
rect 918 2327 919 2331
rect 923 2327 924 2331
rect 918 2326 924 2327
rect 990 2331 996 2332
rect 990 2327 991 2331
rect 995 2327 996 2331
rect 990 2326 996 2327
rect 1062 2331 1068 2332
rect 1062 2327 1063 2331
rect 1067 2327 1068 2331
rect 1062 2326 1068 2327
rect 1240 2309 1242 2341
rect 1280 2313 1282 2345
rect 1328 2336 1330 2345
rect 1384 2336 1386 2345
rect 1440 2336 1442 2345
rect 1504 2336 1506 2345
rect 1576 2336 1578 2345
rect 1648 2336 1650 2345
rect 1720 2336 1722 2345
rect 1800 2336 1802 2345
rect 1880 2336 1882 2345
rect 1968 2336 1970 2345
rect 2064 2336 2066 2345
rect 2168 2336 2170 2345
rect 2272 2336 2274 2345
rect 2360 2336 2362 2345
rect 1326 2335 1332 2336
rect 1326 2331 1327 2335
rect 1331 2331 1332 2335
rect 1326 2330 1332 2331
rect 1382 2335 1388 2336
rect 1382 2331 1383 2335
rect 1387 2331 1388 2335
rect 1382 2330 1388 2331
rect 1438 2335 1444 2336
rect 1438 2331 1439 2335
rect 1443 2331 1444 2335
rect 1438 2330 1444 2331
rect 1502 2335 1508 2336
rect 1502 2331 1503 2335
rect 1507 2331 1508 2335
rect 1502 2330 1508 2331
rect 1574 2335 1580 2336
rect 1574 2331 1575 2335
rect 1579 2331 1580 2335
rect 1574 2330 1580 2331
rect 1646 2335 1652 2336
rect 1646 2331 1647 2335
rect 1651 2331 1652 2335
rect 1646 2330 1652 2331
rect 1718 2335 1724 2336
rect 1718 2331 1719 2335
rect 1723 2331 1724 2335
rect 1718 2330 1724 2331
rect 1798 2335 1804 2336
rect 1798 2331 1799 2335
rect 1803 2331 1804 2335
rect 1798 2330 1804 2331
rect 1878 2335 1884 2336
rect 1878 2331 1879 2335
rect 1883 2331 1884 2335
rect 1878 2330 1884 2331
rect 1966 2335 1972 2336
rect 1966 2331 1967 2335
rect 1971 2331 1972 2335
rect 1966 2330 1972 2331
rect 2062 2335 2068 2336
rect 2062 2331 2063 2335
rect 2067 2331 2068 2335
rect 2062 2330 2068 2331
rect 2166 2335 2172 2336
rect 2166 2331 2167 2335
rect 2171 2331 2172 2335
rect 2166 2330 2172 2331
rect 2270 2335 2276 2336
rect 2270 2331 2271 2335
rect 2275 2331 2276 2335
rect 2270 2330 2276 2331
rect 2358 2335 2364 2336
rect 2358 2331 2359 2335
rect 2363 2331 2364 2335
rect 2358 2330 2364 2331
rect 2408 2313 2410 2345
rect 1278 2312 1284 2313
rect 110 2308 116 2309
rect 110 2304 111 2308
rect 115 2304 116 2308
rect 110 2303 116 2304
rect 1238 2308 1244 2309
rect 1238 2304 1239 2308
rect 1243 2304 1244 2308
rect 1278 2308 1279 2312
rect 1283 2308 1284 2312
rect 1278 2307 1284 2308
rect 2406 2312 2412 2313
rect 2406 2308 2407 2312
rect 2411 2308 2412 2312
rect 2406 2307 2412 2308
rect 1238 2303 1244 2304
rect 1278 2295 1284 2296
rect 110 2291 116 2292
rect 110 2287 111 2291
rect 115 2287 116 2291
rect 110 2286 116 2287
rect 1238 2291 1244 2292
rect 1238 2287 1239 2291
rect 1243 2287 1244 2291
rect 1278 2291 1279 2295
rect 1283 2291 1284 2295
rect 1278 2290 1284 2291
rect 2406 2295 2412 2296
rect 2406 2291 2407 2295
rect 2411 2291 2412 2295
rect 2406 2290 2412 2291
rect 1238 2286 1244 2287
rect 112 2271 114 2286
rect 270 2284 276 2285
rect 270 2280 271 2284
rect 275 2280 276 2284
rect 270 2279 276 2280
rect 326 2284 332 2285
rect 326 2280 327 2284
rect 331 2280 332 2284
rect 326 2279 332 2280
rect 398 2284 404 2285
rect 398 2280 399 2284
rect 403 2280 404 2284
rect 398 2279 404 2280
rect 470 2284 476 2285
rect 470 2280 471 2284
rect 475 2280 476 2284
rect 470 2279 476 2280
rect 550 2284 556 2285
rect 550 2280 551 2284
rect 555 2280 556 2284
rect 550 2279 556 2280
rect 630 2284 636 2285
rect 630 2280 631 2284
rect 635 2280 636 2284
rect 630 2279 636 2280
rect 710 2284 716 2285
rect 710 2280 711 2284
rect 715 2280 716 2284
rect 710 2279 716 2280
rect 782 2284 788 2285
rect 782 2280 783 2284
rect 787 2280 788 2284
rect 782 2279 788 2280
rect 854 2284 860 2285
rect 854 2280 855 2284
rect 859 2280 860 2284
rect 854 2279 860 2280
rect 918 2284 924 2285
rect 918 2280 919 2284
rect 923 2280 924 2284
rect 918 2279 924 2280
rect 990 2284 996 2285
rect 990 2280 991 2284
rect 995 2280 996 2284
rect 990 2279 996 2280
rect 1062 2284 1068 2285
rect 1062 2280 1063 2284
rect 1067 2280 1068 2284
rect 1062 2279 1068 2280
rect 272 2271 274 2279
rect 328 2271 330 2279
rect 400 2271 402 2279
rect 472 2271 474 2279
rect 552 2271 554 2279
rect 632 2271 634 2279
rect 712 2271 714 2279
rect 784 2271 786 2279
rect 856 2271 858 2279
rect 920 2271 922 2279
rect 992 2271 994 2279
rect 1064 2271 1066 2279
rect 1240 2271 1242 2286
rect 1280 2283 1282 2290
rect 1326 2288 1332 2289
rect 1326 2284 1327 2288
rect 1331 2284 1332 2288
rect 1326 2283 1332 2284
rect 1382 2288 1388 2289
rect 1382 2284 1383 2288
rect 1387 2284 1388 2288
rect 1382 2283 1388 2284
rect 1438 2288 1444 2289
rect 1438 2284 1439 2288
rect 1443 2284 1444 2288
rect 1438 2283 1444 2284
rect 1502 2288 1508 2289
rect 1502 2284 1503 2288
rect 1507 2284 1508 2288
rect 1502 2283 1508 2284
rect 1574 2288 1580 2289
rect 1574 2284 1575 2288
rect 1579 2284 1580 2288
rect 1574 2283 1580 2284
rect 1646 2288 1652 2289
rect 1646 2284 1647 2288
rect 1651 2284 1652 2288
rect 1646 2283 1652 2284
rect 1718 2288 1724 2289
rect 1718 2284 1719 2288
rect 1723 2284 1724 2288
rect 1718 2283 1724 2284
rect 1798 2288 1804 2289
rect 1798 2284 1799 2288
rect 1803 2284 1804 2288
rect 1798 2283 1804 2284
rect 1878 2288 1884 2289
rect 1878 2284 1879 2288
rect 1883 2284 1884 2288
rect 1878 2283 1884 2284
rect 1966 2288 1972 2289
rect 1966 2284 1967 2288
rect 1971 2284 1972 2288
rect 1966 2283 1972 2284
rect 2062 2288 2068 2289
rect 2062 2284 2063 2288
rect 2067 2284 2068 2288
rect 2062 2283 2068 2284
rect 2166 2288 2172 2289
rect 2166 2284 2167 2288
rect 2171 2284 2172 2288
rect 2166 2283 2172 2284
rect 2270 2288 2276 2289
rect 2270 2284 2271 2288
rect 2275 2284 2276 2288
rect 2270 2283 2276 2284
rect 2358 2288 2364 2289
rect 2358 2284 2359 2288
rect 2363 2284 2364 2288
rect 2358 2283 2364 2284
rect 2408 2283 2410 2290
rect 1279 2282 1283 2283
rect 1279 2277 1283 2278
rect 1327 2282 1331 2283
rect 1327 2277 1331 2278
rect 1335 2282 1339 2283
rect 1335 2277 1339 2278
rect 1383 2282 1387 2283
rect 1383 2277 1387 2278
rect 1407 2282 1411 2283
rect 1407 2277 1411 2278
rect 1439 2282 1443 2283
rect 1439 2277 1443 2278
rect 1487 2282 1491 2283
rect 1487 2277 1491 2278
rect 1503 2282 1507 2283
rect 1503 2277 1507 2278
rect 1559 2282 1563 2283
rect 1559 2277 1563 2278
rect 1575 2282 1579 2283
rect 1575 2277 1579 2278
rect 1631 2282 1635 2283
rect 1631 2277 1635 2278
rect 1647 2282 1651 2283
rect 1647 2277 1651 2278
rect 1703 2282 1707 2283
rect 1703 2277 1707 2278
rect 1719 2282 1723 2283
rect 1719 2277 1723 2278
rect 1775 2282 1779 2283
rect 1775 2277 1779 2278
rect 1799 2282 1803 2283
rect 1799 2277 1803 2278
rect 1839 2282 1843 2283
rect 1839 2277 1843 2278
rect 1879 2282 1883 2283
rect 1879 2277 1883 2278
rect 1911 2282 1915 2283
rect 1911 2277 1915 2278
rect 1967 2282 1971 2283
rect 1967 2277 1971 2278
rect 1991 2282 1995 2283
rect 1991 2277 1995 2278
rect 2063 2282 2067 2283
rect 2063 2277 2067 2278
rect 2079 2282 2083 2283
rect 2079 2277 2083 2278
rect 2167 2282 2171 2283
rect 2167 2277 2171 2278
rect 2175 2282 2179 2283
rect 2175 2277 2179 2278
rect 2271 2282 2275 2283
rect 2271 2277 2275 2278
rect 2279 2282 2283 2283
rect 2279 2277 2283 2278
rect 2359 2282 2363 2283
rect 2359 2277 2363 2278
rect 2407 2282 2411 2283
rect 2407 2277 2411 2278
rect 111 2270 115 2271
rect 111 2265 115 2266
rect 143 2270 147 2271
rect 143 2265 147 2266
rect 183 2270 187 2271
rect 183 2265 187 2266
rect 223 2270 227 2271
rect 223 2265 227 2266
rect 271 2270 275 2271
rect 271 2265 275 2266
rect 279 2270 283 2271
rect 279 2265 283 2266
rect 327 2270 331 2271
rect 327 2265 331 2266
rect 335 2270 339 2271
rect 335 2265 339 2266
rect 399 2270 403 2271
rect 399 2265 403 2266
rect 407 2270 411 2271
rect 407 2265 411 2266
rect 471 2270 475 2271
rect 471 2265 475 2266
rect 479 2270 483 2271
rect 479 2265 483 2266
rect 551 2270 555 2271
rect 551 2265 555 2266
rect 559 2270 563 2271
rect 559 2265 563 2266
rect 631 2270 635 2271
rect 631 2265 635 2266
rect 647 2270 651 2271
rect 647 2265 651 2266
rect 711 2270 715 2271
rect 711 2265 715 2266
rect 727 2270 731 2271
rect 727 2265 731 2266
rect 783 2270 787 2271
rect 783 2265 787 2266
rect 807 2270 811 2271
rect 807 2265 811 2266
rect 855 2270 859 2271
rect 855 2265 859 2266
rect 887 2270 891 2271
rect 887 2265 891 2266
rect 919 2270 923 2271
rect 919 2265 923 2266
rect 967 2270 971 2271
rect 967 2265 971 2266
rect 991 2270 995 2271
rect 991 2265 995 2266
rect 1047 2270 1051 2271
rect 1047 2265 1051 2266
rect 1063 2270 1067 2271
rect 1063 2265 1067 2266
rect 1127 2270 1131 2271
rect 1127 2265 1131 2266
rect 1239 2270 1243 2271
rect 1280 2270 1282 2277
rect 1334 2276 1340 2277
rect 1334 2272 1335 2276
rect 1339 2272 1340 2276
rect 1334 2271 1340 2272
rect 1406 2276 1412 2277
rect 1406 2272 1407 2276
rect 1411 2272 1412 2276
rect 1406 2271 1412 2272
rect 1486 2276 1492 2277
rect 1486 2272 1487 2276
rect 1491 2272 1492 2276
rect 1486 2271 1492 2272
rect 1558 2276 1564 2277
rect 1558 2272 1559 2276
rect 1563 2272 1564 2276
rect 1558 2271 1564 2272
rect 1630 2276 1636 2277
rect 1630 2272 1631 2276
rect 1635 2272 1636 2276
rect 1630 2271 1636 2272
rect 1702 2276 1708 2277
rect 1702 2272 1703 2276
rect 1707 2272 1708 2276
rect 1702 2271 1708 2272
rect 1774 2276 1780 2277
rect 1774 2272 1775 2276
rect 1779 2272 1780 2276
rect 1774 2271 1780 2272
rect 1838 2276 1844 2277
rect 1838 2272 1839 2276
rect 1843 2272 1844 2276
rect 1838 2271 1844 2272
rect 1910 2276 1916 2277
rect 1910 2272 1911 2276
rect 1915 2272 1916 2276
rect 1910 2271 1916 2272
rect 1990 2276 1996 2277
rect 1990 2272 1991 2276
rect 1995 2272 1996 2276
rect 1990 2271 1996 2272
rect 2078 2276 2084 2277
rect 2078 2272 2079 2276
rect 2083 2272 2084 2276
rect 2078 2271 2084 2272
rect 2174 2276 2180 2277
rect 2174 2272 2175 2276
rect 2179 2272 2180 2276
rect 2174 2271 2180 2272
rect 2278 2276 2284 2277
rect 2278 2272 2279 2276
rect 2283 2272 2284 2276
rect 2278 2271 2284 2272
rect 2358 2276 2364 2277
rect 2358 2272 2359 2276
rect 2363 2272 2364 2276
rect 2358 2271 2364 2272
rect 2408 2270 2410 2277
rect 1239 2265 1243 2266
rect 1278 2269 1284 2270
rect 1278 2265 1279 2269
rect 1283 2265 1284 2269
rect 112 2258 114 2265
rect 142 2264 148 2265
rect 142 2260 143 2264
rect 147 2260 148 2264
rect 142 2259 148 2260
rect 182 2264 188 2265
rect 182 2260 183 2264
rect 187 2260 188 2264
rect 182 2259 188 2260
rect 222 2264 228 2265
rect 222 2260 223 2264
rect 227 2260 228 2264
rect 222 2259 228 2260
rect 278 2264 284 2265
rect 278 2260 279 2264
rect 283 2260 284 2264
rect 278 2259 284 2260
rect 334 2264 340 2265
rect 334 2260 335 2264
rect 339 2260 340 2264
rect 334 2259 340 2260
rect 406 2264 412 2265
rect 406 2260 407 2264
rect 411 2260 412 2264
rect 406 2259 412 2260
rect 478 2264 484 2265
rect 478 2260 479 2264
rect 483 2260 484 2264
rect 478 2259 484 2260
rect 558 2264 564 2265
rect 558 2260 559 2264
rect 563 2260 564 2264
rect 558 2259 564 2260
rect 646 2264 652 2265
rect 646 2260 647 2264
rect 651 2260 652 2264
rect 646 2259 652 2260
rect 726 2264 732 2265
rect 726 2260 727 2264
rect 731 2260 732 2264
rect 726 2259 732 2260
rect 806 2264 812 2265
rect 806 2260 807 2264
rect 811 2260 812 2264
rect 806 2259 812 2260
rect 886 2264 892 2265
rect 886 2260 887 2264
rect 891 2260 892 2264
rect 886 2259 892 2260
rect 966 2264 972 2265
rect 966 2260 967 2264
rect 971 2260 972 2264
rect 966 2259 972 2260
rect 1046 2264 1052 2265
rect 1046 2260 1047 2264
rect 1051 2260 1052 2264
rect 1046 2259 1052 2260
rect 1126 2264 1132 2265
rect 1126 2260 1127 2264
rect 1131 2260 1132 2264
rect 1126 2259 1132 2260
rect 1240 2258 1242 2265
rect 1278 2264 1284 2265
rect 2406 2269 2412 2270
rect 2406 2265 2407 2269
rect 2411 2265 2412 2269
rect 2406 2264 2412 2265
rect 110 2257 116 2258
rect 110 2253 111 2257
rect 115 2253 116 2257
rect 110 2252 116 2253
rect 1238 2257 1244 2258
rect 1238 2253 1239 2257
rect 1243 2253 1244 2257
rect 1238 2252 1244 2253
rect 1278 2252 1284 2253
rect 1278 2248 1279 2252
rect 1283 2248 1284 2252
rect 1278 2247 1284 2248
rect 2406 2252 2412 2253
rect 2406 2248 2407 2252
rect 2411 2248 2412 2252
rect 2406 2247 2412 2248
rect 110 2240 116 2241
rect 110 2236 111 2240
rect 115 2236 116 2240
rect 110 2235 116 2236
rect 1238 2240 1244 2241
rect 1238 2236 1239 2240
rect 1243 2236 1244 2240
rect 1238 2235 1244 2236
rect 112 2203 114 2235
rect 142 2217 148 2218
rect 142 2213 143 2217
rect 147 2213 148 2217
rect 142 2212 148 2213
rect 182 2217 188 2218
rect 182 2213 183 2217
rect 187 2213 188 2217
rect 182 2212 188 2213
rect 222 2217 228 2218
rect 222 2213 223 2217
rect 227 2213 228 2217
rect 222 2212 228 2213
rect 278 2217 284 2218
rect 278 2213 279 2217
rect 283 2213 284 2217
rect 278 2212 284 2213
rect 334 2217 340 2218
rect 334 2213 335 2217
rect 339 2213 340 2217
rect 334 2212 340 2213
rect 406 2217 412 2218
rect 406 2213 407 2217
rect 411 2213 412 2217
rect 406 2212 412 2213
rect 478 2217 484 2218
rect 478 2213 479 2217
rect 483 2213 484 2217
rect 478 2212 484 2213
rect 558 2217 564 2218
rect 558 2213 559 2217
rect 563 2213 564 2217
rect 558 2212 564 2213
rect 646 2217 652 2218
rect 646 2213 647 2217
rect 651 2213 652 2217
rect 646 2212 652 2213
rect 726 2217 732 2218
rect 726 2213 727 2217
rect 731 2213 732 2217
rect 726 2212 732 2213
rect 806 2217 812 2218
rect 806 2213 807 2217
rect 811 2213 812 2217
rect 806 2212 812 2213
rect 886 2217 892 2218
rect 886 2213 887 2217
rect 891 2213 892 2217
rect 886 2212 892 2213
rect 966 2217 972 2218
rect 966 2213 967 2217
rect 971 2213 972 2217
rect 966 2212 972 2213
rect 1046 2217 1052 2218
rect 1046 2213 1047 2217
rect 1051 2213 1052 2217
rect 1046 2212 1052 2213
rect 1126 2217 1132 2218
rect 1126 2213 1127 2217
rect 1131 2213 1132 2217
rect 1126 2212 1132 2213
rect 144 2203 146 2212
rect 184 2203 186 2212
rect 224 2203 226 2212
rect 280 2203 282 2212
rect 336 2203 338 2212
rect 408 2203 410 2212
rect 480 2203 482 2212
rect 560 2203 562 2212
rect 648 2203 650 2212
rect 728 2203 730 2212
rect 808 2203 810 2212
rect 888 2203 890 2212
rect 968 2203 970 2212
rect 1048 2203 1050 2212
rect 1128 2203 1130 2212
rect 1240 2203 1242 2235
rect 1280 2207 1282 2247
rect 1334 2229 1340 2230
rect 1334 2225 1335 2229
rect 1339 2225 1340 2229
rect 1334 2224 1340 2225
rect 1406 2229 1412 2230
rect 1406 2225 1407 2229
rect 1411 2225 1412 2229
rect 1406 2224 1412 2225
rect 1486 2229 1492 2230
rect 1486 2225 1487 2229
rect 1491 2225 1492 2229
rect 1486 2224 1492 2225
rect 1558 2229 1564 2230
rect 1558 2225 1559 2229
rect 1563 2225 1564 2229
rect 1558 2224 1564 2225
rect 1630 2229 1636 2230
rect 1630 2225 1631 2229
rect 1635 2225 1636 2229
rect 1630 2224 1636 2225
rect 1702 2229 1708 2230
rect 1702 2225 1703 2229
rect 1707 2225 1708 2229
rect 1702 2224 1708 2225
rect 1774 2229 1780 2230
rect 1774 2225 1775 2229
rect 1779 2225 1780 2229
rect 1774 2224 1780 2225
rect 1838 2229 1844 2230
rect 1838 2225 1839 2229
rect 1843 2225 1844 2229
rect 1838 2224 1844 2225
rect 1910 2229 1916 2230
rect 1910 2225 1911 2229
rect 1915 2225 1916 2229
rect 1910 2224 1916 2225
rect 1990 2229 1996 2230
rect 1990 2225 1991 2229
rect 1995 2225 1996 2229
rect 1990 2224 1996 2225
rect 2078 2229 2084 2230
rect 2078 2225 2079 2229
rect 2083 2225 2084 2229
rect 2078 2224 2084 2225
rect 2174 2229 2180 2230
rect 2174 2225 2175 2229
rect 2179 2225 2180 2229
rect 2174 2224 2180 2225
rect 2278 2229 2284 2230
rect 2278 2225 2279 2229
rect 2283 2225 2284 2229
rect 2278 2224 2284 2225
rect 2358 2229 2364 2230
rect 2358 2225 2359 2229
rect 2363 2225 2364 2229
rect 2358 2224 2364 2225
rect 1336 2207 1338 2224
rect 1408 2207 1410 2224
rect 1488 2207 1490 2224
rect 1560 2207 1562 2224
rect 1632 2207 1634 2224
rect 1704 2207 1706 2224
rect 1776 2207 1778 2224
rect 1840 2207 1842 2224
rect 1912 2207 1914 2224
rect 1992 2207 1994 2224
rect 2080 2207 2082 2224
rect 2176 2207 2178 2224
rect 2280 2207 2282 2224
rect 2360 2207 2362 2224
rect 2408 2207 2410 2247
rect 1279 2206 1283 2207
rect 111 2202 115 2203
rect 111 2197 115 2198
rect 135 2202 139 2203
rect 135 2197 139 2198
rect 143 2202 147 2203
rect 143 2197 147 2198
rect 183 2202 187 2203
rect 183 2197 187 2198
rect 207 2202 211 2203
rect 207 2197 211 2198
rect 223 2202 227 2203
rect 223 2197 227 2198
rect 279 2202 283 2203
rect 279 2197 283 2198
rect 335 2202 339 2203
rect 335 2197 339 2198
rect 359 2202 363 2203
rect 359 2197 363 2198
rect 407 2202 411 2203
rect 407 2197 411 2198
rect 439 2202 443 2203
rect 439 2197 443 2198
rect 479 2202 483 2203
rect 479 2197 483 2198
rect 519 2202 523 2203
rect 519 2197 523 2198
rect 559 2202 563 2203
rect 559 2197 563 2198
rect 599 2202 603 2203
rect 599 2197 603 2198
rect 647 2202 651 2203
rect 647 2197 651 2198
rect 679 2202 683 2203
rect 679 2197 683 2198
rect 727 2202 731 2203
rect 727 2197 731 2198
rect 759 2202 763 2203
rect 759 2197 763 2198
rect 807 2202 811 2203
rect 807 2197 811 2198
rect 831 2202 835 2203
rect 831 2197 835 2198
rect 887 2202 891 2203
rect 887 2197 891 2198
rect 903 2202 907 2203
rect 903 2197 907 2198
rect 967 2202 971 2203
rect 967 2197 971 2198
rect 975 2202 979 2203
rect 975 2197 979 2198
rect 1047 2202 1051 2203
rect 1047 2197 1051 2198
rect 1119 2202 1123 2203
rect 1119 2197 1123 2198
rect 1127 2202 1131 2203
rect 1127 2197 1131 2198
rect 1239 2202 1243 2203
rect 1279 2201 1283 2202
rect 1335 2206 1339 2207
rect 1335 2201 1339 2202
rect 1375 2206 1379 2207
rect 1375 2201 1379 2202
rect 1407 2206 1411 2207
rect 1407 2201 1411 2202
rect 1439 2206 1443 2207
rect 1439 2201 1443 2202
rect 1487 2206 1491 2207
rect 1487 2201 1491 2202
rect 1511 2206 1515 2207
rect 1511 2201 1515 2202
rect 1559 2206 1563 2207
rect 1559 2201 1563 2202
rect 1591 2206 1595 2207
rect 1591 2201 1595 2202
rect 1631 2206 1635 2207
rect 1631 2201 1635 2202
rect 1671 2206 1675 2207
rect 1671 2201 1675 2202
rect 1703 2206 1707 2207
rect 1703 2201 1707 2202
rect 1751 2206 1755 2207
rect 1751 2201 1755 2202
rect 1775 2206 1779 2207
rect 1775 2201 1779 2202
rect 1831 2206 1835 2207
rect 1831 2201 1835 2202
rect 1839 2206 1843 2207
rect 1839 2201 1843 2202
rect 1903 2206 1907 2207
rect 1903 2201 1907 2202
rect 1911 2206 1915 2207
rect 1911 2201 1915 2202
rect 1967 2206 1971 2207
rect 1967 2201 1971 2202
rect 1991 2206 1995 2207
rect 1991 2201 1995 2202
rect 2031 2206 2035 2207
rect 2031 2201 2035 2202
rect 2079 2206 2083 2207
rect 2079 2201 2083 2202
rect 2095 2206 2099 2207
rect 2095 2201 2099 2202
rect 2167 2206 2171 2207
rect 2167 2201 2171 2202
rect 2175 2206 2179 2207
rect 2175 2201 2179 2202
rect 2239 2206 2243 2207
rect 2239 2201 2243 2202
rect 2279 2206 2283 2207
rect 2279 2201 2283 2202
rect 2311 2206 2315 2207
rect 2311 2201 2315 2202
rect 2359 2206 2363 2207
rect 2359 2201 2363 2202
rect 2407 2206 2411 2207
rect 2407 2201 2411 2202
rect 1239 2197 1243 2198
rect 112 2165 114 2197
rect 136 2188 138 2197
rect 208 2188 210 2197
rect 280 2188 282 2197
rect 360 2188 362 2197
rect 440 2188 442 2197
rect 520 2188 522 2197
rect 600 2188 602 2197
rect 680 2188 682 2197
rect 760 2188 762 2197
rect 832 2188 834 2197
rect 904 2188 906 2197
rect 976 2188 978 2197
rect 1048 2188 1050 2197
rect 1120 2188 1122 2197
rect 134 2187 140 2188
rect 134 2183 135 2187
rect 139 2183 140 2187
rect 134 2182 140 2183
rect 206 2187 212 2188
rect 206 2183 207 2187
rect 211 2183 212 2187
rect 206 2182 212 2183
rect 278 2187 284 2188
rect 278 2183 279 2187
rect 283 2183 284 2187
rect 278 2182 284 2183
rect 358 2187 364 2188
rect 358 2183 359 2187
rect 363 2183 364 2187
rect 358 2182 364 2183
rect 438 2187 444 2188
rect 438 2183 439 2187
rect 443 2183 444 2187
rect 438 2182 444 2183
rect 518 2187 524 2188
rect 518 2183 519 2187
rect 523 2183 524 2187
rect 518 2182 524 2183
rect 598 2187 604 2188
rect 598 2183 599 2187
rect 603 2183 604 2187
rect 598 2182 604 2183
rect 678 2187 684 2188
rect 678 2183 679 2187
rect 683 2183 684 2187
rect 678 2182 684 2183
rect 758 2187 764 2188
rect 758 2183 759 2187
rect 763 2183 764 2187
rect 758 2182 764 2183
rect 830 2187 836 2188
rect 830 2183 831 2187
rect 835 2183 836 2187
rect 830 2182 836 2183
rect 902 2187 908 2188
rect 902 2183 903 2187
rect 907 2183 908 2187
rect 902 2182 908 2183
rect 974 2187 980 2188
rect 974 2183 975 2187
rect 979 2183 980 2187
rect 974 2182 980 2183
rect 1046 2187 1052 2188
rect 1046 2183 1047 2187
rect 1051 2183 1052 2187
rect 1046 2182 1052 2183
rect 1118 2187 1124 2188
rect 1118 2183 1119 2187
rect 1123 2183 1124 2187
rect 1118 2182 1124 2183
rect 1240 2165 1242 2197
rect 1280 2169 1282 2201
rect 1376 2192 1378 2201
rect 1440 2192 1442 2201
rect 1512 2192 1514 2201
rect 1592 2192 1594 2201
rect 1672 2192 1674 2201
rect 1752 2192 1754 2201
rect 1832 2192 1834 2201
rect 1904 2192 1906 2201
rect 1968 2192 1970 2201
rect 2032 2192 2034 2201
rect 2096 2192 2098 2201
rect 2168 2192 2170 2201
rect 2240 2192 2242 2201
rect 2312 2192 2314 2201
rect 2360 2192 2362 2201
rect 1374 2191 1380 2192
rect 1374 2187 1375 2191
rect 1379 2187 1380 2191
rect 1374 2186 1380 2187
rect 1438 2191 1444 2192
rect 1438 2187 1439 2191
rect 1443 2187 1444 2191
rect 1438 2186 1444 2187
rect 1510 2191 1516 2192
rect 1510 2187 1511 2191
rect 1515 2187 1516 2191
rect 1510 2186 1516 2187
rect 1590 2191 1596 2192
rect 1590 2187 1591 2191
rect 1595 2187 1596 2191
rect 1590 2186 1596 2187
rect 1670 2191 1676 2192
rect 1670 2187 1671 2191
rect 1675 2187 1676 2191
rect 1670 2186 1676 2187
rect 1750 2191 1756 2192
rect 1750 2187 1751 2191
rect 1755 2187 1756 2191
rect 1750 2186 1756 2187
rect 1830 2191 1836 2192
rect 1830 2187 1831 2191
rect 1835 2187 1836 2191
rect 1830 2186 1836 2187
rect 1902 2191 1908 2192
rect 1902 2187 1903 2191
rect 1907 2187 1908 2191
rect 1902 2186 1908 2187
rect 1966 2191 1972 2192
rect 1966 2187 1967 2191
rect 1971 2187 1972 2191
rect 1966 2186 1972 2187
rect 2030 2191 2036 2192
rect 2030 2187 2031 2191
rect 2035 2187 2036 2191
rect 2030 2186 2036 2187
rect 2094 2191 2100 2192
rect 2094 2187 2095 2191
rect 2099 2187 2100 2191
rect 2094 2186 2100 2187
rect 2166 2191 2172 2192
rect 2166 2187 2167 2191
rect 2171 2187 2172 2191
rect 2166 2186 2172 2187
rect 2238 2191 2244 2192
rect 2238 2187 2239 2191
rect 2243 2187 2244 2191
rect 2238 2186 2244 2187
rect 2310 2191 2316 2192
rect 2310 2187 2311 2191
rect 2315 2187 2316 2191
rect 2310 2186 2316 2187
rect 2358 2191 2364 2192
rect 2358 2187 2359 2191
rect 2363 2187 2364 2191
rect 2358 2186 2364 2187
rect 2408 2169 2410 2201
rect 1278 2168 1284 2169
rect 110 2164 116 2165
rect 110 2160 111 2164
rect 115 2160 116 2164
rect 110 2159 116 2160
rect 1238 2164 1244 2165
rect 1238 2160 1239 2164
rect 1243 2160 1244 2164
rect 1278 2164 1279 2168
rect 1283 2164 1284 2168
rect 1278 2163 1284 2164
rect 2406 2168 2412 2169
rect 2406 2164 2407 2168
rect 2411 2164 2412 2168
rect 2406 2163 2412 2164
rect 1238 2159 1244 2160
rect 1278 2151 1284 2152
rect 110 2147 116 2148
rect 110 2143 111 2147
rect 115 2143 116 2147
rect 110 2142 116 2143
rect 1238 2147 1244 2148
rect 1238 2143 1239 2147
rect 1243 2143 1244 2147
rect 1278 2147 1279 2151
rect 1283 2147 1284 2151
rect 1278 2146 1284 2147
rect 2406 2151 2412 2152
rect 2406 2147 2407 2151
rect 2411 2147 2412 2151
rect 2406 2146 2412 2147
rect 1238 2142 1244 2143
rect 112 2127 114 2142
rect 134 2140 140 2141
rect 134 2136 135 2140
rect 139 2136 140 2140
rect 134 2135 140 2136
rect 206 2140 212 2141
rect 206 2136 207 2140
rect 211 2136 212 2140
rect 206 2135 212 2136
rect 278 2140 284 2141
rect 278 2136 279 2140
rect 283 2136 284 2140
rect 278 2135 284 2136
rect 358 2140 364 2141
rect 358 2136 359 2140
rect 363 2136 364 2140
rect 358 2135 364 2136
rect 438 2140 444 2141
rect 438 2136 439 2140
rect 443 2136 444 2140
rect 438 2135 444 2136
rect 518 2140 524 2141
rect 518 2136 519 2140
rect 523 2136 524 2140
rect 518 2135 524 2136
rect 598 2140 604 2141
rect 598 2136 599 2140
rect 603 2136 604 2140
rect 598 2135 604 2136
rect 678 2140 684 2141
rect 678 2136 679 2140
rect 683 2136 684 2140
rect 678 2135 684 2136
rect 758 2140 764 2141
rect 758 2136 759 2140
rect 763 2136 764 2140
rect 758 2135 764 2136
rect 830 2140 836 2141
rect 830 2136 831 2140
rect 835 2136 836 2140
rect 830 2135 836 2136
rect 902 2140 908 2141
rect 902 2136 903 2140
rect 907 2136 908 2140
rect 902 2135 908 2136
rect 974 2140 980 2141
rect 974 2136 975 2140
rect 979 2136 980 2140
rect 974 2135 980 2136
rect 1046 2140 1052 2141
rect 1046 2136 1047 2140
rect 1051 2136 1052 2140
rect 1046 2135 1052 2136
rect 1118 2140 1124 2141
rect 1118 2136 1119 2140
rect 1123 2136 1124 2140
rect 1118 2135 1124 2136
rect 136 2127 138 2135
rect 208 2127 210 2135
rect 280 2127 282 2135
rect 360 2127 362 2135
rect 440 2127 442 2135
rect 520 2127 522 2135
rect 600 2127 602 2135
rect 680 2127 682 2135
rect 760 2127 762 2135
rect 832 2127 834 2135
rect 904 2127 906 2135
rect 976 2127 978 2135
rect 1048 2127 1050 2135
rect 1120 2127 1122 2135
rect 1240 2127 1242 2142
rect 1280 2139 1282 2146
rect 1374 2144 1380 2145
rect 1374 2140 1375 2144
rect 1379 2140 1380 2144
rect 1374 2139 1380 2140
rect 1438 2144 1444 2145
rect 1438 2140 1439 2144
rect 1443 2140 1444 2144
rect 1438 2139 1444 2140
rect 1510 2144 1516 2145
rect 1510 2140 1511 2144
rect 1515 2140 1516 2144
rect 1510 2139 1516 2140
rect 1590 2144 1596 2145
rect 1590 2140 1591 2144
rect 1595 2140 1596 2144
rect 1590 2139 1596 2140
rect 1670 2144 1676 2145
rect 1670 2140 1671 2144
rect 1675 2140 1676 2144
rect 1670 2139 1676 2140
rect 1750 2144 1756 2145
rect 1750 2140 1751 2144
rect 1755 2140 1756 2144
rect 1750 2139 1756 2140
rect 1830 2144 1836 2145
rect 1830 2140 1831 2144
rect 1835 2140 1836 2144
rect 1830 2139 1836 2140
rect 1902 2144 1908 2145
rect 1902 2140 1903 2144
rect 1907 2140 1908 2144
rect 1902 2139 1908 2140
rect 1966 2144 1972 2145
rect 1966 2140 1967 2144
rect 1971 2140 1972 2144
rect 1966 2139 1972 2140
rect 2030 2144 2036 2145
rect 2030 2140 2031 2144
rect 2035 2140 2036 2144
rect 2030 2139 2036 2140
rect 2094 2144 2100 2145
rect 2094 2140 2095 2144
rect 2099 2140 2100 2144
rect 2094 2139 2100 2140
rect 2166 2144 2172 2145
rect 2166 2140 2167 2144
rect 2171 2140 2172 2144
rect 2166 2139 2172 2140
rect 2238 2144 2244 2145
rect 2238 2140 2239 2144
rect 2243 2140 2244 2144
rect 2238 2139 2244 2140
rect 2310 2144 2316 2145
rect 2310 2140 2311 2144
rect 2315 2140 2316 2144
rect 2310 2139 2316 2140
rect 2358 2144 2364 2145
rect 2358 2140 2359 2144
rect 2363 2140 2364 2144
rect 2358 2139 2364 2140
rect 2408 2139 2410 2146
rect 1279 2138 1283 2139
rect 1279 2133 1283 2134
rect 1375 2138 1379 2139
rect 1375 2133 1379 2134
rect 1399 2138 1403 2139
rect 1399 2133 1403 2134
rect 1439 2138 1443 2139
rect 1439 2133 1443 2134
rect 1495 2138 1499 2139
rect 1495 2133 1499 2134
rect 1511 2138 1515 2139
rect 1511 2133 1515 2134
rect 1567 2138 1571 2139
rect 1567 2133 1571 2134
rect 1591 2138 1595 2139
rect 1591 2133 1595 2134
rect 1647 2138 1651 2139
rect 1647 2133 1651 2134
rect 1671 2138 1675 2139
rect 1671 2133 1675 2134
rect 1735 2138 1739 2139
rect 1735 2133 1739 2134
rect 1751 2138 1755 2139
rect 1751 2133 1755 2134
rect 1823 2138 1827 2139
rect 1823 2133 1827 2134
rect 1831 2138 1835 2139
rect 1831 2133 1835 2134
rect 1903 2138 1907 2139
rect 1903 2133 1907 2134
rect 1911 2138 1915 2139
rect 1911 2133 1915 2134
rect 1967 2138 1971 2139
rect 1967 2133 1971 2134
rect 1999 2138 2003 2139
rect 1999 2133 2003 2134
rect 2031 2138 2035 2139
rect 2031 2133 2035 2134
rect 2087 2138 2091 2139
rect 2087 2133 2091 2134
rect 2095 2138 2099 2139
rect 2095 2133 2099 2134
rect 2167 2138 2171 2139
rect 2167 2133 2171 2134
rect 2175 2138 2179 2139
rect 2175 2133 2179 2134
rect 2239 2138 2243 2139
rect 2239 2133 2243 2134
rect 2271 2138 2275 2139
rect 2271 2133 2275 2134
rect 2311 2138 2315 2139
rect 2311 2133 2315 2134
rect 2359 2138 2363 2139
rect 2359 2133 2363 2134
rect 2407 2138 2411 2139
rect 2407 2133 2411 2134
rect 111 2126 115 2127
rect 111 2121 115 2122
rect 135 2126 139 2127
rect 135 2121 139 2122
rect 191 2126 195 2127
rect 191 2121 195 2122
rect 207 2126 211 2127
rect 207 2121 211 2122
rect 271 2126 275 2127
rect 271 2121 275 2122
rect 279 2126 283 2127
rect 279 2121 283 2122
rect 343 2126 347 2127
rect 343 2121 347 2122
rect 359 2126 363 2127
rect 359 2121 363 2122
rect 415 2126 419 2127
rect 415 2121 419 2122
rect 439 2126 443 2127
rect 439 2121 443 2122
rect 479 2126 483 2127
rect 479 2121 483 2122
rect 519 2126 523 2127
rect 519 2121 523 2122
rect 543 2126 547 2127
rect 543 2121 547 2122
rect 599 2126 603 2127
rect 599 2121 603 2122
rect 607 2126 611 2127
rect 607 2121 611 2122
rect 671 2126 675 2127
rect 671 2121 675 2122
rect 679 2126 683 2127
rect 679 2121 683 2122
rect 735 2126 739 2127
rect 735 2121 739 2122
rect 759 2126 763 2127
rect 759 2121 763 2122
rect 791 2126 795 2127
rect 791 2121 795 2122
rect 831 2126 835 2127
rect 831 2121 835 2122
rect 839 2126 843 2127
rect 839 2121 843 2122
rect 887 2126 891 2127
rect 887 2121 891 2122
rect 903 2126 907 2127
rect 903 2121 907 2122
rect 935 2126 939 2127
rect 935 2121 939 2122
rect 975 2126 979 2127
rect 975 2121 979 2122
rect 991 2126 995 2127
rect 991 2121 995 2122
rect 1047 2126 1051 2127
rect 1047 2121 1051 2122
rect 1119 2126 1123 2127
rect 1119 2121 1123 2122
rect 1239 2126 1243 2127
rect 1280 2126 1282 2133
rect 1398 2132 1404 2133
rect 1398 2128 1399 2132
rect 1403 2128 1404 2132
rect 1398 2127 1404 2128
rect 1438 2132 1444 2133
rect 1438 2128 1439 2132
rect 1443 2128 1444 2132
rect 1438 2127 1444 2128
rect 1494 2132 1500 2133
rect 1494 2128 1495 2132
rect 1499 2128 1500 2132
rect 1494 2127 1500 2128
rect 1566 2132 1572 2133
rect 1566 2128 1567 2132
rect 1571 2128 1572 2132
rect 1566 2127 1572 2128
rect 1646 2132 1652 2133
rect 1646 2128 1647 2132
rect 1651 2128 1652 2132
rect 1646 2127 1652 2128
rect 1734 2132 1740 2133
rect 1734 2128 1735 2132
rect 1739 2128 1740 2132
rect 1734 2127 1740 2128
rect 1822 2132 1828 2133
rect 1822 2128 1823 2132
rect 1827 2128 1828 2132
rect 1822 2127 1828 2128
rect 1910 2132 1916 2133
rect 1910 2128 1911 2132
rect 1915 2128 1916 2132
rect 1910 2127 1916 2128
rect 1998 2132 2004 2133
rect 1998 2128 1999 2132
rect 2003 2128 2004 2132
rect 1998 2127 2004 2128
rect 2086 2132 2092 2133
rect 2086 2128 2087 2132
rect 2091 2128 2092 2132
rect 2086 2127 2092 2128
rect 2174 2132 2180 2133
rect 2174 2128 2175 2132
rect 2179 2128 2180 2132
rect 2174 2127 2180 2128
rect 2270 2132 2276 2133
rect 2270 2128 2271 2132
rect 2275 2128 2276 2132
rect 2270 2127 2276 2128
rect 2358 2132 2364 2133
rect 2358 2128 2359 2132
rect 2363 2128 2364 2132
rect 2358 2127 2364 2128
rect 2408 2126 2410 2133
rect 1239 2121 1243 2122
rect 1278 2125 1284 2126
rect 1278 2121 1279 2125
rect 1283 2121 1284 2125
rect 112 2114 114 2121
rect 134 2120 140 2121
rect 134 2116 135 2120
rect 139 2116 140 2120
rect 134 2115 140 2116
rect 190 2120 196 2121
rect 190 2116 191 2120
rect 195 2116 196 2120
rect 190 2115 196 2116
rect 270 2120 276 2121
rect 270 2116 271 2120
rect 275 2116 276 2120
rect 270 2115 276 2116
rect 342 2120 348 2121
rect 342 2116 343 2120
rect 347 2116 348 2120
rect 342 2115 348 2116
rect 414 2120 420 2121
rect 414 2116 415 2120
rect 419 2116 420 2120
rect 414 2115 420 2116
rect 478 2120 484 2121
rect 478 2116 479 2120
rect 483 2116 484 2120
rect 478 2115 484 2116
rect 542 2120 548 2121
rect 542 2116 543 2120
rect 547 2116 548 2120
rect 542 2115 548 2116
rect 606 2120 612 2121
rect 606 2116 607 2120
rect 611 2116 612 2120
rect 606 2115 612 2116
rect 670 2120 676 2121
rect 670 2116 671 2120
rect 675 2116 676 2120
rect 670 2115 676 2116
rect 734 2120 740 2121
rect 734 2116 735 2120
rect 739 2116 740 2120
rect 734 2115 740 2116
rect 790 2120 796 2121
rect 790 2116 791 2120
rect 795 2116 796 2120
rect 790 2115 796 2116
rect 838 2120 844 2121
rect 838 2116 839 2120
rect 843 2116 844 2120
rect 838 2115 844 2116
rect 886 2120 892 2121
rect 886 2116 887 2120
rect 891 2116 892 2120
rect 886 2115 892 2116
rect 934 2120 940 2121
rect 934 2116 935 2120
rect 939 2116 940 2120
rect 934 2115 940 2116
rect 990 2120 996 2121
rect 990 2116 991 2120
rect 995 2116 996 2120
rect 990 2115 996 2116
rect 1046 2120 1052 2121
rect 1046 2116 1047 2120
rect 1051 2116 1052 2120
rect 1046 2115 1052 2116
rect 1240 2114 1242 2121
rect 1278 2120 1284 2121
rect 2406 2125 2412 2126
rect 2406 2121 2407 2125
rect 2411 2121 2412 2125
rect 2406 2120 2412 2121
rect 110 2113 116 2114
rect 110 2109 111 2113
rect 115 2109 116 2113
rect 110 2108 116 2109
rect 1238 2113 1244 2114
rect 1238 2109 1239 2113
rect 1243 2109 1244 2113
rect 1238 2108 1244 2109
rect 1278 2108 1284 2109
rect 1278 2104 1279 2108
rect 1283 2104 1284 2108
rect 1278 2103 1284 2104
rect 2406 2108 2412 2109
rect 2406 2104 2407 2108
rect 2411 2104 2412 2108
rect 2406 2103 2412 2104
rect 110 2096 116 2097
rect 110 2092 111 2096
rect 115 2092 116 2096
rect 110 2091 116 2092
rect 1238 2096 1244 2097
rect 1238 2092 1239 2096
rect 1243 2092 1244 2096
rect 1238 2091 1244 2092
rect 112 2055 114 2091
rect 134 2073 140 2074
rect 134 2069 135 2073
rect 139 2069 140 2073
rect 134 2068 140 2069
rect 190 2073 196 2074
rect 190 2069 191 2073
rect 195 2069 196 2073
rect 190 2068 196 2069
rect 270 2073 276 2074
rect 270 2069 271 2073
rect 275 2069 276 2073
rect 270 2068 276 2069
rect 342 2073 348 2074
rect 342 2069 343 2073
rect 347 2069 348 2073
rect 342 2068 348 2069
rect 414 2073 420 2074
rect 414 2069 415 2073
rect 419 2069 420 2073
rect 414 2068 420 2069
rect 478 2073 484 2074
rect 478 2069 479 2073
rect 483 2069 484 2073
rect 478 2068 484 2069
rect 542 2073 548 2074
rect 542 2069 543 2073
rect 547 2069 548 2073
rect 542 2068 548 2069
rect 606 2073 612 2074
rect 606 2069 607 2073
rect 611 2069 612 2073
rect 606 2068 612 2069
rect 670 2073 676 2074
rect 670 2069 671 2073
rect 675 2069 676 2073
rect 670 2068 676 2069
rect 734 2073 740 2074
rect 734 2069 735 2073
rect 739 2069 740 2073
rect 734 2068 740 2069
rect 790 2073 796 2074
rect 790 2069 791 2073
rect 795 2069 796 2073
rect 790 2068 796 2069
rect 838 2073 844 2074
rect 838 2069 839 2073
rect 843 2069 844 2073
rect 838 2068 844 2069
rect 886 2073 892 2074
rect 886 2069 887 2073
rect 891 2069 892 2073
rect 886 2068 892 2069
rect 934 2073 940 2074
rect 934 2069 935 2073
rect 939 2069 940 2073
rect 934 2068 940 2069
rect 990 2073 996 2074
rect 990 2069 991 2073
rect 995 2069 996 2073
rect 990 2068 996 2069
rect 1046 2073 1052 2074
rect 1046 2069 1047 2073
rect 1051 2069 1052 2073
rect 1046 2068 1052 2069
rect 136 2055 138 2068
rect 192 2055 194 2068
rect 272 2055 274 2068
rect 344 2055 346 2068
rect 416 2055 418 2068
rect 480 2055 482 2068
rect 544 2055 546 2068
rect 608 2055 610 2068
rect 672 2055 674 2068
rect 736 2055 738 2068
rect 792 2055 794 2068
rect 840 2055 842 2068
rect 888 2055 890 2068
rect 936 2055 938 2068
rect 992 2055 994 2068
rect 1048 2055 1050 2068
rect 1240 2055 1242 2091
rect 1280 2071 1282 2103
rect 1398 2085 1404 2086
rect 1398 2081 1399 2085
rect 1403 2081 1404 2085
rect 1398 2080 1404 2081
rect 1438 2085 1444 2086
rect 1438 2081 1439 2085
rect 1443 2081 1444 2085
rect 1438 2080 1444 2081
rect 1494 2085 1500 2086
rect 1494 2081 1495 2085
rect 1499 2081 1500 2085
rect 1494 2080 1500 2081
rect 1566 2085 1572 2086
rect 1566 2081 1567 2085
rect 1571 2081 1572 2085
rect 1566 2080 1572 2081
rect 1646 2085 1652 2086
rect 1646 2081 1647 2085
rect 1651 2081 1652 2085
rect 1646 2080 1652 2081
rect 1734 2085 1740 2086
rect 1734 2081 1735 2085
rect 1739 2081 1740 2085
rect 1734 2080 1740 2081
rect 1822 2085 1828 2086
rect 1822 2081 1823 2085
rect 1827 2081 1828 2085
rect 1822 2080 1828 2081
rect 1910 2085 1916 2086
rect 1910 2081 1911 2085
rect 1915 2081 1916 2085
rect 1910 2080 1916 2081
rect 1998 2085 2004 2086
rect 1998 2081 1999 2085
rect 2003 2081 2004 2085
rect 1998 2080 2004 2081
rect 2086 2085 2092 2086
rect 2086 2081 2087 2085
rect 2091 2081 2092 2085
rect 2086 2080 2092 2081
rect 2174 2085 2180 2086
rect 2174 2081 2175 2085
rect 2179 2081 2180 2085
rect 2174 2080 2180 2081
rect 2270 2085 2276 2086
rect 2270 2081 2271 2085
rect 2275 2081 2276 2085
rect 2270 2080 2276 2081
rect 2358 2085 2364 2086
rect 2358 2081 2359 2085
rect 2363 2081 2364 2085
rect 2358 2080 2364 2081
rect 1400 2071 1402 2080
rect 1440 2071 1442 2080
rect 1496 2071 1498 2080
rect 1568 2071 1570 2080
rect 1648 2071 1650 2080
rect 1736 2071 1738 2080
rect 1824 2071 1826 2080
rect 1912 2071 1914 2080
rect 2000 2071 2002 2080
rect 2088 2071 2090 2080
rect 2176 2071 2178 2080
rect 2272 2071 2274 2080
rect 2360 2071 2362 2080
rect 2408 2071 2410 2103
rect 1279 2070 1283 2071
rect 1279 2065 1283 2066
rect 1399 2070 1403 2071
rect 1399 2065 1403 2066
rect 1439 2070 1443 2071
rect 1439 2065 1443 2066
rect 1495 2070 1499 2071
rect 1495 2065 1499 2066
rect 1567 2070 1571 2071
rect 1567 2065 1571 2066
rect 1647 2070 1651 2071
rect 1647 2065 1651 2066
rect 1735 2070 1739 2071
rect 1735 2065 1739 2066
rect 1823 2070 1827 2071
rect 1823 2065 1827 2066
rect 1911 2070 1915 2071
rect 1911 2065 1915 2066
rect 1999 2070 2003 2071
rect 1999 2065 2003 2066
rect 2039 2070 2043 2071
rect 2039 2065 2043 2066
rect 2079 2070 2083 2071
rect 2079 2065 2083 2066
rect 2087 2070 2091 2071
rect 2087 2065 2091 2066
rect 2119 2070 2123 2071
rect 2119 2065 2123 2066
rect 2159 2070 2163 2071
rect 2159 2065 2163 2066
rect 2175 2070 2179 2071
rect 2175 2065 2179 2066
rect 2199 2070 2203 2071
rect 2199 2065 2203 2066
rect 2239 2070 2243 2071
rect 2239 2065 2243 2066
rect 2271 2070 2275 2071
rect 2271 2065 2275 2066
rect 2279 2070 2283 2071
rect 2279 2065 2283 2066
rect 2319 2070 2323 2071
rect 2319 2065 2323 2066
rect 2359 2070 2363 2071
rect 2359 2065 2363 2066
rect 2407 2070 2411 2071
rect 2407 2065 2411 2066
rect 111 2054 115 2055
rect 111 2049 115 2050
rect 135 2054 139 2055
rect 135 2049 139 2050
rect 175 2054 179 2055
rect 175 2049 179 2050
rect 191 2054 195 2055
rect 191 2049 195 2050
rect 215 2054 219 2055
rect 215 2049 219 2050
rect 271 2054 275 2055
rect 271 2049 275 2050
rect 279 2054 283 2055
rect 279 2049 283 2050
rect 343 2054 347 2055
rect 343 2049 347 2050
rect 351 2054 355 2055
rect 351 2049 355 2050
rect 415 2054 419 2055
rect 415 2049 419 2050
rect 423 2054 427 2055
rect 423 2049 427 2050
rect 479 2054 483 2055
rect 479 2049 483 2050
rect 487 2054 491 2055
rect 487 2049 491 2050
rect 543 2054 547 2055
rect 543 2049 547 2050
rect 551 2054 555 2055
rect 551 2049 555 2050
rect 607 2054 611 2055
rect 607 2049 611 2050
rect 615 2054 619 2055
rect 615 2049 619 2050
rect 671 2054 675 2055
rect 671 2049 675 2050
rect 679 2054 683 2055
rect 679 2049 683 2050
rect 735 2054 739 2055
rect 735 2049 739 2050
rect 743 2054 747 2055
rect 743 2049 747 2050
rect 791 2054 795 2055
rect 791 2049 795 2050
rect 815 2054 819 2055
rect 815 2049 819 2050
rect 839 2054 843 2055
rect 839 2049 843 2050
rect 887 2054 891 2055
rect 887 2049 891 2050
rect 935 2054 939 2055
rect 935 2049 939 2050
rect 991 2054 995 2055
rect 991 2049 995 2050
rect 1047 2054 1051 2055
rect 1047 2049 1051 2050
rect 1239 2054 1243 2055
rect 1239 2049 1243 2050
rect 112 2017 114 2049
rect 136 2040 138 2049
rect 176 2040 178 2049
rect 216 2040 218 2049
rect 280 2040 282 2049
rect 352 2040 354 2049
rect 424 2040 426 2049
rect 488 2040 490 2049
rect 552 2040 554 2049
rect 616 2040 618 2049
rect 680 2040 682 2049
rect 744 2040 746 2049
rect 816 2040 818 2049
rect 134 2039 140 2040
rect 134 2035 135 2039
rect 139 2035 140 2039
rect 134 2034 140 2035
rect 174 2039 180 2040
rect 174 2035 175 2039
rect 179 2035 180 2039
rect 174 2034 180 2035
rect 214 2039 220 2040
rect 214 2035 215 2039
rect 219 2035 220 2039
rect 214 2034 220 2035
rect 278 2039 284 2040
rect 278 2035 279 2039
rect 283 2035 284 2039
rect 278 2034 284 2035
rect 350 2039 356 2040
rect 350 2035 351 2039
rect 355 2035 356 2039
rect 350 2034 356 2035
rect 422 2039 428 2040
rect 422 2035 423 2039
rect 427 2035 428 2039
rect 422 2034 428 2035
rect 486 2039 492 2040
rect 486 2035 487 2039
rect 491 2035 492 2039
rect 486 2034 492 2035
rect 550 2039 556 2040
rect 550 2035 551 2039
rect 555 2035 556 2039
rect 550 2034 556 2035
rect 614 2039 620 2040
rect 614 2035 615 2039
rect 619 2035 620 2039
rect 614 2034 620 2035
rect 678 2039 684 2040
rect 678 2035 679 2039
rect 683 2035 684 2039
rect 678 2034 684 2035
rect 742 2039 748 2040
rect 742 2035 743 2039
rect 747 2035 748 2039
rect 742 2034 748 2035
rect 814 2039 820 2040
rect 814 2035 815 2039
rect 819 2035 820 2039
rect 814 2034 820 2035
rect 1240 2017 1242 2049
rect 1280 2033 1282 2065
rect 2040 2056 2042 2065
rect 2080 2056 2082 2065
rect 2120 2056 2122 2065
rect 2160 2056 2162 2065
rect 2200 2056 2202 2065
rect 2240 2056 2242 2065
rect 2280 2056 2282 2065
rect 2320 2056 2322 2065
rect 2360 2056 2362 2065
rect 2038 2055 2044 2056
rect 2038 2051 2039 2055
rect 2043 2051 2044 2055
rect 2038 2050 2044 2051
rect 2078 2055 2084 2056
rect 2078 2051 2079 2055
rect 2083 2051 2084 2055
rect 2078 2050 2084 2051
rect 2118 2055 2124 2056
rect 2118 2051 2119 2055
rect 2123 2051 2124 2055
rect 2118 2050 2124 2051
rect 2158 2055 2164 2056
rect 2158 2051 2159 2055
rect 2163 2051 2164 2055
rect 2158 2050 2164 2051
rect 2198 2055 2204 2056
rect 2198 2051 2199 2055
rect 2203 2051 2204 2055
rect 2198 2050 2204 2051
rect 2238 2055 2244 2056
rect 2238 2051 2239 2055
rect 2243 2051 2244 2055
rect 2238 2050 2244 2051
rect 2278 2055 2284 2056
rect 2278 2051 2279 2055
rect 2283 2051 2284 2055
rect 2278 2050 2284 2051
rect 2318 2055 2324 2056
rect 2318 2051 2319 2055
rect 2323 2051 2324 2055
rect 2318 2050 2324 2051
rect 2358 2055 2364 2056
rect 2358 2051 2359 2055
rect 2363 2051 2364 2055
rect 2358 2050 2364 2051
rect 2408 2033 2410 2065
rect 1278 2032 1284 2033
rect 1278 2028 1279 2032
rect 1283 2028 1284 2032
rect 1278 2027 1284 2028
rect 2406 2032 2412 2033
rect 2406 2028 2407 2032
rect 2411 2028 2412 2032
rect 2406 2027 2412 2028
rect 110 2016 116 2017
rect 110 2012 111 2016
rect 115 2012 116 2016
rect 110 2011 116 2012
rect 1238 2016 1244 2017
rect 1238 2012 1239 2016
rect 1243 2012 1244 2016
rect 1238 2011 1244 2012
rect 1278 2015 1284 2016
rect 1278 2011 1279 2015
rect 1283 2011 1284 2015
rect 1278 2010 1284 2011
rect 2406 2015 2412 2016
rect 2406 2011 2407 2015
rect 2411 2011 2412 2015
rect 2406 2010 2412 2011
rect 1280 2003 1282 2010
rect 2038 2008 2044 2009
rect 2038 2004 2039 2008
rect 2043 2004 2044 2008
rect 2038 2003 2044 2004
rect 2078 2008 2084 2009
rect 2078 2004 2079 2008
rect 2083 2004 2084 2008
rect 2078 2003 2084 2004
rect 2118 2008 2124 2009
rect 2118 2004 2119 2008
rect 2123 2004 2124 2008
rect 2118 2003 2124 2004
rect 2158 2008 2164 2009
rect 2158 2004 2159 2008
rect 2163 2004 2164 2008
rect 2158 2003 2164 2004
rect 2198 2008 2204 2009
rect 2198 2004 2199 2008
rect 2203 2004 2204 2008
rect 2198 2003 2204 2004
rect 2238 2008 2244 2009
rect 2238 2004 2239 2008
rect 2243 2004 2244 2008
rect 2238 2003 2244 2004
rect 2278 2008 2284 2009
rect 2278 2004 2279 2008
rect 2283 2004 2284 2008
rect 2278 2003 2284 2004
rect 2318 2008 2324 2009
rect 2318 2004 2319 2008
rect 2323 2004 2324 2008
rect 2318 2003 2324 2004
rect 2358 2008 2364 2009
rect 2358 2004 2359 2008
rect 2363 2004 2364 2008
rect 2358 2003 2364 2004
rect 2408 2003 2410 2010
rect 1279 2002 1283 2003
rect 110 1999 116 2000
rect 110 1995 111 1999
rect 115 1995 116 1999
rect 110 1994 116 1995
rect 1238 1999 1244 2000
rect 1238 1995 1239 1999
rect 1243 1995 1244 1999
rect 1279 1997 1283 1998
rect 1399 2002 1403 2003
rect 1399 1997 1403 1998
rect 1439 2002 1443 2003
rect 1439 1997 1443 1998
rect 1479 2002 1483 2003
rect 1479 1997 1483 1998
rect 1519 2002 1523 2003
rect 1519 1997 1523 1998
rect 1559 2002 1563 2003
rect 1559 1997 1563 1998
rect 1599 2002 1603 2003
rect 1599 1997 1603 1998
rect 1639 2002 1643 2003
rect 1639 1997 1643 1998
rect 1679 2002 1683 2003
rect 1679 1997 1683 1998
rect 1719 2002 1723 2003
rect 1719 1997 1723 1998
rect 1767 2002 1771 2003
rect 1767 1997 1771 1998
rect 1823 2002 1827 2003
rect 1823 1997 1827 1998
rect 1871 2002 1875 2003
rect 1871 1997 1875 1998
rect 1919 2002 1923 2003
rect 1919 1997 1923 1998
rect 1967 2002 1971 2003
rect 1967 1997 1971 1998
rect 2015 2002 2019 2003
rect 2015 1997 2019 1998
rect 2039 2002 2043 2003
rect 2039 1997 2043 1998
rect 2055 2002 2059 2003
rect 2055 1997 2059 1998
rect 2079 2002 2083 2003
rect 2079 1997 2083 1998
rect 2095 2002 2099 2003
rect 2095 1997 2099 1998
rect 2119 2002 2123 2003
rect 2119 1997 2123 1998
rect 2143 2002 2147 2003
rect 2143 1997 2147 1998
rect 2159 2002 2163 2003
rect 2159 1997 2163 1998
rect 2191 2002 2195 2003
rect 2191 1997 2195 1998
rect 2199 2002 2203 2003
rect 2199 1997 2203 1998
rect 2239 2002 2243 2003
rect 2239 1997 2243 1998
rect 2279 2002 2283 2003
rect 2279 1997 2283 1998
rect 2319 2002 2323 2003
rect 2319 1997 2323 1998
rect 2359 2002 2363 2003
rect 2359 1997 2363 1998
rect 2407 2002 2411 2003
rect 2407 1997 2411 1998
rect 1238 1994 1244 1995
rect 112 1987 114 1994
rect 134 1992 140 1993
rect 134 1988 135 1992
rect 139 1988 140 1992
rect 134 1987 140 1988
rect 174 1992 180 1993
rect 174 1988 175 1992
rect 179 1988 180 1992
rect 174 1987 180 1988
rect 214 1992 220 1993
rect 214 1988 215 1992
rect 219 1988 220 1992
rect 214 1987 220 1988
rect 278 1992 284 1993
rect 278 1988 279 1992
rect 283 1988 284 1992
rect 278 1987 284 1988
rect 350 1992 356 1993
rect 350 1988 351 1992
rect 355 1988 356 1992
rect 350 1987 356 1988
rect 422 1992 428 1993
rect 422 1988 423 1992
rect 427 1988 428 1992
rect 422 1987 428 1988
rect 486 1992 492 1993
rect 486 1988 487 1992
rect 491 1988 492 1992
rect 486 1987 492 1988
rect 550 1992 556 1993
rect 550 1988 551 1992
rect 555 1988 556 1992
rect 550 1987 556 1988
rect 614 1992 620 1993
rect 614 1988 615 1992
rect 619 1988 620 1992
rect 614 1987 620 1988
rect 678 1992 684 1993
rect 678 1988 679 1992
rect 683 1988 684 1992
rect 678 1987 684 1988
rect 742 1992 748 1993
rect 742 1988 743 1992
rect 747 1988 748 1992
rect 742 1987 748 1988
rect 814 1992 820 1993
rect 814 1988 815 1992
rect 819 1988 820 1992
rect 814 1987 820 1988
rect 1240 1987 1242 1994
rect 1280 1990 1282 1997
rect 1398 1996 1404 1997
rect 1398 1992 1399 1996
rect 1403 1992 1404 1996
rect 1398 1991 1404 1992
rect 1438 1996 1444 1997
rect 1438 1992 1439 1996
rect 1443 1992 1444 1996
rect 1438 1991 1444 1992
rect 1478 1996 1484 1997
rect 1478 1992 1479 1996
rect 1483 1992 1484 1996
rect 1478 1991 1484 1992
rect 1518 1996 1524 1997
rect 1518 1992 1519 1996
rect 1523 1992 1524 1996
rect 1518 1991 1524 1992
rect 1558 1996 1564 1997
rect 1558 1992 1559 1996
rect 1563 1992 1564 1996
rect 1558 1991 1564 1992
rect 1598 1996 1604 1997
rect 1598 1992 1599 1996
rect 1603 1992 1604 1996
rect 1598 1991 1604 1992
rect 1638 1996 1644 1997
rect 1638 1992 1639 1996
rect 1643 1992 1644 1996
rect 1638 1991 1644 1992
rect 1678 1996 1684 1997
rect 1678 1992 1679 1996
rect 1683 1992 1684 1996
rect 1678 1991 1684 1992
rect 1718 1996 1724 1997
rect 1718 1992 1719 1996
rect 1723 1992 1724 1996
rect 1718 1991 1724 1992
rect 1766 1996 1772 1997
rect 1766 1992 1767 1996
rect 1771 1992 1772 1996
rect 1766 1991 1772 1992
rect 1822 1996 1828 1997
rect 1822 1992 1823 1996
rect 1827 1992 1828 1996
rect 1822 1991 1828 1992
rect 1870 1996 1876 1997
rect 1870 1992 1871 1996
rect 1875 1992 1876 1996
rect 1870 1991 1876 1992
rect 1918 1996 1924 1997
rect 1918 1992 1919 1996
rect 1923 1992 1924 1996
rect 1918 1991 1924 1992
rect 1966 1996 1972 1997
rect 1966 1992 1967 1996
rect 1971 1992 1972 1996
rect 1966 1991 1972 1992
rect 2014 1996 2020 1997
rect 2014 1992 2015 1996
rect 2019 1992 2020 1996
rect 2014 1991 2020 1992
rect 2054 1996 2060 1997
rect 2054 1992 2055 1996
rect 2059 1992 2060 1996
rect 2054 1991 2060 1992
rect 2094 1996 2100 1997
rect 2094 1992 2095 1996
rect 2099 1992 2100 1996
rect 2094 1991 2100 1992
rect 2142 1996 2148 1997
rect 2142 1992 2143 1996
rect 2147 1992 2148 1996
rect 2142 1991 2148 1992
rect 2190 1996 2196 1997
rect 2190 1992 2191 1996
rect 2195 1992 2196 1996
rect 2190 1991 2196 1992
rect 2238 1996 2244 1997
rect 2238 1992 2239 1996
rect 2243 1992 2244 1996
rect 2238 1991 2244 1992
rect 2278 1996 2284 1997
rect 2278 1992 2279 1996
rect 2283 1992 2284 1996
rect 2278 1991 2284 1992
rect 2318 1996 2324 1997
rect 2318 1992 2319 1996
rect 2323 1992 2324 1996
rect 2318 1991 2324 1992
rect 2358 1996 2364 1997
rect 2358 1992 2359 1996
rect 2363 1992 2364 1996
rect 2358 1991 2364 1992
rect 2408 1990 2410 1997
rect 1278 1989 1284 1990
rect 111 1986 115 1987
rect 111 1981 115 1982
rect 135 1986 139 1987
rect 135 1981 139 1982
rect 175 1986 179 1987
rect 175 1981 179 1982
rect 215 1986 219 1987
rect 215 1981 219 1982
rect 271 1986 275 1987
rect 271 1981 275 1982
rect 279 1986 283 1987
rect 279 1981 283 1982
rect 343 1986 347 1987
rect 343 1981 347 1982
rect 351 1986 355 1987
rect 351 1981 355 1982
rect 415 1986 419 1987
rect 415 1981 419 1982
rect 423 1986 427 1987
rect 423 1981 427 1982
rect 487 1986 491 1987
rect 487 1981 491 1982
rect 495 1986 499 1987
rect 495 1981 499 1982
rect 551 1986 555 1987
rect 551 1981 555 1982
rect 575 1986 579 1987
rect 575 1981 579 1982
rect 615 1986 619 1987
rect 615 1981 619 1982
rect 647 1986 651 1987
rect 647 1981 651 1982
rect 679 1986 683 1987
rect 679 1981 683 1982
rect 719 1986 723 1987
rect 719 1981 723 1982
rect 743 1986 747 1987
rect 743 1981 747 1982
rect 791 1986 795 1987
rect 791 1981 795 1982
rect 815 1986 819 1987
rect 815 1981 819 1982
rect 863 1986 867 1987
rect 863 1981 867 1982
rect 935 1986 939 1987
rect 935 1981 939 1982
rect 1007 1986 1011 1987
rect 1007 1981 1011 1982
rect 1239 1986 1243 1987
rect 1278 1985 1279 1989
rect 1283 1985 1284 1989
rect 1278 1984 1284 1985
rect 2406 1989 2412 1990
rect 2406 1985 2407 1989
rect 2411 1985 2412 1989
rect 2406 1984 2412 1985
rect 1239 1981 1243 1982
rect 112 1974 114 1981
rect 134 1980 140 1981
rect 134 1976 135 1980
rect 139 1976 140 1980
rect 134 1975 140 1976
rect 174 1980 180 1981
rect 174 1976 175 1980
rect 179 1976 180 1980
rect 174 1975 180 1976
rect 214 1980 220 1981
rect 214 1976 215 1980
rect 219 1976 220 1980
rect 214 1975 220 1976
rect 270 1980 276 1981
rect 270 1976 271 1980
rect 275 1976 276 1980
rect 270 1975 276 1976
rect 342 1980 348 1981
rect 342 1976 343 1980
rect 347 1976 348 1980
rect 342 1975 348 1976
rect 414 1980 420 1981
rect 414 1976 415 1980
rect 419 1976 420 1980
rect 414 1975 420 1976
rect 494 1980 500 1981
rect 494 1976 495 1980
rect 499 1976 500 1980
rect 494 1975 500 1976
rect 574 1980 580 1981
rect 574 1976 575 1980
rect 579 1976 580 1980
rect 574 1975 580 1976
rect 646 1980 652 1981
rect 646 1976 647 1980
rect 651 1976 652 1980
rect 646 1975 652 1976
rect 718 1980 724 1981
rect 718 1976 719 1980
rect 723 1976 724 1980
rect 718 1975 724 1976
rect 790 1980 796 1981
rect 790 1976 791 1980
rect 795 1976 796 1980
rect 790 1975 796 1976
rect 862 1980 868 1981
rect 862 1976 863 1980
rect 867 1976 868 1980
rect 862 1975 868 1976
rect 934 1980 940 1981
rect 934 1976 935 1980
rect 939 1976 940 1980
rect 934 1975 940 1976
rect 1006 1980 1012 1981
rect 1006 1976 1007 1980
rect 1011 1976 1012 1980
rect 1006 1975 1012 1976
rect 1240 1974 1242 1981
rect 110 1973 116 1974
rect 110 1969 111 1973
rect 115 1969 116 1973
rect 110 1968 116 1969
rect 1238 1973 1244 1974
rect 1238 1969 1239 1973
rect 1243 1969 1244 1973
rect 1238 1968 1244 1969
rect 1278 1972 1284 1973
rect 1278 1968 1279 1972
rect 1283 1968 1284 1972
rect 1278 1967 1284 1968
rect 2406 1972 2412 1973
rect 2406 1968 2407 1972
rect 2411 1968 2412 1972
rect 2406 1967 2412 1968
rect 110 1956 116 1957
rect 110 1952 111 1956
rect 115 1952 116 1956
rect 110 1951 116 1952
rect 1238 1956 1244 1957
rect 1238 1952 1239 1956
rect 1243 1952 1244 1956
rect 1238 1951 1244 1952
rect 112 1915 114 1951
rect 134 1933 140 1934
rect 134 1929 135 1933
rect 139 1929 140 1933
rect 134 1928 140 1929
rect 174 1933 180 1934
rect 174 1929 175 1933
rect 179 1929 180 1933
rect 174 1928 180 1929
rect 214 1933 220 1934
rect 214 1929 215 1933
rect 219 1929 220 1933
rect 214 1928 220 1929
rect 270 1933 276 1934
rect 270 1929 271 1933
rect 275 1929 276 1933
rect 270 1928 276 1929
rect 342 1933 348 1934
rect 342 1929 343 1933
rect 347 1929 348 1933
rect 342 1928 348 1929
rect 414 1933 420 1934
rect 414 1929 415 1933
rect 419 1929 420 1933
rect 414 1928 420 1929
rect 494 1933 500 1934
rect 494 1929 495 1933
rect 499 1929 500 1933
rect 494 1928 500 1929
rect 574 1933 580 1934
rect 574 1929 575 1933
rect 579 1929 580 1933
rect 574 1928 580 1929
rect 646 1933 652 1934
rect 646 1929 647 1933
rect 651 1929 652 1933
rect 646 1928 652 1929
rect 718 1933 724 1934
rect 718 1929 719 1933
rect 723 1929 724 1933
rect 718 1928 724 1929
rect 790 1933 796 1934
rect 790 1929 791 1933
rect 795 1929 796 1933
rect 790 1928 796 1929
rect 862 1933 868 1934
rect 862 1929 863 1933
rect 867 1929 868 1933
rect 862 1928 868 1929
rect 934 1933 940 1934
rect 934 1929 935 1933
rect 939 1929 940 1933
rect 934 1928 940 1929
rect 1006 1933 1012 1934
rect 1006 1929 1007 1933
rect 1011 1929 1012 1933
rect 1006 1928 1012 1929
rect 136 1915 138 1928
rect 176 1915 178 1928
rect 216 1915 218 1928
rect 272 1915 274 1928
rect 344 1915 346 1928
rect 416 1915 418 1928
rect 496 1915 498 1928
rect 576 1915 578 1928
rect 648 1915 650 1928
rect 720 1915 722 1928
rect 792 1915 794 1928
rect 864 1915 866 1928
rect 936 1915 938 1928
rect 1008 1915 1010 1928
rect 1240 1915 1242 1951
rect 1280 1931 1282 1967
rect 1398 1949 1404 1950
rect 1398 1945 1399 1949
rect 1403 1945 1404 1949
rect 1398 1944 1404 1945
rect 1438 1949 1444 1950
rect 1438 1945 1439 1949
rect 1443 1945 1444 1949
rect 1438 1944 1444 1945
rect 1478 1949 1484 1950
rect 1478 1945 1479 1949
rect 1483 1945 1484 1949
rect 1478 1944 1484 1945
rect 1518 1949 1524 1950
rect 1518 1945 1519 1949
rect 1523 1945 1524 1949
rect 1518 1944 1524 1945
rect 1558 1949 1564 1950
rect 1558 1945 1559 1949
rect 1563 1945 1564 1949
rect 1558 1944 1564 1945
rect 1598 1949 1604 1950
rect 1598 1945 1599 1949
rect 1603 1945 1604 1949
rect 1598 1944 1604 1945
rect 1638 1949 1644 1950
rect 1638 1945 1639 1949
rect 1643 1945 1644 1949
rect 1638 1944 1644 1945
rect 1678 1949 1684 1950
rect 1678 1945 1679 1949
rect 1683 1945 1684 1949
rect 1678 1944 1684 1945
rect 1718 1949 1724 1950
rect 1718 1945 1719 1949
rect 1723 1945 1724 1949
rect 1718 1944 1724 1945
rect 1766 1949 1772 1950
rect 1766 1945 1767 1949
rect 1771 1945 1772 1949
rect 1766 1944 1772 1945
rect 1822 1949 1828 1950
rect 1822 1945 1823 1949
rect 1827 1945 1828 1949
rect 1822 1944 1828 1945
rect 1870 1949 1876 1950
rect 1870 1945 1871 1949
rect 1875 1945 1876 1949
rect 1870 1944 1876 1945
rect 1918 1949 1924 1950
rect 1918 1945 1919 1949
rect 1923 1945 1924 1949
rect 1918 1944 1924 1945
rect 1966 1949 1972 1950
rect 1966 1945 1967 1949
rect 1971 1945 1972 1949
rect 1966 1944 1972 1945
rect 2014 1949 2020 1950
rect 2014 1945 2015 1949
rect 2019 1945 2020 1949
rect 2014 1944 2020 1945
rect 2054 1949 2060 1950
rect 2054 1945 2055 1949
rect 2059 1945 2060 1949
rect 2054 1944 2060 1945
rect 2094 1949 2100 1950
rect 2094 1945 2095 1949
rect 2099 1945 2100 1949
rect 2094 1944 2100 1945
rect 2142 1949 2148 1950
rect 2142 1945 2143 1949
rect 2147 1945 2148 1949
rect 2142 1944 2148 1945
rect 2190 1949 2196 1950
rect 2190 1945 2191 1949
rect 2195 1945 2196 1949
rect 2190 1944 2196 1945
rect 2238 1949 2244 1950
rect 2238 1945 2239 1949
rect 2243 1945 2244 1949
rect 2238 1944 2244 1945
rect 2278 1949 2284 1950
rect 2278 1945 2279 1949
rect 2283 1945 2284 1949
rect 2278 1944 2284 1945
rect 2318 1949 2324 1950
rect 2318 1945 2319 1949
rect 2323 1945 2324 1949
rect 2318 1944 2324 1945
rect 2358 1949 2364 1950
rect 2358 1945 2359 1949
rect 2363 1945 2364 1949
rect 2358 1944 2364 1945
rect 1400 1931 1402 1944
rect 1440 1931 1442 1944
rect 1480 1931 1482 1944
rect 1520 1931 1522 1944
rect 1560 1931 1562 1944
rect 1600 1931 1602 1944
rect 1640 1931 1642 1944
rect 1680 1931 1682 1944
rect 1720 1931 1722 1944
rect 1768 1931 1770 1944
rect 1824 1931 1826 1944
rect 1872 1931 1874 1944
rect 1920 1931 1922 1944
rect 1968 1931 1970 1944
rect 2016 1931 2018 1944
rect 2056 1931 2058 1944
rect 2096 1931 2098 1944
rect 2144 1931 2146 1944
rect 2192 1931 2194 1944
rect 2240 1931 2242 1944
rect 2280 1931 2282 1944
rect 2320 1931 2322 1944
rect 2360 1931 2362 1944
rect 2408 1931 2410 1967
rect 1279 1930 1283 1931
rect 1279 1925 1283 1926
rect 1343 1930 1347 1931
rect 1343 1925 1347 1926
rect 1383 1930 1387 1931
rect 1383 1925 1387 1926
rect 1399 1930 1403 1931
rect 1399 1925 1403 1926
rect 1423 1930 1427 1931
rect 1423 1925 1427 1926
rect 1439 1930 1443 1931
rect 1439 1925 1443 1926
rect 1463 1930 1467 1931
rect 1463 1925 1467 1926
rect 1479 1930 1483 1931
rect 1479 1925 1483 1926
rect 1511 1930 1515 1931
rect 1511 1925 1515 1926
rect 1519 1930 1523 1931
rect 1519 1925 1523 1926
rect 1559 1930 1563 1931
rect 1559 1925 1563 1926
rect 1567 1930 1571 1931
rect 1567 1925 1571 1926
rect 1599 1930 1603 1931
rect 1599 1925 1603 1926
rect 1631 1930 1635 1931
rect 1631 1925 1635 1926
rect 1639 1930 1643 1931
rect 1639 1925 1643 1926
rect 1679 1930 1683 1931
rect 1679 1925 1683 1926
rect 1711 1930 1715 1931
rect 1711 1925 1715 1926
rect 1719 1930 1723 1931
rect 1719 1925 1723 1926
rect 1767 1930 1771 1931
rect 1767 1925 1771 1926
rect 1807 1930 1811 1931
rect 1807 1925 1811 1926
rect 1823 1930 1827 1931
rect 1823 1925 1827 1926
rect 1871 1930 1875 1931
rect 1871 1925 1875 1926
rect 1919 1930 1923 1931
rect 1919 1925 1923 1926
rect 1967 1930 1971 1931
rect 1967 1925 1971 1926
rect 2015 1930 2019 1931
rect 2015 1925 2019 1926
rect 2031 1930 2035 1931
rect 2031 1925 2035 1926
rect 2055 1930 2059 1931
rect 2055 1925 2059 1926
rect 2095 1930 2099 1931
rect 2095 1925 2099 1926
rect 2143 1930 2147 1931
rect 2143 1925 2147 1926
rect 2151 1930 2155 1931
rect 2151 1925 2155 1926
rect 2191 1930 2195 1931
rect 2191 1925 2195 1926
rect 2239 1930 2243 1931
rect 2239 1925 2243 1926
rect 2279 1930 2283 1931
rect 2279 1925 2283 1926
rect 2319 1930 2323 1931
rect 2319 1925 2323 1926
rect 2359 1930 2363 1931
rect 2359 1925 2363 1926
rect 2407 1930 2411 1931
rect 2407 1925 2411 1926
rect 111 1914 115 1915
rect 111 1909 115 1910
rect 135 1914 139 1915
rect 135 1909 139 1910
rect 175 1914 179 1915
rect 175 1909 179 1910
rect 215 1914 219 1915
rect 215 1909 219 1910
rect 247 1914 251 1915
rect 247 1909 251 1910
rect 271 1914 275 1915
rect 271 1909 275 1910
rect 287 1914 291 1915
rect 287 1909 291 1910
rect 327 1914 331 1915
rect 327 1909 331 1910
rect 343 1914 347 1915
rect 343 1909 347 1910
rect 367 1914 371 1915
rect 367 1909 371 1910
rect 415 1914 419 1915
rect 415 1909 419 1910
rect 471 1914 475 1915
rect 471 1909 475 1910
rect 495 1914 499 1915
rect 495 1909 499 1910
rect 535 1914 539 1915
rect 535 1909 539 1910
rect 575 1914 579 1915
rect 575 1909 579 1910
rect 599 1914 603 1915
rect 599 1909 603 1910
rect 647 1914 651 1915
rect 647 1909 651 1910
rect 663 1914 667 1915
rect 663 1909 667 1910
rect 719 1914 723 1915
rect 719 1909 723 1910
rect 727 1914 731 1915
rect 727 1909 731 1910
rect 791 1914 795 1915
rect 791 1909 795 1910
rect 855 1914 859 1915
rect 855 1909 859 1910
rect 863 1914 867 1915
rect 863 1909 867 1910
rect 919 1914 923 1915
rect 919 1909 923 1910
rect 935 1914 939 1915
rect 935 1909 939 1910
rect 983 1914 987 1915
rect 983 1909 987 1910
rect 1007 1914 1011 1915
rect 1007 1909 1011 1910
rect 1055 1914 1059 1915
rect 1055 1909 1059 1910
rect 1127 1914 1131 1915
rect 1127 1909 1131 1910
rect 1239 1914 1243 1915
rect 1239 1909 1243 1910
rect 112 1877 114 1909
rect 248 1900 250 1909
rect 288 1900 290 1909
rect 328 1900 330 1909
rect 368 1900 370 1909
rect 416 1900 418 1909
rect 472 1900 474 1909
rect 536 1900 538 1909
rect 600 1900 602 1909
rect 664 1900 666 1909
rect 728 1900 730 1909
rect 792 1900 794 1909
rect 856 1900 858 1909
rect 920 1900 922 1909
rect 984 1900 986 1909
rect 1056 1900 1058 1909
rect 1128 1900 1130 1909
rect 246 1899 252 1900
rect 246 1895 247 1899
rect 251 1895 252 1899
rect 246 1894 252 1895
rect 286 1899 292 1900
rect 286 1895 287 1899
rect 291 1895 292 1899
rect 286 1894 292 1895
rect 326 1899 332 1900
rect 326 1895 327 1899
rect 331 1895 332 1899
rect 326 1894 332 1895
rect 366 1899 372 1900
rect 366 1895 367 1899
rect 371 1895 372 1899
rect 366 1894 372 1895
rect 414 1899 420 1900
rect 414 1895 415 1899
rect 419 1895 420 1899
rect 414 1894 420 1895
rect 470 1899 476 1900
rect 470 1895 471 1899
rect 475 1895 476 1899
rect 470 1894 476 1895
rect 534 1899 540 1900
rect 534 1895 535 1899
rect 539 1895 540 1899
rect 534 1894 540 1895
rect 598 1899 604 1900
rect 598 1895 599 1899
rect 603 1895 604 1899
rect 598 1894 604 1895
rect 662 1899 668 1900
rect 662 1895 663 1899
rect 667 1895 668 1899
rect 662 1894 668 1895
rect 726 1899 732 1900
rect 726 1895 727 1899
rect 731 1895 732 1899
rect 726 1894 732 1895
rect 790 1899 796 1900
rect 790 1895 791 1899
rect 795 1895 796 1899
rect 790 1894 796 1895
rect 854 1899 860 1900
rect 854 1895 855 1899
rect 859 1895 860 1899
rect 854 1894 860 1895
rect 918 1899 924 1900
rect 918 1895 919 1899
rect 923 1895 924 1899
rect 918 1894 924 1895
rect 982 1899 988 1900
rect 982 1895 983 1899
rect 987 1895 988 1899
rect 982 1894 988 1895
rect 1054 1899 1060 1900
rect 1054 1895 1055 1899
rect 1059 1895 1060 1899
rect 1054 1894 1060 1895
rect 1126 1899 1132 1900
rect 1126 1895 1127 1899
rect 1131 1895 1132 1899
rect 1126 1894 1132 1895
rect 1240 1877 1242 1909
rect 1280 1893 1282 1925
rect 1344 1916 1346 1925
rect 1384 1916 1386 1925
rect 1424 1916 1426 1925
rect 1464 1916 1466 1925
rect 1512 1916 1514 1925
rect 1568 1916 1570 1925
rect 1632 1916 1634 1925
rect 1712 1916 1714 1925
rect 1808 1916 1810 1925
rect 1920 1916 1922 1925
rect 2032 1916 2034 1925
rect 2152 1916 2154 1925
rect 1342 1915 1348 1916
rect 1342 1911 1343 1915
rect 1347 1911 1348 1915
rect 1342 1910 1348 1911
rect 1382 1915 1388 1916
rect 1382 1911 1383 1915
rect 1387 1911 1388 1915
rect 1382 1910 1388 1911
rect 1422 1915 1428 1916
rect 1422 1911 1423 1915
rect 1427 1911 1428 1915
rect 1422 1910 1428 1911
rect 1462 1915 1468 1916
rect 1462 1911 1463 1915
rect 1467 1911 1468 1915
rect 1462 1910 1468 1911
rect 1510 1915 1516 1916
rect 1510 1911 1511 1915
rect 1515 1911 1516 1915
rect 1510 1910 1516 1911
rect 1566 1915 1572 1916
rect 1566 1911 1567 1915
rect 1571 1911 1572 1915
rect 1566 1910 1572 1911
rect 1630 1915 1636 1916
rect 1630 1911 1631 1915
rect 1635 1911 1636 1915
rect 1630 1910 1636 1911
rect 1710 1915 1716 1916
rect 1710 1911 1711 1915
rect 1715 1911 1716 1915
rect 1710 1910 1716 1911
rect 1806 1915 1812 1916
rect 1806 1911 1807 1915
rect 1811 1911 1812 1915
rect 1806 1910 1812 1911
rect 1918 1915 1924 1916
rect 1918 1911 1919 1915
rect 1923 1911 1924 1915
rect 1918 1910 1924 1911
rect 2030 1915 2036 1916
rect 2030 1911 2031 1915
rect 2035 1911 2036 1915
rect 2030 1910 2036 1911
rect 2150 1915 2156 1916
rect 2150 1911 2151 1915
rect 2155 1911 2156 1915
rect 2150 1910 2156 1911
rect 2408 1893 2410 1925
rect 1278 1892 1284 1893
rect 1278 1888 1279 1892
rect 1283 1888 1284 1892
rect 1278 1887 1284 1888
rect 2406 1892 2412 1893
rect 2406 1888 2407 1892
rect 2411 1888 2412 1892
rect 2406 1887 2412 1888
rect 110 1876 116 1877
rect 110 1872 111 1876
rect 115 1872 116 1876
rect 110 1871 116 1872
rect 1238 1876 1244 1877
rect 1238 1872 1239 1876
rect 1243 1872 1244 1876
rect 1238 1871 1244 1872
rect 1278 1875 1284 1876
rect 1278 1871 1279 1875
rect 1283 1871 1284 1875
rect 1278 1870 1284 1871
rect 2406 1875 2412 1876
rect 2406 1871 2407 1875
rect 2411 1871 2412 1875
rect 2406 1870 2412 1871
rect 110 1859 116 1860
rect 110 1855 111 1859
rect 115 1855 116 1859
rect 110 1854 116 1855
rect 1238 1859 1244 1860
rect 1238 1855 1239 1859
rect 1243 1855 1244 1859
rect 1280 1855 1282 1870
rect 1342 1868 1348 1869
rect 1342 1864 1343 1868
rect 1347 1864 1348 1868
rect 1342 1863 1348 1864
rect 1382 1868 1388 1869
rect 1382 1864 1383 1868
rect 1387 1864 1388 1868
rect 1382 1863 1388 1864
rect 1422 1868 1428 1869
rect 1422 1864 1423 1868
rect 1427 1864 1428 1868
rect 1422 1863 1428 1864
rect 1462 1868 1468 1869
rect 1462 1864 1463 1868
rect 1467 1864 1468 1868
rect 1462 1863 1468 1864
rect 1510 1868 1516 1869
rect 1510 1864 1511 1868
rect 1515 1864 1516 1868
rect 1510 1863 1516 1864
rect 1566 1868 1572 1869
rect 1566 1864 1567 1868
rect 1571 1864 1572 1868
rect 1566 1863 1572 1864
rect 1630 1868 1636 1869
rect 1630 1864 1631 1868
rect 1635 1864 1636 1868
rect 1630 1863 1636 1864
rect 1710 1868 1716 1869
rect 1710 1864 1711 1868
rect 1715 1864 1716 1868
rect 1710 1863 1716 1864
rect 1806 1868 1812 1869
rect 1806 1864 1807 1868
rect 1811 1864 1812 1868
rect 1806 1863 1812 1864
rect 1918 1868 1924 1869
rect 1918 1864 1919 1868
rect 1923 1864 1924 1868
rect 1918 1863 1924 1864
rect 2030 1868 2036 1869
rect 2030 1864 2031 1868
rect 2035 1864 2036 1868
rect 2030 1863 2036 1864
rect 2150 1868 2156 1869
rect 2150 1864 2151 1868
rect 2155 1864 2156 1868
rect 2150 1863 2156 1864
rect 1344 1855 1346 1863
rect 1384 1855 1386 1863
rect 1424 1855 1426 1863
rect 1464 1855 1466 1863
rect 1512 1855 1514 1863
rect 1568 1855 1570 1863
rect 1632 1855 1634 1863
rect 1712 1855 1714 1863
rect 1808 1855 1810 1863
rect 1920 1855 1922 1863
rect 2032 1855 2034 1863
rect 2152 1855 2154 1863
rect 2408 1855 2410 1870
rect 1238 1854 1244 1855
rect 1279 1854 1283 1855
rect 112 1843 114 1854
rect 246 1852 252 1853
rect 246 1848 247 1852
rect 251 1848 252 1852
rect 246 1847 252 1848
rect 286 1852 292 1853
rect 286 1848 287 1852
rect 291 1848 292 1852
rect 286 1847 292 1848
rect 326 1852 332 1853
rect 326 1848 327 1852
rect 331 1848 332 1852
rect 326 1847 332 1848
rect 366 1852 372 1853
rect 366 1848 367 1852
rect 371 1848 372 1852
rect 366 1847 372 1848
rect 414 1852 420 1853
rect 414 1848 415 1852
rect 419 1848 420 1852
rect 414 1847 420 1848
rect 470 1852 476 1853
rect 470 1848 471 1852
rect 475 1848 476 1852
rect 470 1847 476 1848
rect 534 1852 540 1853
rect 534 1848 535 1852
rect 539 1848 540 1852
rect 534 1847 540 1848
rect 598 1852 604 1853
rect 598 1848 599 1852
rect 603 1848 604 1852
rect 598 1847 604 1848
rect 662 1852 668 1853
rect 662 1848 663 1852
rect 667 1848 668 1852
rect 662 1847 668 1848
rect 726 1852 732 1853
rect 726 1848 727 1852
rect 731 1848 732 1852
rect 726 1847 732 1848
rect 790 1852 796 1853
rect 790 1848 791 1852
rect 795 1848 796 1852
rect 790 1847 796 1848
rect 854 1852 860 1853
rect 854 1848 855 1852
rect 859 1848 860 1852
rect 854 1847 860 1848
rect 918 1852 924 1853
rect 918 1848 919 1852
rect 923 1848 924 1852
rect 918 1847 924 1848
rect 982 1852 988 1853
rect 982 1848 983 1852
rect 987 1848 988 1852
rect 982 1847 988 1848
rect 1054 1852 1060 1853
rect 1054 1848 1055 1852
rect 1059 1848 1060 1852
rect 1054 1847 1060 1848
rect 1126 1852 1132 1853
rect 1126 1848 1127 1852
rect 1131 1848 1132 1852
rect 1126 1847 1132 1848
rect 248 1843 250 1847
rect 288 1843 290 1847
rect 328 1843 330 1847
rect 368 1843 370 1847
rect 416 1843 418 1847
rect 472 1843 474 1847
rect 536 1843 538 1847
rect 600 1843 602 1847
rect 664 1843 666 1847
rect 728 1843 730 1847
rect 792 1843 794 1847
rect 856 1843 858 1847
rect 920 1843 922 1847
rect 984 1843 986 1847
rect 1056 1843 1058 1847
rect 1128 1843 1130 1847
rect 1240 1843 1242 1854
rect 1279 1849 1283 1850
rect 1343 1854 1347 1855
rect 1343 1849 1347 1850
rect 1359 1854 1363 1855
rect 1359 1849 1363 1850
rect 1383 1854 1387 1855
rect 1383 1849 1387 1850
rect 1399 1854 1403 1855
rect 1399 1849 1403 1850
rect 1423 1854 1427 1855
rect 1423 1849 1427 1850
rect 1447 1854 1451 1855
rect 1447 1849 1451 1850
rect 1463 1854 1467 1855
rect 1463 1849 1467 1850
rect 1503 1854 1507 1855
rect 1503 1849 1507 1850
rect 1511 1854 1515 1855
rect 1511 1849 1515 1850
rect 1559 1854 1563 1855
rect 1559 1849 1563 1850
rect 1567 1854 1571 1855
rect 1567 1849 1571 1850
rect 1615 1854 1619 1855
rect 1615 1849 1619 1850
rect 1631 1854 1635 1855
rect 1631 1849 1635 1850
rect 1671 1854 1675 1855
rect 1671 1849 1675 1850
rect 1711 1854 1715 1855
rect 1711 1849 1715 1850
rect 1727 1854 1731 1855
rect 1727 1849 1731 1850
rect 1783 1854 1787 1855
rect 1783 1849 1787 1850
rect 1807 1854 1811 1855
rect 1807 1849 1811 1850
rect 1839 1854 1843 1855
rect 1839 1849 1843 1850
rect 1895 1854 1899 1855
rect 1895 1849 1899 1850
rect 1919 1854 1923 1855
rect 1919 1849 1923 1850
rect 1951 1854 1955 1855
rect 1951 1849 1955 1850
rect 2031 1854 2035 1855
rect 2031 1849 2035 1850
rect 2151 1854 2155 1855
rect 2151 1849 2155 1850
rect 2407 1854 2411 1855
rect 2407 1849 2411 1850
rect 111 1842 115 1843
rect 111 1837 115 1838
rect 247 1842 251 1843
rect 247 1837 251 1838
rect 287 1842 291 1843
rect 287 1837 291 1838
rect 327 1842 331 1843
rect 327 1837 331 1838
rect 367 1842 371 1843
rect 367 1837 371 1838
rect 399 1842 403 1843
rect 399 1837 403 1838
rect 415 1842 419 1843
rect 415 1837 419 1838
rect 439 1842 443 1843
rect 439 1837 443 1838
rect 471 1842 475 1843
rect 471 1837 475 1838
rect 479 1842 483 1843
rect 479 1837 483 1838
rect 519 1842 523 1843
rect 519 1837 523 1838
rect 535 1842 539 1843
rect 535 1837 539 1838
rect 567 1842 571 1843
rect 567 1837 571 1838
rect 599 1842 603 1843
rect 599 1837 603 1838
rect 623 1842 627 1843
rect 623 1837 627 1838
rect 663 1842 667 1843
rect 663 1837 667 1838
rect 687 1842 691 1843
rect 687 1837 691 1838
rect 727 1842 731 1843
rect 727 1837 731 1838
rect 759 1842 763 1843
rect 759 1837 763 1838
rect 791 1842 795 1843
rect 791 1837 795 1838
rect 831 1842 835 1843
rect 831 1837 835 1838
rect 855 1842 859 1843
rect 855 1837 859 1838
rect 903 1842 907 1843
rect 903 1837 907 1838
rect 919 1842 923 1843
rect 919 1837 923 1838
rect 975 1842 979 1843
rect 975 1837 979 1838
rect 983 1842 987 1843
rect 983 1837 987 1838
rect 1047 1842 1051 1843
rect 1047 1837 1051 1838
rect 1055 1842 1059 1843
rect 1055 1837 1059 1838
rect 1127 1842 1131 1843
rect 1127 1837 1131 1838
rect 1191 1842 1195 1843
rect 1191 1837 1195 1838
rect 1239 1842 1243 1843
rect 1280 1842 1282 1849
rect 1358 1848 1364 1849
rect 1358 1844 1359 1848
rect 1363 1844 1364 1848
rect 1358 1843 1364 1844
rect 1398 1848 1404 1849
rect 1398 1844 1399 1848
rect 1403 1844 1404 1848
rect 1398 1843 1404 1844
rect 1446 1848 1452 1849
rect 1446 1844 1447 1848
rect 1451 1844 1452 1848
rect 1446 1843 1452 1844
rect 1502 1848 1508 1849
rect 1502 1844 1503 1848
rect 1507 1844 1508 1848
rect 1502 1843 1508 1844
rect 1558 1848 1564 1849
rect 1558 1844 1559 1848
rect 1563 1844 1564 1848
rect 1558 1843 1564 1844
rect 1614 1848 1620 1849
rect 1614 1844 1615 1848
rect 1619 1844 1620 1848
rect 1614 1843 1620 1844
rect 1670 1848 1676 1849
rect 1670 1844 1671 1848
rect 1675 1844 1676 1848
rect 1670 1843 1676 1844
rect 1726 1848 1732 1849
rect 1726 1844 1727 1848
rect 1731 1844 1732 1848
rect 1726 1843 1732 1844
rect 1782 1848 1788 1849
rect 1782 1844 1783 1848
rect 1787 1844 1788 1848
rect 1782 1843 1788 1844
rect 1838 1848 1844 1849
rect 1838 1844 1839 1848
rect 1843 1844 1844 1848
rect 1838 1843 1844 1844
rect 1894 1848 1900 1849
rect 1894 1844 1895 1848
rect 1899 1844 1900 1848
rect 1894 1843 1900 1844
rect 1950 1848 1956 1849
rect 1950 1844 1951 1848
rect 1955 1844 1956 1848
rect 1950 1843 1956 1844
rect 2408 1842 2410 1849
rect 1239 1837 1243 1838
rect 1278 1841 1284 1842
rect 1278 1837 1279 1841
rect 1283 1837 1284 1841
rect 112 1830 114 1837
rect 398 1836 404 1837
rect 398 1832 399 1836
rect 403 1832 404 1836
rect 398 1831 404 1832
rect 438 1836 444 1837
rect 438 1832 439 1836
rect 443 1832 444 1836
rect 438 1831 444 1832
rect 478 1836 484 1837
rect 478 1832 479 1836
rect 483 1832 484 1836
rect 478 1831 484 1832
rect 518 1836 524 1837
rect 518 1832 519 1836
rect 523 1832 524 1836
rect 518 1831 524 1832
rect 566 1836 572 1837
rect 566 1832 567 1836
rect 571 1832 572 1836
rect 566 1831 572 1832
rect 622 1836 628 1837
rect 622 1832 623 1836
rect 627 1832 628 1836
rect 622 1831 628 1832
rect 686 1836 692 1837
rect 686 1832 687 1836
rect 691 1832 692 1836
rect 686 1831 692 1832
rect 758 1836 764 1837
rect 758 1832 759 1836
rect 763 1832 764 1836
rect 758 1831 764 1832
rect 830 1836 836 1837
rect 830 1832 831 1836
rect 835 1832 836 1836
rect 830 1831 836 1832
rect 902 1836 908 1837
rect 902 1832 903 1836
rect 907 1832 908 1836
rect 902 1831 908 1832
rect 974 1836 980 1837
rect 974 1832 975 1836
rect 979 1832 980 1836
rect 974 1831 980 1832
rect 1046 1836 1052 1837
rect 1046 1832 1047 1836
rect 1051 1832 1052 1836
rect 1046 1831 1052 1832
rect 1126 1836 1132 1837
rect 1126 1832 1127 1836
rect 1131 1832 1132 1836
rect 1126 1831 1132 1832
rect 1190 1836 1196 1837
rect 1190 1832 1191 1836
rect 1195 1832 1196 1836
rect 1190 1831 1196 1832
rect 1240 1830 1242 1837
rect 1278 1836 1284 1837
rect 2406 1841 2412 1842
rect 2406 1837 2407 1841
rect 2411 1837 2412 1841
rect 2406 1836 2412 1837
rect 110 1829 116 1830
rect 110 1825 111 1829
rect 115 1825 116 1829
rect 110 1824 116 1825
rect 1238 1829 1244 1830
rect 1238 1825 1239 1829
rect 1243 1825 1244 1829
rect 1238 1824 1244 1825
rect 1278 1824 1284 1825
rect 1278 1820 1279 1824
rect 1283 1820 1284 1824
rect 1278 1819 1284 1820
rect 2406 1824 2412 1825
rect 2406 1820 2407 1824
rect 2411 1820 2412 1824
rect 2406 1819 2412 1820
rect 110 1812 116 1813
rect 110 1808 111 1812
rect 115 1808 116 1812
rect 110 1807 116 1808
rect 1238 1812 1244 1813
rect 1238 1808 1239 1812
rect 1243 1808 1244 1812
rect 1238 1807 1244 1808
rect 112 1775 114 1807
rect 398 1789 404 1790
rect 398 1785 399 1789
rect 403 1785 404 1789
rect 398 1784 404 1785
rect 438 1789 444 1790
rect 438 1785 439 1789
rect 443 1785 444 1789
rect 438 1784 444 1785
rect 478 1789 484 1790
rect 478 1785 479 1789
rect 483 1785 484 1789
rect 478 1784 484 1785
rect 518 1789 524 1790
rect 518 1785 519 1789
rect 523 1785 524 1789
rect 518 1784 524 1785
rect 566 1789 572 1790
rect 566 1785 567 1789
rect 571 1785 572 1789
rect 566 1784 572 1785
rect 622 1789 628 1790
rect 622 1785 623 1789
rect 627 1785 628 1789
rect 622 1784 628 1785
rect 686 1789 692 1790
rect 686 1785 687 1789
rect 691 1785 692 1789
rect 686 1784 692 1785
rect 758 1789 764 1790
rect 758 1785 759 1789
rect 763 1785 764 1789
rect 758 1784 764 1785
rect 830 1789 836 1790
rect 830 1785 831 1789
rect 835 1785 836 1789
rect 830 1784 836 1785
rect 902 1789 908 1790
rect 902 1785 903 1789
rect 907 1785 908 1789
rect 902 1784 908 1785
rect 974 1789 980 1790
rect 974 1785 975 1789
rect 979 1785 980 1789
rect 974 1784 980 1785
rect 1046 1789 1052 1790
rect 1046 1785 1047 1789
rect 1051 1785 1052 1789
rect 1046 1784 1052 1785
rect 1126 1789 1132 1790
rect 1126 1785 1127 1789
rect 1131 1785 1132 1789
rect 1126 1784 1132 1785
rect 1190 1789 1196 1790
rect 1190 1785 1191 1789
rect 1195 1785 1196 1789
rect 1190 1784 1196 1785
rect 400 1775 402 1784
rect 440 1775 442 1784
rect 480 1775 482 1784
rect 520 1775 522 1784
rect 568 1775 570 1784
rect 624 1775 626 1784
rect 688 1775 690 1784
rect 760 1775 762 1784
rect 832 1775 834 1784
rect 904 1775 906 1784
rect 976 1775 978 1784
rect 1048 1775 1050 1784
rect 1128 1775 1130 1784
rect 1192 1775 1194 1784
rect 1240 1775 1242 1807
rect 1280 1775 1282 1819
rect 1358 1801 1364 1802
rect 1358 1797 1359 1801
rect 1363 1797 1364 1801
rect 1358 1796 1364 1797
rect 1398 1801 1404 1802
rect 1398 1797 1399 1801
rect 1403 1797 1404 1801
rect 1398 1796 1404 1797
rect 1446 1801 1452 1802
rect 1446 1797 1447 1801
rect 1451 1797 1452 1801
rect 1446 1796 1452 1797
rect 1502 1801 1508 1802
rect 1502 1797 1503 1801
rect 1507 1797 1508 1801
rect 1502 1796 1508 1797
rect 1558 1801 1564 1802
rect 1558 1797 1559 1801
rect 1563 1797 1564 1801
rect 1558 1796 1564 1797
rect 1614 1801 1620 1802
rect 1614 1797 1615 1801
rect 1619 1797 1620 1801
rect 1614 1796 1620 1797
rect 1670 1801 1676 1802
rect 1670 1797 1671 1801
rect 1675 1797 1676 1801
rect 1670 1796 1676 1797
rect 1726 1801 1732 1802
rect 1726 1797 1727 1801
rect 1731 1797 1732 1801
rect 1726 1796 1732 1797
rect 1782 1801 1788 1802
rect 1782 1797 1783 1801
rect 1787 1797 1788 1801
rect 1782 1796 1788 1797
rect 1838 1801 1844 1802
rect 1838 1797 1839 1801
rect 1843 1797 1844 1801
rect 1838 1796 1844 1797
rect 1894 1801 1900 1802
rect 1894 1797 1895 1801
rect 1899 1797 1900 1801
rect 1894 1796 1900 1797
rect 1950 1801 1956 1802
rect 1950 1797 1951 1801
rect 1955 1797 1956 1801
rect 1950 1796 1956 1797
rect 1360 1775 1362 1796
rect 1400 1775 1402 1796
rect 1448 1775 1450 1796
rect 1504 1775 1506 1796
rect 1560 1775 1562 1796
rect 1616 1775 1618 1796
rect 1672 1775 1674 1796
rect 1728 1775 1730 1796
rect 1784 1775 1786 1796
rect 1840 1775 1842 1796
rect 1896 1775 1898 1796
rect 1952 1775 1954 1796
rect 2408 1775 2410 1819
rect 111 1774 115 1775
rect 111 1769 115 1770
rect 399 1774 403 1775
rect 399 1769 403 1770
rect 407 1774 411 1775
rect 407 1769 411 1770
rect 439 1774 443 1775
rect 439 1769 443 1770
rect 447 1774 451 1775
rect 447 1769 451 1770
rect 479 1774 483 1775
rect 479 1769 483 1770
rect 487 1774 491 1775
rect 487 1769 491 1770
rect 519 1774 523 1775
rect 519 1769 523 1770
rect 527 1774 531 1775
rect 527 1769 531 1770
rect 567 1774 571 1775
rect 567 1769 571 1770
rect 607 1774 611 1775
rect 607 1769 611 1770
rect 623 1774 627 1775
rect 623 1769 627 1770
rect 647 1774 651 1775
rect 647 1769 651 1770
rect 687 1774 691 1775
rect 687 1769 691 1770
rect 695 1774 699 1775
rect 695 1769 699 1770
rect 751 1774 755 1775
rect 751 1769 755 1770
rect 759 1774 763 1775
rect 759 1769 763 1770
rect 807 1774 811 1775
rect 807 1769 811 1770
rect 831 1774 835 1775
rect 831 1769 835 1770
rect 871 1774 875 1775
rect 871 1769 875 1770
rect 903 1774 907 1775
rect 903 1769 907 1770
rect 935 1774 939 1775
rect 935 1769 939 1770
rect 975 1774 979 1775
rect 975 1769 979 1770
rect 999 1774 1003 1775
rect 999 1769 1003 1770
rect 1047 1774 1051 1775
rect 1047 1769 1051 1770
rect 1071 1774 1075 1775
rect 1071 1769 1075 1770
rect 1127 1774 1131 1775
rect 1127 1769 1131 1770
rect 1143 1774 1147 1775
rect 1143 1769 1147 1770
rect 1191 1774 1195 1775
rect 1191 1769 1195 1770
rect 1239 1774 1243 1775
rect 1239 1769 1243 1770
rect 1279 1774 1283 1775
rect 1279 1769 1283 1770
rect 1303 1774 1307 1775
rect 1303 1769 1307 1770
rect 1343 1774 1347 1775
rect 1343 1769 1347 1770
rect 1359 1774 1363 1775
rect 1359 1769 1363 1770
rect 1391 1774 1395 1775
rect 1391 1769 1395 1770
rect 1399 1774 1403 1775
rect 1399 1769 1403 1770
rect 1447 1774 1451 1775
rect 1447 1769 1451 1770
rect 1455 1774 1459 1775
rect 1455 1769 1459 1770
rect 1503 1774 1507 1775
rect 1503 1769 1507 1770
rect 1519 1774 1523 1775
rect 1519 1769 1523 1770
rect 1559 1774 1563 1775
rect 1559 1769 1563 1770
rect 1583 1774 1587 1775
rect 1583 1769 1587 1770
rect 1615 1774 1619 1775
rect 1615 1769 1619 1770
rect 1647 1774 1651 1775
rect 1647 1769 1651 1770
rect 1671 1774 1675 1775
rect 1671 1769 1675 1770
rect 1703 1774 1707 1775
rect 1703 1769 1707 1770
rect 1727 1774 1731 1775
rect 1727 1769 1731 1770
rect 1759 1774 1763 1775
rect 1759 1769 1763 1770
rect 1783 1774 1787 1775
rect 1783 1769 1787 1770
rect 1807 1774 1811 1775
rect 1807 1769 1811 1770
rect 1839 1774 1843 1775
rect 1839 1769 1843 1770
rect 1863 1774 1867 1775
rect 1863 1769 1867 1770
rect 1895 1774 1899 1775
rect 1895 1769 1899 1770
rect 1919 1774 1923 1775
rect 1919 1769 1923 1770
rect 1951 1774 1955 1775
rect 1951 1769 1955 1770
rect 1975 1774 1979 1775
rect 1975 1769 1979 1770
rect 2407 1774 2411 1775
rect 2407 1769 2411 1770
rect 112 1737 114 1769
rect 408 1760 410 1769
rect 448 1760 450 1769
rect 488 1760 490 1769
rect 528 1760 530 1769
rect 568 1760 570 1769
rect 608 1760 610 1769
rect 648 1760 650 1769
rect 696 1760 698 1769
rect 752 1760 754 1769
rect 808 1760 810 1769
rect 872 1760 874 1769
rect 936 1760 938 1769
rect 1000 1760 1002 1769
rect 1072 1760 1074 1769
rect 1144 1760 1146 1769
rect 1192 1760 1194 1769
rect 406 1759 412 1760
rect 406 1755 407 1759
rect 411 1755 412 1759
rect 406 1754 412 1755
rect 446 1759 452 1760
rect 446 1755 447 1759
rect 451 1755 452 1759
rect 446 1754 452 1755
rect 486 1759 492 1760
rect 486 1755 487 1759
rect 491 1755 492 1759
rect 486 1754 492 1755
rect 526 1759 532 1760
rect 526 1755 527 1759
rect 531 1755 532 1759
rect 526 1754 532 1755
rect 566 1759 572 1760
rect 566 1755 567 1759
rect 571 1755 572 1759
rect 566 1754 572 1755
rect 606 1759 612 1760
rect 606 1755 607 1759
rect 611 1755 612 1759
rect 606 1754 612 1755
rect 646 1759 652 1760
rect 646 1755 647 1759
rect 651 1755 652 1759
rect 646 1754 652 1755
rect 694 1759 700 1760
rect 694 1755 695 1759
rect 699 1755 700 1759
rect 694 1754 700 1755
rect 750 1759 756 1760
rect 750 1755 751 1759
rect 755 1755 756 1759
rect 750 1754 756 1755
rect 806 1759 812 1760
rect 806 1755 807 1759
rect 811 1755 812 1759
rect 806 1754 812 1755
rect 870 1759 876 1760
rect 870 1755 871 1759
rect 875 1755 876 1759
rect 870 1754 876 1755
rect 934 1759 940 1760
rect 934 1755 935 1759
rect 939 1755 940 1759
rect 934 1754 940 1755
rect 998 1759 1004 1760
rect 998 1755 999 1759
rect 1003 1755 1004 1759
rect 998 1754 1004 1755
rect 1070 1759 1076 1760
rect 1070 1755 1071 1759
rect 1075 1755 1076 1759
rect 1070 1754 1076 1755
rect 1142 1759 1148 1760
rect 1142 1755 1143 1759
rect 1147 1755 1148 1759
rect 1142 1754 1148 1755
rect 1190 1759 1196 1760
rect 1190 1755 1191 1759
rect 1195 1755 1196 1759
rect 1190 1754 1196 1755
rect 1240 1737 1242 1769
rect 1280 1737 1282 1769
rect 1304 1760 1306 1769
rect 1344 1760 1346 1769
rect 1392 1760 1394 1769
rect 1456 1760 1458 1769
rect 1520 1760 1522 1769
rect 1584 1760 1586 1769
rect 1648 1760 1650 1769
rect 1704 1760 1706 1769
rect 1760 1760 1762 1769
rect 1808 1760 1810 1769
rect 1864 1760 1866 1769
rect 1920 1760 1922 1769
rect 1976 1760 1978 1769
rect 1302 1759 1308 1760
rect 1302 1755 1303 1759
rect 1307 1755 1308 1759
rect 1302 1754 1308 1755
rect 1342 1759 1348 1760
rect 1342 1755 1343 1759
rect 1347 1755 1348 1759
rect 1342 1754 1348 1755
rect 1390 1759 1396 1760
rect 1390 1755 1391 1759
rect 1395 1755 1396 1759
rect 1390 1754 1396 1755
rect 1454 1759 1460 1760
rect 1454 1755 1455 1759
rect 1459 1755 1460 1759
rect 1454 1754 1460 1755
rect 1518 1759 1524 1760
rect 1518 1755 1519 1759
rect 1523 1755 1524 1759
rect 1518 1754 1524 1755
rect 1582 1759 1588 1760
rect 1582 1755 1583 1759
rect 1587 1755 1588 1759
rect 1582 1754 1588 1755
rect 1646 1759 1652 1760
rect 1646 1755 1647 1759
rect 1651 1755 1652 1759
rect 1646 1754 1652 1755
rect 1702 1759 1708 1760
rect 1702 1755 1703 1759
rect 1707 1755 1708 1759
rect 1702 1754 1708 1755
rect 1758 1759 1764 1760
rect 1758 1755 1759 1759
rect 1763 1755 1764 1759
rect 1758 1754 1764 1755
rect 1806 1759 1812 1760
rect 1806 1755 1807 1759
rect 1811 1755 1812 1759
rect 1806 1754 1812 1755
rect 1862 1759 1868 1760
rect 1862 1755 1863 1759
rect 1867 1755 1868 1759
rect 1862 1754 1868 1755
rect 1918 1759 1924 1760
rect 1918 1755 1919 1759
rect 1923 1755 1924 1759
rect 1918 1754 1924 1755
rect 1974 1759 1980 1760
rect 1974 1755 1975 1759
rect 1979 1755 1980 1759
rect 1974 1754 1980 1755
rect 2408 1737 2410 1769
rect 110 1736 116 1737
rect 110 1732 111 1736
rect 115 1732 116 1736
rect 110 1731 116 1732
rect 1238 1736 1244 1737
rect 1238 1732 1239 1736
rect 1243 1732 1244 1736
rect 1238 1731 1244 1732
rect 1278 1736 1284 1737
rect 1278 1732 1279 1736
rect 1283 1732 1284 1736
rect 1278 1731 1284 1732
rect 2406 1736 2412 1737
rect 2406 1732 2407 1736
rect 2411 1732 2412 1736
rect 2406 1731 2412 1732
rect 110 1719 116 1720
rect 110 1715 111 1719
rect 115 1715 116 1719
rect 110 1714 116 1715
rect 1238 1719 1244 1720
rect 1238 1715 1239 1719
rect 1243 1715 1244 1719
rect 1238 1714 1244 1715
rect 1278 1719 1284 1720
rect 1278 1715 1279 1719
rect 1283 1715 1284 1719
rect 1278 1714 1284 1715
rect 2406 1719 2412 1720
rect 2406 1715 2407 1719
rect 2411 1715 2412 1719
rect 2406 1714 2412 1715
rect 112 1703 114 1714
rect 406 1712 412 1713
rect 406 1708 407 1712
rect 411 1708 412 1712
rect 406 1707 412 1708
rect 446 1712 452 1713
rect 446 1708 447 1712
rect 451 1708 452 1712
rect 446 1707 452 1708
rect 486 1712 492 1713
rect 486 1708 487 1712
rect 491 1708 492 1712
rect 486 1707 492 1708
rect 526 1712 532 1713
rect 526 1708 527 1712
rect 531 1708 532 1712
rect 526 1707 532 1708
rect 566 1712 572 1713
rect 566 1708 567 1712
rect 571 1708 572 1712
rect 566 1707 572 1708
rect 606 1712 612 1713
rect 606 1708 607 1712
rect 611 1708 612 1712
rect 606 1707 612 1708
rect 646 1712 652 1713
rect 646 1708 647 1712
rect 651 1708 652 1712
rect 646 1707 652 1708
rect 694 1712 700 1713
rect 694 1708 695 1712
rect 699 1708 700 1712
rect 694 1707 700 1708
rect 750 1712 756 1713
rect 750 1708 751 1712
rect 755 1708 756 1712
rect 750 1707 756 1708
rect 806 1712 812 1713
rect 806 1708 807 1712
rect 811 1708 812 1712
rect 806 1707 812 1708
rect 870 1712 876 1713
rect 870 1708 871 1712
rect 875 1708 876 1712
rect 870 1707 876 1708
rect 934 1712 940 1713
rect 934 1708 935 1712
rect 939 1708 940 1712
rect 934 1707 940 1708
rect 998 1712 1004 1713
rect 998 1708 999 1712
rect 1003 1708 1004 1712
rect 998 1707 1004 1708
rect 1070 1712 1076 1713
rect 1070 1708 1071 1712
rect 1075 1708 1076 1712
rect 1070 1707 1076 1708
rect 1142 1712 1148 1713
rect 1142 1708 1143 1712
rect 1147 1708 1148 1712
rect 1142 1707 1148 1708
rect 1190 1712 1196 1713
rect 1190 1708 1191 1712
rect 1195 1708 1196 1712
rect 1190 1707 1196 1708
rect 408 1703 410 1707
rect 448 1703 450 1707
rect 488 1703 490 1707
rect 528 1703 530 1707
rect 568 1703 570 1707
rect 608 1703 610 1707
rect 648 1703 650 1707
rect 696 1703 698 1707
rect 752 1703 754 1707
rect 808 1703 810 1707
rect 872 1703 874 1707
rect 936 1703 938 1707
rect 1000 1703 1002 1707
rect 1072 1703 1074 1707
rect 1144 1703 1146 1707
rect 1192 1703 1194 1707
rect 1240 1703 1242 1714
rect 1280 1703 1282 1714
rect 1302 1712 1308 1713
rect 1302 1708 1303 1712
rect 1307 1708 1308 1712
rect 1302 1707 1308 1708
rect 1342 1712 1348 1713
rect 1342 1708 1343 1712
rect 1347 1708 1348 1712
rect 1342 1707 1348 1708
rect 1390 1712 1396 1713
rect 1390 1708 1391 1712
rect 1395 1708 1396 1712
rect 1390 1707 1396 1708
rect 1454 1712 1460 1713
rect 1454 1708 1455 1712
rect 1459 1708 1460 1712
rect 1454 1707 1460 1708
rect 1518 1712 1524 1713
rect 1518 1708 1519 1712
rect 1523 1708 1524 1712
rect 1518 1707 1524 1708
rect 1582 1712 1588 1713
rect 1582 1708 1583 1712
rect 1587 1708 1588 1712
rect 1582 1707 1588 1708
rect 1646 1712 1652 1713
rect 1646 1708 1647 1712
rect 1651 1708 1652 1712
rect 1646 1707 1652 1708
rect 1702 1712 1708 1713
rect 1702 1708 1703 1712
rect 1707 1708 1708 1712
rect 1702 1707 1708 1708
rect 1758 1712 1764 1713
rect 1758 1708 1759 1712
rect 1763 1708 1764 1712
rect 1758 1707 1764 1708
rect 1806 1712 1812 1713
rect 1806 1708 1807 1712
rect 1811 1708 1812 1712
rect 1806 1707 1812 1708
rect 1862 1712 1868 1713
rect 1862 1708 1863 1712
rect 1867 1708 1868 1712
rect 1862 1707 1868 1708
rect 1918 1712 1924 1713
rect 1918 1708 1919 1712
rect 1923 1708 1924 1712
rect 1918 1707 1924 1708
rect 1974 1712 1980 1713
rect 1974 1708 1975 1712
rect 1979 1708 1980 1712
rect 1974 1707 1980 1708
rect 1304 1703 1306 1707
rect 1344 1703 1346 1707
rect 1392 1703 1394 1707
rect 1456 1703 1458 1707
rect 1520 1703 1522 1707
rect 1584 1703 1586 1707
rect 1648 1703 1650 1707
rect 1704 1703 1706 1707
rect 1760 1703 1762 1707
rect 1808 1703 1810 1707
rect 1864 1703 1866 1707
rect 1920 1703 1922 1707
rect 1976 1703 1978 1707
rect 2408 1703 2410 1714
rect 111 1702 115 1703
rect 111 1697 115 1698
rect 279 1702 283 1703
rect 279 1697 283 1698
rect 319 1702 323 1703
rect 319 1697 323 1698
rect 359 1702 363 1703
rect 359 1697 363 1698
rect 399 1702 403 1703
rect 399 1697 403 1698
rect 407 1702 411 1703
rect 407 1697 411 1698
rect 447 1702 451 1703
rect 447 1697 451 1698
rect 487 1702 491 1703
rect 487 1697 491 1698
rect 495 1702 499 1703
rect 495 1697 499 1698
rect 527 1702 531 1703
rect 527 1697 531 1698
rect 543 1702 547 1703
rect 543 1697 547 1698
rect 567 1702 571 1703
rect 567 1697 571 1698
rect 591 1702 595 1703
rect 591 1697 595 1698
rect 607 1702 611 1703
rect 607 1697 611 1698
rect 639 1702 643 1703
rect 639 1697 643 1698
rect 647 1702 651 1703
rect 647 1697 651 1698
rect 687 1702 691 1703
rect 687 1697 691 1698
rect 695 1702 699 1703
rect 695 1697 699 1698
rect 735 1702 739 1703
rect 735 1697 739 1698
rect 751 1702 755 1703
rect 751 1697 755 1698
rect 783 1702 787 1703
rect 783 1697 787 1698
rect 807 1702 811 1703
rect 807 1697 811 1698
rect 839 1702 843 1703
rect 839 1697 843 1698
rect 871 1702 875 1703
rect 871 1697 875 1698
rect 895 1702 899 1703
rect 895 1697 899 1698
rect 935 1702 939 1703
rect 935 1697 939 1698
rect 999 1702 1003 1703
rect 999 1697 1003 1698
rect 1071 1702 1075 1703
rect 1071 1697 1075 1698
rect 1143 1702 1147 1703
rect 1143 1697 1147 1698
rect 1191 1702 1195 1703
rect 1191 1697 1195 1698
rect 1239 1702 1243 1703
rect 1239 1697 1243 1698
rect 1279 1702 1283 1703
rect 1279 1697 1283 1698
rect 1303 1702 1307 1703
rect 1303 1697 1307 1698
rect 1343 1702 1347 1703
rect 1343 1697 1347 1698
rect 1383 1702 1387 1703
rect 1383 1697 1387 1698
rect 1391 1702 1395 1703
rect 1391 1697 1395 1698
rect 1423 1702 1427 1703
rect 1423 1697 1427 1698
rect 1455 1702 1459 1703
rect 1455 1697 1459 1698
rect 1463 1702 1467 1703
rect 1463 1697 1467 1698
rect 1503 1702 1507 1703
rect 1503 1697 1507 1698
rect 1519 1702 1523 1703
rect 1519 1697 1523 1698
rect 1559 1702 1563 1703
rect 1559 1697 1563 1698
rect 1583 1702 1587 1703
rect 1583 1697 1587 1698
rect 1623 1702 1627 1703
rect 1623 1697 1627 1698
rect 1647 1702 1651 1703
rect 1647 1697 1651 1698
rect 1687 1702 1691 1703
rect 1687 1697 1691 1698
rect 1703 1702 1707 1703
rect 1703 1697 1707 1698
rect 1751 1702 1755 1703
rect 1751 1697 1755 1698
rect 1759 1702 1763 1703
rect 1759 1697 1763 1698
rect 1807 1702 1811 1703
rect 1807 1697 1811 1698
rect 1863 1702 1867 1703
rect 1863 1697 1867 1698
rect 1919 1702 1923 1703
rect 1919 1697 1923 1698
rect 1975 1702 1979 1703
rect 1975 1697 1979 1698
rect 2031 1702 2035 1703
rect 2031 1697 2035 1698
rect 2087 1702 2091 1703
rect 2087 1697 2091 1698
rect 2407 1702 2411 1703
rect 2407 1697 2411 1698
rect 112 1690 114 1697
rect 278 1696 284 1697
rect 278 1692 279 1696
rect 283 1692 284 1696
rect 278 1691 284 1692
rect 318 1696 324 1697
rect 318 1692 319 1696
rect 323 1692 324 1696
rect 318 1691 324 1692
rect 358 1696 364 1697
rect 358 1692 359 1696
rect 363 1692 364 1696
rect 358 1691 364 1692
rect 398 1696 404 1697
rect 398 1692 399 1696
rect 403 1692 404 1696
rect 398 1691 404 1692
rect 446 1696 452 1697
rect 446 1692 447 1696
rect 451 1692 452 1696
rect 446 1691 452 1692
rect 494 1696 500 1697
rect 494 1692 495 1696
rect 499 1692 500 1696
rect 494 1691 500 1692
rect 542 1696 548 1697
rect 542 1692 543 1696
rect 547 1692 548 1696
rect 542 1691 548 1692
rect 590 1696 596 1697
rect 590 1692 591 1696
rect 595 1692 596 1696
rect 590 1691 596 1692
rect 638 1696 644 1697
rect 638 1692 639 1696
rect 643 1692 644 1696
rect 638 1691 644 1692
rect 686 1696 692 1697
rect 686 1692 687 1696
rect 691 1692 692 1696
rect 686 1691 692 1692
rect 734 1696 740 1697
rect 734 1692 735 1696
rect 739 1692 740 1696
rect 734 1691 740 1692
rect 782 1696 788 1697
rect 782 1692 783 1696
rect 787 1692 788 1696
rect 782 1691 788 1692
rect 838 1696 844 1697
rect 838 1692 839 1696
rect 843 1692 844 1696
rect 838 1691 844 1692
rect 894 1696 900 1697
rect 894 1692 895 1696
rect 899 1692 900 1696
rect 894 1691 900 1692
rect 1240 1690 1242 1697
rect 1280 1690 1282 1697
rect 1302 1696 1308 1697
rect 1302 1692 1303 1696
rect 1307 1692 1308 1696
rect 1302 1691 1308 1692
rect 1342 1696 1348 1697
rect 1342 1692 1343 1696
rect 1347 1692 1348 1696
rect 1342 1691 1348 1692
rect 1382 1696 1388 1697
rect 1382 1692 1383 1696
rect 1387 1692 1388 1696
rect 1382 1691 1388 1692
rect 1422 1696 1428 1697
rect 1422 1692 1423 1696
rect 1427 1692 1428 1696
rect 1422 1691 1428 1692
rect 1462 1696 1468 1697
rect 1462 1692 1463 1696
rect 1467 1692 1468 1696
rect 1462 1691 1468 1692
rect 1502 1696 1508 1697
rect 1502 1692 1503 1696
rect 1507 1692 1508 1696
rect 1502 1691 1508 1692
rect 1558 1696 1564 1697
rect 1558 1692 1559 1696
rect 1563 1692 1564 1696
rect 1558 1691 1564 1692
rect 1622 1696 1628 1697
rect 1622 1692 1623 1696
rect 1627 1692 1628 1696
rect 1622 1691 1628 1692
rect 1686 1696 1692 1697
rect 1686 1692 1687 1696
rect 1691 1692 1692 1696
rect 1686 1691 1692 1692
rect 1750 1696 1756 1697
rect 1750 1692 1751 1696
rect 1755 1692 1756 1696
rect 1750 1691 1756 1692
rect 1806 1696 1812 1697
rect 1806 1692 1807 1696
rect 1811 1692 1812 1696
rect 1806 1691 1812 1692
rect 1862 1696 1868 1697
rect 1862 1692 1863 1696
rect 1867 1692 1868 1696
rect 1862 1691 1868 1692
rect 1918 1696 1924 1697
rect 1918 1692 1919 1696
rect 1923 1692 1924 1696
rect 1918 1691 1924 1692
rect 1974 1696 1980 1697
rect 1974 1692 1975 1696
rect 1979 1692 1980 1696
rect 1974 1691 1980 1692
rect 2030 1696 2036 1697
rect 2030 1692 2031 1696
rect 2035 1692 2036 1696
rect 2030 1691 2036 1692
rect 2086 1696 2092 1697
rect 2086 1692 2087 1696
rect 2091 1692 2092 1696
rect 2086 1691 2092 1692
rect 2408 1690 2410 1697
rect 110 1689 116 1690
rect 110 1685 111 1689
rect 115 1685 116 1689
rect 110 1684 116 1685
rect 1238 1689 1244 1690
rect 1238 1685 1239 1689
rect 1243 1685 1244 1689
rect 1238 1684 1244 1685
rect 1278 1689 1284 1690
rect 1278 1685 1279 1689
rect 1283 1685 1284 1689
rect 1278 1684 1284 1685
rect 2406 1689 2412 1690
rect 2406 1685 2407 1689
rect 2411 1685 2412 1689
rect 2406 1684 2412 1685
rect 110 1672 116 1673
rect 110 1668 111 1672
rect 115 1668 116 1672
rect 110 1667 116 1668
rect 1238 1672 1244 1673
rect 1238 1668 1239 1672
rect 1243 1668 1244 1672
rect 1238 1667 1244 1668
rect 1278 1672 1284 1673
rect 1278 1668 1279 1672
rect 1283 1668 1284 1672
rect 1278 1667 1284 1668
rect 2406 1672 2412 1673
rect 2406 1668 2407 1672
rect 2411 1668 2412 1672
rect 2406 1667 2412 1668
rect 112 1631 114 1667
rect 278 1649 284 1650
rect 278 1645 279 1649
rect 283 1645 284 1649
rect 278 1644 284 1645
rect 318 1649 324 1650
rect 318 1645 319 1649
rect 323 1645 324 1649
rect 318 1644 324 1645
rect 358 1649 364 1650
rect 358 1645 359 1649
rect 363 1645 364 1649
rect 358 1644 364 1645
rect 398 1649 404 1650
rect 398 1645 399 1649
rect 403 1645 404 1649
rect 398 1644 404 1645
rect 446 1649 452 1650
rect 446 1645 447 1649
rect 451 1645 452 1649
rect 446 1644 452 1645
rect 494 1649 500 1650
rect 494 1645 495 1649
rect 499 1645 500 1649
rect 494 1644 500 1645
rect 542 1649 548 1650
rect 542 1645 543 1649
rect 547 1645 548 1649
rect 542 1644 548 1645
rect 590 1649 596 1650
rect 590 1645 591 1649
rect 595 1645 596 1649
rect 590 1644 596 1645
rect 638 1649 644 1650
rect 638 1645 639 1649
rect 643 1645 644 1649
rect 638 1644 644 1645
rect 686 1649 692 1650
rect 686 1645 687 1649
rect 691 1645 692 1649
rect 686 1644 692 1645
rect 734 1649 740 1650
rect 734 1645 735 1649
rect 739 1645 740 1649
rect 734 1644 740 1645
rect 782 1649 788 1650
rect 782 1645 783 1649
rect 787 1645 788 1649
rect 782 1644 788 1645
rect 838 1649 844 1650
rect 838 1645 839 1649
rect 843 1645 844 1649
rect 838 1644 844 1645
rect 894 1649 900 1650
rect 894 1645 895 1649
rect 899 1645 900 1649
rect 894 1644 900 1645
rect 280 1631 282 1644
rect 320 1631 322 1644
rect 360 1631 362 1644
rect 400 1631 402 1644
rect 448 1631 450 1644
rect 496 1631 498 1644
rect 544 1631 546 1644
rect 592 1631 594 1644
rect 640 1631 642 1644
rect 688 1631 690 1644
rect 736 1631 738 1644
rect 784 1631 786 1644
rect 840 1631 842 1644
rect 896 1631 898 1644
rect 1240 1631 1242 1667
rect 1280 1631 1282 1667
rect 1302 1649 1308 1650
rect 1302 1645 1303 1649
rect 1307 1645 1308 1649
rect 1302 1644 1308 1645
rect 1342 1649 1348 1650
rect 1342 1645 1343 1649
rect 1347 1645 1348 1649
rect 1342 1644 1348 1645
rect 1382 1649 1388 1650
rect 1382 1645 1383 1649
rect 1387 1645 1388 1649
rect 1382 1644 1388 1645
rect 1422 1649 1428 1650
rect 1422 1645 1423 1649
rect 1427 1645 1428 1649
rect 1422 1644 1428 1645
rect 1462 1649 1468 1650
rect 1462 1645 1463 1649
rect 1467 1645 1468 1649
rect 1462 1644 1468 1645
rect 1502 1649 1508 1650
rect 1502 1645 1503 1649
rect 1507 1645 1508 1649
rect 1502 1644 1508 1645
rect 1558 1649 1564 1650
rect 1558 1645 1559 1649
rect 1563 1645 1564 1649
rect 1558 1644 1564 1645
rect 1622 1649 1628 1650
rect 1622 1645 1623 1649
rect 1627 1645 1628 1649
rect 1622 1644 1628 1645
rect 1686 1649 1692 1650
rect 1686 1645 1687 1649
rect 1691 1645 1692 1649
rect 1686 1644 1692 1645
rect 1750 1649 1756 1650
rect 1750 1645 1751 1649
rect 1755 1645 1756 1649
rect 1750 1644 1756 1645
rect 1806 1649 1812 1650
rect 1806 1645 1807 1649
rect 1811 1645 1812 1649
rect 1806 1644 1812 1645
rect 1862 1649 1868 1650
rect 1862 1645 1863 1649
rect 1867 1645 1868 1649
rect 1862 1644 1868 1645
rect 1918 1649 1924 1650
rect 1918 1645 1919 1649
rect 1923 1645 1924 1649
rect 1918 1644 1924 1645
rect 1974 1649 1980 1650
rect 1974 1645 1975 1649
rect 1979 1645 1980 1649
rect 1974 1644 1980 1645
rect 2030 1649 2036 1650
rect 2030 1645 2031 1649
rect 2035 1645 2036 1649
rect 2030 1644 2036 1645
rect 2086 1649 2092 1650
rect 2086 1645 2087 1649
rect 2091 1645 2092 1649
rect 2086 1644 2092 1645
rect 1304 1631 1306 1644
rect 1344 1631 1346 1644
rect 1384 1631 1386 1644
rect 1424 1631 1426 1644
rect 1464 1631 1466 1644
rect 1504 1631 1506 1644
rect 1560 1631 1562 1644
rect 1624 1631 1626 1644
rect 1688 1631 1690 1644
rect 1752 1631 1754 1644
rect 1808 1631 1810 1644
rect 1864 1631 1866 1644
rect 1920 1631 1922 1644
rect 1976 1631 1978 1644
rect 2032 1631 2034 1644
rect 2088 1631 2090 1644
rect 2408 1631 2410 1667
rect 111 1630 115 1631
rect 111 1625 115 1626
rect 135 1630 139 1631
rect 135 1625 139 1626
rect 175 1630 179 1631
rect 175 1625 179 1626
rect 215 1630 219 1631
rect 215 1625 219 1626
rect 255 1630 259 1631
rect 255 1625 259 1626
rect 279 1630 283 1631
rect 279 1625 283 1626
rect 311 1630 315 1631
rect 311 1625 315 1626
rect 319 1630 323 1631
rect 319 1625 323 1626
rect 359 1630 363 1631
rect 359 1625 363 1626
rect 391 1630 395 1631
rect 391 1625 395 1626
rect 399 1630 403 1631
rect 399 1625 403 1626
rect 447 1630 451 1631
rect 447 1625 451 1626
rect 471 1630 475 1631
rect 471 1625 475 1626
rect 495 1630 499 1631
rect 495 1625 499 1626
rect 543 1630 547 1631
rect 543 1625 547 1626
rect 559 1630 563 1631
rect 559 1625 563 1626
rect 591 1630 595 1631
rect 591 1625 595 1626
rect 639 1630 643 1631
rect 639 1625 643 1626
rect 687 1630 691 1631
rect 687 1625 691 1626
rect 719 1630 723 1631
rect 719 1625 723 1626
rect 735 1630 739 1631
rect 735 1625 739 1626
rect 783 1630 787 1631
rect 783 1625 787 1626
rect 791 1630 795 1631
rect 791 1625 795 1626
rect 839 1630 843 1631
rect 839 1625 843 1626
rect 855 1630 859 1631
rect 855 1625 859 1626
rect 895 1630 899 1631
rect 895 1625 899 1626
rect 919 1630 923 1631
rect 919 1625 923 1626
rect 983 1630 987 1631
rect 983 1625 987 1626
rect 1047 1630 1051 1631
rect 1047 1625 1051 1626
rect 1239 1630 1243 1631
rect 1239 1625 1243 1626
rect 1279 1630 1283 1631
rect 1279 1625 1283 1626
rect 1303 1630 1307 1631
rect 1303 1625 1307 1626
rect 1343 1630 1347 1631
rect 1343 1625 1347 1626
rect 1383 1630 1387 1631
rect 1383 1625 1387 1626
rect 1423 1630 1427 1631
rect 1423 1625 1427 1626
rect 1463 1630 1467 1631
rect 1463 1625 1467 1626
rect 1503 1630 1507 1631
rect 1503 1625 1507 1626
rect 1559 1630 1563 1631
rect 1559 1625 1563 1626
rect 1623 1630 1627 1631
rect 1623 1625 1627 1626
rect 1631 1630 1635 1631
rect 1631 1625 1635 1626
rect 1687 1630 1691 1631
rect 1687 1625 1691 1626
rect 1703 1630 1707 1631
rect 1703 1625 1707 1626
rect 1751 1630 1755 1631
rect 1751 1625 1755 1626
rect 1783 1630 1787 1631
rect 1783 1625 1787 1626
rect 1807 1630 1811 1631
rect 1807 1625 1811 1626
rect 1855 1630 1859 1631
rect 1855 1625 1859 1626
rect 1863 1630 1867 1631
rect 1863 1625 1867 1626
rect 1919 1630 1923 1631
rect 1919 1625 1923 1626
rect 1927 1630 1931 1631
rect 1927 1625 1931 1626
rect 1975 1630 1979 1631
rect 1975 1625 1979 1626
rect 1999 1630 2003 1631
rect 1999 1625 2003 1626
rect 2031 1630 2035 1631
rect 2031 1625 2035 1626
rect 2063 1630 2067 1631
rect 2063 1625 2067 1626
rect 2087 1630 2091 1631
rect 2087 1625 2091 1626
rect 2127 1630 2131 1631
rect 2127 1625 2131 1626
rect 2191 1630 2195 1631
rect 2191 1625 2195 1626
rect 2255 1630 2259 1631
rect 2255 1625 2259 1626
rect 2319 1630 2323 1631
rect 2319 1625 2323 1626
rect 2359 1630 2363 1631
rect 2359 1625 2363 1626
rect 2407 1630 2411 1631
rect 2407 1625 2411 1626
rect 112 1593 114 1625
rect 136 1616 138 1625
rect 176 1616 178 1625
rect 216 1616 218 1625
rect 256 1616 258 1625
rect 312 1616 314 1625
rect 392 1616 394 1625
rect 472 1616 474 1625
rect 560 1616 562 1625
rect 640 1616 642 1625
rect 720 1616 722 1625
rect 792 1616 794 1625
rect 856 1616 858 1625
rect 920 1616 922 1625
rect 984 1616 986 1625
rect 1048 1616 1050 1625
rect 134 1615 140 1616
rect 134 1611 135 1615
rect 139 1611 140 1615
rect 134 1610 140 1611
rect 174 1615 180 1616
rect 174 1611 175 1615
rect 179 1611 180 1615
rect 174 1610 180 1611
rect 214 1615 220 1616
rect 214 1611 215 1615
rect 219 1611 220 1615
rect 214 1610 220 1611
rect 254 1615 260 1616
rect 254 1611 255 1615
rect 259 1611 260 1615
rect 254 1610 260 1611
rect 310 1615 316 1616
rect 310 1611 311 1615
rect 315 1611 316 1615
rect 310 1610 316 1611
rect 390 1615 396 1616
rect 390 1611 391 1615
rect 395 1611 396 1615
rect 390 1610 396 1611
rect 470 1615 476 1616
rect 470 1611 471 1615
rect 475 1611 476 1615
rect 470 1610 476 1611
rect 558 1615 564 1616
rect 558 1611 559 1615
rect 563 1611 564 1615
rect 558 1610 564 1611
rect 638 1615 644 1616
rect 638 1611 639 1615
rect 643 1611 644 1615
rect 638 1610 644 1611
rect 718 1615 724 1616
rect 718 1611 719 1615
rect 723 1611 724 1615
rect 718 1610 724 1611
rect 790 1615 796 1616
rect 790 1611 791 1615
rect 795 1611 796 1615
rect 790 1610 796 1611
rect 854 1615 860 1616
rect 854 1611 855 1615
rect 859 1611 860 1615
rect 854 1610 860 1611
rect 918 1615 924 1616
rect 918 1611 919 1615
rect 923 1611 924 1615
rect 918 1610 924 1611
rect 982 1615 988 1616
rect 982 1611 983 1615
rect 987 1611 988 1615
rect 982 1610 988 1611
rect 1046 1615 1052 1616
rect 1046 1611 1047 1615
rect 1051 1611 1052 1615
rect 1046 1610 1052 1611
rect 1240 1593 1242 1625
rect 1280 1593 1282 1625
rect 1304 1616 1306 1625
rect 1344 1616 1346 1625
rect 1384 1616 1386 1625
rect 1424 1616 1426 1625
rect 1464 1616 1466 1625
rect 1504 1616 1506 1625
rect 1560 1616 1562 1625
rect 1632 1616 1634 1625
rect 1704 1616 1706 1625
rect 1784 1616 1786 1625
rect 1856 1616 1858 1625
rect 1928 1616 1930 1625
rect 2000 1616 2002 1625
rect 2064 1616 2066 1625
rect 2128 1616 2130 1625
rect 2192 1616 2194 1625
rect 2256 1616 2258 1625
rect 2320 1616 2322 1625
rect 2360 1616 2362 1625
rect 1302 1615 1308 1616
rect 1302 1611 1303 1615
rect 1307 1611 1308 1615
rect 1302 1610 1308 1611
rect 1342 1615 1348 1616
rect 1342 1611 1343 1615
rect 1347 1611 1348 1615
rect 1342 1610 1348 1611
rect 1382 1615 1388 1616
rect 1382 1611 1383 1615
rect 1387 1611 1388 1615
rect 1382 1610 1388 1611
rect 1422 1615 1428 1616
rect 1422 1611 1423 1615
rect 1427 1611 1428 1615
rect 1422 1610 1428 1611
rect 1462 1615 1468 1616
rect 1462 1611 1463 1615
rect 1467 1611 1468 1615
rect 1462 1610 1468 1611
rect 1502 1615 1508 1616
rect 1502 1611 1503 1615
rect 1507 1611 1508 1615
rect 1502 1610 1508 1611
rect 1558 1615 1564 1616
rect 1558 1611 1559 1615
rect 1563 1611 1564 1615
rect 1558 1610 1564 1611
rect 1630 1615 1636 1616
rect 1630 1611 1631 1615
rect 1635 1611 1636 1615
rect 1630 1610 1636 1611
rect 1702 1615 1708 1616
rect 1702 1611 1703 1615
rect 1707 1611 1708 1615
rect 1702 1610 1708 1611
rect 1782 1615 1788 1616
rect 1782 1611 1783 1615
rect 1787 1611 1788 1615
rect 1782 1610 1788 1611
rect 1854 1615 1860 1616
rect 1854 1611 1855 1615
rect 1859 1611 1860 1615
rect 1854 1610 1860 1611
rect 1926 1615 1932 1616
rect 1926 1611 1927 1615
rect 1931 1611 1932 1615
rect 1926 1610 1932 1611
rect 1998 1615 2004 1616
rect 1998 1611 1999 1615
rect 2003 1611 2004 1615
rect 1998 1610 2004 1611
rect 2062 1615 2068 1616
rect 2062 1611 2063 1615
rect 2067 1611 2068 1615
rect 2062 1610 2068 1611
rect 2126 1615 2132 1616
rect 2126 1611 2127 1615
rect 2131 1611 2132 1615
rect 2126 1610 2132 1611
rect 2190 1615 2196 1616
rect 2190 1611 2191 1615
rect 2195 1611 2196 1615
rect 2190 1610 2196 1611
rect 2254 1615 2260 1616
rect 2254 1611 2255 1615
rect 2259 1611 2260 1615
rect 2254 1610 2260 1611
rect 2318 1615 2324 1616
rect 2318 1611 2319 1615
rect 2323 1611 2324 1615
rect 2318 1610 2324 1611
rect 2358 1615 2364 1616
rect 2358 1611 2359 1615
rect 2363 1611 2364 1615
rect 2358 1610 2364 1611
rect 2408 1593 2410 1625
rect 110 1592 116 1593
rect 110 1588 111 1592
rect 115 1588 116 1592
rect 110 1587 116 1588
rect 1238 1592 1244 1593
rect 1238 1588 1239 1592
rect 1243 1588 1244 1592
rect 1238 1587 1244 1588
rect 1278 1592 1284 1593
rect 1278 1588 1279 1592
rect 1283 1588 1284 1592
rect 1278 1587 1284 1588
rect 2406 1592 2412 1593
rect 2406 1588 2407 1592
rect 2411 1588 2412 1592
rect 2406 1587 2412 1588
rect 110 1575 116 1576
rect 110 1571 111 1575
rect 115 1571 116 1575
rect 110 1570 116 1571
rect 1238 1575 1244 1576
rect 1238 1571 1239 1575
rect 1243 1571 1244 1575
rect 1238 1570 1244 1571
rect 1278 1575 1284 1576
rect 1278 1571 1279 1575
rect 1283 1571 1284 1575
rect 1278 1570 1284 1571
rect 2406 1575 2412 1576
rect 2406 1571 2407 1575
rect 2411 1571 2412 1575
rect 2406 1570 2412 1571
rect 112 1559 114 1570
rect 134 1568 140 1569
rect 134 1564 135 1568
rect 139 1564 140 1568
rect 134 1563 140 1564
rect 174 1568 180 1569
rect 174 1564 175 1568
rect 179 1564 180 1568
rect 174 1563 180 1564
rect 214 1568 220 1569
rect 214 1564 215 1568
rect 219 1564 220 1568
rect 214 1563 220 1564
rect 254 1568 260 1569
rect 254 1564 255 1568
rect 259 1564 260 1568
rect 254 1563 260 1564
rect 310 1568 316 1569
rect 310 1564 311 1568
rect 315 1564 316 1568
rect 310 1563 316 1564
rect 390 1568 396 1569
rect 390 1564 391 1568
rect 395 1564 396 1568
rect 390 1563 396 1564
rect 470 1568 476 1569
rect 470 1564 471 1568
rect 475 1564 476 1568
rect 470 1563 476 1564
rect 558 1568 564 1569
rect 558 1564 559 1568
rect 563 1564 564 1568
rect 558 1563 564 1564
rect 638 1568 644 1569
rect 638 1564 639 1568
rect 643 1564 644 1568
rect 638 1563 644 1564
rect 718 1568 724 1569
rect 718 1564 719 1568
rect 723 1564 724 1568
rect 718 1563 724 1564
rect 790 1568 796 1569
rect 790 1564 791 1568
rect 795 1564 796 1568
rect 790 1563 796 1564
rect 854 1568 860 1569
rect 854 1564 855 1568
rect 859 1564 860 1568
rect 854 1563 860 1564
rect 918 1568 924 1569
rect 918 1564 919 1568
rect 923 1564 924 1568
rect 918 1563 924 1564
rect 982 1568 988 1569
rect 982 1564 983 1568
rect 987 1564 988 1568
rect 982 1563 988 1564
rect 1046 1568 1052 1569
rect 1046 1564 1047 1568
rect 1051 1564 1052 1568
rect 1046 1563 1052 1564
rect 136 1559 138 1563
rect 176 1559 178 1563
rect 216 1559 218 1563
rect 256 1559 258 1563
rect 312 1559 314 1563
rect 392 1559 394 1563
rect 472 1559 474 1563
rect 560 1559 562 1563
rect 640 1559 642 1563
rect 720 1559 722 1563
rect 792 1559 794 1563
rect 856 1559 858 1563
rect 920 1559 922 1563
rect 984 1559 986 1563
rect 1048 1559 1050 1563
rect 1240 1559 1242 1570
rect 1280 1563 1282 1570
rect 1302 1568 1308 1569
rect 1302 1564 1303 1568
rect 1307 1564 1308 1568
rect 1302 1563 1308 1564
rect 1342 1568 1348 1569
rect 1342 1564 1343 1568
rect 1347 1564 1348 1568
rect 1342 1563 1348 1564
rect 1382 1568 1388 1569
rect 1382 1564 1383 1568
rect 1387 1564 1388 1568
rect 1382 1563 1388 1564
rect 1422 1568 1428 1569
rect 1422 1564 1423 1568
rect 1427 1564 1428 1568
rect 1422 1563 1428 1564
rect 1462 1568 1468 1569
rect 1462 1564 1463 1568
rect 1467 1564 1468 1568
rect 1462 1563 1468 1564
rect 1502 1568 1508 1569
rect 1502 1564 1503 1568
rect 1507 1564 1508 1568
rect 1502 1563 1508 1564
rect 1558 1568 1564 1569
rect 1558 1564 1559 1568
rect 1563 1564 1564 1568
rect 1558 1563 1564 1564
rect 1630 1568 1636 1569
rect 1630 1564 1631 1568
rect 1635 1564 1636 1568
rect 1630 1563 1636 1564
rect 1702 1568 1708 1569
rect 1702 1564 1703 1568
rect 1707 1564 1708 1568
rect 1702 1563 1708 1564
rect 1782 1568 1788 1569
rect 1782 1564 1783 1568
rect 1787 1564 1788 1568
rect 1782 1563 1788 1564
rect 1854 1568 1860 1569
rect 1854 1564 1855 1568
rect 1859 1564 1860 1568
rect 1854 1563 1860 1564
rect 1926 1568 1932 1569
rect 1926 1564 1927 1568
rect 1931 1564 1932 1568
rect 1926 1563 1932 1564
rect 1998 1568 2004 1569
rect 1998 1564 1999 1568
rect 2003 1564 2004 1568
rect 1998 1563 2004 1564
rect 2062 1568 2068 1569
rect 2062 1564 2063 1568
rect 2067 1564 2068 1568
rect 2062 1563 2068 1564
rect 2126 1568 2132 1569
rect 2126 1564 2127 1568
rect 2131 1564 2132 1568
rect 2126 1563 2132 1564
rect 2190 1568 2196 1569
rect 2190 1564 2191 1568
rect 2195 1564 2196 1568
rect 2190 1563 2196 1564
rect 2254 1568 2260 1569
rect 2254 1564 2255 1568
rect 2259 1564 2260 1568
rect 2254 1563 2260 1564
rect 2318 1568 2324 1569
rect 2318 1564 2319 1568
rect 2323 1564 2324 1568
rect 2318 1563 2324 1564
rect 2358 1568 2364 1569
rect 2358 1564 2359 1568
rect 2363 1564 2364 1568
rect 2358 1563 2364 1564
rect 2408 1563 2410 1570
rect 1279 1562 1283 1563
rect 111 1558 115 1559
rect 111 1553 115 1554
rect 135 1558 139 1559
rect 135 1553 139 1554
rect 151 1558 155 1559
rect 151 1553 155 1554
rect 175 1558 179 1559
rect 175 1553 179 1554
rect 199 1558 203 1559
rect 199 1553 203 1554
rect 215 1558 219 1559
rect 215 1553 219 1554
rect 255 1558 259 1559
rect 255 1553 259 1554
rect 263 1558 267 1559
rect 263 1553 267 1554
rect 311 1558 315 1559
rect 311 1553 315 1554
rect 343 1558 347 1559
rect 343 1553 347 1554
rect 391 1558 395 1559
rect 391 1553 395 1554
rect 439 1558 443 1559
rect 439 1553 443 1554
rect 471 1558 475 1559
rect 471 1553 475 1554
rect 535 1558 539 1559
rect 535 1553 539 1554
rect 559 1558 563 1559
rect 559 1553 563 1554
rect 639 1558 643 1559
rect 639 1553 643 1554
rect 719 1558 723 1559
rect 719 1553 723 1554
rect 735 1558 739 1559
rect 735 1553 739 1554
rect 791 1558 795 1559
rect 791 1553 795 1554
rect 823 1558 827 1559
rect 823 1553 827 1554
rect 855 1558 859 1559
rect 855 1553 859 1554
rect 903 1558 907 1559
rect 903 1553 907 1554
rect 919 1558 923 1559
rect 919 1553 923 1554
rect 975 1558 979 1559
rect 975 1553 979 1554
rect 983 1558 987 1559
rect 983 1553 987 1554
rect 1047 1558 1051 1559
rect 1047 1553 1051 1554
rect 1119 1558 1123 1559
rect 1119 1553 1123 1554
rect 1191 1558 1195 1559
rect 1191 1553 1195 1554
rect 1239 1558 1243 1559
rect 1279 1557 1283 1558
rect 1303 1562 1307 1563
rect 1303 1557 1307 1558
rect 1343 1562 1347 1563
rect 1343 1557 1347 1558
rect 1383 1562 1387 1563
rect 1383 1557 1387 1558
rect 1423 1562 1427 1563
rect 1423 1557 1427 1558
rect 1463 1562 1467 1563
rect 1463 1557 1467 1558
rect 1471 1562 1475 1563
rect 1471 1557 1475 1558
rect 1503 1562 1507 1563
rect 1503 1557 1507 1558
rect 1559 1562 1563 1563
rect 1559 1557 1563 1558
rect 1623 1562 1627 1563
rect 1623 1557 1627 1558
rect 1631 1562 1635 1563
rect 1631 1557 1635 1558
rect 1703 1562 1707 1563
rect 1703 1557 1707 1558
rect 1759 1562 1763 1563
rect 1759 1557 1763 1558
rect 1783 1562 1787 1563
rect 1783 1557 1787 1558
rect 1855 1562 1859 1563
rect 1855 1557 1859 1558
rect 1871 1562 1875 1563
rect 1871 1557 1875 1558
rect 1927 1562 1931 1563
rect 1927 1557 1931 1558
rect 1967 1562 1971 1563
rect 1967 1557 1971 1558
rect 1999 1562 2003 1563
rect 1999 1557 2003 1558
rect 2055 1562 2059 1563
rect 2055 1557 2059 1558
rect 2063 1562 2067 1563
rect 2063 1557 2067 1558
rect 2127 1562 2131 1563
rect 2127 1557 2131 1558
rect 2191 1562 2195 1563
rect 2191 1557 2195 1558
rect 2255 1562 2259 1563
rect 2255 1557 2259 1558
rect 2319 1562 2323 1563
rect 2319 1557 2323 1558
rect 2359 1562 2363 1563
rect 2359 1557 2363 1558
rect 2407 1562 2411 1563
rect 2407 1557 2411 1558
rect 1239 1553 1243 1554
rect 112 1546 114 1553
rect 150 1552 156 1553
rect 150 1548 151 1552
rect 155 1548 156 1552
rect 150 1547 156 1548
rect 198 1552 204 1553
rect 198 1548 199 1552
rect 203 1548 204 1552
rect 198 1547 204 1548
rect 262 1552 268 1553
rect 262 1548 263 1552
rect 267 1548 268 1552
rect 262 1547 268 1548
rect 342 1552 348 1553
rect 342 1548 343 1552
rect 347 1548 348 1552
rect 342 1547 348 1548
rect 438 1552 444 1553
rect 438 1548 439 1552
rect 443 1548 444 1552
rect 438 1547 444 1548
rect 534 1552 540 1553
rect 534 1548 535 1552
rect 539 1548 540 1552
rect 534 1547 540 1548
rect 638 1552 644 1553
rect 638 1548 639 1552
rect 643 1548 644 1552
rect 638 1547 644 1548
rect 734 1552 740 1553
rect 734 1548 735 1552
rect 739 1548 740 1552
rect 734 1547 740 1548
rect 822 1552 828 1553
rect 822 1548 823 1552
rect 827 1548 828 1552
rect 822 1547 828 1548
rect 902 1552 908 1553
rect 902 1548 903 1552
rect 907 1548 908 1552
rect 902 1547 908 1548
rect 974 1552 980 1553
rect 974 1548 975 1552
rect 979 1548 980 1552
rect 974 1547 980 1548
rect 1046 1552 1052 1553
rect 1046 1548 1047 1552
rect 1051 1548 1052 1552
rect 1046 1547 1052 1548
rect 1118 1552 1124 1553
rect 1118 1548 1119 1552
rect 1123 1548 1124 1552
rect 1118 1547 1124 1548
rect 1190 1552 1196 1553
rect 1190 1548 1191 1552
rect 1195 1548 1196 1552
rect 1190 1547 1196 1548
rect 1240 1546 1242 1553
rect 1280 1550 1282 1557
rect 1470 1556 1476 1557
rect 1470 1552 1471 1556
rect 1475 1552 1476 1556
rect 1470 1551 1476 1552
rect 1622 1556 1628 1557
rect 1622 1552 1623 1556
rect 1627 1552 1628 1556
rect 1622 1551 1628 1552
rect 1758 1556 1764 1557
rect 1758 1552 1759 1556
rect 1763 1552 1764 1556
rect 1758 1551 1764 1552
rect 1870 1556 1876 1557
rect 1870 1552 1871 1556
rect 1875 1552 1876 1556
rect 1870 1551 1876 1552
rect 1966 1556 1972 1557
rect 1966 1552 1967 1556
rect 1971 1552 1972 1556
rect 1966 1551 1972 1552
rect 2054 1556 2060 1557
rect 2054 1552 2055 1556
rect 2059 1552 2060 1556
rect 2054 1551 2060 1552
rect 2126 1556 2132 1557
rect 2126 1552 2127 1556
rect 2131 1552 2132 1556
rect 2126 1551 2132 1552
rect 2190 1556 2196 1557
rect 2190 1552 2191 1556
rect 2195 1552 2196 1556
rect 2190 1551 2196 1552
rect 2254 1556 2260 1557
rect 2254 1552 2255 1556
rect 2259 1552 2260 1556
rect 2254 1551 2260 1552
rect 2318 1556 2324 1557
rect 2318 1552 2319 1556
rect 2323 1552 2324 1556
rect 2318 1551 2324 1552
rect 2358 1556 2364 1557
rect 2358 1552 2359 1556
rect 2363 1552 2364 1556
rect 2358 1551 2364 1552
rect 2408 1550 2410 1557
rect 1278 1549 1284 1550
rect 110 1545 116 1546
rect 110 1541 111 1545
rect 115 1541 116 1545
rect 110 1540 116 1541
rect 1238 1545 1244 1546
rect 1238 1541 1239 1545
rect 1243 1541 1244 1545
rect 1278 1545 1279 1549
rect 1283 1545 1284 1549
rect 1278 1544 1284 1545
rect 2406 1549 2412 1550
rect 2406 1545 2407 1549
rect 2411 1545 2412 1549
rect 2406 1544 2412 1545
rect 1238 1540 1244 1541
rect 1278 1532 1284 1533
rect 110 1528 116 1529
rect 110 1524 111 1528
rect 115 1524 116 1528
rect 110 1523 116 1524
rect 1238 1528 1244 1529
rect 1238 1524 1239 1528
rect 1243 1524 1244 1528
rect 1278 1528 1279 1532
rect 1283 1528 1284 1532
rect 1278 1527 1284 1528
rect 2406 1532 2412 1533
rect 2406 1528 2407 1532
rect 2411 1528 2412 1532
rect 2406 1527 2412 1528
rect 1238 1523 1244 1524
rect 112 1487 114 1523
rect 150 1505 156 1506
rect 150 1501 151 1505
rect 155 1501 156 1505
rect 150 1500 156 1501
rect 198 1505 204 1506
rect 198 1501 199 1505
rect 203 1501 204 1505
rect 198 1500 204 1501
rect 262 1505 268 1506
rect 262 1501 263 1505
rect 267 1501 268 1505
rect 262 1500 268 1501
rect 342 1505 348 1506
rect 342 1501 343 1505
rect 347 1501 348 1505
rect 342 1500 348 1501
rect 438 1505 444 1506
rect 438 1501 439 1505
rect 443 1501 444 1505
rect 438 1500 444 1501
rect 534 1505 540 1506
rect 534 1501 535 1505
rect 539 1501 540 1505
rect 534 1500 540 1501
rect 638 1505 644 1506
rect 638 1501 639 1505
rect 643 1501 644 1505
rect 638 1500 644 1501
rect 734 1505 740 1506
rect 734 1501 735 1505
rect 739 1501 740 1505
rect 734 1500 740 1501
rect 822 1505 828 1506
rect 822 1501 823 1505
rect 827 1501 828 1505
rect 822 1500 828 1501
rect 902 1505 908 1506
rect 902 1501 903 1505
rect 907 1501 908 1505
rect 902 1500 908 1501
rect 974 1505 980 1506
rect 974 1501 975 1505
rect 979 1501 980 1505
rect 974 1500 980 1501
rect 1046 1505 1052 1506
rect 1046 1501 1047 1505
rect 1051 1501 1052 1505
rect 1046 1500 1052 1501
rect 1118 1505 1124 1506
rect 1118 1501 1119 1505
rect 1123 1501 1124 1505
rect 1118 1500 1124 1501
rect 1190 1505 1196 1506
rect 1190 1501 1191 1505
rect 1195 1501 1196 1505
rect 1190 1500 1196 1501
rect 152 1487 154 1500
rect 200 1487 202 1500
rect 264 1487 266 1500
rect 344 1487 346 1500
rect 440 1487 442 1500
rect 536 1487 538 1500
rect 640 1487 642 1500
rect 736 1487 738 1500
rect 824 1487 826 1500
rect 904 1487 906 1500
rect 976 1487 978 1500
rect 1048 1487 1050 1500
rect 1120 1487 1122 1500
rect 1192 1487 1194 1500
rect 1240 1487 1242 1523
rect 111 1486 115 1487
rect 111 1481 115 1482
rect 151 1486 155 1487
rect 151 1481 155 1482
rect 199 1486 203 1487
rect 199 1481 203 1482
rect 263 1486 267 1487
rect 263 1481 267 1482
rect 319 1486 323 1487
rect 319 1481 323 1482
rect 343 1486 347 1487
rect 343 1481 347 1482
rect 359 1486 363 1487
rect 359 1481 363 1482
rect 399 1486 403 1487
rect 399 1481 403 1482
rect 439 1486 443 1487
rect 439 1481 443 1482
rect 447 1486 451 1487
rect 447 1481 451 1482
rect 503 1486 507 1487
rect 503 1481 507 1482
rect 535 1486 539 1487
rect 535 1481 539 1482
rect 559 1486 563 1487
rect 559 1481 563 1482
rect 615 1486 619 1487
rect 615 1481 619 1482
rect 639 1486 643 1487
rect 639 1481 643 1482
rect 671 1486 675 1487
rect 671 1481 675 1482
rect 735 1486 739 1487
rect 735 1481 739 1482
rect 799 1486 803 1487
rect 799 1481 803 1482
rect 823 1486 827 1487
rect 823 1481 827 1482
rect 855 1486 859 1487
rect 855 1481 859 1482
rect 903 1486 907 1487
rect 903 1481 907 1482
rect 911 1486 915 1487
rect 911 1481 915 1482
rect 967 1486 971 1487
rect 967 1481 971 1482
rect 975 1486 979 1487
rect 975 1481 979 1482
rect 1023 1486 1027 1487
rect 1023 1481 1027 1482
rect 1047 1486 1051 1487
rect 1047 1481 1051 1482
rect 1087 1486 1091 1487
rect 1087 1481 1091 1482
rect 1119 1486 1123 1487
rect 1119 1481 1123 1482
rect 1151 1486 1155 1487
rect 1151 1481 1155 1482
rect 1191 1486 1195 1487
rect 1191 1481 1195 1482
rect 1239 1486 1243 1487
rect 1239 1481 1243 1482
rect 112 1449 114 1481
rect 320 1472 322 1481
rect 360 1472 362 1481
rect 400 1472 402 1481
rect 448 1472 450 1481
rect 504 1472 506 1481
rect 560 1472 562 1481
rect 616 1472 618 1481
rect 672 1472 674 1481
rect 736 1472 738 1481
rect 800 1472 802 1481
rect 856 1472 858 1481
rect 912 1472 914 1481
rect 968 1472 970 1481
rect 1024 1472 1026 1481
rect 1088 1472 1090 1481
rect 1152 1472 1154 1481
rect 1192 1472 1194 1481
rect 318 1471 324 1472
rect 318 1467 319 1471
rect 323 1467 324 1471
rect 318 1466 324 1467
rect 358 1471 364 1472
rect 358 1467 359 1471
rect 363 1467 364 1471
rect 358 1466 364 1467
rect 398 1471 404 1472
rect 398 1467 399 1471
rect 403 1467 404 1471
rect 398 1466 404 1467
rect 446 1471 452 1472
rect 446 1467 447 1471
rect 451 1467 452 1471
rect 446 1466 452 1467
rect 502 1471 508 1472
rect 502 1467 503 1471
rect 507 1467 508 1471
rect 502 1466 508 1467
rect 558 1471 564 1472
rect 558 1467 559 1471
rect 563 1467 564 1471
rect 558 1466 564 1467
rect 614 1471 620 1472
rect 614 1467 615 1471
rect 619 1467 620 1471
rect 614 1466 620 1467
rect 670 1471 676 1472
rect 670 1467 671 1471
rect 675 1467 676 1471
rect 670 1466 676 1467
rect 734 1471 740 1472
rect 734 1467 735 1471
rect 739 1467 740 1471
rect 734 1466 740 1467
rect 798 1471 804 1472
rect 798 1467 799 1471
rect 803 1467 804 1471
rect 798 1466 804 1467
rect 854 1471 860 1472
rect 854 1467 855 1471
rect 859 1467 860 1471
rect 854 1466 860 1467
rect 910 1471 916 1472
rect 910 1467 911 1471
rect 915 1467 916 1471
rect 910 1466 916 1467
rect 966 1471 972 1472
rect 966 1467 967 1471
rect 971 1467 972 1471
rect 966 1466 972 1467
rect 1022 1471 1028 1472
rect 1022 1467 1023 1471
rect 1027 1467 1028 1471
rect 1022 1466 1028 1467
rect 1086 1471 1092 1472
rect 1086 1467 1087 1471
rect 1091 1467 1092 1471
rect 1086 1466 1092 1467
rect 1150 1471 1156 1472
rect 1150 1467 1151 1471
rect 1155 1467 1156 1471
rect 1150 1466 1156 1467
rect 1190 1471 1196 1472
rect 1190 1467 1191 1471
rect 1195 1467 1196 1471
rect 1190 1466 1196 1467
rect 1240 1449 1242 1481
rect 1280 1475 1282 1527
rect 1470 1509 1476 1510
rect 1470 1505 1471 1509
rect 1475 1505 1476 1509
rect 1470 1504 1476 1505
rect 1622 1509 1628 1510
rect 1622 1505 1623 1509
rect 1627 1505 1628 1509
rect 1622 1504 1628 1505
rect 1758 1509 1764 1510
rect 1758 1505 1759 1509
rect 1763 1505 1764 1509
rect 1758 1504 1764 1505
rect 1870 1509 1876 1510
rect 1870 1505 1871 1509
rect 1875 1505 1876 1509
rect 1870 1504 1876 1505
rect 1966 1509 1972 1510
rect 1966 1505 1967 1509
rect 1971 1505 1972 1509
rect 1966 1504 1972 1505
rect 2054 1509 2060 1510
rect 2054 1505 2055 1509
rect 2059 1505 2060 1509
rect 2054 1504 2060 1505
rect 2126 1509 2132 1510
rect 2126 1505 2127 1509
rect 2131 1505 2132 1509
rect 2126 1504 2132 1505
rect 2190 1509 2196 1510
rect 2190 1505 2191 1509
rect 2195 1505 2196 1509
rect 2190 1504 2196 1505
rect 2254 1509 2260 1510
rect 2254 1505 2255 1509
rect 2259 1505 2260 1509
rect 2254 1504 2260 1505
rect 2318 1509 2324 1510
rect 2318 1505 2319 1509
rect 2323 1505 2324 1509
rect 2318 1504 2324 1505
rect 2358 1509 2364 1510
rect 2358 1505 2359 1509
rect 2363 1505 2364 1509
rect 2358 1504 2364 1505
rect 1472 1475 1474 1504
rect 1624 1475 1626 1504
rect 1760 1475 1762 1504
rect 1872 1475 1874 1504
rect 1968 1475 1970 1504
rect 2056 1475 2058 1504
rect 2128 1475 2130 1504
rect 2192 1475 2194 1504
rect 2256 1475 2258 1504
rect 2320 1475 2322 1504
rect 2360 1475 2362 1504
rect 2408 1475 2410 1527
rect 1279 1474 1283 1475
rect 1279 1469 1283 1470
rect 1303 1474 1307 1475
rect 1303 1469 1307 1470
rect 1375 1474 1379 1475
rect 1375 1469 1379 1470
rect 1471 1474 1475 1475
rect 1471 1469 1475 1470
rect 1479 1474 1483 1475
rect 1479 1469 1483 1470
rect 1583 1474 1587 1475
rect 1583 1469 1587 1470
rect 1623 1474 1627 1475
rect 1623 1469 1627 1470
rect 1687 1474 1691 1475
rect 1687 1469 1691 1470
rect 1759 1474 1763 1475
rect 1759 1469 1763 1470
rect 1783 1474 1787 1475
rect 1783 1469 1787 1470
rect 1871 1474 1875 1475
rect 1871 1469 1875 1470
rect 1951 1474 1955 1475
rect 1951 1469 1955 1470
rect 1967 1474 1971 1475
rect 1967 1469 1971 1470
rect 2031 1474 2035 1475
rect 2031 1469 2035 1470
rect 2055 1474 2059 1475
rect 2055 1469 2059 1470
rect 2103 1474 2107 1475
rect 2103 1469 2107 1470
rect 2127 1474 2131 1475
rect 2127 1469 2131 1470
rect 2167 1474 2171 1475
rect 2167 1469 2171 1470
rect 2191 1474 2195 1475
rect 2191 1469 2195 1470
rect 2239 1474 2243 1475
rect 2239 1469 2243 1470
rect 2255 1474 2259 1475
rect 2255 1469 2259 1470
rect 2311 1474 2315 1475
rect 2311 1469 2315 1470
rect 2319 1474 2323 1475
rect 2319 1469 2323 1470
rect 2359 1474 2363 1475
rect 2359 1469 2363 1470
rect 2407 1474 2411 1475
rect 2407 1469 2411 1470
rect 110 1448 116 1449
rect 110 1444 111 1448
rect 115 1444 116 1448
rect 110 1443 116 1444
rect 1238 1448 1244 1449
rect 1238 1444 1239 1448
rect 1243 1444 1244 1448
rect 1238 1443 1244 1444
rect 1280 1437 1282 1469
rect 1304 1460 1306 1469
rect 1376 1460 1378 1469
rect 1480 1460 1482 1469
rect 1584 1460 1586 1469
rect 1688 1460 1690 1469
rect 1784 1460 1786 1469
rect 1872 1460 1874 1469
rect 1952 1460 1954 1469
rect 2032 1460 2034 1469
rect 2104 1460 2106 1469
rect 2168 1460 2170 1469
rect 2240 1460 2242 1469
rect 2312 1460 2314 1469
rect 2360 1460 2362 1469
rect 1302 1459 1308 1460
rect 1302 1455 1303 1459
rect 1307 1455 1308 1459
rect 1302 1454 1308 1455
rect 1374 1459 1380 1460
rect 1374 1455 1375 1459
rect 1379 1455 1380 1459
rect 1374 1454 1380 1455
rect 1478 1459 1484 1460
rect 1478 1455 1479 1459
rect 1483 1455 1484 1459
rect 1478 1454 1484 1455
rect 1582 1459 1588 1460
rect 1582 1455 1583 1459
rect 1587 1455 1588 1459
rect 1582 1454 1588 1455
rect 1686 1459 1692 1460
rect 1686 1455 1687 1459
rect 1691 1455 1692 1459
rect 1686 1454 1692 1455
rect 1782 1459 1788 1460
rect 1782 1455 1783 1459
rect 1787 1455 1788 1459
rect 1782 1454 1788 1455
rect 1870 1459 1876 1460
rect 1870 1455 1871 1459
rect 1875 1455 1876 1459
rect 1870 1454 1876 1455
rect 1950 1459 1956 1460
rect 1950 1455 1951 1459
rect 1955 1455 1956 1459
rect 1950 1454 1956 1455
rect 2030 1459 2036 1460
rect 2030 1455 2031 1459
rect 2035 1455 2036 1459
rect 2030 1454 2036 1455
rect 2102 1459 2108 1460
rect 2102 1455 2103 1459
rect 2107 1455 2108 1459
rect 2102 1454 2108 1455
rect 2166 1459 2172 1460
rect 2166 1455 2167 1459
rect 2171 1455 2172 1459
rect 2166 1454 2172 1455
rect 2238 1459 2244 1460
rect 2238 1455 2239 1459
rect 2243 1455 2244 1459
rect 2238 1454 2244 1455
rect 2310 1459 2316 1460
rect 2310 1455 2311 1459
rect 2315 1455 2316 1459
rect 2310 1454 2316 1455
rect 2358 1459 2364 1460
rect 2358 1455 2359 1459
rect 2363 1455 2364 1459
rect 2358 1454 2364 1455
rect 2408 1437 2410 1469
rect 1278 1436 1284 1437
rect 1278 1432 1279 1436
rect 1283 1432 1284 1436
rect 110 1431 116 1432
rect 110 1427 111 1431
rect 115 1427 116 1431
rect 110 1426 116 1427
rect 1238 1431 1244 1432
rect 1278 1431 1284 1432
rect 2406 1436 2412 1437
rect 2406 1432 2407 1436
rect 2411 1432 2412 1436
rect 2406 1431 2412 1432
rect 1238 1427 1239 1431
rect 1243 1427 1244 1431
rect 1238 1426 1244 1427
rect 112 1415 114 1426
rect 318 1424 324 1425
rect 318 1420 319 1424
rect 323 1420 324 1424
rect 318 1419 324 1420
rect 358 1424 364 1425
rect 358 1420 359 1424
rect 363 1420 364 1424
rect 358 1419 364 1420
rect 398 1424 404 1425
rect 398 1420 399 1424
rect 403 1420 404 1424
rect 398 1419 404 1420
rect 446 1424 452 1425
rect 446 1420 447 1424
rect 451 1420 452 1424
rect 446 1419 452 1420
rect 502 1424 508 1425
rect 502 1420 503 1424
rect 507 1420 508 1424
rect 502 1419 508 1420
rect 558 1424 564 1425
rect 558 1420 559 1424
rect 563 1420 564 1424
rect 558 1419 564 1420
rect 614 1424 620 1425
rect 614 1420 615 1424
rect 619 1420 620 1424
rect 614 1419 620 1420
rect 670 1424 676 1425
rect 670 1420 671 1424
rect 675 1420 676 1424
rect 670 1419 676 1420
rect 734 1424 740 1425
rect 734 1420 735 1424
rect 739 1420 740 1424
rect 734 1419 740 1420
rect 798 1424 804 1425
rect 798 1420 799 1424
rect 803 1420 804 1424
rect 798 1419 804 1420
rect 854 1424 860 1425
rect 854 1420 855 1424
rect 859 1420 860 1424
rect 854 1419 860 1420
rect 910 1424 916 1425
rect 910 1420 911 1424
rect 915 1420 916 1424
rect 910 1419 916 1420
rect 966 1424 972 1425
rect 966 1420 967 1424
rect 971 1420 972 1424
rect 966 1419 972 1420
rect 1022 1424 1028 1425
rect 1022 1420 1023 1424
rect 1027 1420 1028 1424
rect 1022 1419 1028 1420
rect 1086 1424 1092 1425
rect 1086 1420 1087 1424
rect 1091 1420 1092 1424
rect 1086 1419 1092 1420
rect 1150 1424 1156 1425
rect 1150 1420 1151 1424
rect 1155 1420 1156 1424
rect 1150 1419 1156 1420
rect 1190 1424 1196 1425
rect 1190 1420 1191 1424
rect 1195 1420 1196 1424
rect 1190 1419 1196 1420
rect 320 1415 322 1419
rect 360 1415 362 1419
rect 400 1415 402 1419
rect 448 1415 450 1419
rect 504 1415 506 1419
rect 560 1415 562 1419
rect 616 1415 618 1419
rect 672 1415 674 1419
rect 736 1415 738 1419
rect 800 1415 802 1419
rect 856 1415 858 1419
rect 912 1415 914 1419
rect 968 1415 970 1419
rect 1024 1415 1026 1419
rect 1088 1415 1090 1419
rect 1152 1415 1154 1419
rect 1192 1415 1194 1419
rect 1240 1415 1242 1426
rect 1278 1419 1284 1420
rect 1278 1415 1279 1419
rect 1283 1415 1284 1419
rect 111 1414 115 1415
rect 111 1409 115 1410
rect 263 1414 267 1415
rect 263 1409 267 1410
rect 303 1414 307 1415
rect 303 1409 307 1410
rect 319 1414 323 1415
rect 319 1409 323 1410
rect 343 1414 347 1415
rect 343 1409 347 1410
rect 359 1414 363 1415
rect 359 1409 363 1410
rect 391 1414 395 1415
rect 391 1409 395 1410
rect 399 1414 403 1415
rect 399 1409 403 1410
rect 447 1414 451 1415
rect 447 1409 451 1410
rect 503 1414 507 1415
rect 503 1409 507 1410
rect 559 1414 563 1415
rect 559 1409 563 1410
rect 615 1414 619 1415
rect 615 1409 619 1410
rect 623 1414 627 1415
rect 623 1409 627 1410
rect 671 1414 675 1415
rect 671 1409 675 1410
rect 687 1414 691 1415
rect 687 1409 691 1410
rect 735 1414 739 1415
rect 735 1409 739 1410
rect 751 1414 755 1415
rect 751 1409 755 1410
rect 799 1414 803 1415
rect 799 1409 803 1410
rect 815 1414 819 1415
rect 815 1409 819 1410
rect 855 1414 859 1415
rect 855 1409 859 1410
rect 879 1414 883 1415
rect 879 1409 883 1410
rect 911 1414 915 1415
rect 911 1409 915 1410
rect 951 1414 955 1415
rect 951 1409 955 1410
rect 967 1414 971 1415
rect 967 1409 971 1410
rect 1023 1414 1027 1415
rect 1023 1409 1027 1410
rect 1087 1414 1091 1415
rect 1087 1409 1091 1410
rect 1151 1414 1155 1415
rect 1151 1409 1155 1410
rect 1191 1414 1195 1415
rect 1191 1409 1195 1410
rect 1239 1414 1243 1415
rect 1278 1414 1284 1415
rect 2406 1419 2412 1420
rect 2406 1415 2407 1419
rect 2411 1415 2412 1419
rect 2406 1414 2412 1415
rect 1239 1409 1243 1410
rect 112 1402 114 1409
rect 262 1408 268 1409
rect 262 1404 263 1408
rect 267 1404 268 1408
rect 262 1403 268 1404
rect 302 1408 308 1409
rect 302 1404 303 1408
rect 307 1404 308 1408
rect 302 1403 308 1404
rect 342 1408 348 1409
rect 342 1404 343 1408
rect 347 1404 348 1408
rect 342 1403 348 1404
rect 390 1408 396 1409
rect 390 1404 391 1408
rect 395 1404 396 1408
rect 390 1403 396 1404
rect 446 1408 452 1409
rect 446 1404 447 1408
rect 451 1404 452 1408
rect 446 1403 452 1404
rect 502 1408 508 1409
rect 502 1404 503 1408
rect 507 1404 508 1408
rect 502 1403 508 1404
rect 558 1408 564 1409
rect 558 1404 559 1408
rect 563 1404 564 1408
rect 558 1403 564 1404
rect 622 1408 628 1409
rect 622 1404 623 1408
rect 627 1404 628 1408
rect 622 1403 628 1404
rect 686 1408 692 1409
rect 686 1404 687 1408
rect 691 1404 692 1408
rect 686 1403 692 1404
rect 750 1408 756 1409
rect 750 1404 751 1408
rect 755 1404 756 1408
rect 750 1403 756 1404
rect 814 1408 820 1409
rect 814 1404 815 1408
rect 819 1404 820 1408
rect 814 1403 820 1404
rect 878 1408 884 1409
rect 878 1404 879 1408
rect 883 1404 884 1408
rect 878 1403 884 1404
rect 950 1408 956 1409
rect 950 1404 951 1408
rect 955 1404 956 1408
rect 950 1403 956 1404
rect 1022 1408 1028 1409
rect 1022 1404 1023 1408
rect 1027 1404 1028 1408
rect 1022 1403 1028 1404
rect 1240 1402 1242 1409
rect 1280 1407 1282 1414
rect 1302 1412 1308 1413
rect 1302 1408 1303 1412
rect 1307 1408 1308 1412
rect 1302 1407 1308 1408
rect 1374 1412 1380 1413
rect 1374 1408 1375 1412
rect 1379 1408 1380 1412
rect 1374 1407 1380 1408
rect 1478 1412 1484 1413
rect 1478 1408 1479 1412
rect 1483 1408 1484 1412
rect 1478 1407 1484 1408
rect 1582 1412 1588 1413
rect 1582 1408 1583 1412
rect 1587 1408 1588 1412
rect 1582 1407 1588 1408
rect 1686 1412 1692 1413
rect 1686 1408 1687 1412
rect 1691 1408 1692 1412
rect 1686 1407 1692 1408
rect 1782 1412 1788 1413
rect 1782 1408 1783 1412
rect 1787 1408 1788 1412
rect 1782 1407 1788 1408
rect 1870 1412 1876 1413
rect 1870 1408 1871 1412
rect 1875 1408 1876 1412
rect 1870 1407 1876 1408
rect 1950 1412 1956 1413
rect 1950 1408 1951 1412
rect 1955 1408 1956 1412
rect 1950 1407 1956 1408
rect 2030 1412 2036 1413
rect 2030 1408 2031 1412
rect 2035 1408 2036 1412
rect 2030 1407 2036 1408
rect 2102 1412 2108 1413
rect 2102 1408 2103 1412
rect 2107 1408 2108 1412
rect 2102 1407 2108 1408
rect 2166 1412 2172 1413
rect 2166 1408 2167 1412
rect 2171 1408 2172 1412
rect 2166 1407 2172 1408
rect 2238 1412 2244 1413
rect 2238 1408 2239 1412
rect 2243 1408 2244 1412
rect 2238 1407 2244 1408
rect 2310 1412 2316 1413
rect 2310 1408 2311 1412
rect 2315 1408 2316 1412
rect 2310 1407 2316 1408
rect 2358 1412 2364 1413
rect 2358 1408 2359 1412
rect 2363 1408 2364 1412
rect 2358 1407 2364 1408
rect 2408 1407 2410 1414
rect 1279 1406 1283 1407
rect 110 1401 116 1402
rect 110 1397 111 1401
rect 115 1397 116 1401
rect 110 1396 116 1397
rect 1238 1401 1244 1402
rect 1279 1401 1283 1402
rect 1303 1406 1307 1407
rect 1303 1401 1307 1402
rect 1343 1406 1347 1407
rect 1343 1401 1347 1402
rect 1375 1406 1379 1407
rect 1375 1401 1379 1402
rect 1399 1406 1403 1407
rect 1399 1401 1403 1402
rect 1471 1406 1475 1407
rect 1471 1401 1475 1402
rect 1479 1406 1483 1407
rect 1479 1401 1483 1402
rect 1551 1406 1555 1407
rect 1551 1401 1555 1402
rect 1583 1406 1587 1407
rect 1583 1401 1587 1402
rect 1639 1406 1643 1407
rect 1639 1401 1643 1402
rect 1687 1406 1691 1407
rect 1687 1401 1691 1402
rect 1727 1406 1731 1407
rect 1727 1401 1731 1402
rect 1783 1406 1787 1407
rect 1783 1401 1787 1402
rect 1815 1406 1819 1407
rect 1815 1401 1819 1402
rect 1871 1406 1875 1407
rect 1871 1401 1875 1402
rect 1903 1406 1907 1407
rect 1903 1401 1907 1402
rect 1951 1406 1955 1407
rect 1951 1401 1955 1402
rect 1991 1406 1995 1407
rect 1991 1401 1995 1402
rect 2031 1406 2035 1407
rect 2031 1401 2035 1402
rect 2071 1406 2075 1407
rect 2071 1401 2075 1402
rect 2103 1406 2107 1407
rect 2103 1401 2107 1402
rect 2151 1406 2155 1407
rect 2151 1401 2155 1402
rect 2167 1406 2171 1407
rect 2167 1401 2171 1402
rect 2223 1406 2227 1407
rect 2223 1401 2227 1402
rect 2239 1406 2243 1407
rect 2239 1401 2243 1402
rect 2303 1406 2307 1407
rect 2303 1401 2307 1402
rect 2311 1406 2315 1407
rect 2311 1401 2315 1402
rect 2359 1406 2363 1407
rect 2359 1401 2363 1402
rect 2407 1406 2411 1407
rect 2407 1401 2411 1402
rect 1238 1397 1239 1401
rect 1243 1397 1244 1401
rect 1238 1396 1244 1397
rect 1280 1394 1282 1401
rect 1302 1400 1308 1401
rect 1302 1396 1303 1400
rect 1307 1396 1308 1400
rect 1302 1395 1308 1396
rect 1342 1400 1348 1401
rect 1342 1396 1343 1400
rect 1347 1396 1348 1400
rect 1342 1395 1348 1396
rect 1398 1400 1404 1401
rect 1398 1396 1399 1400
rect 1403 1396 1404 1400
rect 1398 1395 1404 1396
rect 1470 1400 1476 1401
rect 1470 1396 1471 1400
rect 1475 1396 1476 1400
rect 1470 1395 1476 1396
rect 1550 1400 1556 1401
rect 1550 1396 1551 1400
rect 1555 1396 1556 1400
rect 1550 1395 1556 1396
rect 1638 1400 1644 1401
rect 1638 1396 1639 1400
rect 1643 1396 1644 1400
rect 1638 1395 1644 1396
rect 1726 1400 1732 1401
rect 1726 1396 1727 1400
rect 1731 1396 1732 1400
rect 1726 1395 1732 1396
rect 1814 1400 1820 1401
rect 1814 1396 1815 1400
rect 1819 1396 1820 1400
rect 1814 1395 1820 1396
rect 1902 1400 1908 1401
rect 1902 1396 1903 1400
rect 1907 1396 1908 1400
rect 1902 1395 1908 1396
rect 1990 1400 1996 1401
rect 1990 1396 1991 1400
rect 1995 1396 1996 1400
rect 1990 1395 1996 1396
rect 2070 1400 2076 1401
rect 2070 1396 2071 1400
rect 2075 1396 2076 1400
rect 2070 1395 2076 1396
rect 2150 1400 2156 1401
rect 2150 1396 2151 1400
rect 2155 1396 2156 1400
rect 2150 1395 2156 1396
rect 2222 1400 2228 1401
rect 2222 1396 2223 1400
rect 2227 1396 2228 1400
rect 2222 1395 2228 1396
rect 2302 1400 2308 1401
rect 2302 1396 2303 1400
rect 2307 1396 2308 1400
rect 2302 1395 2308 1396
rect 2358 1400 2364 1401
rect 2358 1396 2359 1400
rect 2363 1396 2364 1400
rect 2358 1395 2364 1396
rect 2408 1394 2410 1401
rect 1278 1393 1284 1394
rect 1278 1389 1279 1393
rect 1283 1389 1284 1393
rect 1278 1388 1284 1389
rect 2406 1393 2412 1394
rect 2406 1389 2407 1393
rect 2411 1389 2412 1393
rect 2406 1388 2412 1389
rect 110 1384 116 1385
rect 110 1380 111 1384
rect 115 1380 116 1384
rect 110 1379 116 1380
rect 1238 1384 1244 1385
rect 1238 1380 1239 1384
rect 1243 1380 1244 1384
rect 1238 1379 1244 1380
rect 112 1343 114 1379
rect 262 1361 268 1362
rect 262 1357 263 1361
rect 267 1357 268 1361
rect 262 1356 268 1357
rect 302 1361 308 1362
rect 302 1357 303 1361
rect 307 1357 308 1361
rect 302 1356 308 1357
rect 342 1361 348 1362
rect 342 1357 343 1361
rect 347 1357 348 1361
rect 342 1356 348 1357
rect 390 1361 396 1362
rect 390 1357 391 1361
rect 395 1357 396 1361
rect 390 1356 396 1357
rect 446 1361 452 1362
rect 446 1357 447 1361
rect 451 1357 452 1361
rect 446 1356 452 1357
rect 502 1361 508 1362
rect 502 1357 503 1361
rect 507 1357 508 1361
rect 502 1356 508 1357
rect 558 1361 564 1362
rect 558 1357 559 1361
rect 563 1357 564 1361
rect 558 1356 564 1357
rect 622 1361 628 1362
rect 622 1357 623 1361
rect 627 1357 628 1361
rect 622 1356 628 1357
rect 686 1361 692 1362
rect 686 1357 687 1361
rect 691 1357 692 1361
rect 686 1356 692 1357
rect 750 1361 756 1362
rect 750 1357 751 1361
rect 755 1357 756 1361
rect 750 1356 756 1357
rect 814 1361 820 1362
rect 814 1357 815 1361
rect 819 1357 820 1361
rect 814 1356 820 1357
rect 878 1361 884 1362
rect 878 1357 879 1361
rect 883 1357 884 1361
rect 878 1356 884 1357
rect 950 1361 956 1362
rect 950 1357 951 1361
rect 955 1357 956 1361
rect 950 1356 956 1357
rect 1022 1361 1028 1362
rect 1022 1357 1023 1361
rect 1027 1357 1028 1361
rect 1022 1356 1028 1357
rect 264 1343 266 1356
rect 304 1343 306 1356
rect 344 1343 346 1356
rect 392 1343 394 1356
rect 448 1343 450 1356
rect 504 1343 506 1356
rect 560 1343 562 1356
rect 624 1343 626 1356
rect 688 1343 690 1356
rect 752 1343 754 1356
rect 816 1343 818 1356
rect 880 1343 882 1356
rect 952 1343 954 1356
rect 1024 1343 1026 1356
rect 1240 1343 1242 1379
rect 1278 1376 1284 1377
rect 1278 1372 1279 1376
rect 1283 1372 1284 1376
rect 1278 1371 1284 1372
rect 2406 1376 2412 1377
rect 2406 1372 2407 1376
rect 2411 1372 2412 1376
rect 2406 1371 2412 1372
rect 111 1342 115 1343
rect 111 1337 115 1338
rect 135 1342 139 1343
rect 135 1337 139 1338
rect 175 1342 179 1343
rect 175 1337 179 1338
rect 215 1342 219 1343
rect 215 1337 219 1338
rect 255 1342 259 1343
rect 255 1337 259 1338
rect 263 1342 267 1343
rect 263 1337 267 1338
rect 303 1342 307 1343
rect 303 1337 307 1338
rect 327 1342 331 1343
rect 327 1337 331 1338
rect 343 1342 347 1343
rect 343 1337 347 1338
rect 391 1342 395 1343
rect 391 1337 395 1338
rect 407 1342 411 1343
rect 407 1337 411 1338
rect 447 1342 451 1343
rect 447 1337 451 1338
rect 495 1342 499 1343
rect 495 1337 499 1338
rect 503 1342 507 1343
rect 503 1337 507 1338
rect 559 1342 563 1343
rect 559 1337 563 1338
rect 583 1342 587 1343
rect 583 1337 587 1338
rect 623 1342 627 1343
rect 623 1337 627 1338
rect 671 1342 675 1343
rect 671 1337 675 1338
rect 687 1342 691 1343
rect 687 1337 691 1338
rect 751 1342 755 1343
rect 751 1337 755 1338
rect 759 1342 763 1343
rect 759 1337 763 1338
rect 815 1342 819 1343
rect 815 1337 819 1338
rect 839 1342 843 1343
rect 839 1337 843 1338
rect 879 1342 883 1343
rect 879 1337 883 1338
rect 919 1342 923 1343
rect 919 1337 923 1338
rect 951 1342 955 1343
rect 951 1337 955 1338
rect 1007 1342 1011 1343
rect 1007 1337 1011 1338
rect 1023 1342 1027 1343
rect 1023 1337 1027 1338
rect 1095 1342 1099 1343
rect 1095 1337 1099 1338
rect 1239 1342 1243 1343
rect 1239 1337 1243 1338
rect 112 1305 114 1337
rect 136 1328 138 1337
rect 176 1328 178 1337
rect 216 1328 218 1337
rect 256 1328 258 1337
rect 328 1328 330 1337
rect 408 1328 410 1337
rect 496 1328 498 1337
rect 584 1328 586 1337
rect 672 1328 674 1337
rect 760 1328 762 1337
rect 840 1328 842 1337
rect 920 1328 922 1337
rect 1008 1328 1010 1337
rect 1096 1328 1098 1337
rect 134 1327 140 1328
rect 134 1323 135 1327
rect 139 1323 140 1327
rect 134 1322 140 1323
rect 174 1327 180 1328
rect 174 1323 175 1327
rect 179 1323 180 1327
rect 174 1322 180 1323
rect 214 1327 220 1328
rect 214 1323 215 1327
rect 219 1323 220 1327
rect 214 1322 220 1323
rect 254 1327 260 1328
rect 254 1323 255 1327
rect 259 1323 260 1327
rect 254 1322 260 1323
rect 326 1327 332 1328
rect 326 1323 327 1327
rect 331 1323 332 1327
rect 326 1322 332 1323
rect 406 1327 412 1328
rect 406 1323 407 1327
rect 411 1323 412 1327
rect 406 1322 412 1323
rect 494 1327 500 1328
rect 494 1323 495 1327
rect 499 1323 500 1327
rect 494 1322 500 1323
rect 582 1327 588 1328
rect 582 1323 583 1327
rect 587 1323 588 1327
rect 582 1322 588 1323
rect 670 1327 676 1328
rect 670 1323 671 1327
rect 675 1323 676 1327
rect 670 1322 676 1323
rect 758 1327 764 1328
rect 758 1323 759 1327
rect 763 1323 764 1327
rect 758 1322 764 1323
rect 838 1327 844 1328
rect 838 1323 839 1327
rect 843 1323 844 1327
rect 838 1322 844 1323
rect 918 1327 924 1328
rect 918 1323 919 1327
rect 923 1323 924 1327
rect 918 1322 924 1323
rect 1006 1327 1012 1328
rect 1006 1323 1007 1327
rect 1011 1323 1012 1327
rect 1006 1322 1012 1323
rect 1094 1327 1100 1328
rect 1094 1323 1095 1327
rect 1099 1323 1100 1327
rect 1094 1322 1100 1323
rect 1240 1305 1242 1337
rect 1280 1335 1282 1371
rect 1302 1353 1308 1354
rect 1302 1349 1303 1353
rect 1307 1349 1308 1353
rect 1302 1348 1308 1349
rect 1342 1353 1348 1354
rect 1342 1349 1343 1353
rect 1347 1349 1348 1353
rect 1342 1348 1348 1349
rect 1398 1353 1404 1354
rect 1398 1349 1399 1353
rect 1403 1349 1404 1353
rect 1398 1348 1404 1349
rect 1470 1353 1476 1354
rect 1470 1349 1471 1353
rect 1475 1349 1476 1353
rect 1470 1348 1476 1349
rect 1550 1353 1556 1354
rect 1550 1349 1551 1353
rect 1555 1349 1556 1353
rect 1550 1348 1556 1349
rect 1638 1353 1644 1354
rect 1638 1349 1639 1353
rect 1643 1349 1644 1353
rect 1638 1348 1644 1349
rect 1726 1353 1732 1354
rect 1726 1349 1727 1353
rect 1731 1349 1732 1353
rect 1726 1348 1732 1349
rect 1814 1353 1820 1354
rect 1814 1349 1815 1353
rect 1819 1349 1820 1353
rect 1814 1348 1820 1349
rect 1902 1353 1908 1354
rect 1902 1349 1903 1353
rect 1907 1349 1908 1353
rect 1902 1348 1908 1349
rect 1990 1353 1996 1354
rect 1990 1349 1991 1353
rect 1995 1349 1996 1353
rect 1990 1348 1996 1349
rect 2070 1353 2076 1354
rect 2070 1349 2071 1353
rect 2075 1349 2076 1353
rect 2070 1348 2076 1349
rect 2150 1353 2156 1354
rect 2150 1349 2151 1353
rect 2155 1349 2156 1353
rect 2150 1348 2156 1349
rect 2222 1353 2228 1354
rect 2222 1349 2223 1353
rect 2227 1349 2228 1353
rect 2222 1348 2228 1349
rect 2302 1353 2308 1354
rect 2302 1349 2303 1353
rect 2307 1349 2308 1353
rect 2302 1348 2308 1349
rect 2358 1353 2364 1354
rect 2358 1349 2359 1353
rect 2363 1349 2364 1353
rect 2358 1348 2364 1349
rect 1304 1335 1306 1348
rect 1344 1335 1346 1348
rect 1400 1335 1402 1348
rect 1472 1335 1474 1348
rect 1552 1335 1554 1348
rect 1640 1335 1642 1348
rect 1728 1335 1730 1348
rect 1816 1335 1818 1348
rect 1904 1335 1906 1348
rect 1992 1335 1994 1348
rect 2072 1335 2074 1348
rect 2152 1335 2154 1348
rect 2224 1335 2226 1348
rect 2304 1335 2306 1348
rect 2360 1335 2362 1348
rect 2408 1335 2410 1371
rect 1279 1334 1283 1335
rect 1279 1329 1283 1330
rect 1303 1334 1307 1335
rect 1303 1329 1307 1330
rect 1343 1334 1347 1335
rect 1343 1329 1347 1330
rect 1399 1334 1403 1335
rect 1399 1329 1403 1330
rect 1447 1334 1451 1335
rect 1447 1329 1451 1330
rect 1471 1334 1475 1335
rect 1471 1329 1475 1330
rect 1487 1334 1491 1335
rect 1487 1329 1491 1330
rect 1527 1334 1531 1335
rect 1527 1329 1531 1330
rect 1551 1334 1555 1335
rect 1551 1329 1555 1330
rect 1567 1334 1571 1335
rect 1567 1329 1571 1330
rect 1615 1334 1619 1335
rect 1615 1329 1619 1330
rect 1639 1334 1643 1335
rect 1639 1329 1643 1330
rect 1671 1334 1675 1335
rect 1671 1329 1675 1330
rect 1719 1334 1723 1335
rect 1719 1329 1723 1330
rect 1727 1334 1731 1335
rect 1727 1329 1731 1330
rect 1775 1334 1779 1335
rect 1775 1329 1779 1330
rect 1815 1334 1819 1335
rect 1815 1329 1819 1330
rect 1831 1334 1835 1335
rect 1831 1329 1835 1330
rect 1903 1334 1907 1335
rect 1903 1329 1907 1330
rect 1983 1334 1987 1335
rect 1983 1329 1987 1330
rect 1991 1334 1995 1335
rect 1991 1329 1995 1330
rect 2071 1334 2075 1335
rect 2071 1329 2075 1330
rect 2151 1334 2155 1335
rect 2151 1329 2155 1330
rect 2167 1334 2171 1335
rect 2167 1329 2171 1330
rect 2223 1334 2227 1335
rect 2223 1329 2227 1330
rect 2271 1334 2275 1335
rect 2271 1329 2275 1330
rect 2303 1334 2307 1335
rect 2303 1329 2307 1330
rect 2359 1334 2363 1335
rect 2359 1329 2363 1330
rect 2407 1334 2411 1335
rect 2407 1329 2411 1330
rect 110 1304 116 1305
rect 110 1300 111 1304
rect 115 1300 116 1304
rect 110 1299 116 1300
rect 1238 1304 1244 1305
rect 1238 1300 1239 1304
rect 1243 1300 1244 1304
rect 1238 1299 1244 1300
rect 1280 1297 1282 1329
rect 1448 1320 1450 1329
rect 1488 1320 1490 1329
rect 1528 1320 1530 1329
rect 1568 1320 1570 1329
rect 1616 1320 1618 1329
rect 1672 1320 1674 1329
rect 1720 1320 1722 1329
rect 1776 1320 1778 1329
rect 1832 1320 1834 1329
rect 1904 1320 1906 1329
rect 1984 1320 1986 1329
rect 2072 1320 2074 1329
rect 2168 1320 2170 1329
rect 2272 1320 2274 1329
rect 2360 1320 2362 1329
rect 1446 1319 1452 1320
rect 1446 1315 1447 1319
rect 1451 1315 1452 1319
rect 1446 1314 1452 1315
rect 1486 1319 1492 1320
rect 1486 1315 1487 1319
rect 1491 1315 1492 1319
rect 1486 1314 1492 1315
rect 1526 1319 1532 1320
rect 1526 1315 1527 1319
rect 1531 1315 1532 1319
rect 1526 1314 1532 1315
rect 1566 1319 1572 1320
rect 1566 1315 1567 1319
rect 1571 1315 1572 1319
rect 1566 1314 1572 1315
rect 1614 1319 1620 1320
rect 1614 1315 1615 1319
rect 1619 1315 1620 1319
rect 1614 1314 1620 1315
rect 1670 1319 1676 1320
rect 1670 1315 1671 1319
rect 1675 1315 1676 1319
rect 1670 1314 1676 1315
rect 1718 1319 1724 1320
rect 1718 1315 1719 1319
rect 1723 1315 1724 1319
rect 1718 1314 1724 1315
rect 1774 1319 1780 1320
rect 1774 1315 1775 1319
rect 1779 1315 1780 1319
rect 1774 1314 1780 1315
rect 1830 1319 1836 1320
rect 1830 1315 1831 1319
rect 1835 1315 1836 1319
rect 1830 1314 1836 1315
rect 1902 1319 1908 1320
rect 1902 1315 1903 1319
rect 1907 1315 1908 1319
rect 1902 1314 1908 1315
rect 1982 1319 1988 1320
rect 1982 1315 1983 1319
rect 1987 1315 1988 1319
rect 1982 1314 1988 1315
rect 2070 1319 2076 1320
rect 2070 1315 2071 1319
rect 2075 1315 2076 1319
rect 2070 1314 2076 1315
rect 2166 1319 2172 1320
rect 2166 1315 2167 1319
rect 2171 1315 2172 1319
rect 2166 1314 2172 1315
rect 2270 1319 2276 1320
rect 2270 1315 2271 1319
rect 2275 1315 2276 1319
rect 2270 1314 2276 1315
rect 2358 1319 2364 1320
rect 2358 1315 2359 1319
rect 2363 1315 2364 1319
rect 2358 1314 2364 1315
rect 2408 1297 2410 1329
rect 1278 1296 1284 1297
rect 1278 1292 1279 1296
rect 1283 1292 1284 1296
rect 1278 1291 1284 1292
rect 2406 1296 2412 1297
rect 2406 1292 2407 1296
rect 2411 1292 2412 1296
rect 2406 1291 2412 1292
rect 110 1287 116 1288
rect 110 1283 111 1287
rect 115 1283 116 1287
rect 110 1282 116 1283
rect 1238 1287 1244 1288
rect 1238 1283 1239 1287
rect 1243 1283 1244 1287
rect 1238 1282 1244 1283
rect 112 1271 114 1282
rect 134 1280 140 1281
rect 134 1276 135 1280
rect 139 1276 140 1280
rect 134 1275 140 1276
rect 174 1280 180 1281
rect 174 1276 175 1280
rect 179 1276 180 1280
rect 174 1275 180 1276
rect 214 1280 220 1281
rect 214 1276 215 1280
rect 219 1276 220 1280
rect 214 1275 220 1276
rect 254 1280 260 1281
rect 254 1276 255 1280
rect 259 1276 260 1280
rect 254 1275 260 1276
rect 326 1280 332 1281
rect 326 1276 327 1280
rect 331 1276 332 1280
rect 326 1275 332 1276
rect 406 1280 412 1281
rect 406 1276 407 1280
rect 411 1276 412 1280
rect 406 1275 412 1276
rect 494 1280 500 1281
rect 494 1276 495 1280
rect 499 1276 500 1280
rect 494 1275 500 1276
rect 582 1280 588 1281
rect 582 1276 583 1280
rect 587 1276 588 1280
rect 582 1275 588 1276
rect 670 1280 676 1281
rect 670 1276 671 1280
rect 675 1276 676 1280
rect 670 1275 676 1276
rect 758 1280 764 1281
rect 758 1276 759 1280
rect 763 1276 764 1280
rect 758 1275 764 1276
rect 838 1280 844 1281
rect 838 1276 839 1280
rect 843 1276 844 1280
rect 838 1275 844 1276
rect 918 1280 924 1281
rect 918 1276 919 1280
rect 923 1276 924 1280
rect 918 1275 924 1276
rect 1006 1280 1012 1281
rect 1006 1276 1007 1280
rect 1011 1276 1012 1280
rect 1006 1275 1012 1276
rect 1094 1280 1100 1281
rect 1094 1276 1095 1280
rect 1099 1276 1100 1280
rect 1094 1275 1100 1276
rect 136 1271 138 1275
rect 176 1271 178 1275
rect 216 1271 218 1275
rect 256 1271 258 1275
rect 328 1271 330 1275
rect 408 1271 410 1275
rect 496 1271 498 1275
rect 584 1271 586 1275
rect 672 1271 674 1275
rect 760 1271 762 1275
rect 840 1271 842 1275
rect 920 1271 922 1275
rect 1008 1271 1010 1275
rect 1096 1271 1098 1275
rect 1240 1271 1242 1282
rect 1278 1279 1284 1280
rect 1278 1275 1279 1279
rect 1283 1275 1284 1279
rect 1278 1274 1284 1275
rect 2406 1279 2412 1280
rect 2406 1275 2407 1279
rect 2411 1275 2412 1279
rect 2406 1274 2412 1275
rect 111 1270 115 1271
rect 111 1265 115 1266
rect 135 1270 139 1271
rect 135 1265 139 1266
rect 175 1270 179 1271
rect 175 1265 179 1266
rect 215 1270 219 1271
rect 215 1265 219 1266
rect 247 1270 251 1271
rect 247 1265 251 1266
rect 255 1270 259 1271
rect 255 1265 259 1266
rect 327 1270 331 1271
rect 327 1265 331 1266
rect 407 1270 411 1271
rect 407 1265 411 1266
rect 415 1270 419 1271
rect 415 1265 419 1266
rect 495 1270 499 1271
rect 495 1265 499 1266
rect 503 1270 507 1271
rect 503 1265 507 1266
rect 583 1270 587 1271
rect 583 1265 587 1266
rect 591 1270 595 1271
rect 591 1265 595 1266
rect 671 1270 675 1271
rect 671 1265 675 1266
rect 743 1270 747 1271
rect 743 1265 747 1266
rect 759 1270 763 1271
rect 759 1265 763 1266
rect 815 1270 819 1271
rect 815 1265 819 1266
rect 839 1270 843 1271
rect 839 1265 843 1266
rect 879 1270 883 1271
rect 879 1265 883 1266
rect 919 1270 923 1271
rect 919 1265 923 1266
rect 943 1270 947 1271
rect 943 1265 947 1266
rect 1007 1270 1011 1271
rect 1007 1265 1011 1266
rect 1071 1270 1075 1271
rect 1071 1265 1075 1266
rect 1095 1270 1099 1271
rect 1095 1265 1099 1266
rect 1239 1270 1243 1271
rect 1239 1265 1243 1266
rect 112 1258 114 1265
rect 134 1264 140 1265
rect 134 1260 135 1264
rect 139 1260 140 1264
rect 134 1259 140 1260
rect 174 1264 180 1265
rect 174 1260 175 1264
rect 179 1260 180 1264
rect 174 1259 180 1260
rect 246 1264 252 1265
rect 246 1260 247 1264
rect 251 1260 252 1264
rect 246 1259 252 1260
rect 326 1264 332 1265
rect 326 1260 327 1264
rect 331 1260 332 1264
rect 326 1259 332 1260
rect 414 1264 420 1265
rect 414 1260 415 1264
rect 419 1260 420 1264
rect 414 1259 420 1260
rect 502 1264 508 1265
rect 502 1260 503 1264
rect 507 1260 508 1264
rect 502 1259 508 1260
rect 590 1264 596 1265
rect 590 1260 591 1264
rect 595 1260 596 1264
rect 590 1259 596 1260
rect 670 1264 676 1265
rect 670 1260 671 1264
rect 675 1260 676 1264
rect 670 1259 676 1260
rect 742 1264 748 1265
rect 742 1260 743 1264
rect 747 1260 748 1264
rect 742 1259 748 1260
rect 814 1264 820 1265
rect 814 1260 815 1264
rect 819 1260 820 1264
rect 814 1259 820 1260
rect 878 1264 884 1265
rect 878 1260 879 1264
rect 883 1260 884 1264
rect 878 1259 884 1260
rect 942 1264 948 1265
rect 942 1260 943 1264
rect 947 1260 948 1264
rect 942 1259 948 1260
rect 1006 1264 1012 1265
rect 1006 1260 1007 1264
rect 1011 1260 1012 1264
rect 1006 1259 1012 1260
rect 1070 1264 1076 1265
rect 1070 1260 1071 1264
rect 1075 1260 1076 1264
rect 1070 1259 1076 1260
rect 1240 1258 1242 1265
rect 1280 1263 1282 1274
rect 1446 1272 1452 1273
rect 1446 1268 1447 1272
rect 1451 1268 1452 1272
rect 1446 1267 1452 1268
rect 1486 1272 1492 1273
rect 1486 1268 1487 1272
rect 1491 1268 1492 1272
rect 1486 1267 1492 1268
rect 1526 1272 1532 1273
rect 1526 1268 1527 1272
rect 1531 1268 1532 1272
rect 1526 1267 1532 1268
rect 1566 1272 1572 1273
rect 1566 1268 1567 1272
rect 1571 1268 1572 1272
rect 1566 1267 1572 1268
rect 1614 1272 1620 1273
rect 1614 1268 1615 1272
rect 1619 1268 1620 1272
rect 1614 1267 1620 1268
rect 1670 1272 1676 1273
rect 1670 1268 1671 1272
rect 1675 1268 1676 1272
rect 1670 1267 1676 1268
rect 1718 1272 1724 1273
rect 1718 1268 1719 1272
rect 1723 1268 1724 1272
rect 1718 1267 1724 1268
rect 1774 1272 1780 1273
rect 1774 1268 1775 1272
rect 1779 1268 1780 1272
rect 1774 1267 1780 1268
rect 1830 1272 1836 1273
rect 1830 1268 1831 1272
rect 1835 1268 1836 1272
rect 1830 1267 1836 1268
rect 1902 1272 1908 1273
rect 1902 1268 1903 1272
rect 1907 1268 1908 1272
rect 1902 1267 1908 1268
rect 1982 1272 1988 1273
rect 1982 1268 1983 1272
rect 1987 1268 1988 1272
rect 1982 1267 1988 1268
rect 2070 1272 2076 1273
rect 2070 1268 2071 1272
rect 2075 1268 2076 1272
rect 2070 1267 2076 1268
rect 2166 1272 2172 1273
rect 2166 1268 2167 1272
rect 2171 1268 2172 1272
rect 2166 1267 2172 1268
rect 2270 1272 2276 1273
rect 2270 1268 2271 1272
rect 2275 1268 2276 1272
rect 2270 1267 2276 1268
rect 2358 1272 2364 1273
rect 2358 1268 2359 1272
rect 2363 1268 2364 1272
rect 2358 1267 2364 1268
rect 1448 1263 1450 1267
rect 1488 1263 1490 1267
rect 1528 1263 1530 1267
rect 1568 1263 1570 1267
rect 1616 1263 1618 1267
rect 1672 1263 1674 1267
rect 1720 1263 1722 1267
rect 1776 1263 1778 1267
rect 1832 1263 1834 1267
rect 1904 1263 1906 1267
rect 1984 1263 1986 1267
rect 2072 1263 2074 1267
rect 2168 1263 2170 1267
rect 2272 1263 2274 1267
rect 2360 1263 2362 1267
rect 2408 1263 2410 1274
rect 1279 1262 1283 1263
rect 110 1257 116 1258
rect 110 1253 111 1257
rect 115 1253 116 1257
rect 110 1252 116 1253
rect 1238 1257 1244 1258
rect 1279 1257 1283 1258
rect 1447 1262 1451 1263
rect 1447 1257 1451 1258
rect 1487 1262 1491 1263
rect 1487 1257 1491 1258
rect 1511 1262 1515 1263
rect 1511 1257 1515 1258
rect 1527 1262 1531 1263
rect 1527 1257 1531 1258
rect 1551 1262 1555 1263
rect 1551 1257 1555 1258
rect 1567 1262 1571 1263
rect 1567 1257 1571 1258
rect 1591 1262 1595 1263
rect 1591 1257 1595 1258
rect 1615 1262 1619 1263
rect 1615 1257 1619 1258
rect 1631 1262 1635 1263
rect 1631 1257 1635 1258
rect 1671 1262 1675 1263
rect 1671 1257 1675 1258
rect 1711 1262 1715 1263
rect 1711 1257 1715 1258
rect 1719 1262 1723 1263
rect 1719 1257 1723 1258
rect 1751 1262 1755 1263
rect 1751 1257 1755 1258
rect 1775 1262 1779 1263
rect 1775 1257 1779 1258
rect 1791 1262 1795 1263
rect 1791 1257 1795 1258
rect 1831 1262 1835 1263
rect 1831 1257 1835 1258
rect 1839 1262 1843 1263
rect 1839 1257 1843 1258
rect 1903 1262 1907 1263
rect 1903 1257 1907 1258
rect 1967 1262 1971 1263
rect 1967 1257 1971 1258
rect 1983 1262 1987 1263
rect 1983 1257 1987 1258
rect 2039 1262 2043 1263
rect 2039 1257 2043 1258
rect 2071 1262 2075 1263
rect 2071 1257 2075 1258
rect 2119 1262 2123 1263
rect 2119 1257 2123 1258
rect 2167 1262 2171 1263
rect 2167 1257 2171 1258
rect 2207 1262 2211 1263
rect 2207 1257 2211 1258
rect 2271 1262 2275 1263
rect 2271 1257 2275 1258
rect 2295 1262 2299 1263
rect 2295 1257 2299 1258
rect 2359 1262 2363 1263
rect 2359 1257 2363 1258
rect 2407 1262 2411 1263
rect 2407 1257 2411 1258
rect 1238 1253 1239 1257
rect 1243 1253 1244 1257
rect 1238 1252 1244 1253
rect 1280 1250 1282 1257
rect 1510 1256 1516 1257
rect 1510 1252 1511 1256
rect 1515 1252 1516 1256
rect 1510 1251 1516 1252
rect 1550 1256 1556 1257
rect 1550 1252 1551 1256
rect 1555 1252 1556 1256
rect 1550 1251 1556 1252
rect 1590 1256 1596 1257
rect 1590 1252 1591 1256
rect 1595 1252 1596 1256
rect 1590 1251 1596 1252
rect 1630 1256 1636 1257
rect 1630 1252 1631 1256
rect 1635 1252 1636 1256
rect 1630 1251 1636 1252
rect 1670 1256 1676 1257
rect 1670 1252 1671 1256
rect 1675 1252 1676 1256
rect 1670 1251 1676 1252
rect 1710 1256 1716 1257
rect 1710 1252 1711 1256
rect 1715 1252 1716 1256
rect 1710 1251 1716 1252
rect 1750 1256 1756 1257
rect 1750 1252 1751 1256
rect 1755 1252 1756 1256
rect 1750 1251 1756 1252
rect 1790 1256 1796 1257
rect 1790 1252 1791 1256
rect 1795 1252 1796 1256
rect 1790 1251 1796 1252
rect 1838 1256 1844 1257
rect 1838 1252 1839 1256
rect 1843 1252 1844 1256
rect 1838 1251 1844 1252
rect 1902 1256 1908 1257
rect 1902 1252 1903 1256
rect 1907 1252 1908 1256
rect 1902 1251 1908 1252
rect 1966 1256 1972 1257
rect 1966 1252 1967 1256
rect 1971 1252 1972 1256
rect 1966 1251 1972 1252
rect 2038 1256 2044 1257
rect 2038 1252 2039 1256
rect 2043 1252 2044 1256
rect 2038 1251 2044 1252
rect 2118 1256 2124 1257
rect 2118 1252 2119 1256
rect 2123 1252 2124 1256
rect 2118 1251 2124 1252
rect 2206 1256 2212 1257
rect 2206 1252 2207 1256
rect 2211 1252 2212 1256
rect 2206 1251 2212 1252
rect 2294 1256 2300 1257
rect 2294 1252 2295 1256
rect 2299 1252 2300 1256
rect 2294 1251 2300 1252
rect 2358 1256 2364 1257
rect 2358 1252 2359 1256
rect 2363 1252 2364 1256
rect 2358 1251 2364 1252
rect 2408 1250 2410 1257
rect 1278 1249 1284 1250
rect 1278 1245 1279 1249
rect 1283 1245 1284 1249
rect 1278 1244 1284 1245
rect 2406 1249 2412 1250
rect 2406 1245 2407 1249
rect 2411 1245 2412 1249
rect 2406 1244 2412 1245
rect 110 1240 116 1241
rect 110 1236 111 1240
rect 115 1236 116 1240
rect 110 1235 116 1236
rect 1238 1240 1244 1241
rect 1238 1236 1239 1240
rect 1243 1236 1244 1240
rect 1238 1235 1244 1236
rect 112 1195 114 1235
rect 134 1217 140 1218
rect 134 1213 135 1217
rect 139 1213 140 1217
rect 134 1212 140 1213
rect 174 1217 180 1218
rect 174 1213 175 1217
rect 179 1213 180 1217
rect 174 1212 180 1213
rect 246 1217 252 1218
rect 246 1213 247 1217
rect 251 1213 252 1217
rect 246 1212 252 1213
rect 326 1217 332 1218
rect 326 1213 327 1217
rect 331 1213 332 1217
rect 326 1212 332 1213
rect 414 1217 420 1218
rect 414 1213 415 1217
rect 419 1213 420 1217
rect 414 1212 420 1213
rect 502 1217 508 1218
rect 502 1213 503 1217
rect 507 1213 508 1217
rect 502 1212 508 1213
rect 590 1217 596 1218
rect 590 1213 591 1217
rect 595 1213 596 1217
rect 590 1212 596 1213
rect 670 1217 676 1218
rect 670 1213 671 1217
rect 675 1213 676 1217
rect 670 1212 676 1213
rect 742 1217 748 1218
rect 742 1213 743 1217
rect 747 1213 748 1217
rect 742 1212 748 1213
rect 814 1217 820 1218
rect 814 1213 815 1217
rect 819 1213 820 1217
rect 814 1212 820 1213
rect 878 1217 884 1218
rect 878 1213 879 1217
rect 883 1213 884 1217
rect 878 1212 884 1213
rect 942 1217 948 1218
rect 942 1213 943 1217
rect 947 1213 948 1217
rect 942 1212 948 1213
rect 1006 1217 1012 1218
rect 1006 1213 1007 1217
rect 1011 1213 1012 1217
rect 1006 1212 1012 1213
rect 1070 1217 1076 1218
rect 1070 1213 1071 1217
rect 1075 1213 1076 1217
rect 1070 1212 1076 1213
rect 136 1195 138 1212
rect 176 1195 178 1212
rect 248 1195 250 1212
rect 328 1195 330 1212
rect 416 1195 418 1212
rect 504 1195 506 1212
rect 592 1195 594 1212
rect 672 1195 674 1212
rect 744 1195 746 1212
rect 816 1195 818 1212
rect 880 1195 882 1212
rect 944 1195 946 1212
rect 1008 1195 1010 1212
rect 1072 1195 1074 1212
rect 1240 1195 1242 1235
rect 1278 1232 1284 1233
rect 1278 1228 1279 1232
rect 1283 1228 1284 1232
rect 1278 1227 1284 1228
rect 2406 1232 2412 1233
rect 2406 1228 2407 1232
rect 2411 1228 2412 1232
rect 2406 1227 2412 1228
rect 111 1194 115 1195
rect 111 1189 115 1190
rect 135 1194 139 1195
rect 135 1189 139 1190
rect 175 1194 179 1195
rect 175 1189 179 1190
rect 231 1194 235 1195
rect 231 1189 235 1190
rect 247 1194 251 1195
rect 247 1189 251 1190
rect 303 1194 307 1195
rect 303 1189 307 1190
rect 327 1194 331 1195
rect 327 1189 331 1190
rect 383 1194 387 1195
rect 383 1189 387 1190
rect 415 1194 419 1195
rect 415 1189 419 1190
rect 471 1194 475 1195
rect 471 1189 475 1190
rect 503 1194 507 1195
rect 503 1189 507 1190
rect 559 1194 563 1195
rect 559 1189 563 1190
rect 591 1194 595 1195
rect 591 1189 595 1190
rect 639 1194 643 1195
rect 639 1189 643 1190
rect 671 1194 675 1195
rect 671 1189 675 1190
rect 719 1194 723 1195
rect 719 1189 723 1190
rect 743 1194 747 1195
rect 743 1189 747 1190
rect 799 1194 803 1195
rect 799 1189 803 1190
rect 815 1194 819 1195
rect 815 1189 819 1190
rect 871 1194 875 1195
rect 871 1189 875 1190
rect 879 1194 883 1195
rect 879 1189 883 1190
rect 935 1194 939 1195
rect 935 1189 939 1190
rect 943 1194 947 1195
rect 943 1189 947 1190
rect 991 1194 995 1195
rect 991 1189 995 1190
rect 1007 1194 1011 1195
rect 1007 1189 1011 1190
rect 1047 1194 1051 1195
rect 1047 1189 1051 1190
rect 1071 1194 1075 1195
rect 1071 1189 1075 1190
rect 1103 1194 1107 1195
rect 1103 1189 1107 1190
rect 1151 1194 1155 1195
rect 1151 1189 1155 1190
rect 1191 1194 1195 1195
rect 1191 1189 1195 1190
rect 1239 1194 1243 1195
rect 1280 1191 1282 1227
rect 1510 1209 1516 1210
rect 1510 1205 1511 1209
rect 1515 1205 1516 1209
rect 1510 1204 1516 1205
rect 1550 1209 1556 1210
rect 1550 1205 1551 1209
rect 1555 1205 1556 1209
rect 1550 1204 1556 1205
rect 1590 1209 1596 1210
rect 1590 1205 1591 1209
rect 1595 1205 1596 1209
rect 1590 1204 1596 1205
rect 1630 1209 1636 1210
rect 1630 1205 1631 1209
rect 1635 1205 1636 1209
rect 1630 1204 1636 1205
rect 1670 1209 1676 1210
rect 1670 1205 1671 1209
rect 1675 1205 1676 1209
rect 1670 1204 1676 1205
rect 1710 1209 1716 1210
rect 1710 1205 1711 1209
rect 1715 1205 1716 1209
rect 1710 1204 1716 1205
rect 1750 1209 1756 1210
rect 1750 1205 1751 1209
rect 1755 1205 1756 1209
rect 1750 1204 1756 1205
rect 1790 1209 1796 1210
rect 1790 1205 1791 1209
rect 1795 1205 1796 1209
rect 1790 1204 1796 1205
rect 1838 1209 1844 1210
rect 1838 1205 1839 1209
rect 1843 1205 1844 1209
rect 1838 1204 1844 1205
rect 1902 1209 1908 1210
rect 1902 1205 1903 1209
rect 1907 1205 1908 1209
rect 1902 1204 1908 1205
rect 1966 1209 1972 1210
rect 1966 1205 1967 1209
rect 1971 1205 1972 1209
rect 1966 1204 1972 1205
rect 2038 1209 2044 1210
rect 2038 1205 2039 1209
rect 2043 1205 2044 1209
rect 2038 1204 2044 1205
rect 2118 1209 2124 1210
rect 2118 1205 2119 1209
rect 2123 1205 2124 1209
rect 2118 1204 2124 1205
rect 2206 1209 2212 1210
rect 2206 1205 2207 1209
rect 2211 1205 2212 1209
rect 2206 1204 2212 1205
rect 2294 1209 2300 1210
rect 2294 1205 2295 1209
rect 2299 1205 2300 1209
rect 2294 1204 2300 1205
rect 2358 1209 2364 1210
rect 2358 1205 2359 1209
rect 2363 1205 2364 1209
rect 2358 1204 2364 1205
rect 1512 1191 1514 1204
rect 1552 1191 1554 1204
rect 1592 1191 1594 1204
rect 1632 1191 1634 1204
rect 1672 1191 1674 1204
rect 1712 1191 1714 1204
rect 1752 1191 1754 1204
rect 1792 1191 1794 1204
rect 1840 1191 1842 1204
rect 1904 1191 1906 1204
rect 1968 1191 1970 1204
rect 2040 1191 2042 1204
rect 2120 1191 2122 1204
rect 2208 1191 2210 1204
rect 2296 1191 2298 1204
rect 2360 1191 2362 1204
rect 2408 1191 2410 1227
rect 1239 1189 1243 1190
rect 1279 1190 1283 1191
rect 112 1157 114 1189
rect 136 1180 138 1189
rect 176 1180 178 1189
rect 232 1180 234 1189
rect 304 1180 306 1189
rect 384 1180 386 1189
rect 472 1180 474 1189
rect 560 1180 562 1189
rect 640 1180 642 1189
rect 720 1180 722 1189
rect 800 1180 802 1189
rect 872 1180 874 1189
rect 936 1180 938 1189
rect 992 1180 994 1189
rect 1048 1180 1050 1189
rect 1104 1180 1106 1189
rect 1152 1180 1154 1189
rect 1192 1180 1194 1189
rect 134 1179 140 1180
rect 134 1175 135 1179
rect 139 1175 140 1179
rect 134 1174 140 1175
rect 174 1179 180 1180
rect 174 1175 175 1179
rect 179 1175 180 1179
rect 174 1174 180 1175
rect 230 1179 236 1180
rect 230 1175 231 1179
rect 235 1175 236 1179
rect 230 1174 236 1175
rect 302 1179 308 1180
rect 302 1175 303 1179
rect 307 1175 308 1179
rect 302 1174 308 1175
rect 382 1179 388 1180
rect 382 1175 383 1179
rect 387 1175 388 1179
rect 382 1174 388 1175
rect 470 1179 476 1180
rect 470 1175 471 1179
rect 475 1175 476 1179
rect 470 1174 476 1175
rect 558 1179 564 1180
rect 558 1175 559 1179
rect 563 1175 564 1179
rect 558 1174 564 1175
rect 638 1179 644 1180
rect 638 1175 639 1179
rect 643 1175 644 1179
rect 638 1174 644 1175
rect 718 1179 724 1180
rect 718 1175 719 1179
rect 723 1175 724 1179
rect 718 1174 724 1175
rect 798 1179 804 1180
rect 798 1175 799 1179
rect 803 1175 804 1179
rect 798 1174 804 1175
rect 870 1179 876 1180
rect 870 1175 871 1179
rect 875 1175 876 1179
rect 870 1174 876 1175
rect 934 1179 940 1180
rect 934 1175 935 1179
rect 939 1175 940 1179
rect 934 1174 940 1175
rect 990 1179 996 1180
rect 990 1175 991 1179
rect 995 1175 996 1179
rect 990 1174 996 1175
rect 1046 1179 1052 1180
rect 1046 1175 1047 1179
rect 1051 1175 1052 1179
rect 1046 1174 1052 1175
rect 1102 1179 1108 1180
rect 1102 1175 1103 1179
rect 1107 1175 1108 1179
rect 1102 1174 1108 1175
rect 1150 1179 1156 1180
rect 1150 1175 1151 1179
rect 1155 1175 1156 1179
rect 1150 1174 1156 1175
rect 1190 1179 1196 1180
rect 1190 1175 1191 1179
rect 1195 1175 1196 1179
rect 1190 1174 1196 1175
rect 1240 1157 1242 1189
rect 1279 1185 1283 1186
rect 1511 1190 1515 1191
rect 1511 1185 1515 1186
rect 1551 1190 1555 1191
rect 1551 1185 1555 1186
rect 1559 1190 1563 1191
rect 1559 1185 1563 1186
rect 1591 1190 1595 1191
rect 1591 1185 1595 1186
rect 1599 1190 1603 1191
rect 1599 1185 1603 1186
rect 1631 1190 1635 1191
rect 1631 1185 1635 1186
rect 1639 1190 1643 1191
rect 1639 1185 1643 1186
rect 1671 1190 1675 1191
rect 1671 1185 1675 1186
rect 1679 1190 1683 1191
rect 1679 1185 1683 1186
rect 1711 1190 1715 1191
rect 1711 1185 1715 1186
rect 1719 1190 1723 1191
rect 1719 1185 1723 1186
rect 1751 1190 1755 1191
rect 1751 1185 1755 1186
rect 1759 1190 1763 1191
rect 1759 1185 1763 1186
rect 1791 1190 1795 1191
rect 1791 1185 1795 1186
rect 1799 1190 1803 1191
rect 1799 1185 1803 1186
rect 1839 1190 1843 1191
rect 1839 1185 1843 1186
rect 1855 1190 1859 1191
rect 1855 1185 1859 1186
rect 1903 1190 1907 1191
rect 1903 1185 1907 1186
rect 1927 1190 1931 1191
rect 1927 1185 1931 1186
rect 1967 1190 1971 1191
rect 1967 1185 1971 1186
rect 2023 1190 2027 1191
rect 2023 1185 2027 1186
rect 2039 1190 2043 1191
rect 2039 1185 2043 1186
rect 2119 1190 2123 1191
rect 2119 1185 2123 1186
rect 2135 1190 2139 1191
rect 2135 1185 2139 1186
rect 2207 1190 2211 1191
rect 2207 1185 2211 1186
rect 2255 1190 2259 1191
rect 2255 1185 2259 1186
rect 2295 1190 2299 1191
rect 2295 1185 2299 1186
rect 2359 1190 2363 1191
rect 2359 1185 2363 1186
rect 2407 1190 2411 1191
rect 2407 1185 2411 1186
rect 110 1156 116 1157
rect 110 1152 111 1156
rect 115 1152 116 1156
rect 110 1151 116 1152
rect 1238 1156 1244 1157
rect 1238 1152 1239 1156
rect 1243 1152 1244 1156
rect 1280 1153 1282 1185
rect 1560 1176 1562 1185
rect 1600 1176 1602 1185
rect 1640 1176 1642 1185
rect 1680 1176 1682 1185
rect 1720 1176 1722 1185
rect 1760 1176 1762 1185
rect 1800 1176 1802 1185
rect 1856 1176 1858 1185
rect 1928 1176 1930 1185
rect 2024 1176 2026 1185
rect 2136 1176 2138 1185
rect 2256 1176 2258 1185
rect 2360 1176 2362 1185
rect 1558 1175 1564 1176
rect 1558 1171 1559 1175
rect 1563 1171 1564 1175
rect 1558 1170 1564 1171
rect 1598 1175 1604 1176
rect 1598 1171 1599 1175
rect 1603 1171 1604 1175
rect 1598 1170 1604 1171
rect 1638 1175 1644 1176
rect 1638 1171 1639 1175
rect 1643 1171 1644 1175
rect 1638 1170 1644 1171
rect 1678 1175 1684 1176
rect 1678 1171 1679 1175
rect 1683 1171 1684 1175
rect 1678 1170 1684 1171
rect 1718 1175 1724 1176
rect 1718 1171 1719 1175
rect 1723 1171 1724 1175
rect 1718 1170 1724 1171
rect 1758 1175 1764 1176
rect 1758 1171 1759 1175
rect 1763 1171 1764 1175
rect 1758 1170 1764 1171
rect 1798 1175 1804 1176
rect 1798 1171 1799 1175
rect 1803 1171 1804 1175
rect 1798 1170 1804 1171
rect 1854 1175 1860 1176
rect 1854 1171 1855 1175
rect 1859 1171 1860 1175
rect 1854 1170 1860 1171
rect 1926 1175 1932 1176
rect 1926 1171 1927 1175
rect 1931 1171 1932 1175
rect 1926 1170 1932 1171
rect 2022 1175 2028 1176
rect 2022 1171 2023 1175
rect 2027 1171 2028 1175
rect 2022 1170 2028 1171
rect 2134 1175 2140 1176
rect 2134 1171 2135 1175
rect 2139 1171 2140 1175
rect 2134 1170 2140 1171
rect 2254 1175 2260 1176
rect 2254 1171 2255 1175
rect 2259 1171 2260 1175
rect 2254 1170 2260 1171
rect 2358 1175 2364 1176
rect 2358 1171 2359 1175
rect 2363 1171 2364 1175
rect 2358 1170 2364 1171
rect 2408 1153 2410 1185
rect 1238 1151 1244 1152
rect 1278 1152 1284 1153
rect 1278 1148 1279 1152
rect 1283 1148 1284 1152
rect 1278 1147 1284 1148
rect 2406 1152 2412 1153
rect 2406 1148 2407 1152
rect 2411 1148 2412 1152
rect 2406 1147 2412 1148
rect 110 1139 116 1140
rect 110 1135 111 1139
rect 115 1135 116 1139
rect 110 1134 116 1135
rect 1238 1139 1244 1140
rect 1238 1135 1239 1139
rect 1243 1135 1244 1139
rect 1238 1134 1244 1135
rect 1278 1135 1284 1136
rect 112 1127 114 1134
rect 134 1132 140 1133
rect 134 1128 135 1132
rect 139 1128 140 1132
rect 134 1127 140 1128
rect 174 1132 180 1133
rect 174 1128 175 1132
rect 179 1128 180 1132
rect 174 1127 180 1128
rect 230 1132 236 1133
rect 230 1128 231 1132
rect 235 1128 236 1132
rect 230 1127 236 1128
rect 302 1132 308 1133
rect 302 1128 303 1132
rect 307 1128 308 1132
rect 302 1127 308 1128
rect 382 1132 388 1133
rect 382 1128 383 1132
rect 387 1128 388 1132
rect 382 1127 388 1128
rect 470 1132 476 1133
rect 470 1128 471 1132
rect 475 1128 476 1132
rect 470 1127 476 1128
rect 558 1132 564 1133
rect 558 1128 559 1132
rect 563 1128 564 1132
rect 558 1127 564 1128
rect 638 1132 644 1133
rect 638 1128 639 1132
rect 643 1128 644 1132
rect 638 1127 644 1128
rect 718 1132 724 1133
rect 718 1128 719 1132
rect 723 1128 724 1132
rect 718 1127 724 1128
rect 798 1132 804 1133
rect 798 1128 799 1132
rect 803 1128 804 1132
rect 798 1127 804 1128
rect 870 1132 876 1133
rect 870 1128 871 1132
rect 875 1128 876 1132
rect 870 1127 876 1128
rect 934 1132 940 1133
rect 934 1128 935 1132
rect 939 1128 940 1132
rect 934 1127 940 1128
rect 990 1132 996 1133
rect 990 1128 991 1132
rect 995 1128 996 1132
rect 990 1127 996 1128
rect 1046 1132 1052 1133
rect 1046 1128 1047 1132
rect 1051 1128 1052 1132
rect 1046 1127 1052 1128
rect 1102 1132 1108 1133
rect 1102 1128 1103 1132
rect 1107 1128 1108 1132
rect 1102 1127 1108 1128
rect 1150 1132 1156 1133
rect 1150 1128 1151 1132
rect 1155 1128 1156 1132
rect 1150 1127 1156 1128
rect 1190 1132 1196 1133
rect 1190 1128 1191 1132
rect 1195 1128 1196 1132
rect 1190 1127 1196 1128
rect 1240 1127 1242 1134
rect 1278 1131 1279 1135
rect 1283 1131 1284 1135
rect 1278 1130 1284 1131
rect 2406 1135 2412 1136
rect 2406 1131 2407 1135
rect 2411 1131 2412 1135
rect 2406 1130 2412 1131
rect 111 1126 115 1127
rect 111 1121 115 1122
rect 135 1126 139 1127
rect 135 1121 139 1122
rect 175 1126 179 1127
rect 175 1121 179 1122
rect 215 1126 219 1127
rect 215 1121 219 1122
rect 231 1126 235 1127
rect 231 1121 235 1122
rect 303 1126 307 1127
rect 303 1121 307 1122
rect 383 1126 387 1127
rect 383 1121 387 1122
rect 391 1126 395 1127
rect 391 1121 395 1122
rect 471 1126 475 1127
rect 471 1121 475 1122
rect 479 1126 483 1127
rect 479 1121 483 1122
rect 559 1126 563 1127
rect 559 1121 563 1122
rect 639 1126 643 1127
rect 639 1121 643 1122
rect 711 1126 715 1127
rect 711 1121 715 1122
rect 719 1126 723 1127
rect 719 1121 723 1122
rect 775 1126 779 1127
rect 775 1121 779 1122
rect 799 1126 803 1127
rect 799 1121 803 1122
rect 839 1126 843 1127
rect 839 1121 843 1122
rect 871 1126 875 1127
rect 871 1121 875 1122
rect 903 1126 907 1127
rect 903 1121 907 1122
rect 935 1126 939 1127
rect 935 1121 939 1122
rect 959 1126 963 1127
rect 959 1121 963 1122
rect 991 1126 995 1127
rect 991 1121 995 1122
rect 1023 1126 1027 1127
rect 1023 1121 1027 1122
rect 1047 1126 1051 1127
rect 1047 1121 1051 1122
rect 1087 1126 1091 1127
rect 1087 1121 1091 1122
rect 1103 1126 1107 1127
rect 1103 1121 1107 1122
rect 1151 1126 1155 1127
rect 1151 1121 1155 1122
rect 1191 1126 1195 1127
rect 1191 1121 1195 1122
rect 1239 1126 1243 1127
rect 1239 1121 1243 1122
rect 112 1114 114 1121
rect 134 1120 140 1121
rect 134 1116 135 1120
rect 139 1116 140 1120
rect 134 1115 140 1116
rect 214 1120 220 1121
rect 214 1116 215 1120
rect 219 1116 220 1120
rect 214 1115 220 1116
rect 302 1120 308 1121
rect 302 1116 303 1120
rect 307 1116 308 1120
rect 302 1115 308 1116
rect 390 1120 396 1121
rect 390 1116 391 1120
rect 395 1116 396 1120
rect 390 1115 396 1116
rect 478 1120 484 1121
rect 478 1116 479 1120
rect 483 1116 484 1120
rect 478 1115 484 1116
rect 558 1120 564 1121
rect 558 1116 559 1120
rect 563 1116 564 1120
rect 558 1115 564 1116
rect 638 1120 644 1121
rect 638 1116 639 1120
rect 643 1116 644 1120
rect 638 1115 644 1116
rect 710 1120 716 1121
rect 710 1116 711 1120
rect 715 1116 716 1120
rect 710 1115 716 1116
rect 774 1120 780 1121
rect 774 1116 775 1120
rect 779 1116 780 1120
rect 774 1115 780 1116
rect 838 1120 844 1121
rect 838 1116 839 1120
rect 843 1116 844 1120
rect 838 1115 844 1116
rect 902 1120 908 1121
rect 902 1116 903 1120
rect 907 1116 908 1120
rect 902 1115 908 1116
rect 958 1120 964 1121
rect 958 1116 959 1120
rect 963 1116 964 1120
rect 958 1115 964 1116
rect 1022 1120 1028 1121
rect 1022 1116 1023 1120
rect 1027 1116 1028 1120
rect 1022 1115 1028 1116
rect 1086 1120 1092 1121
rect 1086 1116 1087 1120
rect 1091 1116 1092 1120
rect 1086 1115 1092 1116
rect 1150 1120 1156 1121
rect 1150 1116 1151 1120
rect 1155 1116 1156 1120
rect 1150 1115 1156 1116
rect 1190 1120 1196 1121
rect 1190 1116 1191 1120
rect 1195 1116 1196 1120
rect 1190 1115 1196 1116
rect 1240 1114 1242 1121
rect 1280 1115 1282 1130
rect 1558 1128 1564 1129
rect 1558 1124 1559 1128
rect 1563 1124 1564 1128
rect 1558 1123 1564 1124
rect 1598 1128 1604 1129
rect 1598 1124 1599 1128
rect 1603 1124 1604 1128
rect 1598 1123 1604 1124
rect 1638 1128 1644 1129
rect 1638 1124 1639 1128
rect 1643 1124 1644 1128
rect 1638 1123 1644 1124
rect 1678 1128 1684 1129
rect 1678 1124 1679 1128
rect 1683 1124 1684 1128
rect 1678 1123 1684 1124
rect 1718 1128 1724 1129
rect 1718 1124 1719 1128
rect 1723 1124 1724 1128
rect 1718 1123 1724 1124
rect 1758 1128 1764 1129
rect 1758 1124 1759 1128
rect 1763 1124 1764 1128
rect 1758 1123 1764 1124
rect 1798 1128 1804 1129
rect 1798 1124 1799 1128
rect 1803 1124 1804 1128
rect 1798 1123 1804 1124
rect 1854 1128 1860 1129
rect 1854 1124 1855 1128
rect 1859 1124 1860 1128
rect 1854 1123 1860 1124
rect 1926 1128 1932 1129
rect 1926 1124 1927 1128
rect 1931 1124 1932 1128
rect 1926 1123 1932 1124
rect 2022 1128 2028 1129
rect 2022 1124 2023 1128
rect 2027 1124 2028 1128
rect 2022 1123 2028 1124
rect 2134 1128 2140 1129
rect 2134 1124 2135 1128
rect 2139 1124 2140 1128
rect 2134 1123 2140 1124
rect 2254 1128 2260 1129
rect 2254 1124 2255 1128
rect 2259 1124 2260 1128
rect 2254 1123 2260 1124
rect 2358 1128 2364 1129
rect 2358 1124 2359 1128
rect 2363 1124 2364 1128
rect 2358 1123 2364 1124
rect 1560 1115 1562 1123
rect 1600 1115 1602 1123
rect 1640 1115 1642 1123
rect 1680 1115 1682 1123
rect 1720 1115 1722 1123
rect 1760 1115 1762 1123
rect 1800 1115 1802 1123
rect 1856 1115 1858 1123
rect 1928 1115 1930 1123
rect 2024 1115 2026 1123
rect 2136 1115 2138 1123
rect 2256 1115 2258 1123
rect 2360 1115 2362 1123
rect 2408 1115 2410 1130
rect 1279 1114 1283 1115
rect 110 1113 116 1114
rect 110 1109 111 1113
rect 115 1109 116 1113
rect 110 1108 116 1109
rect 1238 1113 1244 1114
rect 1238 1109 1239 1113
rect 1243 1109 1244 1113
rect 1279 1109 1283 1110
rect 1535 1114 1539 1115
rect 1535 1109 1539 1110
rect 1559 1114 1563 1115
rect 1559 1109 1563 1110
rect 1599 1114 1603 1115
rect 1599 1109 1603 1110
rect 1639 1114 1643 1115
rect 1639 1109 1643 1110
rect 1663 1114 1667 1115
rect 1663 1109 1667 1110
rect 1679 1114 1683 1115
rect 1679 1109 1683 1110
rect 1719 1114 1723 1115
rect 1719 1109 1723 1110
rect 1727 1114 1731 1115
rect 1727 1109 1731 1110
rect 1759 1114 1763 1115
rect 1759 1109 1763 1110
rect 1791 1114 1795 1115
rect 1791 1109 1795 1110
rect 1799 1114 1803 1115
rect 1799 1109 1803 1110
rect 1855 1114 1859 1115
rect 1855 1109 1859 1110
rect 1911 1114 1915 1115
rect 1911 1109 1915 1110
rect 1927 1114 1931 1115
rect 1927 1109 1931 1110
rect 1967 1114 1971 1115
rect 1967 1109 1971 1110
rect 2023 1114 2027 1115
rect 2023 1109 2027 1110
rect 2079 1114 2083 1115
rect 2079 1109 2083 1110
rect 2135 1114 2139 1115
rect 2135 1109 2139 1110
rect 2191 1114 2195 1115
rect 2191 1109 2195 1110
rect 2255 1114 2259 1115
rect 2255 1109 2259 1110
rect 2319 1114 2323 1115
rect 2319 1109 2323 1110
rect 2359 1114 2363 1115
rect 2359 1109 2363 1110
rect 2407 1114 2411 1115
rect 2407 1109 2411 1110
rect 1238 1108 1244 1109
rect 1280 1102 1282 1109
rect 1534 1108 1540 1109
rect 1534 1104 1535 1108
rect 1539 1104 1540 1108
rect 1534 1103 1540 1104
rect 1598 1108 1604 1109
rect 1598 1104 1599 1108
rect 1603 1104 1604 1108
rect 1598 1103 1604 1104
rect 1662 1108 1668 1109
rect 1662 1104 1663 1108
rect 1667 1104 1668 1108
rect 1662 1103 1668 1104
rect 1726 1108 1732 1109
rect 1726 1104 1727 1108
rect 1731 1104 1732 1108
rect 1726 1103 1732 1104
rect 1790 1108 1796 1109
rect 1790 1104 1791 1108
rect 1795 1104 1796 1108
rect 1790 1103 1796 1104
rect 1854 1108 1860 1109
rect 1854 1104 1855 1108
rect 1859 1104 1860 1108
rect 1854 1103 1860 1104
rect 1910 1108 1916 1109
rect 1910 1104 1911 1108
rect 1915 1104 1916 1108
rect 1910 1103 1916 1104
rect 1966 1108 1972 1109
rect 1966 1104 1967 1108
rect 1971 1104 1972 1108
rect 1966 1103 1972 1104
rect 2022 1108 2028 1109
rect 2022 1104 2023 1108
rect 2027 1104 2028 1108
rect 2022 1103 2028 1104
rect 2078 1108 2084 1109
rect 2078 1104 2079 1108
rect 2083 1104 2084 1108
rect 2078 1103 2084 1104
rect 2134 1108 2140 1109
rect 2134 1104 2135 1108
rect 2139 1104 2140 1108
rect 2134 1103 2140 1104
rect 2190 1108 2196 1109
rect 2190 1104 2191 1108
rect 2195 1104 2196 1108
rect 2190 1103 2196 1104
rect 2254 1108 2260 1109
rect 2254 1104 2255 1108
rect 2259 1104 2260 1108
rect 2254 1103 2260 1104
rect 2318 1108 2324 1109
rect 2318 1104 2319 1108
rect 2323 1104 2324 1108
rect 2318 1103 2324 1104
rect 2358 1108 2364 1109
rect 2358 1104 2359 1108
rect 2363 1104 2364 1108
rect 2358 1103 2364 1104
rect 2408 1102 2410 1109
rect 1278 1101 1284 1102
rect 1278 1097 1279 1101
rect 1283 1097 1284 1101
rect 110 1096 116 1097
rect 110 1092 111 1096
rect 115 1092 116 1096
rect 110 1091 116 1092
rect 1238 1096 1244 1097
rect 1278 1096 1284 1097
rect 2406 1101 2412 1102
rect 2406 1097 2407 1101
rect 2411 1097 2412 1101
rect 2406 1096 2412 1097
rect 1238 1092 1239 1096
rect 1243 1092 1244 1096
rect 1238 1091 1244 1092
rect 112 1055 114 1091
rect 134 1073 140 1074
rect 134 1069 135 1073
rect 139 1069 140 1073
rect 134 1068 140 1069
rect 214 1073 220 1074
rect 214 1069 215 1073
rect 219 1069 220 1073
rect 214 1068 220 1069
rect 302 1073 308 1074
rect 302 1069 303 1073
rect 307 1069 308 1073
rect 302 1068 308 1069
rect 390 1073 396 1074
rect 390 1069 391 1073
rect 395 1069 396 1073
rect 390 1068 396 1069
rect 478 1073 484 1074
rect 478 1069 479 1073
rect 483 1069 484 1073
rect 478 1068 484 1069
rect 558 1073 564 1074
rect 558 1069 559 1073
rect 563 1069 564 1073
rect 558 1068 564 1069
rect 638 1073 644 1074
rect 638 1069 639 1073
rect 643 1069 644 1073
rect 638 1068 644 1069
rect 710 1073 716 1074
rect 710 1069 711 1073
rect 715 1069 716 1073
rect 710 1068 716 1069
rect 774 1073 780 1074
rect 774 1069 775 1073
rect 779 1069 780 1073
rect 774 1068 780 1069
rect 838 1073 844 1074
rect 838 1069 839 1073
rect 843 1069 844 1073
rect 838 1068 844 1069
rect 902 1073 908 1074
rect 902 1069 903 1073
rect 907 1069 908 1073
rect 902 1068 908 1069
rect 958 1073 964 1074
rect 958 1069 959 1073
rect 963 1069 964 1073
rect 958 1068 964 1069
rect 1022 1073 1028 1074
rect 1022 1069 1023 1073
rect 1027 1069 1028 1073
rect 1022 1068 1028 1069
rect 1086 1073 1092 1074
rect 1086 1069 1087 1073
rect 1091 1069 1092 1073
rect 1086 1068 1092 1069
rect 1150 1073 1156 1074
rect 1150 1069 1151 1073
rect 1155 1069 1156 1073
rect 1150 1068 1156 1069
rect 1190 1073 1196 1074
rect 1190 1069 1191 1073
rect 1195 1069 1196 1073
rect 1190 1068 1196 1069
rect 136 1055 138 1068
rect 216 1055 218 1068
rect 304 1055 306 1068
rect 392 1055 394 1068
rect 480 1055 482 1068
rect 560 1055 562 1068
rect 640 1055 642 1068
rect 712 1055 714 1068
rect 776 1055 778 1068
rect 840 1055 842 1068
rect 904 1055 906 1068
rect 960 1055 962 1068
rect 1024 1055 1026 1068
rect 1088 1055 1090 1068
rect 1152 1055 1154 1068
rect 1192 1055 1194 1068
rect 1240 1055 1242 1091
rect 1278 1084 1284 1085
rect 1278 1080 1279 1084
rect 1283 1080 1284 1084
rect 1278 1079 1284 1080
rect 2406 1084 2412 1085
rect 2406 1080 2407 1084
rect 2411 1080 2412 1084
rect 2406 1079 2412 1080
rect 111 1054 115 1055
rect 111 1049 115 1050
rect 135 1054 139 1055
rect 135 1049 139 1050
rect 199 1054 203 1055
rect 199 1049 203 1050
rect 215 1054 219 1055
rect 215 1049 219 1050
rect 239 1054 243 1055
rect 239 1049 243 1050
rect 287 1054 291 1055
rect 287 1049 291 1050
rect 303 1054 307 1055
rect 303 1049 307 1050
rect 343 1054 347 1055
rect 343 1049 347 1050
rect 391 1054 395 1055
rect 391 1049 395 1050
rect 439 1054 443 1055
rect 439 1049 443 1050
rect 479 1054 483 1055
rect 479 1049 483 1050
rect 487 1054 491 1055
rect 487 1049 491 1050
rect 535 1054 539 1055
rect 535 1049 539 1050
rect 559 1054 563 1055
rect 559 1049 563 1050
rect 583 1054 587 1055
rect 583 1049 587 1050
rect 631 1054 635 1055
rect 631 1049 635 1050
rect 639 1054 643 1055
rect 639 1049 643 1050
rect 679 1054 683 1055
rect 679 1049 683 1050
rect 711 1054 715 1055
rect 711 1049 715 1050
rect 727 1054 731 1055
rect 727 1049 731 1050
rect 775 1054 779 1055
rect 775 1049 779 1050
rect 783 1054 787 1055
rect 783 1049 787 1050
rect 839 1054 843 1055
rect 839 1049 843 1050
rect 895 1054 899 1055
rect 895 1049 899 1050
rect 903 1054 907 1055
rect 903 1049 907 1050
rect 959 1054 963 1055
rect 959 1049 963 1050
rect 1023 1054 1027 1055
rect 1023 1049 1027 1050
rect 1087 1054 1091 1055
rect 1087 1049 1091 1050
rect 1151 1054 1155 1055
rect 1151 1049 1155 1050
rect 1191 1054 1195 1055
rect 1191 1049 1195 1050
rect 1239 1054 1243 1055
rect 1239 1049 1243 1050
rect 112 1017 114 1049
rect 200 1040 202 1049
rect 240 1040 242 1049
rect 288 1040 290 1049
rect 344 1040 346 1049
rect 392 1040 394 1049
rect 440 1040 442 1049
rect 488 1040 490 1049
rect 536 1040 538 1049
rect 584 1040 586 1049
rect 632 1040 634 1049
rect 680 1040 682 1049
rect 728 1040 730 1049
rect 784 1040 786 1049
rect 840 1040 842 1049
rect 896 1040 898 1049
rect 960 1040 962 1049
rect 1024 1040 1026 1049
rect 1088 1040 1090 1049
rect 1152 1040 1154 1049
rect 1192 1040 1194 1049
rect 198 1039 204 1040
rect 198 1035 199 1039
rect 203 1035 204 1039
rect 198 1034 204 1035
rect 238 1039 244 1040
rect 238 1035 239 1039
rect 243 1035 244 1039
rect 238 1034 244 1035
rect 286 1039 292 1040
rect 286 1035 287 1039
rect 291 1035 292 1039
rect 286 1034 292 1035
rect 342 1039 348 1040
rect 342 1035 343 1039
rect 347 1035 348 1039
rect 342 1034 348 1035
rect 390 1039 396 1040
rect 390 1035 391 1039
rect 395 1035 396 1039
rect 390 1034 396 1035
rect 438 1039 444 1040
rect 438 1035 439 1039
rect 443 1035 444 1039
rect 438 1034 444 1035
rect 486 1039 492 1040
rect 486 1035 487 1039
rect 491 1035 492 1039
rect 486 1034 492 1035
rect 534 1039 540 1040
rect 534 1035 535 1039
rect 539 1035 540 1039
rect 534 1034 540 1035
rect 582 1039 588 1040
rect 582 1035 583 1039
rect 587 1035 588 1039
rect 582 1034 588 1035
rect 630 1039 636 1040
rect 630 1035 631 1039
rect 635 1035 636 1039
rect 630 1034 636 1035
rect 678 1039 684 1040
rect 678 1035 679 1039
rect 683 1035 684 1039
rect 678 1034 684 1035
rect 726 1039 732 1040
rect 726 1035 727 1039
rect 731 1035 732 1039
rect 726 1034 732 1035
rect 782 1039 788 1040
rect 782 1035 783 1039
rect 787 1035 788 1039
rect 782 1034 788 1035
rect 838 1039 844 1040
rect 838 1035 839 1039
rect 843 1035 844 1039
rect 838 1034 844 1035
rect 894 1039 900 1040
rect 894 1035 895 1039
rect 899 1035 900 1039
rect 894 1034 900 1035
rect 958 1039 964 1040
rect 958 1035 959 1039
rect 963 1035 964 1039
rect 958 1034 964 1035
rect 1022 1039 1028 1040
rect 1022 1035 1023 1039
rect 1027 1035 1028 1039
rect 1022 1034 1028 1035
rect 1086 1039 1092 1040
rect 1086 1035 1087 1039
rect 1091 1035 1092 1039
rect 1086 1034 1092 1035
rect 1150 1039 1156 1040
rect 1150 1035 1151 1039
rect 1155 1035 1156 1039
rect 1150 1034 1156 1035
rect 1190 1039 1196 1040
rect 1190 1035 1191 1039
rect 1195 1035 1196 1039
rect 1190 1034 1196 1035
rect 1240 1017 1242 1049
rect 1280 1035 1282 1079
rect 1534 1061 1540 1062
rect 1534 1057 1535 1061
rect 1539 1057 1540 1061
rect 1534 1056 1540 1057
rect 1598 1061 1604 1062
rect 1598 1057 1599 1061
rect 1603 1057 1604 1061
rect 1598 1056 1604 1057
rect 1662 1061 1668 1062
rect 1662 1057 1663 1061
rect 1667 1057 1668 1061
rect 1662 1056 1668 1057
rect 1726 1061 1732 1062
rect 1726 1057 1727 1061
rect 1731 1057 1732 1061
rect 1726 1056 1732 1057
rect 1790 1061 1796 1062
rect 1790 1057 1791 1061
rect 1795 1057 1796 1061
rect 1790 1056 1796 1057
rect 1854 1061 1860 1062
rect 1854 1057 1855 1061
rect 1859 1057 1860 1061
rect 1854 1056 1860 1057
rect 1910 1061 1916 1062
rect 1910 1057 1911 1061
rect 1915 1057 1916 1061
rect 1910 1056 1916 1057
rect 1966 1061 1972 1062
rect 1966 1057 1967 1061
rect 1971 1057 1972 1061
rect 1966 1056 1972 1057
rect 2022 1061 2028 1062
rect 2022 1057 2023 1061
rect 2027 1057 2028 1061
rect 2022 1056 2028 1057
rect 2078 1061 2084 1062
rect 2078 1057 2079 1061
rect 2083 1057 2084 1061
rect 2078 1056 2084 1057
rect 2134 1061 2140 1062
rect 2134 1057 2135 1061
rect 2139 1057 2140 1061
rect 2134 1056 2140 1057
rect 2190 1061 2196 1062
rect 2190 1057 2191 1061
rect 2195 1057 2196 1061
rect 2190 1056 2196 1057
rect 2254 1061 2260 1062
rect 2254 1057 2255 1061
rect 2259 1057 2260 1061
rect 2254 1056 2260 1057
rect 2318 1061 2324 1062
rect 2318 1057 2319 1061
rect 2323 1057 2324 1061
rect 2318 1056 2324 1057
rect 2358 1061 2364 1062
rect 2358 1057 2359 1061
rect 2363 1057 2364 1061
rect 2358 1056 2364 1057
rect 1536 1035 1538 1056
rect 1600 1035 1602 1056
rect 1664 1035 1666 1056
rect 1728 1035 1730 1056
rect 1792 1035 1794 1056
rect 1856 1035 1858 1056
rect 1912 1035 1914 1056
rect 1968 1035 1970 1056
rect 2024 1035 2026 1056
rect 2080 1035 2082 1056
rect 2136 1035 2138 1056
rect 2192 1035 2194 1056
rect 2256 1035 2258 1056
rect 2320 1035 2322 1056
rect 2360 1035 2362 1056
rect 2408 1035 2410 1079
rect 1279 1034 1283 1035
rect 1279 1029 1283 1030
rect 1503 1034 1507 1035
rect 1503 1029 1507 1030
rect 1535 1034 1539 1035
rect 1535 1029 1539 1030
rect 1599 1034 1603 1035
rect 1599 1029 1603 1030
rect 1623 1034 1627 1035
rect 1623 1029 1627 1030
rect 1663 1034 1667 1035
rect 1663 1029 1667 1030
rect 1727 1034 1731 1035
rect 1727 1029 1731 1030
rect 1735 1034 1739 1035
rect 1735 1029 1739 1030
rect 1791 1034 1795 1035
rect 1791 1029 1795 1030
rect 1831 1034 1835 1035
rect 1831 1029 1835 1030
rect 1855 1034 1859 1035
rect 1855 1029 1859 1030
rect 1911 1034 1915 1035
rect 1911 1029 1915 1030
rect 1919 1034 1923 1035
rect 1919 1029 1923 1030
rect 1967 1034 1971 1035
rect 1967 1029 1971 1030
rect 1999 1034 2003 1035
rect 1999 1029 2003 1030
rect 2023 1034 2027 1035
rect 2023 1029 2027 1030
rect 2071 1034 2075 1035
rect 2071 1029 2075 1030
rect 2079 1034 2083 1035
rect 2079 1029 2083 1030
rect 2135 1034 2139 1035
rect 2135 1029 2139 1030
rect 2143 1034 2147 1035
rect 2143 1029 2147 1030
rect 2191 1034 2195 1035
rect 2191 1029 2195 1030
rect 2207 1034 2211 1035
rect 2207 1029 2211 1030
rect 2255 1034 2259 1035
rect 2255 1029 2259 1030
rect 2279 1034 2283 1035
rect 2279 1029 2283 1030
rect 2319 1034 2323 1035
rect 2319 1029 2323 1030
rect 2359 1034 2363 1035
rect 2359 1029 2363 1030
rect 2407 1034 2411 1035
rect 2407 1029 2411 1030
rect 110 1016 116 1017
rect 110 1012 111 1016
rect 115 1012 116 1016
rect 110 1011 116 1012
rect 1238 1016 1244 1017
rect 1238 1012 1239 1016
rect 1243 1012 1244 1016
rect 1238 1011 1244 1012
rect 110 999 116 1000
rect 110 995 111 999
rect 115 995 116 999
rect 110 994 116 995
rect 1238 999 1244 1000
rect 1238 995 1239 999
rect 1243 995 1244 999
rect 1280 997 1282 1029
rect 1504 1020 1506 1029
rect 1624 1020 1626 1029
rect 1736 1020 1738 1029
rect 1832 1020 1834 1029
rect 1920 1020 1922 1029
rect 2000 1020 2002 1029
rect 2072 1020 2074 1029
rect 2144 1020 2146 1029
rect 2208 1020 2210 1029
rect 2280 1020 2282 1029
rect 1502 1019 1508 1020
rect 1502 1015 1503 1019
rect 1507 1015 1508 1019
rect 1502 1014 1508 1015
rect 1622 1019 1628 1020
rect 1622 1015 1623 1019
rect 1627 1015 1628 1019
rect 1622 1014 1628 1015
rect 1734 1019 1740 1020
rect 1734 1015 1735 1019
rect 1739 1015 1740 1019
rect 1734 1014 1740 1015
rect 1830 1019 1836 1020
rect 1830 1015 1831 1019
rect 1835 1015 1836 1019
rect 1830 1014 1836 1015
rect 1918 1019 1924 1020
rect 1918 1015 1919 1019
rect 1923 1015 1924 1019
rect 1918 1014 1924 1015
rect 1998 1019 2004 1020
rect 1998 1015 1999 1019
rect 2003 1015 2004 1019
rect 1998 1014 2004 1015
rect 2070 1019 2076 1020
rect 2070 1015 2071 1019
rect 2075 1015 2076 1019
rect 2070 1014 2076 1015
rect 2142 1019 2148 1020
rect 2142 1015 2143 1019
rect 2147 1015 2148 1019
rect 2142 1014 2148 1015
rect 2206 1019 2212 1020
rect 2206 1015 2207 1019
rect 2211 1015 2212 1019
rect 2206 1014 2212 1015
rect 2278 1019 2284 1020
rect 2278 1015 2279 1019
rect 2283 1015 2284 1019
rect 2278 1014 2284 1015
rect 2408 997 2410 1029
rect 1238 994 1244 995
rect 1278 996 1284 997
rect 112 975 114 994
rect 198 992 204 993
rect 198 988 199 992
rect 203 988 204 992
rect 198 987 204 988
rect 238 992 244 993
rect 238 988 239 992
rect 243 988 244 992
rect 238 987 244 988
rect 286 992 292 993
rect 286 988 287 992
rect 291 988 292 992
rect 286 987 292 988
rect 342 992 348 993
rect 342 988 343 992
rect 347 988 348 992
rect 342 987 348 988
rect 390 992 396 993
rect 390 988 391 992
rect 395 988 396 992
rect 390 987 396 988
rect 438 992 444 993
rect 438 988 439 992
rect 443 988 444 992
rect 438 987 444 988
rect 486 992 492 993
rect 486 988 487 992
rect 491 988 492 992
rect 486 987 492 988
rect 534 992 540 993
rect 534 988 535 992
rect 539 988 540 992
rect 534 987 540 988
rect 582 992 588 993
rect 582 988 583 992
rect 587 988 588 992
rect 582 987 588 988
rect 630 992 636 993
rect 630 988 631 992
rect 635 988 636 992
rect 630 987 636 988
rect 678 992 684 993
rect 678 988 679 992
rect 683 988 684 992
rect 678 987 684 988
rect 726 992 732 993
rect 726 988 727 992
rect 731 988 732 992
rect 726 987 732 988
rect 782 992 788 993
rect 782 988 783 992
rect 787 988 788 992
rect 782 987 788 988
rect 838 992 844 993
rect 838 988 839 992
rect 843 988 844 992
rect 838 987 844 988
rect 894 992 900 993
rect 894 988 895 992
rect 899 988 900 992
rect 894 987 900 988
rect 958 992 964 993
rect 958 988 959 992
rect 963 988 964 992
rect 958 987 964 988
rect 1022 992 1028 993
rect 1022 988 1023 992
rect 1027 988 1028 992
rect 1022 987 1028 988
rect 1086 992 1092 993
rect 1086 988 1087 992
rect 1091 988 1092 992
rect 1086 987 1092 988
rect 1150 992 1156 993
rect 1150 988 1151 992
rect 1155 988 1156 992
rect 1150 987 1156 988
rect 1190 992 1196 993
rect 1190 988 1191 992
rect 1195 988 1196 992
rect 1190 987 1196 988
rect 200 975 202 987
rect 240 975 242 987
rect 288 975 290 987
rect 344 975 346 987
rect 392 975 394 987
rect 440 975 442 987
rect 488 975 490 987
rect 536 975 538 987
rect 584 975 586 987
rect 632 975 634 987
rect 680 975 682 987
rect 728 975 730 987
rect 784 975 786 987
rect 840 975 842 987
rect 896 975 898 987
rect 960 975 962 987
rect 1024 975 1026 987
rect 1088 975 1090 987
rect 1152 975 1154 987
rect 1192 975 1194 987
rect 1240 975 1242 994
rect 1278 992 1279 996
rect 1283 992 1284 996
rect 1278 991 1284 992
rect 2406 996 2412 997
rect 2406 992 2407 996
rect 2411 992 2412 996
rect 2406 991 2412 992
rect 1278 979 1284 980
rect 1278 975 1279 979
rect 1283 975 1284 979
rect 111 974 115 975
rect 111 969 115 970
rect 199 974 203 975
rect 199 969 203 970
rect 239 974 243 975
rect 239 969 243 970
rect 287 974 291 975
rect 287 969 291 970
rect 295 974 299 975
rect 295 969 299 970
rect 343 974 347 975
rect 343 969 347 970
rect 391 974 395 975
rect 391 969 395 970
rect 399 974 403 975
rect 399 969 403 970
rect 439 974 443 975
rect 439 969 443 970
rect 471 974 475 975
rect 471 969 475 970
rect 487 974 491 975
rect 487 969 491 970
rect 535 974 539 975
rect 535 969 539 970
rect 551 974 555 975
rect 551 969 555 970
rect 583 974 587 975
rect 583 969 587 970
rect 631 974 635 975
rect 631 969 635 970
rect 639 974 643 975
rect 639 969 643 970
rect 679 974 683 975
rect 679 969 683 970
rect 727 974 731 975
rect 727 969 731 970
rect 783 974 787 975
rect 783 969 787 970
rect 807 974 811 975
rect 807 969 811 970
rect 839 974 843 975
rect 839 969 843 970
rect 887 974 891 975
rect 887 969 891 970
rect 895 974 899 975
rect 895 969 899 970
rect 959 974 963 975
rect 959 969 963 970
rect 1023 974 1027 975
rect 1023 969 1027 970
rect 1087 974 1091 975
rect 1087 969 1091 970
rect 1151 974 1155 975
rect 1151 969 1155 970
rect 1191 974 1195 975
rect 1191 969 1195 970
rect 1239 974 1243 975
rect 1278 974 1284 975
rect 2406 979 2412 980
rect 2406 975 2407 979
rect 2411 975 2412 979
rect 2406 974 2412 975
rect 1239 969 1243 970
rect 112 962 114 969
rect 294 968 300 969
rect 294 964 295 968
rect 299 964 300 968
rect 294 963 300 964
rect 342 968 348 969
rect 342 964 343 968
rect 347 964 348 968
rect 342 963 348 964
rect 398 968 404 969
rect 398 964 399 968
rect 403 964 404 968
rect 398 963 404 964
rect 470 968 476 969
rect 470 964 471 968
rect 475 964 476 968
rect 470 963 476 964
rect 550 968 556 969
rect 550 964 551 968
rect 555 964 556 968
rect 550 963 556 964
rect 638 968 644 969
rect 638 964 639 968
rect 643 964 644 968
rect 638 963 644 964
rect 726 968 732 969
rect 726 964 727 968
rect 731 964 732 968
rect 726 963 732 964
rect 806 968 812 969
rect 806 964 807 968
rect 811 964 812 968
rect 806 963 812 964
rect 886 968 892 969
rect 886 964 887 968
rect 891 964 892 968
rect 886 963 892 964
rect 958 968 964 969
rect 958 964 959 968
rect 963 964 964 968
rect 958 963 964 964
rect 1022 968 1028 969
rect 1022 964 1023 968
rect 1027 964 1028 968
rect 1022 963 1028 964
rect 1086 968 1092 969
rect 1086 964 1087 968
rect 1091 964 1092 968
rect 1086 963 1092 964
rect 1150 968 1156 969
rect 1150 964 1151 968
rect 1155 964 1156 968
rect 1150 963 1156 964
rect 1190 968 1196 969
rect 1190 964 1191 968
rect 1195 964 1196 968
rect 1190 963 1196 964
rect 1240 962 1242 969
rect 110 961 116 962
rect 110 957 111 961
rect 115 957 116 961
rect 110 956 116 957
rect 1238 961 1244 962
rect 1238 957 1239 961
rect 1243 957 1244 961
rect 1280 959 1282 974
rect 1502 972 1508 973
rect 1502 968 1503 972
rect 1507 968 1508 972
rect 1502 967 1508 968
rect 1622 972 1628 973
rect 1622 968 1623 972
rect 1627 968 1628 972
rect 1622 967 1628 968
rect 1734 972 1740 973
rect 1734 968 1735 972
rect 1739 968 1740 972
rect 1734 967 1740 968
rect 1830 972 1836 973
rect 1830 968 1831 972
rect 1835 968 1836 972
rect 1830 967 1836 968
rect 1918 972 1924 973
rect 1918 968 1919 972
rect 1923 968 1924 972
rect 1918 967 1924 968
rect 1998 972 2004 973
rect 1998 968 1999 972
rect 2003 968 2004 972
rect 1998 967 2004 968
rect 2070 972 2076 973
rect 2070 968 2071 972
rect 2075 968 2076 972
rect 2070 967 2076 968
rect 2142 972 2148 973
rect 2142 968 2143 972
rect 2147 968 2148 972
rect 2142 967 2148 968
rect 2206 972 2212 973
rect 2206 968 2207 972
rect 2211 968 2212 972
rect 2206 967 2212 968
rect 2278 972 2284 973
rect 2278 968 2279 972
rect 2283 968 2284 972
rect 2278 967 2284 968
rect 1504 959 1506 967
rect 1624 959 1626 967
rect 1736 959 1738 967
rect 1832 959 1834 967
rect 1920 959 1922 967
rect 2000 959 2002 967
rect 2072 959 2074 967
rect 2144 959 2146 967
rect 2208 959 2210 967
rect 2280 959 2282 967
rect 2408 959 2410 974
rect 1238 956 1244 957
rect 1279 958 1283 959
rect 1279 953 1283 954
rect 1319 958 1323 959
rect 1319 953 1323 954
rect 1359 958 1363 959
rect 1359 953 1363 954
rect 1399 958 1403 959
rect 1399 953 1403 954
rect 1463 958 1467 959
rect 1463 953 1467 954
rect 1503 958 1507 959
rect 1503 953 1507 954
rect 1543 958 1547 959
rect 1543 953 1547 954
rect 1623 958 1627 959
rect 1623 953 1627 954
rect 1639 958 1643 959
rect 1639 953 1643 954
rect 1735 958 1739 959
rect 1735 953 1739 954
rect 1831 958 1835 959
rect 1831 953 1835 954
rect 1839 958 1843 959
rect 1839 953 1843 954
rect 1919 958 1923 959
rect 1919 953 1923 954
rect 1935 958 1939 959
rect 1935 953 1939 954
rect 1999 958 2003 959
rect 1999 953 2003 954
rect 2023 958 2027 959
rect 2023 953 2027 954
rect 2071 958 2075 959
rect 2071 953 2075 954
rect 2103 958 2107 959
rect 2103 953 2107 954
rect 2143 958 2147 959
rect 2143 953 2147 954
rect 2175 958 2179 959
rect 2175 953 2179 954
rect 2207 958 2211 959
rect 2207 953 2211 954
rect 2239 958 2243 959
rect 2239 953 2243 954
rect 2279 958 2283 959
rect 2279 953 2283 954
rect 2311 958 2315 959
rect 2311 953 2315 954
rect 2359 958 2363 959
rect 2359 953 2363 954
rect 2407 958 2411 959
rect 2407 953 2411 954
rect 1280 946 1282 953
rect 1318 952 1324 953
rect 1318 948 1319 952
rect 1323 948 1324 952
rect 1318 947 1324 948
rect 1358 952 1364 953
rect 1358 948 1359 952
rect 1363 948 1364 952
rect 1358 947 1364 948
rect 1398 952 1404 953
rect 1398 948 1399 952
rect 1403 948 1404 952
rect 1398 947 1404 948
rect 1462 952 1468 953
rect 1462 948 1463 952
rect 1467 948 1468 952
rect 1462 947 1468 948
rect 1542 952 1548 953
rect 1542 948 1543 952
rect 1547 948 1548 952
rect 1542 947 1548 948
rect 1638 952 1644 953
rect 1638 948 1639 952
rect 1643 948 1644 952
rect 1638 947 1644 948
rect 1734 952 1740 953
rect 1734 948 1735 952
rect 1739 948 1740 952
rect 1734 947 1740 948
rect 1838 952 1844 953
rect 1838 948 1839 952
rect 1843 948 1844 952
rect 1838 947 1844 948
rect 1934 952 1940 953
rect 1934 948 1935 952
rect 1939 948 1940 952
rect 1934 947 1940 948
rect 2022 952 2028 953
rect 2022 948 2023 952
rect 2027 948 2028 952
rect 2022 947 2028 948
rect 2102 952 2108 953
rect 2102 948 2103 952
rect 2107 948 2108 952
rect 2102 947 2108 948
rect 2174 952 2180 953
rect 2174 948 2175 952
rect 2179 948 2180 952
rect 2174 947 2180 948
rect 2238 952 2244 953
rect 2238 948 2239 952
rect 2243 948 2244 952
rect 2238 947 2244 948
rect 2310 952 2316 953
rect 2310 948 2311 952
rect 2315 948 2316 952
rect 2310 947 2316 948
rect 2358 952 2364 953
rect 2358 948 2359 952
rect 2363 948 2364 952
rect 2358 947 2364 948
rect 2408 946 2410 953
rect 1278 945 1284 946
rect 110 944 116 945
rect 110 940 111 944
rect 115 940 116 944
rect 110 939 116 940
rect 1238 944 1244 945
rect 1238 940 1239 944
rect 1243 940 1244 944
rect 1278 941 1279 945
rect 1283 941 1284 945
rect 1278 940 1284 941
rect 2406 945 2412 946
rect 2406 941 2407 945
rect 2411 941 2412 945
rect 2406 940 2412 941
rect 1238 939 1244 940
rect 112 899 114 939
rect 294 921 300 922
rect 294 917 295 921
rect 299 917 300 921
rect 294 916 300 917
rect 342 921 348 922
rect 342 917 343 921
rect 347 917 348 921
rect 342 916 348 917
rect 398 921 404 922
rect 398 917 399 921
rect 403 917 404 921
rect 398 916 404 917
rect 470 921 476 922
rect 470 917 471 921
rect 475 917 476 921
rect 470 916 476 917
rect 550 921 556 922
rect 550 917 551 921
rect 555 917 556 921
rect 550 916 556 917
rect 638 921 644 922
rect 638 917 639 921
rect 643 917 644 921
rect 638 916 644 917
rect 726 921 732 922
rect 726 917 727 921
rect 731 917 732 921
rect 726 916 732 917
rect 806 921 812 922
rect 806 917 807 921
rect 811 917 812 921
rect 806 916 812 917
rect 886 921 892 922
rect 886 917 887 921
rect 891 917 892 921
rect 886 916 892 917
rect 958 921 964 922
rect 958 917 959 921
rect 963 917 964 921
rect 958 916 964 917
rect 1022 921 1028 922
rect 1022 917 1023 921
rect 1027 917 1028 921
rect 1022 916 1028 917
rect 1086 921 1092 922
rect 1086 917 1087 921
rect 1091 917 1092 921
rect 1086 916 1092 917
rect 1150 921 1156 922
rect 1150 917 1151 921
rect 1155 917 1156 921
rect 1150 916 1156 917
rect 1190 921 1196 922
rect 1190 917 1191 921
rect 1195 917 1196 921
rect 1190 916 1196 917
rect 296 899 298 916
rect 344 899 346 916
rect 400 899 402 916
rect 472 899 474 916
rect 552 899 554 916
rect 640 899 642 916
rect 728 899 730 916
rect 808 899 810 916
rect 888 899 890 916
rect 960 899 962 916
rect 1024 899 1026 916
rect 1088 899 1090 916
rect 1152 899 1154 916
rect 1192 899 1194 916
rect 1240 899 1242 939
rect 1278 928 1284 929
rect 1278 924 1279 928
rect 1283 924 1284 928
rect 1278 923 1284 924
rect 2406 928 2412 929
rect 2406 924 2407 928
rect 2411 924 2412 928
rect 2406 923 2412 924
rect 111 898 115 899
rect 111 893 115 894
rect 255 898 259 899
rect 255 893 259 894
rect 295 898 299 899
rect 295 893 299 894
rect 311 898 315 899
rect 311 893 315 894
rect 343 898 347 899
rect 343 893 347 894
rect 375 898 379 899
rect 375 893 379 894
rect 399 898 403 899
rect 399 893 403 894
rect 455 898 459 899
rect 455 893 459 894
rect 471 898 475 899
rect 471 893 475 894
rect 535 898 539 899
rect 535 893 539 894
rect 551 898 555 899
rect 551 893 555 894
rect 623 898 627 899
rect 623 893 627 894
rect 639 898 643 899
rect 639 893 643 894
rect 711 898 715 899
rect 711 893 715 894
rect 727 898 731 899
rect 727 893 731 894
rect 791 898 795 899
rect 791 893 795 894
rect 807 898 811 899
rect 807 893 811 894
rect 863 898 867 899
rect 863 893 867 894
rect 887 898 891 899
rect 887 893 891 894
rect 935 898 939 899
rect 935 893 939 894
rect 959 898 963 899
rect 959 893 963 894
rect 999 898 1003 899
rect 999 893 1003 894
rect 1023 898 1027 899
rect 1023 893 1027 894
rect 1055 898 1059 899
rect 1055 893 1059 894
rect 1087 898 1091 899
rect 1087 893 1091 894
rect 1119 898 1123 899
rect 1119 893 1123 894
rect 1151 898 1155 899
rect 1151 893 1155 894
rect 1183 898 1187 899
rect 1183 893 1187 894
rect 1191 898 1195 899
rect 1191 893 1195 894
rect 1239 898 1243 899
rect 1239 893 1243 894
rect 112 861 114 893
rect 256 884 258 893
rect 312 884 314 893
rect 376 884 378 893
rect 456 884 458 893
rect 536 884 538 893
rect 624 884 626 893
rect 712 884 714 893
rect 792 884 794 893
rect 864 884 866 893
rect 936 884 938 893
rect 1000 884 1002 893
rect 1056 884 1058 893
rect 1120 884 1122 893
rect 1184 884 1186 893
rect 254 883 260 884
rect 254 879 255 883
rect 259 879 260 883
rect 254 878 260 879
rect 310 883 316 884
rect 310 879 311 883
rect 315 879 316 883
rect 310 878 316 879
rect 374 883 380 884
rect 374 879 375 883
rect 379 879 380 883
rect 374 878 380 879
rect 454 883 460 884
rect 454 879 455 883
rect 459 879 460 883
rect 454 878 460 879
rect 534 883 540 884
rect 534 879 535 883
rect 539 879 540 883
rect 534 878 540 879
rect 622 883 628 884
rect 622 879 623 883
rect 627 879 628 883
rect 622 878 628 879
rect 710 883 716 884
rect 710 879 711 883
rect 715 879 716 883
rect 710 878 716 879
rect 790 883 796 884
rect 790 879 791 883
rect 795 879 796 883
rect 790 878 796 879
rect 862 883 868 884
rect 862 879 863 883
rect 867 879 868 883
rect 862 878 868 879
rect 934 883 940 884
rect 934 879 935 883
rect 939 879 940 883
rect 934 878 940 879
rect 998 883 1004 884
rect 998 879 999 883
rect 1003 879 1004 883
rect 998 878 1004 879
rect 1054 883 1060 884
rect 1054 879 1055 883
rect 1059 879 1060 883
rect 1054 878 1060 879
rect 1118 883 1124 884
rect 1118 879 1119 883
rect 1123 879 1124 883
rect 1118 878 1124 879
rect 1182 883 1188 884
rect 1182 879 1183 883
rect 1187 879 1188 883
rect 1182 878 1188 879
rect 1240 861 1242 893
rect 1280 883 1282 923
rect 1318 905 1324 906
rect 1318 901 1319 905
rect 1323 901 1324 905
rect 1318 900 1324 901
rect 1358 905 1364 906
rect 1358 901 1359 905
rect 1363 901 1364 905
rect 1358 900 1364 901
rect 1398 905 1404 906
rect 1398 901 1399 905
rect 1403 901 1404 905
rect 1398 900 1404 901
rect 1462 905 1468 906
rect 1462 901 1463 905
rect 1467 901 1468 905
rect 1462 900 1468 901
rect 1542 905 1548 906
rect 1542 901 1543 905
rect 1547 901 1548 905
rect 1542 900 1548 901
rect 1638 905 1644 906
rect 1638 901 1639 905
rect 1643 901 1644 905
rect 1638 900 1644 901
rect 1734 905 1740 906
rect 1734 901 1735 905
rect 1739 901 1740 905
rect 1734 900 1740 901
rect 1838 905 1844 906
rect 1838 901 1839 905
rect 1843 901 1844 905
rect 1838 900 1844 901
rect 1934 905 1940 906
rect 1934 901 1935 905
rect 1939 901 1940 905
rect 1934 900 1940 901
rect 2022 905 2028 906
rect 2022 901 2023 905
rect 2027 901 2028 905
rect 2022 900 2028 901
rect 2102 905 2108 906
rect 2102 901 2103 905
rect 2107 901 2108 905
rect 2102 900 2108 901
rect 2174 905 2180 906
rect 2174 901 2175 905
rect 2179 901 2180 905
rect 2174 900 2180 901
rect 2238 905 2244 906
rect 2238 901 2239 905
rect 2243 901 2244 905
rect 2238 900 2244 901
rect 2310 905 2316 906
rect 2310 901 2311 905
rect 2315 901 2316 905
rect 2310 900 2316 901
rect 2358 905 2364 906
rect 2358 901 2359 905
rect 2363 901 2364 905
rect 2358 900 2364 901
rect 1320 883 1322 900
rect 1360 883 1362 900
rect 1400 883 1402 900
rect 1464 883 1466 900
rect 1544 883 1546 900
rect 1640 883 1642 900
rect 1736 883 1738 900
rect 1840 883 1842 900
rect 1936 883 1938 900
rect 2024 883 2026 900
rect 2104 883 2106 900
rect 2176 883 2178 900
rect 2240 883 2242 900
rect 2312 883 2314 900
rect 2360 883 2362 900
rect 2408 883 2410 923
rect 1279 882 1283 883
rect 1279 877 1283 878
rect 1319 882 1323 883
rect 1319 877 1323 878
rect 1335 882 1339 883
rect 1335 877 1339 878
rect 1359 882 1363 883
rect 1359 877 1363 878
rect 1375 882 1379 883
rect 1375 877 1379 878
rect 1399 882 1403 883
rect 1399 877 1403 878
rect 1415 882 1419 883
rect 1415 877 1419 878
rect 1463 882 1467 883
rect 1463 877 1467 878
rect 1471 882 1475 883
rect 1471 877 1475 878
rect 1535 882 1539 883
rect 1535 877 1539 878
rect 1543 882 1547 883
rect 1543 877 1547 878
rect 1607 882 1611 883
rect 1607 877 1611 878
rect 1639 882 1643 883
rect 1639 877 1643 878
rect 1679 882 1683 883
rect 1679 877 1683 878
rect 1735 882 1739 883
rect 1735 877 1739 878
rect 1751 882 1755 883
rect 1751 877 1755 878
rect 1823 882 1827 883
rect 1823 877 1827 878
rect 1839 882 1843 883
rect 1839 877 1843 878
rect 1895 882 1899 883
rect 1895 877 1899 878
rect 1935 882 1939 883
rect 1935 877 1939 878
rect 1959 882 1963 883
rect 1959 877 1963 878
rect 2023 882 2027 883
rect 2023 877 2027 878
rect 2087 882 2091 883
rect 2087 877 2091 878
rect 2103 882 2107 883
rect 2103 877 2107 878
rect 2143 882 2147 883
rect 2143 877 2147 878
rect 2175 882 2179 883
rect 2175 877 2179 878
rect 2199 882 2203 883
rect 2199 877 2203 878
rect 2239 882 2243 883
rect 2239 877 2243 878
rect 2255 882 2259 883
rect 2255 877 2259 878
rect 2311 882 2315 883
rect 2311 877 2315 878
rect 2319 882 2323 883
rect 2319 877 2323 878
rect 2359 882 2363 883
rect 2359 877 2363 878
rect 2407 882 2411 883
rect 2407 877 2411 878
rect 110 860 116 861
rect 110 856 111 860
rect 115 856 116 860
rect 110 855 116 856
rect 1238 860 1244 861
rect 1238 856 1239 860
rect 1243 856 1244 860
rect 1238 855 1244 856
rect 1280 845 1282 877
rect 1336 868 1338 877
rect 1376 868 1378 877
rect 1416 868 1418 877
rect 1472 868 1474 877
rect 1536 868 1538 877
rect 1608 868 1610 877
rect 1680 868 1682 877
rect 1752 868 1754 877
rect 1824 868 1826 877
rect 1896 868 1898 877
rect 1960 868 1962 877
rect 2024 868 2026 877
rect 2088 868 2090 877
rect 2144 868 2146 877
rect 2200 868 2202 877
rect 2256 868 2258 877
rect 2320 868 2322 877
rect 2360 868 2362 877
rect 1334 867 1340 868
rect 1334 863 1335 867
rect 1339 863 1340 867
rect 1334 862 1340 863
rect 1374 867 1380 868
rect 1374 863 1375 867
rect 1379 863 1380 867
rect 1374 862 1380 863
rect 1414 867 1420 868
rect 1414 863 1415 867
rect 1419 863 1420 867
rect 1414 862 1420 863
rect 1470 867 1476 868
rect 1470 863 1471 867
rect 1475 863 1476 867
rect 1470 862 1476 863
rect 1534 867 1540 868
rect 1534 863 1535 867
rect 1539 863 1540 867
rect 1534 862 1540 863
rect 1606 867 1612 868
rect 1606 863 1607 867
rect 1611 863 1612 867
rect 1606 862 1612 863
rect 1678 867 1684 868
rect 1678 863 1679 867
rect 1683 863 1684 867
rect 1678 862 1684 863
rect 1750 867 1756 868
rect 1750 863 1751 867
rect 1755 863 1756 867
rect 1750 862 1756 863
rect 1822 867 1828 868
rect 1822 863 1823 867
rect 1827 863 1828 867
rect 1822 862 1828 863
rect 1894 867 1900 868
rect 1894 863 1895 867
rect 1899 863 1900 867
rect 1894 862 1900 863
rect 1958 867 1964 868
rect 1958 863 1959 867
rect 1963 863 1964 867
rect 1958 862 1964 863
rect 2022 867 2028 868
rect 2022 863 2023 867
rect 2027 863 2028 867
rect 2022 862 2028 863
rect 2086 867 2092 868
rect 2086 863 2087 867
rect 2091 863 2092 867
rect 2086 862 2092 863
rect 2142 867 2148 868
rect 2142 863 2143 867
rect 2147 863 2148 867
rect 2142 862 2148 863
rect 2198 867 2204 868
rect 2198 863 2199 867
rect 2203 863 2204 867
rect 2198 862 2204 863
rect 2254 867 2260 868
rect 2254 863 2255 867
rect 2259 863 2260 867
rect 2254 862 2260 863
rect 2318 867 2324 868
rect 2318 863 2319 867
rect 2323 863 2324 867
rect 2318 862 2324 863
rect 2358 867 2364 868
rect 2358 863 2359 867
rect 2363 863 2364 867
rect 2358 862 2364 863
rect 2408 845 2410 877
rect 1278 844 1284 845
rect 110 843 116 844
rect 110 839 111 843
rect 115 839 116 843
rect 110 838 116 839
rect 1238 843 1244 844
rect 1238 839 1239 843
rect 1243 839 1244 843
rect 1278 840 1279 844
rect 1283 840 1284 844
rect 1278 839 1284 840
rect 2406 844 2412 845
rect 2406 840 2407 844
rect 2411 840 2412 844
rect 2406 839 2412 840
rect 1238 838 1244 839
rect 112 831 114 838
rect 254 836 260 837
rect 254 832 255 836
rect 259 832 260 836
rect 254 831 260 832
rect 310 836 316 837
rect 310 832 311 836
rect 315 832 316 836
rect 310 831 316 832
rect 374 836 380 837
rect 374 832 375 836
rect 379 832 380 836
rect 374 831 380 832
rect 454 836 460 837
rect 454 832 455 836
rect 459 832 460 836
rect 454 831 460 832
rect 534 836 540 837
rect 534 832 535 836
rect 539 832 540 836
rect 534 831 540 832
rect 622 836 628 837
rect 622 832 623 836
rect 627 832 628 836
rect 622 831 628 832
rect 710 836 716 837
rect 710 832 711 836
rect 715 832 716 836
rect 710 831 716 832
rect 790 836 796 837
rect 790 832 791 836
rect 795 832 796 836
rect 790 831 796 832
rect 862 836 868 837
rect 862 832 863 836
rect 867 832 868 836
rect 862 831 868 832
rect 934 836 940 837
rect 934 832 935 836
rect 939 832 940 836
rect 934 831 940 832
rect 998 836 1004 837
rect 998 832 999 836
rect 1003 832 1004 836
rect 998 831 1004 832
rect 1054 836 1060 837
rect 1054 832 1055 836
rect 1059 832 1060 836
rect 1054 831 1060 832
rect 1118 836 1124 837
rect 1118 832 1119 836
rect 1123 832 1124 836
rect 1118 831 1124 832
rect 1182 836 1188 837
rect 1182 832 1183 836
rect 1187 832 1188 836
rect 1182 831 1188 832
rect 1240 831 1242 838
rect 111 830 115 831
rect 111 825 115 826
rect 191 830 195 831
rect 191 825 195 826
rect 247 830 251 831
rect 247 825 251 826
rect 255 830 259 831
rect 255 825 259 826
rect 311 830 315 831
rect 311 825 315 826
rect 375 830 379 831
rect 375 825 379 826
rect 383 830 387 831
rect 383 825 387 826
rect 455 830 459 831
rect 455 825 459 826
rect 463 830 467 831
rect 463 825 467 826
rect 535 830 539 831
rect 535 825 539 826
rect 543 830 547 831
rect 543 825 547 826
rect 615 830 619 831
rect 615 825 619 826
rect 623 830 627 831
rect 623 825 627 826
rect 687 830 691 831
rect 687 825 691 826
rect 711 830 715 831
rect 711 825 715 826
rect 751 830 755 831
rect 751 825 755 826
rect 791 830 795 831
rect 791 825 795 826
rect 815 830 819 831
rect 815 825 819 826
rect 863 830 867 831
rect 863 825 867 826
rect 871 830 875 831
rect 871 825 875 826
rect 927 830 931 831
rect 927 825 931 826
rect 935 830 939 831
rect 935 825 939 826
rect 983 830 987 831
rect 983 825 987 826
rect 999 830 1003 831
rect 999 825 1003 826
rect 1047 830 1051 831
rect 1047 825 1051 826
rect 1055 830 1059 831
rect 1055 825 1059 826
rect 1119 830 1123 831
rect 1119 825 1123 826
rect 1183 830 1187 831
rect 1183 825 1187 826
rect 1239 830 1243 831
rect 1239 825 1243 826
rect 1278 827 1284 828
rect 112 818 114 825
rect 190 824 196 825
rect 190 820 191 824
rect 195 820 196 824
rect 190 819 196 820
rect 246 824 252 825
rect 246 820 247 824
rect 251 820 252 824
rect 246 819 252 820
rect 310 824 316 825
rect 310 820 311 824
rect 315 820 316 824
rect 310 819 316 820
rect 382 824 388 825
rect 382 820 383 824
rect 387 820 388 824
rect 382 819 388 820
rect 462 824 468 825
rect 462 820 463 824
rect 467 820 468 824
rect 462 819 468 820
rect 542 824 548 825
rect 542 820 543 824
rect 547 820 548 824
rect 542 819 548 820
rect 614 824 620 825
rect 614 820 615 824
rect 619 820 620 824
rect 614 819 620 820
rect 686 824 692 825
rect 686 820 687 824
rect 691 820 692 824
rect 686 819 692 820
rect 750 824 756 825
rect 750 820 751 824
rect 755 820 756 824
rect 750 819 756 820
rect 814 824 820 825
rect 814 820 815 824
rect 819 820 820 824
rect 814 819 820 820
rect 870 824 876 825
rect 870 820 871 824
rect 875 820 876 824
rect 870 819 876 820
rect 926 824 932 825
rect 926 820 927 824
rect 931 820 932 824
rect 926 819 932 820
rect 982 824 988 825
rect 982 820 983 824
rect 987 820 988 824
rect 982 819 988 820
rect 1046 824 1052 825
rect 1046 820 1047 824
rect 1051 820 1052 824
rect 1046 819 1052 820
rect 1240 818 1242 825
rect 1278 823 1279 827
rect 1283 823 1284 827
rect 1278 822 1284 823
rect 2406 827 2412 828
rect 2406 823 2407 827
rect 2411 823 2412 827
rect 2406 822 2412 823
rect 110 817 116 818
rect 110 813 111 817
rect 115 813 116 817
rect 110 812 116 813
rect 1238 817 1244 818
rect 1238 813 1239 817
rect 1243 813 1244 817
rect 1238 812 1244 813
rect 1280 811 1282 822
rect 1334 820 1340 821
rect 1334 816 1335 820
rect 1339 816 1340 820
rect 1334 815 1340 816
rect 1374 820 1380 821
rect 1374 816 1375 820
rect 1379 816 1380 820
rect 1374 815 1380 816
rect 1414 820 1420 821
rect 1414 816 1415 820
rect 1419 816 1420 820
rect 1414 815 1420 816
rect 1470 820 1476 821
rect 1470 816 1471 820
rect 1475 816 1476 820
rect 1470 815 1476 816
rect 1534 820 1540 821
rect 1534 816 1535 820
rect 1539 816 1540 820
rect 1534 815 1540 816
rect 1606 820 1612 821
rect 1606 816 1607 820
rect 1611 816 1612 820
rect 1606 815 1612 816
rect 1678 820 1684 821
rect 1678 816 1679 820
rect 1683 816 1684 820
rect 1678 815 1684 816
rect 1750 820 1756 821
rect 1750 816 1751 820
rect 1755 816 1756 820
rect 1750 815 1756 816
rect 1822 820 1828 821
rect 1822 816 1823 820
rect 1827 816 1828 820
rect 1822 815 1828 816
rect 1894 820 1900 821
rect 1894 816 1895 820
rect 1899 816 1900 820
rect 1894 815 1900 816
rect 1958 820 1964 821
rect 1958 816 1959 820
rect 1963 816 1964 820
rect 1958 815 1964 816
rect 2022 820 2028 821
rect 2022 816 2023 820
rect 2027 816 2028 820
rect 2022 815 2028 816
rect 2086 820 2092 821
rect 2086 816 2087 820
rect 2091 816 2092 820
rect 2086 815 2092 816
rect 2142 820 2148 821
rect 2142 816 2143 820
rect 2147 816 2148 820
rect 2142 815 2148 816
rect 2198 820 2204 821
rect 2198 816 2199 820
rect 2203 816 2204 820
rect 2198 815 2204 816
rect 2254 820 2260 821
rect 2254 816 2255 820
rect 2259 816 2260 820
rect 2254 815 2260 816
rect 2318 820 2324 821
rect 2318 816 2319 820
rect 2323 816 2324 820
rect 2318 815 2324 816
rect 2358 820 2364 821
rect 2358 816 2359 820
rect 2363 816 2364 820
rect 2358 815 2364 816
rect 1336 811 1338 815
rect 1376 811 1378 815
rect 1416 811 1418 815
rect 1472 811 1474 815
rect 1536 811 1538 815
rect 1608 811 1610 815
rect 1680 811 1682 815
rect 1752 811 1754 815
rect 1824 811 1826 815
rect 1896 811 1898 815
rect 1960 811 1962 815
rect 2024 811 2026 815
rect 2088 811 2090 815
rect 2144 811 2146 815
rect 2200 811 2202 815
rect 2256 811 2258 815
rect 2320 811 2322 815
rect 2360 811 2362 815
rect 2408 811 2410 822
rect 1279 810 1283 811
rect 1279 805 1283 806
rect 1303 810 1307 811
rect 1303 805 1307 806
rect 1335 810 1339 811
rect 1335 805 1339 806
rect 1343 810 1347 811
rect 1343 805 1347 806
rect 1375 810 1379 811
rect 1375 805 1379 806
rect 1407 810 1411 811
rect 1407 805 1411 806
rect 1415 810 1419 811
rect 1415 805 1419 806
rect 1471 810 1475 811
rect 1471 805 1475 806
rect 1479 810 1483 811
rect 1479 805 1483 806
rect 1535 810 1539 811
rect 1535 805 1539 806
rect 1551 810 1555 811
rect 1551 805 1555 806
rect 1607 810 1611 811
rect 1607 805 1611 806
rect 1623 810 1627 811
rect 1623 805 1627 806
rect 1679 810 1683 811
rect 1679 805 1683 806
rect 1695 810 1699 811
rect 1695 805 1699 806
rect 1751 810 1755 811
rect 1751 805 1755 806
rect 1759 810 1763 811
rect 1759 805 1763 806
rect 1823 810 1827 811
rect 1823 805 1827 806
rect 1887 810 1891 811
rect 1887 805 1891 806
rect 1895 810 1899 811
rect 1895 805 1899 806
rect 1951 810 1955 811
rect 1951 805 1955 806
rect 1959 810 1963 811
rect 1959 805 1963 806
rect 2023 810 2027 811
rect 2023 805 2027 806
rect 2087 810 2091 811
rect 2087 805 2091 806
rect 2103 810 2107 811
rect 2103 805 2107 806
rect 2143 810 2147 811
rect 2143 805 2147 806
rect 2191 810 2195 811
rect 2191 805 2195 806
rect 2199 810 2203 811
rect 2199 805 2203 806
rect 2255 810 2259 811
rect 2255 805 2259 806
rect 2279 810 2283 811
rect 2279 805 2283 806
rect 2319 810 2323 811
rect 2319 805 2323 806
rect 2359 810 2363 811
rect 2359 805 2363 806
rect 2407 810 2411 811
rect 2407 805 2411 806
rect 110 800 116 801
rect 110 796 111 800
rect 115 796 116 800
rect 110 795 116 796
rect 1238 800 1244 801
rect 1238 796 1239 800
rect 1243 796 1244 800
rect 1280 798 1282 805
rect 1302 804 1308 805
rect 1302 800 1303 804
rect 1307 800 1308 804
rect 1302 799 1308 800
rect 1342 804 1348 805
rect 1342 800 1343 804
rect 1347 800 1348 804
rect 1342 799 1348 800
rect 1406 804 1412 805
rect 1406 800 1407 804
rect 1411 800 1412 804
rect 1406 799 1412 800
rect 1478 804 1484 805
rect 1478 800 1479 804
rect 1483 800 1484 804
rect 1478 799 1484 800
rect 1550 804 1556 805
rect 1550 800 1551 804
rect 1555 800 1556 804
rect 1550 799 1556 800
rect 1622 804 1628 805
rect 1622 800 1623 804
rect 1627 800 1628 804
rect 1622 799 1628 800
rect 1694 804 1700 805
rect 1694 800 1695 804
rect 1699 800 1700 804
rect 1694 799 1700 800
rect 1758 804 1764 805
rect 1758 800 1759 804
rect 1763 800 1764 804
rect 1758 799 1764 800
rect 1822 804 1828 805
rect 1822 800 1823 804
rect 1827 800 1828 804
rect 1822 799 1828 800
rect 1886 804 1892 805
rect 1886 800 1887 804
rect 1891 800 1892 804
rect 1886 799 1892 800
rect 1950 804 1956 805
rect 1950 800 1951 804
rect 1955 800 1956 804
rect 1950 799 1956 800
rect 2022 804 2028 805
rect 2022 800 2023 804
rect 2027 800 2028 804
rect 2022 799 2028 800
rect 2102 804 2108 805
rect 2102 800 2103 804
rect 2107 800 2108 804
rect 2102 799 2108 800
rect 2190 804 2196 805
rect 2190 800 2191 804
rect 2195 800 2196 804
rect 2190 799 2196 800
rect 2278 804 2284 805
rect 2278 800 2279 804
rect 2283 800 2284 804
rect 2278 799 2284 800
rect 2358 804 2364 805
rect 2358 800 2359 804
rect 2363 800 2364 804
rect 2358 799 2364 800
rect 2408 798 2410 805
rect 1238 795 1244 796
rect 1278 797 1284 798
rect 112 763 114 795
rect 190 777 196 778
rect 190 773 191 777
rect 195 773 196 777
rect 190 772 196 773
rect 246 777 252 778
rect 246 773 247 777
rect 251 773 252 777
rect 246 772 252 773
rect 310 777 316 778
rect 310 773 311 777
rect 315 773 316 777
rect 310 772 316 773
rect 382 777 388 778
rect 382 773 383 777
rect 387 773 388 777
rect 382 772 388 773
rect 462 777 468 778
rect 462 773 463 777
rect 467 773 468 777
rect 462 772 468 773
rect 542 777 548 778
rect 542 773 543 777
rect 547 773 548 777
rect 542 772 548 773
rect 614 777 620 778
rect 614 773 615 777
rect 619 773 620 777
rect 614 772 620 773
rect 686 777 692 778
rect 686 773 687 777
rect 691 773 692 777
rect 686 772 692 773
rect 750 777 756 778
rect 750 773 751 777
rect 755 773 756 777
rect 750 772 756 773
rect 814 777 820 778
rect 814 773 815 777
rect 819 773 820 777
rect 814 772 820 773
rect 870 777 876 778
rect 870 773 871 777
rect 875 773 876 777
rect 870 772 876 773
rect 926 777 932 778
rect 926 773 927 777
rect 931 773 932 777
rect 926 772 932 773
rect 982 777 988 778
rect 982 773 983 777
rect 987 773 988 777
rect 982 772 988 773
rect 1046 777 1052 778
rect 1046 773 1047 777
rect 1051 773 1052 777
rect 1046 772 1052 773
rect 192 763 194 772
rect 248 763 250 772
rect 312 763 314 772
rect 384 763 386 772
rect 464 763 466 772
rect 544 763 546 772
rect 616 763 618 772
rect 688 763 690 772
rect 752 763 754 772
rect 816 763 818 772
rect 872 763 874 772
rect 928 763 930 772
rect 984 763 986 772
rect 1048 763 1050 772
rect 1240 763 1242 795
rect 1278 793 1279 797
rect 1283 793 1284 797
rect 1278 792 1284 793
rect 2406 797 2412 798
rect 2406 793 2407 797
rect 2411 793 2412 797
rect 2406 792 2412 793
rect 1278 780 1284 781
rect 1278 776 1279 780
rect 1283 776 1284 780
rect 1278 775 1284 776
rect 2406 780 2412 781
rect 2406 776 2407 780
rect 2411 776 2412 780
rect 2406 775 2412 776
rect 111 762 115 763
rect 111 757 115 758
rect 135 762 139 763
rect 135 757 139 758
rect 175 762 179 763
rect 175 757 179 758
rect 191 762 195 763
rect 191 757 195 758
rect 215 762 219 763
rect 215 757 219 758
rect 247 762 251 763
rect 247 757 251 758
rect 279 762 283 763
rect 279 757 283 758
rect 311 762 315 763
rect 311 757 315 758
rect 351 762 355 763
rect 351 757 355 758
rect 383 762 387 763
rect 383 757 387 758
rect 423 762 427 763
rect 423 757 427 758
rect 463 762 467 763
rect 463 757 467 758
rect 495 762 499 763
rect 495 757 499 758
rect 543 762 547 763
rect 543 757 547 758
rect 559 762 563 763
rect 559 757 563 758
rect 615 762 619 763
rect 615 757 619 758
rect 623 762 627 763
rect 623 757 627 758
rect 687 762 691 763
rect 687 757 691 758
rect 695 762 699 763
rect 695 757 699 758
rect 751 762 755 763
rect 751 757 755 758
rect 783 762 787 763
rect 783 757 787 758
rect 815 762 819 763
rect 815 757 819 758
rect 871 762 875 763
rect 871 757 875 758
rect 879 762 883 763
rect 879 757 883 758
rect 927 762 931 763
rect 927 757 931 758
rect 983 762 987 763
rect 983 757 987 758
rect 1047 762 1051 763
rect 1047 757 1051 758
rect 1095 762 1099 763
rect 1095 757 1099 758
rect 1191 762 1195 763
rect 1191 757 1195 758
rect 1239 762 1243 763
rect 1239 757 1243 758
rect 112 725 114 757
rect 136 748 138 757
rect 176 748 178 757
rect 216 748 218 757
rect 280 748 282 757
rect 352 748 354 757
rect 424 748 426 757
rect 496 748 498 757
rect 560 748 562 757
rect 624 748 626 757
rect 696 748 698 757
rect 784 748 786 757
rect 880 748 882 757
rect 984 748 986 757
rect 1096 748 1098 757
rect 1192 748 1194 757
rect 134 747 140 748
rect 134 743 135 747
rect 139 743 140 747
rect 134 742 140 743
rect 174 747 180 748
rect 174 743 175 747
rect 179 743 180 747
rect 174 742 180 743
rect 214 747 220 748
rect 214 743 215 747
rect 219 743 220 747
rect 214 742 220 743
rect 278 747 284 748
rect 278 743 279 747
rect 283 743 284 747
rect 278 742 284 743
rect 350 747 356 748
rect 350 743 351 747
rect 355 743 356 747
rect 350 742 356 743
rect 422 747 428 748
rect 422 743 423 747
rect 427 743 428 747
rect 422 742 428 743
rect 494 747 500 748
rect 494 743 495 747
rect 499 743 500 747
rect 494 742 500 743
rect 558 747 564 748
rect 558 743 559 747
rect 563 743 564 747
rect 558 742 564 743
rect 622 747 628 748
rect 622 743 623 747
rect 627 743 628 747
rect 622 742 628 743
rect 694 747 700 748
rect 694 743 695 747
rect 699 743 700 747
rect 694 742 700 743
rect 782 747 788 748
rect 782 743 783 747
rect 787 743 788 747
rect 782 742 788 743
rect 878 747 884 748
rect 878 743 879 747
rect 883 743 884 747
rect 878 742 884 743
rect 982 747 988 748
rect 982 743 983 747
rect 987 743 988 747
rect 982 742 988 743
rect 1094 747 1100 748
rect 1094 743 1095 747
rect 1099 743 1100 747
rect 1094 742 1100 743
rect 1190 747 1196 748
rect 1190 743 1191 747
rect 1195 743 1196 747
rect 1190 742 1196 743
rect 1240 725 1242 757
rect 1280 743 1282 775
rect 1302 757 1308 758
rect 1302 753 1303 757
rect 1307 753 1308 757
rect 1302 752 1308 753
rect 1342 757 1348 758
rect 1342 753 1343 757
rect 1347 753 1348 757
rect 1342 752 1348 753
rect 1406 757 1412 758
rect 1406 753 1407 757
rect 1411 753 1412 757
rect 1406 752 1412 753
rect 1478 757 1484 758
rect 1478 753 1479 757
rect 1483 753 1484 757
rect 1478 752 1484 753
rect 1550 757 1556 758
rect 1550 753 1551 757
rect 1555 753 1556 757
rect 1550 752 1556 753
rect 1622 757 1628 758
rect 1622 753 1623 757
rect 1627 753 1628 757
rect 1622 752 1628 753
rect 1694 757 1700 758
rect 1694 753 1695 757
rect 1699 753 1700 757
rect 1694 752 1700 753
rect 1758 757 1764 758
rect 1758 753 1759 757
rect 1763 753 1764 757
rect 1758 752 1764 753
rect 1822 757 1828 758
rect 1822 753 1823 757
rect 1827 753 1828 757
rect 1822 752 1828 753
rect 1886 757 1892 758
rect 1886 753 1887 757
rect 1891 753 1892 757
rect 1886 752 1892 753
rect 1950 757 1956 758
rect 1950 753 1951 757
rect 1955 753 1956 757
rect 1950 752 1956 753
rect 2022 757 2028 758
rect 2022 753 2023 757
rect 2027 753 2028 757
rect 2022 752 2028 753
rect 2102 757 2108 758
rect 2102 753 2103 757
rect 2107 753 2108 757
rect 2102 752 2108 753
rect 2190 757 2196 758
rect 2190 753 2191 757
rect 2195 753 2196 757
rect 2190 752 2196 753
rect 2278 757 2284 758
rect 2278 753 2279 757
rect 2283 753 2284 757
rect 2278 752 2284 753
rect 2358 757 2364 758
rect 2358 753 2359 757
rect 2363 753 2364 757
rect 2358 752 2364 753
rect 1304 743 1306 752
rect 1344 743 1346 752
rect 1408 743 1410 752
rect 1480 743 1482 752
rect 1552 743 1554 752
rect 1624 743 1626 752
rect 1696 743 1698 752
rect 1760 743 1762 752
rect 1824 743 1826 752
rect 1888 743 1890 752
rect 1952 743 1954 752
rect 2024 743 2026 752
rect 2104 743 2106 752
rect 2192 743 2194 752
rect 2280 743 2282 752
rect 2360 743 2362 752
rect 2408 743 2410 775
rect 1279 742 1283 743
rect 1279 737 1283 738
rect 1303 742 1307 743
rect 1303 737 1307 738
rect 1343 742 1347 743
rect 1343 737 1347 738
rect 1367 742 1371 743
rect 1367 737 1371 738
rect 1407 742 1411 743
rect 1407 737 1411 738
rect 1455 742 1459 743
rect 1455 737 1459 738
rect 1479 742 1483 743
rect 1479 737 1483 738
rect 1535 742 1539 743
rect 1535 737 1539 738
rect 1551 742 1555 743
rect 1551 737 1555 738
rect 1615 742 1619 743
rect 1615 737 1619 738
rect 1623 742 1627 743
rect 1623 737 1627 738
rect 1695 742 1699 743
rect 1695 737 1699 738
rect 1759 742 1763 743
rect 1759 737 1763 738
rect 1775 742 1779 743
rect 1775 737 1779 738
rect 1823 742 1827 743
rect 1823 737 1827 738
rect 1855 742 1859 743
rect 1855 737 1859 738
rect 1887 742 1891 743
rect 1887 737 1891 738
rect 1943 742 1947 743
rect 1943 737 1947 738
rect 1951 742 1955 743
rect 1951 737 1955 738
rect 2023 742 2027 743
rect 2023 737 2027 738
rect 2031 742 2035 743
rect 2031 737 2035 738
rect 2103 742 2107 743
rect 2103 737 2107 738
rect 2119 742 2123 743
rect 2119 737 2123 738
rect 2191 742 2195 743
rect 2191 737 2195 738
rect 2207 742 2211 743
rect 2207 737 2211 738
rect 2279 742 2283 743
rect 2279 737 2283 738
rect 2295 742 2299 743
rect 2295 737 2299 738
rect 2359 742 2363 743
rect 2359 737 2363 738
rect 2407 742 2411 743
rect 2407 737 2411 738
rect 110 724 116 725
rect 110 720 111 724
rect 115 720 116 724
rect 110 719 116 720
rect 1238 724 1244 725
rect 1238 720 1239 724
rect 1243 720 1244 724
rect 1238 719 1244 720
rect 110 707 116 708
rect 110 703 111 707
rect 115 703 116 707
rect 110 702 116 703
rect 1238 707 1244 708
rect 1238 703 1239 707
rect 1243 703 1244 707
rect 1280 705 1282 737
rect 1304 728 1306 737
rect 1368 728 1370 737
rect 1456 728 1458 737
rect 1536 728 1538 737
rect 1616 728 1618 737
rect 1696 728 1698 737
rect 1776 728 1778 737
rect 1856 728 1858 737
rect 1944 728 1946 737
rect 2032 728 2034 737
rect 2120 728 2122 737
rect 2208 728 2210 737
rect 2296 728 2298 737
rect 2360 728 2362 737
rect 1302 727 1308 728
rect 1302 723 1303 727
rect 1307 723 1308 727
rect 1302 722 1308 723
rect 1366 727 1372 728
rect 1366 723 1367 727
rect 1371 723 1372 727
rect 1366 722 1372 723
rect 1454 727 1460 728
rect 1454 723 1455 727
rect 1459 723 1460 727
rect 1454 722 1460 723
rect 1534 727 1540 728
rect 1534 723 1535 727
rect 1539 723 1540 727
rect 1534 722 1540 723
rect 1614 727 1620 728
rect 1614 723 1615 727
rect 1619 723 1620 727
rect 1614 722 1620 723
rect 1694 727 1700 728
rect 1694 723 1695 727
rect 1699 723 1700 727
rect 1694 722 1700 723
rect 1774 727 1780 728
rect 1774 723 1775 727
rect 1779 723 1780 727
rect 1774 722 1780 723
rect 1854 727 1860 728
rect 1854 723 1855 727
rect 1859 723 1860 727
rect 1854 722 1860 723
rect 1942 727 1948 728
rect 1942 723 1943 727
rect 1947 723 1948 727
rect 1942 722 1948 723
rect 2030 727 2036 728
rect 2030 723 2031 727
rect 2035 723 2036 727
rect 2030 722 2036 723
rect 2118 727 2124 728
rect 2118 723 2119 727
rect 2123 723 2124 727
rect 2118 722 2124 723
rect 2206 727 2212 728
rect 2206 723 2207 727
rect 2211 723 2212 727
rect 2206 722 2212 723
rect 2294 727 2300 728
rect 2294 723 2295 727
rect 2299 723 2300 727
rect 2294 722 2300 723
rect 2358 727 2364 728
rect 2358 723 2359 727
rect 2363 723 2364 727
rect 2358 722 2364 723
rect 2408 705 2410 737
rect 1238 702 1244 703
rect 1278 704 1284 705
rect 112 687 114 702
rect 134 700 140 701
rect 134 696 135 700
rect 139 696 140 700
rect 134 695 140 696
rect 174 700 180 701
rect 174 696 175 700
rect 179 696 180 700
rect 174 695 180 696
rect 214 700 220 701
rect 214 696 215 700
rect 219 696 220 700
rect 214 695 220 696
rect 278 700 284 701
rect 278 696 279 700
rect 283 696 284 700
rect 278 695 284 696
rect 350 700 356 701
rect 350 696 351 700
rect 355 696 356 700
rect 350 695 356 696
rect 422 700 428 701
rect 422 696 423 700
rect 427 696 428 700
rect 422 695 428 696
rect 494 700 500 701
rect 494 696 495 700
rect 499 696 500 700
rect 494 695 500 696
rect 558 700 564 701
rect 558 696 559 700
rect 563 696 564 700
rect 558 695 564 696
rect 622 700 628 701
rect 622 696 623 700
rect 627 696 628 700
rect 622 695 628 696
rect 694 700 700 701
rect 694 696 695 700
rect 699 696 700 700
rect 694 695 700 696
rect 782 700 788 701
rect 782 696 783 700
rect 787 696 788 700
rect 782 695 788 696
rect 878 700 884 701
rect 878 696 879 700
rect 883 696 884 700
rect 878 695 884 696
rect 982 700 988 701
rect 982 696 983 700
rect 987 696 988 700
rect 982 695 988 696
rect 1094 700 1100 701
rect 1094 696 1095 700
rect 1099 696 1100 700
rect 1094 695 1100 696
rect 1190 700 1196 701
rect 1190 696 1191 700
rect 1195 696 1196 700
rect 1190 695 1196 696
rect 136 687 138 695
rect 176 687 178 695
rect 216 687 218 695
rect 280 687 282 695
rect 352 687 354 695
rect 424 687 426 695
rect 496 687 498 695
rect 560 687 562 695
rect 624 687 626 695
rect 696 687 698 695
rect 784 687 786 695
rect 880 687 882 695
rect 984 687 986 695
rect 1096 687 1098 695
rect 1192 687 1194 695
rect 1240 687 1242 702
rect 1278 700 1279 704
rect 1283 700 1284 704
rect 1278 699 1284 700
rect 2406 704 2412 705
rect 2406 700 2407 704
rect 2411 700 2412 704
rect 2406 699 2412 700
rect 1278 687 1284 688
rect 111 686 115 687
rect 111 681 115 682
rect 135 686 139 687
rect 135 681 139 682
rect 175 686 179 687
rect 175 681 179 682
rect 215 686 219 687
rect 215 681 219 682
rect 231 686 235 687
rect 231 681 235 682
rect 279 686 283 687
rect 279 681 283 682
rect 287 686 291 687
rect 287 681 291 682
rect 343 686 347 687
rect 343 681 347 682
rect 351 686 355 687
rect 351 681 355 682
rect 399 686 403 687
rect 399 681 403 682
rect 423 686 427 687
rect 423 681 427 682
rect 455 686 459 687
rect 455 681 459 682
rect 495 686 499 687
rect 495 681 499 682
rect 503 686 507 687
rect 503 681 507 682
rect 559 686 563 687
rect 559 681 563 682
rect 623 686 627 687
rect 623 681 627 682
rect 695 686 699 687
rect 695 681 699 682
rect 767 686 771 687
rect 767 681 771 682
rect 783 686 787 687
rect 783 681 787 682
rect 839 686 843 687
rect 839 681 843 682
rect 879 686 883 687
rect 879 681 883 682
rect 903 686 907 687
rect 903 681 907 682
rect 967 686 971 687
rect 967 681 971 682
rect 983 686 987 687
rect 983 681 987 682
rect 1023 686 1027 687
rect 1023 681 1027 682
rect 1087 686 1091 687
rect 1087 681 1091 682
rect 1095 686 1099 687
rect 1095 681 1099 682
rect 1151 686 1155 687
rect 1151 681 1155 682
rect 1191 686 1195 687
rect 1191 681 1195 682
rect 1239 686 1243 687
rect 1278 683 1279 687
rect 1283 683 1284 687
rect 1278 682 1284 683
rect 2406 687 2412 688
rect 2406 683 2407 687
rect 2411 683 2412 687
rect 2406 682 2412 683
rect 1239 681 1243 682
rect 112 674 114 681
rect 134 680 140 681
rect 134 676 135 680
rect 139 676 140 680
rect 134 675 140 676
rect 174 680 180 681
rect 174 676 175 680
rect 179 676 180 680
rect 174 675 180 676
rect 230 680 236 681
rect 230 676 231 680
rect 235 676 236 680
rect 230 675 236 676
rect 286 680 292 681
rect 286 676 287 680
rect 291 676 292 680
rect 286 675 292 676
rect 342 680 348 681
rect 342 676 343 680
rect 347 676 348 680
rect 342 675 348 676
rect 398 680 404 681
rect 398 676 399 680
rect 403 676 404 680
rect 398 675 404 676
rect 454 680 460 681
rect 454 676 455 680
rect 459 676 460 680
rect 454 675 460 676
rect 502 680 508 681
rect 502 676 503 680
rect 507 676 508 680
rect 502 675 508 676
rect 558 680 564 681
rect 558 676 559 680
rect 563 676 564 680
rect 558 675 564 676
rect 622 680 628 681
rect 622 676 623 680
rect 627 676 628 680
rect 622 675 628 676
rect 694 680 700 681
rect 694 676 695 680
rect 699 676 700 680
rect 694 675 700 676
rect 766 680 772 681
rect 766 676 767 680
rect 771 676 772 680
rect 766 675 772 676
rect 838 680 844 681
rect 838 676 839 680
rect 843 676 844 680
rect 838 675 844 676
rect 902 680 908 681
rect 902 676 903 680
rect 907 676 908 680
rect 902 675 908 676
rect 966 680 972 681
rect 966 676 967 680
rect 971 676 972 680
rect 966 675 972 676
rect 1022 680 1028 681
rect 1022 676 1023 680
rect 1027 676 1028 680
rect 1022 675 1028 676
rect 1086 680 1092 681
rect 1086 676 1087 680
rect 1091 676 1092 680
rect 1086 675 1092 676
rect 1150 680 1156 681
rect 1150 676 1151 680
rect 1155 676 1156 680
rect 1150 675 1156 676
rect 1190 680 1196 681
rect 1190 676 1191 680
rect 1195 676 1196 680
rect 1190 675 1196 676
rect 1240 674 1242 681
rect 1280 675 1282 682
rect 1302 680 1308 681
rect 1302 676 1303 680
rect 1307 676 1308 680
rect 1302 675 1308 676
rect 1366 680 1372 681
rect 1366 676 1367 680
rect 1371 676 1372 680
rect 1366 675 1372 676
rect 1454 680 1460 681
rect 1454 676 1455 680
rect 1459 676 1460 680
rect 1454 675 1460 676
rect 1534 680 1540 681
rect 1534 676 1535 680
rect 1539 676 1540 680
rect 1534 675 1540 676
rect 1614 680 1620 681
rect 1614 676 1615 680
rect 1619 676 1620 680
rect 1614 675 1620 676
rect 1694 680 1700 681
rect 1694 676 1695 680
rect 1699 676 1700 680
rect 1694 675 1700 676
rect 1774 680 1780 681
rect 1774 676 1775 680
rect 1779 676 1780 680
rect 1774 675 1780 676
rect 1854 680 1860 681
rect 1854 676 1855 680
rect 1859 676 1860 680
rect 1854 675 1860 676
rect 1942 680 1948 681
rect 1942 676 1943 680
rect 1947 676 1948 680
rect 1942 675 1948 676
rect 2030 680 2036 681
rect 2030 676 2031 680
rect 2035 676 2036 680
rect 2030 675 2036 676
rect 2118 680 2124 681
rect 2118 676 2119 680
rect 2123 676 2124 680
rect 2118 675 2124 676
rect 2206 680 2212 681
rect 2206 676 2207 680
rect 2211 676 2212 680
rect 2206 675 2212 676
rect 2294 680 2300 681
rect 2294 676 2295 680
rect 2299 676 2300 680
rect 2294 675 2300 676
rect 2358 680 2364 681
rect 2358 676 2359 680
rect 2363 676 2364 680
rect 2358 675 2364 676
rect 2408 675 2410 682
rect 1279 674 1283 675
rect 110 673 116 674
rect 110 669 111 673
rect 115 669 116 673
rect 110 668 116 669
rect 1238 673 1244 674
rect 1238 669 1239 673
rect 1243 669 1244 673
rect 1279 669 1283 670
rect 1303 674 1307 675
rect 1303 669 1307 670
rect 1367 674 1371 675
rect 1367 669 1371 670
rect 1455 674 1459 675
rect 1455 669 1459 670
rect 1535 674 1539 675
rect 1535 669 1539 670
rect 1591 674 1595 675
rect 1591 669 1595 670
rect 1615 674 1619 675
rect 1615 669 1619 670
rect 1639 674 1643 675
rect 1639 669 1643 670
rect 1687 674 1691 675
rect 1687 669 1691 670
rect 1695 674 1699 675
rect 1695 669 1699 670
rect 1743 674 1747 675
rect 1743 669 1747 670
rect 1775 674 1779 675
rect 1775 669 1779 670
rect 1799 674 1803 675
rect 1799 669 1803 670
rect 1855 674 1859 675
rect 1855 669 1859 670
rect 1871 674 1875 675
rect 1871 669 1875 670
rect 1943 674 1947 675
rect 1943 669 1947 670
rect 1951 674 1955 675
rect 1951 669 1955 670
rect 2031 674 2035 675
rect 2031 669 2035 670
rect 2047 674 2051 675
rect 2047 669 2051 670
rect 2119 674 2123 675
rect 2119 669 2123 670
rect 2151 674 2155 675
rect 2151 669 2155 670
rect 2207 674 2211 675
rect 2207 669 2211 670
rect 2263 674 2267 675
rect 2263 669 2267 670
rect 2295 674 2299 675
rect 2295 669 2299 670
rect 2359 674 2363 675
rect 2359 669 2363 670
rect 2407 674 2411 675
rect 2407 669 2411 670
rect 1238 668 1244 669
rect 1280 662 1282 669
rect 1590 668 1596 669
rect 1590 664 1591 668
rect 1595 664 1596 668
rect 1590 663 1596 664
rect 1638 668 1644 669
rect 1638 664 1639 668
rect 1643 664 1644 668
rect 1638 663 1644 664
rect 1686 668 1692 669
rect 1686 664 1687 668
rect 1691 664 1692 668
rect 1686 663 1692 664
rect 1742 668 1748 669
rect 1742 664 1743 668
rect 1747 664 1748 668
rect 1742 663 1748 664
rect 1798 668 1804 669
rect 1798 664 1799 668
rect 1803 664 1804 668
rect 1798 663 1804 664
rect 1870 668 1876 669
rect 1870 664 1871 668
rect 1875 664 1876 668
rect 1870 663 1876 664
rect 1950 668 1956 669
rect 1950 664 1951 668
rect 1955 664 1956 668
rect 1950 663 1956 664
rect 2046 668 2052 669
rect 2046 664 2047 668
rect 2051 664 2052 668
rect 2046 663 2052 664
rect 2150 668 2156 669
rect 2150 664 2151 668
rect 2155 664 2156 668
rect 2150 663 2156 664
rect 2262 668 2268 669
rect 2262 664 2263 668
rect 2267 664 2268 668
rect 2262 663 2268 664
rect 2358 668 2364 669
rect 2358 664 2359 668
rect 2363 664 2364 668
rect 2358 663 2364 664
rect 2408 662 2410 669
rect 1278 661 1284 662
rect 1278 657 1279 661
rect 1283 657 1284 661
rect 110 656 116 657
rect 110 652 111 656
rect 115 652 116 656
rect 110 651 116 652
rect 1238 656 1244 657
rect 1278 656 1284 657
rect 2406 661 2412 662
rect 2406 657 2407 661
rect 2411 657 2412 661
rect 2406 656 2412 657
rect 1238 652 1239 656
rect 1243 652 1244 656
rect 1238 651 1244 652
rect 112 619 114 651
rect 134 633 140 634
rect 134 629 135 633
rect 139 629 140 633
rect 134 628 140 629
rect 174 633 180 634
rect 174 629 175 633
rect 179 629 180 633
rect 174 628 180 629
rect 230 633 236 634
rect 230 629 231 633
rect 235 629 236 633
rect 230 628 236 629
rect 286 633 292 634
rect 286 629 287 633
rect 291 629 292 633
rect 286 628 292 629
rect 342 633 348 634
rect 342 629 343 633
rect 347 629 348 633
rect 342 628 348 629
rect 398 633 404 634
rect 398 629 399 633
rect 403 629 404 633
rect 398 628 404 629
rect 454 633 460 634
rect 454 629 455 633
rect 459 629 460 633
rect 454 628 460 629
rect 502 633 508 634
rect 502 629 503 633
rect 507 629 508 633
rect 502 628 508 629
rect 558 633 564 634
rect 558 629 559 633
rect 563 629 564 633
rect 558 628 564 629
rect 622 633 628 634
rect 622 629 623 633
rect 627 629 628 633
rect 622 628 628 629
rect 694 633 700 634
rect 694 629 695 633
rect 699 629 700 633
rect 694 628 700 629
rect 766 633 772 634
rect 766 629 767 633
rect 771 629 772 633
rect 766 628 772 629
rect 838 633 844 634
rect 838 629 839 633
rect 843 629 844 633
rect 838 628 844 629
rect 902 633 908 634
rect 902 629 903 633
rect 907 629 908 633
rect 902 628 908 629
rect 966 633 972 634
rect 966 629 967 633
rect 971 629 972 633
rect 966 628 972 629
rect 1022 633 1028 634
rect 1022 629 1023 633
rect 1027 629 1028 633
rect 1022 628 1028 629
rect 1086 633 1092 634
rect 1086 629 1087 633
rect 1091 629 1092 633
rect 1086 628 1092 629
rect 1150 633 1156 634
rect 1150 629 1151 633
rect 1155 629 1156 633
rect 1150 628 1156 629
rect 1190 633 1196 634
rect 1190 629 1191 633
rect 1195 629 1196 633
rect 1190 628 1196 629
rect 136 619 138 628
rect 176 619 178 628
rect 232 619 234 628
rect 288 619 290 628
rect 344 619 346 628
rect 400 619 402 628
rect 456 619 458 628
rect 504 619 506 628
rect 560 619 562 628
rect 624 619 626 628
rect 696 619 698 628
rect 768 619 770 628
rect 840 619 842 628
rect 904 619 906 628
rect 968 619 970 628
rect 1024 619 1026 628
rect 1088 619 1090 628
rect 1152 619 1154 628
rect 1192 619 1194 628
rect 1240 619 1242 651
rect 1278 644 1284 645
rect 1278 640 1279 644
rect 1283 640 1284 644
rect 1278 639 1284 640
rect 2406 644 2412 645
rect 2406 640 2407 644
rect 2411 640 2412 644
rect 2406 639 2412 640
rect 111 618 115 619
rect 111 613 115 614
rect 135 618 139 619
rect 135 613 139 614
rect 175 618 179 619
rect 175 613 179 614
rect 183 618 187 619
rect 183 613 187 614
rect 231 618 235 619
rect 231 613 235 614
rect 255 618 259 619
rect 255 613 259 614
rect 287 618 291 619
rect 287 613 291 614
rect 327 618 331 619
rect 327 613 331 614
rect 343 618 347 619
rect 343 613 347 614
rect 399 618 403 619
rect 399 613 403 614
rect 455 618 459 619
rect 455 613 459 614
rect 479 618 483 619
rect 479 613 483 614
rect 503 618 507 619
rect 503 613 507 614
rect 559 618 563 619
rect 559 613 563 614
rect 623 618 627 619
rect 623 613 627 614
rect 639 618 643 619
rect 639 613 643 614
rect 695 618 699 619
rect 695 613 699 614
rect 719 618 723 619
rect 719 613 723 614
rect 767 618 771 619
rect 767 613 771 614
rect 799 618 803 619
rect 799 613 803 614
rect 839 618 843 619
rect 839 613 843 614
rect 879 618 883 619
rect 879 613 883 614
rect 903 618 907 619
rect 903 613 907 614
rect 951 618 955 619
rect 951 613 955 614
rect 967 618 971 619
rect 967 613 971 614
rect 1015 618 1019 619
rect 1015 613 1019 614
rect 1023 618 1027 619
rect 1023 613 1027 614
rect 1079 618 1083 619
rect 1079 613 1083 614
rect 1087 618 1091 619
rect 1087 613 1091 614
rect 1143 618 1147 619
rect 1143 613 1147 614
rect 1151 618 1155 619
rect 1151 613 1155 614
rect 1191 618 1195 619
rect 1191 613 1195 614
rect 1239 618 1243 619
rect 1239 613 1243 614
rect 112 581 114 613
rect 136 604 138 613
rect 184 604 186 613
rect 256 604 258 613
rect 328 604 330 613
rect 400 604 402 613
rect 480 604 482 613
rect 560 604 562 613
rect 640 604 642 613
rect 720 604 722 613
rect 800 604 802 613
rect 880 604 882 613
rect 952 604 954 613
rect 1016 604 1018 613
rect 1080 604 1082 613
rect 1144 604 1146 613
rect 1192 604 1194 613
rect 134 603 140 604
rect 134 599 135 603
rect 139 599 140 603
rect 134 598 140 599
rect 182 603 188 604
rect 182 599 183 603
rect 187 599 188 603
rect 182 598 188 599
rect 254 603 260 604
rect 254 599 255 603
rect 259 599 260 603
rect 254 598 260 599
rect 326 603 332 604
rect 326 599 327 603
rect 331 599 332 603
rect 326 598 332 599
rect 398 603 404 604
rect 398 599 399 603
rect 403 599 404 603
rect 398 598 404 599
rect 478 603 484 604
rect 478 599 479 603
rect 483 599 484 603
rect 478 598 484 599
rect 558 603 564 604
rect 558 599 559 603
rect 563 599 564 603
rect 558 598 564 599
rect 638 603 644 604
rect 638 599 639 603
rect 643 599 644 603
rect 638 598 644 599
rect 718 603 724 604
rect 718 599 719 603
rect 723 599 724 603
rect 718 598 724 599
rect 798 603 804 604
rect 798 599 799 603
rect 803 599 804 603
rect 798 598 804 599
rect 878 603 884 604
rect 878 599 879 603
rect 883 599 884 603
rect 878 598 884 599
rect 950 603 956 604
rect 950 599 951 603
rect 955 599 956 603
rect 950 598 956 599
rect 1014 603 1020 604
rect 1014 599 1015 603
rect 1019 599 1020 603
rect 1014 598 1020 599
rect 1078 603 1084 604
rect 1078 599 1079 603
rect 1083 599 1084 603
rect 1078 598 1084 599
rect 1142 603 1148 604
rect 1142 599 1143 603
rect 1147 599 1148 603
rect 1142 598 1148 599
rect 1190 603 1196 604
rect 1190 599 1191 603
rect 1195 599 1196 603
rect 1190 598 1196 599
rect 1240 581 1242 613
rect 1280 599 1282 639
rect 1590 621 1596 622
rect 1590 617 1591 621
rect 1595 617 1596 621
rect 1590 616 1596 617
rect 1638 621 1644 622
rect 1638 617 1639 621
rect 1643 617 1644 621
rect 1638 616 1644 617
rect 1686 621 1692 622
rect 1686 617 1687 621
rect 1691 617 1692 621
rect 1686 616 1692 617
rect 1742 621 1748 622
rect 1742 617 1743 621
rect 1747 617 1748 621
rect 1742 616 1748 617
rect 1798 621 1804 622
rect 1798 617 1799 621
rect 1803 617 1804 621
rect 1798 616 1804 617
rect 1870 621 1876 622
rect 1870 617 1871 621
rect 1875 617 1876 621
rect 1870 616 1876 617
rect 1950 621 1956 622
rect 1950 617 1951 621
rect 1955 617 1956 621
rect 1950 616 1956 617
rect 2046 621 2052 622
rect 2046 617 2047 621
rect 2051 617 2052 621
rect 2046 616 2052 617
rect 2150 621 2156 622
rect 2150 617 2151 621
rect 2155 617 2156 621
rect 2150 616 2156 617
rect 2262 621 2268 622
rect 2262 617 2263 621
rect 2267 617 2268 621
rect 2262 616 2268 617
rect 2358 621 2364 622
rect 2358 617 2359 621
rect 2363 617 2364 621
rect 2358 616 2364 617
rect 1592 599 1594 616
rect 1640 599 1642 616
rect 1688 599 1690 616
rect 1744 599 1746 616
rect 1800 599 1802 616
rect 1872 599 1874 616
rect 1952 599 1954 616
rect 2048 599 2050 616
rect 2152 599 2154 616
rect 2264 599 2266 616
rect 2360 599 2362 616
rect 2408 599 2410 639
rect 1279 598 1283 599
rect 1279 593 1283 594
rect 1559 598 1563 599
rect 1559 593 1563 594
rect 1591 598 1595 599
rect 1591 593 1595 594
rect 1599 598 1603 599
rect 1599 593 1603 594
rect 1639 598 1643 599
rect 1639 593 1643 594
rect 1679 598 1683 599
rect 1679 593 1683 594
rect 1687 598 1691 599
rect 1687 593 1691 594
rect 1719 598 1723 599
rect 1719 593 1723 594
rect 1743 598 1747 599
rect 1743 593 1747 594
rect 1759 598 1763 599
rect 1759 593 1763 594
rect 1799 598 1803 599
rect 1799 593 1803 594
rect 1807 598 1811 599
rect 1807 593 1811 594
rect 1855 598 1859 599
rect 1855 593 1859 594
rect 1871 598 1875 599
rect 1871 593 1875 594
rect 1911 598 1915 599
rect 1911 593 1915 594
rect 1951 598 1955 599
rect 1951 593 1955 594
rect 1967 598 1971 599
rect 1967 593 1971 594
rect 2031 598 2035 599
rect 2031 593 2035 594
rect 2047 598 2051 599
rect 2047 593 2051 594
rect 2095 598 2099 599
rect 2095 593 2099 594
rect 2151 598 2155 599
rect 2151 593 2155 594
rect 2167 598 2171 599
rect 2167 593 2171 594
rect 2239 598 2243 599
rect 2239 593 2243 594
rect 2263 598 2267 599
rect 2263 593 2267 594
rect 2311 598 2315 599
rect 2311 593 2315 594
rect 2359 598 2363 599
rect 2359 593 2363 594
rect 2407 598 2411 599
rect 2407 593 2411 594
rect 110 580 116 581
rect 110 576 111 580
rect 115 576 116 580
rect 110 575 116 576
rect 1238 580 1244 581
rect 1238 576 1239 580
rect 1243 576 1244 580
rect 1238 575 1244 576
rect 110 563 116 564
rect 110 559 111 563
rect 115 559 116 563
rect 110 558 116 559
rect 1238 563 1244 564
rect 1238 559 1239 563
rect 1243 559 1244 563
rect 1280 561 1282 593
rect 1560 584 1562 593
rect 1600 584 1602 593
rect 1640 584 1642 593
rect 1680 584 1682 593
rect 1720 584 1722 593
rect 1760 584 1762 593
rect 1808 584 1810 593
rect 1856 584 1858 593
rect 1912 584 1914 593
rect 1968 584 1970 593
rect 2032 584 2034 593
rect 2096 584 2098 593
rect 2168 584 2170 593
rect 2240 584 2242 593
rect 2312 584 2314 593
rect 2360 584 2362 593
rect 1558 583 1564 584
rect 1558 579 1559 583
rect 1563 579 1564 583
rect 1558 578 1564 579
rect 1598 583 1604 584
rect 1598 579 1599 583
rect 1603 579 1604 583
rect 1598 578 1604 579
rect 1638 583 1644 584
rect 1638 579 1639 583
rect 1643 579 1644 583
rect 1638 578 1644 579
rect 1678 583 1684 584
rect 1678 579 1679 583
rect 1683 579 1684 583
rect 1678 578 1684 579
rect 1718 583 1724 584
rect 1718 579 1719 583
rect 1723 579 1724 583
rect 1718 578 1724 579
rect 1758 583 1764 584
rect 1758 579 1759 583
rect 1763 579 1764 583
rect 1758 578 1764 579
rect 1806 583 1812 584
rect 1806 579 1807 583
rect 1811 579 1812 583
rect 1806 578 1812 579
rect 1854 583 1860 584
rect 1854 579 1855 583
rect 1859 579 1860 583
rect 1854 578 1860 579
rect 1910 583 1916 584
rect 1910 579 1911 583
rect 1915 579 1916 583
rect 1910 578 1916 579
rect 1966 583 1972 584
rect 1966 579 1967 583
rect 1971 579 1972 583
rect 1966 578 1972 579
rect 2030 583 2036 584
rect 2030 579 2031 583
rect 2035 579 2036 583
rect 2030 578 2036 579
rect 2094 583 2100 584
rect 2094 579 2095 583
rect 2099 579 2100 583
rect 2094 578 2100 579
rect 2166 583 2172 584
rect 2166 579 2167 583
rect 2171 579 2172 583
rect 2166 578 2172 579
rect 2238 583 2244 584
rect 2238 579 2239 583
rect 2243 579 2244 583
rect 2238 578 2244 579
rect 2310 583 2316 584
rect 2310 579 2311 583
rect 2315 579 2316 583
rect 2310 578 2316 579
rect 2358 583 2364 584
rect 2358 579 2359 583
rect 2363 579 2364 583
rect 2358 578 2364 579
rect 2408 561 2410 593
rect 1238 558 1244 559
rect 1278 560 1284 561
rect 112 547 114 558
rect 134 556 140 557
rect 134 552 135 556
rect 139 552 140 556
rect 134 551 140 552
rect 182 556 188 557
rect 182 552 183 556
rect 187 552 188 556
rect 182 551 188 552
rect 254 556 260 557
rect 254 552 255 556
rect 259 552 260 556
rect 254 551 260 552
rect 326 556 332 557
rect 326 552 327 556
rect 331 552 332 556
rect 326 551 332 552
rect 398 556 404 557
rect 398 552 399 556
rect 403 552 404 556
rect 398 551 404 552
rect 478 556 484 557
rect 478 552 479 556
rect 483 552 484 556
rect 478 551 484 552
rect 558 556 564 557
rect 558 552 559 556
rect 563 552 564 556
rect 558 551 564 552
rect 638 556 644 557
rect 638 552 639 556
rect 643 552 644 556
rect 638 551 644 552
rect 718 556 724 557
rect 718 552 719 556
rect 723 552 724 556
rect 718 551 724 552
rect 798 556 804 557
rect 798 552 799 556
rect 803 552 804 556
rect 798 551 804 552
rect 878 556 884 557
rect 878 552 879 556
rect 883 552 884 556
rect 878 551 884 552
rect 950 556 956 557
rect 950 552 951 556
rect 955 552 956 556
rect 950 551 956 552
rect 1014 556 1020 557
rect 1014 552 1015 556
rect 1019 552 1020 556
rect 1014 551 1020 552
rect 1078 556 1084 557
rect 1078 552 1079 556
rect 1083 552 1084 556
rect 1078 551 1084 552
rect 1142 556 1148 557
rect 1142 552 1143 556
rect 1147 552 1148 556
rect 1142 551 1148 552
rect 1190 556 1196 557
rect 1190 552 1191 556
rect 1195 552 1196 556
rect 1190 551 1196 552
rect 136 547 138 551
rect 184 547 186 551
rect 256 547 258 551
rect 328 547 330 551
rect 400 547 402 551
rect 480 547 482 551
rect 560 547 562 551
rect 640 547 642 551
rect 720 547 722 551
rect 800 547 802 551
rect 880 547 882 551
rect 952 547 954 551
rect 1016 547 1018 551
rect 1080 547 1082 551
rect 1144 547 1146 551
rect 1192 547 1194 551
rect 1240 547 1242 558
rect 1278 556 1279 560
rect 1283 556 1284 560
rect 1278 555 1284 556
rect 2406 560 2412 561
rect 2406 556 2407 560
rect 2411 556 2412 560
rect 2406 555 2412 556
rect 111 546 115 547
rect 111 541 115 542
rect 135 546 139 547
rect 135 541 139 542
rect 151 546 155 547
rect 151 541 155 542
rect 183 546 187 547
rect 183 541 187 542
rect 223 546 227 547
rect 223 541 227 542
rect 255 546 259 547
rect 255 541 259 542
rect 287 546 291 547
rect 287 541 291 542
rect 327 546 331 547
rect 327 541 331 542
rect 351 546 355 547
rect 351 541 355 542
rect 399 546 403 547
rect 399 541 403 542
rect 415 546 419 547
rect 415 541 419 542
rect 479 546 483 547
rect 479 541 483 542
rect 551 546 555 547
rect 551 541 555 542
rect 559 546 563 547
rect 559 541 563 542
rect 623 546 627 547
rect 623 541 627 542
rect 639 546 643 547
rect 639 541 643 542
rect 695 546 699 547
rect 695 541 699 542
rect 719 546 723 547
rect 719 541 723 542
rect 767 546 771 547
rect 767 541 771 542
rect 799 546 803 547
rect 799 541 803 542
rect 839 546 843 547
rect 839 541 843 542
rect 879 546 883 547
rect 879 541 883 542
rect 919 546 923 547
rect 919 541 923 542
rect 951 546 955 547
rect 951 541 955 542
rect 999 546 1003 547
rect 999 541 1003 542
rect 1015 546 1019 547
rect 1015 541 1019 542
rect 1079 546 1083 547
rect 1079 541 1083 542
rect 1143 546 1147 547
rect 1143 541 1147 542
rect 1191 546 1195 547
rect 1191 541 1195 542
rect 1239 546 1243 547
rect 1239 541 1243 542
rect 1278 543 1284 544
rect 112 534 114 541
rect 150 540 156 541
rect 150 536 151 540
rect 155 536 156 540
rect 150 535 156 536
rect 222 540 228 541
rect 222 536 223 540
rect 227 536 228 540
rect 222 535 228 536
rect 286 540 292 541
rect 286 536 287 540
rect 291 536 292 540
rect 286 535 292 536
rect 350 540 356 541
rect 350 536 351 540
rect 355 536 356 540
rect 350 535 356 536
rect 414 540 420 541
rect 414 536 415 540
rect 419 536 420 540
rect 414 535 420 536
rect 478 540 484 541
rect 478 536 479 540
rect 483 536 484 540
rect 478 535 484 536
rect 550 540 556 541
rect 550 536 551 540
rect 555 536 556 540
rect 550 535 556 536
rect 622 540 628 541
rect 622 536 623 540
rect 627 536 628 540
rect 622 535 628 536
rect 694 540 700 541
rect 694 536 695 540
rect 699 536 700 540
rect 694 535 700 536
rect 766 540 772 541
rect 766 536 767 540
rect 771 536 772 540
rect 766 535 772 536
rect 838 540 844 541
rect 838 536 839 540
rect 843 536 844 540
rect 838 535 844 536
rect 918 540 924 541
rect 918 536 919 540
rect 923 536 924 540
rect 918 535 924 536
rect 998 540 1004 541
rect 998 536 999 540
rect 1003 536 1004 540
rect 998 535 1004 536
rect 1078 540 1084 541
rect 1078 536 1079 540
rect 1083 536 1084 540
rect 1078 535 1084 536
rect 1240 534 1242 541
rect 1278 539 1279 543
rect 1283 539 1284 543
rect 1278 538 1284 539
rect 2406 543 2412 544
rect 2406 539 2407 543
rect 2411 539 2412 543
rect 2406 538 2412 539
rect 110 533 116 534
rect 110 529 111 533
rect 115 529 116 533
rect 110 528 116 529
rect 1238 533 1244 534
rect 1238 529 1239 533
rect 1243 529 1244 533
rect 1280 531 1282 538
rect 1558 536 1564 537
rect 1558 532 1559 536
rect 1563 532 1564 536
rect 1558 531 1564 532
rect 1598 536 1604 537
rect 1598 532 1599 536
rect 1603 532 1604 536
rect 1598 531 1604 532
rect 1638 536 1644 537
rect 1638 532 1639 536
rect 1643 532 1644 536
rect 1638 531 1644 532
rect 1678 536 1684 537
rect 1678 532 1679 536
rect 1683 532 1684 536
rect 1678 531 1684 532
rect 1718 536 1724 537
rect 1718 532 1719 536
rect 1723 532 1724 536
rect 1718 531 1724 532
rect 1758 536 1764 537
rect 1758 532 1759 536
rect 1763 532 1764 536
rect 1758 531 1764 532
rect 1806 536 1812 537
rect 1806 532 1807 536
rect 1811 532 1812 536
rect 1806 531 1812 532
rect 1854 536 1860 537
rect 1854 532 1855 536
rect 1859 532 1860 536
rect 1854 531 1860 532
rect 1910 536 1916 537
rect 1910 532 1911 536
rect 1915 532 1916 536
rect 1910 531 1916 532
rect 1966 536 1972 537
rect 1966 532 1967 536
rect 1971 532 1972 536
rect 1966 531 1972 532
rect 2030 536 2036 537
rect 2030 532 2031 536
rect 2035 532 2036 536
rect 2030 531 2036 532
rect 2094 536 2100 537
rect 2094 532 2095 536
rect 2099 532 2100 536
rect 2094 531 2100 532
rect 2166 536 2172 537
rect 2166 532 2167 536
rect 2171 532 2172 536
rect 2166 531 2172 532
rect 2238 536 2244 537
rect 2238 532 2239 536
rect 2243 532 2244 536
rect 2238 531 2244 532
rect 2310 536 2316 537
rect 2310 532 2311 536
rect 2315 532 2316 536
rect 2310 531 2316 532
rect 2358 536 2364 537
rect 2358 532 2359 536
rect 2363 532 2364 536
rect 2358 531 2364 532
rect 2408 531 2410 538
rect 1238 528 1244 529
rect 1279 530 1283 531
rect 1279 525 1283 526
rect 1407 530 1411 531
rect 1407 525 1411 526
rect 1447 530 1451 531
rect 1447 525 1451 526
rect 1487 530 1491 531
rect 1487 525 1491 526
rect 1535 530 1539 531
rect 1535 525 1539 526
rect 1559 530 1563 531
rect 1559 525 1563 526
rect 1591 530 1595 531
rect 1591 525 1595 526
rect 1599 530 1603 531
rect 1599 525 1603 526
rect 1639 530 1643 531
rect 1639 525 1643 526
rect 1647 530 1651 531
rect 1647 525 1651 526
rect 1679 530 1683 531
rect 1679 525 1683 526
rect 1711 530 1715 531
rect 1711 525 1715 526
rect 1719 530 1723 531
rect 1719 525 1723 526
rect 1759 530 1763 531
rect 1759 525 1763 526
rect 1783 530 1787 531
rect 1783 525 1787 526
rect 1807 530 1811 531
rect 1807 525 1811 526
rect 1855 530 1859 531
rect 1855 525 1859 526
rect 1863 530 1867 531
rect 1863 525 1867 526
rect 1911 530 1915 531
rect 1911 525 1915 526
rect 1943 530 1947 531
rect 1943 525 1947 526
rect 1967 530 1971 531
rect 1967 525 1971 526
rect 2023 530 2027 531
rect 2023 525 2027 526
rect 2031 530 2035 531
rect 2031 525 2035 526
rect 2095 530 2099 531
rect 2095 525 2099 526
rect 2103 530 2107 531
rect 2103 525 2107 526
rect 2167 530 2171 531
rect 2167 525 2171 526
rect 2191 530 2195 531
rect 2191 525 2195 526
rect 2239 530 2243 531
rect 2239 525 2243 526
rect 2287 530 2291 531
rect 2287 525 2291 526
rect 2311 530 2315 531
rect 2311 525 2315 526
rect 2359 530 2363 531
rect 2359 525 2363 526
rect 2407 530 2411 531
rect 2407 525 2411 526
rect 1280 518 1282 525
rect 1406 524 1412 525
rect 1406 520 1407 524
rect 1411 520 1412 524
rect 1406 519 1412 520
rect 1446 524 1452 525
rect 1446 520 1447 524
rect 1451 520 1452 524
rect 1446 519 1452 520
rect 1486 524 1492 525
rect 1486 520 1487 524
rect 1491 520 1492 524
rect 1486 519 1492 520
rect 1534 524 1540 525
rect 1534 520 1535 524
rect 1539 520 1540 524
rect 1534 519 1540 520
rect 1590 524 1596 525
rect 1590 520 1591 524
rect 1595 520 1596 524
rect 1590 519 1596 520
rect 1646 524 1652 525
rect 1646 520 1647 524
rect 1651 520 1652 524
rect 1646 519 1652 520
rect 1710 524 1716 525
rect 1710 520 1711 524
rect 1715 520 1716 524
rect 1710 519 1716 520
rect 1782 524 1788 525
rect 1782 520 1783 524
rect 1787 520 1788 524
rect 1782 519 1788 520
rect 1862 524 1868 525
rect 1862 520 1863 524
rect 1867 520 1868 524
rect 1862 519 1868 520
rect 1942 524 1948 525
rect 1942 520 1943 524
rect 1947 520 1948 524
rect 1942 519 1948 520
rect 2022 524 2028 525
rect 2022 520 2023 524
rect 2027 520 2028 524
rect 2022 519 2028 520
rect 2102 524 2108 525
rect 2102 520 2103 524
rect 2107 520 2108 524
rect 2102 519 2108 520
rect 2190 524 2196 525
rect 2190 520 2191 524
rect 2195 520 2196 524
rect 2190 519 2196 520
rect 2286 524 2292 525
rect 2286 520 2287 524
rect 2291 520 2292 524
rect 2286 519 2292 520
rect 2358 524 2364 525
rect 2358 520 2359 524
rect 2363 520 2364 524
rect 2358 519 2364 520
rect 2408 518 2410 525
rect 1278 517 1284 518
rect 110 516 116 517
rect 110 512 111 516
rect 115 512 116 516
rect 110 511 116 512
rect 1238 516 1244 517
rect 1238 512 1239 516
rect 1243 512 1244 516
rect 1278 513 1279 517
rect 1283 513 1284 517
rect 1278 512 1284 513
rect 2406 517 2412 518
rect 2406 513 2407 517
rect 2411 513 2412 517
rect 2406 512 2412 513
rect 1238 511 1244 512
rect 112 479 114 511
rect 150 493 156 494
rect 150 489 151 493
rect 155 489 156 493
rect 150 488 156 489
rect 222 493 228 494
rect 222 489 223 493
rect 227 489 228 493
rect 222 488 228 489
rect 286 493 292 494
rect 286 489 287 493
rect 291 489 292 493
rect 286 488 292 489
rect 350 493 356 494
rect 350 489 351 493
rect 355 489 356 493
rect 350 488 356 489
rect 414 493 420 494
rect 414 489 415 493
rect 419 489 420 493
rect 414 488 420 489
rect 478 493 484 494
rect 478 489 479 493
rect 483 489 484 493
rect 478 488 484 489
rect 550 493 556 494
rect 550 489 551 493
rect 555 489 556 493
rect 550 488 556 489
rect 622 493 628 494
rect 622 489 623 493
rect 627 489 628 493
rect 622 488 628 489
rect 694 493 700 494
rect 694 489 695 493
rect 699 489 700 493
rect 694 488 700 489
rect 766 493 772 494
rect 766 489 767 493
rect 771 489 772 493
rect 766 488 772 489
rect 838 493 844 494
rect 838 489 839 493
rect 843 489 844 493
rect 838 488 844 489
rect 918 493 924 494
rect 918 489 919 493
rect 923 489 924 493
rect 918 488 924 489
rect 998 493 1004 494
rect 998 489 999 493
rect 1003 489 1004 493
rect 998 488 1004 489
rect 1078 493 1084 494
rect 1078 489 1079 493
rect 1083 489 1084 493
rect 1078 488 1084 489
rect 152 479 154 488
rect 224 479 226 488
rect 288 479 290 488
rect 352 479 354 488
rect 416 479 418 488
rect 480 479 482 488
rect 552 479 554 488
rect 624 479 626 488
rect 696 479 698 488
rect 768 479 770 488
rect 840 479 842 488
rect 920 479 922 488
rect 1000 479 1002 488
rect 1080 479 1082 488
rect 1240 479 1242 511
rect 1278 500 1284 501
rect 1278 496 1279 500
rect 1283 496 1284 500
rect 1278 495 1284 496
rect 2406 500 2412 501
rect 2406 496 2407 500
rect 2411 496 2412 500
rect 2406 495 2412 496
rect 111 478 115 479
rect 111 473 115 474
rect 151 478 155 479
rect 151 473 155 474
rect 223 478 227 479
rect 223 473 227 474
rect 239 478 243 479
rect 239 473 243 474
rect 279 478 283 479
rect 279 473 283 474
rect 287 478 291 479
rect 287 473 291 474
rect 327 478 331 479
rect 327 473 331 474
rect 351 478 355 479
rect 351 473 355 474
rect 383 478 387 479
rect 383 473 387 474
rect 415 478 419 479
rect 415 473 419 474
rect 439 478 443 479
rect 439 473 443 474
rect 479 478 483 479
rect 479 473 483 474
rect 503 478 507 479
rect 503 473 507 474
rect 551 478 555 479
rect 551 473 555 474
rect 567 478 571 479
rect 567 473 571 474
rect 623 478 627 479
rect 623 473 627 474
rect 631 478 635 479
rect 631 473 635 474
rect 695 478 699 479
rect 695 473 699 474
rect 759 478 763 479
rect 759 473 763 474
rect 767 478 771 479
rect 767 473 771 474
rect 823 478 827 479
rect 823 473 827 474
rect 839 478 843 479
rect 839 473 843 474
rect 887 478 891 479
rect 887 473 891 474
rect 919 478 923 479
rect 919 473 923 474
rect 951 478 955 479
rect 951 473 955 474
rect 999 478 1003 479
rect 999 473 1003 474
rect 1015 478 1019 479
rect 1015 473 1019 474
rect 1079 478 1083 479
rect 1079 473 1083 474
rect 1239 478 1243 479
rect 1239 473 1243 474
rect 112 441 114 473
rect 240 464 242 473
rect 280 464 282 473
rect 328 464 330 473
rect 384 464 386 473
rect 440 464 442 473
rect 504 464 506 473
rect 568 464 570 473
rect 632 464 634 473
rect 696 464 698 473
rect 760 464 762 473
rect 824 464 826 473
rect 888 464 890 473
rect 952 464 954 473
rect 1016 464 1018 473
rect 238 463 244 464
rect 238 459 239 463
rect 243 459 244 463
rect 238 458 244 459
rect 278 463 284 464
rect 278 459 279 463
rect 283 459 284 463
rect 278 458 284 459
rect 326 463 332 464
rect 326 459 327 463
rect 331 459 332 463
rect 326 458 332 459
rect 382 463 388 464
rect 382 459 383 463
rect 387 459 388 463
rect 382 458 388 459
rect 438 463 444 464
rect 438 459 439 463
rect 443 459 444 463
rect 438 458 444 459
rect 502 463 508 464
rect 502 459 503 463
rect 507 459 508 463
rect 502 458 508 459
rect 566 463 572 464
rect 566 459 567 463
rect 571 459 572 463
rect 566 458 572 459
rect 630 463 636 464
rect 630 459 631 463
rect 635 459 636 463
rect 630 458 636 459
rect 694 463 700 464
rect 694 459 695 463
rect 699 459 700 463
rect 694 458 700 459
rect 758 463 764 464
rect 758 459 759 463
rect 763 459 764 463
rect 758 458 764 459
rect 822 463 828 464
rect 822 459 823 463
rect 827 459 828 463
rect 822 458 828 459
rect 886 463 892 464
rect 886 459 887 463
rect 891 459 892 463
rect 886 458 892 459
rect 950 463 956 464
rect 950 459 951 463
rect 955 459 956 463
rect 950 458 956 459
rect 1014 463 1020 464
rect 1014 459 1015 463
rect 1019 459 1020 463
rect 1014 458 1020 459
rect 1240 441 1242 473
rect 1280 463 1282 495
rect 1406 477 1412 478
rect 1406 473 1407 477
rect 1411 473 1412 477
rect 1406 472 1412 473
rect 1446 477 1452 478
rect 1446 473 1447 477
rect 1451 473 1452 477
rect 1446 472 1452 473
rect 1486 477 1492 478
rect 1486 473 1487 477
rect 1491 473 1492 477
rect 1486 472 1492 473
rect 1534 477 1540 478
rect 1534 473 1535 477
rect 1539 473 1540 477
rect 1534 472 1540 473
rect 1590 477 1596 478
rect 1590 473 1591 477
rect 1595 473 1596 477
rect 1590 472 1596 473
rect 1646 477 1652 478
rect 1646 473 1647 477
rect 1651 473 1652 477
rect 1646 472 1652 473
rect 1710 477 1716 478
rect 1710 473 1711 477
rect 1715 473 1716 477
rect 1710 472 1716 473
rect 1782 477 1788 478
rect 1782 473 1783 477
rect 1787 473 1788 477
rect 1782 472 1788 473
rect 1862 477 1868 478
rect 1862 473 1863 477
rect 1867 473 1868 477
rect 1862 472 1868 473
rect 1942 477 1948 478
rect 1942 473 1943 477
rect 1947 473 1948 477
rect 1942 472 1948 473
rect 2022 477 2028 478
rect 2022 473 2023 477
rect 2027 473 2028 477
rect 2022 472 2028 473
rect 2102 477 2108 478
rect 2102 473 2103 477
rect 2107 473 2108 477
rect 2102 472 2108 473
rect 2190 477 2196 478
rect 2190 473 2191 477
rect 2195 473 2196 477
rect 2190 472 2196 473
rect 2286 477 2292 478
rect 2286 473 2287 477
rect 2291 473 2292 477
rect 2286 472 2292 473
rect 2358 477 2364 478
rect 2358 473 2359 477
rect 2363 473 2364 477
rect 2358 472 2364 473
rect 1408 463 1410 472
rect 1448 463 1450 472
rect 1488 463 1490 472
rect 1536 463 1538 472
rect 1592 463 1594 472
rect 1648 463 1650 472
rect 1712 463 1714 472
rect 1784 463 1786 472
rect 1864 463 1866 472
rect 1944 463 1946 472
rect 2024 463 2026 472
rect 2104 463 2106 472
rect 2192 463 2194 472
rect 2288 463 2290 472
rect 2360 463 2362 472
rect 2408 463 2410 495
rect 1279 462 1283 463
rect 1279 457 1283 458
rect 1303 462 1307 463
rect 1303 457 1307 458
rect 1343 462 1347 463
rect 1343 457 1347 458
rect 1383 462 1387 463
rect 1383 457 1387 458
rect 1407 462 1411 463
rect 1407 457 1411 458
rect 1447 462 1451 463
rect 1447 457 1451 458
rect 1487 462 1491 463
rect 1487 457 1491 458
rect 1535 462 1539 463
rect 1535 457 1539 458
rect 1591 462 1595 463
rect 1591 457 1595 458
rect 1631 462 1635 463
rect 1631 457 1635 458
rect 1647 462 1651 463
rect 1647 457 1651 458
rect 1711 462 1715 463
rect 1711 457 1715 458
rect 1735 462 1739 463
rect 1735 457 1739 458
rect 1783 462 1787 463
rect 1783 457 1787 458
rect 1831 462 1835 463
rect 1831 457 1835 458
rect 1863 462 1867 463
rect 1863 457 1867 458
rect 1919 462 1923 463
rect 1919 457 1923 458
rect 1943 462 1947 463
rect 1943 457 1947 458
rect 1999 462 2003 463
rect 1999 457 2003 458
rect 2023 462 2027 463
rect 2023 457 2027 458
rect 2071 462 2075 463
rect 2071 457 2075 458
rect 2103 462 2107 463
rect 2103 457 2107 458
rect 2135 462 2139 463
rect 2135 457 2139 458
rect 2191 462 2195 463
rect 2191 457 2195 458
rect 2199 462 2203 463
rect 2199 457 2203 458
rect 2255 462 2259 463
rect 2255 457 2259 458
rect 2287 462 2291 463
rect 2287 457 2291 458
rect 2319 462 2323 463
rect 2319 457 2323 458
rect 2359 462 2363 463
rect 2359 457 2363 458
rect 2407 462 2411 463
rect 2407 457 2411 458
rect 110 440 116 441
rect 110 436 111 440
rect 115 436 116 440
rect 110 435 116 436
rect 1238 440 1244 441
rect 1238 436 1239 440
rect 1243 436 1244 440
rect 1238 435 1244 436
rect 1280 425 1282 457
rect 1304 448 1306 457
rect 1344 448 1346 457
rect 1384 448 1386 457
rect 1448 448 1450 457
rect 1536 448 1538 457
rect 1632 448 1634 457
rect 1736 448 1738 457
rect 1832 448 1834 457
rect 1920 448 1922 457
rect 2000 448 2002 457
rect 2072 448 2074 457
rect 2136 448 2138 457
rect 2200 448 2202 457
rect 2256 448 2258 457
rect 2320 448 2322 457
rect 2360 448 2362 457
rect 1302 447 1308 448
rect 1302 443 1303 447
rect 1307 443 1308 447
rect 1302 442 1308 443
rect 1342 447 1348 448
rect 1342 443 1343 447
rect 1347 443 1348 447
rect 1342 442 1348 443
rect 1382 447 1388 448
rect 1382 443 1383 447
rect 1387 443 1388 447
rect 1382 442 1388 443
rect 1446 447 1452 448
rect 1446 443 1447 447
rect 1451 443 1452 447
rect 1446 442 1452 443
rect 1534 447 1540 448
rect 1534 443 1535 447
rect 1539 443 1540 447
rect 1534 442 1540 443
rect 1630 447 1636 448
rect 1630 443 1631 447
rect 1635 443 1636 447
rect 1630 442 1636 443
rect 1734 447 1740 448
rect 1734 443 1735 447
rect 1739 443 1740 447
rect 1734 442 1740 443
rect 1830 447 1836 448
rect 1830 443 1831 447
rect 1835 443 1836 447
rect 1830 442 1836 443
rect 1918 447 1924 448
rect 1918 443 1919 447
rect 1923 443 1924 447
rect 1918 442 1924 443
rect 1998 447 2004 448
rect 1998 443 1999 447
rect 2003 443 2004 447
rect 1998 442 2004 443
rect 2070 447 2076 448
rect 2070 443 2071 447
rect 2075 443 2076 447
rect 2070 442 2076 443
rect 2134 447 2140 448
rect 2134 443 2135 447
rect 2139 443 2140 447
rect 2134 442 2140 443
rect 2198 447 2204 448
rect 2198 443 2199 447
rect 2203 443 2204 447
rect 2198 442 2204 443
rect 2254 447 2260 448
rect 2254 443 2255 447
rect 2259 443 2260 447
rect 2254 442 2260 443
rect 2318 447 2324 448
rect 2318 443 2319 447
rect 2323 443 2324 447
rect 2318 442 2324 443
rect 2358 447 2364 448
rect 2358 443 2359 447
rect 2363 443 2364 447
rect 2358 442 2364 443
rect 2408 425 2410 457
rect 1278 424 1284 425
rect 110 423 116 424
rect 110 419 111 423
rect 115 419 116 423
rect 110 418 116 419
rect 1238 423 1244 424
rect 1238 419 1239 423
rect 1243 419 1244 423
rect 1278 420 1279 424
rect 1283 420 1284 424
rect 1278 419 1284 420
rect 2406 424 2412 425
rect 2406 420 2407 424
rect 2411 420 2412 424
rect 2406 419 2412 420
rect 1238 418 1244 419
rect 112 407 114 418
rect 238 416 244 417
rect 238 412 239 416
rect 243 412 244 416
rect 238 411 244 412
rect 278 416 284 417
rect 278 412 279 416
rect 283 412 284 416
rect 278 411 284 412
rect 326 416 332 417
rect 326 412 327 416
rect 331 412 332 416
rect 326 411 332 412
rect 382 416 388 417
rect 382 412 383 416
rect 387 412 388 416
rect 382 411 388 412
rect 438 416 444 417
rect 438 412 439 416
rect 443 412 444 416
rect 438 411 444 412
rect 502 416 508 417
rect 502 412 503 416
rect 507 412 508 416
rect 502 411 508 412
rect 566 416 572 417
rect 566 412 567 416
rect 571 412 572 416
rect 566 411 572 412
rect 630 416 636 417
rect 630 412 631 416
rect 635 412 636 416
rect 630 411 636 412
rect 694 416 700 417
rect 694 412 695 416
rect 699 412 700 416
rect 694 411 700 412
rect 758 416 764 417
rect 758 412 759 416
rect 763 412 764 416
rect 758 411 764 412
rect 822 416 828 417
rect 822 412 823 416
rect 827 412 828 416
rect 822 411 828 412
rect 886 416 892 417
rect 886 412 887 416
rect 891 412 892 416
rect 886 411 892 412
rect 950 416 956 417
rect 950 412 951 416
rect 955 412 956 416
rect 950 411 956 412
rect 1014 416 1020 417
rect 1014 412 1015 416
rect 1019 412 1020 416
rect 1014 411 1020 412
rect 240 407 242 411
rect 280 407 282 411
rect 328 407 330 411
rect 384 407 386 411
rect 440 407 442 411
rect 504 407 506 411
rect 568 407 570 411
rect 632 407 634 411
rect 696 407 698 411
rect 760 407 762 411
rect 824 407 826 411
rect 888 407 890 411
rect 952 407 954 411
rect 1016 407 1018 411
rect 1240 407 1242 418
rect 1278 407 1284 408
rect 111 406 115 407
rect 111 401 115 402
rect 143 406 147 407
rect 143 401 147 402
rect 183 406 187 407
rect 183 401 187 402
rect 223 406 227 407
rect 223 401 227 402
rect 239 406 243 407
rect 239 401 243 402
rect 271 406 275 407
rect 271 401 275 402
rect 279 406 283 407
rect 279 401 283 402
rect 327 406 331 407
rect 327 401 331 402
rect 335 406 339 407
rect 335 401 339 402
rect 383 406 387 407
rect 383 401 387 402
rect 399 406 403 407
rect 399 401 403 402
rect 439 406 443 407
rect 439 401 443 402
rect 471 406 475 407
rect 471 401 475 402
rect 503 406 507 407
rect 503 401 507 402
rect 543 406 547 407
rect 543 401 547 402
rect 567 406 571 407
rect 567 401 571 402
rect 615 406 619 407
rect 615 401 619 402
rect 631 406 635 407
rect 631 401 635 402
rect 687 406 691 407
rect 687 401 691 402
rect 695 406 699 407
rect 695 401 699 402
rect 751 406 755 407
rect 751 401 755 402
rect 759 406 763 407
rect 759 401 763 402
rect 807 406 811 407
rect 807 401 811 402
rect 823 406 827 407
rect 823 401 827 402
rect 863 406 867 407
rect 863 401 867 402
rect 887 406 891 407
rect 887 401 891 402
rect 919 406 923 407
rect 919 401 923 402
rect 951 406 955 407
rect 951 401 955 402
rect 975 406 979 407
rect 975 401 979 402
rect 1015 406 1019 407
rect 1015 401 1019 402
rect 1031 406 1035 407
rect 1031 401 1035 402
rect 1239 406 1243 407
rect 1278 403 1279 407
rect 1283 403 1284 407
rect 1278 402 1284 403
rect 2406 407 2412 408
rect 2406 403 2407 407
rect 2411 403 2412 407
rect 2406 402 2412 403
rect 1239 401 1243 402
rect 112 394 114 401
rect 142 400 148 401
rect 142 396 143 400
rect 147 396 148 400
rect 142 395 148 396
rect 182 400 188 401
rect 182 396 183 400
rect 187 396 188 400
rect 182 395 188 396
rect 222 400 228 401
rect 222 396 223 400
rect 227 396 228 400
rect 222 395 228 396
rect 270 400 276 401
rect 270 396 271 400
rect 275 396 276 400
rect 270 395 276 396
rect 334 400 340 401
rect 334 396 335 400
rect 339 396 340 400
rect 334 395 340 396
rect 398 400 404 401
rect 398 396 399 400
rect 403 396 404 400
rect 398 395 404 396
rect 470 400 476 401
rect 470 396 471 400
rect 475 396 476 400
rect 470 395 476 396
rect 542 400 548 401
rect 542 396 543 400
rect 547 396 548 400
rect 542 395 548 396
rect 614 400 620 401
rect 614 396 615 400
rect 619 396 620 400
rect 614 395 620 396
rect 686 400 692 401
rect 686 396 687 400
rect 691 396 692 400
rect 686 395 692 396
rect 750 400 756 401
rect 750 396 751 400
rect 755 396 756 400
rect 750 395 756 396
rect 806 400 812 401
rect 806 396 807 400
rect 811 396 812 400
rect 806 395 812 396
rect 862 400 868 401
rect 862 396 863 400
rect 867 396 868 400
rect 862 395 868 396
rect 918 400 924 401
rect 918 396 919 400
rect 923 396 924 400
rect 918 395 924 396
rect 974 400 980 401
rect 974 396 975 400
rect 979 396 980 400
rect 974 395 980 396
rect 1030 400 1036 401
rect 1030 396 1031 400
rect 1035 396 1036 400
rect 1030 395 1036 396
rect 1240 394 1242 401
rect 1280 395 1282 402
rect 1302 400 1308 401
rect 1302 396 1303 400
rect 1307 396 1308 400
rect 1302 395 1308 396
rect 1342 400 1348 401
rect 1342 396 1343 400
rect 1347 396 1348 400
rect 1342 395 1348 396
rect 1382 400 1388 401
rect 1382 396 1383 400
rect 1387 396 1388 400
rect 1382 395 1388 396
rect 1446 400 1452 401
rect 1446 396 1447 400
rect 1451 396 1452 400
rect 1446 395 1452 396
rect 1534 400 1540 401
rect 1534 396 1535 400
rect 1539 396 1540 400
rect 1534 395 1540 396
rect 1630 400 1636 401
rect 1630 396 1631 400
rect 1635 396 1636 400
rect 1630 395 1636 396
rect 1734 400 1740 401
rect 1734 396 1735 400
rect 1739 396 1740 400
rect 1734 395 1740 396
rect 1830 400 1836 401
rect 1830 396 1831 400
rect 1835 396 1836 400
rect 1830 395 1836 396
rect 1918 400 1924 401
rect 1918 396 1919 400
rect 1923 396 1924 400
rect 1918 395 1924 396
rect 1998 400 2004 401
rect 1998 396 1999 400
rect 2003 396 2004 400
rect 1998 395 2004 396
rect 2070 400 2076 401
rect 2070 396 2071 400
rect 2075 396 2076 400
rect 2070 395 2076 396
rect 2134 400 2140 401
rect 2134 396 2135 400
rect 2139 396 2140 400
rect 2134 395 2140 396
rect 2198 400 2204 401
rect 2198 396 2199 400
rect 2203 396 2204 400
rect 2198 395 2204 396
rect 2254 400 2260 401
rect 2254 396 2255 400
rect 2259 396 2260 400
rect 2254 395 2260 396
rect 2318 400 2324 401
rect 2318 396 2319 400
rect 2323 396 2324 400
rect 2318 395 2324 396
rect 2358 400 2364 401
rect 2358 396 2359 400
rect 2363 396 2364 400
rect 2358 395 2364 396
rect 2408 395 2410 402
rect 1279 394 1283 395
rect 110 393 116 394
rect 110 389 111 393
rect 115 389 116 393
rect 110 388 116 389
rect 1238 393 1244 394
rect 1238 389 1239 393
rect 1243 389 1244 393
rect 1279 389 1283 390
rect 1303 394 1307 395
rect 1303 389 1307 390
rect 1343 394 1347 395
rect 1343 389 1347 390
rect 1359 394 1363 395
rect 1359 389 1363 390
rect 1383 394 1387 395
rect 1383 389 1387 390
rect 1399 394 1403 395
rect 1399 389 1403 390
rect 1439 394 1443 395
rect 1439 389 1443 390
rect 1447 394 1451 395
rect 1447 389 1451 390
rect 1487 394 1491 395
rect 1487 389 1491 390
rect 1535 394 1539 395
rect 1535 389 1539 390
rect 1543 394 1547 395
rect 1543 389 1547 390
rect 1607 394 1611 395
rect 1607 389 1611 390
rect 1631 394 1635 395
rect 1631 389 1635 390
rect 1679 394 1683 395
rect 1679 389 1683 390
rect 1735 394 1739 395
rect 1735 389 1739 390
rect 1759 394 1763 395
rect 1759 389 1763 390
rect 1831 394 1835 395
rect 1831 389 1835 390
rect 1839 394 1843 395
rect 1839 389 1843 390
rect 1919 394 1923 395
rect 1919 389 1923 390
rect 1999 394 2003 395
rect 1999 389 2003 390
rect 2071 394 2075 395
rect 2071 389 2075 390
rect 2079 394 2083 395
rect 2079 389 2083 390
rect 2135 394 2139 395
rect 2135 389 2139 390
rect 2159 394 2163 395
rect 2159 389 2163 390
rect 2199 394 2203 395
rect 2199 389 2203 390
rect 2247 394 2251 395
rect 2247 389 2251 390
rect 2255 394 2259 395
rect 2255 389 2259 390
rect 2319 394 2323 395
rect 2319 389 2323 390
rect 2335 394 2339 395
rect 2335 389 2339 390
rect 2359 394 2363 395
rect 2359 389 2363 390
rect 2407 394 2411 395
rect 2407 389 2411 390
rect 1238 388 1244 389
rect 1280 382 1282 389
rect 1358 388 1364 389
rect 1358 384 1359 388
rect 1363 384 1364 388
rect 1358 383 1364 384
rect 1398 388 1404 389
rect 1398 384 1399 388
rect 1403 384 1404 388
rect 1398 383 1404 384
rect 1438 388 1444 389
rect 1438 384 1439 388
rect 1443 384 1444 388
rect 1438 383 1444 384
rect 1486 388 1492 389
rect 1486 384 1487 388
rect 1491 384 1492 388
rect 1486 383 1492 384
rect 1542 388 1548 389
rect 1542 384 1543 388
rect 1547 384 1548 388
rect 1542 383 1548 384
rect 1606 388 1612 389
rect 1606 384 1607 388
rect 1611 384 1612 388
rect 1606 383 1612 384
rect 1678 388 1684 389
rect 1678 384 1679 388
rect 1683 384 1684 388
rect 1678 383 1684 384
rect 1758 388 1764 389
rect 1758 384 1759 388
rect 1763 384 1764 388
rect 1758 383 1764 384
rect 1838 388 1844 389
rect 1838 384 1839 388
rect 1843 384 1844 388
rect 1838 383 1844 384
rect 1918 388 1924 389
rect 1918 384 1919 388
rect 1923 384 1924 388
rect 1918 383 1924 384
rect 1998 388 2004 389
rect 1998 384 1999 388
rect 2003 384 2004 388
rect 1998 383 2004 384
rect 2078 388 2084 389
rect 2078 384 2079 388
rect 2083 384 2084 388
rect 2078 383 2084 384
rect 2158 388 2164 389
rect 2158 384 2159 388
rect 2163 384 2164 388
rect 2158 383 2164 384
rect 2246 388 2252 389
rect 2246 384 2247 388
rect 2251 384 2252 388
rect 2246 383 2252 384
rect 2334 388 2340 389
rect 2334 384 2335 388
rect 2339 384 2340 388
rect 2334 383 2340 384
rect 2408 382 2410 389
rect 1278 381 1284 382
rect 1278 377 1279 381
rect 1283 377 1284 381
rect 110 376 116 377
rect 110 372 111 376
rect 115 372 116 376
rect 110 371 116 372
rect 1238 376 1244 377
rect 1278 376 1284 377
rect 2406 381 2412 382
rect 2406 377 2407 381
rect 2411 377 2412 381
rect 2406 376 2412 377
rect 1238 372 1239 376
rect 1243 372 1244 376
rect 1238 371 1244 372
rect 112 331 114 371
rect 142 353 148 354
rect 142 349 143 353
rect 147 349 148 353
rect 142 348 148 349
rect 182 353 188 354
rect 182 349 183 353
rect 187 349 188 353
rect 182 348 188 349
rect 222 353 228 354
rect 222 349 223 353
rect 227 349 228 353
rect 222 348 228 349
rect 270 353 276 354
rect 270 349 271 353
rect 275 349 276 353
rect 270 348 276 349
rect 334 353 340 354
rect 334 349 335 353
rect 339 349 340 353
rect 334 348 340 349
rect 398 353 404 354
rect 398 349 399 353
rect 403 349 404 353
rect 398 348 404 349
rect 470 353 476 354
rect 470 349 471 353
rect 475 349 476 353
rect 470 348 476 349
rect 542 353 548 354
rect 542 349 543 353
rect 547 349 548 353
rect 542 348 548 349
rect 614 353 620 354
rect 614 349 615 353
rect 619 349 620 353
rect 614 348 620 349
rect 686 353 692 354
rect 686 349 687 353
rect 691 349 692 353
rect 686 348 692 349
rect 750 353 756 354
rect 750 349 751 353
rect 755 349 756 353
rect 750 348 756 349
rect 806 353 812 354
rect 806 349 807 353
rect 811 349 812 353
rect 806 348 812 349
rect 862 353 868 354
rect 862 349 863 353
rect 867 349 868 353
rect 862 348 868 349
rect 918 353 924 354
rect 918 349 919 353
rect 923 349 924 353
rect 918 348 924 349
rect 974 353 980 354
rect 974 349 975 353
rect 979 349 980 353
rect 974 348 980 349
rect 1030 353 1036 354
rect 1030 349 1031 353
rect 1035 349 1036 353
rect 1030 348 1036 349
rect 144 331 146 348
rect 184 331 186 348
rect 224 331 226 348
rect 272 331 274 348
rect 336 331 338 348
rect 400 331 402 348
rect 472 331 474 348
rect 544 331 546 348
rect 616 331 618 348
rect 688 331 690 348
rect 752 331 754 348
rect 808 331 810 348
rect 864 331 866 348
rect 920 331 922 348
rect 976 331 978 348
rect 1032 331 1034 348
rect 1240 331 1242 371
rect 1278 364 1284 365
rect 1278 360 1279 364
rect 1283 360 1284 364
rect 1278 359 1284 360
rect 2406 364 2412 365
rect 2406 360 2407 364
rect 2411 360 2412 364
rect 2406 359 2412 360
rect 111 330 115 331
rect 111 325 115 326
rect 135 330 139 331
rect 135 325 139 326
rect 143 330 147 331
rect 143 325 147 326
rect 175 330 179 331
rect 175 325 179 326
rect 183 330 187 331
rect 183 325 187 326
rect 215 330 219 331
rect 215 325 219 326
rect 223 330 227 331
rect 223 325 227 326
rect 255 330 259 331
rect 255 325 259 326
rect 271 330 275 331
rect 271 325 275 326
rect 295 330 299 331
rect 295 325 299 326
rect 335 330 339 331
rect 335 325 339 326
rect 391 330 395 331
rect 391 325 395 326
rect 399 330 403 331
rect 399 325 403 326
rect 447 330 451 331
rect 447 325 451 326
rect 471 330 475 331
rect 471 325 475 326
rect 495 330 499 331
rect 495 325 499 326
rect 543 330 547 331
rect 543 325 547 326
rect 591 330 595 331
rect 591 325 595 326
rect 615 330 619 331
rect 615 325 619 326
rect 639 330 643 331
rect 639 325 643 326
rect 687 330 691 331
rect 687 325 691 326
rect 735 330 739 331
rect 735 325 739 326
rect 751 330 755 331
rect 751 325 755 326
rect 783 330 787 331
rect 783 325 787 326
rect 807 330 811 331
rect 807 325 811 326
rect 839 330 843 331
rect 839 325 843 326
rect 863 330 867 331
rect 863 325 867 326
rect 919 330 923 331
rect 919 325 923 326
rect 975 330 979 331
rect 975 325 979 326
rect 1031 330 1035 331
rect 1031 325 1035 326
rect 1239 330 1243 331
rect 1239 325 1243 326
rect 112 293 114 325
rect 136 316 138 325
rect 176 316 178 325
rect 216 316 218 325
rect 256 316 258 325
rect 296 316 298 325
rect 336 316 338 325
rect 392 316 394 325
rect 448 316 450 325
rect 496 316 498 325
rect 544 316 546 325
rect 592 316 594 325
rect 640 316 642 325
rect 688 316 690 325
rect 736 316 738 325
rect 784 316 786 325
rect 840 316 842 325
rect 134 315 140 316
rect 134 311 135 315
rect 139 311 140 315
rect 134 310 140 311
rect 174 315 180 316
rect 174 311 175 315
rect 179 311 180 315
rect 174 310 180 311
rect 214 315 220 316
rect 214 311 215 315
rect 219 311 220 315
rect 214 310 220 311
rect 254 315 260 316
rect 254 311 255 315
rect 259 311 260 315
rect 254 310 260 311
rect 294 315 300 316
rect 294 311 295 315
rect 299 311 300 315
rect 294 310 300 311
rect 334 315 340 316
rect 334 311 335 315
rect 339 311 340 315
rect 334 310 340 311
rect 390 315 396 316
rect 390 311 391 315
rect 395 311 396 315
rect 390 310 396 311
rect 446 315 452 316
rect 446 311 447 315
rect 451 311 452 315
rect 446 310 452 311
rect 494 315 500 316
rect 494 311 495 315
rect 499 311 500 315
rect 494 310 500 311
rect 542 315 548 316
rect 542 311 543 315
rect 547 311 548 315
rect 542 310 548 311
rect 590 315 596 316
rect 590 311 591 315
rect 595 311 596 315
rect 590 310 596 311
rect 638 315 644 316
rect 638 311 639 315
rect 643 311 644 315
rect 638 310 644 311
rect 686 315 692 316
rect 686 311 687 315
rect 691 311 692 315
rect 686 310 692 311
rect 734 315 740 316
rect 734 311 735 315
rect 739 311 740 315
rect 734 310 740 311
rect 782 315 788 316
rect 782 311 783 315
rect 787 311 788 315
rect 782 310 788 311
rect 838 315 844 316
rect 838 311 839 315
rect 843 311 844 315
rect 838 310 844 311
rect 1240 293 1242 325
rect 1280 319 1282 359
rect 1358 341 1364 342
rect 1358 337 1359 341
rect 1363 337 1364 341
rect 1358 336 1364 337
rect 1398 341 1404 342
rect 1398 337 1399 341
rect 1403 337 1404 341
rect 1398 336 1404 337
rect 1438 341 1444 342
rect 1438 337 1439 341
rect 1443 337 1444 341
rect 1438 336 1444 337
rect 1486 341 1492 342
rect 1486 337 1487 341
rect 1491 337 1492 341
rect 1486 336 1492 337
rect 1542 341 1548 342
rect 1542 337 1543 341
rect 1547 337 1548 341
rect 1542 336 1548 337
rect 1606 341 1612 342
rect 1606 337 1607 341
rect 1611 337 1612 341
rect 1606 336 1612 337
rect 1678 341 1684 342
rect 1678 337 1679 341
rect 1683 337 1684 341
rect 1678 336 1684 337
rect 1758 341 1764 342
rect 1758 337 1759 341
rect 1763 337 1764 341
rect 1758 336 1764 337
rect 1838 341 1844 342
rect 1838 337 1839 341
rect 1843 337 1844 341
rect 1838 336 1844 337
rect 1918 341 1924 342
rect 1918 337 1919 341
rect 1923 337 1924 341
rect 1918 336 1924 337
rect 1998 341 2004 342
rect 1998 337 1999 341
rect 2003 337 2004 341
rect 1998 336 2004 337
rect 2078 341 2084 342
rect 2078 337 2079 341
rect 2083 337 2084 341
rect 2078 336 2084 337
rect 2158 341 2164 342
rect 2158 337 2159 341
rect 2163 337 2164 341
rect 2158 336 2164 337
rect 2246 341 2252 342
rect 2246 337 2247 341
rect 2251 337 2252 341
rect 2246 336 2252 337
rect 2334 341 2340 342
rect 2334 337 2335 341
rect 2339 337 2340 341
rect 2334 336 2340 337
rect 1360 319 1362 336
rect 1400 319 1402 336
rect 1440 319 1442 336
rect 1488 319 1490 336
rect 1544 319 1546 336
rect 1608 319 1610 336
rect 1680 319 1682 336
rect 1760 319 1762 336
rect 1840 319 1842 336
rect 1920 319 1922 336
rect 2000 319 2002 336
rect 2080 319 2082 336
rect 2160 319 2162 336
rect 2248 319 2250 336
rect 2336 319 2338 336
rect 2408 319 2410 359
rect 1279 318 1283 319
rect 1279 313 1283 314
rect 1359 318 1363 319
rect 1359 313 1363 314
rect 1399 318 1403 319
rect 1399 313 1403 314
rect 1439 318 1443 319
rect 1439 313 1443 314
rect 1487 318 1491 319
rect 1487 313 1491 314
rect 1511 318 1515 319
rect 1511 313 1515 314
rect 1543 318 1547 319
rect 1543 313 1547 314
rect 1551 318 1555 319
rect 1551 313 1555 314
rect 1591 318 1595 319
rect 1591 313 1595 314
rect 1607 318 1611 319
rect 1607 313 1611 314
rect 1631 318 1635 319
rect 1631 313 1635 314
rect 1671 318 1675 319
rect 1671 313 1675 314
rect 1679 318 1683 319
rect 1679 313 1683 314
rect 1711 318 1715 319
rect 1711 313 1715 314
rect 1751 318 1755 319
rect 1751 313 1755 314
rect 1759 318 1763 319
rect 1759 313 1763 314
rect 1791 318 1795 319
rect 1791 313 1795 314
rect 1839 318 1843 319
rect 1839 313 1843 314
rect 1903 318 1907 319
rect 1903 313 1907 314
rect 1919 318 1923 319
rect 1919 313 1923 314
rect 1967 318 1971 319
rect 1967 313 1971 314
rect 1999 318 2003 319
rect 1999 313 2003 314
rect 2039 318 2043 319
rect 2039 313 2043 314
rect 2079 318 2083 319
rect 2079 313 2083 314
rect 2119 318 2123 319
rect 2119 313 2123 314
rect 2159 318 2163 319
rect 2159 313 2163 314
rect 2199 318 2203 319
rect 2199 313 2203 314
rect 2247 318 2251 319
rect 2247 313 2251 314
rect 2279 318 2283 319
rect 2279 313 2283 314
rect 2335 318 2339 319
rect 2335 313 2339 314
rect 2359 318 2363 319
rect 2359 313 2363 314
rect 2407 318 2411 319
rect 2407 313 2411 314
rect 110 292 116 293
rect 110 288 111 292
rect 115 288 116 292
rect 110 287 116 288
rect 1238 292 1244 293
rect 1238 288 1239 292
rect 1243 288 1244 292
rect 1238 287 1244 288
rect 1280 281 1282 313
rect 1512 304 1514 313
rect 1552 304 1554 313
rect 1592 304 1594 313
rect 1632 304 1634 313
rect 1672 304 1674 313
rect 1712 304 1714 313
rect 1752 304 1754 313
rect 1792 304 1794 313
rect 1840 304 1842 313
rect 1904 304 1906 313
rect 1968 304 1970 313
rect 2040 304 2042 313
rect 2120 304 2122 313
rect 2200 304 2202 313
rect 2280 304 2282 313
rect 2360 304 2362 313
rect 1510 303 1516 304
rect 1510 299 1511 303
rect 1515 299 1516 303
rect 1510 298 1516 299
rect 1550 303 1556 304
rect 1550 299 1551 303
rect 1555 299 1556 303
rect 1550 298 1556 299
rect 1590 303 1596 304
rect 1590 299 1591 303
rect 1595 299 1596 303
rect 1590 298 1596 299
rect 1630 303 1636 304
rect 1630 299 1631 303
rect 1635 299 1636 303
rect 1630 298 1636 299
rect 1670 303 1676 304
rect 1670 299 1671 303
rect 1675 299 1676 303
rect 1670 298 1676 299
rect 1710 303 1716 304
rect 1710 299 1711 303
rect 1715 299 1716 303
rect 1710 298 1716 299
rect 1750 303 1756 304
rect 1750 299 1751 303
rect 1755 299 1756 303
rect 1750 298 1756 299
rect 1790 303 1796 304
rect 1790 299 1791 303
rect 1795 299 1796 303
rect 1790 298 1796 299
rect 1838 303 1844 304
rect 1838 299 1839 303
rect 1843 299 1844 303
rect 1838 298 1844 299
rect 1902 303 1908 304
rect 1902 299 1903 303
rect 1907 299 1908 303
rect 1902 298 1908 299
rect 1966 303 1972 304
rect 1966 299 1967 303
rect 1971 299 1972 303
rect 1966 298 1972 299
rect 2038 303 2044 304
rect 2038 299 2039 303
rect 2043 299 2044 303
rect 2038 298 2044 299
rect 2118 303 2124 304
rect 2118 299 2119 303
rect 2123 299 2124 303
rect 2118 298 2124 299
rect 2198 303 2204 304
rect 2198 299 2199 303
rect 2203 299 2204 303
rect 2198 298 2204 299
rect 2278 303 2284 304
rect 2278 299 2279 303
rect 2283 299 2284 303
rect 2278 298 2284 299
rect 2358 303 2364 304
rect 2358 299 2359 303
rect 2363 299 2364 303
rect 2358 298 2364 299
rect 2408 281 2410 313
rect 1278 280 1284 281
rect 1278 276 1279 280
rect 1283 276 1284 280
rect 110 275 116 276
rect 110 271 111 275
rect 115 271 116 275
rect 110 270 116 271
rect 1238 275 1244 276
rect 1278 275 1284 276
rect 2406 280 2412 281
rect 2406 276 2407 280
rect 2411 276 2412 280
rect 2406 275 2412 276
rect 1238 271 1239 275
rect 1243 271 1244 275
rect 1238 270 1244 271
rect 112 255 114 270
rect 134 268 140 269
rect 134 264 135 268
rect 139 264 140 268
rect 134 263 140 264
rect 174 268 180 269
rect 174 264 175 268
rect 179 264 180 268
rect 174 263 180 264
rect 214 268 220 269
rect 214 264 215 268
rect 219 264 220 268
rect 214 263 220 264
rect 254 268 260 269
rect 254 264 255 268
rect 259 264 260 268
rect 254 263 260 264
rect 294 268 300 269
rect 294 264 295 268
rect 299 264 300 268
rect 294 263 300 264
rect 334 268 340 269
rect 334 264 335 268
rect 339 264 340 268
rect 334 263 340 264
rect 390 268 396 269
rect 390 264 391 268
rect 395 264 396 268
rect 390 263 396 264
rect 446 268 452 269
rect 446 264 447 268
rect 451 264 452 268
rect 446 263 452 264
rect 494 268 500 269
rect 494 264 495 268
rect 499 264 500 268
rect 494 263 500 264
rect 542 268 548 269
rect 542 264 543 268
rect 547 264 548 268
rect 542 263 548 264
rect 590 268 596 269
rect 590 264 591 268
rect 595 264 596 268
rect 590 263 596 264
rect 638 268 644 269
rect 638 264 639 268
rect 643 264 644 268
rect 638 263 644 264
rect 686 268 692 269
rect 686 264 687 268
rect 691 264 692 268
rect 686 263 692 264
rect 734 268 740 269
rect 734 264 735 268
rect 739 264 740 268
rect 734 263 740 264
rect 782 268 788 269
rect 782 264 783 268
rect 787 264 788 268
rect 782 263 788 264
rect 838 268 844 269
rect 838 264 839 268
rect 843 264 844 268
rect 838 263 844 264
rect 136 255 138 263
rect 176 255 178 263
rect 216 255 218 263
rect 256 255 258 263
rect 296 255 298 263
rect 336 255 338 263
rect 392 255 394 263
rect 448 255 450 263
rect 496 255 498 263
rect 544 255 546 263
rect 592 255 594 263
rect 640 255 642 263
rect 688 255 690 263
rect 736 255 738 263
rect 784 255 786 263
rect 840 255 842 263
rect 1240 255 1242 270
rect 1278 263 1284 264
rect 1278 259 1279 263
rect 1283 259 1284 263
rect 1278 258 1284 259
rect 2406 263 2412 264
rect 2406 259 2407 263
rect 2411 259 2412 263
rect 2406 258 2412 259
rect 111 254 115 255
rect 111 249 115 250
rect 135 254 139 255
rect 135 249 139 250
rect 175 254 179 255
rect 175 249 179 250
rect 215 254 219 255
rect 215 249 219 250
rect 223 254 227 255
rect 223 249 227 250
rect 255 254 259 255
rect 255 249 259 250
rect 295 254 299 255
rect 295 249 299 250
rect 311 254 315 255
rect 311 249 315 250
rect 335 254 339 255
rect 335 249 339 250
rect 391 254 395 255
rect 391 249 395 250
rect 447 254 451 255
rect 447 249 451 250
rect 463 254 467 255
rect 463 249 467 250
rect 495 254 499 255
rect 495 249 499 250
rect 527 254 531 255
rect 527 249 531 250
rect 543 254 547 255
rect 543 249 547 250
rect 591 254 595 255
rect 591 249 595 250
rect 639 254 643 255
rect 639 249 643 250
rect 647 254 651 255
rect 647 249 651 250
rect 687 254 691 255
rect 687 249 691 250
rect 695 254 699 255
rect 695 249 699 250
rect 735 254 739 255
rect 735 249 739 250
rect 783 254 787 255
rect 783 249 787 250
rect 831 254 835 255
rect 831 249 835 250
rect 839 254 843 255
rect 839 249 843 250
rect 879 254 883 255
rect 879 249 883 250
rect 927 254 931 255
rect 927 249 931 250
rect 975 254 979 255
rect 975 249 979 250
rect 1023 254 1027 255
rect 1023 249 1027 250
rect 1239 254 1243 255
rect 1239 249 1243 250
rect 112 242 114 249
rect 134 248 140 249
rect 134 244 135 248
rect 139 244 140 248
rect 134 243 140 244
rect 222 248 228 249
rect 222 244 223 248
rect 227 244 228 248
rect 222 243 228 244
rect 310 248 316 249
rect 310 244 311 248
rect 315 244 316 248
rect 310 243 316 244
rect 390 248 396 249
rect 390 244 391 248
rect 395 244 396 248
rect 390 243 396 244
rect 462 248 468 249
rect 462 244 463 248
rect 467 244 468 248
rect 462 243 468 244
rect 526 248 532 249
rect 526 244 527 248
rect 531 244 532 248
rect 526 243 532 244
rect 590 248 596 249
rect 590 244 591 248
rect 595 244 596 248
rect 590 243 596 244
rect 646 248 652 249
rect 646 244 647 248
rect 651 244 652 248
rect 646 243 652 244
rect 694 248 700 249
rect 694 244 695 248
rect 699 244 700 248
rect 694 243 700 244
rect 734 248 740 249
rect 734 244 735 248
rect 739 244 740 248
rect 734 243 740 244
rect 782 248 788 249
rect 782 244 783 248
rect 787 244 788 248
rect 782 243 788 244
rect 830 248 836 249
rect 830 244 831 248
rect 835 244 836 248
rect 830 243 836 244
rect 878 248 884 249
rect 878 244 879 248
rect 883 244 884 248
rect 878 243 884 244
rect 926 248 932 249
rect 926 244 927 248
rect 931 244 932 248
rect 926 243 932 244
rect 974 248 980 249
rect 974 244 975 248
rect 979 244 980 248
rect 974 243 980 244
rect 1022 248 1028 249
rect 1022 244 1023 248
rect 1027 244 1028 248
rect 1022 243 1028 244
rect 1240 242 1242 249
rect 1280 247 1282 258
rect 1510 256 1516 257
rect 1510 252 1511 256
rect 1515 252 1516 256
rect 1510 251 1516 252
rect 1550 256 1556 257
rect 1550 252 1551 256
rect 1555 252 1556 256
rect 1550 251 1556 252
rect 1590 256 1596 257
rect 1590 252 1591 256
rect 1595 252 1596 256
rect 1590 251 1596 252
rect 1630 256 1636 257
rect 1630 252 1631 256
rect 1635 252 1636 256
rect 1630 251 1636 252
rect 1670 256 1676 257
rect 1670 252 1671 256
rect 1675 252 1676 256
rect 1670 251 1676 252
rect 1710 256 1716 257
rect 1710 252 1711 256
rect 1715 252 1716 256
rect 1710 251 1716 252
rect 1750 256 1756 257
rect 1750 252 1751 256
rect 1755 252 1756 256
rect 1750 251 1756 252
rect 1790 256 1796 257
rect 1790 252 1791 256
rect 1795 252 1796 256
rect 1790 251 1796 252
rect 1838 256 1844 257
rect 1838 252 1839 256
rect 1843 252 1844 256
rect 1838 251 1844 252
rect 1902 256 1908 257
rect 1902 252 1903 256
rect 1907 252 1908 256
rect 1902 251 1908 252
rect 1966 256 1972 257
rect 1966 252 1967 256
rect 1971 252 1972 256
rect 1966 251 1972 252
rect 2038 256 2044 257
rect 2038 252 2039 256
rect 2043 252 2044 256
rect 2038 251 2044 252
rect 2118 256 2124 257
rect 2118 252 2119 256
rect 2123 252 2124 256
rect 2118 251 2124 252
rect 2198 256 2204 257
rect 2198 252 2199 256
rect 2203 252 2204 256
rect 2198 251 2204 252
rect 2278 256 2284 257
rect 2278 252 2279 256
rect 2283 252 2284 256
rect 2278 251 2284 252
rect 2358 256 2364 257
rect 2358 252 2359 256
rect 2363 252 2364 256
rect 2358 251 2364 252
rect 1512 247 1514 251
rect 1552 247 1554 251
rect 1592 247 1594 251
rect 1632 247 1634 251
rect 1672 247 1674 251
rect 1712 247 1714 251
rect 1752 247 1754 251
rect 1792 247 1794 251
rect 1840 247 1842 251
rect 1904 247 1906 251
rect 1968 247 1970 251
rect 2040 247 2042 251
rect 2120 247 2122 251
rect 2200 247 2202 251
rect 2280 247 2282 251
rect 2360 247 2362 251
rect 2408 247 2410 258
rect 1279 246 1283 247
rect 110 241 116 242
rect 110 237 111 241
rect 115 237 116 241
rect 110 236 116 237
rect 1238 241 1244 242
rect 1279 241 1283 242
rect 1367 246 1371 247
rect 1367 241 1371 242
rect 1407 246 1411 247
rect 1407 241 1411 242
rect 1455 246 1459 247
rect 1455 241 1459 242
rect 1511 246 1515 247
rect 1511 241 1515 242
rect 1551 246 1555 247
rect 1551 241 1555 242
rect 1567 246 1571 247
rect 1567 241 1571 242
rect 1591 246 1595 247
rect 1591 241 1595 242
rect 1631 246 1635 247
rect 1631 241 1635 242
rect 1671 246 1675 247
rect 1671 241 1675 242
rect 1703 246 1707 247
rect 1703 241 1707 242
rect 1711 246 1715 247
rect 1711 241 1715 242
rect 1751 246 1755 247
rect 1751 241 1755 242
rect 1775 246 1779 247
rect 1775 241 1779 242
rect 1791 246 1795 247
rect 1791 241 1795 242
rect 1839 246 1843 247
rect 1839 241 1843 242
rect 1855 246 1859 247
rect 1855 241 1859 242
rect 1903 246 1907 247
rect 1903 241 1907 242
rect 1943 246 1947 247
rect 1943 241 1947 242
rect 1967 246 1971 247
rect 1967 241 1971 242
rect 2031 246 2035 247
rect 2031 241 2035 242
rect 2039 246 2043 247
rect 2039 241 2043 242
rect 2119 246 2123 247
rect 2119 241 2123 242
rect 2199 246 2203 247
rect 2199 241 2203 242
rect 2207 246 2211 247
rect 2207 241 2211 242
rect 2279 246 2283 247
rect 2279 241 2283 242
rect 2295 246 2299 247
rect 2295 241 2299 242
rect 2359 246 2363 247
rect 2359 241 2363 242
rect 2407 246 2411 247
rect 2407 241 2411 242
rect 1238 237 1239 241
rect 1243 237 1244 241
rect 1238 236 1244 237
rect 1280 234 1282 241
rect 1366 240 1372 241
rect 1366 236 1367 240
rect 1371 236 1372 240
rect 1366 235 1372 236
rect 1406 240 1412 241
rect 1406 236 1407 240
rect 1411 236 1412 240
rect 1406 235 1412 236
rect 1454 240 1460 241
rect 1454 236 1455 240
rect 1459 236 1460 240
rect 1454 235 1460 236
rect 1510 240 1516 241
rect 1510 236 1511 240
rect 1515 236 1516 240
rect 1510 235 1516 236
rect 1566 240 1572 241
rect 1566 236 1567 240
rect 1571 236 1572 240
rect 1566 235 1572 236
rect 1630 240 1636 241
rect 1630 236 1631 240
rect 1635 236 1636 240
rect 1630 235 1636 236
rect 1702 240 1708 241
rect 1702 236 1703 240
rect 1707 236 1708 240
rect 1702 235 1708 236
rect 1774 240 1780 241
rect 1774 236 1775 240
rect 1779 236 1780 240
rect 1774 235 1780 236
rect 1854 240 1860 241
rect 1854 236 1855 240
rect 1859 236 1860 240
rect 1854 235 1860 236
rect 1942 240 1948 241
rect 1942 236 1943 240
rect 1947 236 1948 240
rect 1942 235 1948 236
rect 2030 240 2036 241
rect 2030 236 2031 240
rect 2035 236 2036 240
rect 2030 235 2036 236
rect 2118 240 2124 241
rect 2118 236 2119 240
rect 2123 236 2124 240
rect 2118 235 2124 236
rect 2206 240 2212 241
rect 2206 236 2207 240
rect 2211 236 2212 240
rect 2206 235 2212 236
rect 2294 240 2300 241
rect 2294 236 2295 240
rect 2299 236 2300 240
rect 2294 235 2300 236
rect 2358 240 2364 241
rect 2358 236 2359 240
rect 2363 236 2364 240
rect 2358 235 2364 236
rect 2408 234 2410 241
rect 1278 233 1284 234
rect 1278 229 1279 233
rect 1283 229 1284 233
rect 1278 228 1284 229
rect 2406 233 2412 234
rect 2406 229 2407 233
rect 2411 229 2412 233
rect 2406 228 2412 229
rect 110 224 116 225
rect 110 220 111 224
rect 115 220 116 224
rect 110 219 116 220
rect 1238 224 1244 225
rect 1238 220 1239 224
rect 1243 220 1244 224
rect 1238 219 1244 220
rect 112 155 114 219
rect 134 201 140 202
rect 134 197 135 201
rect 139 197 140 201
rect 134 196 140 197
rect 222 201 228 202
rect 222 197 223 201
rect 227 197 228 201
rect 222 196 228 197
rect 310 201 316 202
rect 310 197 311 201
rect 315 197 316 201
rect 310 196 316 197
rect 390 201 396 202
rect 390 197 391 201
rect 395 197 396 201
rect 390 196 396 197
rect 462 201 468 202
rect 462 197 463 201
rect 467 197 468 201
rect 462 196 468 197
rect 526 201 532 202
rect 526 197 527 201
rect 531 197 532 201
rect 526 196 532 197
rect 590 201 596 202
rect 590 197 591 201
rect 595 197 596 201
rect 590 196 596 197
rect 646 201 652 202
rect 646 197 647 201
rect 651 197 652 201
rect 646 196 652 197
rect 694 201 700 202
rect 694 197 695 201
rect 699 197 700 201
rect 694 196 700 197
rect 734 201 740 202
rect 734 197 735 201
rect 739 197 740 201
rect 734 196 740 197
rect 782 201 788 202
rect 782 197 783 201
rect 787 197 788 201
rect 782 196 788 197
rect 830 201 836 202
rect 830 197 831 201
rect 835 197 836 201
rect 830 196 836 197
rect 878 201 884 202
rect 878 197 879 201
rect 883 197 884 201
rect 878 196 884 197
rect 926 201 932 202
rect 926 197 927 201
rect 931 197 932 201
rect 926 196 932 197
rect 974 201 980 202
rect 974 197 975 201
rect 979 197 980 201
rect 974 196 980 197
rect 1022 201 1028 202
rect 1022 197 1023 201
rect 1027 197 1028 201
rect 1022 196 1028 197
rect 136 155 138 196
rect 224 155 226 196
rect 312 155 314 196
rect 392 155 394 196
rect 464 155 466 196
rect 528 155 530 196
rect 592 155 594 196
rect 648 155 650 196
rect 696 155 698 196
rect 736 155 738 196
rect 784 155 786 196
rect 832 155 834 196
rect 880 155 882 196
rect 928 155 930 196
rect 976 155 978 196
rect 1024 155 1026 196
rect 1240 155 1242 219
rect 1278 216 1284 217
rect 1278 212 1279 216
rect 1283 212 1284 216
rect 1278 211 1284 212
rect 2406 216 2412 217
rect 2406 212 2407 216
rect 2411 212 2412 216
rect 2406 211 2412 212
rect 1280 171 1282 211
rect 1366 193 1372 194
rect 1366 189 1367 193
rect 1371 189 1372 193
rect 1366 188 1372 189
rect 1406 193 1412 194
rect 1406 189 1407 193
rect 1411 189 1412 193
rect 1406 188 1412 189
rect 1454 193 1460 194
rect 1454 189 1455 193
rect 1459 189 1460 193
rect 1454 188 1460 189
rect 1510 193 1516 194
rect 1510 189 1511 193
rect 1515 189 1516 193
rect 1510 188 1516 189
rect 1566 193 1572 194
rect 1566 189 1567 193
rect 1571 189 1572 193
rect 1566 188 1572 189
rect 1630 193 1636 194
rect 1630 189 1631 193
rect 1635 189 1636 193
rect 1630 188 1636 189
rect 1702 193 1708 194
rect 1702 189 1703 193
rect 1707 189 1708 193
rect 1702 188 1708 189
rect 1774 193 1780 194
rect 1774 189 1775 193
rect 1779 189 1780 193
rect 1774 188 1780 189
rect 1854 193 1860 194
rect 1854 189 1855 193
rect 1859 189 1860 193
rect 1854 188 1860 189
rect 1942 193 1948 194
rect 1942 189 1943 193
rect 1947 189 1948 193
rect 1942 188 1948 189
rect 2030 193 2036 194
rect 2030 189 2031 193
rect 2035 189 2036 193
rect 2030 188 2036 189
rect 2118 193 2124 194
rect 2118 189 2119 193
rect 2123 189 2124 193
rect 2118 188 2124 189
rect 2206 193 2212 194
rect 2206 189 2207 193
rect 2211 189 2212 193
rect 2206 188 2212 189
rect 2294 193 2300 194
rect 2294 189 2295 193
rect 2299 189 2300 193
rect 2294 188 2300 189
rect 2358 193 2364 194
rect 2358 189 2359 193
rect 2363 189 2364 193
rect 2358 188 2364 189
rect 1368 171 1370 188
rect 1408 171 1410 188
rect 1456 171 1458 188
rect 1512 171 1514 188
rect 1568 171 1570 188
rect 1632 171 1634 188
rect 1704 171 1706 188
rect 1776 171 1778 188
rect 1856 171 1858 188
rect 1944 171 1946 188
rect 2032 171 2034 188
rect 2120 171 2122 188
rect 2208 171 2210 188
rect 2296 171 2298 188
rect 2360 171 2362 188
rect 2408 171 2410 211
rect 1279 170 1283 171
rect 1279 165 1283 166
rect 1303 170 1307 171
rect 1303 165 1307 166
rect 1343 170 1347 171
rect 1343 165 1347 166
rect 1367 170 1371 171
rect 1367 165 1371 166
rect 1383 170 1387 171
rect 1383 165 1387 166
rect 1407 170 1411 171
rect 1407 165 1411 166
rect 1423 170 1427 171
rect 1423 165 1427 166
rect 1455 170 1459 171
rect 1455 165 1459 166
rect 1463 170 1467 171
rect 1463 165 1467 166
rect 1511 170 1515 171
rect 1511 165 1515 166
rect 1519 170 1523 171
rect 1519 165 1523 166
rect 1567 170 1571 171
rect 1567 165 1571 166
rect 1583 170 1587 171
rect 1583 165 1587 166
rect 1631 170 1635 171
rect 1631 165 1635 166
rect 1647 170 1651 171
rect 1647 165 1651 166
rect 1703 170 1707 171
rect 1703 165 1707 166
rect 1711 170 1715 171
rect 1711 165 1715 166
rect 1775 170 1779 171
rect 1775 165 1779 166
rect 1831 170 1835 171
rect 1831 165 1835 166
rect 1855 170 1859 171
rect 1855 165 1859 166
rect 1887 170 1891 171
rect 1887 165 1891 166
rect 1935 170 1939 171
rect 1935 165 1939 166
rect 1943 170 1947 171
rect 1943 165 1947 166
rect 1975 170 1979 171
rect 1975 165 1979 166
rect 2015 170 2019 171
rect 2015 165 2019 166
rect 2031 170 2035 171
rect 2031 165 2035 166
rect 2055 170 2059 171
rect 2055 165 2059 166
rect 2095 170 2099 171
rect 2095 165 2099 166
rect 2119 170 2123 171
rect 2119 165 2123 166
rect 2143 170 2147 171
rect 2143 165 2147 166
rect 2191 170 2195 171
rect 2191 165 2195 166
rect 2207 170 2211 171
rect 2207 165 2211 166
rect 2239 170 2243 171
rect 2239 165 2243 166
rect 2279 170 2283 171
rect 2279 165 2283 166
rect 2295 170 2299 171
rect 2295 165 2299 166
rect 2319 170 2323 171
rect 2319 165 2323 166
rect 2359 170 2363 171
rect 2359 165 2363 166
rect 2407 170 2411 171
rect 2407 165 2411 166
rect 111 154 115 155
rect 111 149 115 150
rect 135 154 139 155
rect 135 149 139 150
rect 151 154 155 155
rect 151 149 155 150
rect 191 154 195 155
rect 191 149 195 150
rect 223 154 227 155
rect 223 149 227 150
rect 231 154 235 155
rect 231 149 235 150
rect 271 154 275 155
rect 271 149 275 150
rect 311 154 315 155
rect 311 149 315 150
rect 351 154 355 155
rect 351 149 355 150
rect 391 154 395 155
rect 391 149 395 150
rect 431 154 435 155
rect 431 149 435 150
rect 463 154 467 155
rect 463 149 467 150
rect 471 154 475 155
rect 471 149 475 150
rect 511 154 515 155
rect 511 149 515 150
rect 527 154 531 155
rect 527 149 531 150
rect 551 154 555 155
rect 551 149 555 150
rect 591 154 595 155
rect 591 149 595 150
rect 631 154 635 155
rect 631 149 635 150
rect 647 154 651 155
rect 647 149 651 150
rect 671 154 675 155
rect 671 149 675 150
rect 695 154 699 155
rect 695 149 699 150
rect 711 154 715 155
rect 711 149 715 150
rect 735 154 739 155
rect 735 149 739 150
rect 751 154 755 155
rect 751 149 755 150
rect 783 154 787 155
rect 783 149 787 150
rect 791 154 795 155
rect 791 149 795 150
rect 831 154 835 155
rect 831 149 835 150
rect 871 154 875 155
rect 871 149 875 150
rect 879 154 883 155
rect 879 149 883 150
rect 911 154 915 155
rect 911 149 915 150
rect 927 154 931 155
rect 927 149 931 150
rect 951 154 955 155
rect 951 149 955 150
rect 975 154 979 155
rect 975 149 979 150
rect 991 154 995 155
rect 991 149 995 150
rect 1023 154 1027 155
rect 1023 149 1027 150
rect 1031 154 1035 155
rect 1031 149 1035 150
rect 1071 154 1075 155
rect 1071 149 1075 150
rect 1111 154 1115 155
rect 1111 149 1115 150
rect 1151 154 1155 155
rect 1151 149 1155 150
rect 1191 154 1195 155
rect 1191 149 1195 150
rect 1239 154 1243 155
rect 1239 149 1243 150
rect 112 117 114 149
rect 152 140 154 149
rect 192 140 194 149
rect 232 140 234 149
rect 272 140 274 149
rect 312 140 314 149
rect 352 140 354 149
rect 392 140 394 149
rect 432 140 434 149
rect 472 140 474 149
rect 512 140 514 149
rect 552 140 554 149
rect 592 140 594 149
rect 632 140 634 149
rect 672 140 674 149
rect 712 140 714 149
rect 752 140 754 149
rect 792 140 794 149
rect 832 140 834 149
rect 872 140 874 149
rect 912 140 914 149
rect 952 140 954 149
rect 992 140 994 149
rect 1032 140 1034 149
rect 1072 140 1074 149
rect 1112 140 1114 149
rect 1152 140 1154 149
rect 1192 140 1194 149
rect 150 139 156 140
rect 150 135 151 139
rect 155 135 156 139
rect 150 134 156 135
rect 190 139 196 140
rect 190 135 191 139
rect 195 135 196 139
rect 190 134 196 135
rect 230 139 236 140
rect 230 135 231 139
rect 235 135 236 139
rect 230 134 236 135
rect 270 139 276 140
rect 270 135 271 139
rect 275 135 276 139
rect 270 134 276 135
rect 310 139 316 140
rect 310 135 311 139
rect 315 135 316 139
rect 310 134 316 135
rect 350 139 356 140
rect 350 135 351 139
rect 355 135 356 139
rect 350 134 356 135
rect 390 139 396 140
rect 390 135 391 139
rect 395 135 396 139
rect 390 134 396 135
rect 430 139 436 140
rect 430 135 431 139
rect 435 135 436 139
rect 430 134 436 135
rect 470 139 476 140
rect 470 135 471 139
rect 475 135 476 139
rect 470 134 476 135
rect 510 139 516 140
rect 510 135 511 139
rect 515 135 516 139
rect 510 134 516 135
rect 550 139 556 140
rect 550 135 551 139
rect 555 135 556 139
rect 550 134 556 135
rect 590 139 596 140
rect 590 135 591 139
rect 595 135 596 139
rect 590 134 596 135
rect 630 139 636 140
rect 630 135 631 139
rect 635 135 636 139
rect 630 134 636 135
rect 670 139 676 140
rect 670 135 671 139
rect 675 135 676 139
rect 670 134 676 135
rect 710 139 716 140
rect 710 135 711 139
rect 715 135 716 139
rect 710 134 716 135
rect 750 139 756 140
rect 750 135 751 139
rect 755 135 756 139
rect 750 134 756 135
rect 790 139 796 140
rect 790 135 791 139
rect 795 135 796 139
rect 790 134 796 135
rect 830 139 836 140
rect 830 135 831 139
rect 835 135 836 139
rect 830 134 836 135
rect 870 139 876 140
rect 870 135 871 139
rect 875 135 876 139
rect 870 134 876 135
rect 910 139 916 140
rect 910 135 911 139
rect 915 135 916 139
rect 910 134 916 135
rect 950 139 956 140
rect 950 135 951 139
rect 955 135 956 139
rect 950 134 956 135
rect 990 139 996 140
rect 990 135 991 139
rect 995 135 996 139
rect 990 134 996 135
rect 1030 139 1036 140
rect 1030 135 1031 139
rect 1035 135 1036 139
rect 1030 134 1036 135
rect 1070 139 1076 140
rect 1070 135 1071 139
rect 1075 135 1076 139
rect 1070 134 1076 135
rect 1110 139 1116 140
rect 1110 135 1111 139
rect 1115 135 1116 139
rect 1110 134 1116 135
rect 1150 139 1156 140
rect 1150 135 1151 139
rect 1155 135 1156 139
rect 1150 134 1156 135
rect 1190 139 1196 140
rect 1190 135 1191 139
rect 1195 135 1196 139
rect 1190 134 1196 135
rect 1240 117 1242 149
rect 1280 133 1282 165
rect 1304 156 1306 165
rect 1344 156 1346 165
rect 1384 156 1386 165
rect 1424 156 1426 165
rect 1464 156 1466 165
rect 1520 156 1522 165
rect 1584 156 1586 165
rect 1648 156 1650 165
rect 1712 156 1714 165
rect 1776 156 1778 165
rect 1832 156 1834 165
rect 1888 156 1890 165
rect 1936 156 1938 165
rect 1976 156 1978 165
rect 2016 156 2018 165
rect 2056 156 2058 165
rect 2096 156 2098 165
rect 2144 156 2146 165
rect 2192 156 2194 165
rect 2240 156 2242 165
rect 2280 156 2282 165
rect 2320 156 2322 165
rect 2360 156 2362 165
rect 1302 155 1308 156
rect 1302 151 1303 155
rect 1307 151 1308 155
rect 1302 150 1308 151
rect 1342 155 1348 156
rect 1342 151 1343 155
rect 1347 151 1348 155
rect 1342 150 1348 151
rect 1382 155 1388 156
rect 1382 151 1383 155
rect 1387 151 1388 155
rect 1382 150 1388 151
rect 1422 155 1428 156
rect 1422 151 1423 155
rect 1427 151 1428 155
rect 1422 150 1428 151
rect 1462 155 1468 156
rect 1462 151 1463 155
rect 1467 151 1468 155
rect 1462 150 1468 151
rect 1518 155 1524 156
rect 1518 151 1519 155
rect 1523 151 1524 155
rect 1518 150 1524 151
rect 1582 155 1588 156
rect 1582 151 1583 155
rect 1587 151 1588 155
rect 1582 150 1588 151
rect 1646 155 1652 156
rect 1646 151 1647 155
rect 1651 151 1652 155
rect 1646 150 1652 151
rect 1710 155 1716 156
rect 1710 151 1711 155
rect 1715 151 1716 155
rect 1710 150 1716 151
rect 1774 155 1780 156
rect 1774 151 1775 155
rect 1779 151 1780 155
rect 1774 150 1780 151
rect 1830 155 1836 156
rect 1830 151 1831 155
rect 1835 151 1836 155
rect 1830 150 1836 151
rect 1886 155 1892 156
rect 1886 151 1887 155
rect 1891 151 1892 155
rect 1886 150 1892 151
rect 1934 155 1940 156
rect 1934 151 1935 155
rect 1939 151 1940 155
rect 1934 150 1940 151
rect 1974 155 1980 156
rect 1974 151 1975 155
rect 1979 151 1980 155
rect 1974 150 1980 151
rect 2014 155 2020 156
rect 2014 151 2015 155
rect 2019 151 2020 155
rect 2014 150 2020 151
rect 2054 155 2060 156
rect 2054 151 2055 155
rect 2059 151 2060 155
rect 2054 150 2060 151
rect 2094 155 2100 156
rect 2094 151 2095 155
rect 2099 151 2100 155
rect 2094 150 2100 151
rect 2142 155 2148 156
rect 2142 151 2143 155
rect 2147 151 2148 155
rect 2142 150 2148 151
rect 2190 155 2196 156
rect 2190 151 2191 155
rect 2195 151 2196 155
rect 2190 150 2196 151
rect 2238 155 2244 156
rect 2238 151 2239 155
rect 2243 151 2244 155
rect 2238 150 2244 151
rect 2278 155 2284 156
rect 2278 151 2279 155
rect 2283 151 2284 155
rect 2278 150 2284 151
rect 2318 155 2324 156
rect 2318 151 2319 155
rect 2323 151 2324 155
rect 2318 150 2324 151
rect 2358 155 2364 156
rect 2358 151 2359 155
rect 2363 151 2364 155
rect 2358 150 2364 151
rect 2408 133 2410 165
rect 1278 132 1284 133
rect 1278 128 1279 132
rect 1283 128 1284 132
rect 1278 127 1284 128
rect 2406 132 2412 133
rect 2406 128 2407 132
rect 2411 128 2412 132
rect 2406 127 2412 128
rect 110 116 116 117
rect 110 112 111 116
rect 115 112 116 116
rect 110 111 116 112
rect 1238 116 1244 117
rect 1238 112 1239 116
rect 1243 112 1244 116
rect 1238 111 1244 112
rect 1278 115 1284 116
rect 1278 111 1279 115
rect 1283 111 1284 115
rect 1278 110 1284 111
rect 2406 115 2412 116
rect 2406 111 2407 115
rect 2411 111 2412 115
rect 2406 110 2412 111
rect 1280 103 1282 110
rect 1302 108 1308 109
rect 1302 104 1303 108
rect 1307 104 1308 108
rect 1302 103 1308 104
rect 1342 108 1348 109
rect 1342 104 1343 108
rect 1347 104 1348 108
rect 1342 103 1348 104
rect 1382 108 1388 109
rect 1382 104 1383 108
rect 1387 104 1388 108
rect 1382 103 1388 104
rect 1422 108 1428 109
rect 1422 104 1423 108
rect 1427 104 1428 108
rect 1422 103 1428 104
rect 1462 108 1468 109
rect 1462 104 1463 108
rect 1467 104 1468 108
rect 1462 103 1468 104
rect 1518 108 1524 109
rect 1518 104 1519 108
rect 1523 104 1524 108
rect 1518 103 1524 104
rect 1582 108 1588 109
rect 1582 104 1583 108
rect 1587 104 1588 108
rect 1582 103 1588 104
rect 1646 108 1652 109
rect 1646 104 1647 108
rect 1651 104 1652 108
rect 1646 103 1652 104
rect 1710 108 1716 109
rect 1710 104 1711 108
rect 1715 104 1716 108
rect 1710 103 1716 104
rect 1774 108 1780 109
rect 1774 104 1775 108
rect 1779 104 1780 108
rect 1774 103 1780 104
rect 1830 108 1836 109
rect 1830 104 1831 108
rect 1835 104 1836 108
rect 1830 103 1836 104
rect 1886 108 1892 109
rect 1886 104 1887 108
rect 1891 104 1892 108
rect 1886 103 1892 104
rect 1934 108 1940 109
rect 1934 104 1935 108
rect 1939 104 1940 108
rect 1934 103 1940 104
rect 1974 108 1980 109
rect 1974 104 1975 108
rect 1979 104 1980 108
rect 1974 103 1980 104
rect 2014 108 2020 109
rect 2014 104 2015 108
rect 2019 104 2020 108
rect 2014 103 2020 104
rect 2054 108 2060 109
rect 2054 104 2055 108
rect 2059 104 2060 108
rect 2054 103 2060 104
rect 2094 108 2100 109
rect 2094 104 2095 108
rect 2099 104 2100 108
rect 2094 103 2100 104
rect 2142 108 2148 109
rect 2142 104 2143 108
rect 2147 104 2148 108
rect 2142 103 2148 104
rect 2190 108 2196 109
rect 2190 104 2191 108
rect 2195 104 2196 108
rect 2190 103 2196 104
rect 2238 108 2244 109
rect 2238 104 2239 108
rect 2243 104 2244 108
rect 2238 103 2244 104
rect 2278 108 2284 109
rect 2278 104 2279 108
rect 2283 104 2284 108
rect 2278 103 2284 104
rect 2318 108 2324 109
rect 2318 104 2319 108
rect 2323 104 2324 108
rect 2318 103 2324 104
rect 2358 108 2364 109
rect 2358 104 2359 108
rect 2363 104 2364 108
rect 2358 103 2364 104
rect 2408 103 2410 110
rect 1279 102 1283 103
rect 110 99 116 100
rect 110 95 111 99
rect 115 95 116 99
rect 110 94 116 95
rect 1238 99 1244 100
rect 1238 95 1239 99
rect 1243 95 1244 99
rect 1279 97 1283 98
rect 1303 102 1307 103
rect 1303 97 1307 98
rect 1343 102 1347 103
rect 1343 97 1347 98
rect 1383 102 1387 103
rect 1383 97 1387 98
rect 1423 102 1427 103
rect 1423 97 1427 98
rect 1463 102 1467 103
rect 1463 97 1467 98
rect 1519 102 1523 103
rect 1519 97 1523 98
rect 1583 102 1587 103
rect 1583 97 1587 98
rect 1647 102 1651 103
rect 1647 97 1651 98
rect 1711 102 1715 103
rect 1711 97 1715 98
rect 1775 102 1779 103
rect 1775 97 1779 98
rect 1831 102 1835 103
rect 1831 97 1835 98
rect 1887 102 1891 103
rect 1887 97 1891 98
rect 1935 102 1939 103
rect 1935 97 1939 98
rect 1975 102 1979 103
rect 1975 97 1979 98
rect 2015 102 2019 103
rect 2015 97 2019 98
rect 2055 102 2059 103
rect 2055 97 2059 98
rect 2095 102 2099 103
rect 2095 97 2099 98
rect 2143 102 2147 103
rect 2143 97 2147 98
rect 2191 102 2195 103
rect 2191 97 2195 98
rect 2239 102 2243 103
rect 2239 97 2243 98
rect 2279 102 2283 103
rect 2279 97 2283 98
rect 2319 102 2323 103
rect 2319 97 2323 98
rect 2359 102 2363 103
rect 2359 97 2363 98
rect 2407 102 2411 103
rect 2407 97 2411 98
rect 1238 94 1244 95
rect 112 87 114 94
rect 150 92 156 93
rect 150 88 151 92
rect 155 88 156 92
rect 150 87 156 88
rect 190 92 196 93
rect 190 88 191 92
rect 195 88 196 92
rect 190 87 196 88
rect 230 92 236 93
rect 230 88 231 92
rect 235 88 236 92
rect 230 87 236 88
rect 270 92 276 93
rect 270 88 271 92
rect 275 88 276 92
rect 270 87 276 88
rect 310 92 316 93
rect 310 88 311 92
rect 315 88 316 92
rect 310 87 316 88
rect 350 92 356 93
rect 350 88 351 92
rect 355 88 356 92
rect 350 87 356 88
rect 390 92 396 93
rect 390 88 391 92
rect 395 88 396 92
rect 390 87 396 88
rect 430 92 436 93
rect 430 88 431 92
rect 435 88 436 92
rect 430 87 436 88
rect 470 92 476 93
rect 470 88 471 92
rect 475 88 476 92
rect 470 87 476 88
rect 510 92 516 93
rect 510 88 511 92
rect 515 88 516 92
rect 510 87 516 88
rect 550 92 556 93
rect 550 88 551 92
rect 555 88 556 92
rect 550 87 556 88
rect 590 92 596 93
rect 590 88 591 92
rect 595 88 596 92
rect 590 87 596 88
rect 630 92 636 93
rect 630 88 631 92
rect 635 88 636 92
rect 630 87 636 88
rect 670 92 676 93
rect 670 88 671 92
rect 675 88 676 92
rect 670 87 676 88
rect 710 92 716 93
rect 710 88 711 92
rect 715 88 716 92
rect 710 87 716 88
rect 750 92 756 93
rect 750 88 751 92
rect 755 88 756 92
rect 750 87 756 88
rect 790 92 796 93
rect 790 88 791 92
rect 795 88 796 92
rect 790 87 796 88
rect 830 92 836 93
rect 830 88 831 92
rect 835 88 836 92
rect 830 87 836 88
rect 870 92 876 93
rect 870 88 871 92
rect 875 88 876 92
rect 870 87 876 88
rect 910 92 916 93
rect 910 88 911 92
rect 915 88 916 92
rect 910 87 916 88
rect 950 92 956 93
rect 950 88 951 92
rect 955 88 956 92
rect 950 87 956 88
rect 990 92 996 93
rect 990 88 991 92
rect 995 88 996 92
rect 990 87 996 88
rect 1030 92 1036 93
rect 1030 88 1031 92
rect 1035 88 1036 92
rect 1030 87 1036 88
rect 1070 92 1076 93
rect 1070 88 1071 92
rect 1075 88 1076 92
rect 1070 87 1076 88
rect 1110 92 1116 93
rect 1110 88 1111 92
rect 1115 88 1116 92
rect 1110 87 1116 88
rect 1150 92 1156 93
rect 1150 88 1151 92
rect 1155 88 1156 92
rect 1150 87 1156 88
rect 1190 92 1196 93
rect 1190 88 1191 92
rect 1195 88 1196 92
rect 1190 87 1196 88
rect 1240 87 1242 94
rect 111 86 115 87
rect 111 81 115 82
rect 151 86 155 87
rect 151 81 155 82
rect 191 86 195 87
rect 191 81 195 82
rect 231 86 235 87
rect 231 81 235 82
rect 271 86 275 87
rect 271 81 275 82
rect 311 86 315 87
rect 311 81 315 82
rect 351 86 355 87
rect 351 81 355 82
rect 391 86 395 87
rect 391 81 395 82
rect 431 86 435 87
rect 431 81 435 82
rect 471 86 475 87
rect 471 81 475 82
rect 511 86 515 87
rect 511 81 515 82
rect 551 86 555 87
rect 551 81 555 82
rect 591 86 595 87
rect 591 81 595 82
rect 631 86 635 87
rect 631 81 635 82
rect 671 86 675 87
rect 671 81 675 82
rect 711 86 715 87
rect 711 81 715 82
rect 751 86 755 87
rect 751 81 755 82
rect 791 86 795 87
rect 791 81 795 82
rect 831 86 835 87
rect 831 81 835 82
rect 871 86 875 87
rect 871 81 875 82
rect 911 86 915 87
rect 911 81 915 82
rect 951 86 955 87
rect 951 81 955 82
rect 991 86 995 87
rect 991 81 995 82
rect 1031 86 1035 87
rect 1031 81 1035 82
rect 1071 86 1075 87
rect 1071 81 1075 82
rect 1111 86 1115 87
rect 1111 81 1115 82
rect 1151 86 1155 87
rect 1151 81 1155 82
rect 1191 86 1195 87
rect 1191 81 1195 82
rect 1239 86 1243 87
rect 1239 81 1243 82
<< m4c >>
rect 111 2490 115 2494
rect 231 2490 235 2494
rect 271 2490 275 2494
rect 311 2490 315 2494
rect 351 2490 355 2494
rect 399 2490 403 2494
rect 455 2490 459 2494
rect 511 2490 515 2494
rect 575 2490 579 2494
rect 639 2490 643 2494
rect 703 2490 707 2494
rect 767 2490 771 2494
rect 823 2490 827 2494
rect 879 2490 883 2494
rect 927 2490 931 2494
rect 975 2490 979 2494
rect 1023 2490 1027 2494
rect 1071 2490 1075 2494
rect 1111 2490 1115 2494
rect 1151 2490 1155 2494
rect 1191 2490 1195 2494
rect 1239 2490 1243 2494
rect 1279 2486 1283 2490
rect 1303 2486 1307 2490
rect 1343 2486 1347 2490
rect 1383 2486 1387 2490
rect 1439 2486 1443 2490
rect 1511 2486 1515 2490
rect 1583 2486 1587 2490
rect 1663 2486 1667 2490
rect 1735 2486 1739 2490
rect 1807 2486 1811 2490
rect 1887 2486 1891 2490
rect 1967 2486 1971 2490
rect 2063 2486 2067 2490
rect 2167 2486 2171 2490
rect 2271 2486 2275 2490
rect 2359 2486 2363 2490
rect 2407 2486 2411 2490
rect 111 2414 115 2418
rect 199 2414 203 2418
rect 231 2414 235 2418
rect 263 2414 267 2418
rect 271 2414 275 2418
rect 311 2414 315 2418
rect 327 2414 331 2418
rect 351 2414 355 2418
rect 399 2414 403 2418
rect 455 2414 459 2418
rect 471 2414 475 2418
rect 511 2414 515 2418
rect 543 2414 547 2418
rect 575 2414 579 2418
rect 615 2414 619 2418
rect 639 2414 643 2418
rect 687 2414 691 2418
rect 703 2414 707 2418
rect 751 2414 755 2418
rect 767 2414 771 2418
rect 823 2414 827 2418
rect 879 2414 883 2418
rect 895 2414 899 2418
rect 927 2414 931 2418
rect 967 2414 971 2418
rect 975 2414 979 2418
rect 1023 2414 1027 2418
rect 1071 2414 1075 2418
rect 1111 2414 1115 2418
rect 1151 2414 1155 2418
rect 1191 2414 1195 2418
rect 1239 2414 1243 2418
rect 1279 2418 1283 2422
rect 1303 2418 1307 2422
rect 1343 2418 1347 2422
rect 1375 2418 1379 2422
rect 1383 2418 1387 2422
rect 1415 2418 1419 2422
rect 1439 2418 1443 2422
rect 1455 2418 1459 2422
rect 1503 2418 1507 2422
rect 1511 2418 1515 2422
rect 1559 2418 1563 2422
rect 1583 2418 1587 2422
rect 1615 2418 1619 2422
rect 1663 2418 1667 2422
rect 1679 2418 1683 2422
rect 1735 2418 1739 2422
rect 1799 2418 1803 2422
rect 1807 2418 1811 2422
rect 1871 2418 1875 2422
rect 1887 2418 1891 2422
rect 1951 2418 1955 2422
rect 1967 2418 1971 2422
rect 2047 2418 2051 2422
rect 2063 2418 2067 2422
rect 2151 2418 2155 2422
rect 2167 2418 2171 2422
rect 2263 2418 2267 2422
rect 2271 2418 2275 2422
rect 2359 2418 2363 2422
rect 2407 2418 2411 2422
rect 111 2342 115 2346
rect 199 2342 203 2346
rect 263 2342 267 2346
rect 271 2342 275 2346
rect 327 2342 331 2346
rect 399 2342 403 2346
rect 471 2342 475 2346
rect 543 2342 547 2346
rect 551 2342 555 2346
rect 615 2342 619 2346
rect 631 2342 635 2346
rect 687 2342 691 2346
rect 711 2342 715 2346
rect 751 2342 755 2346
rect 783 2342 787 2346
rect 823 2342 827 2346
rect 855 2342 859 2346
rect 895 2342 899 2346
rect 919 2342 923 2346
rect 967 2342 971 2346
rect 991 2342 995 2346
rect 1063 2342 1067 2346
rect 1239 2342 1243 2346
rect 1279 2346 1283 2350
rect 1327 2346 1331 2350
rect 1375 2346 1379 2350
rect 1383 2346 1387 2350
rect 1415 2346 1419 2350
rect 1439 2346 1443 2350
rect 1455 2346 1459 2350
rect 1503 2346 1507 2350
rect 1559 2346 1563 2350
rect 1575 2346 1579 2350
rect 1615 2346 1619 2350
rect 1647 2346 1651 2350
rect 1679 2346 1683 2350
rect 1719 2346 1723 2350
rect 1735 2346 1739 2350
rect 1799 2346 1803 2350
rect 1871 2346 1875 2350
rect 1879 2346 1883 2350
rect 1951 2346 1955 2350
rect 1967 2346 1971 2350
rect 2047 2346 2051 2350
rect 2063 2346 2067 2350
rect 2151 2346 2155 2350
rect 2167 2346 2171 2350
rect 2263 2346 2267 2350
rect 2271 2346 2275 2350
rect 2359 2346 2363 2350
rect 2407 2346 2411 2350
rect 1279 2278 1283 2282
rect 1327 2278 1331 2282
rect 1335 2278 1339 2282
rect 1383 2278 1387 2282
rect 1407 2278 1411 2282
rect 1439 2278 1443 2282
rect 1487 2278 1491 2282
rect 1503 2278 1507 2282
rect 1559 2278 1563 2282
rect 1575 2278 1579 2282
rect 1631 2278 1635 2282
rect 1647 2278 1651 2282
rect 1703 2278 1707 2282
rect 1719 2278 1723 2282
rect 1775 2278 1779 2282
rect 1799 2278 1803 2282
rect 1839 2278 1843 2282
rect 1879 2278 1883 2282
rect 1911 2278 1915 2282
rect 1967 2278 1971 2282
rect 1991 2278 1995 2282
rect 2063 2278 2067 2282
rect 2079 2278 2083 2282
rect 2167 2278 2171 2282
rect 2175 2278 2179 2282
rect 2271 2278 2275 2282
rect 2279 2278 2283 2282
rect 2359 2278 2363 2282
rect 2407 2278 2411 2282
rect 111 2266 115 2270
rect 143 2266 147 2270
rect 183 2266 187 2270
rect 223 2266 227 2270
rect 271 2266 275 2270
rect 279 2266 283 2270
rect 327 2266 331 2270
rect 335 2266 339 2270
rect 399 2266 403 2270
rect 407 2266 411 2270
rect 471 2266 475 2270
rect 479 2266 483 2270
rect 551 2266 555 2270
rect 559 2266 563 2270
rect 631 2266 635 2270
rect 647 2266 651 2270
rect 711 2266 715 2270
rect 727 2266 731 2270
rect 783 2266 787 2270
rect 807 2266 811 2270
rect 855 2266 859 2270
rect 887 2266 891 2270
rect 919 2266 923 2270
rect 967 2266 971 2270
rect 991 2266 995 2270
rect 1047 2266 1051 2270
rect 1063 2266 1067 2270
rect 1127 2266 1131 2270
rect 1239 2266 1243 2270
rect 111 2198 115 2202
rect 135 2198 139 2202
rect 143 2198 147 2202
rect 183 2198 187 2202
rect 207 2198 211 2202
rect 223 2198 227 2202
rect 279 2198 283 2202
rect 335 2198 339 2202
rect 359 2198 363 2202
rect 407 2198 411 2202
rect 439 2198 443 2202
rect 479 2198 483 2202
rect 519 2198 523 2202
rect 559 2198 563 2202
rect 599 2198 603 2202
rect 647 2198 651 2202
rect 679 2198 683 2202
rect 727 2198 731 2202
rect 759 2198 763 2202
rect 807 2198 811 2202
rect 831 2198 835 2202
rect 887 2198 891 2202
rect 903 2198 907 2202
rect 967 2198 971 2202
rect 975 2198 979 2202
rect 1047 2198 1051 2202
rect 1119 2198 1123 2202
rect 1127 2198 1131 2202
rect 1239 2198 1243 2202
rect 1279 2202 1283 2206
rect 1335 2202 1339 2206
rect 1375 2202 1379 2206
rect 1407 2202 1411 2206
rect 1439 2202 1443 2206
rect 1487 2202 1491 2206
rect 1511 2202 1515 2206
rect 1559 2202 1563 2206
rect 1591 2202 1595 2206
rect 1631 2202 1635 2206
rect 1671 2202 1675 2206
rect 1703 2202 1707 2206
rect 1751 2202 1755 2206
rect 1775 2202 1779 2206
rect 1831 2202 1835 2206
rect 1839 2202 1843 2206
rect 1903 2202 1907 2206
rect 1911 2202 1915 2206
rect 1967 2202 1971 2206
rect 1991 2202 1995 2206
rect 2031 2202 2035 2206
rect 2079 2202 2083 2206
rect 2095 2202 2099 2206
rect 2167 2202 2171 2206
rect 2175 2202 2179 2206
rect 2239 2202 2243 2206
rect 2279 2202 2283 2206
rect 2311 2202 2315 2206
rect 2359 2202 2363 2206
rect 2407 2202 2411 2206
rect 1279 2134 1283 2138
rect 1375 2134 1379 2138
rect 1399 2134 1403 2138
rect 1439 2134 1443 2138
rect 1495 2134 1499 2138
rect 1511 2134 1515 2138
rect 1567 2134 1571 2138
rect 1591 2134 1595 2138
rect 1647 2134 1651 2138
rect 1671 2134 1675 2138
rect 1735 2134 1739 2138
rect 1751 2134 1755 2138
rect 1823 2134 1827 2138
rect 1831 2134 1835 2138
rect 1903 2134 1907 2138
rect 1911 2134 1915 2138
rect 1967 2134 1971 2138
rect 1999 2134 2003 2138
rect 2031 2134 2035 2138
rect 2087 2134 2091 2138
rect 2095 2134 2099 2138
rect 2167 2134 2171 2138
rect 2175 2134 2179 2138
rect 2239 2134 2243 2138
rect 2271 2134 2275 2138
rect 2311 2134 2315 2138
rect 2359 2134 2363 2138
rect 2407 2134 2411 2138
rect 111 2122 115 2126
rect 135 2122 139 2126
rect 191 2122 195 2126
rect 207 2122 211 2126
rect 271 2122 275 2126
rect 279 2122 283 2126
rect 343 2122 347 2126
rect 359 2122 363 2126
rect 415 2122 419 2126
rect 439 2122 443 2126
rect 479 2122 483 2126
rect 519 2122 523 2126
rect 543 2122 547 2126
rect 599 2122 603 2126
rect 607 2122 611 2126
rect 671 2122 675 2126
rect 679 2122 683 2126
rect 735 2122 739 2126
rect 759 2122 763 2126
rect 791 2122 795 2126
rect 831 2122 835 2126
rect 839 2122 843 2126
rect 887 2122 891 2126
rect 903 2122 907 2126
rect 935 2122 939 2126
rect 975 2122 979 2126
rect 991 2122 995 2126
rect 1047 2122 1051 2126
rect 1119 2122 1123 2126
rect 1239 2122 1243 2126
rect 1279 2066 1283 2070
rect 1399 2066 1403 2070
rect 1439 2066 1443 2070
rect 1495 2066 1499 2070
rect 1567 2066 1571 2070
rect 1647 2066 1651 2070
rect 1735 2066 1739 2070
rect 1823 2066 1827 2070
rect 1911 2066 1915 2070
rect 1999 2066 2003 2070
rect 2039 2066 2043 2070
rect 2079 2066 2083 2070
rect 2087 2066 2091 2070
rect 2119 2066 2123 2070
rect 2159 2066 2163 2070
rect 2175 2066 2179 2070
rect 2199 2066 2203 2070
rect 2239 2066 2243 2070
rect 2271 2066 2275 2070
rect 2279 2066 2283 2070
rect 2319 2066 2323 2070
rect 2359 2066 2363 2070
rect 2407 2066 2411 2070
rect 111 2050 115 2054
rect 135 2050 139 2054
rect 175 2050 179 2054
rect 191 2050 195 2054
rect 215 2050 219 2054
rect 271 2050 275 2054
rect 279 2050 283 2054
rect 343 2050 347 2054
rect 351 2050 355 2054
rect 415 2050 419 2054
rect 423 2050 427 2054
rect 479 2050 483 2054
rect 487 2050 491 2054
rect 543 2050 547 2054
rect 551 2050 555 2054
rect 607 2050 611 2054
rect 615 2050 619 2054
rect 671 2050 675 2054
rect 679 2050 683 2054
rect 735 2050 739 2054
rect 743 2050 747 2054
rect 791 2050 795 2054
rect 815 2050 819 2054
rect 839 2050 843 2054
rect 887 2050 891 2054
rect 935 2050 939 2054
rect 991 2050 995 2054
rect 1047 2050 1051 2054
rect 1239 2050 1243 2054
rect 1279 1998 1283 2002
rect 1399 1998 1403 2002
rect 1439 1998 1443 2002
rect 1479 1998 1483 2002
rect 1519 1998 1523 2002
rect 1559 1998 1563 2002
rect 1599 1998 1603 2002
rect 1639 1998 1643 2002
rect 1679 1998 1683 2002
rect 1719 1998 1723 2002
rect 1767 1998 1771 2002
rect 1823 1998 1827 2002
rect 1871 1998 1875 2002
rect 1919 1998 1923 2002
rect 1967 1998 1971 2002
rect 2015 1998 2019 2002
rect 2039 1998 2043 2002
rect 2055 1998 2059 2002
rect 2079 1998 2083 2002
rect 2095 1998 2099 2002
rect 2119 1998 2123 2002
rect 2143 1998 2147 2002
rect 2159 1998 2163 2002
rect 2191 1998 2195 2002
rect 2199 1998 2203 2002
rect 2239 1998 2243 2002
rect 2279 1998 2283 2002
rect 2319 1998 2323 2002
rect 2359 1998 2363 2002
rect 2407 1998 2411 2002
rect 111 1982 115 1986
rect 135 1982 139 1986
rect 175 1982 179 1986
rect 215 1982 219 1986
rect 271 1982 275 1986
rect 279 1982 283 1986
rect 343 1982 347 1986
rect 351 1982 355 1986
rect 415 1982 419 1986
rect 423 1982 427 1986
rect 487 1982 491 1986
rect 495 1982 499 1986
rect 551 1982 555 1986
rect 575 1982 579 1986
rect 615 1982 619 1986
rect 647 1982 651 1986
rect 679 1982 683 1986
rect 719 1982 723 1986
rect 743 1982 747 1986
rect 791 1982 795 1986
rect 815 1982 819 1986
rect 863 1982 867 1986
rect 935 1982 939 1986
rect 1007 1982 1011 1986
rect 1239 1982 1243 1986
rect 1279 1926 1283 1930
rect 1343 1926 1347 1930
rect 1383 1926 1387 1930
rect 1399 1926 1403 1930
rect 1423 1926 1427 1930
rect 1439 1926 1443 1930
rect 1463 1926 1467 1930
rect 1479 1926 1483 1930
rect 1511 1926 1515 1930
rect 1519 1926 1523 1930
rect 1559 1926 1563 1930
rect 1567 1926 1571 1930
rect 1599 1926 1603 1930
rect 1631 1926 1635 1930
rect 1639 1926 1643 1930
rect 1679 1926 1683 1930
rect 1711 1926 1715 1930
rect 1719 1926 1723 1930
rect 1767 1926 1771 1930
rect 1807 1926 1811 1930
rect 1823 1926 1827 1930
rect 1871 1926 1875 1930
rect 1919 1926 1923 1930
rect 1967 1926 1971 1930
rect 2015 1926 2019 1930
rect 2031 1926 2035 1930
rect 2055 1926 2059 1930
rect 2095 1926 2099 1930
rect 2143 1926 2147 1930
rect 2151 1926 2155 1930
rect 2191 1926 2195 1930
rect 2239 1926 2243 1930
rect 2279 1926 2283 1930
rect 2319 1926 2323 1930
rect 2359 1926 2363 1930
rect 2407 1926 2411 1930
rect 111 1910 115 1914
rect 135 1910 139 1914
rect 175 1910 179 1914
rect 215 1910 219 1914
rect 247 1910 251 1914
rect 271 1910 275 1914
rect 287 1910 291 1914
rect 327 1910 331 1914
rect 343 1910 347 1914
rect 367 1910 371 1914
rect 415 1910 419 1914
rect 471 1910 475 1914
rect 495 1910 499 1914
rect 535 1910 539 1914
rect 575 1910 579 1914
rect 599 1910 603 1914
rect 647 1910 651 1914
rect 663 1910 667 1914
rect 719 1910 723 1914
rect 727 1910 731 1914
rect 791 1910 795 1914
rect 855 1910 859 1914
rect 863 1910 867 1914
rect 919 1910 923 1914
rect 935 1910 939 1914
rect 983 1910 987 1914
rect 1007 1910 1011 1914
rect 1055 1910 1059 1914
rect 1127 1910 1131 1914
rect 1239 1910 1243 1914
rect 1279 1850 1283 1854
rect 1343 1850 1347 1854
rect 1359 1850 1363 1854
rect 1383 1850 1387 1854
rect 1399 1850 1403 1854
rect 1423 1850 1427 1854
rect 1447 1850 1451 1854
rect 1463 1850 1467 1854
rect 1503 1850 1507 1854
rect 1511 1850 1515 1854
rect 1559 1850 1563 1854
rect 1567 1850 1571 1854
rect 1615 1850 1619 1854
rect 1631 1850 1635 1854
rect 1671 1850 1675 1854
rect 1711 1850 1715 1854
rect 1727 1850 1731 1854
rect 1783 1850 1787 1854
rect 1807 1850 1811 1854
rect 1839 1850 1843 1854
rect 1895 1850 1899 1854
rect 1919 1850 1923 1854
rect 1951 1850 1955 1854
rect 2031 1850 2035 1854
rect 2151 1850 2155 1854
rect 2407 1850 2411 1854
rect 111 1838 115 1842
rect 247 1838 251 1842
rect 287 1838 291 1842
rect 327 1838 331 1842
rect 367 1838 371 1842
rect 399 1838 403 1842
rect 415 1838 419 1842
rect 439 1838 443 1842
rect 471 1838 475 1842
rect 479 1838 483 1842
rect 519 1838 523 1842
rect 535 1838 539 1842
rect 567 1838 571 1842
rect 599 1838 603 1842
rect 623 1838 627 1842
rect 663 1838 667 1842
rect 687 1838 691 1842
rect 727 1838 731 1842
rect 759 1838 763 1842
rect 791 1838 795 1842
rect 831 1838 835 1842
rect 855 1838 859 1842
rect 903 1838 907 1842
rect 919 1838 923 1842
rect 975 1838 979 1842
rect 983 1838 987 1842
rect 1047 1838 1051 1842
rect 1055 1838 1059 1842
rect 1127 1838 1131 1842
rect 1191 1838 1195 1842
rect 1239 1838 1243 1842
rect 111 1770 115 1774
rect 399 1770 403 1774
rect 407 1770 411 1774
rect 439 1770 443 1774
rect 447 1770 451 1774
rect 479 1770 483 1774
rect 487 1770 491 1774
rect 519 1770 523 1774
rect 527 1770 531 1774
rect 567 1770 571 1774
rect 607 1770 611 1774
rect 623 1770 627 1774
rect 647 1770 651 1774
rect 687 1770 691 1774
rect 695 1770 699 1774
rect 751 1770 755 1774
rect 759 1770 763 1774
rect 807 1770 811 1774
rect 831 1770 835 1774
rect 871 1770 875 1774
rect 903 1770 907 1774
rect 935 1770 939 1774
rect 975 1770 979 1774
rect 999 1770 1003 1774
rect 1047 1770 1051 1774
rect 1071 1770 1075 1774
rect 1127 1770 1131 1774
rect 1143 1770 1147 1774
rect 1191 1770 1195 1774
rect 1239 1770 1243 1774
rect 1279 1770 1283 1774
rect 1303 1770 1307 1774
rect 1343 1770 1347 1774
rect 1359 1770 1363 1774
rect 1391 1770 1395 1774
rect 1399 1770 1403 1774
rect 1447 1770 1451 1774
rect 1455 1770 1459 1774
rect 1503 1770 1507 1774
rect 1519 1770 1523 1774
rect 1559 1770 1563 1774
rect 1583 1770 1587 1774
rect 1615 1770 1619 1774
rect 1647 1770 1651 1774
rect 1671 1770 1675 1774
rect 1703 1770 1707 1774
rect 1727 1770 1731 1774
rect 1759 1770 1763 1774
rect 1783 1770 1787 1774
rect 1807 1770 1811 1774
rect 1839 1770 1843 1774
rect 1863 1770 1867 1774
rect 1895 1770 1899 1774
rect 1919 1770 1923 1774
rect 1951 1770 1955 1774
rect 1975 1770 1979 1774
rect 2407 1770 2411 1774
rect 111 1698 115 1702
rect 279 1698 283 1702
rect 319 1698 323 1702
rect 359 1698 363 1702
rect 399 1698 403 1702
rect 407 1698 411 1702
rect 447 1698 451 1702
rect 487 1698 491 1702
rect 495 1698 499 1702
rect 527 1698 531 1702
rect 543 1698 547 1702
rect 567 1698 571 1702
rect 591 1698 595 1702
rect 607 1698 611 1702
rect 639 1698 643 1702
rect 647 1698 651 1702
rect 687 1698 691 1702
rect 695 1698 699 1702
rect 735 1698 739 1702
rect 751 1698 755 1702
rect 783 1698 787 1702
rect 807 1698 811 1702
rect 839 1698 843 1702
rect 871 1698 875 1702
rect 895 1698 899 1702
rect 935 1698 939 1702
rect 999 1698 1003 1702
rect 1071 1698 1075 1702
rect 1143 1698 1147 1702
rect 1191 1698 1195 1702
rect 1239 1698 1243 1702
rect 1279 1698 1283 1702
rect 1303 1698 1307 1702
rect 1343 1698 1347 1702
rect 1383 1698 1387 1702
rect 1391 1698 1395 1702
rect 1423 1698 1427 1702
rect 1455 1698 1459 1702
rect 1463 1698 1467 1702
rect 1503 1698 1507 1702
rect 1519 1698 1523 1702
rect 1559 1698 1563 1702
rect 1583 1698 1587 1702
rect 1623 1698 1627 1702
rect 1647 1698 1651 1702
rect 1687 1698 1691 1702
rect 1703 1698 1707 1702
rect 1751 1698 1755 1702
rect 1759 1698 1763 1702
rect 1807 1698 1811 1702
rect 1863 1698 1867 1702
rect 1919 1698 1923 1702
rect 1975 1698 1979 1702
rect 2031 1698 2035 1702
rect 2087 1698 2091 1702
rect 2407 1698 2411 1702
rect 111 1626 115 1630
rect 135 1626 139 1630
rect 175 1626 179 1630
rect 215 1626 219 1630
rect 255 1626 259 1630
rect 279 1626 283 1630
rect 311 1626 315 1630
rect 319 1626 323 1630
rect 359 1626 363 1630
rect 391 1626 395 1630
rect 399 1626 403 1630
rect 447 1626 451 1630
rect 471 1626 475 1630
rect 495 1626 499 1630
rect 543 1626 547 1630
rect 559 1626 563 1630
rect 591 1626 595 1630
rect 639 1626 643 1630
rect 687 1626 691 1630
rect 719 1626 723 1630
rect 735 1626 739 1630
rect 783 1626 787 1630
rect 791 1626 795 1630
rect 839 1626 843 1630
rect 855 1626 859 1630
rect 895 1626 899 1630
rect 919 1626 923 1630
rect 983 1626 987 1630
rect 1047 1626 1051 1630
rect 1239 1626 1243 1630
rect 1279 1626 1283 1630
rect 1303 1626 1307 1630
rect 1343 1626 1347 1630
rect 1383 1626 1387 1630
rect 1423 1626 1427 1630
rect 1463 1626 1467 1630
rect 1503 1626 1507 1630
rect 1559 1626 1563 1630
rect 1623 1626 1627 1630
rect 1631 1626 1635 1630
rect 1687 1626 1691 1630
rect 1703 1626 1707 1630
rect 1751 1626 1755 1630
rect 1783 1626 1787 1630
rect 1807 1626 1811 1630
rect 1855 1626 1859 1630
rect 1863 1626 1867 1630
rect 1919 1626 1923 1630
rect 1927 1626 1931 1630
rect 1975 1626 1979 1630
rect 1999 1626 2003 1630
rect 2031 1626 2035 1630
rect 2063 1626 2067 1630
rect 2087 1626 2091 1630
rect 2127 1626 2131 1630
rect 2191 1626 2195 1630
rect 2255 1626 2259 1630
rect 2319 1626 2323 1630
rect 2359 1626 2363 1630
rect 2407 1626 2411 1630
rect 111 1554 115 1558
rect 135 1554 139 1558
rect 151 1554 155 1558
rect 175 1554 179 1558
rect 199 1554 203 1558
rect 215 1554 219 1558
rect 255 1554 259 1558
rect 263 1554 267 1558
rect 311 1554 315 1558
rect 343 1554 347 1558
rect 391 1554 395 1558
rect 439 1554 443 1558
rect 471 1554 475 1558
rect 535 1554 539 1558
rect 559 1554 563 1558
rect 639 1554 643 1558
rect 719 1554 723 1558
rect 735 1554 739 1558
rect 791 1554 795 1558
rect 823 1554 827 1558
rect 855 1554 859 1558
rect 903 1554 907 1558
rect 919 1554 923 1558
rect 975 1554 979 1558
rect 983 1554 987 1558
rect 1047 1554 1051 1558
rect 1119 1554 1123 1558
rect 1191 1554 1195 1558
rect 1239 1554 1243 1558
rect 1279 1558 1283 1562
rect 1303 1558 1307 1562
rect 1343 1558 1347 1562
rect 1383 1558 1387 1562
rect 1423 1558 1427 1562
rect 1463 1558 1467 1562
rect 1471 1558 1475 1562
rect 1503 1558 1507 1562
rect 1559 1558 1563 1562
rect 1623 1558 1627 1562
rect 1631 1558 1635 1562
rect 1703 1558 1707 1562
rect 1759 1558 1763 1562
rect 1783 1558 1787 1562
rect 1855 1558 1859 1562
rect 1871 1558 1875 1562
rect 1927 1558 1931 1562
rect 1967 1558 1971 1562
rect 1999 1558 2003 1562
rect 2055 1558 2059 1562
rect 2063 1558 2067 1562
rect 2127 1558 2131 1562
rect 2191 1558 2195 1562
rect 2255 1558 2259 1562
rect 2319 1558 2323 1562
rect 2359 1558 2363 1562
rect 2407 1558 2411 1562
rect 111 1482 115 1486
rect 151 1482 155 1486
rect 199 1482 203 1486
rect 263 1482 267 1486
rect 319 1482 323 1486
rect 343 1482 347 1486
rect 359 1482 363 1486
rect 399 1482 403 1486
rect 439 1482 443 1486
rect 447 1482 451 1486
rect 503 1482 507 1486
rect 535 1482 539 1486
rect 559 1482 563 1486
rect 615 1482 619 1486
rect 639 1482 643 1486
rect 671 1482 675 1486
rect 735 1482 739 1486
rect 799 1482 803 1486
rect 823 1482 827 1486
rect 855 1482 859 1486
rect 903 1482 907 1486
rect 911 1482 915 1486
rect 967 1482 971 1486
rect 975 1482 979 1486
rect 1023 1482 1027 1486
rect 1047 1482 1051 1486
rect 1087 1482 1091 1486
rect 1119 1482 1123 1486
rect 1151 1482 1155 1486
rect 1191 1482 1195 1486
rect 1239 1482 1243 1486
rect 1279 1470 1283 1474
rect 1303 1470 1307 1474
rect 1375 1470 1379 1474
rect 1471 1470 1475 1474
rect 1479 1470 1483 1474
rect 1583 1470 1587 1474
rect 1623 1470 1627 1474
rect 1687 1470 1691 1474
rect 1759 1470 1763 1474
rect 1783 1470 1787 1474
rect 1871 1470 1875 1474
rect 1951 1470 1955 1474
rect 1967 1470 1971 1474
rect 2031 1470 2035 1474
rect 2055 1470 2059 1474
rect 2103 1470 2107 1474
rect 2127 1470 2131 1474
rect 2167 1470 2171 1474
rect 2191 1470 2195 1474
rect 2239 1470 2243 1474
rect 2255 1470 2259 1474
rect 2311 1470 2315 1474
rect 2319 1470 2323 1474
rect 2359 1470 2363 1474
rect 2407 1470 2411 1474
rect 111 1410 115 1414
rect 263 1410 267 1414
rect 303 1410 307 1414
rect 319 1410 323 1414
rect 343 1410 347 1414
rect 359 1410 363 1414
rect 391 1410 395 1414
rect 399 1410 403 1414
rect 447 1410 451 1414
rect 503 1410 507 1414
rect 559 1410 563 1414
rect 615 1410 619 1414
rect 623 1410 627 1414
rect 671 1410 675 1414
rect 687 1410 691 1414
rect 735 1410 739 1414
rect 751 1410 755 1414
rect 799 1410 803 1414
rect 815 1410 819 1414
rect 855 1410 859 1414
rect 879 1410 883 1414
rect 911 1410 915 1414
rect 951 1410 955 1414
rect 967 1410 971 1414
rect 1023 1410 1027 1414
rect 1087 1410 1091 1414
rect 1151 1410 1155 1414
rect 1191 1410 1195 1414
rect 1239 1410 1243 1414
rect 1279 1402 1283 1406
rect 1303 1402 1307 1406
rect 1343 1402 1347 1406
rect 1375 1402 1379 1406
rect 1399 1402 1403 1406
rect 1471 1402 1475 1406
rect 1479 1402 1483 1406
rect 1551 1402 1555 1406
rect 1583 1402 1587 1406
rect 1639 1402 1643 1406
rect 1687 1402 1691 1406
rect 1727 1402 1731 1406
rect 1783 1402 1787 1406
rect 1815 1402 1819 1406
rect 1871 1402 1875 1406
rect 1903 1402 1907 1406
rect 1951 1402 1955 1406
rect 1991 1402 1995 1406
rect 2031 1402 2035 1406
rect 2071 1402 2075 1406
rect 2103 1402 2107 1406
rect 2151 1402 2155 1406
rect 2167 1402 2171 1406
rect 2223 1402 2227 1406
rect 2239 1402 2243 1406
rect 2303 1402 2307 1406
rect 2311 1402 2315 1406
rect 2359 1402 2363 1406
rect 2407 1402 2411 1406
rect 111 1338 115 1342
rect 135 1338 139 1342
rect 175 1338 179 1342
rect 215 1338 219 1342
rect 255 1338 259 1342
rect 263 1338 267 1342
rect 303 1338 307 1342
rect 327 1338 331 1342
rect 343 1338 347 1342
rect 391 1338 395 1342
rect 407 1338 411 1342
rect 447 1338 451 1342
rect 495 1338 499 1342
rect 503 1338 507 1342
rect 559 1338 563 1342
rect 583 1338 587 1342
rect 623 1338 627 1342
rect 671 1338 675 1342
rect 687 1338 691 1342
rect 751 1338 755 1342
rect 759 1338 763 1342
rect 815 1338 819 1342
rect 839 1338 843 1342
rect 879 1338 883 1342
rect 919 1338 923 1342
rect 951 1338 955 1342
rect 1007 1338 1011 1342
rect 1023 1338 1027 1342
rect 1095 1338 1099 1342
rect 1239 1338 1243 1342
rect 1279 1330 1283 1334
rect 1303 1330 1307 1334
rect 1343 1330 1347 1334
rect 1399 1330 1403 1334
rect 1447 1330 1451 1334
rect 1471 1330 1475 1334
rect 1487 1330 1491 1334
rect 1527 1330 1531 1334
rect 1551 1330 1555 1334
rect 1567 1330 1571 1334
rect 1615 1330 1619 1334
rect 1639 1330 1643 1334
rect 1671 1330 1675 1334
rect 1719 1330 1723 1334
rect 1727 1330 1731 1334
rect 1775 1330 1779 1334
rect 1815 1330 1819 1334
rect 1831 1330 1835 1334
rect 1903 1330 1907 1334
rect 1983 1330 1987 1334
rect 1991 1330 1995 1334
rect 2071 1330 2075 1334
rect 2151 1330 2155 1334
rect 2167 1330 2171 1334
rect 2223 1330 2227 1334
rect 2271 1330 2275 1334
rect 2303 1330 2307 1334
rect 2359 1330 2363 1334
rect 2407 1330 2411 1334
rect 111 1266 115 1270
rect 135 1266 139 1270
rect 175 1266 179 1270
rect 215 1266 219 1270
rect 247 1266 251 1270
rect 255 1266 259 1270
rect 327 1266 331 1270
rect 407 1266 411 1270
rect 415 1266 419 1270
rect 495 1266 499 1270
rect 503 1266 507 1270
rect 583 1266 587 1270
rect 591 1266 595 1270
rect 671 1266 675 1270
rect 743 1266 747 1270
rect 759 1266 763 1270
rect 815 1266 819 1270
rect 839 1266 843 1270
rect 879 1266 883 1270
rect 919 1266 923 1270
rect 943 1266 947 1270
rect 1007 1266 1011 1270
rect 1071 1266 1075 1270
rect 1095 1266 1099 1270
rect 1239 1266 1243 1270
rect 1279 1258 1283 1262
rect 1447 1258 1451 1262
rect 1487 1258 1491 1262
rect 1511 1258 1515 1262
rect 1527 1258 1531 1262
rect 1551 1258 1555 1262
rect 1567 1258 1571 1262
rect 1591 1258 1595 1262
rect 1615 1258 1619 1262
rect 1631 1258 1635 1262
rect 1671 1258 1675 1262
rect 1711 1258 1715 1262
rect 1719 1258 1723 1262
rect 1751 1258 1755 1262
rect 1775 1258 1779 1262
rect 1791 1258 1795 1262
rect 1831 1258 1835 1262
rect 1839 1258 1843 1262
rect 1903 1258 1907 1262
rect 1967 1258 1971 1262
rect 1983 1258 1987 1262
rect 2039 1258 2043 1262
rect 2071 1258 2075 1262
rect 2119 1258 2123 1262
rect 2167 1258 2171 1262
rect 2207 1258 2211 1262
rect 2271 1258 2275 1262
rect 2295 1258 2299 1262
rect 2359 1258 2363 1262
rect 2407 1258 2411 1262
rect 111 1190 115 1194
rect 135 1190 139 1194
rect 175 1190 179 1194
rect 231 1190 235 1194
rect 247 1190 251 1194
rect 303 1190 307 1194
rect 327 1190 331 1194
rect 383 1190 387 1194
rect 415 1190 419 1194
rect 471 1190 475 1194
rect 503 1190 507 1194
rect 559 1190 563 1194
rect 591 1190 595 1194
rect 639 1190 643 1194
rect 671 1190 675 1194
rect 719 1190 723 1194
rect 743 1190 747 1194
rect 799 1190 803 1194
rect 815 1190 819 1194
rect 871 1190 875 1194
rect 879 1190 883 1194
rect 935 1190 939 1194
rect 943 1190 947 1194
rect 991 1190 995 1194
rect 1007 1190 1011 1194
rect 1047 1190 1051 1194
rect 1071 1190 1075 1194
rect 1103 1190 1107 1194
rect 1151 1190 1155 1194
rect 1191 1190 1195 1194
rect 1239 1190 1243 1194
rect 1279 1186 1283 1190
rect 1511 1186 1515 1190
rect 1551 1186 1555 1190
rect 1559 1186 1563 1190
rect 1591 1186 1595 1190
rect 1599 1186 1603 1190
rect 1631 1186 1635 1190
rect 1639 1186 1643 1190
rect 1671 1186 1675 1190
rect 1679 1186 1683 1190
rect 1711 1186 1715 1190
rect 1719 1186 1723 1190
rect 1751 1186 1755 1190
rect 1759 1186 1763 1190
rect 1791 1186 1795 1190
rect 1799 1186 1803 1190
rect 1839 1186 1843 1190
rect 1855 1186 1859 1190
rect 1903 1186 1907 1190
rect 1927 1186 1931 1190
rect 1967 1186 1971 1190
rect 2023 1186 2027 1190
rect 2039 1186 2043 1190
rect 2119 1186 2123 1190
rect 2135 1186 2139 1190
rect 2207 1186 2211 1190
rect 2255 1186 2259 1190
rect 2295 1186 2299 1190
rect 2359 1186 2363 1190
rect 2407 1186 2411 1190
rect 111 1122 115 1126
rect 135 1122 139 1126
rect 175 1122 179 1126
rect 215 1122 219 1126
rect 231 1122 235 1126
rect 303 1122 307 1126
rect 383 1122 387 1126
rect 391 1122 395 1126
rect 471 1122 475 1126
rect 479 1122 483 1126
rect 559 1122 563 1126
rect 639 1122 643 1126
rect 711 1122 715 1126
rect 719 1122 723 1126
rect 775 1122 779 1126
rect 799 1122 803 1126
rect 839 1122 843 1126
rect 871 1122 875 1126
rect 903 1122 907 1126
rect 935 1122 939 1126
rect 959 1122 963 1126
rect 991 1122 995 1126
rect 1023 1122 1027 1126
rect 1047 1122 1051 1126
rect 1087 1122 1091 1126
rect 1103 1122 1107 1126
rect 1151 1122 1155 1126
rect 1191 1122 1195 1126
rect 1239 1122 1243 1126
rect 1279 1110 1283 1114
rect 1535 1110 1539 1114
rect 1559 1110 1563 1114
rect 1599 1110 1603 1114
rect 1639 1110 1643 1114
rect 1663 1110 1667 1114
rect 1679 1110 1683 1114
rect 1719 1110 1723 1114
rect 1727 1110 1731 1114
rect 1759 1110 1763 1114
rect 1791 1110 1795 1114
rect 1799 1110 1803 1114
rect 1855 1110 1859 1114
rect 1911 1110 1915 1114
rect 1927 1110 1931 1114
rect 1967 1110 1971 1114
rect 2023 1110 2027 1114
rect 2079 1110 2083 1114
rect 2135 1110 2139 1114
rect 2191 1110 2195 1114
rect 2255 1110 2259 1114
rect 2319 1110 2323 1114
rect 2359 1110 2363 1114
rect 2407 1110 2411 1114
rect 111 1050 115 1054
rect 135 1050 139 1054
rect 199 1050 203 1054
rect 215 1050 219 1054
rect 239 1050 243 1054
rect 287 1050 291 1054
rect 303 1050 307 1054
rect 343 1050 347 1054
rect 391 1050 395 1054
rect 439 1050 443 1054
rect 479 1050 483 1054
rect 487 1050 491 1054
rect 535 1050 539 1054
rect 559 1050 563 1054
rect 583 1050 587 1054
rect 631 1050 635 1054
rect 639 1050 643 1054
rect 679 1050 683 1054
rect 711 1050 715 1054
rect 727 1050 731 1054
rect 775 1050 779 1054
rect 783 1050 787 1054
rect 839 1050 843 1054
rect 895 1050 899 1054
rect 903 1050 907 1054
rect 959 1050 963 1054
rect 1023 1050 1027 1054
rect 1087 1050 1091 1054
rect 1151 1050 1155 1054
rect 1191 1050 1195 1054
rect 1239 1050 1243 1054
rect 1279 1030 1283 1034
rect 1503 1030 1507 1034
rect 1535 1030 1539 1034
rect 1599 1030 1603 1034
rect 1623 1030 1627 1034
rect 1663 1030 1667 1034
rect 1727 1030 1731 1034
rect 1735 1030 1739 1034
rect 1791 1030 1795 1034
rect 1831 1030 1835 1034
rect 1855 1030 1859 1034
rect 1911 1030 1915 1034
rect 1919 1030 1923 1034
rect 1967 1030 1971 1034
rect 1999 1030 2003 1034
rect 2023 1030 2027 1034
rect 2071 1030 2075 1034
rect 2079 1030 2083 1034
rect 2135 1030 2139 1034
rect 2143 1030 2147 1034
rect 2191 1030 2195 1034
rect 2207 1030 2211 1034
rect 2255 1030 2259 1034
rect 2279 1030 2283 1034
rect 2319 1030 2323 1034
rect 2359 1030 2363 1034
rect 2407 1030 2411 1034
rect 111 970 115 974
rect 199 970 203 974
rect 239 970 243 974
rect 287 970 291 974
rect 295 970 299 974
rect 343 970 347 974
rect 391 970 395 974
rect 399 970 403 974
rect 439 970 443 974
rect 471 970 475 974
rect 487 970 491 974
rect 535 970 539 974
rect 551 970 555 974
rect 583 970 587 974
rect 631 970 635 974
rect 639 970 643 974
rect 679 970 683 974
rect 727 970 731 974
rect 783 970 787 974
rect 807 970 811 974
rect 839 970 843 974
rect 887 970 891 974
rect 895 970 899 974
rect 959 970 963 974
rect 1023 970 1027 974
rect 1087 970 1091 974
rect 1151 970 1155 974
rect 1191 970 1195 974
rect 1239 970 1243 974
rect 1279 954 1283 958
rect 1319 954 1323 958
rect 1359 954 1363 958
rect 1399 954 1403 958
rect 1463 954 1467 958
rect 1503 954 1507 958
rect 1543 954 1547 958
rect 1623 954 1627 958
rect 1639 954 1643 958
rect 1735 954 1739 958
rect 1831 954 1835 958
rect 1839 954 1843 958
rect 1919 954 1923 958
rect 1935 954 1939 958
rect 1999 954 2003 958
rect 2023 954 2027 958
rect 2071 954 2075 958
rect 2103 954 2107 958
rect 2143 954 2147 958
rect 2175 954 2179 958
rect 2207 954 2211 958
rect 2239 954 2243 958
rect 2279 954 2283 958
rect 2311 954 2315 958
rect 2359 954 2363 958
rect 2407 954 2411 958
rect 111 894 115 898
rect 255 894 259 898
rect 295 894 299 898
rect 311 894 315 898
rect 343 894 347 898
rect 375 894 379 898
rect 399 894 403 898
rect 455 894 459 898
rect 471 894 475 898
rect 535 894 539 898
rect 551 894 555 898
rect 623 894 627 898
rect 639 894 643 898
rect 711 894 715 898
rect 727 894 731 898
rect 791 894 795 898
rect 807 894 811 898
rect 863 894 867 898
rect 887 894 891 898
rect 935 894 939 898
rect 959 894 963 898
rect 999 894 1003 898
rect 1023 894 1027 898
rect 1055 894 1059 898
rect 1087 894 1091 898
rect 1119 894 1123 898
rect 1151 894 1155 898
rect 1183 894 1187 898
rect 1191 894 1195 898
rect 1239 894 1243 898
rect 1279 878 1283 882
rect 1319 878 1323 882
rect 1335 878 1339 882
rect 1359 878 1363 882
rect 1375 878 1379 882
rect 1399 878 1403 882
rect 1415 878 1419 882
rect 1463 878 1467 882
rect 1471 878 1475 882
rect 1535 878 1539 882
rect 1543 878 1547 882
rect 1607 878 1611 882
rect 1639 878 1643 882
rect 1679 878 1683 882
rect 1735 878 1739 882
rect 1751 878 1755 882
rect 1823 878 1827 882
rect 1839 878 1843 882
rect 1895 878 1899 882
rect 1935 878 1939 882
rect 1959 878 1963 882
rect 2023 878 2027 882
rect 2087 878 2091 882
rect 2103 878 2107 882
rect 2143 878 2147 882
rect 2175 878 2179 882
rect 2199 878 2203 882
rect 2239 878 2243 882
rect 2255 878 2259 882
rect 2311 878 2315 882
rect 2319 878 2323 882
rect 2359 878 2363 882
rect 2407 878 2411 882
rect 111 826 115 830
rect 191 826 195 830
rect 247 826 251 830
rect 255 826 259 830
rect 311 826 315 830
rect 375 826 379 830
rect 383 826 387 830
rect 455 826 459 830
rect 463 826 467 830
rect 535 826 539 830
rect 543 826 547 830
rect 615 826 619 830
rect 623 826 627 830
rect 687 826 691 830
rect 711 826 715 830
rect 751 826 755 830
rect 791 826 795 830
rect 815 826 819 830
rect 863 826 867 830
rect 871 826 875 830
rect 927 826 931 830
rect 935 826 939 830
rect 983 826 987 830
rect 999 826 1003 830
rect 1047 826 1051 830
rect 1055 826 1059 830
rect 1119 826 1123 830
rect 1183 826 1187 830
rect 1239 826 1243 830
rect 1279 806 1283 810
rect 1303 806 1307 810
rect 1335 806 1339 810
rect 1343 806 1347 810
rect 1375 806 1379 810
rect 1407 806 1411 810
rect 1415 806 1419 810
rect 1471 806 1475 810
rect 1479 806 1483 810
rect 1535 806 1539 810
rect 1551 806 1555 810
rect 1607 806 1611 810
rect 1623 806 1627 810
rect 1679 806 1683 810
rect 1695 806 1699 810
rect 1751 806 1755 810
rect 1759 806 1763 810
rect 1823 806 1827 810
rect 1887 806 1891 810
rect 1895 806 1899 810
rect 1951 806 1955 810
rect 1959 806 1963 810
rect 2023 806 2027 810
rect 2087 806 2091 810
rect 2103 806 2107 810
rect 2143 806 2147 810
rect 2191 806 2195 810
rect 2199 806 2203 810
rect 2255 806 2259 810
rect 2279 806 2283 810
rect 2319 806 2323 810
rect 2359 806 2363 810
rect 2407 806 2411 810
rect 111 758 115 762
rect 135 758 139 762
rect 175 758 179 762
rect 191 758 195 762
rect 215 758 219 762
rect 247 758 251 762
rect 279 758 283 762
rect 311 758 315 762
rect 351 758 355 762
rect 383 758 387 762
rect 423 758 427 762
rect 463 758 467 762
rect 495 758 499 762
rect 543 758 547 762
rect 559 758 563 762
rect 615 758 619 762
rect 623 758 627 762
rect 687 758 691 762
rect 695 758 699 762
rect 751 758 755 762
rect 783 758 787 762
rect 815 758 819 762
rect 871 758 875 762
rect 879 758 883 762
rect 927 758 931 762
rect 983 758 987 762
rect 1047 758 1051 762
rect 1095 758 1099 762
rect 1191 758 1195 762
rect 1239 758 1243 762
rect 1279 738 1283 742
rect 1303 738 1307 742
rect 1343 738 1347 742
rect 1367 738 1371 742
rect 1407 738 1411 742
rect 1455 738 1459 742
rect 1479 738 1483 742
rect 1535 738 1539 742
rect 1551 738 1555 742
rect 1615 738 1619 742
rect 1623 738 1627 742
rect 1695 738 1699 742
rect 1759 738 1763 742
rect 1775 738 1779 742
rect 1823 738 1827 742
rect 1855 738 1859 742
rect 1887 738 1891 742
rect 1943 738 1947 742
rect 1951 738 1955 742
rect 2023 738 2027 742
rect 2031 738 2035 742
rect 2103 738 2107 742
rect 2119 738 2123 742
rect 2191 738 2195 742
rect 2207 738 2211 742
rect 2279 738 2283 742
rect 2295 738 2299 742
rect 2359 738 2363 742
rect 2407 738 2411 742
rect 111 682 115 686
rect 135 682 139 686
rect 175 682 179 686
rect 215 682 219 686
rect 231 682 235 686
rect 279 682 283 686
rect 287 682 291 686
rect 343 682 347 686
rect 351 682 355 686
rect 399 682 403 686
rect 423 682 427 686
rect 455 682 459 686
rect 495 682 499 686
rect 503 682 507 686
rect 559 682 563 686
rect 623 682 627 686
rect 695 682 699 686
rect 767 682 771 686
rect 783 682 787 686
rect 839 682 843 686
rect 879 682 883 686
rect 903 682 907 686
rect 967 682 971 686
rect 983 682 987 686
rect 1023 682 1027 686
rect 1087 682 1091 686
rect 1095 682 1099 686
rect 1151 682 1155 686
rect 1191 682 1195 686
rect 1239 682 1243 686
rect 1279 670 1283 674
rect 1303 670 1307 674
rect 1367 670 1371 674
rect 1455 670 1459 674
rect 1535 670 1539 674
rect 1591 670 1595 674
rect 1615 670 1619 674
rect 1639 670 1643 674
rect 1687 670 1691 674
rect 1695 670 1699 674
rect 1743 670 1747 674
rect 1775 670 1779 674
rect 1799 670 1803 674
rect 1855 670 1859 674
rect 1871 670 1875 674
rect 1943 670 1947 674
rect 1951 670 1955 674
rect 2031 670 2035 674
rect 2047 670 2051 674
rect 2119 670 2123 674
rect 2151 670 2155 674
rect 2207 670 2211 674
rect 2263 670 2267 674
rect 2295 670 2299 674
rect 2359 670 2363 674
rect 2407 670 2411 674
rect 111 614 115 618
rect 135 614 139 618
rect 175 614 179 618
rect 183 614 187 618
rect 231 614 235 618
rect 255 614 259 618
rect 287 614 291 618
rect 327 614 331 618
rect 343 614 347 618
rect 399 614 403 618
rect 455 614 459 618
rect 479 614 483 618
rect 503 614 507 618
rect 559 614 563 618
rect 623 614 627 618
rect 639 614 643 618
rect 695 614 699 618
rect 719 614 723 618
rect 767 614 771 618
rect 799 614 803 618
rect 839 614 843 618
rect 879 614 883 618
rect 903 614 907 618
rect 951 614 955 618
rect 967 614 971 618
rect 1015 614 1019 618
rect 1023 614 1027 618
rect 1079 614 1083 618
rect 1087 614 1091 618
rect 1143 614 1147 618
rect 1151 614 1155 618
rect 1191 614 1195 618
rect 1239 614 1243 618
rect 1279 594 1283 598
rect 1559 594 1563 598
rect 1591 594 1595 598
rect 1599 594 1603 598
rect 1639 594 1643 598
rect 1679 594 1683 598
rect 1687 594 1691 598
rect 1719 594 1723 598
rect 1743 594 1747 598
rect 1759 594 1763 598
rect 1799 594 1803 598
rect 1807 594 1811 598
rect 1855 594 1859 598
rect 1871 594 1875 598
rect 1911 594 1915 598
rect 1951 594 1955 598
rect 1967 594 1971 598
rect 2031 594 2035 598
rect 2047 594 2051 598
rect 2095 594 2099 598
rect 2151 594 2155 598
rect 2167 594 2171 598
rect 2239 594 2243 598
rect 2263 594 2267 598
rect 2311 594 2315 598
rect 2359 594 2363 598
rect 2407 594 2411 598
rect 111 542 115 546
rect 135 542 139 546
rect 151 542 155 546
rect 183 542 187 546
rect 223 542 227 546
rect 255 542 259 546
rect 287 542 291 546
rect 327 542 331 546
rect 351 542 355 546
rect 399 542 403 546
rect 415 542 419 546
rect 479 542 483 546
rect 551 542 555 546
rect 559 542 563 546
rect 623 542 627 546
rect 639 542 643 546
rect 695 542 699 546
rect 719 542 723 546
rect 767 542 771 546
rect 799 542 803 546
rect 839 542 843 546
rect 879 542 883 546
rect 919 542 923 546
rect 951 542 955 546
rect 999 542 1003 546
rect 1015 542 1019 546
rect 1079 542 1083 546
rect 1143 542 1147 546
rect 1191 542 1195 546
rect 1239 542 1243 546
rect 1279 526 1283 530
rect 1407 526 1411 530
rect 1447 526 1451 530
rect 1487 526 1491 530
rect 1535 526 1539 530
rect 1559 526 1563 530
rect 1591 526 1595 530
rect 1599 526 1603 530
rect 1639 526 1643 530
rect 1647 526 1651 530
rect 1679 526 1683 530
rect 1711 526 1715 530
rect 1719 526 1723 530
rect 1759 526 1763 530
rect 1783 526 1787 530
rect 1807 526 1811 530
rect 1855 526 1859 530
rect 1863 526 1867 530
rect 1911 526 1915 530
rect 1943 526 1947 530
rect 1967 526 1971 530
rect 2023 526 2027 530
rect 2031 526 2035 530
rect 2095 526 2099 530
rect 2103 526 2107 530
rect 2167 526 2171 530
rect 2191 526 2195 530
rect 2239 526 2243 530
rect 2287 526 2291 530
rect 2311 526 2315 530
rect 2359 526 2363 530
rect 2407 526 2411 530
rect 111 474 115 478
rect 151 474 155 478
rect 223 474 227 478
rect 239 474 243 478
rect 279 474 283 478
rect 287 474 291 478
rect 327 474 331 478
rect 351 474 355 478
rect 383 474 387 478
rect 415 474 419 478
rect 439 474 443 478
rect 479 474 483 478
rect 503 474 507 478
rect 551 474 555 478
rect 567 474 571 478
rect 623 474 627 478
rect 631 474 635 478
rect 695 474 699 478
rect 759 474 763 478
rect 767 474 771 478
rect 823 474 827 478
rect 839 474 843 478
rect 887 474 891 478
rect 919 474 923 478
rect 951 474 955 478
rect 999 474 1003 478
rect 1015 474 1019 478
rect 1079 474 1083 478
rect 1239 474 1243 478
rect 1279 458 1283 462
rect 1303 458 1307 462
rect 1343 458 1347 462
rect 1383 458 1387 462
rect 1407 458 1411 462
rect 1447 458 1451 462
rect 1487 458 1491 462
rect 1535 458 1539 462
rect 1591 458 1595 462
rect 1631 458 1635 462
rect 1647 458 1651 462
rect 1711 458 1715 462
rect 1735 458 1739 462
rect 1783 458 1787 462
rect 1831 458 1835 462
rect 1863 458 1867 462
rect 1919 458 1923 462
rect 1943 458 1947 462
rect 1999 458 2003 462
rect 2023 458 2027 462
rect 2071 458 2075 462
rect 2103 458 2107 462
rect 2135 458 2139 462
rect 2191 458 2195 462
rect 2199 458 2203 462
rect 2255 458 2259 462
rect 2287 458 2291 462
rect 2319 458 2323 462
rect 2359 458 2363 462
rect 2407 458 2411 462
rect 111 402 115 406
rect 143 402 147 406
rect 183 402 187 406
rect 223 402 227 406
rect 239 402 243 406
rect 271 402 275 406
rect 279 402 283 406
rect 327 402 331 406
rect 335 402 339 406
rect 383 402 387 406
rect 399 402 403 406
rect 439 402 443 406
rect 471 402 475 406
rect 503 402 507 406
rect 543 402 547 406
rect 567 402 571 406
rect 615 402 619 406
rect 631 402 635 406
rect 687 402 691 406
rect 695 402 699 406
rect 751 402 755 406
rect 759 402 763 406
rect 807 402 811 406
rect 823 402 827 406
rect 863 402 867 406
rect 887 402 891 406
rect 919 402 923 406
rect 951 402 955 406
rect 975 402 979 406
rect 1015 402 1019 406
rect 1031 402 1035 406
rect 1239 402 1243 406
rect 1279 390 1283 394
rect 1303 390 1307 394
rect 1343 390 1347 394
rect 1359 390 1363 394
rect 1383 390 1387 394
rect 1399 390 1403 394
rect 1439 390 1443 394
rect 1447 390 1451 394
rect 1487 390 1491 394
rect 1535 390 1539 394
rect 1543 390 1547 394
rect 1607 390 1611 394
rect 1631 390 1635 394
rect 1679 390 1683 394
rect 1735 390 1739 394
rect 1759 390 1763 394
rect 1831 390 1835 394
rect 1839 390 1843 394
rect 1919 390 1923 394
rect 1999 390 2003 394
rect 2071 390 2075 394
rect 2079 390 2083 394
rect 2135 390 2139 394
rect 2159 390 2163 394
rect 2199 390 2203 394
rect 2247 390 2251 394
rect 2255 390 2259 394
rect 2319 390 2323 394
rect 2335 390 2339 394
rect 2359 390 2363 394
rect 2407 390 2411 394
rect 111 326 115 330
rect 135 326 139 330
rect 143 326 147 330
rect 175 326 179 330
rect 183 326 187 330
rect 215 326 219 330
rect 223 326 227 330
rect 255 326 259 330
rect 271 326 275 330
rect 295 326 299 330
rect 335 326 339 330
rect 391 326 395 330
rect 399 326 403 330
rect 447 326 451 330
rect 471 326 475 330
rect 495 326 499 330
rect 543 326 547 330
rect 591 326 595 330
rect 615 326 619 330
rect 639 326 643 330
rect 687 326 691 330
rect 735 326 739 330
rect 751 326 755 330
rect 783 326 787 330
rect 807 326 811 330
rect 839 326 843 330
rect 863 326 867 330
rect 919 326 923 330
rect 975 326 979 330
rect 1031 326 1035 330
rect 1239 326 1243 330
rect 1279 314 1283 318
rect 1359 314 1363 318
rect 1399 314 1403 318
rect 1439 314 1443 318
rect 1487 314 1491 318
rect 1511 314 1515 318
rect 1543 314 1547 318
rect 1551 314 1555 318
rect 1591 314 1595 318
rect 1607 314 1611 318
rect 1631 314 1635 318
rect 1671 314 1675 318
rect 1679 314 1683 318
rect 1711 314 1715 318
rect 1751 314 1755 318
rect 1759 314 1763 318
rect 1791 314 1795 318
rect 1839 314 1843 318
rect 1903 314 1907 318
rect 1919 314 1923 318
rect 1967 314 1971 318
rect 1999 314 2003 318
rect 2039 314 2043 318
rect 2079 314 2083 318
rect 2119 314 2123 318
rect 2159 314 2163 318
rect 2199 314 2203 318
rect 2247 314 2251 318
rect 2279 314 2283 318
rect 2335 314 2339 318
rect 2359 314 2363 318
rect 2407 314 2411 318
rect 111 250 115 254
rect 135 250 139 254
rect 175 250 179 254
rect 215 250 219 254
rect 223 250 227 254
rect 255 250 259 254
rect 295 250 299 254
rect 311 250 315 254
rect 335 250 339 254
rect 391 250 395 254
rect 447 250 451 254
rect 463 250 467 254
rect 495 250 499 254
rect 527 250 531 254
rect 543 250 547 254
rect 591 250 595 254
rect 639 250 643 254
rect 647 250 651 254
rect 687 250 691 254
rect 695 250 699 254
rect 735 250 739 254
rect 783 250 787 254
rect 831 250 835 254
rect 839 250 843 254
rect 879 250 883 254
rect 927 250 931 254
rect 975 250 979 254
rect 1023 250 1027 254
rect 1239 250 1243 254
rect 1279 242 1283 246
rect 1367 242 1371 246
rect 1407 242 1411 246
rect 1455 242 1459 246
rect 1511 242 1515 246
rect 1551 242 1555 246
rect 1567 242 1571 246
rect 1591 242 1595 246
rect 1631 242 1635 246
rect 1671 242 1675 246
rect 1703 242 1707 246
rect 1711 242 1715 246
rect 1751 242 1755 246
rect 1775 242 1779 246
rect 1791 242 1795 246
rect 1839 242 1843 246
rect 1855 242 1859 246
rect 1903 242 1907 246
rect 1943 242 1947 246
rect 1967 242 1971 246
rect 2031 242 2035 246
rect 2039 242 2043 246
rect 2119 242 2123 246
rect 2199 242 2203 246
rect 2207 242 2211 246
rect 2279 242 2283 246
rect 2295 242 2299 246
rect 2359 242 2363 246
rect 2407 242 2411 246
rect 1279 166 1283 170
rect 1303 166 1307 170
rect 1343 166 1347 170
rect 1367 166 1371 170
rect 1383 166 1387 170
rect 1407 166 1411 170
rect 1423 166 1427 170
rect 1455 166 1459 170
rect 1463 166 1467 170
rect 1511 166 1515 170
rect 1519 166 1523 170
rect 1567 166 1571 170
rect 1583 166 1587 170
rect 1631 166 1635 170
rect 1647 166 1651 170
rect 1703 166 1707 170
rect 1711 166 1715 170
rect 1775 166 1779 170
rect 1831 166 1835 170
rect 1855 166 1859 170
rect 1887 166 1891 170
rect 1935 166 1939 170
rect 1943 166 1947 170
rect 1975 166 1979 170
rect 2015 166 2019 170
rect 2031 166 2035 170
rect 2055 166 2059 170
rect 2095 166 2099 170
rect 2119 166 2123 170
rect 2143 166 2147 170
rect 2191 166 2195 170
rect 2207 166 2211 170
rect 2239 166 2243 170
rect 2279 166 2283 170
rect 2295 166 2299 170
rect 2319 166 2323 170
rect 2359 166 2363 170
rect 2407 166 2411 170
rect 111 150 115 154
rect 135 150 139 154
rect 151 150 155 154
rect 191 150 195 154
rect 223 150 227 154
rect 231 150 235 154
rect 271 150 275 154
rect 311 150 315 154
rect 351 150 355 154
rect 391 150 395 154
rect 431 150 435 154
rect 463 150 467 154
rect 471 150 475 154
rect 511 150 515 154
rect 527 150 531 154
rect 551 150 555 154
rect 591 150 595 154
rect 631 150 635 154
rect 647 150 651 154
rect 671 150 675 154
rect 695 150 699 154
rect 711 150 715 154
rect 735 150 739 154
rect 751 150 755 154
rect 783 150 787 154
rect 791 150 795 154
rect 831 150 835 154
rect 871 150 875 154
rect 879 150 883 154
rect 911 150 915 154
rect 927 150 931 154
rect 951 150 955 154
rect 975 150 979 154
rect 991 150 995 154
rect 1023 150 1027 154
rect 1031 150 1035 154
rect 1071 150 1075 154
rect 1111 150 1115 154
rect 1151 150 1155 154
rect 1191 150 1195 154
rect 1239 150 1243 154
rect 1279 98 1283 102
rect 1303 98 1307 102
rect 1343 98 1347 102
rect 1383 98 1387 102
rect 1423 98 1427 102
rect 1463 98 1467 102
rect 1519 98 1523 102
rect 1583 98 1587 102
rect 1647 98 1651 102
rect 1711 98 1715 102
rect 1775 98 1779 102
rect 1831 98 1835 102
rect 1887 98 1891 102
rect 1935 98 1939 102
rect 1975 98 1979 102
rect 2015 98 2019 102
rect 2055 98 2059 102
rect 2095 98 2099 102
rect 2143 98 2147 102
rect 2191 98 2195 102
rect 2239 98 2243 102
rect 2279 98 2283 102
rect 2319 98 2323 102
rect 2359 98 2363 102
rect 2407 98 2411 102
rect 111 82 115 86
rect 151 82 155 86
rect 191 82 195 86
rect 231 82 235 86
rect 271 82 275 86
rect 311 82 315 86
rect 351 82 355 86
rect 391 82 395 86
rect 431 82 435 86
rect 471 82 475 86
rect 511 82 515 86
rect 551 82 555 86
rect 591 82 595 86
rect 631 82 635 86
rect 671 82 675 86
rect 711 82 715 86
rect 751 82 755 86
rect 791 82 795 86
rect 831 82 835 86
rect 871 82 875 86
rect 911 82 915 86
rect 951 82 955 86
rect 991 82 995 86
rect 1031 82 1035 86
rect 1071 82 1075 86
rect 1111 82 1115 86
rect 1151 82 1155 86
rect 1191 82 1195 86
rect 1239 82 1243 86
<< m4 >>
rect 96 2489 97 2495
rect 103 2494 1263 2495
rect 103 2490 111 2494
rect 115 2490 231 2494
rect 235 2490 271 2494
rect 275 2490 311 2494
rect 315 2490 351 2494
rect 355 2490 399 2494
rect 403 2490 455 2494
rect 459 2490 511 2494
rect 515 2490 575 2494
rect 579 2490 639 2494
rect 643 2490 703 2494
rect 707 2490 767 2494
rect 771 2490 823 2494
rect 827 2490 879 2494
rect 883 2490 927 2494
rect 931 2490 975 2494
rect 979 2490 1023 2494
rect 1027 2490 1071 2494
rect 1075 2490 1111 2494
rect 1115 2490 1151 2494
rect 1155 2490 1191 2494
rect 1195 2490 1239 2494
rect 1243 2490 1263 2494
rect 103 2489 1263 2490
rect 1269 2491 1270 2495
rect 1269 2490 2454 2491
rect 1269 2489 1279 2490
rect 1262 2486 1279 2489
rect 1283 2486 1303 2490
rect 1307 2486 1343 2490
rect 1347 2486 1383 2490
rect 1387 2486 1439 2490
rect 1443 2486 1511 2490
rect 1515 2486 1583 2490
rect 1587 2486 1663 2490
rect 1667 2486 1735 2490
rect 1739 2486 1807 2490
rect 1811 2486 1887 2490
rect 1891 2486 1967 2490
rect 1971 2486 2063 2490
rect 2067 2486 2167 2490
rect 2171 2486 2271 2490
rect 2275 2486 2359 2490
rect 2363 2486 2407 2490
rect 2411 2486 2454 2490
rect 1262 2485 2454 2486
rect 1250 2422 2442 2423
rect 1250 2419 1279 2422
rect 84 2413 85 2419
rect 91 2418 1251 2419
rect 91 2414 111 2418
rect 115 2414 199 2418
rect 203 2414 231 2418
rect 235 2414 263 2418
rect 267 2414 271 2418
rect 275 2414 311 2418
rect 315 2414 327 2418
rect 331 2414 351 2418
rect 355 2414 399 2418
rect 403 2414 455 2418
rect 459 2414 471 2418
rect 475 2414 511 2418
rect 515 2414 543 2418
rect 547 2414 575 2418
rect 579 2414 615 2418
rect 619 2414 639 2418
rect 643 2414 687 2418
rect 691 2414 703 2418
rect 707 2414 751 2418
rect 755 2414 767 2418
rect 771 2414 823 2418
rect 827 2414 879 2418
rect 883 2414 895 2418
rect 899 2414 927 2418
rect 931 2414 967 2418
rect 971 2414 975 2418
rect 979 2414 1023 2418
rect 1027 2414 1071 2418
rect 1075 2414 1111 2418
rect 1115 2414 1151 2418
rect 1155 2414 1191 2418
rect 1195 2414 1239 2418
rect 1243 2414 1251 2418
rect 91 2413 1251 2414
rect 1257 2418 1279 2419
rect 1283 2418 1303 2422
rect 1307 2418 1343 2422
rect 1347 2418 1375 2422
rect 1379 2418 1383 2422
rect 1387 2418 1415 2422
rect 1419 2418 1439 2422
rect 1443 2418 1455 2422
rect 1459 2418 1503 2422
rect 1507 2418 1511 2422
rect 1515 2418 1559 2422
rect 1563 2418 1583 2422
rect 1587 2418 1615 2422
rect 1619 2418 1663 2422
rect 1667 2418 1679 2422
rect 1683 2418 1735 2422
rect 1739 2418 1799 2422
rect 1803 2418 1807 2422
rect 1811 2418 1871 2422
rect 1875 2418 1887 2422
rect 1891 2418 1951 2422
rect 1955 2418 1967 2422
rect 1971 2418 2047 2422
rect 2051 2418 2063 2422
rect 2067 2418 2151 2422
rect 2155 2418 2167 2422
rect 2171 2418 2263 2422
rect 2267 2418 2271 2422
rect 2275 2418 2359 2422
rect 2363 2418 2407 2422
rect 2411 2418 2442 2422
rect 1257 2417 2442 2418
rect 1257 2413 1258 2417
rect 1262 2350 2454 2351
rect 1262 2347 1279 2350
rect 96 2341 97 2347
rect 103 2346 1263 2347
rect 103 2342 111 2346
rect 115 2342 199 2346
rect 203 2342 263 2346
rect 267 2342 271 2346
rect 275 2342 327 2346
rect 331 2342 399 2346
rect 403 2342 471 2346
rect 475 2342 543 2346
rect 547 2342 551 2346
rect 555 2342 615 2346
rect 619 2342 631 2346
rect 635 2342 687 2346
rect 691 2342 711 2346
rect 715 2342 751 2346
rect 755 2342 783 2346
rect 787 2342 823 2346
rect 827 2342 855 2346
rect 859 2342 895 2346
rect 899 2342 919 2346
rect 923 2342 967 2346
rect 971 2342 991 2346
rect 995 2342 1063 2346
rect 1067 2342 1239 2346
rect 1243 2342 1263 2346
rect 103 2341 1263 2342
rect 1269 2346 1279 2347
rect 1283 2346 1327 2350
rect 1331 2346 1375 2350
rect 1379 2346 1383 2350
rect 1387 2346 1415 2350
rect 1419 2346 1439 2350
rect 1443 2346 1455 2350
rect 1459 2346 1503 2350
rect 1507 2346 1559 2350
rect 1563 2346 1575 2350
rect 1579 2346 1615 2350
rect 1619 2346 1647 2350
rect 1651 2346 1679 2350
rect 1683 2346 1719 2350
rect 1723 2346 1735 2350
rect 1739 2346 1799 2350
rect 1803 2346 1871 2350
rect 1875 2346 1879 2350
rect 1883 2346 1951 2350
rect 1955 2346 1967 2350
rect 1971 2346 2047 2350
rect 2051 2346 2063 2350
rect 2067 2346 2151 2350
rect 2155 2346 2167 2350
rect 2171 2346 2263 2350
rect 2267 2346 2271 2350
rect 2275 2346 2359 2350
rect 2363 2346 2407 2350
rect 2411 2346 2454 2350
rect 1269 2345 2454 2346
rect 1269 2341 1270 2345
rect 1250 2277 1251 2283
rect 1257 2282 2435 2283
rect 1257 2278 1279 2282
rect 1283 2278 1327 2282
rect 1331 2278 1335 2282
rect 1339 2278 1383 2282
rect 1387 2278 1407 2282
rect 1411 2278 1439 2282
rect 1443 2278 1487 2282
rect 1491 2278 1503 2282
rect 1507 2278 1559 2282
rect 1563 2278 1575 2282
rect 1579 2278 1631 2282
rect 1635 2278 1647 2282
rect 1651 2278 1703 2282
rect 1707 2278 1719 2282
rect 1723 2278 1775 2282
rect 1779 2278 1799 2282
rect 1803 2278 1839 2282
rect 1843 2278 1879 2282
rect 1883 2278 1911 2282
rect 1915 2278 1967 2282
rect 1971 2278 1991 2282
rect 1995 2278 2063 2282
rect 2067 2278 2079 2282
rect 2083 2278 2167 2282
rect 2171 2278 2175 2282
rect 2179 2278 2271 2282
rect 2275 2278 2279 2282
rect 2283 2278 2359 2282
rect 2363 2278 2407 2282
rect 2411 2278 2435 2282
rect 1257 2277 2435 2278
rect 2441 2277 2442 2283
rect 84 2265 85 2271
rect 91 2270 1251 2271
rect 91 2266 111 2270
rect 115 2266 143 2270
rect 147 2266 183 2270
rect 187 2266 223 2270
rect 227 2266 271 2270
rect 275 2266 279 2270
rect 283 2266 327 2270
rect 331 2266 335 2270
rect 339 2266 399 2270
rect 403 2266 407 2270
rect 411 2266 471 2270
rect 475 2266 479 2270
rect 483 2266 551 2270
rect 555 2266 559 2270
rect 563 2266 631 2270
rect 635 2266 647 2270
rect 651 2266 711 2270
rect 715 2266 727 2270
rect 731 2266 783 2270
rect 787 2266 807 2270
rect 811 2266 855 2270
rect 859 2266 887 2270
rect 891 2266 919 2270
rect 923 2266 967 2270
rect 971 2266 991 2270
rect 995 2266 1047 2270
rect 1051 2266 1063 2270
rect 1067 2266 1127 2270
rect 1131 2266 1239 2270
rect 1243 2266 1251 2270
rect 91 2265 1251 2266
rect 1257 2265 1258 2271
rect 1262 2206 2454 2207
rect 1262 2203 1279 2206
rect 96 2197 97 2203
rect 103 2202 1263 2203
rect 103 2198 111 2202
rect 115 2198 135 2202
rect 139 2198 143 2202
rect 147 2198 183 2202
rect 187 2198 207 2202
rect 211 2198 223 2202
rect 227 2198 279 2202
rect 283 2198 335 2202
rect 339 2198 359 2202
rect 363 2198 407 2202
rect 411 2198 439 2202
rect 443 2198 479 2202
rect 483 2198 519 2202
rect 523 2198 559 2202
rect 563 2198 599 2202
rect 603 2198 647 2202
rect 651 2198 679 2202
rect 683 2198 727 2202
rect 731 2198 759 2202
rect 763 2198 807 2202
rect 811 2198 831 2202
rect 835 2198 887 2202
rect 891 2198 903 2202
rect 907 2198 967 2202
rect 971 2198 975 2202
rect 979 2198 1047 2202
rect 1051 2198 1119 2202
rect 1123 2198 1127 2202
rect 1131 2198 1239 2202
rect 1243 2198 1263 2202
rect 103 2197 1263 2198
rect 1269 2202 1279 2203
rect 1283 2202 1335 2206
rect 1339 2202 1375 2206
rect 1379 2202 1407 2206
rect 1411 2202 1439 2206
rect 1443 2202 1487 2206
rect 1491 2202 1511 2206
rect 1515 2202 1559 2206
rect 1563 2202 1591 2206
rect 1595 2202 1631 2206
rect 1635 2202 1671 2206
rect 1675 2202 1703 2206
rect 1707 2202 1751 2206
rect 1755 2202 1775 2206
rect 1779 2202 1831 2206
rect 1835 2202 1839 2206
rect 1843 2202 1903 2206
rect 1907 2202 1911 2206
rect 1915 2202 1967 2206
rect 1971 2202 1991 2206
rect 1995 2202 2031 2206
rect 2035 2202 2079 2206
rect 2083 2202 2095 2206
rect 2099 2202 2167 2206
rect 2171 2202 2175 2206
rect 2179 2202 2239 2206
rect 2243 2202 2279 2206
rect 2283 2202 2311 2206
rect 2315 2202 2359 2206
rect 2363 2202 2407 2206
rect 2411 2202 2454 2206
rect 1269 2201 2454 2202
rect 1269 2197 1270 2201
rect 1250 2133 1251 2139
rect 1257 2138 2435 2139
rect 1257 2134 1279 2138
rect 1283 2134 1375 2138
rect 1379 2134 1399 2138
rect 1403 2134 1439 2138
rect 1443 2134 1495 2138
rect 1499 2134 1511 2138
rect 1515 2134 1567 2138
rect 1571 2134 1591 2138
rect 1595 2134 1647 2138
rect 1651 2134 1671 2138
rect 1675 2134 1735 2138
rect 1739 2134 1751 2138
rect 1755 2134 1823 2138
rect 1827 2134 1831 2138
rect 1835 2134 1903 2138
rect 1907 2134 1911 2138
rect 1915 2134 1967 2138
rect 1971 2134 1999 2138
rect 2003 2134 2031 2138
rect 2035 2134 2087 2138
rect 2091 2134 2095 2138
rect 2099 2134 2167 2138
rect 2171 2134 2175 2138
rect 2179 2134 2239 2138
rect 2243 2134 2271 2138
rect 2275 2134 2311 2138
rect 2315 2134 2359 2138
rect 2363 2134 2407 2138
rect 2411 2134 2435 2138
rect 1257 2133 2435 2134
rect 2441 2133 2442 2139
rect 84 2121 85 2127
rect 91 2126 1251 2127
rect 91 2122 111 2126
rect 115 2122 135 2126
rect 139 2122 191 2126
rect 195 2122 207 2126
rect 211 2122 271 2126
rect 275 2122 279 2126
rect 283 2122 343 2126
rect 347 2122 359 2126
rect 363 2122 415 2126
rect 419 2122 439 2126
rect 443 2122 479 2126
rect 483 2122 519 2126
rect 523 2122 543 2126
rect 547 2122 599 2126
rect 603 2122 607 2126
rect 611 2122 671 2126
rect 675 2122 679 2126
rect 683 2122 735 2126
rect 739 2122 759 2126
rect 763 2122 791 2126
rect 795 2122 831 2126
rect 835 2122 839 2126
rect 843 2122 887 2126
rect 891 2122 903 2126
rect 907 2122 935 2126
rect 939 2122 975 2126
rect 979 2122 991 2126
rect 995 2122 1047 2126
rect 1051 2122 1119 2126
rect 1123 2122 1239 2126
rect 1243 2122 1251 2126
rect 91 2121 1251 2122
rect 1257 2121 1258 2127
rect 1262 2065 1263 2071
rect 1269 2070 2447 2071
rect 1269 2066 1279 2070
rect 1283 2066 1399 2070
rect 1403 2066 1439 2070
rect 1443 2066 1495 2070
rect 1499 2066 1567 2070
rect 1571 2066 1647 2070
rect 1651 2066 1735 2070
rect 1739 2066 1823 2070
rect 1827 2066 1911 2070
rect 1915 2066 1999 2070
rect 2003 2066 2039 2070
rect 2043 2066 2079 2070
rect 2083 2066 2087 2070
rect 2091 2066 2119 2070
rect 2123 2066 2159 2070
rect 2163 2066 2175 2070
rect 2179 2066 2199 2070
rect 2203 2066 2239 2070
rect 2243 2066 2271 2070
rect 2275 2066 2279 2070
rect 2283 2066 2319 2070
rect 2323 2066 2359 2070
rect 2363 2066 2407 2070
rect 2411 2066 2447 2070
rect 1269 2065 2447 2066
rect 2453 2065 2454 2071
rect 96 2049 97 2055
rect 103 2054 1263 2055
rect 103 2050 111 2054
rect 115 2050 135 2054
rect 139 2050 175 2054
rect 179 2050 191 2054
rect 195 2050 215 2054
rect 219 2050 271 2054
rect 275 2050 279 2054
rect 283 2050 343 2054
rect 347 2050 351 2054
rect 355 2050 415 2054
rect 419 2050 423 2054
rect 427 2050 479 2054
rect 483 2050 487 2054
rect 491 2050 543 2054
rect 547 2050 551 2054
rect 555 2050 607 2054
rect 611 2050 615 2054
rect 619 2050 671 2054
rect 675 2050 679 2054
rect 683 2050 735 2054
rect 739 2050 743 2054
rect 747 2050 791 2054
rect 795 2050 815 2054
rect 819 2050 839 2054
rect 843 2050 887 2054
rect 891 2050 935 2054
rect 939 2050 991 2054
rect 995 2050 1047 2054
rect 1051 2050 1239 2054
rect 1243 2050 1263 2054
rect 103 2049 1263 2050
rect 1269 2049 1270 2055
rect 1250 1997 1251 2003
rect 1257 2002 2435 2003
rect 1257 1998 1279 2002
rect 1283 1998 1399 2002
rect 1403 1998 1439 2002
rect 1443 1998 1479 2002
rect 1483 1998 1519 2002
rect 1523 1998 1559 2002
rect 1563 1998 1599 2002
rect 1603 1998 1639 2002
rect 1643 1998 1679 2002
rect 1683 1998 1719 2002
rect 1723 1998 1767 2002
rect 1771 1998 1823 2002
rect 1827 1998 1871 2002
rect 1875 1998 1919 2002
rect 1923 1998 1967 2002
rect 1971 1998 2015 2002
rect 2019 1998 2039 2002
rect 2043 1998 2055 2002
rect 2059 1998 2079 2002
rect 2083 1998 2095 2002
rect 2099 1998 2119 2002
rect 2123 1998 2143 2002
rect 2147 1998 2159 2002
rect 2163 1998 2191 2002
rect 2195 1998 2199 2002
rect 2203 1998 2239 2002
rect 2243 1998 2279 2002
rect 2283 1998 2319 2002
rect 2323 1998 2359 2002
rect 2363 1998 2407 2002
rect 2411 1998 2435 2002
rect 1257 1997 2435 1998
rect 2441 1997 2442 2003
rect 84 1981 85 1987
rect 91 1986 1251 1987
rect 91 1982 111 1986
rect 115 1982 135 1986
rect 139 1982 175 1986
rect 179 1982 215 1986
rect 219 1982 271 1986
rect 275 1982 279 1986
rect 283 1982 343 1986
rect 347 1982 351 1986
rect 355 1982 415 1986
rect 419 1982 423 1986
rect 427 1982 487 1986
rect 491 1982 495 1986
rect 499 1982 551 1986
rect 555 1982 575 1986
rect 579 1982 615 1986
rect 619 1982 647 1986
rect 651 1982 679 1986
rect 683 1982 719 1986
rect 723 1982 743 1986
rect 747 1982 791 1986
rect 795 1982 815 1986
rect 819 1982 863 1986
rect 867 1982 935 1986
rect 939 1982 1007 1986
rect 1011 1982 1239 1986
rect 1243 1982 1251 1986
rect 91 1981 1251 1982
rect 1257 1981 1258 1987
rect 1262 1925 1263 1931
rect 1269 1930 2447 1931
rect 1269 1926 1279 1930
rect 1283 1926 1343 1930
rect 1347 1926 1383 1930
rect 1387 1926 1399 1930
rect 1403 1926 1423 1930
rect 1427 1926 1439 1930
rect 1443 1926 1463 1930
rect 1467 1926 1479 1930
rect 1483 1926 1511 1930
rect 1515 1926 1519 1930
rect 1523 1926 1559 1930
rect 1563 1926 1567 1930
rect 1571 1926 1599 1930
rect 1603 1926 1631 1930
rect 1635 1926 1639 1930
rect 1643 1926 1679 1930
rect 1683 1926 1711 1930
rect 1715 1926 1719 1930
rect 1723 1926 1767 1930
rect 1771 1926 1807 1930
rect 1811 1926 1823 1930
rect 1827 1926 1871 1930
rect 1875 1926 1919 1930
rect 1923 1926 1967 1930
rect 1971 1926 2015 1930
rect 2019 1926 2031 1930
rect 2035 1926 2055 1930
rect 2059 1926 2095 1930
rect 2099 1926 2143 1930
rect 2147 1926 2151 1930
rect 2155 1926 2191 1930
rect 2195 1926 2239 1930
rect 2243 1926 2279 1930
rect 2283 1926 2319 1930
rect 2323 1926 2359 1930
rect 2363 1926 2407 1930
rect 2411 1926 2447 1930
rect 1269 1925 2447 1926
rect 2453 1925 2454 1931
rect 96 1909 97 1915
rect 103 1914 1263 1915
rect 103 1910 111 1914
rect 115 1910 135 1914
rect 139 1910 175 1914
rect 179 1910 215 1914
rect 219 1910 247 1914
rect 251 1910 271 1914
rect 275 1910 287 1914
rect 291 1910 327 1914
rect 331 1910 343 1914
rect 347 1910 367 1914
rect 371 1910 415 1914
rect 419 1910 471 1914
rect 475 1910 495 1914
rect 499 1910 535 1914
rect 539 1910 575 1914
rect 579 1910 599 1914
rect 603 1910 647 1914
rect 651 1910 663 1914
rect 667 1910 719 1914
rect 723 1910 727 1914
rect 731 1910 791 1914
rect 795 1910 855 1914
rect 859 1910 863 1914
rect 867 1910 919 1914
rect 923 1910 935 1914
rect 939 1910 983 1914
rect 987 1910 1007 1914
rect 1011 1910 1055 1914
rect 1059 1910 1127 1914
rect 1131 1910 1239 1914
rect 1243 1910 1263 1914
rect 103 1909 1263 1910
rect 1269 1909 1270 1915
rect 1250 1849 1251 1855
rect 1257 1854 2435 1855
rect 1257 1850 1279 1854
rect 1283 1850 1343 1854
rect 1347 1850 1359 1854
rect 1363 1850 1383 1854
rect 1387 1850 1399 1854
rect 1403 1850 1423 1854
rect 1427 1850 1447 1854
rect 1451 1850 1463 1854
rect 1467 1850 1503 1854
rect 1507 1850 1511 1854
rect 1515 1850 1559 1854
rect 1563 1850 1567 1854
rect 1571 1850 1615 1854
rect 1619 1850 1631 1854
rect 1635 1850 1671 1854
rect 1675 1850 1711 1854
rect 1715 1850 1727 1854
rect 1731 1850 1783 1854
rect 1787 1850 1807 1854
rect 1811 1850 1839 1854
rect 1843 1850 1895 1854
rect 1899 1850 1919 1854
rect 1923 1850 1951 1854
rect 1955 1850 2031 1854
rect 2035 1850 2151 1854
rect 2155 1850 2407 1854
rect 2411 1850 2435 1854
rect 1257 1849 2435 1850
rect 2441 1849 2442 1855
rect 84 1837 85 1843
rect 91 1842 1251 1843
rect 91 1838 111 1842
rect 115 1838 247 1842
rect 251 1838 287 1842
rect 291 1838 327 1842
rect 331 1838 367 1842
rect 371 1838 399 1842
rect 403 1838 415 1842
rect 419 1838 439 1842
rect 443 1838 471 1842
rect 475 1838 479 1842
rect 483 1838 519 1842
rect 523 1838 535 1842
rect 539 1838 567 1842
rect 571 1838 599 1842
rect 603 1838 623 1842
rect 627 1838 663 1842
rect 667 1838 687 1842
rect 691 1838 727 1842
rect 731 1838 759 1842
rect 763 1838 791 1842
rect 795 1838 831 1842
rect 835 1838 855 1842
rect 859 1838 903 1842
rect 907 1838 919 1842
rect 923 1838 975 1842
rect 979 1838 983 1842
rect 987 1838 1047 1842
rect 1051 1838 1055 1842
rect 1059 1838 1127 1842
rect 1131 1838 1191 1842
rect 1195 1838 1239 1842
rect 1243 1838 1251 1842
rect 91 1837 1251 1838
rect 1257 1837 1258 1843
rect 96 1769 97 1775
rect 103 1774 1263 1775
rect 103 1770 111 1774
rect 115 1770 399 1774
rect 403 1770 407 1774
rect 411 1770 439 1774
rect 443 1770 447 1774
rect 451 1770 479 1774
rect 483 1770 487 1774
rect 491 1770 519 1774
rect 523 1770 527 1774
rect 531 1770 567 1774
rect 571 1770 607 1774
rect 611 1770 623 1774
rect 627 1770 647 1774
rect 651 1770 687 1774
rect 691 1770 695 1774
rect 699 1770 751 1774
rect 755 1770 759 1774
rect 763 1770 807 1774
rect 811 1770 831 1774
rect 835 1770 871 1774
rect 875 1770 903 1774
rect 907 1770 935 1774
rect 939 1770 975 1774
rect 979 1770 999 1774
rect 1003 1770 1047 1774
rect 1051 1770 1071 1774
rect 1075 1770 1127 1774
rect 1131 1770 1143 1774
rect 1147 1770 1191 1774
rect 1195 1770 1239 1774
rect 1243 1770 1263 1774
rect 103 1769 1263 1770
rect 1269 1774 2454 1775
rect 1269 1770 1279 1774
rect 1283 1770 1303 1774
rect 1307 1770 1343 1774
rect 1347 1770 1359 1774
rect 1363 1770 1391 1774
rect 1395 1770 1399 1774
rect 1403 1770 1447 1774
rect 1451 1770 1455 1774
rect 1459 1770 1503 1774
rect 1507 1770 1519 1774
rect 1523 1770 1559 1774
rect 1563 1770 1583 1774
rect 1587 1770 1615 1774
rect 1619 1770 1647 1774
rect 1651 1770 1671 1774
rect 1675 1770 1703 1774
rect 1707 1770 1727 1774
rect 1731 1770 1759 1774
rect 1763 1770 1783 1774
rect 1787 1770 1807 1774
rect 1811 1770 1839 1774
rect 1843 1770 1863 1774
rect 1867 1770 1895 1774
rect 1899 1770 1919 1774
rect 1923 1770 1951 1774
rect 1955 1770 1975 1774
rect 1979 1770 2407 1774
rect 2411 1770 2454 1774
rect 1269 1769 2454 1770
rect 84 1697 85 1703
rect 91 1702 1251 1703
rect 91 1698 111 1702
rect 115 1698 279 1702
rect 283 1698 319 1702
rect 323 1698 359 1702
rect 363 1698 399 1702
rect 403 1698 407 1702
rect 411 1698 447 1702
rect 451 1698 487 1702
rect 491 1698 495 1702
rect 499 1698 527 1702
rect 531 1698 543 1702
rect 547 1698 567 1702
rect 571 1698 591 1702
rect 595 1698 607 1702
rect 611 1698 639 1702
rect 643 1698 647 1702
rect 651 1698 687 1702
rect 691 1698 695 1702
rect 699 1698 735 1702
rect 739 1698 751 1702
rect 755 1698 783 1702
rect 787 1698 807 1702
rect 811 1698 839 1702
rect 843 1698 871 1702
rect 875 1698 895 1702
rect 899 1698 935 1702
rect 939 1698 999 1702
rect 1003 1698 1071 1702
rect 1075 1698 1143 1702
rect 1147 1698 1191 1702
rect 1195 1698 1239 1702
rect 1243 1698 1251 1702
rect 91 1697 1251 1698
rect 1257 1702 2442 1703
rect 1257 1698 1279 1702
rect 1283 1698 1303 1702
rect 1307 1698 1343 1702
rect 1347 1698 1383 1702
rect 1387 1698 1391 1702
rect 1395 1698 1423 1702
rect 1427 1698 1455 1702
rect 1459 1698 1463 1702
rect 1467 1698 1503 1702
rect 1507 1698 1519 1702
rect 1523 1698 1559 1702
rect 1563 1698 1583 1702
rect 1587 1698 1623 1702
rect 1627 1698 1647 1702
rect 1651 1698 1687 1702
rect 1691 1698 1703 1702
rect 1707 1698 1751 1702
rect 1755 1698 1759 1702
rect 1763 1698 1807 1702
rect 1811 1698 1863 1702
rect 1867 1698 1919 1702
rect 1923 1698 1975 1702
rect 1979 1698 2031 1702
rect 2035 1698 2087 1702
rect 2091 1698 2407 1702
rect 2411 1698 2442 1702
rect 1257 1697 2442 1698
rect 96 1625 97 1631
rect 103 1630 1263 1631
rect 103 1626 111 1630
rect 115 1626 135 1630
rect 139 1626 175 1630
rect 179 1626 215 1630
rect 219 1626 255 1630
rect 259 1626 279 1630
rect 283 1626 311 1630
rect 315 1626 319 1630
rect 323 1626 359 1630
rect 363 1626 391 1630
rect 395 1626 399 1630
rect 403 1626 447 1630
rect 451 1626 471 1630
rect 475 1626 495 1630
rect 499 1626 543 1630
rect 547 1626 559 1630
rect 563 1626 591 1630
rect 595 1626 639 1630
rect 643 1626 687 1630
rect 691 1626 719 1630
rect 723 1626 735 1630
rect 739 1626 783 1630
rect 787 1626 791 1630
rect 795 1626 839 1630
rect 843 1626 855 1630
rect 859 1626 895 1630
rect 899 1626 919 1630
rect 923 1626 983 1630
rect 987 1626 1047 1630
rect 1051 1626 1239 1630
rect 1243 1626 1263 1630
rect 103 1625 1263 1626
rect 1269 1630 2454 1631
rect 1269 1626 1279 1630
rect 1283 1626 1303 1630
rect 1307 1626 1343 1630
rect 1347 1626 1383 1630
rect 1387 1626 1423 1630
rect 1427 1626 1463 1630
rect 1467 1626 1503 1630
rect 1507 1626 1559 1630
rect 1563 1626 1623 1630
rect 1627 1626 1631 1630
rect 1635 1626 1687 1630
rect 1691 1626 1703 1630
rect 1707 1626 1751 1630
rect 1755 1626 1783 1630
rect 1787 1626 1807 1630
rect 1811 1626 1855 1630
rect 1859 1626 1863 1630
rect 1867 1626 1919 1630
rect 1923 1626 1927 1630
rect 1931 1626 1975 1630
rect 1979 1626 1999 1630
rect 2003 1626 2031 1630
rect 2035 1626 2063 1630
rect 2067 1626 2087 1630
rect 2091 1626 2127 1630
rect 2131 1626 2191 1630
rect 2195 1626 2255 1630
rect 2259 1626 2319 1630
rect 2323 1626 2359 1630
rect 2363 1626 2407 1630
rect 2411 1626 2454 1630
rect 1269 1625 2454 1626
rect 1250 1562 2442 1563
rect 1250 1559 1279 1562
rect 84 1553 85 1559
rect 91 1558 1251 1559
rect 91 1554 111 1558
rect 115 1554 135 1558
rect 139 1554 151 1558
rect 155 1554 175 1558
rect 179 1554 199 1558
rect 203 1554 215 1558
rect 219 1554 255 1558
rect 259 1554 263 1558
rect 267 1554 311 1558
rect 315 1554 343 1558
rect 347 1554 391 1558
rect 395 1554 439 1558
rect 443 1554 471 1558
rect 475 1554 535 1558
rect 539 1554 559 1558
rect 563 1554 639 1558
rect 643 1554 719 1558
rect 723 1554 735 1558
rect 739 1554 791 1558
rect 795 1554 823 1558
rect 827 1554 855 1558
rect 859 1554 903 1558
rect 907 1554 919 1558
rect 923 1554 975 1558
rect 979 1554 983 1558
rect 987 1554 1047 1558
rect 1051 1554 1119 1558
rect 1123 1554 1191 1558
rect 1195 1554 1239 1558
rect 1243 1554 1251 1558
rect 91 1553 1251 1554
rect 1257 1558 1279 1559
rect 1283 1558 1303 1562
rect 1307 1558 1343 1562
rect 1347 1558 1383 1562
rect 1387 1558 1423 1562
rect 1427 1558 1463 1562
rect 1467 1558 1471 1562
rect 1475 1558 1503 1562
rect 1507 1558 1559 1562
rect 1563 1558 1623 1562
rect 1627 1558 1631 1562
rect 1635 1558 1703 1562
rect 1707 1558 1759 1562
rect 1763 1558 1783 1562
rect 1787 1558 1855 1562
rect 1859 1558 1871 1562
rect 1875 1558 1927 1562
rect 1931 1558 1967 1562
rect 1971 1558 1999 1562
rect 2003 1558 2055 1562
rect 2059 1558 2063 1562
rect 2067 1558 2127 1562
rect 2131 1558 2191 1562
rect 2195 1558 2255 1562
rect 2259 1558 2319 1562
rect 2323 1558 2359 1562
rect 2363 1558 2407 1562
rect 2411 1558 2442 1562
rect 1257 1557 2442 1558
rect 1257 1553 1258 1557
rect 96 1481 97 1487
rect 103 1486 1263 1487
rect 103 1482 111 1486
rect 115 1482 151 1486
rect 155 1482 199 1486
rect 203 1482 263 1486
rect 267 1482 319 1486
rect 323 1482 343 1486
rect 347 1482 359 1486
rect 363 1482 399 1486
rect 403 1482 439 1486
rect 443 1482 447 1486
rect 451 1482 503 1486
rect 507 1482 535 1486
rect 539 1482 559 1486
rect 563 1482 615 1486
rect 619 1482 639 1486
rect 643 1482 671 1486
rect 675 1482 735 1486
rect 739 1482 799 1486
rect 803 1482 823 1486
rect 827 1482 855 1486
rect 859 1482 903 1486
rect 907 1482 911 1486
rect 915 1482 967 1486
rect 971 1482 975 1486
rect 979 1482 1023 1486
rect 1027 1482 1047 1486
rect 1051 1482 1087 1486
rect 1091 1482 1119 1486
rect 1123 1482 1151 1486
rect 1155 1482 1191 1486
rect 1195 1482 1239 1486
rect 1243 1482 1263 1486
rect 103 1481 1263 1482
rect 1269 1481 1270 1487
rect 1262 1469 1263 1475
rect 1269 1474 2447 1475
rect 1269 1470 1279 1474
rect 1283 1470 1303 1474
rect 1307 1470 1375 1474
rect 1379 1470 1471 1474
rect 1475 1470 1479 1474
rect 1483 1470 1583 1474
rect 1587 1470 1623 1474
rect 1627 1470 1687 1474
rect 1691 1470 1759 1474
rect 1763 1470 1783 1474
rect 1787 1470 1871 1474
rect 1875 1470 1951 1474
rect 1955 1470 1967 1474
rect 1971 1470 2031 1474
rect 2035 1470 2055 1474
rect 2059 1470 2103 1474
rect 2107 1470 2127 1474
rect 2131 1470 2167 1474
rect 2171 1470 2191 1474
rect 2195 1470 2239 1474
rect 2243 1470 2255 1474
rect 2259 1470 2311 1474
rect 2315 1470 2319 1474
rect 2323 1470 2359 1474
rect 2363 1470 2407 1474
rect 2411 1470 2447 1474
rect 1269 1469 2447 1470
rect 2453 1469 2454 1475
rect 84 1409 85 1415
rect 91 1414 1251 1415
rect 91 1410 111 1414
rect 115 1410 263 1414
rect 267 1410 303 1414
rect 307 1410 319 1414
rect 323 1410 343 1414
rect 347 1410 359 1414
rect 363 1410 391 1414
rect 395 1410 399 1414
rect 403 1410 447 1414
rect 451 1410 503 1414
rect 507 1410 559 1414
rect 563 1410 615 1414
rect 619 1410 623 1414
rect 627 1410 671 1414
rect 675 1410 687 1414
rect 691 1410 735 1414
rect 739 1410 751 1414
rect 755 1410 799 1414
rect 803 1410 815 1414
rect 819 1410 855 1414
rect 859 1410 879 1414
rect 883 1410 911 1414
rect 915 1410 951 1414
rect 955 1410 967 1414
rect 971 1410 1023 1414
rect 1027 1410 1087 1414
rect 1091 1410 1151 1414
rect 1155 1410 1191 1414
rect 1195 1410 1239 1414
rect 1243 1410 1251 1414
rect 91 1409 1251 1410
rect 1257 1409 1258 1415
rect 1250 1407 1258 1409
rect 1250 1401 1251 1407
rect 1257 1406 2435 1407
rect 1257 1402 1279 1406
rect 1283 1402 1303 1406
rect 1307 1402 1343 1406
rect 1347 1402 1375 1406
rect 1379 1402 1399 1406
rect 1403 1402 1471 1406
rect 1475 1402 1479 1406
rect 1483 1402 1551 1406
rect 1555 1402 1583 1406
rect 1587 1402 1639 1406
rect 1643 1402 1687 1406
rect 1691 1402 1727 1406
rect 1731 1402 1783 1406
rect 1787 1402 1815 1406
rect 1819 1402 1871 1406
rect 1875 1402 1903 1406
rect 1907 1402 1951 1406
rect 1955 1402 1991 1406
rect 1995 1402 2031 1406
rect 2035 1402 2071 1406
rect 2075 1402 2103 1406
rect 2107 1402 2151 1406
rect 2155 1402 2167 1406
rect 2171 1402 2223 1406
rect 2227 1402 2239 1406
rect 2243 1402 2303 1406
rect 2307 1402 2311 1406
rect 2315 1402 2359 1406
rect 2363 1402 2407 1406
rect 2411 1402 2435 1406
rect 1257 1401 2435 1402
rect 2441 1401 2442 1407
rect 96 1337 97 1343
rect 103 1342 1263 1343
rect 103 1338 111 1342
rect 115 1338 135 1342
rect 139 1338 175 1342
rect 179 1338 215 1342
rect 219 1338 255 1342
rect 259 1338 263 1342
rect 267 1338 303 1342
rect 307 1338 327 1342
rect 331 1338 343 1342
rect 347 1338 391 1342
rect 395 1338 407 1342
rect 411 1338 447 1342
rect 451 1338 495 1342
rect 499 1338 503 1342
rect 507 1338 559 1342
rect 563 1338 583 1342
rect 587 1338 623 1342
rect 627 1338 671 1342
rect 675 1338 687 1342
rect 691 1338 751 1342
rect 755 1338 759 1342
rect 763 1338 815 1342
rect 819 1338 839 1342
rect 843 1338 879 1342
rect 883 1338 919 1342
rect 923 1338 951 1342
rect 955 1338 1007 1342
rect 1011 1338 1023 1342
rect 1027 1338 1095 1342
rect 1099 1338 1239 1342
rect 1243 1338 1263 1342
rect 103 1337 1263 1338
rect 1269 1337 1270 1343
rect 1262 1335 1270 1337
rect 1262 1329 1263 1335
rect 1269 1334 2447 1335
rect 1269 1330 1279 1334
rect 1283 1330 1303 1334
rect 1307 1330 1343 1334
rect 1347 1330 1399 1334
rect 1403 1330 1447 1334
rect 1451 1330 1471 1334
rect 1475 1330 1487 1334
rect 1491 1330 1527 1334
rect 1531 1330 1551 1334
rect 1555 1330 1567 1334
rect 1571 1330 1615 1334
rect 1619 1330 1639 1334
rect 1643 1330 1671 1334
rect 1675 1330 1719 1334
rect 1723 1330 1727 1334
rect 1731 1330 1775 1334
rect 1779 1330 1815 1334
rect 1819 1330 1831 1334
rect 1835 1330 1903 1334
rect 1907 1330 1983 1334
rect 1987 1330 1991 1334
rect 1995 1330 2071 1334
rect 2075 1330 2151 1334
rect 2155 1330 2167 1334
rect 2171 1330 2223 1334
rect 2227 1330 2271 1334
rect 2275 1330 2303 1334
rect 2307 1330 2359 1334
rect 2363 1330 2407 1334
rect 2411 1330 2447 1334
rect 1269 1329 2447 1330
rect 2453 1329 2454 1335
rect 84 1265 85 1271
rect 91 1270 1251 1271
rect 91 1266 111 1270
rect 115 1266 135 1270
rect 139 1266 175 1270
rect 179 1266 215 1270
rect 219 1266 247 1270
rect 251 1266 255 1270
rect 259 1266 327 1270
rect 331 1266 407 1270
rect 411 1266 415 1270
rect 419 1266 495 1270
rect 499 1266 503 1270
rect 507 1266 583 1270
rect 587 1266 591 1270
rect 595 1266 671 1270
rect 675 1266 743 1270
rect 747 1266 759 1270
rect 763 1266 815 1270
rect 819 1266 839 1270
rect 843 1266 879 1270
rect 883 1266 919 1270
rect 923 1266 943 1270
rect 947 1266 1007 1270
rect 1011 1266 1071 1270
rect 1075 1266 1095 1270
rect 1099 1266 1239 1270
rect 1243 1266 1251 1270
rect 91 1265 1251 1266
rect 1257 1265 1258 1271
rect 1250 1263 1258 1265
rect 1250 1257 1251 1263
rect 1257 1262 2435 1263
rect 1257 1258 1279 1262
rect 1283 1258 1447 1262
rect 1451 1258 1487 1262
rect 1491 1258 1511 1262
rect 1515 1258 1527 1262
rect 1531 1258 1551 1262
rect 1555 1258 1567 1262
rect 1571 1258 1591 1262
rect 1595 1258 1615 1262
rect 1619 1258 1631 1262
rect 1635 1258 1671 1262
rect 1675 1258 1711 1262
rect 1715 1258 1719 1262
rect 1723 1258 1751 1262
rect 1755 1258 1775 1262
rect 1779 1258 1791 1262
rect 1795 1258 1831 1262
rect 1835 1258 1839 1262
rect 1843 1258 1903 1262
rect 1907 1258 1967 1262
rect 1971 1258 1983 1262
rect 1987 1258 2039 1262
rect 2043 1258 2071 1262
rect 2075 1258 2119 1262
rect 2123 1258 2167 1262
rect 2171 1258 2207 1262
rect 2211 1258 2271 1262
rect 2275 1258 2295 1262
rect 2299 1258 2359 1262
rect 2363 1258 2407 1262
rect 2411 1258 2435 1262
rect 1257 1257 2435 1258
rect 2441 1257 2442 1263
rect 96 1189 97 1195
rect 103 1194 1263 1195
rect 103 1190 111 1194
rect 115 1190 135 1194
rect 139 1190 175 1194
rect 179 1190 231 1194
rect 235 1190 247 1194
rect 251 1190 303 1194
rect 307 1190 327 1194
rect 331 1190 383 1194
rect 387 1190 415 1194
rect 419 1190 471 1194
rect 475 1190 503 1194
rect 507 1190 559 1194
rect 563 1190 591 1194
rect 595 1190 639 1194
rect 643 1190 671 1194
rect 675 1190 719 1194
rect 723 1190 743 1194
rect 747 1190 799 1194
rect 803 1190 815 1194
rect 819 1190 871 1194
rect 875 1190 879 1194
rect 883 1190 935 1194
rect 939 1190 943 1194
rect 947 1190 991 1194
rect 995 1190 1007 1194
rect 1011 1190 1047 1194
rect 1051 1190 1071 1194
rect 1075 1190 1103 1194
rect 1107 1190 1151 1194
rect 1155 1190 1191 1194
rect 1195 1190 1239 1194
rect 1243 1190 1263 1194
rect 103 1189 1263 1190
rect 1269 1191 1270 1195
rect 1269 1190 2454 1191
rect 1269 1189 1279 1190
rect 1262 1186 1279 1189
rect 1283 1186 1511 1190
rect 1515 1186 1551 1190
rect 1555 1186 1559 1190
rect 1563 1186 1591 1190
rect 1595 1186 1599 1190
rect 1603 1186 1631 1190
rect 1635 1186 1639 1190
rect 1643 1186 1671 1190
rect 1675 1186 1679 1190
rect 1683 1186 1711 1190
rect 1715 1186 1719 1190
rect 1723 1186 1751 1190
rect 1755 1186 1759 1190
rect 1763 1186 1791 1190
rect 1795 1186 1799 1190
rect 1803 1186 1839 1190
rect 1843 1186 1855 1190
rect 1859 1186 1903 1190
rect 1907 1186 1927 1190
rect 1931 1186 1967 1190
rect 1971 1186 2023 1190
rect 2027 1186 2039 1190
rect 2043 1186 2119 1190
rect 2123 1186 2135 1190
rect 2139 1186 2207 1190
rect 2211 1186 2255 1190
rect 2259 1186 2295 1190
rect 2299 1186 2359 1190
rect 2363 1186 2407 1190
rect 2411 1186 2454 1190
rect 1262 1185 2454 1186
rect 84 1121 85 1127
rect 91 1126 1251 1127
rect 91 1122 111 1126
rect 115 1122 135 1126
rect 139 1122 175 1126
rect 179 1122 215 1126
rect 219 1122 231 1126
rect 235 1122 303 1126
rect 307 1122 383 1126
rect 387 1122 391 1126
rect 395 1122 471 1126
rect 475 1122 479 1126
rect 483 1122 559 1126
rect 563 1122 639 1126
rect 643 1122 711 1126
rect 715 1122 719 1126
rect 723 1122 775 1126
rect 779 1122 799 1126
rect 803 1122 839 1126
rect 843 1122 871 1126
rect 875 1122 903 1126
rect 907 1122 935 1126
rect 939 1122 959 1126
rect 963 1122 991 1126
rect 995 1122 1023 1126
rect 1027 1122 1047 1126
rect 1051 1122 1087 1126
rect 1091 1122 1103 1126
rect 1107 1122 1151 1126
rect 1155 1122 1191 1126
rect 1195 1122 1239 1126
rect 1243 1122 1251 1126
rect 91 1121 1251 1122
rect 1257 1121 1258 1127
rect 1250 1109 1251 1115
rect 1257 1114 2435 1115
rect 1257 1110 1279 1114
rect 1283 1110 1535 1114
rect 1539 1110 1559 1114
rect 1563 1110 1599 1114
rect 1603 1110 1639 1114
rect 1643 1110 1663 1114
rect 1667 1110 1679 1114
rect 1683 1110 1719 1114
rect 1723 1110 1727 1114
rect 1731 1110 1759 1114
rect 1763 1110 1791 1114
rect 1795 1110 1799 1114
rect 1803 1110 1855 1114
rect 1859 1110 1911 1114
rect 1915 1110 1927 1114
rect 1931 1110 1967 1114
rect 1971 1110 2023 1114
rect 2027 1110 2079 1114
rect 2083 1110 2135 1114
rect 2139 1110 2191 1114
rect 2195 1110 2255 1114
rect 2259 1110 2319 1114
rect 2323 1110 2359 1114
rect 2363 1110 2407 1114
rect 2411 1110 2435 1114
rect 1257 1109 2435 1110
rect 2441 1109 2442 1115
rect 96 1049 97 1055
rect 103 1054 1263 1055
rect 103 1050 111 1054
rect 115 1050 135 1054
rect 139 1050 199 1054
rect 203 1050 215 1054
rect 219 1050 239 1054
rect 243 1050 287 1054
rect 291 1050 303 1054
rect 307 1050 343 1054
rect 347 1050 391 1054
rect 395 1050 439 1054
rect 443 1050 479 1054
rect 483 1050 487 1054
rect 491 1050 535 1054
rect 539 1050 559 1054
rect 563 1050 583 1054
rect 587 1050 631 1054
rect 635 1050 639 1054
rect 643 1050 679 1054
rect 683 1050 711 1054
rect 715 1050 727 1054
rect 731 1050 775 1054
rect 779 1050 783 1054
rect 787 1050 839 1054
rect 843 1050 895 1054
rect 899 1050 903 1054
rect 907 1050 959 1054
rect 963 1050 1023 1054
rect 1027 1050 1087 1054
rect 1091 1050 1151 1054
rect 1155 1050 1191 1054
rect 1195 1050 1239 1054
rect 1243 1050 1263 1054
rect 103 1049 1263 1050
rect 1269 1049 1270 1055
rect 1262 1029 1263 1035
rect 1269 1034 2447 1035
rect 1269 1030 1279 1034
rect 1283 1030 1503 1034
rect 1507 1030 1535 1034
rect 1539 1030 1599 1034
rect 1603 1030 1623 1034
rect 1627 1030 1663 1034
rect 1667 1030 1727 1034
rect 1731 1030 1735 1034
rect 1739 1030 1791 1034
rect 1795 1030 1831 1034
rect 1835 1030 1855 1034
rect 1859 1030 1911 1034
rect 1915 1030 1919 1034
rect 1923 1030 1967 1034
rect 1971 1030 1999 1034
rect 2003 1030 2023 1034
rect 2027 1030 2071 1034
rect 2075 1030 2079 1034
rect 2083 1030 2135 1034
rect 2139 1030 2143 1034
rect 2147 1030 2191 1034
rect 2195 1030 2207 1034
rect 2211 1030 2255 1034
rect 2259 1030 2279 1034
rect 2283 1030 2319 1034
rect 2323 1030 2359 1034
rect 2363 1030 2407 1034
rect 2411 1030 2447 1034
rect 1269 1029 2447 1030
rect 2453 1029 2454 1035
rect 84 969 85 975
rect 91 974 1251 975
rect 91 970 111 974
rect 115 970 199 974
rect 203 970 239 974
rect 243 970 287 974
rect 291 970 295 974
rect 299 970 343 974
rect 347 970 391 974
rect 395 970 399 974
rect 403 970 439 974
rect 443 970 471 974
rect 475 970 487 974
rect 491 970 535 974
rect 539 970 551 974
rect 555 970 583 974
rect 587 970 631 974
rect 635 970 639 974
rect 643 970 679 974
rect 683 970 727 974
rect 731 970 783 974
rect 787 970 807 974
rect 811 970 839 974
rect 843 970 887 974
rect 891 970 895 974
rect 899 970 959 974
rect 963 970 1023 974
rect 1027 970 1087 974
rect 1091 970 1151 974
rect 1155 970 1191 974
rect 1195 970 1239 974
rect 1243 970 1251 974
rect 91 969 1251 970
rect 1257 969 1258 975
rect 1250 953 1251 959
rect 1257 958 2435 959
rect 1257 954 1279 958
rect 1283 954 1319 958
rect 1323 954 1359 958
rect 1363 954 1399 958
rect 1403 954 1463 958
rect 1467 954 1503 958
rect 1507 954 1543 958
rect 1547 954 1623 958
rect 1627 954 1639 958
rect 1643 954 1735 958
rect 1739 954 1831 958
rect 1835 954 1839 958
rect 1843 954 1919 958
rect 1923 954 1935 958
rect 1939 954 1999 958
rect 2003 954 2023 958
rect 2027 954 2071 958
rect 2075 954 2103 958
rect 2107 954 2143 958
rect 2147 954 2175 958
rect 2179 954 2207 958
rect 2211 954 2239 958
rect 2243 954 2279 958
rect 2283 954 2311 958
rect 2315 954 2359 958
rect 2363 954 2407 958
rect 2411 954 2435 958
rect 1257 953 2435 954
rect 2441 953 2442 959
rect 96 893 97 899
rect 103 898 1263 899
rect 103 894 111 898
rect 115 894 255 898
rect 259 894 295 898
rect 299 894 311 898
rect 315 894 343 898
rect 347 894 375 898
rect 379 894 399 898
rect 403 894 455 898
rect 459 894 471 898
rect 475 894 535 898
rect 539 894 551 898
rect 555 894 623 898
rect 627 894 639 898
rect 643 894 711 898
rect 715 894 727 898
rect 731 894 791 898
rect 795 894 807 898
rect 811 894 863 898
rect 867 894 887 898
rect 891 894 935 898
rect 939 894 959 898
rect 963 894 999 898
rect 1003 894 1023 898
rect 1027 894 1055 898
rect 1059 894 1087 898
rect 1091 894 1119 898
rect 1123 894 1151 898
rect 1155 894 1183 898
rect 1187 894 1191 898
rect 1195 894 1239 898
rect 1243 894 1263 898
rect 103 893 1263 894
rect 1269 893 1270 899
rect 1262 877 1263 883
rect 1269 882 2447 883
rect 1269 878 1279 882
rect 1283 878 1319 882
rect 1323 878 1335 882
rect 1339 878 1359 882
rect 1363 878 1375 882
rect 1379 878 1399 882
rect 1403 878 1415 882
rect 1419 878 1463 882
rect 1467 878 1471 882
rect 1475 878 1535 882
rect 1539 878 1543 882
rect 1547 878 1607 882
rect 1611 878 1639 882
rect 1643 878 1679 882
rect 1683 878 1735 882
rect 1739 878 1751 882
rect 1755 878 1823 882
rect 1827 878 1839 882
rect 1843 878 1895 882
rect 1899 878 1935 882
rect 1939 878 1959 882
rect 1963 878 2023 882
rect 2027 878 2087 882
rect 2091 878 2103 882
rect 2107 878 2143 882
rect 2147 878 2175 882
rect 2179 878 2199 882
rect 2203 878 2239 882
rect 2243 878 2255 882
rect 2259 878 2311 882
rect 2315 878 2319 882
rect 2323 878 2359 882
rect 2363 878 2407 882
rect 2411 878 2447 882
rect 1269 877 2447 878
rect 2453 877 2454 883
rect 84 825 85 831
rect 91 830 1251 831
rect 91 826 111 830
rect 115 826 191 830
rect 195 826 247 830
rect 251 826 255 830
rect 259 826 311 830
rect 315 826 375 830
rect 379 826 383 830
rect 387 826 455 830
rect 459 826 463 830
rect 467 826 535 830
rect 539 826 543 830
rect 547 826 615 830
rect 619 826 623 830
rect 627 826 687 830
rect 691 826 711 830
rect 715 826 751 830
rect 755 826 791 830
rect 795 826 815 830
rect 819 826 863 830
rect 867 826 871 830
rect 875 826 927 830
rect 931 826 935 830
rect 939 826 983 830
rect 987 826 999 830
rect 1003 826 1047 830
rect 1051 826 1055 830
rect 1059 826 1119 830
rect 1123 826 1183 830
rect 1187 826 1239 830
rect 1243 826 1251 830
rect 91 825 1251 826
rect 1257 825 1258 831
rect 1250 805 1251 811
rect 1257 810 2435 811
rect 1257 806 1279 810
rect 1283 806 1303 810
rect 1307 806 1335 810
rect 1339 806 1343 810
rect 1347 806 1375 810
rect 1379 806 1407 810
rect 1411 806 1415 810
rect 1419 806 1471 810
rect 1475 806 1479 810
rect 1483 806 1535 810
rect 1539 806 1551 810
rect 1555 806 1607 810
rect 1611 806 1623 810
rect 1627 806 1679 810
rect 1683 806 1695 810
rect 1699 806 1751 810
rect 1755 806 1759 810
rect 1763 806 1823 810
rect 1827 806 1887 810
rect 1891 806 1895 810
rect 1899 806 1951 810
rect 1955 806 1959 810
rect 1963 806 2023 810
rect 2027 806 2087 810
rect 2091 806 2103 810
rect 2107 806 2143 810
rect 2147 806 2191 810
rect 2195 806 2199 810
rect 2203 806 2255 810
rect 2259 806 2279 810
rect 2283 806 2319 810
rect 2323 806 2359 810
rect 2363 806 2407 810
rect 2411 806 2435 810
rect 1257 805 2435 806
rect 2441 805 2442 811
rect 96 757 97 763
rect 103 762 1263 763
rect 103 758 111 762
rect 115 758 135 762
rect 139 758 175 762
rect 179 758 191 762
rect 195 758 215 762
rect 219 758 247 762
rect 251 758 279 762
rect 283 758 311 762
rect 315 758 351 762
rect 355 758 383 762
rect 387 758 423 762
rect 427 758 463 762
rect 467 758 495 762
rect 499 758 543 762
rect 547 758 559 762
rect 563 758 615 762
rect 619 758 623 762
rect 627 758 687 762
rect 691 758 695 762
rect 699 758 751 762
rect 755 758 783 762
rect 787 758 815 762
rect 819 758 871 762
rect 875 758 879 762
rect 883 758 927 762
rect 931 758 983 762
rect 987 758 1047 762
rect 1051 758 1095 762
rect 1099 758 1191 762
rect 1195 758 1239 762
rect 1243 758 1263 762
rect 103 757 1263 758
rect 1269 757 1270 763
rect 1262 737 1263 743
rect 1269 742 2447 743
rect 1269 738 1279 742
rect 1283 738 1303 742
rect 1307 738 1343 742
rect 1347 738 1367 742
rect 1371 738 1407 742
rect 1411 738 1455 742
rect 1459 738 1479 742
rect 1483 738 1535 742
rect 1539 738 1551 742
rect 1555 738 1615 742
rect 1619 738 1623 742
rect 1627 738 1695 742
rect 1699 738 1759 742
rect 1763 738 1775 742
rect 1779 738 1823 742
rect 1827 738 1855 742
rect 1859 738 1887 742
rect 1891 738 1943 742
rect 1947 738 1951 742
rect 1955 738 2023 742
rect 2027 738 2031 742
rect 2035 738 2103 742
rect 2107 738 2119 742
rect 2123 738 2191 742
rect 2195 738 2207 742
rect 2211 738 2279 742
rect 2283 738 2295 742
rect 2299 738 2359 742
rect 2363 738 2407 742
rect 2411 738 2447 742
rect 1269 737 2447 738
rect 2453 737 2454 743
rect 84 681 85 687
rect 91 686 1251 687
rect 91 682 111 686
rect 115 682 135 686
rect 139 682 175 686
rect 179 682 215 686
rect 219 682 231 686
rect 235 682 279 686
rect 283 682 287 686
rect 291 682 343 686
rect 347 682 351 686
rect 355 682 399 686
rect 403 682 423 686
rect 427 682 455 686
rect 459 682 495 686
rect 499 682 503 686
rect 507 682 559 686
rect 563 682 623 686
rect 627 682 695 686
rect 699 682 767 686
rect 771 682 783 686
rect 787 682 839 686
rect 843 682 879 686
rect 883 682 903 686
rect 907 682 967 686
rect 971 682 983 686
rect 987 682 1023 686
rect 1027 682 1087 686
rect 1091 682 1095 686
rect 1099 682 1151 686
rect 1155 682 1191 686
rect 1195 682 1239 686
rect 1243 682 1251 686
rect 91 681 1251 682
rect 1257 681 1258 687
rect 1250 669 1251 675
rect 1257 674 2435 675
rect 1257 670 1279 674
rect 1283 670 1303 674
rect 1307 670 1367 674
rect 1371 670 1455 674
rect 1459 670 1535 674
rect 1539 670 1591 674
rect 1595 670 1615 674
rect 1619 670 1639 674
rect 1643 670 1687 674
rect 1691 670 1695 674
rect 1699 670 1743 674
rect 1747 670 1775 674
rect 1779 670 1799 674
rect 1803 670 1855 674
rect 1859 670 1871 674
rect 1875 670 1943 674
rect 1947 670 1951 674
rect 1955 670 2031 674
rect 2035 670 2047 674
rect 2051 670 2119 674
rect 2123 670 2151 674
rect 2155 670 2207 674
rect 2211 670 2263 674
rect 2267 670 2295 674
rect 2299 670 2359 674
rect 2363 670 2407 674
rect 2411 670 2435 674
rect 1257 669 2435 670
rect 2441 669 2442 675
rect 96 613 97 619
rect 103 618 1263 619
rect 103 614 111 618
rect 115 614 135 618
rect 139 614 175 618
rect 179 614 183 618
rect 187 614 231 618
rect 235 614 255 618
rect 259 614 287 618
rect 291 614 327 618
rect 331 614 343 618
rect 347 614 399 618
rect 403 614 455 618
rect 459 614 479 618
rect 483 614 503 618
rect 507 614 559 618
rect 563 614 623 618
rect 627 614 639 618
rect 643 614 695 618
rect 699 614 719 618
rect 723 614 767 618
rect 771 614 799 618
rect 803 614 839 618
rect 843 614 879 618
rect 883 614 903 618
rect 907 614 951 618
rect 955 614 967 618
rect 971 614 1015 618
rect 1019 614 1023 618
rect 1027 614 1079 618
rect 1083 614 1087 618
rect 1091 614 1143 618
rect 1147 614 1151 618
rect 1155 614 1191 618
rect 1195 614 1239 618
rect 1243 614 1263 618
rect 103 613 1263 614
rect 1269 613 1270 619
rect 1262 593 1263 599
rect 1269 598 2447 599
rect 1269 594 1279 598
rect 1283 594 1559 598
rect 1563 594 1591 598
rect 1595 594 1599 598
rect 1603 594 1639 598
rect 1643 594 1679 598
rect 1683 594 1687 598
rect 1691 594 1719 598
rect 1723 594 1743 598
rect 1747 594 1759 598
rect 1763 594 1799 598
rect 1803 594 1807 598
rect 1811 594 1855 598
rect 1859 594 1871 598
rect 1875 594 1911 598
rect 1915 594 1951 598
rect 1955 594 1967 598
rect 1971 594 2031 598
rect 2035 594 2047 598
rect 2051 594 2095 598
rect 2099 594 2151 598
rect 2155 594 2167 598
rect 2171 594 2239 598
rect 2243 594 2263 598
rect 2267 594 2311 598
rect 2315 594 2359 598
rect 2363 594 2407 598
rect 2411 594 2447 598
rect 1269 593 2447 594
rect 2453 593 2454 599
rect 84 541 85 547
rect 91 546 1251 547
rect 91 542 111 546
rect 115 542 135 546
rect 139 542 151 546
rect 155 542 183 546
rect 187 542 223 546
rect 227 542 255 546
rect 259 542 287 546
rect 291 542 327 546
rect 331 542 351 546
rect 355 542 399 546
rect 403 542 415 546
rect 419 542 479 546
rect 483 542 551 546
rect 555 542 559 546
rect 563 542 623 546
rect 627 542 639 546
rect 643 542 695 546
rect 699 542 719 546
rect 723 542 767 546
rect 771 542 799 546
rect 803 542 839 546
rect 843 542 879 546
rect 883 542 919 546
rect 923 542 951 546
rect 955 542 999 546
rect 1003 542 1015 546
rect 1019 542 1079 546
rect 1083 542 1143 546
rect 1147 542 1191 546
rect 1195 542 1239 546
rect 1243 542 1251 546
rect 91 541 1251 542
rect 1257 541 1258 547
rect 1250 525 1251 531
rect 1257 530 2435 531
rect 1257 526 1279 530
rect 1283 526 1407 530
rect 1411 526 1447 530
rect 1451 526 1487 530
rect 1491 526 1535 530
rect 1539 526 1559 530
rect 1563 526 1591 530
rect 1595 526 1599 530
rect 1603 526 1639 530
rect 1643 526 1647 530
rect 1651 526 1679 530
rect 1683 526 1711 530
rect 1715 526 1719 530
rect 1723 526 1759 530
rect 1763 526 1783 530
rect 1787 526 1807 530
rect 1811 526 1855 530
rect 1859 526 1863 530
rect 1867 526 1911 530
rect 1915 526 1943 530
rect 1947 526 1967 530
rect 1971 526 2023 530
rect 2027 526 2031 530
rect 2035 526 2095 530
rect 2099 526 2103 530
rect 2107 526 2167 530
rect 2171 526 2191 530
rect 2195 526 2239 530
rect 2243 526 2287 530
rect 2291 526 2311 530
rect 2315 526 2359 530
rect 2363 526 2407 530
rect 2411 526 2435 530
rect 1257 525 2435 526
rect 2441 525 2442 531
rect 96 473 97 479
rect 103 478 1263 479
rect 103 474 111 478
rect 115 474 151 478
rect 155 474 223 478
rect 227 474 239 478
rect 243 474 279 478
rect 283 474 287 478
rect 291 474 327 478
rect 331 474 351 478
rect 355 474 383 478
rect 387 474 415 478
rect 419 474 439 478
rect 443 474 479 478
rect 483 474 503 478
rect 507 474 551 478
rect 555 474 567 478
rect 571 474 623 478
rect 627 474 631 478
rect 635 474 695 478
rect 699 474 759 478
rect 763 474 767 478
rect 771 474 823 478
rect 827 474 839 478
rect 843 474 887 478
rect 891 474 919 478
rect 923 474 951 478
rect 955 474 999 478
rect 1003 474 1015 478
rect 1019 474 1079 478
rect 1083 474 1239 478
rect 1243 474 1263 478
rect 103 473 1263 474
rect 1269 473 1270 479
rect 1262 457 1263 463
rect 1269 462 2447 463
rect 1269 458 1279 462
rect 1283 458 1303 462
rect 1307 458 1343 462
rect 1347 458 1383 462
rect 1387 458 1407 462
rect 1411 458 1447 462
rect 1451 458 1487 462
rect 1491 458 1535 462
rect 1539 458 1591 462
rect 1595 458 1631 462
rect 1635 458 1647 462
rect 1651 458 1711 462
rect 1715 458 1735 462
rect 1739 458 1783 462
rect 1787 458 1831 462
rect 1835 458 1863 462
rect 1867 458 1919 462
rect 1923 458 1943 462
rect 1947 458 1999 462
rect 2003 458 2023 462
rect 2027 458 2071 462
rect 2075 458 2103 462
rect 2107 458 2135 462
rect 2139 458 2191 462
rect 2195 458 2199 462
rect 2203 458 2255 462
rect 2259 458 2287 462
rect 2291 458 2319 462
rect 2323 458 2359 462
rect 2363 458 2407 462
rect 2411 458 2447 462
rect 1269 457 2447 458
rect 2453 457 2454 463
rect 84 401 85 407
rect 91 406 1251 407
rect 91 402 111 406
rect 115 402 143 406
rect 147 402 183 406
rect 187 402 223 406
rect 227 402 239 406
rect 243 402 271 406
rect 275 402 279 406
rect 283 402 327 406
rect 331 402 335 406
rect 339 402 383 406
rect 387 402 399 406
rect 403 402 439 406
rect 443 402 471 406
rect 475 402 503 406
rect 507 402 543 406
rect 547 402 567 406
rect 571 402 615 406
rect 619 402 631 406
rect 635 402 687 406
rect 691 402 695 406
rect 699 402 751 406
rect 755 402 759 406
rect 763 402 807 406
rect 811 402 823 406
rect 827 402 863 406
rect 867 402 887 406
rect 891 402 919 406
rect 923 402 951 406
rect 955 402 975 406
rect 979 402 1015 406
rect 1019 402 1031 406
rect 1035 402 1239 406
rect 1243 402 1251 406
rect 91 401 1251 402
rect 1257 401 1258 407
rect 1250 389 1251 395
rect 1257 394 2435 395
rect 1257 390 1279 394
rect 1283 390 1303 394
rect 1307 390 1343 394
rect 1347 390 1359 394
rect 1363 390 1383 394
rect 1387 390 1399 394
rect 1403 390 1439 394
rect 1443 390 1447 394
rect 1451 390 1487 394
rect 1491 390 1535 394
rect 1539 390 1543 394
rect 1547 390 1607 394
rect 1611 390 1631 394
rect 1635 390 1679 394
rect 1683 390 1735 394
rect 1739 390 1759 394
rect 1763 390 1831 394
rect 1835 390 1839 394
rect 1843 390 1919 394
rect 1923 390 1999 394
rect 2003 390 2071 394
rect 2075 390 2079 394
rect 2083 390 2135 394
rect 2139 390 2159 394
rect 2163 390 2199 394
rect 2203 390 2247 394
rect 2251 390 2255 394
rect 2259 390 2319 394
rect 2323 390 2335 394
rect 2339 390 2359 394
rect 2363 390 2407 394
rect 2411 390 2435 394
rect 1257 389 2435 390
rect 2441 389 2442 395
rect 96 325 97 331
rect 103 330 1263 331
rect 103 326 111 330
rect 115 326 135 330
rect 139 326 143 330
rect 147 326 175 330
rect 179 326 183 330
rect 187 326 215 330
rect 219 326 223 330
rect 227 326 255 330
rect 259 326 271 330
rect 275 326 295 330
rect 299 326 335 330
rect 339 326 391 330
rect 395 326 399 330
rect 403 326 447 330
rect 451 326 471 330
rect 475 326 495 330
rect 499 326 543 330
rect 547 326 591 330
rect 595 326 615 330
rect 619 326 639 330
rect 643 326 687 330
rect 691 326 735 330
rect 739 326 751 330
rect 755 326 783 330
rect 787 326 807 330
rect 811 326 839 330
rect 843 326 863 330
rect 867 326 919 330
rect 923 326 975 330
rect 979 326 1031 330
rect 1035 326 1239 330
rect 1243 326 1263 330
rect 103 325 1263 326
rect 1269 325 1270 331
rect 1262 313 1263 319
rect 1269 318 2447 319
rect 1269 314 1279 318
rect 1283 314 1359 318
rect 1363 314 1399 318
rect 1403 314 1439 318
rect 1443 314 1487 318
rect 1491 314 1511 318
rect 1515 314 1543 318
rect 1547 314 1551 318
rect 1555 314 1591 318
rect 1595 314 1607 318
rect 1611 314 1631 318
rect 1635 314 1671 318
rect 1675 314 1679 318
rect 1683 314 1711 318
rect 1715 314 1751 318
rect 1755 314 1759 318
rect 1763 314 1791 318
rect 1795 314 1839 318
rect 1843 314 1903 318
rect 1907 314 1919 318
rect 1923 314 1967 318
rect 1971 314 1999 318
rect 2003 314 2039 318
rect 2043 314 2079 318
rect 2083 314 2119 318
rect 2123 314 2159 318
rect 2163 314 2199 318
rect 2203 314 2247 318
rect 2251 314 2279 318
rect 2283 314 2335 318
rect 2339 314 2359 318
rect 2363 314 2407 318
rect 2411 314 2447 318
rect 1269 313 2447 314
rect 2453 313 2454 319
rect 84 249 85 255
rect 91 254 1251 255
rect 91 250 111 254
rect 115 250 135 254
rect 139 250 175 254
rect 179 250 215 254
rect 219 250 223 254
rect 227 250 255 254
rect 259 250 295 254
rect 299 250 311 254
rect 315 250 335 254
rect 339 250 391 254
rect 395 250 447 254
rect 451 250 463 254
rect 467 250 495 254
rect 499 250 527 254
rect 531 250 543 254
rect 547 250 591 254
rect 595 250 639 254
rect 643 250 647 254
rect 651 250 687 254
rect 691 250 695 254
rect 699 250 735 254
rect 739 250 783 254
rect 787 250 831 254
rect 835 250 839 254
rect 843 250 879 254
rect 883 250 927 254
rect 931 250 975 254
rect 979 250 1023 254
rect 1027 250 1239 254
rect 1243 250 1251 254
rect 91 249 1251 250
rect 1257 249 1258 255
rect 1250 247 1258 249
rect 1250 241 1251 247
rect 1257 246 2435 247
rect 1257 242 1279 246
rect 1283 242 1367 246
rect 1371 242 1407 246
rect 1411 242 1455 246
rect 1459 242 1511 246
rect 1515 242 1551 246
rect 1555 242 1567 246
rect 1571 242 1591 246
rect 1595 242 1631 246
rect 1635 242 1671 246
rect 1675 242 1703 246
rect 1707 242 1711 246
rect 1715 242 1751 246
rect 1755 242 1775 246
rect 1779 242 1791 246
rect 1795 242 1839 246
rect 1843 242 1855 246
rect 1859 242 1903 246
rect 1907 242 1943 246
rect 1947 242 1967 246
rect 1971 242 2031 246
rect 2035 242 2039 246
rect 2043 242 2119 246
rect 2123 242 2199 246
rect 2203 242 2207 246
rect 2211 242 2279 246
rect 2283 242 2295 246
rect 2299 242 2359 246
rect 2363 242 2407 246
rect 2411 242 2435 246
rect 1257 241 2435 242
rect 2441 241 2442 247
rect 1262 165 1263 171
rect 1269 170 2447 171
rect 1269 166 1279 170
rect 1283 166 1303 170
rect 1307 166 1343 170
rect 1347 166 1367 170
rect 1371 166 1383 170
rect 1387 166 1407 170
rect 1411 166 1423 170
rect 1427 166 1455 170
rect 1459 166 1463 170
rect 1467 166 1511 170
rect 1515 166 1519 170
rect 1523 166 1567 170
rect 1571 166 1583 170
rect 1587 166 1631 170
rect 1635 166 1647 170
rect 1651 166 1703 170
rect 1707 166 1711 170
rect 1715 166 1775 170
rect 1779 166 1831 170
rect 1835 166 1855 170
rect 1859 166 1887 170
rect 1891 166 1935 170
rect 1939 166 1943 170
rect 1947 166 1975 170
rect 1979 166 2015 170
rect 2019 166 2031 170
rect 2035 166 2055 170
rect 2059 166 2095 170
rect 2099 166 2119 170
rect 2123 166 2143 170
rect 2147 166 2191 170
rect 2195 166 2207 170
rect 2211 166 2239 170
rect 2243 166 2279 170
rect 2283 166 2295 170
rect 2299 166 2319 170
rect 2323 166 2359 170
rect 2363 166 2407 170
rect 2411 166 2447 170
rect 1269 165 2447 166
rect 2453 165 2454 171
rect 96 149 97 155
rect 103 154 1263 155
rect 103 150 111 154
rect 115 150 135 154
rect 139 150 151 154
rect 155 150 191 154
rect 195 150 223 154
rect 227 150 231 154
rect 235 150 271 154
rect 275 150 311 154
rect 315 150 351 154
rect 355 150 391 154
rect 395 150 431 154
rect 435 150 463 154
rect 467 150 471 154
rect 475 150 511 154
rect 515 150 527 154
rect 531 150 551 154
rect 555 150 591 154
rect 595 150 631 154
rect 635 150 647 154
rect 651 150 671 154
rect 675 150 695 154
rect 699 150 711 154
rect 715 150 735 154
rect 739 150 751 154
rect 755 150 783 154
rect 787 150 791 154
rect 795 150 831 154
rect 835 150 871 154
rect 875 150 879 154
rect 883 150 911 154
rect 915 150 927 154
rect 931 150 951 154
rect 955 150 975 154
rect 979 150 991 154
rect 995 150 1023 154
rect 1027 150 1031 154
rect 1035 150 1071 154
rect 1075 150 1111 154
rect 1115 150 1151 154
rect 1155 150 1191 154
rect 1195 150 1239 154
rect 1243 150 1263 154
rect 103 149 1263 150
rect 1269 149 1270 155
rect 1250 97 1251 103
rect 1257 102 2435 103
rect 1257 98 1279 102
rect 1283 98 1303 102
rect 1307 98 1343 102
rect 1347 98 1383 102
rect 1387 98 1423 102
rect 1427 98 1463 102
rect 1467 98 1519 102
rect 1523 98 1583 102
rect 1587 98 1647 102
rect 1651 98 1711 102
rect 1715 98 1775 102
rect 1779 98 1831 102
rect 1835 98 1887 102
rect 1891 98 1935 102
rect 1939 98 1975 102
rect 1979 98 2015 102
rect 2019 98 2055 102
rect 2059 98 2095 102
rect 2099 98 2143 102
rect 2147 98 2191 102
rect 2195 98 2239 102
rect 2243 98 2279 102
rect 2283 98 2319 102
rect 2323 98 2359 102
rect 2363 98 2407 102
rect 2411 98 2435 102
rect 1257 97 2435 98
rect 2441 97 2442 103
rect 84 81 85 87
rect 91 86 1251 87
rect 91 82 111 86
rect 115 82 151 86
rect 155 82 191 86
rect 195 82 231 86
rect 235 82 271 86
rect 275 82 311 86
rect 315 82 351 86
rect 355 82 391 86
rect 395 82 431 86
rect 435 82 471 86
rect 475 82 511 86
rect 515 82 551 86
rect 555 82 591 86
rect 595 82 631 86
rect 635 82 671 86
rect 675 82 711 86
rect 715 82 751 86
rect 755 82 791 86
rect 795 82 831 86
rect 835 82 871 86
rect 875 82 911 86
rect 915 82 951 86
rect 955 82 991 86
rect 995 82 1031 86
rect 1035 82 1071 86
rect 1075 82 1111 86
rect 1115 82 1151 86
rect 1155 82 1191 86
rect 1195 82 1239 86
rect 1243 82 1251 86
rect 91 81 1251 82
rect 1257 81 1258 87
<< m5c >>
rect 97 2489 103 2495
rect 1263 2489 1269 2495
rect 85 2413 91 2419
rect 1251 2413 1257 2419
rect 97 2341 103 2347
rect 1263 2341 1269 2347
rect 1251 2277 1257 2283
rect 2435 2277 2441 2283
rect 85 2265 91 2271
rect 1251 2265 1257 2271
rect 97 2197 103 2203
rect 1263 2197 1269 2203
rect 1251 2133 1257 2139
rect 2435 2133 2441 2139
rect 85 2121 91 2127
rect 1251 2121 1257 2127
rect 1263 2065 1269 2071
rect 2447 2065 2453 2071
rect 97 2049 103 2055
rect 1263 2049 1269 2055
rect 1251 1997 1257 2003
rect 2435 1997 2441 2003
rect 85 1981 91 1987
rect 1251 1981 1257 1987
rect 1263 1925 1269 1931
rect 2447 1925 2453 1931
rect 97 1909 103 1915
rect 1263 1909 1269 1915
rect 1251 1849 1257 1855
rect 2435 1849 2441 1855
rect 85 1837 91 1843
rect 1251 1837 1257 1843
rect 97 1769 103 1775
rect 1263 1769 1269 1775
rect 85 1697 91 1703
rect 1251 1697 1257 1703
rect 97 1625 103 1631
rect 1263 1625 1269 1631
rect 85 1553 91 1559
rect 1251 1553 1257 1559
rect 97 1481 103 1487
rect 1263 1481 1269 1487
rect 1263 1469 1269 1475
rect 2447 1469 2453 1475
rect 85 1409 91 1415
rect 1251 1409 1257 1415
rect 1251 1401 1257 1407
rect 2435 1401 2441 1407
rect 97 1337 103 1343
rect 1263 1337 1269 1343
rect 1263 1329 1269 1335
rect 2447 1329 2453 1335
rect 85 1265 91 1271
rect 1251 1265 1257 1271
rect 1251 1257 1257 1263
rect 2435 1257 2441 1263
rect 97 1189 103 1195
rect 1263 1189 1269 1195
rect 85 1121 91 1127
rect 1251 1121 1257 1127
rect 1251 1109 1257 1115
rect 2435 1109 2441 1115
rect 97 1049 103 1055
rect 1263 1049 1269 1055
rect 1263 1029 1269 1035
rect 2447 1029 2453 1035
rect 85 969 91 975
rect 1251 969 1257 975
rect 1251 953 1257 959
rect 2435 953 2441 959
rect 97 893 103 899
rect 1263 893 1269 899
rect 1263 877 1269 883
rect 2447 877 2453 883
rect 85 825 91 831
rect 1251 825 1257 831
rect 1251 805 1257 811
rect 2435 805 2441 811
rect 97 757 103 763
rect 1263 757 1269 763
rect 1263 737 1269 743
rect 2447 737 2453 743
rect 85 681 91 687
rect 1251 681 1257 687
rect 1251 669 1257 675
rect 2435 669 2441 675
rect 97 613 103 619
rect 1263 613 1269 619
rect 1263 593 1269 599
rect 2447 593 2453 599
rect 85 541 91 547
rect 1251 541 1257 547
rect 1251 525 1257 531
rect 2435 525 2441 531
rect 97 473 103 479
rect 1263 473 1269 479
rect 1263 457 1269 463
rect 2447 457 2453 463
rect 85 401 91 407
rect 1251 401 1257 407
rect 1251 389 1257 395
rect 2435 389 2441 395
rect 97 325 103 331
rect 1263 325 1269 331
rect 1263 313 1269 319
rect 2447 313 2453 319
rect 85 249 91 255
rect 1251 249 1257 255
rect 1251 241 1257 247
rect 2435 241 2441 247
rect 1263 165 1269 171
rect 2447 165 2453 171
rect 97 149 103 155
rect 1263 149 1269 155
rect 1251 97 1257 103
rect 2435 97 2441 103
rect 85 81 91 87
rect 1251 81 1257 87
<< m5 >>
rect 84 2419 92 2520
rect 84 2413 85 2419
rect 91 2413 92 2419
rect 84 2271 92 2413
rect 84 2265 85 2271
rect 91 2265 92 2271
rect 84 2127 92 2265
rect 84 2121 85 2127
rect 91 2121 92 2127
rect 84 1987 92 2121
rect 84 1981 85 1987
rect 91 1981 92 1987
rect 84 1843 92 1981
rect 84 1837 85 1843
rect 91 1837 92 1843
rect 84 1703 92 1837
rect 84 1697 85 1703
rect 91 1697 92 1703
rect 84 1559 92 1697
rect 84 1553 85 1559
rect 91 1553 92 1559
rect 84 1415 92 1553
rect 84 1409 85 1415
rect 91 1409 92 1415
rect 84 1271 92 1409
rect 84 1265 85 1271
rect 91 1265 92 1271
rect 84 1127 92 1265
rect 84 1121 85 1127
rect 91 1121 92 1127
rect 84 975 92 1121
rect 84 969 85 975
rect 91 969 92 975
rect 84 831 92 969
rect 84 825 85 831
rect 91 825 92 831
rect 84 687 92 825
rect 84 681 85 687
rect 91 681 92 687
rect 84 547 92 681
rect 84 541 85 547
rect 91 541 92 547
rect 84 407 92 541
rect 84 401 85 407
rect 91 401 92 407
rect 84 255 92 401
rect 84 249 85 255
rect 91 249 92 255
rect 84 87 92 249
rect 84 81 85 87
rect 91 81 92 87
rect 84 72 92 81
rect 96 2495 104 2520
rect 96 2489 97 2495
rect 103 2489 104 2495
rect 96 2347 104 2489
rect 96 2341 97 2347
rect 103 2341 104 2347
rect 96 2203 104 2341
rect 96 2197 97 2203
rect 103 2197 104 2203
rect 96 2055 104 2197
rect 96 2049 97 2055
rect 103 2049 104 2055
rect 96 1915 104 2049
rect 96 1909 97 1915
rect 103 1909 104 1915
rect 96 1775 104 1909
rect 96 1769 97 1775
rect 103 1769 104 1775
rect 96 1631 104 1769
rect 96 1625 97 1631
rect 103 1625 104 1631
rect 96 1487 104 1625
rect 96 1481 97 1487
rect 103 1481 104 1487
rect 96 1343 104 1481
rect 96 1337 97 1343
rect 103 1337 104 1343
rect 96 1195 104 1337
rect 96 1189 97 1195
rect 103 1189 104 1195
rect 96 1055 104 1189
rect 96 1049 97 1055
rect 103 1049 104 1055
rect 96 899 104 1049
rect 96 893 97 899
rect 103 893 104 899
rect 96 763 104 893
rect 96 757 97 763
rect 103 757 104 763
rect 96 619 104 757
rect 96 613 97 619
rect 103 613 104 619
rect 96 479 104 613
rect 96 473 97 479
rect 103 473 104 479
rect 96 331 104 473
rect 96 325 97 331
rect 103 325 104 331
rect 96 155 104 325
rect 96 149 97 155
rect 103 149 104 155
rect 96 72 104 149
rect 1250 2419 1258 2520
rect 1250 2413 1251 2419
rect 1257 2413 1258 2419
rect 1250 2283 1258 2413
rect 1250 2277 1251 2283
rect 1257 2277 1258 2283
rect 1250 2271 1258 2277
rect 1250 2265 1251 2271
rect 1257 2265 1258 2271
rect 1250 2139 1258 2265
rect 1250 2133 1251 2139
rect 1257 2133 1258 2139
rect 1250 2127 1258 2133
rect 1250 2121 1251 2127
rect 1257 2121 1258 2127
rect 1250 2003 1258 2121
rect 1250 1997 1251 2003
rect 1257 1997 1258 2003
rect 1250 1987 1258 1997
rect 1250 1981 1251 1987
rect 1257 1981 1258 1987
rect 1250 1855 1258 1981
rect 1250 1849 1251 1855
rect 1257 1849 1258 1855
rect 1250 1843 1258 1849
rect 1250 1837 1251 1843
rect 1257 1837 1258 1843
rect 1250 1703 1258 1837
rect 1250 1697 1251 1703
rect 1257 1697 1258 1703
rect 1250 1559 1258 1697
rect 1250 1553 1251 1559
rect 1257 1553 1258 1559
rect 1250 1415 1258 1553
rect 1250 1409 1251 1415
rect 1257 1409 1258 1415
rect 1250 1407 1258 1409
rect 1250 1401 1251 1407
rect 1257 1401 1258 1407
rect 1250 1271 1258 1401
rect 1250 1265 1251 1271
rect 1257 1265 1258 1271
rect 1250 1263 1258 1265
rect 1250 1257 1251 1263
rect 1257 1257 1258 1263
rect 1250 1127 1258 1257
rect 1250 1121 1251 1127
rect 1257 1121 1258 1127
rect 1250 1115 1258 1121
rect 1250 1109 1251 1115
rect 1257 1109 1258 1115
rect 1250 975 1258 1109
rect 1250 969 1251 975
rect 1257 969 1258 975
rect 1250 959 1258 969
rect 1250 953 1251 959
rect 1257 953 1258 959
rect 1250 831 1258 953
rect 1250 825 1251 831
rect 1257 825 1258 831
rect 1250 811 1258 825
rect 1250 805 1251 811
rect 1257 805 1258 811
rect 1250 687 1258 805
rect 1250 681 1251 687
rect 1257 681 1258 687
rect 1250 675 1258 681
rect 1250 669 1251 675
rect 1257 669 1258 675
rect 1250 547 1258 669
rect 1250 541 1251 547
rect 1257 541 1258 547
rect 1250 531 1258 541
rect 1250 525 1251 531
rect 1257 525 1258 531
rect 1250 407 1258 525
rect 1250 401 1251 407
rect 1257 401 1258 407
rect 1250 395 1258 401
rect 1250 389 1251 395
rect 1257 389 1258 395
rect 1250 255 1258 389
rect 1250 249 1251 255
rect 1257 249 1258 255
rect 1250 247 1258 249
rect 1250 241 1251 247
rect 1257 241 1258 247
rect 1250 103 1258 241
rect 1250 97 1251 103
rect 1257 97 1258 103
rect 1250 87 1258 97
rect 1250 81 1251 87
rect 1257 81 1258 87
rect 1250 72 1258 81
rect 1262 2495 1270 2520
rect 1262 2489 1263 2495
rect 1269 2489 1270 2495
rect 1262 2347 1270 2489
rect 1262 2341 1263 2347
rect 1269 2341 1270 2347
rect 1262 2203 1270 2341
rect 1262 2197 1263 2203
rect 1269 2197 1270 2203
rect 1262 2071 1270 2197
rect 1262 2065 1263 2071
rect 1269 2065 1270 2071
rect 1262 2055 1270 2065
rect 1262 2049 1263 2055
rect 1269 2049 1270 2055
rect 1262 1931 1270 2049
rect 1262 1925 1263 1931
rect 1269 1925 1270 1931
rect 1262 1915 1270 1925
rect 1262 1909 1263 1915
rect 1269 1909 1270 1915
rect 1262 1775 1270 1909
rect 1262 1769 1263 1775
rect 1269 1769 1270 1775
rect 1262 1631 1270 1769
rect 1262 1625 1263 1631
rect 1269 1625 1270 1631
rect 1262 1487 1270 1625
rect 1262 1481 1263 1487
rect 1269 1481 1270 1487
rect 1262 1475 1270 1481
rect 1262 1469 1263 1475
rect 1269 1469 1270 1475
rect 1262 1343 1270 1469
rect 1262 1337 1263 1343
rect 1269 1337 1270 1343
rect 1262 1335 1270 1337
rect 1262 1329 1263 1335
rect 1269 1329 1270 1335
rect 1262 1195 1270 1329
rect 1262 1189 1263 1195
rect 1269 1189 1270 1195
rect 1262 1055 1270 1189
rect 1262 1049 1263 1055
rect 1269 1049 1270 1055
rect 1262 1035 1270 1049
rect 1262 1029 1263 1035
rect 1269 1029 1270 1035
rect 1262 899 1270 1029
rect 1262 893 1263 899
rect 1269 893 1270 899
rect 1262 883 1270 893
rect 1262 877 1263 883
rect 1269 877 1270 883
rect 1262 763 1270 877
rect 1262 757 1263 763
rect 1269 757 1270 763
rect 1262 743 1270 757
rect 1262 737 1263 743
rect 1269 737 1270 743
rect 1262 619 1270 737
rect 1262 613 1263 619
rect 1269 613 1270 619
rect 1262 599 1270 613
rect 1262 593 1263 599
rect 1269 593 1270 599
rect 1262 479 1270 593
rect 1262 473 1263 479
rect 1269 473 1270 479
rect 1262 463 1270 473
rect 1262 457 1263 463
rect 1269 457 1270 463
rect 1262 331 1270 457
rect 1262 325 1263 331
rect 1269 325 1270 331
rect 1262 319 1270 325
rect 1262 313 1263 319
rect 1269 313 1270 319
rect 1262 171 1270 313
rect 1262 165 1263 171
rect 1269 165 1270 171
rect 1262 155 1270 165
rect 1262 149 1263 155
rect 1269 149 1270 155
rect 1262 72 1270 149
rect 2434 2283 2442 2520
rect 2434 2277 2435 2283
rect 2441 2277 2442 2283
rect 2434 2139 2442 2277
rect 2434 2133 2435 2139
rect 2441 2133 2442 2139
rect 2434 2003 2442 2133
rect 2434 1997 2435 2003
rect 2441 1997 2442 2003
rect 2434 1855 2442 1997
rect 2434 1849 2435 1855
rect 2441 1849 2442 1855
rect 2434 1407 2442 1849
rect 2434 1401 2435 1407
rect 2441 1401 2442 1407
rect 2434 1263 2442 1401
rect 2434 1257 2435 1263
rect 2441 1257 2442 1263
rect 2434 1115 2442 1257
rect 2434 1109 2435 1115
rect 2441 1109 2442 1115
rect 2434 959 2442 1109
rect 2434 953 2435 959
rect 2441 953 2442 959
rect 2434 811 2442 953
rect 2434 805 2435 811
rect 2441 805 2442 811
rect 2434 675 2442 805
rect 2434 669 2435 675
rect 2441 669 2442 675
rect 2434 531 2442 669
rect 2434 525 2435 531
rect 2441 525 2442 531
rect 2434 395 2442 525
rect 2434 389 2435 395
rect 2441 389 2442 395
rect 2434 247 2442 389
rect 2434 241 2435 247
rect 2441 241 2442 247
rect 2434 103 2442 241
rect 2434 97 2435 103
rect 2441 97 2442 103
rect 2434 72 2442 97
rect 2446 2071 2454 2520
rect 2446 2065 2447 2071
rect 2453 2065 2454 2071
rect 2446 1931 2454 2065
rect 2446 1925 2447 1931
rect 2453 1925 2454 1931
rect 2446 1475 2454 1925
rect 2446 1469 2447 1475
rect 2453 1469 2454 1475
rect 2446 1335 2454 1469
rect 2446 1329 2447 1335
rect 2453 1329 2454 1335
rect 2446 1035 2454 1329
rect 2446 1029 2447 1035
rect 2453 1029 2454 1035
rect 2446 883 2454 1029
rect 2446 877 2447 883
rect 2453 877 2454 883
rect 2446 743 2454 877
rect 2446 737 2447 743
rect 2453 737 2454 743
rect 2446 599 2454 737
rect 2446 593 2447 599
rect 2453 593 2454 599
rect 2446 463 2454 593
rect 2446 457 2447 463
rect 2453 457 2454 463
rect 2446 319 2454 457
rect 2446 313 2447 319
rect 2453 313 2454 319
rect 2446 171 2454 313
rect 2446 165 2447 171
rect 2453 165 2454 171
rect 2446 72 2454 165
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__131
timestamp 1731220637
transform 1 0 2400 0 1 2428
box 7 3 12 24
use welltap_svt  __well_tap__130
timestamp 1731220637
transform 1 0 1272 0 1 2428
box 7 3 12 24
use welltap_svt  __well_tap__129
timestamp 1731220637
transform 1 0 2400 0 -1 2412
box 7 3 12 24
use welltap_svt  __well_tap__128
timestamp 1731220637
transform 1 0 1272 0 -1 2412
box 7 3 12 24
use welltap_svt  __well_tap__127
timestamp 1731220637
transform 1 0 2400 0 1 2288
box 7 3 12 24
use welltap_svt  __well_tap__126
timestamp 1731220637
transform 1 0 1272 0 1 2288
box 7 3 12 24
use welltap_svt  __well_tap__125
timestamp 1731220637
transform 1 0 2400 0 -1 2272
box 7 3 12 24
use welltap_svt  __well_tap__124
timestamp 1731220637
transform 1 0 1272 0 -1 2272
box 7 3 12 24
use welltap_svt  __well_tap__123
timestamp 1731220637
transform 1 0 2400 0 1 2144
box 7 3 12 24
use welltap_svt  __well_tap__122
timestamp 1731220637
transform 1 0 1272 0 1 2144
box 7 3 12 24
use welltap_svt  __well_tap__121
timestamp 1731220637
transform 1 0 2400 0 -1 2128
box 7 3 12 24
use welltap_svt  __well_tap__120
timestamp 1731220637
transform 1 0 1272 0 -1 2128
box 7 3 12 24
use welltap_svt  __well_tap__119
timestamp 1731220637
transform 1 0 2400 0 1 2008
box 7 3 12 24
use welltap_svt  __well_tap__118
timestamp 1731220637
transform 1 0 1272 0 1 2008
box 7 3 12 24
use welltap_svt  __well_tap__117
timestamp 1731220637
transform 1 0 2400 0 -1 1992
box 7 3 12 24
use welltap_svt  __well_tap__116
timestamp 1731220637
transform 1 0 1272 0 -1 1992
box 7 3 12 24
use welltap_svt  __well_tap__115
timestamp 1731220637
transform 1 0 2400 0 1 1868
box 7 3 12 24
use welltap_svt  __well_tap__114
timestamp 1731220637
transform 1 0 1272 0 1 1868
box 7 3 12 24
use welltap_svt  __well_tap__113
timestamp 1731220637
transform 1 0 2400 0 -1 1844
box 7 3 12 24
use welltap_svt  __well_tap__112
timestamp 1731220637
transform 1 0 1272 0 -1 1844
box 7 3 12 24
use welltap_svt  __well_tap__111
timestamp 1731220637
transform 1 0 2400 0 1 1712
box 7 3 12 24
use welltap_svt  __well_tap__110
timestamp 1731220637
transform 1 0 1272 0 1 1712
box 7 3 12 24
use welltap_svt  __well_tap__109
timestamp 1731220637
transform 1 0 2400 0 -1 1692
box 7 3 12 24
use welltap_svt  __well_tap__108
timestamp 1731220637
transform 1 0 1272 0 -1 1692
box 7 3 12 24
use welltap_svt  __well_tap__107
timestamp 1731220637
transform 1 0 2400 0 1 1568
box 7 3 12 24
use welltap_svt  __well_tap__106
timestamp 1731220637
transform 1 0 1272 0 1 1568
box 7 3 12 24
use welltap_svt  __well_tap__105
timestamp 1731220637
transform 1 0 2400 0 -1 1552
box 7 3 12 24
use welltap_svt  __well_tap__104
timestamp 1731220637
transform 1 0 1272 0 -1 1552
box 7 3 12 24
use welltap_svt  __well_tap__103
timestamp 1731220637
transform 1 0 2400 0 1 1412
box 7 3 12 24
use welltap_svt  __well_tap__102
timestamp 1731220637
transform 1 0 1272 0 1 1412
box 7 3 12 24
use welltap_svt  __well_tap__101
timestamp 1731220637
transform 1 0 2400 0 -1 1396
box 7 3 12 24
use welltap_svt  __well_tap__100
timestamp 1731220637
transform 1 0 1272 0 -1 1396
box 7 3 12 24
use welltap_svt  __well_tap__99
timestamp 1731220637
transform 1 0 2400 0 1 1272
box 7 3 12 24
use welltap_svt  __well_tap__98
timestamp 1731220637
transform 1 0 1272 0 1 1272
box 7 3 12 24
use welltap_svt  __well_tap__97
timestamp 1731220637
transform 1 0 2400 0 -1 1252
box 7 3 12 24
use welltap_svt  __well_tap__96
timestamp 1731220637
transform 1 0 1272 0 -1 1252
box 7 3 12 24
use welltap_svt  __well_tap__95
timestamp 1731220637
transform 1 0 2400 0 1 1128
box 7 3 12 24
use welltap_svt  __well_tap__94
timestamp 1731220637
transform 1 0 1272 0 1 1128
box 7 3 12 24
use welltap_svt  __well_tap__93
timestamp 1731220637
transform 1 0 2400 0 -1 1104
box 7 3 12 24
use welltap_svt  __well_tap__92
timestamp 1731220637
transform 1 0 1272 0 -1 1104
box 7 3 12 24
use welltap_svt  __well_tap__91
timestamp 1731220637
transform 1 0 2400 0 1 972
box 7 3 12 24
use welltap_svt  __well_tap__90
timestamp 1731220637
transform 1 0 1272 0 1 972
box 7 3 12 24
use welltap_svt  __well_tap__89
timestamp 1731220637
transform 1 0 2400 0 -1 948
box 7 3 12 24
use welltap_svt  __well_tap__88
timestamp 1731220637
transform 1 0 1272 0 -1 948
box 7 3 12 24
use welltap_svt  __well_tap__87
timestamp 1731220637
transform 1 0 2400 0 1 820
box 7 3 12 24
use welltap_svt  __well_tap__86
timestamp 1731220637
transform 1 0 1272 0 1 820
box 7 3 12 24
use welltap_svt  __well_tap__85
timestamp 1731220637
transform 1 0 2400 0 -1 800
box 7 3 12 24
use welltap_svt  __well_tap__84
timestamp 1731220637
transform 1 0 1272 0 -1 800
box 7 3 12 24
use welltap_svt  __well_tap__83
timestamp 1731220637
transform 1 0 2400 0 1 680
box 7 3 12 24
use welltap_svt  __well_tap__82
timestamp 1731220637
transform 1 0 1272 0 1 680
box 7 3 12 24
use welltap_svt  __well_tap__81
timestamp 1731220637
transform 1 0 2400 0 -1 664
box 7 3 12 24
use welltap_svt  __well_tap__80
timestamp 1731220637
transform 1 0 1272 0 -1 664
box 7 3 12 24
use welltap_svt  __well_tap__79
timestamp 1731220637
transform 1 0 2400 0 1 536
box 7 3 12 24
use welltap_svt  __well_tap__78
timestamp 1731220637
transform 1 0 1272 0 1 536
box 7 3 12 24
use welltap_svt  __well_tap__77
timestamp 1731220637
transform 1 0 2400 0 -1 520
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220637
transform 1 0 1272 0 -1 520
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220637
transform 1 0 2400 0 1 400
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220637
transform 1 0 1272 0 1 400
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220637
transform 1 0 2400 0 -1 384
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220637
transform 1 0 1272 0 -1 384
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220637
transform 1 0 2400 0 1 256
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220637
transform 1 0 1272 0 1 256
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220637
transform 1 0 2400 0 -1 236
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220637
transform 1 0 1272 0 -1 236
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220637
transform 1 0 2400 0 1 108
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220637
transform 1 0 1272 0 1 108
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220637
transform 1 0 1232 0 1 2432
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220637
transform 1 0 104 0 1 2432
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220637
transform 1 0 1232 0 -1 2408
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220637
transform 1 0 104 0 -1 2408
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220637
transform 1 0 1232 0 1 2284
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220637
transform 1 0 104 0 1 2284
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220637
transform 1 0 1232 0 -1 2260
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220637
transform 1 0 104 0 -1 2260
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220637
transform 1 0 1232 0 1 2140
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220637
transform 1 0 104 0 1 2140
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220637
transform 1 0 1232 0 -1 2116
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220637
transform 1 0 104 0 -1 2116
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220637
transform 1 0 1232 0 1 1992
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220637
transform 1 0 104 0 1 1992
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220637
transform 1 0 1232 0 -1 1976
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220637
transform 1 0 104 0 -1 1976
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220637
transform 1 0 1232 0 1 1852
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220637
transform 1 0 104 0 1 1852
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220637
transform 1 0 1232 0 -1 1832
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220637
transform 1 0 104 0 -1 1832
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220637
transform 1 0 1232 0 1 1712
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220637
transform 1 0 104 0 1 1712
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220637
transform 1 0 1232 0 -1 1692
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220637
transform 1 0 104 0 -1 1692
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220637
transform 1 0 1232 0 1 1568
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220637
transform 1 0 104 0 1 1568
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220637
transform 1 0 1232 0 -1 1548
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220637
transform 1 0 104 0 -1 1548
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220637
transform 1 0 1232 0 1 1424
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220637
transform 1 0 104 0 1 1424
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220637
transform 1 0 1232 0 -1 1404
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220637
transform 1 0 104 0 -1 1404
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220637
transform 1 0 1232 0 1 1280
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220637
transform 1 0 104 0 1 1280
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220637
transform 1 0 1232 0 -1 1260
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220637
transform 1 0 104 0 -1 1260
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220637
transform 1 0 1232 0 1 1132
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220637
transform 1 0 104 0 1 1132
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220637
transform 1 0 1232 0 -1 1116
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220637
transform 1 0 104 0 -1 1116
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220637
transform 1 0 1232 0 1 992
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220637
transform 1 0 104 0 1 992
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220637
transform 1 0 1232 0 -1 964
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220637
transform 1 0 104 0 -1 964
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220637
transform 1 0 1232 0 1 836
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220637
transform 1 0 104 0 1 836
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220637
transform 1 0 1232 0 -1 820
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220637
transform 1 0 104 0 -1 820
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220637
transform 1 0 1232 0 1 700
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220637
transform 1 0 104 0 1 700
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220637
transform 1 0 1232 0 -1 676
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220637
transform 1 0 104 0 -1 676
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220637
transform 1 0 1232 0 1 556
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220637
transform 1 0 104 0 1 556
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220637
transform 1 0 1232 0 -1 536
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220637
transform 1 0 104 0 -1 536
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220637
transform 1 0 1232 0 1 416
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220637
transform 1 0 104 0 1 416
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220637
transform 1 0 1232 0 -1 396
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220637
transform 1 0 104 0 -1 396
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220637
transform 1 0 1232 0 1 268
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220637
transform 1 0 104 0 1 268
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220637
transform 1 0 1232 0 -1 244
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220637
transform 1 0 104 0 -1 244
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220637
transform 1 0 1232 0 1 92
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220637
transform 1 0 104 0 1 92
box 7 3 12 24
use _0_0std_0_0cells_0_0NOR2X2  tst_5999_6
timestamp 1731220637
transform 1 0 144 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5998_6
timestamp 1731220637
transform 1 0 184 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5997_6
timestamp 1731220637
transform 1 0 224 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5996_6
timestamp 1731220637
transform 1 0 264 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5995_6
timestamp 1731220637
transform 1 0 304 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5994_6
timestamp 1731220637
transform 1 0 344 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5993_6
timestamp 1731220637
transform 1 0 384 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5992_6
timestamp 1731220637
transform 1 0 424 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5991_6
timestamp 1731220637
transform 1 0 464 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5990_6
timestamp 1731220637
transform 1 0 504 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5989_6
timestamp 1731220637
transform 1 0 544 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5988_6
timestamp 1731220637
transform 1 0 584 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5987_6
timestamp 1731220637
transform 1 0 216 0 -1 252
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5986_6
timestamp 1731220637
transform 1 0 304 0 -1 252
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5985_6
timestamp 1731220637
transform 1 0 384 0 -1 252
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5984_6
timestamp 1731220637
transform 1 0 456 0 -1 252
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5983_6
timestamp 1731220637
transform 1 0 520 0 -1 252
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5982_6
timestamp 1731220637
transform 1 0 584 0 -1 252
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5981_6
timestamp 1731220637
transform 1 0 640 0 -1 252
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5980_6
timestamp 1731220637
transform 1 0 488 0 1 260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5979_6
timestamp 1731220637
transform 1 0 536 0 1 260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5978_6
timestamp 1731220637
transform 1 0 832 0 1 260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5977_6
timestamp 1731220637
transform 1 0 912 0 -1 404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5976_6
timestamp 1731220637
transform 1 0 968 0 -1 404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5975_6
timestamp 1731220637
transform 1 0 1024 0 -1 404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5974_6
timestamp 1731220637
transform 1 0 1008 0 1 408
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5973_6
timestamp 1731220637
transform 1 0 944 0 1 408
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5972_6
timestamp 1731220637
transform 1 0 912 0 -1 544
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5971_6
timestamp 1731220637
transform 1 0 992 0 -1 544
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5970_6
timestamp 1731220637
transform 1 0 1072 0 -1 544
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5969_6
timestamp 1731220637
transform 1 0 1008 0 1 548
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5968_6
timestamp 1731220637
transform 1 0 944 0 1 548
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5967_6
timestamp 1731220637
transform 1 0 872 0 1 548
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5966_6
timestamp 1731220637
transform 1 0 896 0 -1 684
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5965_6
timestamp 1731220637
transform 1 0 960 0 -1 684
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5964_6
timestamp 1731220637
transform 1 0 1016 0 -1 684
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5963_6
timestamp 1731220637
transform 1 0 1072 0 1 548
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5962_6
timestamp 1731220637
transform 1 0 1136 0 1 548
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5961_6
timestamp 1731220637
transform 1 0 1184 0 1 548
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5960_6
timestamp 1731220637
transform 1 0 1184 0 -1 684
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5959_6
timestamp 1731220637
transform 1 0 1080 0 -1 684
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5958_6
timestamp 1731220637
transform 1 0 1144 0 -1 684
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5957_6
timestamp 1731220637
transform 1 0 1184 0 1 692
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5956_6
timestamp 1731220637
transform 1 0 1296 0 1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5955_6
timestamp 1731220637
transform 1 0 1360 0 1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5954_6
timestamp 1731220637
transform 1 0 1400 0 -1 808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5953_6
timestamp 1731220637
transform 1 0 1336 0 -1 808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5952_6
timestamp 1731220637
transform 1 0 1296 0 -1 808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5951_6
timestamp 1731220637
transform 1 0 1328 0 1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5950_6
timestamp 1731220637
transform 1 0 1368 0 1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5949_6
timestamp 1731220637
transform 1 0 1408 0 1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5948_6
timestamp 1731220637
transform 1 0 1312 0 -1 956
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5947_6
timestamp 1731220637
transform 1 0 1352 0 -1 956
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5946_6
timestamp 1731220637
transform 1 0 1392 0 -1 956
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5945_6
timestamp 1731220637
transform 1 0 1536 0 -1 956
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5944_6
timestamp 1731220637
transform 1 0 1632 0 -1 956
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5943_6
timestamp 1731220637
transform 1 0 1728 0 -1 956
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5942_6
timestamp 1731220637
transform 1 0 1832 0 -1 956
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5941_6
timestamp 1731220637
transform 1 0 1744 0 1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5940_6
timestamp 1731220637
transform 1 0 1672 0 1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5939_6
timestamp 1731220637
transform 1 0 1600 0 1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5938_6
timestamp 1731220637
transform 1 0 1616 0 -1 808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5937_6
timestamp 1731220637
transform 1 0 1688 0 -1 808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5936_6
timestamp 1731220637
transform 1 0 1688 0 1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5935_6
timestamp 1731220637
transform 1 0 1608 0 1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5934_6
timestamp 1731220637
transform 1 0 1632 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5933_6
timestamp 1731220637
transform 1 0 1680 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5932_6
timestamp 1731220637
transform 1 0 1736 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5931_6
timestamp 1731220637
transform 1 0 1792 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5930_6
timestamp 1731220637
transform 1 0 1864 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5929_6
timestamp 1731220637
transform 1 0 1848 0 1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5928_6
timestamp 1731220637
transform 1 0 1904 0 1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5927_6
timestamp 1731220637
transform 1 0 1936 0 -1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5926_6
timestamp 1731220637
transform 1 0 1856 0 -1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5925_6
timestamp 1731220637
transform 1 0 1776 0 -1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5924_6
timestamp 1731220637
transform 1 0 1824 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5923_6
timestamp 1731220637
transform 1 0 1912 0 -1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5922_6
timestamp 1731220637
transform 1 0 1992 0 -1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5921_6
timestamp 1731220637
transform 1 0 1832 0 -1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5920_6
timestamp 1731220637
transform 1 0 1752 0 -1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5919_6
timestamp 1731220637
transform 1 0 1832 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5918_6
timestamp 1731220637
transform 1 0 1896 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5917_6
timestamp 1731220637
transform 1 0 1960 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5916_6
timestamp 1731220637
transform 1 0 2032 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5915_6
timestamp 1731220637
transform 1 0 2112 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5914_6
timestamp 1731220637
transform 1 0 1768 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5913_6
timestamp 1731220637
transform 1 0 1848 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5912_6
timestamp 1731220637
transform 1 0 1936 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5911_6
timestamp 1731220637
transform 1 0 2024 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5910_6
timestamp 1731220637
transform 1 0 2112 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5909_6
timestamp 1731220637
transform 1 0 1704 0 1 100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5908_6
timestamp 1731220637
transform 1 0 1768 0 1 100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5907_6
timestamp 1731220637
transform 1 0 1824 0 1 100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5906_6
timestamp 1731220637
transform 1 0 1880 0 1 100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5905_6
timestamp 1731220637
transform 1 0 1928 0 1 100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5904_6
timestamp 1731220637
transform 1 0 1968 0 1 100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5903_6
timestamp 1731220637
transform 1 0 2008 0 1 100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5902_6
timestamp 1731220637
transform 1 0 2048 0 1 100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5901_6
timestamp 1731220637
transform 1 0 2088 0 1 100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5900_6
timestamp 1731220637
transform 1 0 2136 0 1 100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5899_6
timestamp 1731220637
transform 1 0 2184 0 1 100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5898_6
timestamp 1731220637
transform 1 0 2200 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5897_6
timestamp 1731220637
transform 1 0 2232 0 1 100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5896_6
timestamp 1731220637
transform 1 0 2272 0 1 100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5895_6
timestamp 1731220637
transform 1 0 2312 0 1 100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5894_6
timestamp 1731220637
transform 1 0 2352 0 1 100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5893_6
timestamp 1731220637
transform 1 0 2352 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5892_6
timestamp 1731220637
transform 1 0 2288 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5891_6
timestamp 1731220637
transform 1 0 2352 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5890_6
timestamp 1731220637
transform 1 0 2272 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5889_6
timestamp 1731220637
transform 1 0 2192 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5888_6
timestamp 1731220637
transform 1 0 2240 0 -1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5887_6
timestamp 1731220637
transform 1 0 2152 0 -1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5886_6
timestamp 1731220637
transform 1 0 2072 0 -1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5885_6
timestamp 1731220637
transform 1 0 1912 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5884_6
timestamp 1731220637
transform 1 0 1992 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5883_6
timestamp 1731220637
transform 1 0 2016 0 -1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5882_6
timestamp 1731220637
transform 1 0 2096 0 -1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5881_6
timestamp 1731220637
transform 1 0 2088 0 1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5880_6
timestamp 1731220637
transform 1 0 2024 0 1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5879_6
timestamp 1731220637
transform 1 0 1960 0 1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5878_6
timestamp 1731220637
transform 1 0 1944 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5877_6
timestamp 1731220637
transform 1 0 2040 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5876_6
timestamp 1731220637
transform 1 0 2144 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5875_6
timestamp 1731220637
transform 1 0 2024 0 1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5874_6
timestamp 1731220637
transform 1 0 1936 0 1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5873_6
timestamp 1731220637
transform 1 0 1848 0 1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5872_6
timestamp 1731220637
transform 1 0 1768 0 1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5871_6
timestamp 1731220637
transform 1 0 1752 0 -1 808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5870_6
timestamp 1731220637
transform 1 0 1816 0 -1 808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5869_6
timestamp 1731220637
transform 1 0 1880 0 -1 808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5868_6
timestamp 1731220637
transform 1 0 1944 0 -1 808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5867_6
timestamp 1731220637
transform 1 0 2016 0 -1 808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5866_6
timestamp 1731220637
transform 1 0 1816 0 1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5865_6
timestamp 1731220637
transform 1 0 1888 0 1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5864_6
timestamp 1731220637
transform 1 0 1952 0 1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5863_6
timestamp 1731220637
transform 1 0 2016 0 1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5862_6
timestamp 1731220637
transform 1 0 2080 0 1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5861_6
timestamp 1731220637
transform 1 0 2136 0 1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5860_6
timestamp 1731220637
transform 1 0 2184 0 -1 808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5859_6
timestamp 1731220637
transform 1 0 2272 0 -1 808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5858_6
timestamp 1731220637
transform 1 0 2096 0 -1 808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5857_6
timestamp 1731220637
transform 1 0 2112 0 1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5856_6
timestamp 1731220637
transform 1 0 2200 0 1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5855_6
timestamp 1731220637
transform 1 0 2256 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5854_6
timestamp 1731220637
transform 1 0 2160 0 1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5853_6
timestamp 1731220637
transform 1 0 2232 0 1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5852_6
timestamp 1731220637
transform 1 0 2280 0 -1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5851_6
timestamp 1731220637
transform 1 0 2184 0 -1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5850_6
timestamp 1731220637
transform 1 0 2064 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5849_6
timestamp 1731220637
transform 1 0 2128 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5848_6
timestamp 1731220637
transform 1 0 2192 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5847_6
timestamp 1731220637
transform 1 0 2248 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5846_6
timestamp 1731220637
transform 1 0 2328 0 -1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5845_6
timestamp 1731220637
transform 1 0 2312 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5844_6
timestamp 1731220637
transform 1 0 2352 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5843_6
timestamp 1731220637
transform 1 0 2352 0 -1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5842_6
timestamp 1731220637
transform 1 0 2304 0 1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5841_6
timestamp 1731220637
transform 1 0 2352 0 1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5840_6
timestamp 1731220637
transform 1 0 2352 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5839_6
timestamp 1731220637
transform 1 0 2352 0 1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5838_6
timestamp 1731220637
transform 1 0 2288 0 1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5837_6
timestamp 1731220637
transform 1 0 2352 0 -1 808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5836_6
timestamp 1731220637
transform 1 0 2192 0 1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5835_6
timestamp 1731220637
transform 1 0 2248 0 1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5834_6
timestamp 1731220637
transform 1 0 2312 0 1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5833_6
timestamp 1731220637
transform 1 0 2352 0 1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5832_6
timestamp 1731220637
transform 1 0 2352 0 -1 956
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5831_6
timestamp 1731220637
transform 1 0 2304 0 -1 956
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5830_6
timestamp 1731220637
transform 1 0 2232 0 -1 956
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5829_6
timestamp 1731220637
transform 1 0 2168 0 -1 956
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5828_6
timestamp 1731220637
transform 1 0 1928 0 -1 956
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5827_6
timestamp 1731220637
transform 1 0 2016 0 -1 956
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5826_6
timestamp 1731220637
transform 1 0 2096 0 -1 956
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5825_6
timestamp 1731220637
transform 1 0 2136 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5824_6
timestamp 1731220637
transform 1 0 2200 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5823_6
timestamp 1731220637
transform 1 0 2272 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5822_6
timestamp 1731220637
transform 1 0 2064 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5821_6
timestamp 1731220637
transform 1 0 1824 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5820_6
timestamp 1731220637
transform 1 0 1912 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5819_6
timestamp 1731220637
transform 1 0 1992 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5818_6
timestamp 1731220637
transform 1 0 2016 0 -1 1112
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5817_6
timestamp 1731220637
transform 1 0 2072 0 -1 1112
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5816_6
timestamp 1731220637
transform 1 0 2128 0 -1 1112
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5815_6
timestamp 1731220637
transform 1 0 1960 0 -1 1112
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5814_6
timestamp 1731220637
transform 1 0 1784 0 -1 1112
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5813_6
timestamp 1731220637
transform 1 0 1848 0 -1 1112
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5812_6
timestamp 1731220637
transform 1 0 1904 0 -1 1112
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5811_6
timestamp 1731220637
transform 1 0 2016 0 1 1120
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5810_6
timestamp 1731220637
transform 1 0 2128 0 1 1120
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5809_6
timestamp 1731220637
transform 1 0 2248 0 1 1120
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5808_6
timestamp 1731220637
transform 1 0 1920 0 1 1120
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5807_6
timestamp 1731220637
transform 1 0 1848 0 1 1120
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5806_6
timestamp 1731220637
transform 1 0 1792 0 1 1120
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5805_6
timestamp 1731220637
transform 1 0 1752 0 1 1120
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5804_6
timestamp 1731220637
transform 1 0 1784 0 -1 1260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5803_6
timestamp 1731220637
transform 1 0 1832 0 -1 1260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5802_6
timestamp 1731220637
transform 1 0 1896 0 -1 1260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5801_6
timestamp 1731220637
transform 1 0 1960 0 -1 1260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5800_6
timestamp 1731220637
transform 1 0 2032 0 -1 1260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5799_6
timestamp 1731220637
transform 1 0 2112 0 -1 1260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5798_6
timestamp 1731220637
transform 1 0 1768 0 1 1264
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5797_6
timestamp 1731220637
transform 1 0 1824 0 1 1264
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5796_6
timestamp 1731220637
transform 1 0 1896 0 1 1264
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5795_6
timestamp 1731220637
transform 1 0 1976 0 1 1264
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5794_6
timestamp 1731220637
transform 1 0 2064 0 1 1264
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5793_6
timestamp 1731220637
transform 1 0 2160 0 1 1264
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5792_6
timestamp 1731220637
transform 1 0 1808 0 -1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5791_6
timestamp 1731220637
transform 1 0 1896 0 -1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5790_6
timestamp 1731220637
transform 1 0 1984 0 -1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5789_6
timestamp 1731220637
transform 1 0 2064 0 -1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5788_6
timestamp 1731220637
transform 1 0 1776 0 1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5787_6
timestamp 1731220637
transform 1 0 1864 0 1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5786_6
timestamp 1731220637
transform 1 0 1944 0 1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5785_6
timestamp 1731220637
transform 1 0 2024 0 1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5784_6
timestamp 1731220637
transform 1 0 2096 0 1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5783_6
timestamp 1731220637
transform 1 0 2160 0 1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5782_6
timestamp 1731220637
transform 1 0 2232 0 1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5781_6
timestamp 1731220637
transform 1 0 2304 0 1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5780_6
timestamp 1731220637
transform 1 0 2144 0 -1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5779_6
timestamp 1731220637
transform 1 0 2216 0 -1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5778_6
timestamp 1731220637
transform 1 0 2264 0 1 1264
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5777_6
timestamp 1731220637
transform 1 0 2200 0 -1 1260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5776_6
timestamp 1731220637
transform 1 0 2184 0 -1 1112
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5775_6
timestamp 1731220637
transform 1 0 2248 0 -1 1112
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5774_6
timestamp 1731220637
transform 1 0 2312 0 -1 1112
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5773_6
timestamp 1731220637
transform 1 0 2352 0 -1 1112
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5772_6
timestamp 1731220637
transform 1 0 2352 0 1 1120
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5771_6
timestamp 1731220637
transform 1 0 2288 0 -1 1260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5770_6
timestamp 1731220637
transform 1 0 2352 0 -1 1260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5769_6
timestamp 1731220637
transform 1 0 2352 0 1 1264
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5768_6
timestamp 1731220637
transform 1 0 2352 0 -1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5767_6
timestamp 1731220637
transform 1 0 2296 0 -1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5766_6
timestamp 1731220637
transform 1 0 2352 0 1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5765_6
timestamp 1731220637
transform 1 0 2352 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5764_6
timestamp 1731220637
transform 1 0 2312 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5763_6
timestamp 1731220637
transform 1 0 2352 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5762_6
timestamp 1731220637
transform 1 0 2312 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5761_6
timestamp 1731220637
transform 1 0 2248 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5760_6
timestamp 1731220637
transform 1 0 2248 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5759_6
timestamp 1731220637
transform 1 0 2184 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5758_6
timestamp 1731220637
transform 1 0 2120 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5757_6
timestamp 1731220637
transform 1 0 2048 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5756_6
timestamp 1731220637
transform 1 0 1752 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5755_6
timestamp 1731220637
transform 1 0 1864 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5754_6
timestamp 1731220637
transform 1 0 1960 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5753_6
timestamp 1731220637
transform 1 0 2056 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5752_6
timestamp 1731220637
transform 1 0 2120 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5751_6
timestamp 1731220637
transform 1 0 2184 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5750_6
timestamp 1731220637
transform 1 0 1992 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5749_6
timestamp 1731220637
transform 1 0 1848 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5748_6
timestamp 1731220637
transform 1 0 1920 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5747_6
timestamp 1731220637
transform 1 0 1968 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5746_6
timestamp 1731220637
transform 1 0 2024 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5745_6
timestamp 1731220637
transform 1 0 2080 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5744_6
timestamp 1731220637
transform 1 0 1912 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5743_6
timestamp 1731220637
transform 1 0 1744 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5742_6
timestamp 1731220637
transform 1 0 1800 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5741_6
timestamp 1731220637
transform 1 0 1856 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5740_6
timestamp 1731220637
transform 1 0 1912 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5739_6
timestamp 1731220637
transform 1 0 1968 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5738_6
timestamp 1731220637
transform 1 0 1800 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5737_6
timestamp 1731220637
transform 1 0 1640 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5736_6
timestamp 1731220637
transform 1 0 1696 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5735_6
timestamp 1731220637
transform 1 0 1752 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5734_6
timestamp 1731220637
transform 1 0 1856 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5733_6
timestamp 1731220637
transform 1 0 1888 0 -1 1852
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5732_6
timestamp 1731220637
transform 1 0 1944 0 -1 1852
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5731_6
timestamp 1731220637
transform 1 0 1832 0 -1 1852
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5730_6
timestamp 1731220637
transform 1 0 1776 0 -1 1852
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5729_6
timestamp 1731220637
transform 1 0 1720 0 -1 1852
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5728_6
timestamp 1731220637
transform 1 0 1664 0 -1 1852
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5727_6
timestamp 1731220637
transform 1 0 1704 0 1 1860
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5726_6
timestamp 1731220637
transform 1 0 1800 0 1 1860
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5725_6
timestamp 1731220637
transform 1 0 1912 0 1 1860
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5724_6
timestamp 1731220637
transform 1 0 2024 0 1 1860
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5723_6
timestamp 1731220637
transform 1 0 1864 0 -1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5722_6
timestamp 1731220637
transform 1 0 1816 0 -1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5721_6
timestamp 1731220637
transform 1 0 1760 0 -1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5720_6
timestamp 1731220637
transform 1 0 1712 0 -1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5719_6
timestamp 1731220637
transform 1 0 1672 0 -1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5718_6
timestamp 1731220637
transform 1 0 1632 0 -1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5717_6
timestamp 1731220637
transform 1 0 1592 0 -1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5716_6
timestamp 1731220637
transform 1 0 1552 0 -1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5715_6
timestamp 1731220637
transform 1 0 1512 0 -1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5714_6
timestamp 1731220637
transform 1 0 1392 0 -1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5713_6
timestamp 1731220637
transform 1 0 1432 0 -1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5712_6
timestamp 1731220637
transform 1 0 1472 0 -1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5711_6
timestamp 1731220637
transform 1 0 1504 0 1 1860
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5710_6
timestamp 1731220637
transform 1 0 1560 0 1 1860
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5709_6
timestamp 1731220637
transform 1 0 1624 0 1 1860
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5708_6
timestamp 1731220637
transform 1 0 1456 0 1 1860
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5707_6
timestamp 1731220637
transform 1 0 1416 0 1 1860
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5706_6
timestamp 1731220637
transform 1 0 1376 0 1 1860
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5705_6
timestamp 1731220637
transform 1 0 1336 0 1 1860
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5704_6
timestamp 1731220637
transform 1 0 1352 0 -1 1852
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5703_6
timestamp 1731220637
transform 1 0 1392 0 -1 1852
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5702_6
timestamp 1731220637
transform 1 0 1440 0 -1 1852
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5701_6
timestamp 1731220637
transform 1 0 1496 0 -1 1852
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5700_6
timestamp 1731220637
transform 1 0 1552 0 -1 1852
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5699_6
timestamp 1731220637
transform 1 0 1608 0 -1 1852
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5698_6
timestamp 1731220637
transform 1 0 1384 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5697_6
timestamp 1731220637
transform 1 0 1448 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5696_6
timestamp 1731220637
transform 1 0 1512 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5695_6
timestamp 1731220637
transform 1 0 1576 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5694_6
timestamp 1731220637
transform 1 0 1496 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5693_6
timestamp 1731220637
transform 1 0 1552 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5692_6
timestamp 1731220637
transform 1 0 1616 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5691_6
timestamp 1731220637
transform 1 0 1680 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5690_6
timestamp 1731220637
transform 1 0 1552 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5689_6
timestamp 1731220637
transform 1 0 1624 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5688_6
timestamp 1731220637
transform 1 0 1696 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5687_6
timestamp 1731220637
transform 1 0 1776 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5686_6
timestamp 1731220637
transform 1 0 1616 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5685_6
timestamp 1731220637
transform 1 0 1464 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5684_6
timestamp 1731220637
transform 1 0 1496 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5683_6
timestamp 1731220637
transform 1 0 1456 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5682_6
timestamp 1731220637
transform 1 0 1416 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5681_6
timestamp 1731220637
transform 1 0 1296 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5680_6
timestamp 1731220637
transform 1 0 1336 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5679_6
timestamp 1731220637
transform 1 0 1376 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5678_6
timestamp 1731220637
transform 1 0 1416 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5677_6
timestamp 1731220637
transform 1 0 1456 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5676_6
timestamp 1731220637
transform 1 0 1376 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5675_6
timestamp 1731220637
transform 1 0 1296 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5674_6
timestamp 1731220637
transform 1 0 1336 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5673_6
timestamp 1731220637
transform 1 0 1336 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5672_6
timestamp 1731220637
transform 1 0 1296 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5671_6
timestamp 1731220637
transform 1 0 1184 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5670_6
timestamp 1731220637
transform 1 0 992 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5669_6
timestamp 1731220637
transform 1 0 1064 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5668_6
timestamp 1731220637
transform 1 0 1136 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5667_6
timestamp 1731220637
transform 1 0 1184 0 -1 1840
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5666_6
timestamp 1731220637
transform 1 0 1120 0 -1 1840
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5665_6
timestamp 1731220637
transform 1 0 968 0 -1 1840
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5664_6
timestamp 1731220637
transform 1 0 1040 0 -1 1840
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5663_6
timestamp 1731220637
transform 1 0 1048 0 1 1844
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5662_6
timestamp 1731220637
transform 1 0 1120 0 1 1844
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5661_6
timestamp 1731220637
transform 1 0 912 0 1 1844
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5660_6
timestamp 1731220637
transform 1 0 976 0 1 1844
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5659_6
timestamp 1731220637
transform 1 0 1000 0 -1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5658_6
timestamp 1731220637
transform 1 0 928 0 -1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5657_6
timestamp 1731220637
transform 1 0 856 0 -1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5656_6
timestamp 1731220637
transform 1 0 784 0 -1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5655_6
timestamp 1731220637
transform 1 0 808 0 1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5654_6
timestamp 1731220637
transform 1 0 736 0 1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5653_6
timestamp 1731220637
transform 1 0 544 0 1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5652_6
timestamp 1731220637
transform 1 0 480 0 1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5651_6
timestamp 1731220637
transform 1 0 472 0 -1 2124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5650_6
timestamp 1731220637
transform 1 0 336 0 -1 2124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5649_6
timestamp 1731220637
transform 1 0 408 0 -1 2124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5648_6
timestamp 1731220637
transform 1 0 432 0 1 2132
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5647_6
timestamp 1731220637
transform 1 0 272 0 1 2132
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5646_6
timestamp 1731220637
transform 1 0 352 0 1 2132
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5645_6
timestamp 1731220637
transform 1 0 400 0 -1 2268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5644_6
timestamp 1731220637
transform 1 0 328 0 -1 2268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5643_6
timestamp 1731220637
transform 1 0 272 0 -1 2268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5642_6
timestamp 1731220637
transform 1 0 216 0 -1 2268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5641_6
timestamp 1731220637
transform 1 0 176 0 -1 2268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5640_6
timestamp 1731220637
transform 1 0 136 0 -1 2268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5639_6
timestamp 1731220637
transform 1 0 128 0 1 2132
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5638_6
timestamp 1731220637
transform 1 0 200 0 1 2132
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5637_6
timestamp 1731220637
transform 1 0 264 0 -1 2124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5636_6
timestamp 1731220637
transform 1 0 184 0 -1 2124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5635_6
timestamp 1731220637
transform 1 0 128 0 -1 2124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5634_6
timestamp 1731220637
transform 1 0 128 0 1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5633_6
timestamp 1731220637
transform 1 0 168 0 1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5632_6
timestamp 1731220637
transform 1 0 208 0 1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5631_6
timestamp 1731220637
transform 1 0 272 0 1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5630_6
timestamp 1731220637
transform 1 0 344 0 1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5629_6
timestamp 1731220637
transform 1 0 416 0 1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5628_6
timestamp 1731220637
transform 1 0 128 0 -1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5627_6
timestamp 1731220637
transform 1 0 168 0 -1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5626_6
timestamp 1731220637
transform 1 0 208 0 -1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5625_6
timestamp 1731220637
transform 1 0 264 0 -1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5624_6
timestamp 1731220637
transform 1 0 336 0 -1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5623_6
timestamp 1731220637
transform 1 0 408 0 -1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5622_6
timestamp 1731220637
transform 1 0 488 0 -1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5621_6
timestamp 1731220637
transform 1 0 240 0 1 1844
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5620_6
timestamp 1731220637
transform 1 0 280 0 1 1844
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5619_6
timestamp 1731220637
transform 1 0 320 0 1 1844
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5618_6
timestamp 1731220637
transform 1 0 360 0 1 1844
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5617_6
timestamp 1731220637
transform 1 0 408 0 1 1844
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5616_6
timestamp 1731220637
transform 1 0 464 0 1 1844
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5615_6
timestamp 1731220637
transform 1 0 528 0 1 1844
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5614_6
timestamp 1731220637
transform 1 0 592 0 1 1844
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5613_6
timestamp 1731220637
transform 1 0 392 0 -1 1840
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5612_6
timestamp 1731220637
transform 1 0 432 0 -1 1840
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5611_6
timestamp 1731220637
transform 1 0 472 0 -1 1840
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5610_6
timestamp 1731220637
transform 1 0 512 0 -1 1840
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5609_6
timestamp 1731220637
transform 1 0 560 0 -1 1840
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5608_6
timestamp 1731220637
transform 1 0 616 0 -1 1840
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5607_6
timestamp 1731220637
transform 1 0 680 0 -1 1840
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5606_6
timestamp 1731220637
transform 1 0 640 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5605_6
timestamp 1731220637
transform 1 0 600 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5604_6
timestamp 1731220637
transform 1 0 560 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5603_6
timestamp 1731220637
transform 1 0 520 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5602_6
timestamp 1731220637
transform 1 0 480 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5601_6
timestamp 1731220637
transform 1 0 440 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5600_6
timestamp 1731220637
transform 1 0 400 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5599_6
timestamp 1731220637
transform 1 0 440 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5598_6
timestamp 1731220637
transform 1 0 488 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5597_6
timestamp 1731220637
transform 1 0 536 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5596_6
timestamp 1731220637
transform 1 0 392 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5595_6
timestamp 1731220637
transform 1 0 272 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5594_6
timestamp 1731220637
transform 1 0 312 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5593_6
timestamp 1731220637
transform 1 0 352 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5592_6
timestamp 1731220637
transform 1 0 384 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5591_6
timestamp 1731220637
transform 1 0 464 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5590_6
timestamp 1731220637
transform 1 0 552 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5589_6
timestamp 1731220637
transform 1 0 304 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5588_6
timestamp 1731220637
transform 1 0 248 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5587_6
timestamp 1731220637
transform 1 0 208 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5586_6
timestamp 1731220637
transform 1 0 128 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5585_6
timestamp 1731220637
transform 1 0 168 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5584_6
timestamp 1731220637
transform 1 0 144 0 -1 1556
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5583_6
timestamp 1731220637
transform 1 0 192 0 -1 1556
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5582_6
timestamp 1731220637
transform 1 0 256 0 -1 1556
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5581_6
timestamp 1731220637
transform 1 0 336 0 -1 1556
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5580_6
timestamp 1731220637
transform 1 0 432 0 -1 1556
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5579_6
timestamp 1731220637
transform 1 0 528 0 -1 1556
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5578_6
timestamp 1731220637
transform 1 0 632 0 -1 1556
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5577_6
timestamp 1731220637
transform 1 0 312 0 1 1416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5576_6
timestamp 1731220637
transform 1 0 352 0 1 1416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5575_6
timestamp 1731220637
transform 1 0 392 0 1 1416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5574_6
timestamp 1731220637
transform 1 0 440 0 1 1416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5573_6
timestamp 1731220637
transform 1 0 496 0 1 1416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5572_6
timestamp 1731220637
transform 1 0 552 0 1 1416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5571_6
timestamp 1731220637
transform 1 0 608 0 1 1416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5570_6
timestamp 1731220637
transform 1 0 552 0 -1 1412
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5569_6
timestamp 1731220637
transform 1 0 496 0 -1 1412
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5568_6
timestamp 1731220637
transform 1 0 440 0 -1 1412
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5567_6
timestamp 1731220637
transform 1 0 384 0 -1 1412
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5566_6
timestamp 1731220637
transform 1 0 336 0 -1 1412
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5565_6
timestamp 1731220637
transform 1 0 256 0 -1 1412
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5564_6
timestamp 1731220637
transform 1 0 296 0 -1 1412
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5563_6
timestamp 1731220637
transform 1 0 320 0 1 1272
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5562_6
timestamp 1731220637
transform 1 0 400 0 1 1272
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5561_6
timestamp 1731220637
transform 1 0 488 0 1 1272
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5560_6
timestamp 1731220637
transform 1 0 248 0 1 1272
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5559_6
timestamp 1731220637
transform 1 0 128 0 1 1272
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5558_6
timestamp 1731220637
transform 1 0 168 0 1 1272
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5557_6
timestamp 1731220637
transform 1 0 208 0 1 1272
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5556_6
timestamp 1731220637
transform 1 0 240 0 -1 1268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5555_6
timestamp 1731220637
transform 1 0 320 0 -1 1268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5554_6
timestamp 1731220637
transform 1 0 408 0 -1 1268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5553_6
timestamp 1731220637
transform 1 0 168 0 -1 1268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5552_6
timestamp 1731220637
transform 1 0 128 0 -1 1268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5551_6
timestamp 1731220637
transform 1 0 128 0 1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5550_6
timestamp 1731220637
transform 1 0 168 0 1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5549_6
timestamp 1731220637
transform 1 0 224 0 1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5548_6
timestamp 1731220637
transform 1 0 296 0 1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5547_6
timestamp 1731220637
transform 1 0 376 0 1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5546_6
timestamp 1731220637
transform 1 0 128 0 -1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5545_6
timestamp 1731220637
transform 1 0 208 0 -1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5544_6
timestamp 1731220637
transform 1 0 296 0 -1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5543_6
timestamp 1731220637
transform 1 0 384 0 -1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5542_6
timestamp 1731220637
transform 1 0 192 0 1 984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5541_6
timestamp 1731220637
transform 1 0 232 0 1 984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5540_6
timestamp 1731220637
transform 1 0 280 0 1 984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5539_6
timestamp 1731220637
transform 1 0 336 0 1 984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5538_6
timestamp 1731220637
transform 1 0 384 0 1 984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5537_6
timestamp 1731220637
transform 1 0 288 0 -1 972
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5536_6
timestamp 1731220637
transform 1 0 336 0 -1 972
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5535_6
timestamp 1731220637
transform 1 0 392 0 -1 972
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5534_6
timestamp 1731220637
transform 1 0 464 0 -1 972
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5533_6
timestamp 1731220637
transform 1 0 528 0 1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5532_6
timestamp 1731220637
transform 1 0 448 0 1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5531_6
timestamp 1731220637
transform 1 0 368 0 1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5530_6
timestamp 1731220637
transform 1 0 248 0 1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5529_6
timestamp 1731220637
transform 1 0 304 0 1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5528_6
timestamp 1731220637
transform 1 0 304 0 -1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5527_6
timestamp 1731220637
transform 1 0 376 0 -1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5526_6
timestamp 1731220637
transform 1 0 184 0 -1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5525_6
timestamp 1731220637
transform 1 0 240 0 -1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5524_6
timestamp 1731220637
transform 1 0 272 0 1 692
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5523_6
timestamp 1731220637
transform 1 0 344 0 1 692
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5522_6
timestamp 1731220637
transform 1 0 208 0 1 692
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5521_6
timestamp 1731220637
transform 1 0 128 0 1 692
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5520_6
timestamp 1731220637
transform 1 0 168 0 1 692
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5519_6
timestamp 1731220637
transform 1 0 168 0 -1 684
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5518_6
timestamp 1731220637
transform 1 0 224 0 -1 684
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5517_6
timestamp 1731220637
transform 1 0 280 0 -1 684
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5516_6
timestamp 1731220637
transform 1 0 128 0 -1 684
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5515_6
timestamp 1731220637
transform 1 0 128 0 1 548
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5514_6
timestamp 1731220637
transform 1 0 176 0 1 548
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5513_6
timestamp 1731220637
transform 1 0 248 0 1 548
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5512_6
timestamp 1731220637
transform 1 0 320 0 1 548
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5511_6
timestamp 1731220637
transform 1 0 280 0 -1 544
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5510_6
timestamp 1731220637
transform 1 0 144 0 -1 544
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5509_6
timestamp 1731220637
transform 1 0 216 0 -1 544
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5508_6
timestamp 1731220637
transform 1 0 232 0 1 408
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5507_6
timestamp 1731220637
transform 1 0 272 0 1 408
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5506_6
timestamp 1731220637
transform 1 0 320 0 1 408
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5505_6
timestamp 1731220637
transform 1 0 376 0 1 408
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5504_6
timestamp 1731220637
transform 1 0 264 0 -1 404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5503_6
timestamp 1731220637
transform 1 0 216 0 -1 404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5502_6
timestamp 1731220637
transform 1 0 176 0 -1 404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5501_6
timestamp 1731220637
transform 1 0 136 0 -1 404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5500_6
timestamp 1731220637
transform 1 0 168 0 1 260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5499_6
timestamp 1731220637
transform 1 0 208 0 1 260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5498_6
timestamp 1731220637
transform 1 0 248 0 1 260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5497_6
timestamp 1731220637
transform 1 0 128 0 1 260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5496_6
timestamp 1731220637
transform 1 0 128 0 -1 252
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5495_6
timestamp 1731220637
transform 1 0 288 0 1 260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5494_6
timestamp 1731220637
transform 1 0 328 0 1 260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5493_6
timestamp 1731220637
transform 1 0 384 0 1 260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5492_6
timestamp 1731220637
transform 1 0 440 0 1 260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5491_6
timestamp 1731220637
transform 1 0 328 0 -1 404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5490_6
timestamp 1731220637
transform 1 0 392 0 -1 404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5489_6
timestamp 1731220637
transform 1 0 464 0 -1 404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5488_6
timestamp 1731220637
transform 1 0 536 0 -1 404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5487_6
timestamp 1731220637
transform 1 0 560 0 1 408
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5486_6
timestamp 1731220637
transform 1 0 496 0 1 408
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5485_6
timestamp 1731220637
transform 1 0 432 0 1 408
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5484_6
timestamp 1731220637
transform 1 0 344 0 -1 544
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5483_6
timestamp 1731220637
transform 1 0 408 0 -1 544
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5482_6
timestamp 1731220637
transform 1 0 472 0 -1 544
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5481_6
timestamp 1731220637
transform 1 0 544 0 -1 544
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5480_6
timestamp 1731220637
transform 1 0 552 0 1 548
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5479_6
timestamp 1731220637
transform 1 0 392 0 1 548
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5478_6
timestamp 1731220637
transform 1 0 472 0 1 548
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5477_6
timestamp 1731220637
transform 1 0 496 0 -1 684
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5476_6
timestamp 1731220637
transform 1 0 448 0 -1 684
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5475_6
timestamp 1731220637
transform 1 0 336 0 -1 684
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5474_6
timestamp 1731220637
transform 1 0 392 0 -1 684
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5473_6
timestamp 1731220637
transform 1 0 416 0 1 692
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5472_6
timestamp 1731220637
transform 1 0 488 0 1 692
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5471_6
timestamp 1731220637
transform 1 0 456 0 -1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5470_6
timestamp 1731220637
transform 1 0 536 0 -1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5469_6
timestamp 1731220637
transform 1 0 608 0 -1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5468_6
timestamp 1731220637
transform 1 0 616 0 1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5467_6
timestamp 1731220637
transform 1 0 704 0 1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5466_6
timestamp 1731220637
transform 1 0 720 0 -1 972
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5465_6
timestamp 1731220637
transform 1 0 632 0 -1 972
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5464_6
timestamp 1731220637
transform 1 0 544 0 -1 972
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5463_6
timestamp 1731220637
transform 1 0 432 0 1 984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5462_6
timestamp 1731220637
transform 1 0 480 0 1 984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5461_6
timestamp 1731220637
transform 1 0 528 0 1 984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5460_6
timestamp 1731220637
transform 1 0 552 0 -1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5459_6
timestamp 1731220637
transform 1 0 472 0 -1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5458_6
timestamp 1731220637
transform 1 0 464 0 1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5457_6
timestamp 1731220637
transform 1 0 552 0 1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5456_6
timestamp 1731220637
transform 1 0 632 0 1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5455_6
timestamp 1731220637
transform 1 0 664 0 -1 1268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5454_6
timestamp 1731220637
transform 1 0 584 0 -1 1268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5453_6
timestamp 1731220637
transform 1 0 496 0 -1 1268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5452_6
timestamp 1731220637
transform 1 0 576 0 1 1272
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5451_6
timestamp 1731220637
transform 1 0 664 0 1 1272
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5450_6
timestamp 1731220637
transform 1 0 752 0 1 1272
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5449_6
timestamp 1731220637
transform 1 0 616 0 -1 1412
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5448_6
timestamp 1731220637
transform 1 0 680 0 -1 1412
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5447_6
timestamp 1731220637
transform 1 0 744 0 -1 1412
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5446_6
timestamp 1731220637
transform 1 0 808 0 -1 1412
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5445_6
timestamp 1731220637
transform 1 0 664 0 1 1416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5444_6
timestamp 1731220637
transform 1 0 728 0 1 1416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5443_6
timestamp 1731220637
transform 1 0 792 0 1 1416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5442_6
timestamp 1731220637
transform 1 0 848 0 1 1416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5441_6
timestamp 1731220637
transform 1 0 904 0 1 1416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5440_6
timestamp 1731220637
transform 1 0 960 0 1 1416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5439_6
timestamp 1731220637
transform 1 0 1016 0 -1 1412
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5438_6
timestamp 1731220637
transform 1 0 944 0 -1 1412
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5437_6
timestamp 1731220637
transform 1 0 872 0 -1 1412
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5436_6
timestamp 1731220637
transform 1 0 832 0 1 1272
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5435_6
timestamp 1731220637
transform 1 0 912 0 1 1272
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5434_6
timestamp 1731220637
transform 1 0 1000 0 1 1272
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5433_6
timestamp 1731220637
transform 1 0 1088 0 1 1272
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5432_6
timestamp 1731220637
transform 1 0 1064 0 -1 1268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5431_6
timestamp 1731220637
transform 1 0 1000 0 -1 1268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5430_6
timestamp 1731220637
transform 1 0 936 0 -1 1268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5429_6
timestamp 1731220637
transform 1 0 872 0 -1 1268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5428_6
timestamp 1731220637
transform 1 0 736 0 -1 1268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5427_6
timestamp 1731220637
transform 1 0 808 0 -1 1268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5426_6
timestamp 1731220637
transform 1 0 864 0 1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5425_6
timestamp 1731220637
transform 1 0 792 0 1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5424_6
timestamp 1731220637
transform 1 0 712 0 1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5423_6
timestamp 1731220637
transform 1 0 704 0 -1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5422_6
timestamp 1731220637
transform 1 0 632 0 -1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5421_6
timestamp 1731220637
transform 1 0 576 0 1 984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5420_6
timestamp 1731220637
transform 1 0 624 0 1 984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5419_6
timestamp 1731220637
transform 1 0 672 0 1 984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5418_6
timestamp 1731220637
transform 1 0 720 0 1 984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5417_6
timestamp 1731220637
transform 1 0 776 0 1 984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5416_6
timestamp 1731220637
transform 1 0 832 0 1 984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5415_6
timestamp 1731220637
transform 1 0 888 0 1 984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5414_6
timestamp 1731220637
transform 1 0 952 0 1 984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5413_6
timestamp 1731220637
transform 1 0 768 0 -1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5412_6
timestamp 1731220637
transform 1 0 832 0 -1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5411_6
timestamp 1731220637
transform 1 0 896 0 -1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5410_6
timestamp 1731220637
transform 1 0 952 0 -1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5409_6
timestamp 1731220637
transform 1 0 1016 0 -1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5408_6
timestamp 1731220637
transform 1 0 928 0 1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5407_6
timestamp 1731220637
transform 1 0 984 0 1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5406_6
timestamp 1731220637
transform 1 0 1040 0 1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5405_6
timestamp 1731220637
transform 1 0 1096 0 1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5404_6
timestamp 1731220637
transform 1 0 1144 0 1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5403_6
timestamp 1731220637
transform 1 0 1184 0 1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5402_6
timestamp 1731220637
transform 1 0 1080 0 -1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5401_6
timestamp 1731220637
transform 1 0 1144 0 -1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5400_6
timestamp 1731220637
transform 1 0 1184 0 -1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5399_6
timestamp 1731220637
transform 1 0 1184 0 1 984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5398_6
timestamp 1731220637
transform 1 0 1144 0 1 984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5397_6
timestamp 1731220637
transform 1 0 1016 0 1 984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5396_6
timestamp 1731220637
transform 1 0 1080 0 1 984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5395_6
timestamp 1731220637
transform 1 0 1080 0 -1 972
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5394_6
timestamp 1731220637
transform 1 0 1144 0 -1 972
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5393_6
timestamp 1731220637
transform 1 0 1184 0 -1 972
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5392_6
timestamp 1731220637
transform 1 0 800 0 -1 972
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5391_6
timestamp 1731220637
transform 1 0 880 0 -1 972
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5390_6
timestamp 1731220637
transform 1 0 952 0 -1 972
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5389_6
timestamp 1731220637
transform 1 0 1016 0 -1 972
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5388_6
timestamp 1731220637
transform 1 0 1048 0 1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5387_6
timestamp 1731220637
transform 1 0 1112 0 1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5386_6
timestamp 1731220637
transform 1 0 1176 0 1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5385_6
timestamp 1731220637
transform 1 0 992 0 1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5384_6
timestamp 1731220637
transform 1 0 928 0 1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5383_6
timestamp 1731220637
transform 1 0 784 0 1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5382_6
timestamp 1731220637
transform 1 0 856 0 1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5381_6
timestamp 1731220637
transform 1 0 920 0 -1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5380_6
timestamp 1731220637
transform 1 0 976 0 -1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5379_6
timestamp 1731220637
transform 1 0 1040 0 -1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5378_6
timestamp 1731220637
transform 1 0 864 0 -1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5377_6
timestamp 1731220637
transform 1 0 680 0 -1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5376_6
timestamp 1731220637
transform 1 0 744 0 -1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5375_6
timestamp 1731220637
transform 1 0 808 0 -1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5374_6
timestamp 1731220637
transform 1 0 872 0 1 692
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5373_6
timestamp 1731220637
transform 1 0 976 0 1 692
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5372_6
timestamp 1731220637
transform 1 0 1088 0 1 692
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5371_6
timestamp 1731220637
transform 1 0 776 0 1 692
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5370_6
timestamp 1731220637
transform 1 0 552 0 1 692
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5369_6
timestamp 1731220637
transform 1 0 616 0 1 692
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5368_6
timestamp 1731220637
transform 1 0 688 0 1 692
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5367_6
timestamp 1731220637
transform 1 0 760 0 -1 684
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5366_6
timestamp 1731220637
transform 1 0 832 0 -1 684
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5365_6
timestamp 1731220637
transform 1 0 688 0 -1 684
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5364_6
timestamp 1731220637
transform 1 0 552 0 -1 684
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5363_6
timestamp 1731220637
transform 1 0 616 0 -1 684
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5362_6
timestamp 1731220637
transform 1 0 632 0 1 548
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5361_6
timestamp 1731220637
transform 1 0 712 0 1 548
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5360_6
timestamp 1731220637
transform 1 0 792 0 1 548
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5359_6
timestamp 1731220637
transform 1 0 616 0 -1 544
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5358_6
timestamp 1731220637
transform 1 0 688 0 -1 544
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5357_6
timestamp 1731220637
transform 1 0 760 0 -1 544
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5356_6
timestamp 1731220637
transform 1 0 832 0 -1 544
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5355_6
timestamp 1731220637
transform 1 0 624 0 1 408
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5354_6
timestamp 1731220637
transform 1 0 688 0 1 408
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5353_6
timestamp 1731220637
transform 1 0 752 0 1 408
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5352_6
timestamp 1731220637
transform 1 0 816 0 1 408
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5351_6
timestamp 1731220637
transform 1 0 880 0 1 408
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5350_6
timestamp 1731220637
transform 1 0 856 0 -1 404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5349_6
timestamp 1731220637
transform 1 0 800 0 -1 404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5348_6
timestamp 1731220637
transform 1 0 744 0 -1 404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5347_6
timestamp 1731220637
transform 1 0 680 0 -1 404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5346_6
timestamp 1731220637
transform 1 0 608 0 -1 404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5345_6
timestamp 1731220637
transform 1 0 584 0 1 260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5344_6
timestamp 1731220637
transform 1 0 632 0 1 260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5343_6
timestamp 1731220637
transform 1 0 680 0 1 260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5342_6
timestamp 1731220637
transform 1 0 728 0 1 260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5341_6
timestamp 1731220637
transform 1 0 776 0 1 260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5340_6
timestamp 1731220637
transform 1 0 688 0 -1 252
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5339_6
timestamp 1731220637
transform 1 0 728 0 -1 252
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5338_6
timestamp 1731220637
transform 1 0 776 0 -1 252
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5337_6
timestamp 1731220637
transform 1 0 824 0 -1 252
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5336_6
timestamp 1731220637
transform 1 0 872 0 -1 252
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5335_6
timestamp 1731220637
transform 1 0 920 0 -1 252
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5334_6
timestamp 1731220637
transform 1 0 968 0 -1 252
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5333_6
timestamp 1731220637
transform 1 0 1016 0 -1 252
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5332_6
timestamp 1731220637
transform 1 0 624 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5331_6
timestamp 1731220637
transform 1 0 664 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5330_6
timestamp 1731220637
transform 1 0 704 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5329_6
timestamp 1731220637
transform 1 0 744 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5328_6
timestamp 1731220637
transform 1 0 784 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5327_6
timestamp 1731220637
transform 1 0 824 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5326_6
timestamp 1731220637
transform 1 0 864 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5325_6
timestamp 1731220637
transform 1 0 904 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5324_6
timestamp 1731220637
transform 1 0 944 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5323_6
timestamp 1731220637
transform 1 0 984 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5322_6
timestamp 1731220637
transform 1 0 1024 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5321_6
timestamp 1731220637
transform 1 0 1064 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5320_6
timestamp 1731220637
transform 1 0 1104 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5319_6
timestamp 1731220637
transform 1 0 1144 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5318_6
timestamp 1731220637
transform 1 0 1184 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5317_6
timestamp 1731220637
transform 1 0 1296 0 1 100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5316_6
timestamp 1731220637
transform 1 0 1336 0 1 100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5315_6
timestamp 1731220637
transform 1 0 1376 0 1 100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5314_6
timestamp 1731220637
transform 1 0 1416 0 1 100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5313_6
timestamp 1731220637
transform 1 0 1456 0 1 100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5312_6
timestamp 1731220637
transform 1 0 1512 0 1 100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5311_6
timestamp 1731220637
transform 1 0 1576 0 1 100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5310_6
timestamp 1731220637
transform 1 0 1640 0 1 100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5309_6
timestamp 1731220637
transform 1 0 1360 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5308_6
timestamp 1731220637
transform 1 0 1400 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5307_6
timestamp 1731220637
transform 1 0 1448 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5306_6
timestamp 1731220637
transform 1 0 1504 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5305_6
timestamp 1731220637
transform 1 0 1560 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5304_6
timestamp 1731220637
transform 1 0 1624 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5303_6
timestamp 1731220637
transform 1 0 1696 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5302_6
timestamp 1731220637
transform 1 0 1624 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5301_6
timestamp 1731220637
transform 1 0 1664 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5300_6
timestamp 1731220637
transform 1 0 1704 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5299_6
timestamp 1731220637
transform 1 0 1744 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5298_6
timestamp 1731220637
transform 1 0 1784 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5297_6
timestamp 1731220637
transform 1 0 1504 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5296_6
timestamp 1731220637
transform 1 0 1544 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5295_6
timestamp 1731220637
transform 1 0 1584 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5294_6
timestamp 1731220637
transform 1 0 1600 0 -1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5293_6
timestamp 1731220637
transform 1 0 1672 0 -1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5292_6
timestamp 1731220637
transform 1 0 1536 0 -1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5291_6
timestamp 1731220637
transform 1 0 1480 0 -1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5290_6
timestamp 1731220637
transform 1 0 1432 0 -1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5289_6
timestamp 1731220637
transform 1 0 1392 0 -1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5288_6
timestamp 1731220637
transform 1 0 1352 0 -1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5287_6
timestamp 1731220637
transform 1 0 1296 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5286_6
timestamp 1731220637
transform 1 0 1336 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5285_6
timestamp 1731220637
transform 1 0 1376 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5284_6
timestamp 1731220637
transform 1 0 1440 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5283_6
timestamp 1731220637
transform 1 0 1528 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5282_6
timestamp 1731220637
transform 1 0 1624 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5281_6
timestamp 1731220637
transform 1 0 1728 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5280_6
timestamp 1731220637
transform 1 0 1400 0 -1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5279_6
timestamp 1731220637
transform 1 0 1440 0 -1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5278_6
timestamp 1731220637
transform 1 0 1480 0 -1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5277_6
timestamp 1731220637
transform 1 0 1528 0 -1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5276_6
timestamp 1731220637
transform 1 0 1584 0 -1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5275_6
timestamp 1731220637
transform 1 0 1640 0 -1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5274_6
timestamp 1731220637
transform 1 0 1704 0 -1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5273_6
timestamp 1731220637
transform 1 0 1672 0 1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5272_6
timestamp 1731220637
transform 1 0 1712 0 1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5271_6
timestamp 1731220637
transform 1 0 1752 0 1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5270_6
timestamp 1731220637
transform 1 0 1800 0 1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5269_6
timestamp 1731220637
transform 1 0 1632 0 1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5268_6
timestamp 1731220637
transform 1 0 1592 0 1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5267_6
timestamp 1731220637
transform 1 0 1552 0 1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5266_6
timestamp 1731220637
transform 1 0 1584 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5265_6
timestamp 1731220637
transform 1 0 1528 0 1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5264_6
timestamp 1731220637
transform 1 0 1448 0 1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5263_6
timestamp 1731220637
transform 1 0 1472 0 -1 808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5262_6
timestamp 1731220637
transform 1 0 1544 0 -1 808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5261_6
timestamp 1731220637
transform 1 0 1528 0 1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5260_6
timestamp 1731220637
transform 1 0 1464 0 1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5259_6
timestamp 1731220637
transform 1 0 1456 0 -1 956
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5258_6
timestamp 1731220637
transform 1 0 1496 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5257_6
timestamp 1731220637
transform 1 0 1616 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5256_6
timestamp 1731220637
transform 1 0 1728 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5255_6
timestamp 1731220637
transform 1 0 1528 0 -1 1112
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5254_6
timestamp 1731220637
transform 1 0 1592 0 -1 1112
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5253_6
timestamp 1731220637
transform 1 0 1656 0 -1 1112
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5252_6
timestamp 1731220637
transform 1 0 1720 0 -1 1112
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5251_6
timestamp 1731220637
transform 1 0 1552 0 1 1120
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5250_6
timestamp 1731220637
transform 1 0 1592 0 1 1120
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5249_6
timestamp 1731220637
transform 1 0 1632 0 1 1120
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5248_6
timestamp 1731220637
transform 1 0 1672 0 1 1120
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5247_6
timestamp 1731220637
transform 1 0 1712 0 1 1120
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5246_6
timestamp 1731220637
transform 1 0 1744 0 -1 1260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5245_6
timestamp 1731220637
transform 1 0 1704 0 -1 1260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5244_6
timestamp 1731220637
transform 1 0 1664 0 -1 1260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5243_6
timestamp 1731220637
transform 1 0 1624 0 -1 1260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5242_6
timestamp 1731220637
transform 1 0 1504 0 -1 1260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5241_6
timestamp 1731220637
transform 1 0 1544 0 -1 1260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5240_6
timestamp 1731220637
transform 1 0 1584 0 -1 1260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5239_6
timestamp 1731220637
transform 1 0 1608 0 1 1264
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5238_6
timestamp 1731220637
transform 1 0 1664 0 1 1264
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5237_6
timestamp 1731220637
transform 1 0 1712 0 1 1264
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5236_6
timestamp 1731220637
transform 1 0 1560 0 1 1264
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5235_6
timestamp 1731220637
transform 1 0 1440 0 1 1264
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5234_6
timestamp 1731220637
transform 1 0 1480 0 1 1264
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5233_6
timestamp 1731220637
transform 1 0 1520 0 1 1264
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5232_6
timestamp 1731220637
transform 1 0 1544 0 -1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5231_6
timestamp 1731220637
transform 1 0 1632 0 -1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5230_6
timestamp 1731220637
transform 1 0 1720 0 -1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5229_6
timestamp 1731220637
transform 1 0 1464 0 -1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5228_6
timestamp 1731220637
transform 1 0 1296 0 -1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5227_6
timestamp 1731220637
transform 1 0 1336 0 -1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5226_6
timestamp 1731220637
transform 1 0 1392 0 -1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5225_6
timestamp 1731220637
transform 1 0 1472 0 1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5224_6
timestamp 1731220637
transform 1 0 1576 0 1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5223_6
timestamp 1731220637
transform 1 0 1680 0 1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5222_6
timestamp 1731220637
transform 1 0 1368 0 1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5221_6
timestamp 1731220637
transform 1 0 1296 0 1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5220_6
timestamp 1731220637
transform 1 0 1184 0 1 1416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5219_6
timestamp 1731220637
transform 1 0 1016 0 1 1416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5218_6
timestamp 1731220637
transform 1 0 1080 0 1 1416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5217_6
timestamp 1731220637
transform 1 0 1144 0 1 1416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5216_6
timestamp 1731220637
transform 1 0 1184 0 -1 1556
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5215_6
timestamp 1731220637
transform 1 0 1112 0 -1 1556
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5214_6
timestamp 1731220637
transform 1 0 1040 0 -1 1556
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5213_6
timestamp 1731220637
transform 1 0 968 0 -1 1556
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5212_6
timestamp 1731220637
transform 1 0 728 0 -1 1556
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5211_6
timestamp 1731220637
transform 1 0 816 0 -1 1556
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5210_6
timestamp 1731220637
transform 1 0 896 0 -1 1556
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5209_6
timestamp 1731220637
transform 1 0 912 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5208_6
timestamp 1731220637
transform 1 0 976 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5207_6
timestamp 1731220637
transform 1 0 1040 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5206_6
timestamp 1731220637
transform 1 0 848 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5205_6
timestamp 1731220637
transform 1 0 632 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5204_6
timestamp 1731220637
transform 1 0 712 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5203_6
timestamp 1731220637
transform 1 0 784 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5202_6
timestamp 1731220637
transform 1 0 832 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5201_6
timestamp 1731220637
transform 1 0 888 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5200_6
timestamp 1731220637
transform 1 0 776 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5199_6
timestamp 1731220637
transform 1 0 728 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5198_6
timestamp 1731220637
transform 1 0 680 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5197_6
timestamp 1731220637
transform 1 0 584 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5196_6
timestamp 1731220637
transform 1 0 632 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5195_6
timestamp 1731220637
transform 1 0 688 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5194_6
timestamp 1731220637
transform 1 0 744 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5193_6
timestamp 1731220637
transform 1 0 800 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5192_6
timestamp 1731220637
transform 1 0 864 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5191_6
timestamp 1731220637
transform 1 0 928 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5190_6
timestamp 1731220637
transform 1 0 896 0 -1 1840
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5189_6
timestamp 1731220637
transform 1 0 752 0 -1 1840
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5188_6
timestamp 1731220637
transform 1 0 824 0 -1 1840
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5187_6
timestamp 1731220637
transform 1 0 848 0 1 1844
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5186_6
timestamp 1731220637
transform 1 0 784 0 1 1844
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5185_6
timestamp 1731220637
transform 1 0 720 0 1 1844
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5184_6
timestamp 1731220637
transform 1 0 656 0 1 1844
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5183_6
timestamp 1731220637
transform 1 0 712 0 -1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5182_6
timestamp 1731220637
transform 1 0 640 0 -1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5181_6
timestamp 1731220637
transform 1 0 568 0 -1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5180_6
timestamp 1731220637
transform 1 0 608 0 1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5179_6
timestamp 1731220637
transform 1 0 672 0 1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5178_6
timestamp 1731220637
transform 1 0 664 0 -1 2124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5177_6
timestamp 1731220637
transform 1 0 600 0 -1 2124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5176_6
timestamp 1731220637
transform 1 0 536 0 -1 2124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5175_6
timestamp 1731220637
transform 1 0 592 0 1 2132
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5174_6
timestamp 1731220637
transform 1 0 512 0 1 2132
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5173_6
timestamp 1731220637
transform 1 0 472 0 -1 2268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5172_6
timestamp 1731220637
transform 1 0 552 0 -1 2268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5171_6
timestamp 1731220637
transform 1 0 544 0 1 2276
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5170_6
timestamp 1731220637
transform 1 0 464 0 1 2276
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5169_6
timestamp 1731220637
transform 1 0 264 0 1 2276
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5168_6
timestamp 1731220637
transform 1 0 320 0 1 2276
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5167_6
timestamp 1731220637
transform 1 0 392 0 1 2276
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5166_6
timestamp 1731220637
transform 1 0 392 0 -1 2416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5165_6
timestamp 1731220637
transform 1 0 320 0 -1 2416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5164_6
timestamp 1731220637
transform 1 0 256 0 -1 2416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5163_6
timestamp 1731220637
transform 1 0 192 0 -1 2416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5162_6
timestamp 1731220637
transform 1 0 224 0 1 2424
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5161_6
timestamp 1731220637
transform 1 0 264 0 1 2424
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5160_6
timestamp 1731220637
transform 1 0 304 0 1 2424
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5159_6
timestamp 1731220637
transform 1 0 344 0 1 2424
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5158_6
timestamp 1731220637
transform 1 0 392 0 1 2424
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5157_6
timestamp 1731220637
transform 1 0 448 0 1 2424
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5156_6
timestamp 1731220637
transform 1 0 504 0 1 2424
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5155_6
timestamp 1731220637
transform 1 0 568 0 1 2424
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5154_6
timestamp 1731220637
transform 1 0 632 0 1 2424
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5153_6
timestamp 1731220637
transform 1 0 464 0 -1 2416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5152_6
timestamp 1731220637
transform 1 0 536 0 -1 2416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5151_6
timestamp 1731220637
transform 1 0 608 0 -1 2416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5150_6
timestamp 1731220637
transform 1 0 680 0 -1 2416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5149_6
timestamp 1731220637
transform 1 0 704 0 1 2276
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5148_6
timestamp 1731220637
transform 1 0 624 0 1 2276
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5147_6
timestamp 1731220637
transform 1 0 640 0 -1 2268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5146_6
timestamp 1731220637
transform 1 0 720 0 -1 2268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5145_6
timestamp 1731220637
transform 1 0 800 0 -1 2268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5144_6
timestamp 1731220637
transform 1 0 824 0 1 2132
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5143_6
timestamp 1731220637
transform 1 0 752 0 1 2132
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5142_6
timestamp 1731220637
transform 1 0 672 0 1 2132
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5141_6
timestamp 1731220637
transform 1 0 728 0 -1 2124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5140_6
timestamp 1731220637
transform 1 0 784 0 -1 2124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5139_6
timestamp 1731220637
transform 1 0 832 0 -1 2124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5138_6
timestamp 1731220637
transform 1 0 880 0 -1 2124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5137_6
timestamp 1731220637
transform 1 0 928 0 -1 2124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5136_6
timestamp 1731220637
transform 1 0 984 0 -1 2124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5135_6
timestamp 1731220637
transform 1 0 1040 0 -1 2124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5134_6
timestamp 1731220637
transform 1 0 896 0 1 2132
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5133_6
timestamp 1731220637
transform 1 0 968 0 1 2132
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5132_6
timestamp 1731220637
transform 1 0 1040 0 1 2132
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5131_6
timestamp 1731220637
transform 1 0 1112 0 1 2132
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5130_6
timestamp 1731220637
transform 1 0 1120 0 -1 2268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5129_6
timestamp 1731220637
transform 1 0 1040 0 -1 2268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5128_6
timestamp 1731220637
transform 1 0 880 0 -1 2268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5127_6
timestamp 1731220637
transform 1 0 960 0 -1 2268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5126_6
timestamp 1731220637
transform 1 0 984 0 1 2276
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5125_6
timestamp 1731220637
transform 1 0 1056 0 1 2276
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5124_6
timestamp 1731220637
transform 1 0 912 0 1 2276
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5123_6
timestamp 1731220637
transform 1 0 776 0 1 2276
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5122_6
timestamp 1731220637
transform 1 0 848 0 1 2276
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5121_6
timestamp 1731220637
transform 1 0 888 0 -1 2416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5120_6
timestamp 1731220637
transform 1 0 960 0 -1 2416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5119_6
timestamp 1731220637
transform 1 0 816 0 -1 2416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5118_6
timestamp 1731220637
transform 1 0 744 0 -1 2416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5117_6
timestamp 1731220637
transform 1 0 696 0 1 2424
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5116_6
timestamp 1731220637
transform 1 0 760 0 1 2424
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5115_6
timestamp 1731220637
transform 1 0 816 0 1 2424
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5114_6
timestamp 1731220637
transform 1 0 872 0 1 2424
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5113_6
timestamp 1731220637
transform 1 0 920 0 1 2424
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5112_6
timestamp 1731220637
transform 1 0 968 0 1 2424
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5111_6
timestamp 1731220637
transform 1 0 1016 0 1 2424
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5110_6
timestamp 1731220637
transform 1 0 1064 0 1 2424
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5109_6
timestamp 1731220637
transform 1 0 1104 0 1 2424
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5108_6
timestamp 1731220637
transform 1 0 1144 0 1 2424
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5107_6
timestamp 1731220637
transform 1 0 1184 0 1 2424
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5106_6
timestamp 1731220637
transform 1 0 1296 0 1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5105_6
timestamp 1731220637
transform 1 0 1336 0 1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5104_6
timestamp 1731220637
transform 1 0 1376 0 1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5103_6
timestamp 1731220637
transform 1 0 1432 0 1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5102_6
timestamp 1731220637
transform 1 0 1504 0 1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5101_6
timestamp 1731220637
transform 1 0 1576 0 1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5100_6
timestamp 1731220637
transform 1 0 1656 0 1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_599_6
timestamp 1731220637
transform 1 0 1368 0 -1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_598_6
timestamp 1731220637
transform 1 0 1408 0 -1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_597_6
timestamp 1731220637
transform 1 0 1448 0 -1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_596_6
timestamp 1731220637
transform 1 0 1496 0 -1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_595_6
timestamp 1731220637
transform 1 0 1552 0 -1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_594_6
timestamp 1731220637
transform 1 0 1608 0 -1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_593_6
timestamp 1731220637
transform 1 0 1672 0 -1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_592_6
timestamp 1731220637
transform 1 0 1568 0 1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_591_6
timestamp 1731220637
transform 1 0 1496 0 1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_590_6
timestamp 1731220637
transform 1 0 1432 0 1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_589_6
timestamp 1731220637
transform 1 0 1376 0 1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_588_6
timestamp 1731220637
transform 1 0 1320 0 1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_587_6
timestamp 1731220637
transform 1 0 1328 0 -1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_586_6
timestamp 1731220637
transform 1 0 1400 0 -1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_585_6
timestamp 1731220637
transform 1 0 1480 0 -1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_584_6
timestamp 1731220637
transform 1 0 1504 0 1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_583_6
timestamp 1731220637
transform 1 0 1432 0 1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_582_6
timestamp 1731220637
transform 1 0 1368 0 1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_581_6
timestamp 1731220637
transform 1 0 1392 0 -1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_580_6
timestamp 1731220637
transform 1 0 1432 0 -1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_579_6
timestamp 1731220637
transform 1 0 1488 0 -1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_578_6
timestamp 1731220637
transform 1 0 1560 0 -1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_577_6
timestamp 1731220637
transform 1 0 1640 0 -1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_576_6
timestamp 1731220637
transform 1 0 1728 0 -1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_575_6
timestamp 1731220637
transform 1 0 1816 0 -1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_574_6
timestamp 1731220637
transform 1 0 1744 0 1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_573_6
timestamp 1731220637
transform 1 0 1664 0 1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_572_6
timestamp 1731220637
transform 1 0 1584 0 1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_571_6
timestamp 1731220637
transform 1 0 1552 0 -1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_570_6
timestamp 1731220637
transform 1 0 1624 0 -1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_569_6
timestamp 1731220637
transform 1 0 1696 0 -1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_568_6
timestamp 1731220637
transform 1 0 1768 0 -1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_567_6
timestamp 1731220637
transform 1 0 1640 0 1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_566_6
timestamp 1731220637
transform 1 0 1712 0 1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_565_6
timestamp 1731220637
transform 1 0 1792 0 1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_564_6
timestamp 1731220637
transform 1 0 1872 0 1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_563_6
timestamp 1731220637
transform 1 0 1728 0 -1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_562_6
timestamp 1731220637
transform 1 0 1792 0 -1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_561_6
timestamp 1731220637
transform 1 0 1864 0 -1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_560_6
timestamp 1731220637
transform 1 0 1944 0 -1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_559_6
timestamp 1731220637
transform 1 0 1728 0 1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_558_6
timestamp 1731220637
transform 1 0 1800 0 1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_557_6
timestamp 1731220637
transform 1 0 1880 0 1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_556_6
timestamp 1731220637
transform 1 0 1960 0 1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_555_6
timestamp 1731220637
transform 1 0 2056 0 1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_554_6
timestamp 1731220637
transform 1 0 2160 0 1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_553_6
timestamp 1731220637
transform 1 0 2264 0 1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_552_6
timestamp 1731220637
transform 1 0 2256 0 -1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_551_6
timestamp 1731220637
transform 1 0 2040 0 -1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_550_6
timestamp 1731220637
transform 1 0 2144 0 -1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_549_6
timestamp 1731220637
transform 1 0 2160 0 1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_548_6
timestamp 1731220637
transform 1 0 2056 0 1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_547_6
timestamp 1731220637
transform 1 0 1960 0 1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_546_6
timestamp 1731220637
transform 1 0 1832 0 -1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_545_6
timestamp 1731220637
transform 1 0 1904 0 -1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_544_6
timestamp 1731220637
transform 1 0 1984 0 -1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_543_6
timestamp 1731220637
transform 1 0 2072 0 -1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_542_6
timestamp 1731220637
transform 1 0 2168 0 -1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_541_6
timestamp 1731220637
transform 1 0 2272 0 -1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_540_6
timestamp 1731220637
transform 1 0 1824 0 1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_539_6
timestamp 1731220637
transform 1 0 1896 0 1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_538_6
timestamp 1731220637
transform 1 0 1960 0 1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_537_6
timestamp 1731220637
transform 1 0 2024 0 1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_536_6
timestamp 1731220637
transform 1 0 2088 0 1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_535_6
timestamp 1731220637
transform 1 0 2160 0 1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_534_6
timestamp 1731220637
transform 1 0 2232 0 1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_533_6
timestamp 1731220637
transform 1 0 1904 0 -1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_532_6
timestamp 1731220637
transform 1 0 1992 0 -1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_531_6
timestamp 1731220637
transform 1 0 2080 0 -1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_530_6
timestamp 1731220637
transform 1 0 2168 0 -1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_529_6
timestamp 1731220637
transform 1 0 2264 0 -1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_528_6
timestamp 1731220637
transform 1 0 2072 0 1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_527_6
timestamp 1731220637
transform 1 0 2032 0 1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_526_6
timestamp 1731220637
transform 1 0 1912 0 -1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_525_6
timestamp 1731220637
transform 1 0 1960 0 -1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_524_6
timestamp 1731220637
transform 1 0 2008 0 -1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_523_6
timestamp 1731220637
transform 1 0 2144 0 1 1860
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_522_6
timestamp 1731220637
transform 1 0 2048 0 -1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_521_6
timestamp 1731220637
transform 1 0 2088 0 -1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_520_6
timestamp 1731220637
transform 1 0 2136 0 -1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_519_6
timestamp 1731220637
transform 1 0 2184 0 -1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_518_6
timestamp 1731220637
transform 1 0 2112 0 1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_517_6
timestamp 1731220637
transform 1 0 2152 0 1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_516_6
timestamp 1731220637
transform 1 0 2192 0 1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_515_6
timestamp 1731220637
transform 1 0 2232 0 1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_514_6
timestamp 1731220637
transform 1 0 2272 0 1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_513_6
timestamp 1731220637
transform 1 0 2232 0 -1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_512_6
timestamp 1731220637
transform 1 0 2272 0 -1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_511_6
timestamp 1731220637
transform 1 0 2312 0 -1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_510_6
timestamp 1731220637
transform 1 0 2352 0 -1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_59_6
timestamp 1731220637
transform 1 0 2352 0 1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_58_6
timestamp 1731220637
transform 1 0 2312 0 1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_57_6
timestamp 1731220637
transform 1 0 2352 0 -1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_56_6
timestamp 1731220637
transform 1 0 2304 0 1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_55_6
timestamp 1731220637
transform 1 0 2352 0 1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_54_6
timestamp 1731220637
transform 1 0 2352 0 -1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_53_6
timestamp 1731220637
transform 1 0 2264 0 1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_52_6
timestamp 1731220637
transform 1 0 2352 0 1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_51_6
timestamp 1731220637
transform 1 0 2352 0 -1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_50_6
timestamp 1731220637
transform 1 0 2352 0 1 2420
box 4 6 36 64
<< end >>
