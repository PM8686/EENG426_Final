magic
tech sky130l
timestamp 1730593976
<< m1 >>
rect 368 763 372 795
rect 472 651 476 683
rect 680 539 684 563
rect 288 483 292 515
rect 384 303 388 327
rect 448 207 452 271
rect 232 175 236 199
rect 496 175 500 199
rect 568 111 572 155
<< m2c >>
rect 138 851 142 855
rect 186 851 190 855
rect 111 841 115 845
rect 775 841 779 845
rect 111 823 115 827
rect 775 823 779 827
rect 368 795 372 799
rect 111 781 115 785
rect 111 763 115 767
rect 775 781 779 785
rect 775 763 779 767
rect 368 759 372 763
rect 139 751 143 755
rect 184 751 188 755
rect 232 751 236 755
rect 280 751 284 755
rect 328 751 332 755
rect 376 751 380 755
rect 274 743 278 747
rect 322 739 326 743
rect 370 739 374 743
rect 426 739 430 743
rect 490 739 494 743
rect 562 739 566 743
rect 642 739 646 743
rect 722 739 726 743
rect 111 729 115 733
rect 775 729 779 733
rect 111 711 115 715
rect 775 711 779 715
rect 472 683 476 687
rect 111 669 115 673
rect 111 651 115 655
rect 775 669 779 673
rect 775 651 779 655
rect 472 647 476 651
rect 336 639 340 643
rect 384 639 388 643
rect 432 639 436 643
rect 480 639 484 643
rect 531 639 535 643
rect 576 639 580 643
rect 624 639 628 643
rect 675 639 679 643
rect 720 639 724 643
rect 482 631 486 635
rect 722 631 726 635
rect 138 627 142 631
rect 186 627 190 631
rect 258 627 262 631
rect 362 627 366 631
rect 610 627 614 631
rect 111 617 115 621
rect 775 617 779 621
rect 111 599 115 603
rect 775 599 779 603
rect 680 563 684 567
rect 111 557 115 561
rect 111 539 115 543
rect 775 557 779 561
rect 775 539 779 543
rect 680 535 684 539
rect 139 527 143 531
rect 184 527 188 531
rect 264 527 268 531
rect 352 527 356 531
rect 448 527 452 531
rect 544 527 548 531
rect 640 527 644 531
rect 723 527 727 531
rect 194 519 198 523
rect 722 519 726 523
rect 250 515 254 519
rect 288 515 292 519
rect 314 515 318 519
rect 386 515 390 519
rect 466 515 470 519
rect 554 515 558 519
rect 650 515 654 519
rect 111 505 115 509
rect 111 487 115 491
rect 775 505 779 509
rect 775 487 779 491
rect 288 479 292 483
rect 111 445 115 449
rect 775 445 779 449
rect 111 427 115 431
rect 775 427 779 431
rect 352 415 356 419
rect 400 415 404 419
rect 448 415 452 419
rect 496 415 500 419
rect 544 415 548 419
rect 600 415 604 419
rect 664 415 668 419
rect 723 415 727 419
rect 586 403 590 407
rect 722 403 726 407
rect 322 399 326 403
rect 370 399 374 403
rect 418 399 422 403
rect 466 399 470 403
rect 522 399 526 403
rect 650 399 654 403
rect 111 389 115 393
rect 775 389 779 393
rect 111 371 115 375
rect 775 371 779 375
rect 384 327 388 331
rect 111 321 115 325
rect 111 303 115 307
rect 775 321 779 325
rect 775 303 779 307
rect 384 299 388 303
rect 136 291 140 295
rect 200 291 204 295
rect 272 291 276 295
rect 344 291 348 295
rect 427 291 431 295
rect 512 291 516 295
rect 608 291 612 295
rect 707 291 711 295
rect 138 275 142 279
rect 722 275 726 279
rect 194 271 198 275
rect 282 271 286 275
rect 370 271 374 275
rect 448 271 452 275
rect 458 271 462 275
rect 546 271 550 275
rect 642 271 646 275
rect 111 261 115 265
rect 111 243 115 247
rect 775 261 779 265
rect 775 243 779 247
rect 448 203 452 207
rect 232 199 236 203
rect 111 193 115 197
rect 111 175 115 179
rect 232 171 236 175
rect 496 199 500 203
rect 775 193 779 197
rect 775 175 779 179
rect 496 171 500 175
rect 192 163 196 167
rect 280 163 284 167
rect 371 163 375 167
rect 456 163 460 167
rect 552 163 556 167
rect 651 163 655 167
rect 720 163 724 167
rect 568 155 572 159
rect 194 147 198 151
rect 242 143 246 147
rect 290 143 294 147
rect 338 143 342 147
rect 386 143 390 147
rect 434 143 438 147
rect 482 143 486 147
rect 530 143 534 147
rect 111 133 115 137
rect 111 115 115 119
rect 722 147 726 151
rect 578 143 582 147
rect 626 143 630 147
rect 674 143 678 147
rect 775 133 779 137
rect 775 115 779 119
rect 568 107 572 111
<< m2 >>
rect 154 857 160 858
rect 137 855 143 856
rect 137 851 138 855
rect 142 854 143 855
rect 142 852 150 854
rect 154 853 155 857
rect 159 853 160 857
rect 202 857 208 858
rect 154 852 160 853
rect 185 855 191 856
rect 142 851 143 852
rect 137 850 143 851
rect 148 850 150 852
rect 174 851 180 852
rect 174 850 175 851
rect 148 848 175 850
rect 174 847 175 848
rect 179 847 180 851
rect 185 851 186 855
rect 190 854 191 855
rect 190 852 198 854
rect 202 853 203 857
rect 207 853 208 857
rect 202 852 208 853
rect 250 857 256 858
rect 250 853 251 857
rect 255 853 256 857
rect 250 852 256 853
rect 190 851 191 852
rect 185 850 191 851
rect 196 850 198 852
rect 222 851 228 852
rect 222 850 223 851
rect 196 848 223 850
rect 174 846 180 847
rect 222 847 223 848
rect 227 847 228 851
rect 222 846 228 847
rect 110 845 116 846
rect 110 841 111 845
rect 115 841 116 845
rect 110 840 116 841
rect 774 845 780 846
rect 774 841 775 845
rect 779 841 780 845
rect 774 840 780 841
rect 110 827 116 828
rect 110 823 111 827
rect 115 823 116 827
rect 110 822 116 823
rect 134 827 140 828
rect 134 823 135 827
rect 139 823 140 827
rect 134 822 140 823
rect 182 827 188 828
rect 182 823 183 827
rect 187 823 188 827
rect 182 822 188 823
rect 230 827 236 828
rect 230 823 231 827
rect 235 823 236 827
rect 230 822 236 823
rect 774 827 780 828
rect 774 823 775 827
rect 779 823 780 827
rect 774 822 780 823
rect 142 819 148 820
rect 142 815 143 819
rect 147 815 148 819
rect 142 814 148 815
rect 174 819 180 820
rect 174 815 175 819
rect 179 818 180 819
rect 222 819 228 820
rect 179 816 185 818
rect 179 815 180 816
rect 174 814 180 815
rect 222 815 223 819
rect 227 818 228 819
rect 227 816 233 818
rect 227 815 228 816
rect 222 814 228 815
rect 367 799 373 800
rect 367 795 368 799
rect 372 798 373 799
rect 372 796 378 798
rect 372 795 373 796
rect 367 794 373 795
rect 376 793 378 796
rect 174 791 180 792
rect 174 790 175 791
rect 169 788 175 790
rect 174 787 175 788
rect 179 787 180 791
rect 222 791 228 792
rect 222 790 223 791
rect 217 788 223 790
rect 174 786 180 787
rect 222 787 223 788
rect 227 787 228 791
rect 270 791 276 792
rect 270 790 271 791
rect 265 788 271 790
rect 222 786 228 787
rect 270 787 271 788
rect 275 787 276 791
rect 318 791 324 792
rect 318 790 319 791
rect 313 788 319 790
rect 270 786 276 787
rect 318 787 319 788
rect 323 787 324 791
rect 366 791 372 792
rect 366 790 367 791
rect 361 788 367 790
rect 318 786 324 787
rect 366 787 367 788
rect 371 787 372 791
rect 366 786 372 787
rect 110 785 116 786
rect 110 781 111 785
rect 115 781 116 785
rect 110 780 116 781
rect 134 785 140 786
rect 134 781 135 785
rect 139 781 140 785
rect 134 780 140 781
rect 182 785 188 786
rect 182 781 183 785
rect 187 781 188 785
rect 182 780 188 781
rect 230 785 236 786
rect 230 781 231 785
rect 235 781 236 785
rect 230 780 236 781
rect 278 785 284 786
rect 278 781 279 785
rect 283 781 284 785
rect 278 780 284 781
rect 326 785 332 786
rect 326 781 327 785
rect 331 781 332 785
rect 326 780 332 781
rect 374 785 380 786
rect 374 781 375 785
rect 379 781 380 785
rect 374 780 380 781
rect 774 785 780 786
rect 774 781 775 785
rect 779 781 780 785
rect 774 780 780 781
rect 110 767 116 768
rect 110 763 111 767
rect 115 763 116 767
rect 774 767 780 768
rect 110 762 116 763
rect 278 763 284 764
rect 278 759 279 763
rect 283 762 284 763
rect 367 763 373 764
rect 367 762 368 763
rect 283 760 368 762
rect 283 759 284 760
rect 278 758 284 759
rect 367 759 368 760
rect 372 759 373 763
rect 774 763 775 767
rect 779 763 780 767
rect 774 762 780 763
rect 367 758 373 759
rect 138 755 148 756
rect 138 751 139 755
rect 147 751 148 755
rect 138 750 148 751
rect 154 755 160 756
rect 154 751 155 755
rect 159 751 160 755
rect 154 750 160 751
rect 174 755 180 756
rect 174 751 175 755
rect 179 754 180 755
rect 183 755 189 756
rect 183 754 184 755
rect 179 752 184 754
rect 179 751 180 752
rect 174 750 180 751
rect 183 751 184 752
rect 188 751 189 755
rect 183 750 189 751
rect 202 755 208 756
rect 202 751 203 755
rect 207 751 208 755
rect 202 750 208 751
rect 222 755 228 756
rect 222 751 223 755
rect 227 754 228 755
rect 231 755 237 756
rect 231 754 232 755
rect 227 752 232 754
rect 227 751 228 752
rect 222 750 228 751
rect 231 751 232 752
rect 236 751 237 755
rect 231 750 237 751
rect 250 755 256 756
rect 250 751 251 755
rect 255 751 256 755
rect 250 750 256 751
rect 270 755 276 756
rect 270 751 271 755
rect 275 754 276 755
rect 279 755 285 756
rect 279 754 280 755
rect 275 752 280 754
rect 275 751 276 752
rect 270 750 276 751
rect 279 751 280 752
rect 284 751 285 755
rect 279 750 285 751
rect 298 755 304 756
rect 298 751 299 755
rect 303 751 304 755
rect 298 750 304 751
rect 318 755 324 756
rect 318 751 319 755
rect 323 754 324 755
rect 327 755 333 756
rect 327 754 328 755
rect 323 752 328 754
rect 323 751 324 752
rect 318 750 324 751
rect 327 751 328 752
rect 332 751 333 755
rect 327 750 333 751
rect 346 755 352 756
rect 346 751 347 755
rect 351 751 352 755
rect 346 750 352 751
rect 366 755 372 756
rect 366 751 367 755
rect 371 754 372 755
rect 375 755 381 756
rect 375 754 376 755
rect 371 752 376 754
rect 371 751 372 752
rect 366 750 372 751
rect 375 751 376 752
rect 380 751 381 755
rect 375 750 381 751
rect 394 755 400 756
rect 394 751 395 755
rect 399 751 400 755
rect 394 750 400 751
rect 273 747 284 748
rect 273 743 274 747
rect 278 743 279 747
rect 283 743 284 747
rect 273 742 284 743
rect 290 745 296 746
rect 290 741 291 745
rect 295 741 296 745
rect 338 745 344 746
rect 290 740 296 741
rect 310 743 316 744
rect 310 739 311 743
rect 315 742 316 743
rect 321 743 327 744
rect 321 742 322 743
rect 315 740 322 742
rect 315 739 316 740
rect 310 738 316 739
rect 321 739 322 740
rect 326 739 327 743
rect 338 741 339 745
rect 343 741 344 745
rect 386 745 392 746
rect 338 740 344 741
rect 358 743 364 744
rect 321 738 327 739
rect 358 739 359 743
rect 363 742 364 743
rect 369 743 375 744
rect 369 742 370 743
rect 363 740 370 742
rect 363 739 364 740
rect 358 738 364 739
rect 369 739 370 740
rect 374 739 375 743
rect 386 741 387 745
rect 391 741 392 745
rect 442 745 448 746
rect 386 740 392 741
rect 406 743 412 744
rect 369 738 375 739
rect 406 739 407 743
rect 411 742 412 743
rect 425 743 431 744
rect 425 742 426 743
rect 411 740 426 742
rect 411 739 412 740
rect 406 738 412 739
rect 425 739 426 740
rect 430 739 431 743
rect 442 741 443 745
rect 447 741 448 745
rect 506 745 512 746
rect 442 740 448 741
rect 454 743 460 744
rect 425 738 431 739
rect 454 739 455 743
rect 459 742 460 743
rect 489 743 495 744
rect 489 742 490 743
rect 459 740 490 742
rect 459 739 460 740
rect 454 738 460 739
rect 489 739 490 740
rect 494 739 495 743
rect 506 741 507 745
rect 511 741 512 745
rect 578 745 584 746
rect 506 740 512 741
rect 518 743 524 744
rect 489 738 495 739
rect 518 739 519 743
rect 523 742 524 743
rect 561 743 567 744
rect 561 742 562 743
rect 523 740 562 742
rect 523 739 524 740
rect 518 738 524 739
rect 561 739 562 740
rect 566 739 567 743
rect 578 741 579 745
rect 583 741 584 745
rect 658 745 664 746
rect 578 740 584 741
rect 641 743 652 744
rect 561 738 567 739
rect 641 739 642 743
rect 646 739 647 743
rect 651 739 652 743
rect 658 741 659 745
rect 663 741 664 745
rect 738 745 744 746
rect 658 740 664 741
rect 670 743 676 744
rect 641 738 652 739
rect 670 739 671 743
rect 675 742 676 743
rect 721 743 727 744
rect 721 742 722 743
rect 675 740 722 742
rect 675 739 676 740
rect 670 738 676 739
rect 721 739 722 740
rect 726 739 727 743
rect 738 741 739 745
rect 743 741 744 745
rect 738 740 744 741
rect 721 738 727 739
rect 110 733 116 734
rect 110 729 111 733
rect 115 729 116 733
rect 110 728 116 729
rect 774 733 780 734
rect 774 729 775 733
rect 779 729 780 733
rect 774 728 780 729
rect 110 715 116 716
rect 110 711 111 715
rect 115 711 116 715
rect 110 710 116 711
rect 270 715 276 716
rect 270 711 271 715
rect 275 711 276 715
rect 270 710 276 711
rect 318 715 324 716
rect 318 711 319 715
rect 323 711 324 715
rect 318 710 324 711
rect 366 715 372 716
rect 366 711 367 715
rect 371 711 372 715
rect 366 710 372 711
rect 422 715 428 716
rect 422 711 423 715
rect 427 711 428 715
rect 422 710 428 711
rect 486 715 492 716
rect 486 711 487 715
rect 491 711 492 715
rect 486 710 492 711
rect 558 715 564 716
rect 558 711 559 715
rect 563 711 564 715
rect 558 710 564 711
rect 638 715 644 716
rect 638 711 639 715
rect 643 711 644 715
rect 638 710 644 711
rect 718 715 724 716
rect 718 711 719 715
rect 723 711 724 715
rect 718 710 724 711
rect 774 715 780 716
rect 774 711 775 715
rect 779 711 780 715
rect 774 710 780 711
rect 310 707 316 708
rect 310 706 311 707
rect 305 704 311 706
rect 310 703 311 704
rect 315 703 316 707
rect 358 707 364 708
rect 358 706 359 707
rect 353 704 359 706
rect 310 702 316 703
rect 358 703 359 704
rect 363 703 364 707
rect 406 707 412 708
rect 406 706 407 707
rect 401 704 407 706
rect 358 702 364 703
rect 406 703 407 704
rect 411 703 412 707
rect 406 702 412 703
rect 454 707 460 708
rect 454 703 455 707
rect 459 703 460 707
rect 454 702 460 703
rect 518 707 524 708
rect 518 703 519 707
rect 523 703 524 707
rect 518 702 524 703
rect 534 707 540 708
rect 534 703 535 707
rect 539 706 540 707
rect 670 707 676 708
rect 539 704 561 706
rect 539 703 540 704
rect 534 702 540 703
rect 670 703 671 707
rect 675 703 676 707
rect 670 702 676 703
rect 678 707 684 708
rect 678 703 679 707
rect 683 706 684 707
rect 683 704 721 706
rect 683 703 684 704
rect 678 702 684 703
rect 471 687 477 688
rect 366 683 372 684
rect 366 679 367 683
rect 371 679 372 683
rect 471 683 472 687
rect 476 686 477 687
rect 476 684 482 686
rect 476 683 477 684
rect 471 682 477 683
rect 480 681 482 684
rect 654 683 660 684
rect 366 678 372 679
rect 422 679 428 680
rect 422 678 423 679
rect 417 676 423 678
rect 422 675 423 676
rect 427 675 428 679
rect 470 679 476 680
rect 470 678 471 679
rect 465 676 471 678
rect 422 674 428 675
rect 470 675 471 676
rect 475 675 476 679
rect 470 674 476 675
rect 518 679 524 680
rect 518 675 519 679
rect 523 678 524 679
rect 614 679 620 680
rect 614 678 615 679
rect 523 676 529 678
rect 609 676 615 678
rect 523 675 524 676
rect 518 674 524 675
rect 614 675 615 676
rect 619 675 620 679
rect 654 679 655 683
rect 659 679 660 683
rect 654 678 660 679
rect 702 683 708 684
rect 702 679 703 683
rect 707 679 708 683
rect 702 678 708 679
rect 710 679 716 680
rect 614 674 620 675
rect 710 675 711 679
rect 715 678 716 679
rect 715 676 721 678
rect 715 675 716 676
rect 710 674 716 675
rect 110 673 116 674
rect 110 669 111 673
rect 115 669 116 673
rect 110 668 116 669
rect 334 673 340 674
rect 334 669 335 673
rect 339 669 340 673
rect 334 668 340 669
rect 382 673 388 674
rect 382 669 383 673
rect 387 669 388 673
rect 382 668 388 669
rect 430 673 436 674
rect 430 669 431 673
rect 435 669 436 673
rect 430 668 436 669
rect 478 673 484 674
rect 478 669 479 673
rect 483 669 484 673
rect 478 668 484 669
rect 526 673 532 674
rect 526 669 527 673
rect 531 669 532 673
rect 526 668 532 669
rect 574 673 580 674
rect 574 669 575 673
rect 579 669 580 673
rect 574 668 580 669
rect 622 673 628 674
rect 622 669 623 673
rect 627 669 628 673
rect 622 668 628 669
rect 670 673 676 674
rect 670 669 671 673
rect 675 669 676 673
rect 670 668 676 669
rect 718 673 724 674
rect 718 669 719 673
rect 723 669 724 673
rect 718 668 724 669
rect 774 673 780 674
rect 774 669 775 673
rect 779 669 780 673
rect 774 668 780 669
rect 110 655 116 656
rect 110 651 111 655
rect 115 651 116 655
rect 774 655 780 656
rect 110 650 116 651
rect 471 651 477 652
rect 471 650 472 651
rect 348 648 472 650
rect 335 643 341 644
rect 335 639 336 643
rect 340 642 341 643
rect 348 642 350 648
rect 471 647 472 648
rect 476 647 477 651
rect 518 651 524 652
rect 518 650 519 651
rect 471 646 477 647
rect 484 648 519 650
rect 484 644 486 648
rect 518 647 519 648
rect 523 647 524 651
rect 774 651 775 655
rect 779 651 780 655
rect 774 650 780 651
rect 518 646 524 647
rect 340 640 350 642
rect 354 643 360 644
rect 340 639 341 640
rect 335 638 341 639
rect 354 639 355 643
rect 359 639 360 643
rect 354 638 360 639
rect 366 643 372 644
rect 366 639 367 643
rect 371 642 372 643
rect 383 643 389 644
rect 383 642 384 643
rect 371 640 384 642
rect 371 639 372 640
rect 366 638 372 639
rect 383 639 384 640
rect 388 639 389 643
rect 383 638 389 639
rect 402 643 408 644
rect 402 639 403 643
rect 407 639 408 643
rect 402 638 408 639
rect 422 643 428 644
rect 422 639 423 643
rect 427 642 428 643
rect 431 643 437 644
rect 431 642 432 643
rect 427 640 432 642
rect 427 639 428 640
rect 422 638 428 639
rect 431 639 432 640
rect 436 639 437 643
rect 431 638 437 639
rect 450 643 456 644
rect 450 639 451 643
rect 455 639 456 643
rect 450 638 456 639
rect 479 643 486 644
rect 479 639 480 643
rect 484 640 486 643
rect 498 643 504 644
rect 484 639 485 640
rect 479 638 485 639
rect 498 639 499 643
rect 503 639 504 643
rect 498 638 504 639
rect 530 643 540 644
rect 530 639 531 643
rect 539 639 540 643
rect 530 638 540 639
rect 546 643 552 644
rect 546 639 547 643
rect 551 639 552 643
rect 546 638 552 639
rect 574 643 581 644
rect 574 639 575 643
rect 580 639 581 643
rect 574 638 581 639
rect 594 643 600 644
rect 594 639 595 643
rect 599 639 600 643
rect 594 638 600 639
rect 614 643 620 644
rect 614 639 615 643
rect 619 642 620 643
rect 623 643 629 644
rect 623 642 624 643
rect 619 640 624 642
rect 619 639 620 640
rect 614 638 620 639
rect 623 639 624 640
rect 628 639 629 643
rect 623 638 629 639
rect 642 643 648 644
rect 642 639 643 643
rect 647 639 648 643
rect 642 638 648 639
rect 674 643 684 644
rect 674 639 675 643
rect 683 639 684 643
rect 674 638 684 639
rect 690 643 696 644
rect 690 639 691 643
rect 695 639 696 643
rect 690 638 696 639
rect 702 643 708 644
rect 702 639 703 643
rect 707 642 708 643
rect 719 643 725 644
rect 719 642 720 643
rect 707 640 720 642
rect 707 639 708 640
rect 702 638 708 639
rect 719 639 720 640
rect 724 639 725 643
rect 719 638 725 639
rect 738 643 744 644
rect 738 639 739 643
rect 743 639 744 643
rect 738 638 744 639
rect 470 635 476 636
rect 154 633 160 634
rect 137 631 143 632
rect 137 627 138 631
rect 142 630 143 631
rect 142 628 150 630
rect 154 629 155 633
rect 159 629 160 633
rect 202 633 208 634
rect 154 628 160 629
rect 185 631 191 632
rect 142 627 143 628
rect 137 626 143 627
rect 148 626 150 628
rect 174 627 180 628
rect 174 626 175 627
rect 148 624 175 626
rect 174 623 175 624
rect 179 623 180 627
rect 185 627 186 631
rect 190 630 191 631
rect 190 628 198 630
rect 202 629 203 633
rect 207 629 208 633
rect 274 633 280 634
rect 202 628 208 629
rect 257 631 263 632
rect 190 627 191 628
rect 185 626 191 627
rect 196 626 198 628
rect 222 627 228 628
rect 222 626 223 627
rect 196 624 223 626
rect 174 622 180 623
rect 222 623 223 624
rect 227 623 228 627
rect 257 627 258 631
rect 262 630 263 631
rect 262 628 270 630
rect 274 629 275 633
rect 279 629 280 633
rect 378 633 384 634
rect 274 628 280 629
rect 361 631 367 632
rect 262 627 263 628
rect 257 626 263 627
rect 268 626 270 628
rect 310 627 316 628
rect 310 626 311 627
rect 268 624 311 626
rect 222 622 228 623
rect 310 623 311 624
rect 315 623 316 627
rect 361 627 362 631
rect 366 630 367 631
rect 366 628 374 630
rect 378 629 379 633
rect 383 629 384 633
rect 470 631 471 635
rect 475 634 476 635
rect 481 635 487 636
rect 481 634 482 635
rect 475 632 482 634
rect 475 631 476 632
rect 470 630 476 631
rect 481 631 482 632
rect 486 631 487 635
rect 710 635 716 636
rect 481 630 487 631
rect 498 633 504 634
rect 378 628 384 629
rect 498 629 499 633
rect 503 629 504 633
rect 626 633 632 634
rect 498 628 504 629
rect 510 631 516 632
rect 366 627 367 628
rect 361 626 367 627
rect 310 622 316 623
rect 372 622 374 628
rect 510 627 511 631
rect 515 630 516 631
rect 609 631 615 632
rect 609 630 610 631
rect 515 628 610 630
rect 515 627 516 628
rect 510 626 516 627
rect 609 627 610 628
rect 614 627 615 631
rect 626 629 627 633
rect 631 629 632 633
rect 710 631 711 635
rect 715 634 716 635
rect 721 635 727 636
rect 721 634 722 635
rect 715 632 722 634
rect 715 631 716 632
rect 710 630 716 631
rect 721 631 722 632
rect 726 631 727 635
rect 721 630 727 631
rect 738 633 744 634
rect 626 628 632 629
rect 738 629 739 633
rect 743 629 744 633
rect 738 628 744 629
rect 609 626 615 627
rect 518 623 524 624
rect 518 622 519 623
rect 110 621 116 622
rect 110 617 111 621
rect 115 617 116 621
rect 372 620 519 622
rect 518 619 519 620
rect 523 619 524 623
rect 518 618 524 619
rect 774 621 780 622
rect 110 616 116 617
rect 774 617 775 621
rect 779 617 780 621
rect 774 616 780 617
rect 110 603 116 604
rect 110 599 111 603
rect 115 599 116 603
rect 110 598 116 599
rect 134 603 140 604
rect 134 599 135 603
rect 139 599 140 603
rect 134 598 140 599
rect 182 603 188 604
rect 182 599 183 603
rect 187 599 188 603
rect 182 598 188 599
rect 254 603 260 604
rect 254 599 255 603
rect 259 599 260 603
rect 254 598 260 599
rect 358 603 364 604
rect 358 599 359 603
rect 363 599 364 603
rect 358 598 364 599
rect 478 603 484 604
rect 478 599 479 603
rect 483 599 484 603
rect 478 598 484 599
rect 606 603 612 604
rect 606 599 607 603
rect 611 599 612 603
rect 606 598 612 599
rect 718 603 724 604
rect 718 599 719 603
rect 723 599 724 603
rect 718 598 724 599
rect 774 603 780 604
rect 774 599 775 603
rect 779 599 780 603
rect 774 598 780 599
rect 142 595 148 596
rect 142 591 143 595
rect 147 591 148 595
rect 142 590 148 591
rect 174 595 180 596
rect 174 591 175 595
rect 179 594 180 595
rect 222 595 228 596
rect 179 592 185 594
rect 179 591 180 592
rect 174 590 180 591
rect 222 591 223 595
rect 227 594 228 595
rect 310 595 316 596
rect 227 592 257 594
rect 227 591 228 592
rect 222 590 228 591
rect 310 591 311 595
rect 315 594 316 595
rect 510 595 516 596
rect 315 592 361 594
rect 315 591 316 592
rect 310 590 316 591
rect 510 591 511 595
rect 515 591 516 595
rect 510 590 516 591
rect 518 595 524 596
rect 518 591 519 595
rect 523 594 524 595
rect 726 595 732 596
rect 523 592 609 594
rect 523 591 524 592
rect 518 590 524 591
rect 726 591 727 595
rect 731 591 732 595
rect 726 590 732 591
rect 390 575 396 576
rect 390 571 391 575
rect 395 574 396 575
rect 395 572 450 574
rect 395 571 396 572
rect 390 570 396 571
rect 448 569 450 572
rect 574 571 580 572
rect 174 567 180 568
rect 174 566 175 567
rect 169 564 175 566
rect 174 563 175 564
rect 179 563 180 567
rect 222 567 228 568
rect 222 566 223 567
rect 217 564 223 566
rect 174 562 180 563
rect 222 563 223 564
rect 227 563 228 567
rect 342 567 348 568
rect 342 566 343 567
rect 297 564 343 566
rect 222 562 228 563
rect 342 563 343 564
rect 347 563 348 567
rect 438 567 444 568
rect 438 566 439 567
rect 385 564 439 566
rect 342 562 348 563
rect 438 563 439 564
rect 443 563 444 567
rect 574 567 575 571
rect 579 567 580 571
rect 574 566 580 567
rect 670 571 676 572
rect 670 567 671 571
rect 675 567 676 571
rect 670 566 676 567
rect 679 567 685 568
rect 438 562 444 563
rect 679 563 680 567
rect 684 566 685 567
rect 684 564 721 566
rect 684 563 685 564
rect 679 562 685 563
rect 110 561 116 562
rect 110 557 111 561
rect 115 557 116 561
rect 110 556 116 557
rect 134 561 140 562
rect 134 557 135 561
rect 139 557 140 561
rect 134 556 140 557
rect 182 561 188 562
rect 182 557 183 561
rect 187 557 188 561
rect 182 556 188 557
rect 262 561 268 562
rect 262 557 263 561
rect 267 557 268 561
rect 262 556 268 557
rect 350 561 356 562
rect 350 557 351 561
rect 355 557 356 561
rect 350 556 356 557
rect 446 561 452 562
rect 446 557 447 561
rect 451 557 452 561
rect 446 556 452 557
rect 542 561 548 562
rect 542 557 543 561
rect 547 557 548 561
rect 542 556 548 557
rect 638 561 644 562
rect 638 557 639 561
rect 643 557 644 561
rect 638 556 644 557
rect 718 561 724 562
rect 718 557 719 561
rect 723 557 724 561
rect 718 556 724 557
rect 774 561 780 562
rect 774 557 775 561
rect 779 557 780 561
rect 774 556 780 557
rect 110 543 116 544
rect 110 539 111 543
rect 115 539 116 543
rect 774 543 780 544
rect 110 538 116 539
rect 390 539 396 540
rect 390 538 391 539
rect 196 536 391 538
rect 138 531 148 532
rect 138 527 139 531
rect 147 527 148 531
rect 138 526 148 527
rect 154 531 160 532
rect 154 527 155 531
rect 159 527 160 531
rect 154 526 160 527
rect 174 531 180 532
rect 174 527 175 531
rect 179 530 180 531
rect 183 531 189 532
rect 183 530 184 531
rect 179 528 184 530
rect 179 527 180 528
rect 174 526 180 527
rect 183 527 184 528
rect 188 527 189 531
rect 183 526 189 527
rect 196 524 198 536
rect 390 535 391 536
rect 395 535 396 539
rect 590 539 596 540
rect 590 538 591 539
rect 390 534 396 535
rect 556 536 591 538
rect 202 531 208 532
rect 202 527 203 531
rect 207 527 208 531
rect 202 526 208 527
rect 222 531 228 532
rect 222 527 223 531
rect 227 530 228 531
rect 263 531 269 532
rect 263 530 264 531
rect 227 528 264 530
rect 227 527 228 528
rect 222 526 228 527
rect 263 527 264 528
rect 268 527 269 531
rect 263 526 269 527
rect 282 531 288 532
rect 282 527 283 531
rect 287 527 288 531
rect 282 526 288 527
rect 342 531 348 532
rect 342 527 343 531
rect 347 530 348 531
rect 351 531 357 532
rect 351 530 352 531
rect 347 528 352 530
rect 347 527 348 528
rect 342 526 348 527
rect 351 527 352 528
rect 356 527 357 531
rect 351 526 357 527
rect 370 531 376 532
rect 370 527 371 531
rect 375 527 376 531
rect 370 526 376 527
rect 438 531 444 532
rect 438 527 439 531
rect 443 530 444 531
rect 447 531 453 532
rect 447 530 448 531
rect 443 528 448 530
rect 443 527 444 528
rect 438 526 444 527
rect 447 527 448 528
rect 452 527 453 531
rect 447 526 453 527
rect 466 531 472 532
rect 466 527 467 531
rect 471 527 472 531
rect 466 526 472 527
rect 543 531 549 532
rect 543 527 544 531
rect 548 530 549 531
rect 556 530 558 536
rect 590 535 591 536
rect 595 535 596 539
rect 679 539 685 540
rect 679 538 680 539
rect 590 534 596 535
rect 644 536 680 538
rect 644 532 646 536
rect 679 535 680 536
rect 684 535 685 539
rect 774 539 775 543
rect 779 539 780 543
rect 774 538 780 539
rect 679 534 685 535
rect 548 528 558 530
rect 562 531 568 532
rect 548 527 549 528
rect 543 526 549 527
rect 562 527 563 531
rect 567 527 568 531
rect 562 526 568 527
rect 639 531 646 532
rect 639 527 640 531
rect 644 528 646 531
rect 658 531 664 532
rect 644 527 645 528
rect 639 526 645 527
rect 658 527 659 531
rect 663 527 664 531
rect 658 526 664 527
rect 722 531 732 532
rect 722 527 723 531
rect 731 527 732 531
rect 722 526 732 527
rect 738 531 744 532
rect 738 527 739 531
rect 743 527 744 531
rect 738 526 744 527
rect 193 523 199 524
rect 193 519 194 523
rect 198 519 199 523
rect 674 523 680 524
rect 193 518 199 519
rect 210 521 216 522
rect 210 517 211 521
rect 215 517 216 521
rect 266 521 272 522
rect 210 516 216 517
rect 222 519 228 520
rect 222 515 223 519
rect 227 518 228 519
rect 249 519 255 520
rect 249 518 250 519
rect 227 516 250 518
rect 227 515 228 516
rect 222 514 228 515
rect 249 515 250 516
rect 254 515 255 519
rect 266 517 267 521
rect 271 517 272 521
rect 330 521 336 522
rect 266 516 272 517
rect 287 519 293 520
rect 249 514 255 515
rect 287 515 288 519
rect 292 518 293 519
rect 313 519 319 520
rect 313 518 314 519
rect 292 516 314 518
rect 292 515 293 516
rect 287 514 293 515
rect 313 515 314 516
rect 318 515 319 519
rect 330 517 331 521
rect 335 517 336 521
rect 402 521 408 522
rect 330 516 336 517
rect 342 519 348 520
rect 313 514 319 515
rect 342 515 343 519
rect 347 518 348 519
rect 385 519 391 520
rect 385 518 386 519
rect 347 516 386 518
rect 347 515 348 516
rect 342 514 348 515
rect 385 515 386 516
rect 390 515 391 519
rect 402 517 403 521
rect 407 517 408 521
rect 482 521 488 522
rect 402 516 408 517
rect 414 519 420 520
rect 385 514 391 515
rect 414 515 415 519
rect 419 518 420 519
rect 465 519 471 520
rect 465 518 466 519
rect 419 516 466 518
rect 419 515 420 516
rect 414 514 420 515
rect 465 515 466 516
rect 470 515 471 519
rect 482 517 483 521
rect 487 517 488 521
rect 570 521 576 522
rect 482 516 488 517
rect 494 519 500 520
rect 465 514 471 515
rect 494 515 495 519
rect 499 518 500 519
rect 553 519 559 520
rect 553 518 554 519
rect 499 516 554 518
rect 499 515 500 516
rect 494 514 500 515
rect 553 515 554 516
rect 558 515 559 519
rect 570 517 571 521
rect 575 517 576 521
rect 666 521 672 522
rect 570 516 576 517
rect 649 519 655 520
rect 553 514 559 515
rect 649 515 650 519
rect 654 518 655 519
rect 654 516 658 518
rect 666 517 667 521
rect 671 517 672 521
rect 674 519 675 523
rect 679 522 680 523
rect 721 523 727 524
rect 721 522 722 523
rect 679 520 722 522
rect 679 519 680 520
rect 674 518 680 519
rect 721 519 722 520
rect 726 519 727 523
rect 721 518 727 519
rect 738 521 744 522
rect 666 516 672 517
rect 738 517 739 521
rect 743 517 744 521
rect 738 516 744 517
rect 654 515 660 516
rect 649 514 655 515
rect 654 511 655 514
rect 659 511 660 515
rect 654 510 660 511
rect 110 509 116 510
rect 110 505 111 509
rect 115 505 116 509
rect 110 504 116 505
rect 774 509 780 510
rect 774 505 775 509
rect 779 505 780 509
rect 774 504 780 505
rect 110 491 116 492
rect 110 487 111 491
rect 115 487 116 491
rect 110 486 116 487
rect 190 491 196 492
rect 190 487 191 491
rect 195 487 196 491
rect 190 486 196 487
rect 246 491 252 492
rect 246 487 247 491
rect 251 487 252 491
rect 246 486 252 487
rect 310 491 316 492
rect 310 487 311 491
rect 315 487 316 491
rect 310 486 316 487
rect 382 491 388 492
rect 382 487 383 491
rect 387 487 388 491
rect 382 486 388 487
rect 462 491 468 492
rect 462 487 463 491
rect 467 487 468 491
rect 462 486 468 487
rect 550 491 556 492
rect 550 487 551 491
rect 555 487 556 491
rect 550 486 556 487
rect 646 491 652 492
rect 646 487 647 491
rect 651 487 652 491
rect 646 486 652 487
rect 718 491 724 492
rect 718 487 719 491
rect 723 487 724 491
rect 718 486 724 487
rect 774 491 780 492
rect 774 487 775 491
rect 779 487 780 491
rect 774 486 780 487
rect 222 483 228 484
rect 222 479 223 483
rect 227 479 228 483
rect 287 483 293 484
rect 287 482 288 483
rect 281 480 288 482
rect 222 478 228 479
rect 287 479 288 480
rect 292 479 293 483
rect 287 478 293 479
rect 342 483 348 484
rect 342 479 343 483
rect 347 479 348 483
rect 342 478 348 479
rect 414 483 420 484
rect 414 479 415 483
rect 419 479 420 483
rect 414 478 420 479
rect 494 483 500 484
rect 494 479 495 483
rect 499 479 500 483
rect 494 478 500 479
rect 502 483 508 484
rect 502 479 503 483
rect 507 482 508 483
rect 590 483 596 484
rect 507 480 553 482
rect 507 479 508 480
rect 502 478 508 479
rect 590 479 591 483
rect 595 482 596 483
rect 726 483 732 484
rect 595 480 649 482
rect 595 479 596 480
rect 590 478 596 479
rect 726 479 727 483
rect 731 479 732 483
rect 726 478 732 479
rect 574 459 580 460
rect 390 455 396 456
rect 390 454 391 455
rect 385 452 391 454
rect 390 451 391 452
rect 395 451 396 455
rect 438 455 444 456
rect 438 454 439 455
rect 433 452 439 454
rect 390 450 396 451
rect 438 451 439 452
rect 443 451 444 455
rect 486 455 492 456
rect 486 454 487 455
rect 481 452 487 454
rect 438 450 444 451
rect 486 451 487 452
rect 491 451 492 455
rect 534 455 540 456
rect 534 454 535 455
rect 529 452 535 454
rect 486 450 492 451
rect 534 451 535 452
rect 539 451 540 455
rect 574 455 575 459
rect 579 455 580 459
rect 654 459 660 460
rect 574 454 580 455
rect 586 455 592 456
rect 534 450 540 451
rect 586 451 587 455
rect 591 454 592 455
rect 654 455 655 459
rect 659 458 660 459
rect 659 456 665 458
rect 659 455 660 456
rect 654 454 660 455
rect 710 455 716 456
rect 591 452 601 454
rect 591 451 592 452
rect 586 450 592 451
rect 710 451 711 455
rect 715 454 716 455
rect 715 452 721 454
rect 715 451 716 452
rect 710 450 716 451
rect 110 449 116 450
rect 110 445 111 449
rect 115 445 116 449
rect 110 444 116 445
rect 350 449 356 450
rect 350 445 351 449
rect 355 445 356 449
rect 350 444 356 445
rect 398 449 404 450
rect 398 445 399 449
rect 403 445 404 449
rect 398 444 404 445
rect 446 449 452 450
rect 446 445 447 449
rect 451 445 452 449
rect 446 444 452 445
rect 494 449 500 450
rect 494 445 495 449
rect 499 445 500 449
rect 494 444 500 445
rect 542 449 548 450
rect 542 445 543 449
rect 547 445 548 449
rect 542 444 548 445
rect 598 449 604 450
rect 598 445 599 449
rect 603 445 604 449
rect 598 444 604 445
rect 662 449 668 450
rect 662 445 663 449
rect 667 445 668 449
rect 662 444 668 445
rect 718 449 724 450
rect 718 445 719 449
rect 723 445 724 449
rect 718 444 724 445
rect 774 449 780 450
rect 774 445 775 449
rect 779 445 780 449
rect 774 444 780 445
rect 110 431 116 432
rect 110 427 111 431
rect 115 427 116 431
rect 774 431 780 432
rect 110 426 116 427
rect 502 427 508 428
rect 502 426 503 427
rect 364 424 503 426
rect 351 419 357 420
rect 351 415 352 419
rect 356 418 357 419
rect 364 418 366 424
rect 502 423 503 424
rect 507 423 508 427
rect 774 427 775 431
rect 779 427 780 431
rect 774 426 780 427
rect 502 422 508 423
rect 356 416 366 418
rect 370 419 376 420
rect 356 415 357 416
rect 351 414 357 415
rect 370 415 371 419
rect 375 415 376 419
rect 370 414 376 415
rect 390 419 396 420
rect 390 415 391 419
rect 395 418 396 419
rect 399 419 405 420
rect 399 418 400 419
rect 395 416 400 418
rect 395 415 396 416
rect 390 414 396 415
rect 399 415 400 416
rect 404 415 405 419
rect 399 414 405 415
rect 418 419 424 420
rect 418 415 419 419
rect 423 415 424 419
rect 418 414 424 415
rect 438 419 444 420
rect 438 415 439 419
rect 443 418 444 419
rect 447 419 453 420
rect 447 418 448 419
rect 443 416 448 418
rect 443 415 444 416
rect 438 414 444 415
rect 447 415 448 416
rect 452 415 453 419
rect 447 414 453 415
rect 466 419 472 420
rect 466 415 467 419
rect 471 415 472 419
rect 466 414 472 415
rect 486 419 492 420
rect 486 415 487 419
rect 491 418 492 419
rect 495 419 501 420
rect 495 418 496 419
rect 491 416 496 418
rect 491 415 492 416
rect 486 414 492 415
rect 495 415 496 416
rect 500 415 501 419
rect 495 414 501 415
rect 514 419 520 420
rect 514 415 515 419
rect 519 415 520 419
rect 514 414 520 415
rect 534 419 540 420
rect 534 415 535 419
rect 539 418 540 419
rect 543 419 549 420
rect 543 418 544 419
rect 539 416 544 418
rect 539 415 540 416
rect 534 414 540 415
rect 543 415 544 416
rect 548 415 549 419
rect 543 414 549 415
rect 562 419 568 420
rect 562 415 563 419
rect 567 415 568 419
rect 562 414 568 415
rect 574 419 580 420
rect 574 415 575 419
rect 579 418 580 419
rect 599 419 605 420
rect 599 418 600 419
rect 579 416 600 418
rect 579 415 580 416
rect 574 414 580 415
rect 599 415 600 416
rect 604 415 605 419
rect 599 414 605 415
rect 618 419 624 420
rect 618 415 619 419
rect 623 415 624 419
rect 618 414 624 415
rect 658 419 669 420
rect 658 415 659 419
rect 663 415 664 419
rect 668 415 669 419
rect 658 414 669 415
rect 682 419 688 420
rect 682 415 683 419
rect 687 415 688 419
rect 682 414 688 415
rect 722 419 732 420
rect 722 415 723 419
rect 731 415 732 419
rect 722 414 732 415
rect 738 419 744 420
rect 738 415 739 419
rect 743 415 744 419
rect 738 414 744 415
rect 585 407 592 408
rect 338 405 344 406
rect 321 403 327 404
rect 321 399 322 403
rect 326 402 327 403
rect 326 400 334 402
rect 338 401 339 405
rect 343 401 344 405
rect 386 405 392 406
rect 338 400 344 401
rect 350 403 356 404
rect 326 399 327 400
rect 321 398 327 399
rect 332 394 334 400
rect 350 399 351 403
rect 355 402 356 403
rect 369 403 375 404
rect 369 402 370 403
rect 355 400 370 402
rect 355 399 356 400
rect 350 398 356 399
rect 369 399 370 400
rect 374 399 375 403
rect 386 401 387 405
rect 391 401 392 405
rect 434 405 440 406
rect 386 400 392 401
rect 398 403 404 404
rect 369 398 375 399
rect 398 399 399 403
rect 403 402 404 403
rect 417 403 423 404
rect 417 402 418 403
rect 403 400 418 402
rect 403 399 404 400
rect 398 398 404 399
rect 417 399 418 400
rect 422 399 423 403
rect 434 401 435 405
rect 439 401 440 405
rect 482 405 488 406
rect 434 400 440 401
rect 465 403 471 404
rect 417 398 423 399
rect 465 399 466 403
rect 470 402 471 403
rect 470 400 478 402
rect 482 401 483 405
rect 487 401 488 405
rect 538 405 544 406
rect 482 400 488 401
rect 521 403 527 404
rect 470 399 471 400
rect 465 398 471 399
rect 476 398 478 400
rect 502 399 508 400
rect 502 398 503 399
rect 476 396 503 398
rect 454 395 460 396
rect 454 394 455 395
rect 110 393 116 394
rect 110 389 111 393
rect 115 389 116 393
rect 332 392 455 394
rect 454 391 455 392
rect 459 391 460 395
rect 502 395 503 396
rect 507 395 508 399
rect 521 399 522 403
rect 526 402 527 403
rect 526 400 534 402
rect 538 401 539 405
rect 543 401 544 405
rect 585 403 586 407
rect 591 403 592 407
rect 710 407 716 408
rect 585 402 592 403
rect 602 405 608 406
rect 538 400 544 401
rect 602 401 603 405
rect 607 401 608 405
rect 666 405 672 406
rect 602 400 608 401
rect 638 403 644 404
rect 526 399 527 400
rect 521 398 527 399
rect 532 398 534 400
rect 558 399 564 400
rect 558 398 559 399
rect 532 396 559 398
rect 502 394 508 395
rect 558 395 559 396
rect 563 395 564 399
rect 638 399 639 403
rect 643 402 644 403
rect 649 403 655 404
rect 649 402 650 403
rect 643 400 650 402
rect 643 399 644 400
rect 638 398 644 399
rect 649 399 650 400
rect 654 399 655 403
rect 666 401 667 405
rect 671 401 672 405
rect 710 403 711 407
rect 715 406 716 407
rect 721 407 727 408
rect 721 406 722 407
rect 715 404 722 406
rect 715 403 716 404
rect 710 402 716 403
rect 721 403 722 404
rect 726 403 727 407
rect 721 402 727 403
rect 738 405 744 406
rect 666 400 672 401
rect 738 401 739 405
rect 743 401 744 405
rect 738 400 744 401
rect 649 398 655 399
rect 558 394 564 395
rect 454 390 460 391
rect 774 393 780 394
rect 110 388 116 389
rect 774 389 775 393
rect 779 389 780 393
rect 774 388 780 389
rect 110 375 116 376
rect 110 371 111 375
rect 115 371 116 375
rect 110 370 116 371
rect 318 375 324 376
rect 318 371 319 375
rect 323 371 324 375
rect 318 370 324 371
rect 366 375 372 376
rect 366 371 367 375
rect 371 371 372 375
rect 366 370 372 371
rect 414 375 420 376
rect 414 371 415 375
rect 419 371 420 375
rect 414 370 420 371
rect 462 375 468 376
rect 462 371 463 375
rect 467 371 468 375
rect 462 370 468 371
rect 518 375 524 376
rect 518 371 519 375
rect 523 371 524 375
rect 518 370 524 371
rect 582 375 588 376
rect 582 371 583 375
rect 587 371 588 375
rect 582 370 588 371
rect 646 375 652 376
rect 646 371 647 375
rect 651 371 652 375
rect 646 370 652 371
rect 718 375 724 376
rect 718 371 719 375
rect 723 371 724 375
rect 718 370 724 371
rect 774 375 780 376
rect 774 371 775 375
rect 779 371 780 375
rect 774 370 780 371
rect 350 367 356 368
rect 350 363 351 367
rect 355 363 356 367
rect 350 362 356 363
rect 398 367 404 368
rect 398 363 399 367
rect 403 363 404 367
rect 398 362 404 363
rect 430 367 436 368
rect 430 363 431 367
rect 435 363 436 367
rect 430 362 436 363
rect 454 367 460 368
rect 454 363 455 367
rect 459 366 460 367
rect 502 367 508 368
rect 459 364 465 366
rect 459 363 460 364
rect 454 362 460 363
rect 502 363 503 367
rect 507 366 508 367
rect 558 367 564 368
rect 507 364 521 366
rect 507 363 508 364
rect 502 362 508 363
rect 558 363 559 367
rect 563 366 564 367
rect 658 367 664 368
rect 563 364 585 366
rect 563 363 564 364
rect 558 362 564 363
rect 658 363 659 367
rect 663 363 664 367
rect 658 362 664 363
rect 710 367 716 368
rect 710 363 711 367
rect 715 366 716 367
rect 715 364 721 366
rect 715 363 716 364
rect 710 362 716 363
rect 638 335 644 336
rect 126 331 132 332
rect 126 327 127 331
rect 131 330 132 331
rect 174 331 180 332
rect 131 328 137 330
rect 131 327 132 328
rect 126 326 132 327
rect 174 327 175 331
rect 179 330 180 331
rect 238 331 244 332
rect 179 328 201 330
rect 179 327 180 328
rect 174 326 180 327
rect 238 327 239 331
rect 243 330 244 331
rect 310 331 316 332
rect 243 328 273 330
rect 243 327 244 328
rect 238 326 244 327
rect 310 327 311 331
rect 315 330 316 331
rect 383 331 389 332
rect 315 328 345 330
rect 315 327 316 328
rect 310 326 316 327
rect 383 327 384 331
rect 388 330 389 331
rect 598 331 604 332
rect 598 330 599 331
rect 388 328 425 330
rect 545 328 599 330
rect 388 327 389 328
rect 383 326 389 327
rect 598 327 599 328
rect 603 327 604 331
rect 638 331 639 335
rect 643 331 644 335
rect 638 330 644 331
rect 694 331 700 332
rect 598 326 604 327
rect 694 327 695 331
rect 699 330 700 331
rect 699 328 705 330
rect 699 327 700 328
rect 694 326 700 327
rect 110 325 116 326
rect 110 321 111 325
rect 115 321 116 325
rect 110 320 116 321
rect 134 325 140 326
rect 134 321 135 325
rect 139 321 140 325
rect 134 320 140 321
rect 198 325 204 326
rect 198 321 199 325
rect 203 321 204 325
rect 198 320 204 321
rect 270 325 276 326
rect 270 321 271 325
rect 275 321 276 325
rect 270 320 276 321
rect 342 325 348 326
rect 342 321 343 325
rect 347 321 348 325
rect 342 320 348 321
rect 422 325 428 326
rect 422 321 423 325
rect 427 321 428 325
rect 422 320 428 321
rect 510 325 516 326
rect 510 321 511 325
rect 515 321 516 325
rect 510 320 516 321
rect 606 325 612 326
rect 606 321 607 325
rect 611 321 612 325
rect 606 320 612 321
rect 702 325 708 326
rect 702 321 703 325
rect 707 321 708 325
rect 702 320 708 321
rect 774 325 780 326
rect 774 321 775 325
rect 779 321 780 325
rect 774 320 780 321
rect 110 307 116 308
rect 110 303 111 307
rect 115 303 116 307
rect 774 307 780 308
rect 110 302 116 303
rect 174 303 180 304
rect 174 302 175 303
rect 140 300 175 302
rect 140 296 142 300
rect 174 299 175 300
rect 179 299 180 303
rect 238 303 244 304
rect 238 302 239 303
rect 174 298 180 299
rect 204 300 239 302
rect 204 296 206 300
rect 238 299 239 300
rect 243 299 244 303
rect 310 303 316 304
rect 310 302 311 303
rect 238 298 244 299
rect 276 300 311 302
rect 276 296 278 300
rect 310 299 311 300
rect 315 299 316 303
rect 383 303 389 304
rect 383 302 384 303
rect 310 298 316 299
rect 356 300 384 302
rect 135 295 142 296
rect 135 291 136 295
rect 140 292 142 295
rect 154 295 160 296
rect 140 291 141 292
rect 135 290 141 291
rect 154 291 155 295
rect 159 291 160 295
rect 154 290 160 291
rect 199 295 206 296
rect 199 291 200 295
rect 204 292 206 295
rect 218 295 224 296
rect 204 291 205 292
rect 199 290 205 291
rect 218 291 219 295
rect 223 291 224 295
rect 218 290 224 291
rect 271 295 278 296
rect 271 291 272 295
rect 276 292 278 295
rect 290 295 296 296
rect 276 291 277 292
rect 271 290 277 291
rect 290 291 291 295
rect 295 291 296 295
rect 290 290 296 291
rect 343 295 349 296
rect 343 291 344 295
rect 348 294 349 295
rect 356 294 358 300
rect 383 299 384 300
rect 388 299 389 303
rect 774 303 775 307
rect 779 303 780 307
rect 774 302 780 303
rect 383 298 389 299
rect 348 292 358 294
rect 362 295 368 296
rect 348 291 349 292
rect 343 290 349 291
rect 362 291 363 295
rect 367 291 368 295
rect 362 290 368 291
rect 426 295 436 296
rect 426 291 427 295
rect 435 291 436 295
rect 426 290 436 291
rect 442 295 448 296
rect 442 291 443 295
rect 447 291 448 295
rect 442 290 448 291
rect 510 295 517 296
rect 510 291 511 295
rect 516 291 517 295
rect 510 290 517 291
rect 530 295 536 296
rect 530 291 531 295
rect 535 291 536 295
rect 530 290 536 291
rect 598 295 604 296
rect 598 291 599 295
rect 603 294 604 295
rect 607 295 613 296
rect 607 294 608 295
rect 603 292 608 294
rect 603 291 604 292
rect 598 290 604 291
rect 607 291 608 292
rect 612 291 613 295
rect 607 290 613 291
rect 626 295 632 296
rect 626 291 627 295
rect 631 291 632 295
rect 626 290 632 291
rect 706 295 716 296
rect 706 291 707 295
rect 715 291 716 295
rect 706 290 716 291
rect 722 295 728 296
rect 722 291 723 295
rect 727 291 728 295
rect 722 290 728 291
rect 126 279 132 280
rect 126 275 127 279
rect 131 278 132 279
rect 137 279 143 280
rect 137 278 138 279
rect 131 276 138 278
rect 131 275 132 276
rect 126 274 132 275
rect 137 275 138 276
rect 142 275 143 279
rect 694 279 700 280
rect 137 274 143 275
rect 154 277 160 278
rect 154 273 155 277
rect 159 273 160 277
rect 210 277 216 278
rect 154 272 160 273
rect 166 275 172 276
rect 166 271 167 275
rect 171 274 172 275
rect 193 275 199 276
rect 193 274 194 275
rect 171 272 194 274
rect 171 271 172 272
rect 166 270 172 271
rect 193 271 194 272
rect 198 271 199 275
rect 210 273 211 277
rect 215 273 216 277
rect 298 277 304 278
rect 210 272 216 273
rect 234 275 240 276
rect 193 270 199 271
rect 234 271 235 275
rect 239 274 240 275
rect 281 275 287 276
rect 281 274 282 275
rect 239 272 282 274
rect 239 271 240 272
rect 234 270 240 271
rect 281 271 282 272
rect 286 271 287 275
rect 298 273 299 277
rect 303 273 304 277
rect 386 277 392 278
rect 298 272 304 273
rect 310 275 316 276
rect 281 270 287 271
rect 310 271 311 275
rect 315 274 316 275
rect 369 275 375 276
rect 369 274 370 275
rect 315 272 370 274
rect 315 271 316 272
rect 310 270 316 271
rect 369 271 370 272
rect 374 271 375 275
rect 386 273 387 277
rect 391 273 392 277
rect 474 277 480 278
rect 386 272 392 273
rect 447 275 453 276
rect 369 270 375 271
rect 447 271 448 275
rect 452 274 453 275
rect 457 275 463 276
rect 457 274 458 275
rect 452 272 458 274
rect 452 271 453 272
rect 447 270 453 271
rect 457 271 458 272
rect 462 271 463 275
rect 474 273 475 277
rect 479 273 480 277
rect 562 277 568 278
rect 474 272 480 273
rect 486 275 492 276
rect 457 270 463 271
rect 486 271 487 275
rect 491 274 492 275
rect 545 275 551 276
rect 545 274 546 275
rect 491 272 546 274
rect 491 271 492 272
rect 486 270 492 271
rect 545 271 546 272
rect 550 271 551 275
rect 562 273 563 277
rect 567 273 568 277
rect 658 277 664 278
rect 562 272 568 273
rect 641 275 647 276
rect 545 270 551 271
rect 641 271 642 275
rect 646 274 647 275
rect 646 272 654 274
rect 658 273 659 277
rect 663 273 664 277
rect 694 275 695 279
rect 699 278 700 279
rect 721 279 727 280
rect 721 278 722 279
rect 699 276 722 278
rect 699 275 700 276
rect 694 274 700 275
rect 721 275 722 276
rect 726 275 727 279
rect 721 274 727 275
rect 738 277 744 278
rect 658 272 664 273
rect 738 273 739 277
rect 743 273 744 277
rect 738 272 744 273
rect 646 271 647 272
rect 641 270 647 271
rect 652 270 654 272
rect 682 271 688 272
rect 682 270 683 271
rect 652 268 683 270
rect 682 267 683 268
rect 687 267 688 271
rect 682 266 688 267
rect 110 265 116 266
rect 110 261 111 265
rect 115 261 116 265
rect 110 260 116 261
rect 774 265 780 266
rect 774 261 775 265
rect 779 261 780 265
rect 774 260 780 261
rect 110 247 116 248
rect 110 243 111 247
rect 115 243 116 247
rect 110 242 116 243
rect 134 247 140 248
rect 134 243 135 247
rect 139 243 140 247
rect 134 242 140 243
rect 190 247 196 248
rect 190 243 191 247
rect 195 243 196 247
rect 190 242 196 243
rect 278 247 284 248
rect 278 243 279 247
rect 283 243 284 247
rect 278 242 284 243
rect 366 247 372 248
rect 366 243 367 247
rect 371 243 372 247
rect 366 242 372 243
rect 454 247 460 248
rect 454 243 455 247
rect 459 243 460 247
rect 454 242 460 243
rect 542 247 548 248
rect 542 243 543 247
rect 547 243 548 247
rect 542 242 548 243
rect 638 247 644 248
rect 638 243 639 247
rect 643 243 644 247
rect 638 242 644 243
rect 718 247 724 248
rect 718 243 719 247
rect 723 243 724 247
rect 718 242 724 243
rect 774 247 780 248
rect 774 243 775 247
rect 779 243 780 247
rect 774 242 780 243
rect 166 239 172 240
rect 166 235 167 239
rect 171 235 172 239
rect 234 239 240 240
rect 234 238 235 239
rect 225 236 235 238
rect 166 234 172 235
rect 234 235 235 236
rect 239 235 240 239
rect 234 234 240 235
rect 310 239 316 240
rect 310 235 311 239
rect 315 235 316 239
rect 310 234 316 235
rect 374 239 380 240
rect 374 235 375 239
rect 379 235 380 239
rect 374 234 380 235
rect 486 239 492 240
rect 486 235 487 239
rect 491 235 492 239
rect 486 234 492 235
rect 510 239 516 240
rect 510 235 511 239
rect 515 238 516 239
rect 654 239 660 240
rect 515 236 545 238
rect 515 235 516 236
rect 510 234 516 235
rect 654 235 655 239
rect 659 235 660 239
rect 654 234 660 235
rect 682 239 688 240
rect 682 235 683 239
rect 687 238 688 239
rect 687 236 721 238
rect 687 235 688 236
rect 682 234 688 235
rect 447 207 453 208
rect 182 203 188 204
rect 182 199 183 203
rect 187 202 188 203
rect 231 203 237 204
rect 187 200 193 202
rect 187 199 188 200
rect 182 198 188 199
rect 231 199 232 203
rect 236 202 237 203
rect 326 203 332 204
rect 236 200 281 202
rect 236 199 237 200
rect 231 198 237 199
rect 326 199 327 203
rect 331 202 332 203
rect 447 203 448 207
rect 452 206 453 207
rect 452 204 457 206
rect 452 203 453 204
rect 447 202 453 203
rect 495 203 501 204
rect 331 200 369 202
rect 331 199 332 200
rect 326 198 332 199
rect 495 199 496 203
rect 500 202 501 203
rect 702 203 708 204
rect 702 202 703 203
rect 500 200 553 202
rect 681 200 703 202
rect 500 199 501 200
rect 495 198 501 199
rect 702 199 703 200
rect 707 199 708 203
rect 702 198 708 199
rect 710 203 716 204
rect 710 199 711 203
rect 715 202 716 203
rect 715 200 721 202
rect 715 199 716 200
rect 710 198 716 199
rect 110 197 116 198
rect 110 193 111 197
rect 115 193 116 197
rect 110 192 116 193
rect 190 197 196 198
rect 190 193 191 197
rect 195 193 196 197
rect 190 192 196 193
rect 278 197 284 198
rect 278 193 279 197
rect 283 193 284 197
rect 278 192 284 193
rect 366 197 372 198
rect 366 193 367 197
rect 371 193 372 197
rect 366 192 372 193
rect 454 197 460 198
rect 454 193 455 197
rect 459 193 460 197
rect 454 192 460 193
rect 550 197 556 198
rect 550 193 551 197
rect 555 193 556 197
rect 550 192 556 193
rect 646 197 652 198
rect 646 193 647 197
rect 651 193 652 197
rect 646 192 652 193
rect 718 197 724 198
rect 718 193 719 197
rect 723 193 724 197
rect 718 192 724 193
rect 774 197 780 198
rect 774 193 775 197
rect 779 193 780 197
rect 774 192 780 193
rect 110 179 116 180
rect 110 175 111 179
rect 115 175 116 179
rect 774 179 780 180
rect 110 174 116 175
rect 231 175 237 176
rect 231 174 232 175
rect 204 172 232 174
rect 191 167 197 168
rect 191 163 192 167
rect 196 166 197 167
rect 204 166 206 172
rect 231 171 232 172
rect 236 171 237 175
rect 326 175 332 176
rect 326 174 327 175
rect 231 170 237 171
rect 284 172 327 174
rect 284 168 286 172
rect 326 171 327 172
rect 331 171 332 175
rect 495 175 501 176
rect 495 174 496 175
rect 326 170 332 171
rect 460 172 496 174
rect 460 168 462 172
rect 495 171 496 172
rect 500 171 501 175
rect 774 175 775 179
rect 779 175 780 179
rect 774 174 780 175
rect 495 170 501 171
rect 196 164 206 166
rect 210 167 216 168
rect 196 163 197 164
rect 191 162 197 163
rect 210 163 211 167
rect 215 163 216 167
rect 210 162 216 163
rect 279 167 286 168
rect 279 163 280 167
rect 284 164 286 167
rect 298 167 304 168
rect 284 163 285 164
rect 279 162 285 163
rect 298 163 299 167
rect 303 163 304 167
rect 298 162 304 163
rect 370 167 380 168
rect 370 163 371 167
rect 379 163 380 167
rect 370 162 380 163
rect 386 167 392 168
rect 386 163 387 167
rect 391 163 392 167
rect 386 162 392 163
rect 455 167 462 168
rect 455 163 456 167
rect 460 164 462 167
rect 474 167 480 168
rect 460 163 461 164
rect 455 162 461 163
rect 474 163 475 167
rect 479 163 480 167
rect 474 162 480 163
rect 551 167 557 168
rect 551 163 552 167
rect 556 166 557 167
rect 570 167 576 168
rect 556 163 558 166
rect 551 162 558 163
rect 570 163 571 167
rect 575 163 576 167
rect 570 162 576 163
rect 650 167 660 168
rect 650 163 651 167
rect 659 163 660 167
rect 650 162 660 163
rect 666 167 672 168
rect 666 163 667 167
rect 671 163 672 167
rect 666 162 672 163
rect 702 167 708 168
rect 702 163 703 167
rect 707 166 708 167
rect 719 167 725 168
rect 719 166 720 167
rect 707 164 720 166
rect 707 163 708 164
rect 702 162 708 163
rect 719 163 720 164
rect 724 163 725 167
rect 719 162 725 163
rect 738 167 744 168
rect 738 163 739 167
rect 743 163 744 167
rect 738 162 744 163
rect 556 158 558 162
rect 567 159 573 160
rect 567 158 568 159
rect 556 156 568 158
rect 567 155 568 156
rect 572 155 573 159
rect 567 154 573 155
rect 182 151 188 152
rect 182 147 183 151
rect 187 150 188 151
rect 193 151 199 152
rect 193 150 194 151
rect 187 148 194 150
rect 187 147 188 148
rect 182 146 188 147
rect 193 147 194 148
rect 198 147 199 151
rect 710 151 716 152
rect 193 146 199 147
rect 210 149 216 150
rect 210 145 211 149
rect 215 145 216 149
rect 258 149 264 150
rect 210 144 216 145
rect 222 147 228 148
rect 222 143 223 147
rect 227 146 228 147
rect 241 147 247 148
rect 241 146 242 147
rect 227 144 242 146
rect 227 143 228 144
rect 222 142 228 143
rect 241 143 242 144
rect 246 143 247 147
rect 258 145 259 149
rect 263 145 264 149
rect 306 149 312 150
rect 258 144 264 145
rect 270 147 276 148
rect 241 142 247 143
rect 270 143 271 147
rect 275 146 276 147
rect 289 147 295 148
rect 289 146 290 147
rect 275 144 290 146
rect 275 143 276 144
rect 270 142 276 143
rect 289 143 290 144
rect 294 143 295 147
rect 306 145 307 149
rect 311 145 312 149
rect 354 149 360 150
rect 306 144 312 145
rect 318 147 324 148
rect 289 142 295 143
rect 318 143 319 147
rect 323 146 324 147
rect 337 147 343 148
rect 337 146 338 147
rect 323 144 338 146
rect 323 143 324 144
rect 318 142 324 143
rect 337 143 338 144
rect 342 143 343 147
rect 354 145 355 149
rect 359 145 360 149
rect 402 149 408 150
rect 354 144 360 145
rect 366 147 372 148
rect 337 142 343 143
rect 366 143 367 147
rect 371 146 372 147
rect 385 147 391 148
rect 385 146 386 147
rect 371 144 386 146
rect 371 143 372 144
rect 366 142 372 143
rect 385 143 386 144
rect 390 143 391 147
rect 402 145 403 149
rect 407 145 408 149
rect 450 149 456 150
rect 402 144 408 145
rect 414 147 420 148
rect 385 142 391 143
rect 414 143 415 147
rect 419 146 420 147
rect 433 147 439 148
rect 433 146 434 147
rect 419 144 434 146
rect 419 143 420 144
rect 414 142 420 143
rect 433 143 434 144
rect 438 143 439 147
rect 450 145 451 149
rect 455 145 456 149
rect 498 149 504 150
rect 450 144 456 145
rect 462 147 468 148
rect 433 142 439 143
rect 462 143 463 147
rect 467 146 468 147
rect 481 147 487 148
rect 481 146 482 147
rect 467 144 482 146
rect 467 143 468 144
rect 462 142 468 143
rect 481 143 482 144
rect 486 143 487 147
rect 498 145 499 149
rect 503 145 504 149
rect 546 149 552 150
rect 498 144 504 145
rect 510 147 516 148
rect 481 142 487 143
rect 510 143 511 147
rect 515 146 516 147
rect 529 147 535 148
rect 529 146 530 147
rect 515 144 530 146
rect 515 143 516 144
rect 510 142 516 143
rect 529 143 530 144
rect 534 143 535 147
rect 546 145 547 149
rect 551 145 552 149
rect 594 149 600 150
rect 546 144 552 145
rect 558 147 564 148
rect 529 142 535 143
rect 558 143 559 147
rect 563 146 564 147
rect 577 147 583 148
rect 577 146 578 147
rect 563 144 578 146
rect 563 143 564 144
rect 558 142 564 143
rect 577 143 578 144
rect 582 143 583 147
rect 594 145 595 149
rect 599 145 600 149
rect 642 149 648 150
rect 594 144 600 145
rect 625 147 631 148
rect 577 142 583 143
rect 625 143 626 147
rect 630 146 631 147
rect 630 144 638 146
rect 642 145 643 149
rect 647 145 648 149
rect 690 149 696 150
rect 642 144 648 145
rect 673 147 679 148
rect 630 143 631 144
rect 625 142 631 143
rect 636 142 638 144
rect 662 143 668 144
rect 662 142 663 143
rect 636 140 663 142
rect 662 139 663 140
rect 667 139 668 143
rect 673 143 674 147
rect 678 146 679 147
rect 678 144 686 146
rect 690 145 691 149
rect 695 145 696 149
rect 710 147 711 151
rect 715 150 716 151
rect 721 151 727 152
rect 721 150 722 151
rect 715 148 722 150
rect 715 147 716 148
rect 710 146 716 147
rect 721 147 722 148
rect 726 147 727 151
rect 721 146 727 147
rect 738 149 744 150
rect 690 144 696 145
rect 738 145 739 149
rect 743 145 744 149
rect 738 144 744 145
rect 678 143 679 144
rect 673 142 679 143
rect 684 142 686 144
rect 710 143 716 144
rect 710 142 711 143
rect 684 140 711 142
rect 662 138 668 139
rect 710 139 711 140
rect 715 139 716 143
rect 710 138 716 139
rect 110 137 116 138
rect 110 133 111 137
rect 115 133 116 137
rect 110 132 116 133
rect 774 137 780 138
rect 774 133 775 137
rect 779 133 780 137
rect 774 132 780 133
rect 110 119 116 120
rect 110 115 111 119
rect 115 115 116 119
rect 110 114 116 115
rect 190 119 196 120
rect 190 115 191 119
rect 195 115 196 119
rect 190 114 196 115
rect 238 119 244 120
rect 238 115 239 119
rect 243 115 244 119
rect 238 114 244 115
rect 286 119 292 120
rect 286 115 287 119
rect 291 115 292 119
rect 286 114 292 115
rect 334 119 340 120
rect 334 115 335 119
rect 339 115 340 119
rect 334 114 340 115
rect 382 119 388 120
rect 382 115 383 119
rect 387 115 388 119
rect 382 114 388 115
rect 430 119 436 120
rect 430 115 431 119
rect 435 115 436 119
rect 430 114 436 115
rect 478 119 484 120
rect 478 115 479 119
rect 483 115 484 119
rect 478 114 484 115
rect 526 119 532 120
rect 526 115 527 119
rect 531 115 532 119
rect 526 114 532 115
rect 574 119 580 120
rect 574 115 575 119
rect 579 115 580 119
rect 574 114 580 115
rect 622 119 628 120
rect 622 115 623 119
rect 627 115 628 119
rect 622 114 628 115
rect 670 119 676 120
rect 670 115 671 119
rect 675 115 676 119
rect 670 114 676 115
rect 718 119 724 120
rect 718 115 719 119
rect 723 115 724 119
rect 718 114 724 115
rect 774 119 780 120
rect 774 115 775 119
rect 779 115 780 119
rect 774 114 780 115
rect 222 111 228 112
rect 222 107 223 111
rect 227 107 228 111
rect 222 106 228 107
rect 270 111 276 112
rect 270 107 271 111
rect 275 107 276 111
rect 270 106 276 107
rect 318 111 324 112
rect 318 107 319 111
rect 323 107 324 111
rect 318 106 324 107
rect 366 111 372 112
rect 366 107 367 111
rect 371 107 372 111
rect 366 106 372 107
rect 414 111 420 112
rect 414 107 415 111
rect 419 107 420 111
rect 414 106 420 107
rect 462 111 468 112
rect 462 107 463 111
rect 467 107 468 111
rect 462 106 468 107
rect 510 111 516 112
rect 510 107 511 111
rect 515 107 516 111
rect 510 106 516 107
rect 558 111 564 112
rect 558 107 559 111
rect 563 107 564 111
rect 558 106 564 107
rect 567 111 573 112
rect 567 107 568 111
rect 572 110 573 111
rect 662 111 668 112
rect 572 108 577 110
rect 572 107 573 108
rect 567 106 573 107
rect 662 107 663 111
rect 667 110 668 111
rect 710 111 716 112
rect 667 108 673 110
rect 667 107 668 108
rect 662 106 668 107
rect 710 107 711 111
rect 715 110 716 111
rect 715 108 721 110
rect 715 107 716 108
rect 710 106 716 107
<< m3c >>
rect 155 853 159 857
rect 175 847 179 851
rect 203 853 207 857
rect 251 853 255 857
rect 223 847 227 851
rect 111 841 115 845
rect 775 841 779 845
rect 111 823 115 827
rect 135 823 139 827
rect 183 823 187 827
rect 231 823 235 827
rect 775 823 779 827
rect 143 815 147 819
rect 175 815 179 819
rect 223 815 227 819
rect 175 787 179 791
rect 223 787 227 791
rect 271 787 275 791
rect 319 787 323 791
rect 367 787 371 791
rect 111 781 115 785
rect 135 781 139 785
rect 183 781 187 785
rect 231 781 235 785
rect 279 781 283 785
rect 327 781 331 785
rect 375 781 379 785
rect 775 781 779 785
rect 111 763 115 767
rect 279 759 283 763
rect 775 763 779 767
rect 143 751 147 755
rect 155 751 159 755
rect 175 751 179 755
rect 203 751 207 755
rect 223 751 227 755
rect 251 751 255 755
rect 271 751 275 755
rect 299 751 303 755
rect 319 751 323 755
rect 347 751 351 755
rect 367 751 371 755
rect 395 751 399 755
rect 279 743 283 747
rect 291 741 295 745
rect 311 739 315 743
rect 339 741 343 745
rect 359 739 363 743
rect 387 741 391 745
rect 407 739 411 743
rect 443 741 447 745
rect 455 739 459 743
rect 507 741 511 745
rect 519 739 523 743
rect 579 741 583 745
rect 647 739 651 743
rect 659 741 663 745
rect 671 739 675 743
rect 739 741 743 745
rect 111 729 115 733
rect 775 729 779 733
rect 111 711 115 715
rect 271 711 275 715
rect 319 711 323 715
rect 367 711 371 715
rect 423 711 427 715
rect 487 711 491 715
rect 559 711 563 715
rect 639 711 643 715
rect 719 711 723 715
rect 775 711 779 715
rect 311 703 315 707
rect 359 703 363 707
rect 407 703 411 707
rect 455 703 459 707
rect 519 703 523 707
rect 535 703 539 707
rect 671 703 675 707
rect 679 703 683 707
rect 367 679 371 683
rect 423 675 427 679
rect 471 675 475 679
rect 519 675 523 679
rect 615 675 619 679
rect 655 679 659 683
rect 703 679 707 683
rect 711 675 715 679
rect 111 669 115 673
rect 335 669 339 673
rect 383 669 387 673
rect 431 669 435 673
rect 479 669 483 673
rect 527 669 531 673
rect 575 669 579 673
rect 623 669 627 673
rect 671 669 675 673
rect 719 669 723 673
rect 775 669 779 673
rect 111 651 115 655
rect 519 647 523 651
rect 775 651 779 655
rect 355 639 359 643
rect 367 639 371 643
rect 403 639 407 643
rect 423 639 427 643
rect 451 639 455 643
rect 499 639 503 643
rect 535 639 539 643
rect 547 639 551 643
rect 575 639 576 643
rect 576 639 579 643
rect 595 639 599 643
rect 615 639 619 643
rect 643 639 647 643
rect 679 639 683 643
rect 691 639 695 643
rect 703 639 707 643
rect 739 639 743 643
rect 155 629 159 633
rect 175 623 179 627
rect 203 629 207 633
rect 223 623 227 627
rect 275 629 279 633
rect 311 623 315 627
rect 379 629 383 633
rect 471 631 475 635
rect 499 629 503 633
rect 511 627 515 631
rect 627 629 631 633
rect 711 631 715 635
rect 739 629 743 633
rect 111 617 115 621
rect 519 619 523 623
rect 775 617 779 621
rect 111 599 115 603
rect 135 599 139 603
rect 183 599 187 603
rect 255 599 259 603
rect 359 599 363 603
rect 479 599 483 603
rect 607 599 611 603
rect 719 599 723 603
rect 775 599 779 603
rect 143 591 147 595
rect 175 591 179 595
rect 223 591 227 595
rect 311 591 315 595
rect 511 591 515 595
rect 519 591 523 595
rect 727 591 731 595
rect 391 571 395 575
rect 175 563 179 567
rect 223 563 227 567
rect 343 563 347 567
rect 439 563 443 567
rect 575 567 579 571
rect 671 567 675 571
rect 111 557 115 561
rect 135 557 139 561
rect 183 557 187 561
rect 263 557 267 561
rect 351 557 355 561
rect 447 557 451 561
rect 543 557 547 561
rect 639 557 643 561
rect 719 557 723 561
rect 775 557 779 561
rect 111 539 115 543
rect 143 527 147 531
rect 155 527 159 531
rect 175 527 179 531
rect 391 535 395 539
rect 203 527 207 531
rect 223 527 227 531
rect 283 527 287 531
rect 343 527 347 531
rect 371 527 375 531
rect 439 527 443 531
rect 467 527 471 531
rect 591 535 595 539
rect 775 539 779 543
rect 563 527 567 531
rect 659 527 663 531
rect 727 527 731 531
rect 739 527 743 531
rect 211 517 215 521
rect 223 515 227 519
rect 267 517 271 521
rect 331 517 335 521
rect 343 515 347 519
rect 403 517 407 521
rect 415 515 419 519
rect 483 517 487 521
rect 495 515 499 519
rect 571 517 575 521
rect 667 517 671 521
rect 675 519 679 523
rect 739 517 743 521
rect 655 511 659 515
rect 111 505 115 509
rect 775 505 779 509
rect 111 487 115 491
rect 191 487 195 491
rect 247 487 251 491
rect 311 487 315 491
rect 383 487 387 491
rect 463 487 467 491
rect 551 487 555 491
rect 647 487 651 491
rect 719 487 723 491
rect 775 487 779 491
rect 223 479 227 483
rect 343 479 347 483
rect 415 479 419 483
rect 495 479 499 483
rect 503 479 507 483
rect 591 479 595 483
rect 727 479 731 483
rect 391 451 395 455
rect 439 451 443 455
rect 487 451 491 455
rect 535 451 539 455
rect 575 455 579 459
rect 587 451 591 455
rect 655 455 659 459
rect 711 451 715 455
rect 111 445 115 449
rect 351 445 355 449
rect 399 445 403 449
rect 447 445 451 449
rect 495 445 499 449
rect 543 445 547 449
rect 599 445 603 449
rect 663 445 667 449
rect 719 445 723 449
rect 775 445 779 449
rect 111 427 115 431
rect 503 423 507 427
rect 775 427 779 431
rect 371 415 375 419
rect 391 415 395 419
rect 419 415 423 419
rect 439 415 443 419
rect 467 415 471 419
rect 487 415 491 419
rect 515 415 519 419
rect 535 415 539 419
rect 563 415 567 419
rect 575 415 579 419
rect 619 415 623 419
rect 659 415 663 419
rect 683 415 687 419
rect 727 415 731 419
rect 739 415 743 419
rect 339 401 343 405
rect 351 399 355 403
rect 387 401 391 405
rect 399 399 403 403
rect 435 401 439 405
rect 483 401 487 405
rect 111 389 115 393
rect 455 391 459 395
rect 503 395 507 399
rect 539 401 543 405
rect 587 403 590 407
rect 590 403 591 407
rect 603 401 607 405
rect 559 395 563 399
rect 639 399 643 403
rect 667 401 671 405
rect 711 403 715 407
rect 739 401 743 405
rect 775 389 779 393
rect 111 371 115 375
rect 319 371 323 375
rect 367 371 371 375
rect 415 371 419 375
rect 463 371 467 375
rect 519 371 523 375
rect 583 371 587 375
rect 647 371 651 375
rect 719 371 723 375
rect 775 371 779 375
rect 351 363 355 367
rect 399 363 403 367
rect 431 363 435 367
rect 455 363 459 367
rect 503 363 507 367
rect 559 363 563 367
rect 659 363 663 367
rect 711 363 715 367
rect 127 327 131 331
rect 175 327 179 331
rect 239 327 243 331
rect 311 327 315 331
rect 599 327 603 331
rect 639 331 643 335
rect 695 327 699 331
rect 111 321 115 325
rect 135 321 139 325
rect 199 321 203 325
rect 271 321 275 325
rect 343 321 347 325
rect 423 321 427 325
rect 511 321 515 325
rect 607 321 611 325
rect 703 321 707 325
rect 775 321 779 325
rect 111 303 115 307
rect 175 299 179 303
rect 239 299 243 303
rect 311 299 315 303
rect 155 291 159 295
rect 219 291 223 295
rect 291 291 295 295
rect 775 303 779 307
rect 363 291 367 295
rect 431 291 435 295
rect 443 291 447 295
rect 511 291 512 295
rect 512 291 515 295
rect 531 291 535 295
rect 599 291 603 295
rect 627 291 631 295
rect 711 291 715 295
rect 723 291 727 295
rect 127 275 131 279
rect 155 273 159 277
rect 167 271 171 275
rect 211 273 215 277
rect 235 271 239 275
rect 299 273 303 277
rect 311 271 315 275
rect 387 273 391 277
rect 475 273 479 277
rect 487 271 491 275
rect 563 273 567 277
rect 659 273 663 277
rect 695 275 699 279
rect 739 273 743 277
rect 683 267 687 271
rect 111 261 115 265
rect 775 261 779 265
rect 111 243 115 247
rect 135 243 139 247
rect 191 243 195 247
rect 279 243 283 247
rect 367 243 371 247
rect 455 243 459 247
rect 543 243 547 247
rect 639 243 643 247
rect 719 243 723 247
rect 775 243 779 247
rect 167 235 171 239
rect 235 235 239 239
rect 311 235 315 239
rect 375 235 379 239
rect 487 235 491 239
rect 511 235 515 239
rect 655 235 659 239
rect 683 235 687 239
rect 183 199 187 203
rect 327 199 331 203
rect 703 199 707 203
rect 711 199 715 203
rect 111 193 115 197
rect 191 193 195 197
rect 279 193 283 197
rect 367 193 371 197
rect 455 193 459 197
rect 551 193 555 197
rect 647 193 651 197
rect 719 193 723 197
rect 775 193 779 197
rect 111 175 115 179
rect 327 171 331 175
rect 775 175 779 179
rect 211 163 215 167
rect 299 163 303 167
rect 375 163 379 167
rect 387 163 391 167
rect 475 163 479 167
rect 571 163 575 167
rect 655 163 659 167
rect 667 163 671 167
rect 703 163 707 167
rect 739 163 743 167
rect 183 147 187 151
rect 211 145 215 149
rect 223 143 227 147
rect 259 145 263 149
rect 271 143 275 147
rect 307 145 311 149
rect 319 143 323 147
rect 355 145 359 149
rect 367 143 371 147
rect 403 145 407 149
rect 415 143 419 147
rect 451 145 455 149
rect 463 143 467 147
rect 499 145 503 149
rect 511 143 515 147
rect 547 145 551 149
rect 559 143 563 147
rect 595 145 599 149
rect 643 145 647 149
rect 663 139 667 143
rect 691 145 695 149
rect 711 147 715 151
rect 739 145 743 149
rect 711 139 715 143
rect 111 133 115 137
rect 775 133 779 137
rect 111 115 115 119
rect 191 115 195 119
rect 239 115 243 119
rect 287 115 291 119
rect 335 115 339 119
rect 383 115 387 119
rect 431 115 435 119
rect 479 115 483 119
rect 527 115 531 119
rect 575 115 579 119
rect 623 115 627 119
rect 671 115 675 119
rect 719 115 723 119
rect 775 115 779 119
rect 223 107 227 111
rect 271 107 275 111
rect 319 107 323 111
rect 367 107 371 111
rect 415 107 419 111
rect 463 107 467 111
rect 511 107 515 111
rect 559 107 563 111
rect 663 107 667 111
rect 711 107 715 111
<< m3 >>
rect 111 862 115 863
rect 155 862 159 863
rect 203 862 207 863
rect 251 862 255 863
rect 775 862 779 863
rect 111 857 115 858
rect 154 857 160 858
rect 112 846 114 857
rect 154 853 155 857
rect 159 853 160 857
rect 154 852 160 853
rect 202 857 208 858
rect 202 853 203 857
rect 207 853 208 857
rect 202 852 208 853
rect 250 857 256 858
rect 775 857 779 858
rect 250 853 251 857
rect 255 853 256 857
rect 250 852 256 853
rect 174 851 180 852
rect 174 847 175 851
rect 179 847 180 851
rect 174 846 180 847
rect 222 851 228 852
rect 222 847 223 851
rect 227 847 228 851
rect 222 846 228 847
rect 776 846 778 857
rect 110 845 116 846
rect 110 841 111 845
rect 115 841 116 845
rect 110 840 116 841
rect 110 827 116 828
rect 110 823 111 827
rect 115 823 116 827
rect 110 822 116 823
rect 134 827 140 828
rect 134 823 135 827
rect 139 823 140 827
rect 134 822 140 823
rect 112 807 114 822
rect 136 807 138 822
rect 176 820 178 846
rect 182 827 188 828
rect 182 823 183 827
rect 187 823 188 827
rect 182 822 188 823
rect 142 819 148 820
rect 142 815 143 819
rect 147 815 148 819
rect 142 814 148 815
rect 174 819 180 820
rect 174 815 175 819
rect 179 815 180 819
rect 174 814 180 815
rect 111 806 115 807
rect 111 801 115 802
rect 135 806 139 807
rect 135 801 139 802
rect 112 786 114 801
rect 136 786 138 801
rect 110 785 116 786
rect 110 781 111 785
rect 115 781 116 785
rect 110 780 116 781
rect 134 785 140 786
rect 134 781 135 785
rect 139 781 140 785
rect 134 780 140 781
rect 110 767 116 768
rect 110 763 111 767
rect 115 763 116 767
rect 110 762 116 763
rect 112 751 114 762
rect 144 756 146 814
rect 184 807 186 822
rect 224 820 226 846
rect 774 845 780 846
rect 774 841 775 845
rect 779 841 780 845
rect 774 840 780 841
rect 230 827 236 828
rect 230 823 231 827
rect 235 823 236 827
rect 230 822 236 823
rect 774 827 780 828
rect 774 823 775 827
rect 779 823 780 827
rect 774 822 780 823
rect 222 819 228 820
rect 222 815 223 819
rect 227 815 228 819
rect 222 814 228 815
rect 232 807 234 822
rect 776 807 778 822
rect 183 806 187 807
rect 183 801 187 802
rect 231 806 235 807
rect 231 801 235 802
rect 279 806 283 807
rect 279 801 283 802
rect 327 806 331 807
rect 327 801 331 802
rect 375 806 379 807
rect 375 801 379 802
rect 775 806 779 807
rect 775 801 779 802
rect 174 791 180 792
rect 174 787 175 791
rect 179 787 180 791
rect 174 786 180 787
rect 184 786 186 801
rect 222 791 228 792
rect 222 787 223 791
rect 227 787 228 791
rect 222 786 228 787
rect 232 786 234 801
rect 270 791 276 792
rect 270 787 271 791
rect 275 787 276 791
rect 270 786 276 787
rect 280 786 282 801
rect 318 791 324 792
rect 318 787 319 791
rect 323 787 324 791
rect 318 786 324 787
rect 328 786 330 801
rect 366 791 372 792
rect 366 787 367 791
rect 371 787 372 791
rect 366 786 372 787
rect 376 786 378 801
rect 776 786 778 801
rect 176 756 178 786
rect 182 785 188 786
rect 182 781 183 785
rect 187 781 188 785
rect 182 780 188 781
rect 224 756 226 786
rect 230 785 236 786
rect 230 781 231 785
rect 235 781 236 785
rect 230 780 236 781
rect 272 756 274 786
rect 278 785 284 786
rect 278 781 279 785
rect 283 781 284 785
rect 278 780 284 781
rect 278 763 284 764
rect 278 759 279 763
rect 283 759 284 763
rect 278 758 284 759
rect 142 755 148 756
rect 142 751 143 755
rect 147 751 148 755
rect 111 750 115 751
rect 142 750 148 751
rect 154 755 160 756
rect 154 751 155 755
rect 159 751 160 755
rect 154 750 160 751
rect 174 755 180 756
rect 174 751 175 755
rect 179 751 180 755
rect 174 750 180 751
rect 202 755 208 756
rect 202 751 203 755
rect 207 751 208 755
rect 202 750 208 751
rect 222 755 228 756
rect 222 751 223 755
rect 227 751 228 755
rect 222 750 228 751
rect 250 755 256 756
rect 250 751 251 755
rect 255 751 256 755
rect 250 750 256 751
rect 270 755 276 756
rect 270 751 271 755
rect 275 751 276 755
rect 270 750 276 751
rect 111 745 115 746
rect 155 745 159 746
rect 203 745 207 746
rect 280 748 282 758
rect 320 756 322 786
rect 326 785 332 786
rect 326 781 327 785
rect 331 781 332 785
rect 326 780 332 781
rect 368 756 370 786
rect 374 785 380 786
rect 374 781 375 785
rect 379 781 380 785
rect 374 780 380 781
rect 774 785 780 786
rect 774 781 775 785
rect 779 781 780 785
rect 774 780 780 781
rect 774 767 780 768
rect 774 763 775 767
rect 779 763 780 767
rect 774 762 780 763
rect 298 755 304 756
rect 298 751 299 755
rect 303 751 304 755
rect 291 750 295 751
rect 298 750 304 751
rect 318 755 324 756
rect 318 751 319 755
rect 323 751 324 755
rect 346 755 352 756
rect 346 751 347 755
rect 351 751 352 755
rect 318 750 324 751
rect 339 750 343 751
rect 346 750 352 751
rect 366 755 372 756
rect 366 751 367 755
rect 371 751 372 755
rect 394 755 400 756
rect 394 751 395 755
rect 399 751 400 755
rect 776 751 778 762
rect 366 750 372 751
rect 387 750 391 751
rect 394 750 400 751
rect 443 750 447 751
rect 251 745 255 746
rect 278 747 284 748
rect 112 734 114 745
rect 278 743 279 747
rect 283 743 284 747
rect 507 750 511 751
rect 579 750 583 751
rect 659 750 663 751
rect 739 750 743 751
rect 775 750 779 751
rect 278 742 284 743
rect 290 745 296 746
rect 299 745 303 746
rect 338 745 344 746
rect 347 745 351 746
rect 386 745 392 746
rect 395 745 399 746
rect 442 745 448 746
rect 290 741 291 745
rect 295 741 296 745
rect 290 740 296 741
rect 310 743 316 744
rect 310 739 311 743
rect 315 739 316 743
rect 338 741 339 745
rect 343 741 344 745
rect 338 740 344 741
rect 358 743 364 744
rect 310 738 316 739
rect 358 739 359 743
rect 363 739 364 743
rect 386 741 387 745
rect 391 741 392 745
rect 386 740 392 741
rect 406 743 412 744
rect 358 738 364 739
rect 406 739 407 743
rect 411 739 412 743
rect 442 741 443 745
rect 447 741 448 745
rect 506 745 512 746
rect 442 740 448 741
rect 454 743 460 744
rect 406 738 412 739
rect 454 739 455 743
rect 459 739 460 743
rect 506 741 507 745
rect 511 741 512 745
rect 578 745 584 746
rect 506 740 512 741
rect 518 743 524 744
rect 454 738 460 739
rect 518 739 519 743
rect 523 739 524 743
rect 578 741 579 745
rect 583 741 584 745
rect 658 745 664 746
rect 578 740 584 741
rect 646 743 652 744
rect 518 738 524 739
rect 646 739 647 743
rect 651 739 652 743
rect 658 741 659 745
rect 663 741 664 745
rect 738 745 744 746
rect 775 745 779 746
rect 658 740 664 741
rect 670 743 676 744
rect 646 738 652 739
rect 670 739 671 743
rect 675 739 676 743
rect 738 741 739 745
rect 743 741 744 745
rect 738 740 744 741
rect 670 738 676 739
rect 110 733 116 734
rect 110 729 111 733
rect 115 729 116 733
rect 110 728 116 729
rect 110 715 116 716
rect 110 711 111 715
rect 115 711 116 715
rect 110 710 116 711
rect 270 715 276 716
rect 270 711 271 715
rect 275 711 276 715
rect 270 710 276 711
rect 112 695 114 710
rect 272 695 274 710
rect 312 708 314 738
rect 318 715 324 716
rect 318 711 319 715
rect 323 711 324 715
rect 318 710 324 711
rect 310 707 316 708
rect 310 703 311 707
rect 315 703 316 707
rect 310 702 316 703
rect 320 695 322 710
rect 360 708 362 738
rect 366 715 372 716
rect 366 711 367 715
rect 371 711 372 715
rect 366 710 372 711
rect 358 707 364 708
rect 358 703 359 707
rect 363 703 364 707
rect 358 702 364 703
rect 368 695 370 710
rect 408 708 410 738
rect 422 715 428 716
rect 422 711 423 715
rect 427 711 428 715
rect 422 710 428 711
rect 406 707 412 708
rect 406 703 407 707
rect 411 703 412 707
rect 406 702 412 703
rect 424 695 426 710
rect 456 708 458 738
rect 486 715 492 716
rect 486 711 487 715
rect 491 711 492 715
rect 486 710 492 711
rect 454 707 460 708
rect 454 703 455 707
rect 459 703 460 707
rect 454 702 460 703
rect 488 695 490 710
rect 520 708 522 738
rect 648 731 650 738
rect 648 729 658 731
rect 558 715 564 716
rect 558 711 559 715
rect 563 711 564 715
rect 558 710 564 711
rect 638 715 644 716
rect 638 711 639 715
rect 643 711 644 715
rect 638 710 644 711
rect 518 707 524 708
rect 518 703 519 707
rect 523 703 524 707
rect 518 702 524 703
rect 534 707 540 708
rect 534 703 535 707
rect 539 703 540 707
rect 534 702 540 703
rect 111 694 115 695
rect 111 689 115 690
rect 271 694 275 695
rect 271 689 275 690
rect 319 694 323 695
rect 319 689 323 690
rect 335 694 339 695
rect 335 689 339 690
rect 367 694 371 695
rect 367 689 371 690
rect 383 694 387 695
rect 383 689 387 690
rect 423 694 427 695
rect 423 689 427 690
rect 431 694 435 695
rect 431 689 435 690
rect 479 694 483 695
rect 479 689 483 690
rect 487 694 491 695
rect 487 689 491 690
rect 527 694 531 695
rect 527 689 531 690
rect 112 674 114 689
rect 336 674 338 689
rect 366 683 372 684
rect 366 679 367 683
rect 371 679 372 683
rect 366 678 372 679
rect 110 673 116 674
rect 110 669 111 673
rect 115 669 116 673
rect 110 668 116 669
rect 334 673 340 674
rect 334 669 335 673
rect 339 669 340 673
rect 334 668 340 669
rect 110 655 116 656
rect 110 651 111 655
rect 115 651 116 655
rect 110 650 116 651
rect 112 639 114 650
rect 368 644 370 678
rect 384 674 386 689
rect 422 679 428 680
rect 422 675 423 679
rect 427 675 428 679
rect 422 674 428 675
rect 432 674 434 689
rect 470 679 476 680
rect 470 675 471 679
rect 475 675 476 679
rect 470 674 476 675
rect 480 674 482 689
rect 518 679 524 680
rect 518 675 519 679
rect 523 675 524 679
rect 518 674 524 675
rect 528 674 530 689
rect 382 673 388 674
rect 382 669 383 673
rect 387 669 388 673
rect 382 668 388 669
rect 424 644 426 674
rect 430 673 436 674
rect 430 669 431 673
rect 435 669 436 673
rect 430 668 436 669
rect 354 643 360 644
rect 354 639 355 643
rect 359 639 360 643
rect 111 638 115 639
rect 155 638 159 639
rect 203 638 207 639
rect 275 638 279 639
rect 354 638 360 639
rect 366 643 372 644
rect 366 639 367 643
rect 371 639 372 643
rect 402 643 408 644
rect 402 639 403 643
rect 407 639 408 643
rect 366 638 372 639
rect 379 638 383 639
rect 402 638 408 639
rect 422 643 428 644
rect 422 639 423 643
rect 427 639 428 643
rect 422 638 428 639
rect 450 643 456 644
rect 450 639 451 643
rect 455 639 456 643
rect 450 638 456 639
rect 111 633 115 634
rect 154 633 160 634
rect 112 622 114 633
rect 154 629 155 633
rect 159 629 160 633
rect 154 628 160 629
rect 202 633 208 634
rect 202 629 203 633
rect 207 629 208 633
rect 202 628 208 629
rect 274 633 280 634
rect 355 633 359 634
rect 378 633 384 634
rect 403 633 407 634
rect 472 636 474 674
rect 478 673 484 674
rect 478 669 479 673
rect 483 669 484 673
rect 478 668 484 669
rect 520 652 522 674
rect 526 673 532 674
rect 526 669 527 673
rect 531 669 532 673
rect 526 668 532 669
rect 518 651 524 652
rect 518 647 519 651
rect 523 647 524 651
rect 518 646 524 647
rect 536 644 538 702
rect 560 695 562 710
rect 640 695 642 710
rect 559 694 563 695
rect 559 689 563 690
rect 575 694 579 695
rect 575 689 579 690
rect 623 694 627 695
rect 623 689 627 690
rect 639 694 643 695
rect 639 689 643 690
rect 576 674 578 689
rect 614 679 620 680
rect 614 675 615 679
rect 619 675 620 679
rect 614 674 620 675
rect 624 674 626 689
rect 656 684 658 729
rect 672 708 674 738
rect 776 734 778 745
rect 774 733 780 734
rect 774 729 775 733
rect 779 729 780 733
rect 774 728 780 729
rect 718 715 724 716
rect 718 711 719 715
rect 723 711 724 715
rect 718 710 724 711
rect 774 715 780 716
rect 774 711 775 715
rect 779 711 780 715
rect 774 710 780 711
rect 670 707 676 708
rect 670 703 671 707
rect 675 703 676 707
rect 670 702 676 703
rect 678 707 684 708
rect 678 703 679 707
rect 683 703 684 707
rect 678 702 684 703
rect 671 694 675 695
rect 671 689 675 690
rect 654 683 660 684
rect 654 679 655 683
rect 659 679 660 683
rect 654 678 660 679
rect 672 674 674 689
rect 574 673 580 674
rect 574 669 575 673
rect 579 669 580 673
rect 574 668 580 669
rect 616 644 618 674
rect 622 673 628 674
rect 622 669 623 673
rect 627 669 628 673
rect 622 668 628 669
rect 670 673 676 674
rect 670 669 671 673
rect 675 669 676 673
rect 670 668 676 669
rect 680 644 682 702
rect 720 695 722 710
rect 776 695 778 710
rect 719 694 723 695
rect 719 689 723 690
rect 775 694 779 695
rect 775 689 779 690
rect 702 683 708 684
rect 702 679 703 683
rect 707 679 708 683
rect 702 678 708 679
rect 710 679 716 680
rect 704 644 706 678
rect 710 675 711 679
rect 715 675 716 679
rect 710 674 716 675
rect 720 674 722 689
rect 776 674 778 689
rect 498 643 504 644
rect 498 639 499 643
rect 503 639 504 643
rect 498 638 504 639
rect 534 643 540 644
rect 534 639 535 643
rect 539 639 540 643
rect 534 638 540 639
rect 546 643 552 644
rect 546 639 547 643
rect 551 639 552 643
rect 546 638 552 639
rect 574 643 580 644
rect 574 639 575 643
rect 579 639 580 643
rect 574 638 580 639
rect 594 643 600 644
rect 594 639 595 643
rect 599 639 600 643
rect 594 638 600 639
rect 614 643 620 644
rect 614 639 615 643
rect 619 639 620 643
rect 642 643 648 644
rect 642 639 643 643
rect 647 639 648 643
rect 614 638 620 639
rect 627 638 631 639
rect 642 638 648 639
rect 678 643 684 644
rect 678 639 679 643
rect 683 639 684 643
rect 678 638 684 639
rect 690 643 696 644
rect 690 639 691 643
rect 695 639 696 643
rect 690 638 696 639
rect 702 643 708 644
rect 702 639 703 643
rect 707 639 708 643
rect 702 638 708 639
rect 451 633 455 634
rect 470 635 476 636
rect 274 629 275 633
rect 279 629 280 633
rect 274 628 280 629
rect 378 629 379 633
rect 383 629 384 633
rect 470 631 471 635
rect 475 631 476 635
rect 470 630 476 631
rect 498 633 504 634
rect 547 633 551 634
rect 378 628 384 629
rect 498 629 499 633
rect 503 629 504 633
rect 498 628 504 629
rect 510 631 516 632
rect 174 627 180 628
rect 174 623 175 627
rect 179 623 180 627
rect 174 622 180 623
rect 222 627 228 628
rect 222 623 223 627
rect 227 623 228 627
rect 222 622 228 623
rect 310 627 316 628
rect 310 623 311 627
rect 315 623 316 627
rect 510 627 511 631
rect 515 627 516 631
rect 510 626 516 627
rect 310 622 316 623
rect 110 621 116 622
rect 110 617 111 621
rect 115 617 116 621
rect 110 616 116 617
rect 110 603 116 604
rect 110 599 111 603
rect 115 599 116 603
rect 110 598 116 599
rect 134 603 140 604
rect 134 599 135 603
rect 139 599 140 603
rect 134 598 140 599
rect 112 583 114 598
rect 136 583 138 598
rect 176 596 178 622
rect 182 603 188 604
rect 182 599 183 603
rect 187 599 188 603
rect 182 598 188 599
rect 142 595 148 596
rect 142 591 143 595
rect 147 591 148 595
rect 142 590 148 591
rect 174 595 180 596
rect 174 591 175 595
rect 179 591 180 595
rect 174 590 180 591
rect 111 582 115 583
rect 111 577 115 578
rect 135 582 139 583
rect 135 577 139 578
rect 112 562 114 577
rect 136 562 138 577
rect 110 561 116 562
rect 110 557 111 561
rect 115 557 116 561
rect 110 556 116 557
rect 134 561 140 562
rect 134 557 135 561
rect 139 557 140 561
rect 134 556 140 557
rect 110 543 116 544
rect 110 539 111 543
rect 115 539 116 543
rect 110 538 116 539
rect 112 527 114 538
rect 144 532 146 590
rect 184 583 186 598
rect 224 596 226 622
rect 254 603 260 604
rect 254 599 255 603
rect 259 599 260 603
rect 254 598 260 599
rect 222 595 228 596
rect 222 591 223 595
rect 227 591 228 595
rect 222 590 228 591
rect 256 583 258 598
rect 312 596 314 622
rect 358 603 364 604
rect 358 599 359 603
rect 363 599 364 603
rect 358 598 364 599
rect 478 603 484 604
rect 478 599 479 603
rect 483 599 484 603
rect 478 598 484 599
rect 310 595 316 596
rect 310 591 311 595
rect 315 591 316 595
rect 310 590 316 591
rect 360 583 362 598
rect 480 583 482 598
rect 512 596 514 626
rect 518 623 524 624
rect 518 619 519 623
rect 523 619 524 623
rect 518 618 524 619
rect 520 596 522 618
rect 510 595 516 596
rect 510 591 511 595
rect 515 591 516 595
rect 510 590 516 591
rect 518 595 524 596
rect 518 591 519 595
rect 523 591 524 595
rect 518 590 524 591
rect 183 582 187 583
rect 183 577 187 578
rect 255 582 259 583
rect 255 577 259 578
rect 263 582 267 583
rect 263 577 267 578
rect 351 582 355 583
rect 351 577 355 578
rect 359 582 363 583
rect 359 577 363 578
rect 447 582 451 583
rect 447 577 451 578
rect 479 582 483 583
rect 479 577 483 578
rect 543 582 547 583
rect 543 577 547 578
rect 174 567 180 568
rect 174 563 175 567
rect 179 563 180 567
rect 174 562 180 563
rect 184 562 186 577
rect 222 567 228 568
rect 222 563 223 567
rect 227 563 228 567
rect 222 562 228 563
rect 264 562 266 577
rect 342 567 348 568
rect 342 563 343 567
rect 347 563 348 567
rect 342 562 348 563
rect 352 562 354 577
rect 390 575 396 576
rect 390 571 391 575
rect 395 571 396 575
rect 390 570 396 571
rect 176 532 178 562
rect 182 561 188 562
rect 182 557 183 561
rect 187 557 188 561
rect 182 556 188 557
rect 224 532 226 562
rect 262 561 268 562
rect 262 557 263 561
rect 267 557 268 561
rect 262 556 268 557
rect 344 532 346 562
rect 350 561 356 562
rect 350 557 351 561
rect 355 557 356 561
rect 350 556 356 557
rect 392 540 394 570
rect 438 567 444 568
rect 438 563 439 567
rect 443 563 444 567
rect 438 562 444 563
rect 448 562 450 577
rect 544 562 546 577
rect 576 572 578 638
rect 595 633 599 634
rect 626 633 632 634
rect 643 633 647 634
rect 712 636 714 674
rect 718 673 724 674
rect 718 669 719 673
rect 723 669 724 673
rect 718 668 724 669
rect 774 673 780 674
rect 774 669 775 673
rect 779 669 780 673
rect 774 668 780 669
rect 774 655 780 656
rect 774 651 775 655
rect 779 651 780 655
rect 774 650 780 651
rect 738 643 744 644
rect 738 639 739 643
rect 743 639 744 643
rect 776 639 778 650
rect 738 638 744 639
rect 775 638 779 639
rect 691 633 695 634
rect 710 635 716 636
rect 626 629 627 633
rect 631 629 632 633
rect 710 631 711 635
rect 715 631 716 635
rect 710 630 716 631
rect 738 633 744 634
rect 775 633 779 634
rect 626 628 632 629
rect 738 629 739 633
rect 743 629 744 633
rect 738 628 744 629
rect 776 622 778 633
rect 774 621 780 622
rect 774 617 775 621
rect 779 617 780 621
rect 774 616 780 617
rect 606 603 612 604
rect 606 599 607 603
rect 611 599 612 603
rect 606 598 612 599
rect 718 603 724 604
rect 718 599 719 603
rect 723 599 724 603
rect 718 598 724 599
rect 774 603 780 604
rect 774 599 775 603
rect 779 599 780 603
rect 774 598 780 599
rect 608 583 610 598
rect 720 583 722 598
rect 726 595 732 596
rect 726 591 727 595
rect 731 591 732 595
rect 726 590 732 591
rect 607 582 611 583
rect 607 577 611 578
rect 639 582 643 583
rect 639 577 643 578
rect 719 582 723 583
rect 719 577 723 578
rect 574 571 580 572
rect 574 567 575 571
rect 579 567 580 571
rect 574 566 580 567
rect 640 562 642 577
rect 670 571 676 572
rect 670 567 671 571
rect 675 567 676 571
rect 670 566 676 567
rect 390 539 396 540
rect 390 535 391 539
rect 395 535 396 539
rect 390 534 396 535
rect 440 532 442 562
rect 446 561 452 562
rect 446 557 447 561
rect 451 557 452 561
rect 446 556 452 557
rect 542 561 548 562
rect 542 557 543 561
rect 547 557 548 561
rect 542 556 548 557
rect 638 561 644 562
rect 638 557 639 561
rect 643 557 644 561
rect 638 556 644 557
rect 590 539 596 540
rect 590 535 591 539
rect 595 535 596 539
rect 590 534 596 535
rect 142 531 148 532
rect 142 527 143 531
rect 147 527 148 531
rect 111 526 115 527
rect 142 526 148 527
rect 154 531 160 532
rect 154 527 155 531
rect 159 527 160 531
rect 154 526 160 527
rect 174 531 180 532
rect 174 527 175 531
rect 179 527 180 531
rect 174 526 180 527
rect 202 531 208 532
rect 202 527 203 531
rect 207 527 208 531
rect 222 531 228 532
rect 222 527 223 531
rect 227 527 228 531
rect 282 531 288 532
rect 282 527 283 531
rect 287 527 288 531
rect 342 531 348 532
rect 342 527 343 531
rect 347 527 348 531
rect 202 526 208 527
rect 211 526 215 527
rect 222 526 228 527
rect 267 526 271 527
rect 282 526 288 527
rect 331 526 335 527
rect 342 526 348 527
rect 370 531 376 532
rect 370 527 371 531
rect 375 527 376 531
rect 438 531 444 532
rect 438 527 439 531
rect 443 527 444 531
rect 370 526 376 527
rect 403 526 407 527
rect 438 526 444 527
rect 466 531 472 532
rect 466 527 467 531
rect 471 527 472 531
rect 562 531 568 532
rect 562 527 563 531
rect 567 527 568 531
rect 466 526 472 527
rect 483 526 487 527
rect 562 526 568 527
rect 571 526 575 527
rect 111 521 115 522
rect 155 521 159 522
rect 203 521 207 522
rect 210 521 216 522
rect 112 510 114 521
rect 210 517 211 521
rect 215 517 216 521
rect 266 521 272 522
rect 283 521 287 522
rect 330 521 336 522
rect 371 521 375 522
rect 402 521 408 522
rect 467 521 471 522
rect 482 521 488 522
rect 563 521 567 522
rect 570 521 576 522
rect 210 516 216 517
rect 222 519 228 520
rect 222 515 223 519
rect 227 515 228 519
rect 266 517 267 521
rect 271 517 272 521
rect 266 516 272 517
rect 330 517 331 521
rect 335 517 336 521
rect 330 516 336 517
rect 342 519 348 520
rect 222 514 228 515
rect 342 515 343 519
rect 347 515 348 519
rect 402 517 403 521
rect 407 517 408 521
rect 402 516 408 517
rect 414 519 420 520
rect 342 514 348 515
rect 414 515 415 519
rect 419 515 420 519
rect 482 517 483 521
rect 487 517 488 521
rect 482 516 488 517
rect 494 519 500 520
rect 414 514 420 515
rect 494 515 495 519
rect 499 515 500 519
rect 570 517 571 521
rect 575 517 576 521
rect 570 516 576 517
rect 494 514 500 515
rect 110 509 116 510
rect 110 505 111 509
rect 115 505 116 509
rect 110 504 116 505
rect 110 491 116 492
rect 110 487 111 491
rect 115 487 116 491
rect 110 486 116 487
rect 190 491 196 492
rect 190 487 191 491
rect 195 487 196 491
rect 190 486 196 487
rect 112 471 114 486
rect 192 471 194 486
rect 224 484 226 514
rect 246 491 252 492
rect 246 487 247 491
rect 251 487 252 491
rect 246 486 252 487
rect 310 491 316 492
rect 310 487 311 491
rect 315 487 316 491
rect 310 486 316 487
rect 222 483 228 484
rect 222 479 223 483
rect 227 479 228 483
rect 222 478 228 479
rect 248 471 250 486
rect 312 471 314 486
rect 344 484 346 514
rect 382 491 388 492
rect 382 487 383 491
rect 387 487 388 491
rect 382 486 388 487
rect 342 483 348 484
rect 342 479 343 483
rect 347 479 348 483
rect 342 478 348 479
rect 384 471 386 486
rect 416 484 418 514
rect 462 491 468 492
rect 462 487 463 491
rect 467 487 468 491
rect 462 486 468 487
rect 414 483 420 484
rect 414 479 415 483
rect 419 479 420 483
rect 414 478 420 479
rect 464 471 466 486
rect 496 484 498 514
rect 550 491 556 492
rect 550 487 551 491
rect 555 487 556 491
rect 550 486 556 487
rect 494 483 500 484
rect 494 479 495 483
rect 499 479 500 483
rect 494 478 500 479
rect 502 483 508 484
rect 502 479 503 483
rect 507 479 508 483
rect 502 478 508 479
rect 111 470 115 471
rect 111 465 115 466
rect 191 470 195 471
rect 191 465 195 466
rect 247 470 251 471
rect 247 465 251 466
rect 311 470 315 471
rect 311 465 315 466
rect 351 470 355 471
rect 351 465 355 466
rect 383 470 387 471
rect 383 465 387 466
rect 399 470 403 471
rect 399 465 403 466
rect 447 470 451 471
rect 447 465 451 466
rect 463 470 467 471
rect 463 465 467 466
rect 495 470 499 471
rect 495 465 499 466
rect 112 450 114 465
rect 352 450 354 465
rect 390 455 396 456
rect 390 451 391 455
rect 395 451 396 455
rect 390 450 396 451
rect 400 450 402 465
rect 438 455 444 456
rect 438 451 439 455
rect 443 451 444 455
rect 438 450 444 451
rect 448 450 450 465
rect 486 455 492 456
rect 486 451 487 455
rect 491 451 492 455
rect 486 450 492 451
rect 496 450 498 465
rect 110 449 116 450
rect 110 445 111 449
rect 115 445 116 449
rect 110 444 116 445
rect 350 449 356 450
rect 350 445 351 449
rect 355 445 356 449
rect 350 444 356 445
rect 110 431 116 432
rect 110 427 111 431
rect 115 427 116 431
rect 110 426 116 427
rect 112 411 114 426
rect 392 420 394 450
rect 398 449 404 450
rect 398 445 399 449
rect 403 445 404 449
rect 398 444 404 445
rect 440 420 442 450
rect 446 449 452 450
rect 446 445 447 449
rect 451 445 452 449
rect 446 444 452 445
rect 488 420 490 450
rect 494 449 500 450
rect 494 445 495 449
rect 499 445 500 449
rect 494 444 500 445
rect 504 428 506 478
rect 552 471 554 486
rect 592 484 594 534
rect 658 531 664 532
rect 658 527 659 531
rect 663 527 664 531
rect 672 531 674 566
rect 720 562 722 577
rect 718 561 724 562
rect 718 557 719 561
rect 723 557 724 561
rect 718 556 724 557
rect 728 532 730 590
rect 776 583 778 598
rect 775 582 779 583
rect 775 577 779 578
rect 776 562 778 577
rect 774 561 780 562
rect 774 557 775 561
rect 779 557 780 561
rect 774 556 780 557
rect 774 543 780 544
rect 774 539 775 543
rect 779 539 780 543
rect 774 538 780 539
rect 726 531 732 532
rect 672 529 678 531
rect 658 526 664 527
rect 667 526 671 527
rect 676 524 678 529
rect 726 527 727 531
rect 731 527 732 531
rect 726 526 732 527
rect 738 531 744 532
rect 738 527 739 531
rect 743 527 744 531
rect 776 527 778 538
rect 738 526 744 527
rect 775 526 779 527
rect 674 523 680 524
rect 659 521 663 522
rect 666 521 672 522
rect 666 517 667 521
rect 671 517 672 521
rect 674 519 675 523
rect 679 519 680 523
rect 674 518 680 519
rect 738 521 744 522
rect 775 521 779 522
rect 666 516 672 517
rect 738 517 739 521
rect 743 517 744 521
rect 738 516 744 517
rect 654 515 660 516
rect 654 511 655 515
rect 659 511 660 515
rect 654 510 660 511
rect 776 510 778 521
rect 646 491 652 492
rect 646 487 647 491
rect 651 487 652 491
rect 646 486 652 487
rect 590 483 596 484
rect 590 479 591 483
rect 595 479 596 483
rect 590 478 596 479
rect 648 471 650 486
rect 543 470 547 471
rect 543 465 547 466
rect 551 470 555 471
rect 551 465 555 466
rect 599 470 603 471
rect 599 465 603 466
rect 647 470 651 471
rect 647 465 651 466
rect 534 455 540 456
rect 534 451 535 455
rect 539 451 540 455
rect 534 450 540 451
rect 544 450 546 465
rect 574 459 580 460
rect 574 455 575 459
rect 579 455 580 459
rect 574 454 580 455
rect 586 455 592 456
rect 502 427 508 428
rect 502 423 503 427
rect 507 423 508 427
rect 502 422 508 423
rect 536 420 538 450
rect 542 449 548 450
rect 542 445 543 449
rect 547 445 548 449
rect 542 444 548 445
rect 576 420 578 454
rect 586 451 587 455
rect 591 451 592 455
rect 586 450 592 451
rect 600 450 602 465
rect 656 460 658 510
rect 774 509 780 510
rect 774 505 775 509
rect 779 505 780 509
rect 774 504 780 505
rect 718 491 724 492
rect 718 487 719 491
rect 723 487 724 491
rect 718 486 724 487
rect 774 491 780 492
rect 774 487 775 491
rect 779 487 780 491
rect 774 486 780 487
rect 720 471 722 486
rect 726 483 732 484
rect 726 479 727 483
rect 731 479 732 483
rect 726 478 732 479
rect 663 470 667 471
rect 663 465 667 466
rect 719 470 723 471
rect 719 465 723 466
rect 654 459 660 460
rect 654 455 655 459
rect 659 455 660 459
rect 654 454 660 455
rect 664 450 666 465
rect 710 455 716 456
rect 710 451 711 455
rect 715 451 716 455
rect 710 450 716 451
rect 720 450 722 465
rect 370 419 376 420
rect 370 415 371 419
rect 375 415 376 419
rect 370 414 376 415
rect 390 419 396 420
rect 390 415 391 419
rect 395 415 396 419
rect 390 414 396 415
rect 418 419 424 420
rect 418 415 419 419
rect 423 415 424 419
rect 418 414 424 415
rect 438 419 444 420
rect 438 415 439 419
rect 443 415 444 419
rect 438 414 444 415
rect 466 419 472 420
rect 466 415 467 419
rect 471 415 472 419
rect 466 414 472 415
rect 486 419 492 420
rect 486 415 487 419
rect 491 415 492 419
rect 486 414 492 415
rect 514 419 520 420
rect 514 415 515 419
rect 519 415 520 419
rect 514 414 520 415
rect 534 419 540 420
rect 534 415 535 419
rect 539 415 540 419
rect 534 414 540 415
rect 562 419 568 420
rect 562 415 563 419
rect 567 415 568 419
rect 562 414 568 415
rect 574 419 580 420
rect 574 415 575 419
rect 579 415 580 419
rect 574 414 580 415
rect 372 411 374 414
rect 420 411 422 414
rect 468 411 470 414
rect 516 411 518 414
rect 564 411 566 414
rect 111 410 115 411
rect 339 410 343 411
rect 371 410 375 411
rect 387 410 391 411
rect 419 410 423 411
rect 435 410 439 411
rect 467 410 471 411
rect 483 410 487 411
rect 515 410 519 411
rect 539 410 543 411
rect 563 410 567 411
rect 588 408 590 450
rect 598 449 604 450
rect 598 445 599 449
rect 603 445 604 449
rect 598 444 604 445
rect 662 449 668 450
rect 662 445 663 449
rect 667 445 668 449
rect 662 444 668 445
rect 618 419 624 420
rect 618 415 619 419
rect 623 415 624 419
rect 618 414 624 415
rect 658 419 664 420
rect 658 415 659 419
rect 663 415 664 419
rect 658 414 664 415
rect 682 419 688 420
rect 682 415 683 419
rect 687 415 688 419
rect 682 414 688 415
rect 620 411 622 414
rect 603 410 607 411
rect 111 405 115 406
rect 338 405 344 406
rect 371 405 375 406
rect 386 405 392 406
rect 419 405 423 406
rect 434 405 440 406
rect 467 405 471 406
rect 482 405 488 406
rect 515 405 519 406
rect 538 405 544 406
rect 563 405 567 406
rect 586 407 592 408
rect 112 394 114 405
rect 338 401 339 405
rect 343 401 344 405
rect 338 400 344 401
rect 350 403 356 404
rect 350 399 351 403
rect 355 399 356 403
rect 386 401 387 405
rect 391 401 392 405
rect 386 400 392 401
rect 398 403 404 404
rect 350 398 356 399
rect 398 399 399 403
rect 403 399 404 403
rect 434 401 435 405
rect 439 401 440 405
rect 434 400 440 401
rect 482 401 483 405
rect 487 401 488 405
rect 482 400 488 401
rect 538 401 539 405
rect 543 401 544 405
rect 586 403 587 407
rect 591 403 592 407
rect 619 410 623 411
rect 586 402 592 403
rect 602 405 608 406
rect 619 405 623 406
rect 538 400 544 401
rect 602 401 603 405
rect 607 401 608 405
rect 602 400 608 401
rect 638 403 644 404
rect 398 398 404 399
rect 502 399 508 400
rect 110 393 116 394
rect 110 389 111 393
rect 115 389 116 393
rect 110 388 116 389
rect 110 375 116 376
rect 110 371 111 375
rect 115 371 116 375
rect 110 370 116 371
rect 318 375 324 376
rect 318 371 319 375
rect 323 371 324 375
rect 318 370 324 371
rect 112 347 114 370
rect 320 347 322 370
rect 352 368 354 398
rect 366 375 372 376
rect 366 371 367 375
rect 371 371 372 375
rect 366 370 372 371
rect 350 367 356 368
rect 350 363 351 367
rect 355 363 356 367
rect 350 362 356 363
rect 368 347 370 370
rect 400 368 402 398
rect 454 395 460 396
rect 454 391 455 395
rect 459 391 460 395
rect 502 395 503 399
rect 507 395 508 399
rect 502 394 508 395
rect 558 399 564 400
rect 558 395 559 399
rect 563 395 564 399
rect 638 399 639 403
rect 643 399 644 403
rect 638 398 644 399
rect 558 394 564 395
rect 454 390 460 391
rect 414 375 420 376
rect 414 371 415 375
rect 419 371 420 375
rect 414 370 420 371
rect 398 367 404 368
rect 398 363 399 367
rect 403 363 404 367
rect 398 362 404 363
rect 416 347 418 370
rect 456 368 458 390
rect 462 375 468 376
rect 462 371 463 375
rect 467 371 468 375
rect 462 370 468 371
rect 430 367 436 368
rect 430 363 431 367
rect 435 363 436 367
rect 430 362 436 363
rect 454 367 460 368
rect 454 363 455 367
rect 459 363 460 367
rect 454 362 460 363
rect 111 346 115 347
rect 111 341 115 342
rect 135 346 139 347
rect 135 341 139 342
rect 199 346 203 347
rect 199 341 203 342
rect 271 346 275 347
rect 271 341 275 342
rect 319 346 323 347
rect 319 341 323 342
rect 343 346 347 347
rect 343 341 347 342
rect 367 346 371 347
rect 367 341 371 342
rect 415 346 419 347
rect 415 341 419 342
rect 423 346 427 347
rect 423 341 427 342
rect 112 326 114 341
rect 126 331 132 332
rect 126 327 127 331
rect 131 327 132 331
rect 126 326 132 327
rect 136 326 138 341
rect 174 331 180 332
rect 174 327 175 331
rect 179 327 180 331
rect 174 326 180 327
rect 200 326 202 341
rect 238 331 244 332
rect 238 327 239 331
rect 243 327 244 331
rect 238 326 244 327
rect 272 326 274 341
rect 310 331 316 332
rect 310 327 311 331
rect 315 327 316 331
rect 310 326 316 327
rect 344 326 346 341
rect 424 326 426 341
rect 110 325 116 326
rect 110 321 111 325
rect 115 321 116 325
rect 110 320 116 321
rect 110 307 116 308
rect 110 303 111 307
rect 115 303 116 307
rect 110 302 116 303
rect 112 283 114 302
rect 111 282 115 283
rect 128 280 130 326
rect 134 325 140 326
rect 134 321 135 325
rect 139 321 140 325
rect 134 320 140 321
rect 176 304 178 326
rect 198 325 204 326
rect 198 321 199 325
rect 203 321 204 325
rect 198 320 204 321
rect 240 304 242 326
rect 270 325 276 326
rect 270 321 271 325
rect 275 321 276 325
rect 270 320 276 321
rect 312 304 314 326
rect 342 325 348 326
rect 342 321 343 325
rect 347 321 348 325
rect 342 320 348 321
rect 422 325 428 326
rect 422 321 423 325
rect 427 321 428 325
rect 422 320 428 321
rect 174 303 180 304
rect 174 299 175 303
rect 179 299 180 303
rect 174 298 180 299
rect 238 303 244 304
rect 238 299 239 303
rect 243 299 244 303
rect 238 298 244 299
rect 310 303 316 304
rect 310 299 311 303
rect 315 299 316 303
rect 310 298 316 299
rect 432 296 434 362
rect 464 347 466 370
rect 504 368 506 394
rect 518 375 524 376
rect 518 371 519 375
rect 523 371 524 375
rect 518 370 524 371
rect 502 367 508 368
rect 502 363 503 367
rect 507 363 508 367
rect 502 362 508 363
rect 520 347 522 370
rect 560 368 562 394
rect 582 375 588 376
rect 582 371 583 375
rect 587 371 588 375
rect 582 370 588 371
rect 558 367 564 368
rect 558 363 559 367
rect 563 363 564 367
rect 558 362 564 363
rect 584 347 586 370
rect 463 346 467 347
rect 463 341 467 342
rect 511 346 515 347
rect 511 341 515 342
rect 519 346 523 347
rect 519 341 523 342
rect 583 346 587 347
rect 583 341 587 342
rect 607 346 611 347
rect 607 341 611 342
rect 512 326 514 341
rect 598 331 604 332
rect 598 327 599 331
rect 603 327 604 331
rect 598 326 604 327
rect 608 326 610 341
rect 640 336 642 398
rect 646 375 652 376
rect 646 371 647 375
rect 651 371 652 375
rect 646 370 652 371
rect 648 347 650 370
rect 660 368 662 414
rect 684 411 686 414
rect 667 410 671 411
rect 683 410 687 411
rect 712 408 714 450
rect 718 449 724 450
rect 718 445 719 449
rect 723 445 724 449
rect 718 444 724 445
rect 728 420 730 478
rect 776 471 778 486
rect 775 470 779 471
rect 775 465 779 466
rect 776 450 778 465
rect 774 449 780 450
rect 774 445 775 449
rect 779 445 780 449
rect 774 444 780 445
rect 774 431 780 432
rect 774 427 775 431
rect 779 427 780 431
rect 774 426 780 427
rect 726 419 732 420
rect 726 415 727 419
rect 731 415 732 419
rect 726 414 732 415
rect 738 419 744 420
rect 738 415 739 419
rect 743 415 744 419
rect 738 414 744 415
rect 740 411 742 414
rect 776 411 778 426
rect 739 410 743 411
rect 666 405 672 406
rect 683 405 687 406
rect 710 407 716 408
rect 666 401 667 405
rect 671 401 672 405
rect 710 403 711 407
rect 715 403 716 407
rect 775 410 779 411
rect 710 402 716 403
rect 738 405 744 406
rect 775 405 779 406
rect 666 400 672 401
rect 738 401 739 405
rect 743 401 744 405
rect 738 400 744 401
rect 776 394 778 405
rect 774 393 780 394
rect 774 389 775 393
rect 779 389 780 393
rect 774 388 780 389
rect 718 375 724 376
rect 718 371 719 375
rect 723 371 724 375
rect 718 370 724 371
rect 774 375 780 376
rect 774 371 775 375
rect 779 371 780 375
rect 774 370 780 371
rect 658 367 664 368
rect 658 363 659 367
rect 663 363 664 367
rect 658 362 664 363
rect 710 367 716 368
rect 710 363 711 367
rect 715 363 716 367
rect 710 362 716 363
rect 647 346 651 347
rect 647 341 651 342
rect 703 346 707 347
rect 703 341 707 342
rect 638 335 644 336
rect 638 331 639 335
rect 643 331 644 335
rect 638 330 644 331
rect 694 331 700 332
rect 694 327 695 331
rect 699 327 700 331
rect 694 326 700 327
rect 704 326 706 341
rect 510 325 516 326
rect 510 321 511 325
rect 515 321 516 325
rect 510 320 516 321
rect 600 296 602 326
rect 606 325 612 326
rect 606 321 607 325
rect 611 321 612 325
rect 606 320 612 321
rect 154 295 160 296
rect 154 291 155 295
rect 159 291 160 295
rect 154 290 160 291
rect 218 295 224 296
rect 218 291 219 295
rect 223 291 224 295
rect 218 290 224 291
rect 290 295 296 296
rect 290 291 291 295
rect 295 291 296 295
rect 290 290 296 291
rect 362 295 368 296
rect 362 291 363 295
rect 367 291 368 295
rect 362 290 368 291
rect 430 295 436 296
rect 430 291 431 295
rect 435 291 436 295
rect 430 290 436 291
rect 442 295 448 296
rect 442 291 443 295
rect 447 291 448 295
rect 442 290 448 291
rect 510 295 516 296
rect 510 291 511 295
rect 515 291 516 295
rect 510 290 516 291
rect 530 295 536 296
rect 530 291 531 295
rect 535 291 536 295
rect 530 290 536 291
rect 598 295 604 296
rect 598 291 599 295
rect 603 291 604 295
rect 598 290 604 291
rect 626 295 632 296
rect 626 291 627 295
rect 631 291 632 295
rect 626 290 632 291
rect 156 283 158 290
rect 220 283 222 290
rect 292 283 294 290
rect 364 283 366 290
rect 444 283 446 290
rect 155 282 159 283
rect 111 277 115 278
rect 126 279 132 280
rect 112 266 114 277
rect 126 275 127 279
rect 131 275 132 279
rect 211 282 215 283
rect 219 282 223 283
rect 126 274 132 275
rect 154 277 160 278
rect 154 273 155 277
rect 159 273 160 277
rect 210 277 216 278
rect 219 277 223 278
rect 291 282 295 283
rect 299 282 303 283
rect 363 282 367 283
rect 387 282 391 283
rect 443 282 447 283
rect 475 282 479 283
rect 291 277 295 278
rect 298 277 304 278
rect 363 277 367 278
rect 386 277 392 278
rect 443 277 447 278
rect 474 277 480 278
rect 154 272 160 273
rect 166 275 172 276
rect 166 271 167 275
rect 171 271 172 275
rect 210 273 211 277
rect 215 273 216 277
rect 210 272 216 273
rect 234 275 240 276
rect 166 270 172 271
rect 234 271 235 275
rect 239 271 240 275
rect 298 273 299 277
rect 303 273 304 277
rect 298 272 304 273
rect 310 275 316 276
rect 234 270 240 271
rect 310 271 311 275
rect 315 271 316 275
rect 386 273 387 277
rect 391 273 392 277
rect 386 272 392 273
rect 474 273 475 277
rect 479 273 480 277
rect 474 272 480 273
rect 486 275 492 276
rect 310 270 316 271
rect 486 271 487 275
rect 491 271 492 275
rect 486 270 492 271
rect 110 265 116 266
rect 110 261 111 265
rect 115 261 116 265
rect 110 260 116 261
rect 110 247 116 248
rect 110 243 111 247
rect 115 243 116 247
rect 110 242 116 243
rect 134 247 140 248
rect 134 243 135 247
rect 139 243 140 247
rect 134 242 140 243
rect 112 219 114 242
rect 136 219 138 242
rect 168 240 170 270
rect 190 247 196 248
rect 190 243 191 247
rect 195 243 196 247
rect 190 242 196 243
rect 166 239 172 240
rect 166 235 167 239
rect 171 235 172 239
rect 166 234 172 235
rect 192 219 194 242
rect 236 240 238 270
rect 278 247 284 248
rect 278 243 279 247
rect 283 243 284 247
rect 278 242 284 243
rect 234 239 240 240
rect 234 235 235 239
rect 239 235 240 239
rect 234 234 240 235
rect 280 219 282 242
rect 312 240 314 270
rect 366 247 372 248
rect 366 243 367 247
rect 371 243 372 247
rect 366 242 372 243
rect 454 247 460 248
rect 454 243 455 247
rect 459 243 460 247
rect 454 242 460 243
rect 310 239 316 240
rect 310 235 311 239
rect 315 235 316 239
rect 310 234 316 235
rect 368 219 370 242
rect 374 239 380 240
rect 374 235 375 239
rect 379 235 380 239
rect 374 234 380 235
rect 111 218 115 219
rect 111 213 115 214
rect 135 218 139 219
rect 135 213 139 214
rect 191 218 195 219
rect 191 213 195 214
rect 279 218 283 219
rect 279 213 283 214
rect 367 218 371 219
rect 367 213 371 214
rect 112 198 114 213
rect 182 203 188 204
rect 182 199 183 203
rect 187 199 188 203
rect 182 198 188 199
rect 192 198 194 213
rect 280 198 282 213
rect 326 203 332 204
rect 326 199 327 203
rect 331 199 332 203
rect 326 198 332 199
rect 368 198 370 213
rect 110 197 116 198
rect 110 193 111 197
rect 115 193 116 197
rect 110 192 116 193
rect 110 179 116 180
rect 110 175 111 179
rect 115 175 116 179
rect 110 174 116 175
rect 112 155 114 174
rect 111 154 115 155
rect 184 152 186 198
rect 190 197 196 198
rect 190 193 191 197
rect 195 193 196 197
rect 190 192 196 193
rect 278 197 284 198
rect 278 193 279 197
rect 283 193 284 197
rect 278 192 284 193
rect 328 176 330 198
rect 366 197 372 198
rect 366 193 367 197
rect 371 193 372 197
rect 366 192 372 193
rect 326 175 332 176
rect 326 171 327 175
rect 331 171 332 175
rect 326 170 332 171
rect 376 168 378 234
rect 456 219 458 242
rect 488 240 490 270
rect 512 240 514 290
rect 532 283 534 290
rect 628 283 630 290
rect 531 282 535 283
rect 563 282 567 283
rect 627 282 631 283
rect 659 282 663 283
rect 696 280 698 326
rect 702 325 708 326
rect 702 321 703 325
rect 707 321 708 325
rect 702 320 708 321
rect 712 296 714 362
rect 720 347 722 370
rect 776 347 778 370
rect 719 346 723 347
rect 719 341 723 342
rect 775 346 779 347
rect 775 341 779 342
rect 776 326 778 341
rect 774 325 780 326
rect 774 321 775 325
rect 779 321 780 325
rect 774 320 780 321
rect 774 307 780 308
rect 774 303 775 307
rect 779 303 780 307
rect 774 302 780 303
rect 710 295 716 296
rect 710 291 711 295
rect 715 291 716 295
rect 710 290 716 291
rect 722 295 728 296
rect 722 291 723 295
rect 727 291 728 295
rect 722 290 728 291
rect 724 283 726 290
rect 776 283 778 302
rect 723 282 727 283
rect 694 279 700 280
rect 531 277 535 278
rect 562 277 568 278
rect 627 277 631 278
rect 658 277 664 278
rect 562 273 563 277
rect 567 273 568 277
rect 562 272 568 273
rect 658 273 659 277
rect 663 273 664 277
rect 694 275 695 279
rect 699 275 700 279
rect 739 282 743 283
rect 775 282 779 283
rect 723 277 727 278
rect 738 277 744 278
rect 775 277 779 278
rect 694 274 700 275
rect 658 272 664 273
rect 738 273 739 277
rect 743 273 744 277
rect 738 272 744 273
rect 682 271 688 272
rect 682 267 683 271
rect 687 267 688 271
rect 682 266 688 267
rect 776 266 778 277
rect 542 247 548 248
rect 542 243 543 247
rect 547 243 548 247
rect 542 242 548 243
rect 638 247 644 248
rect 638 243 639 247
rect 643 243 644 247
rect 638 242 644 243
rect 486 239 492 240
rect 486 235 487 239
rect 491 235 492 239
rect 486 234 492 235
rect 510 239 516 240
rect 510 235 511 239
rect 515 235 516 239
rect 510 234 516 235
rect 544 219 546 242
rect 640 219 642 242
rect 684 240 686 266
rect 774 265 780 266
rect 774 261 775 265
rect 779 261 780 265
rect 774 260 780 261
rect 718 247 724 248
rect 718 243 719 247
rect 723 243 724 247
rect 718 242 724 243
rect 774 247 780 248
rect 774 243 775 247
rect 779 243 780 247
rect 774 242 780 243
rect 654 239 660 240
rect 654 235 655 239
rect 659 235 660 239
rect 654 234 660 235
rect 682 239 688 240
rect 682 235 683 239
rect 687 235 688 239
rect 682 234 688 235
rect 455 218 459 219
rect 455 213 459 214
rect 543 218 547 219
rect 543 213 547 214
rect 551 218 555 219
rect 551 213 555 214
rect 639 218 643 219
rect 639 213 643 214
rect 647 218 651 219
rect 647 213 651 214
rect 456 198 458 213
rect 552 198 554 213
rect 648 198 650 213
rect 454 197 460 198
rect 454 193 455 197
rect 459 193 460 197
rect 454 192 460 193
rect 550 197 556 198
rect 550 193 551 197
rect 555 193 556 197
rect 550 192 556 193
rect 646 197 652 198
rect 646 193 647 197
rect 651 193 652 197
rect 646 192 652 193
rect 656 168 658 234
rect 720 219 722 242
rect 776 219 778 242
rect 719 218 723 219
rect 719 213 723 214
rect 775 218 779 219
rect 775 213 779 214
rect 702 203 708 204
rect 702 199 703 203
rect 707 199 708 203
rect 702 198 708 199
rect 710 203 716 204
rect 710 199 711 203
rect 715 199 716 203
rect 710 198 716 199
rect 720 198 722 213
rect 776 198 778 213
rect 704 168 706 198
rect 210 167 216 168
rect 210 163 211 167
rect 215 163 216 167
rect 210 162 216 163
rect 298 167 304 168
rect 298 163 299 167
rect 303 163 304 167
rect 298 162 304 163
rect 374 167 380 168
rect 374 163 375 167
rect 379 163 380 167
rect 374 162 380 163
rect 386 167 392 168
rect 386 163 387 167
rect 391 163 392 167
rect 386 162 392 163
rect 474 167 480 168
rect 474 163 475 167
rect 479 163 480 167
rect 474 162 480 163
rect 570 167 576 168
rect 570 163 571 167
rect 575 163 576 167
rect 570 162 576 163
rect 654 167 660 168
rect 654 163 655 167
rect 659 163 660 167
rect 654 162 660 163
rect 666 167 672 168
rect 666 163 667 167
rect 671 163 672 167
rect 666 162 672 163
rect 702 167 708 168
rect 702 163 703 167
rect 707 163 708 167
rect 702 162 708 163
rect 212 155 214 162
rect 300 155 302 162
rect 388 155 390 162
rect 476 155 478 162
rect 572 155 574 162
rect 668 155 670 162
rect 211 154 215 155
rect 111 149 115 150
rect 182 151 188 152
rect 112 138 114 149
rect 182 147 183 151
rect 187 147 188 151
rect 259 154 263 155
rect 299 154 303 155
rect 307 154 311 155
rect 355 154 359 155
rect 387 154 391 155
rect 403 154 407 155
rect 451 154 455 155
rect 475 154 479 155
rect 499 154 503 155
rect 547 154 551 155
rect 571 154 575 155
rect 595 154 599 155
rect 643 154 647 155
rect 667 154 671 155
rect 691 154 695 155
rect 712 152 714 198
rect 718 197 724 198
rect 718 193 719 197
rect 723 193 724 197
rect 718 192 724 193
rect 774 197 780 198
rect 774 193 775 197
rect 779 193 780 197
rect 774 192 780 193
rect 774 179 780 180
rect 774 175 775 179
rect 779 175 780 179
rect 774 174 780 175
rect 738 167 744 168
rect 738 163 739 167
rect 743 163 744 167
rect 738 162 744 163
rect 740 155 742 162
rect 776 155 778 174
rect 739 154 743 155
rect 710 151 716 152
rect 182 146 188 147
rect 210 149 216 150
rect 210 145 211 149
rect 215 145 216 149
rect 258 149 264 150
rect 299 149 303 150
rect 306 149 312 150
rect 210 144 216 145
rect 222 147 228 148
rect 222 143 223 147
rect 227 143 228 147
rect 258 145 259 149
rect 263 145 264 149
rect 258 144 264 145
rect 270 147 276 148
rect 222 142 228 143
rect 270 143 271 147
rect 275 143 276 147
rect 306 145 307 149
rect 311 145 312 149
rect 354 149 360 150
rect 387 149 391 150
rect 402 149 408 150
rect 306 144 312 145
rect 318 147 324 148
rect 270 142 276 143
rect 318 143 319 147
rect 323 143 324 147
rect 354 145 355 149
rect 359 145 360 149
rect 354 144 360 145
rect 366 147 372 148
rect 318 142 324 143
rect 366 143 367 147
rect 371 143 372 147
rect 402 145 403 149
rect 407 145 408 149
rect 450 149 456 150
rect 475 149 479 150
rect 498 149 504 150
rect 402 144 408 145
rect 414 147 420 148
rect 366 142 372 143
rect 414 143 415 147
rect 419 143 420 147
rect 450 145 451 149
rect 455 145 456 149
rect 450 144 456 145
rect 462 147 468 148
rect 414 142 420 143
rect 462 143 463 147
rect 467 143 468 147
rect 498 145 499 149
rect 503 145 504 149
rect 546 149 552 150
rect 571 149 575 150
rect 594 149 600 150
rect 498 144 504 145
rect 510 147 516 148
rect 462 142 468 143
rect 510 143 511 147
rect 515 143 516 147
rect 546 145 547 149
rect 551 145 552 149
rect 546 144 552 145
rect 558 147 564 148
rect 510 142 516 143
rect 558 143 559 147
rect 563 143 564 147
rect 594 145 595 149
rect 599 145 600 149
rect 594 144 600 145
rect 642 149 648 150
rect 667 149 671 150
rect 690 149 696 150
rect 642 145 643 149
rect 647 145 648 149
rect 642 144 648 145
rect 690 145 691 149
rect 695 145 696 149
rect 710 147 711 151
rect 715 147 716 151
rect 775 154 779 155
rect 710 146 716 147
rect 738 149 744 150
rect 775 149 779 150
rect 690 144 696 145
rect 738 145 739 149
rect 743 145 744 149
rect 738 144 744 145
rect 558 142 564 143
rect 662 143 668 144
rect 110 137 116 138
rect 110 133 111 137
rect 115 133 116 137
rect 110 132 116 133
rect 110 119 116 120
rect 110 115 111 119
rect 115 115 116 119
rect 110 114 116 115
rect 190 119 196 120
rect 190 115 191 119
rect 195 115 196 119
rect 190 114 196 115
rect 112 99 114 114
rect 192 99 194 114
rect 224 112 226 142
rect 238 119 244 120
rect 238 115 239 119
rect 243 115 244 119
rect 238 114 244 115
rect 222 111 228 112
rect 222 107 223 111
rect 227 107 228 111
rect 222 106 228 107
rect 240 99 242 114
rect 272 112 274 142
rect 286 119 292 120
rect 286 115 287 119
rect 291 115 292 119
rect 286 114 292 115
rect 270 111 276 112
rect 270 107 271 111
rect 275 107 276 111
rect 270 106 276 107
rect 288 99 290 114
rect 320 112 322 142
rect 334 119 340 120
rect 334 115 335 119
rect 339 115 340 119
rect 334 114 340 115
rect 318 111 324 112
rect 318 107 319 111
rect 323 107 324 111
rect 318 106 324 107
rect 336 99 338 114
rect 368 112 370 142
rect 382 119 388 120
rect 382 115 383 119
rect 387 115 388 119
rect 382 114 388 115
rect 366 111 372 112
rect 366 107 367 111
rect 371 107 372 111
rect 366 106 372 107
rect 384 99 386 114
rect 416 112 418 142
rect 430 119 436 120
rect 430 115 431 119
rect 435 115 436 119
rect 430 114 436 115
rect 414 111 420 112
rect 414 107 415 111
rect 419 107 420 111
rect 414 106 420 107
rect 432 99 434 114
rect 464 112 466 142
rect 478 119 484 120
rect 478 115 479 119
rect 483 115 484 119
rect 478 114 484 115
rect 462 111 468 112
rect 462 107 463 111
rect 467 107 468 111
rect 462 106 468 107
rect 480 99 482 114
rect 512 112 514 142
rect 526 119 532 120
rect 526 115 527 119
rect 531 115 532 119
rect 526 114 532 115
rect 510 111 516 112
rect 510 107 511 111
rect 515 107 516 111
rect 510 106 516 107
rect 528 99 530 114
rect 560 112 562 142
rect 662 139 663 143
rect 667 139 668 143
rect 662 138 668 139
rect 710 143 716 144
rect 710 139 711 143
rect 715 139 716 143
rect 710 138 716 139
rect 776 138 778 149
rect 574 119 580 120
rect 574 115 575 119
rect 579 115 580 119
rect 574 114 580 115
rect 622 119 628 120
rect 622 115 623 119
rect 627 115 628 119
rect 622 114 628 115
rect 558 111 564 112
rect 558 107 559 111
rect 563 107 564 111
rect 558 106 564 107
rect 576 99 578 114
rect 624 99 626 114
rect 664 112 666 138
rect 670 119 676 120
rect 670 115 671 119
rect 675 115 676 119
rect 670 114 676 115
rect 662 111 668 112
rect 662 107 663 111
rect 667 107 668 111
rect 662 106 668 107
rect 672 99 674 114
rect 712 112 714 138
rect 774 137 780 138
rect 774 133 775 137
rect 779 133 780 137
rect 774 132 780 133
rect 718 119 724 120
rect 718 115 719 119
rect 723 115 724 119
rect 718 114 724 115
rect 774 119 780 120
rect 774 115 775 119
rect 779 115 780 119
rect 774 114 780 115
rect 710 111 716 112
rect 710 107 711 111
rect 715 107 716 111
rect 710 106 716 107
rect 720 99 722 114
rect 776 99 778 114
rect 111 98 115 99
rect 111 93 115 94
rect 191 98 195 99
rect 191 93 195 94
rect 239 98 243 99
rect 239 93 243 94
rect 287 98 291 99
rect 287 93 291 94
rect 335 98 339 99
rect 335 93 339 94
rect 383 98 387 99
rect 383 93 387 94
rect 431 98 435 99
rect 431 93 435 94
rect 479 98 483 99
rect 479 93 483 94
rect 527 98 531 99
rect 527 93 531 94
rect 575 98 579 99
rect 575 93 579 94
rect 623 98 627 99
rect 623 93 627 94
rect 671 98 675 99
rect 671 93 675 94
rect 719 98 723 99
rect 719 93 723 94
rect 775 98 779 99
rect 775 93 779 94
<< m4c >>
rect 111 858 115 862
rect 155 858 159 862
rect 203 858 207 862
rect 251 858 255 862
rect 775 858 779 862
rect 111 802 115 806
rect 135 802 139 806
rect 183 802 187 806
rect 231 802 235 806
rect 279 802 283 806
rect 327 802 331 806
rect 375 802 379 806
rect 775 802 779 806
rect 111 746 115 750
rect 155 746 159 750
rect 203 746 207 750
rect 251 746 255 750
rect 291 746 295 750
rect 299 746 303 750
rect 339 746 343 750
rect 347 746 351 750
rect 387 746 391 750
rect 395 746 399 750
rect 443 746 447 750
rect 507 746 511 750
rect 579 746 583 750
rect 659 746 663 750
rect 739 746 743 750
rect 775 746 779 750
rect 111 690 115 694
rect 271 690 275 694
rect 319 690 323 694
rect 335 690 339 694
rect 367 690 371 694
rect 383 690 387 694
rect 423 690 427 694
rect 431 690 435 694
rect 479 690 483 694
rect 487 690 491 694
rect 527 690 531 694
rect 111 634 115 638
rect 155 634 159 638
rect 203 634 207 638
rect 275 634 279 638
rect 355 634 359 638
rect 379 634 383 638
rect 403 634 407 638
rect 451 634 455 638
rect 559 690 563 694
rect 575 690 579 694
rect 623 690 627 694
rect 639 690 643 694
rect 671 690 675 694
rect 719 690 723 694
rect 775 690 779 694
rect 499 634 503 638
rect 547 634 551 638
rect 111 578 115 582
rect 135 578 139 582
rect 183 578 187 582
rect 255 578 259 582
rect 263 578 267 582
rect 351 578 355 582
rect 359 578 363 582
rect 447 578 451 582
rect 479 578 483 582
rect 543 578 547 582
rect 595 634 599 638
rect 627 634 631 638
rect 643 634 647 638
rect 691 634 695 638
rect 739 634 743 638
rect 775 634 779 638
rect 607 578 611 582
rect 639 578 643 582
rect 719 578 723 582
rect 111 522 115 526
rect 155 522 159 526
rect 203 522 207 526
rect 211 522 215 526
rect 267 522 271 526
rect 283 522 287 526
rect 331 522 335 526
rect 371 522 375 526
rect 403 522 407 526
rect 467 522 471 526
rect 483 522 487 526
rect 563 522 567 526
rect 571 522 575 526
rect 111 466 115 470
rect 191 466 195 470
rect 247 466 251 470
rect 311 466 315 470
rect 351 466 355 470
rect 383 466 387 470
rect 399 466 403 470
rect 447 466 451 470
rect 463 466 467 470
rect 495 466 499 470
rect 775 578 779 582
rect 659 522 663 526
rect 667 522 671 526
rect 739 522 743 526
rect 775 522 779 526
rect 543 466 547 470
rect 551 466 555 470
rect 599 466 603 470
rect 647 466 651 470
rect 663 466 667 470
rect 719 466 723 470
rect 111 406 115 410
rect 339 406 343 410
rect 371 406 375 410
rect 387 406 391 410
rect 419 406 423 410
rect 435 406 439 410
rect 467 406 471 410
rect 483 406 487 410
rect 515 406 519 410
rect 539 406 543 410
rect 563 406 567 410
rect 603 406 607 410
rect 619 406 623 410
rect 111 342 115 346
rect 135 342 139 346
rect 199 342 203 346
rect 271 342 275 346
rect 319 342 323 346
rect 343 342 347 346
rect 367 342 371 346
rect 415 342 419 346
rect 423 342 427 346
rect 111 278 115 282
rect 463 342 467 346
rect 511 342 515 346
rect 519 342 523 346
rect 583 342 587 346
rect 607 342 611 346
rect 667 406 671 410
rect 683 406 687 410
rect 775 466 779 470
rect 739 406 743 410
rect 775 406 779 410
rect 647 342 651 346
rect 703 342 707 346
rect 155 278 159 282
rect 211 278 215 282
rect 219 278 223 282
rect 291 278 295 282
rect 299 278 303 282
rect 363 278 367 282
rect 387 278 391 282
rect 443 278 447 282
rect 475 278 479 282
rect 111 214 115 218
rect 135 214 139 218
rect 191 214 195 218
rect 279 214 283 218
rect 367 214 371 218
rect 111 150 115 154
rect 531 278 535 282
rect 563 278 567 282
rect 627 278 631 282
rect 659 278 663 282
rect 719 342 723 346
rect 775 342 779 346
rect 723 278 727 282
rect 739 278 743 282
rect 775 278 779 282
rect 455 214 459 218
rect 543 214 547 218
rect 551 214 555 218
rect 639 214 643 218
rect 647 214 651 218
rect 719 214 723 218
rect 775 214 779 218
rect 211 150 215 154
rect 259 150 263 154
rect 299 150 303 154
rect 307 150 311 154
rect 355 150 359 154
rect 387 150 391 154
rect 403 150 407 154
rect 451 150 455 154
rect 475 150 479 154
rect 499 150 503 154
rect 547 150 551 154
rect 571 150 575 154
rect 595 150 599 154
rect 643 150 647 154
rect 667 150 671 154
rect 691 150 695 154
rect 739 150 743 154
rect 775 150 779 154
rect 111 94 115 98
rect 191 94 195 98
rect 239 94 243 98
rect 287 94 291 98
rect 335 94 339 98
rect 383 94 387 98
rect 431 94 435 98
rect 479 94 483 98
rect 527 94 531 98
rect 575 94 579 98
rect 623 94 627 98
rect 671 94 675 98
rect 719 94 723 98
rect 775 94 779 98
<< m4 >>
rect 96 857 97 863
rect 103 862 811 863
rect 103 858 111 862
rect 115 858 155 862
rect 159 858 203 862
rect 207 858 251 862
rect 255 858 775 862
rect 779 858 811 862
rect 103 857 811 858
rect 817 857 818 863
rect 84 801 85 807
rect 91 806 799 807
rect 91 802 111 806
rect 115 802 135 806
rect 139 802 183 806
rect 187 802 231 806
rect 235 802 279 806
rect 283 802 327 806
rect 331 802 375 806
rect 379 802 775 806
rect 779 802 799 806
rect 91 801 799 802
rect 805 801 806 807
rect 96 745 97 751
rect 103 750 811 751
rect 103 746 111 750
rect 115 746 155 750
rect 159 746 203 750
rect 207 746 251 750
rect 255 746 291 750
rect 295 746 299 750
rect 303 746 339 750
rect 343 746 347 750
rect 351 746 387 750
rect 391 746 395 750
rect 399 746 443 750
rect 447 746 507 750
rect 511 746 579 750
rect 583 746 659 750
rect 663 746 739 750
rect 743 746 775 750
rect 779 746 811 750
rect 103 745 811 746
rect 817 745 818 751
rect 84 689 85 695
rect 91 694 799 695
rect 91 690 111 694
rect 115 690 271 694
rect 275 690 319 694
rect 323 690 335 694
rect 339 690 367 694
rect 371 690 383 694
rect 387 690 423 694
rect 427 690 431 694
rect 435 690 479 694
rect 483 690 487 694
rect 491 690 527 694
rect 531 690 559 694
rect 563 690 575 694
rect 579 690 623 694
rect 627 690 639 694
rect 643 690 671 694
rect 675 690 719 694
rect 723 690 775 694
rect 779 690 799 694
rect 91 689 799 690
rect 805 689 806 695
rect 96 633 97 639
rect 103 638 811 639
rect 103 634 111 638
rect 115 634 155 638
rect 159 634 203 638
rect 207 634 275 638
rect 279 634 355 638
rect 359 634 379 638
rect 383 634 403 638
rect 407 634 451 638
rect 455 634 499 638
rect 503 634 547 638
rect 551 634 595 638
rect 599 634 627 638
rect 631 634 643 638
rect 647 634 691 638
rect 695 634 739 638
rect 743 634 775 638
rect 779 634 811 638
rect 103 633 811 634
rect 817 633 818 639
rect 84 577 85 583
rect 91 582 799 583
rect 91 578 111 582
rect 115 578 135 582
rect 139 578 183 582
rect 187 578 255 582
rect 259 578 263 582
rect 267 578 351 582
rect 355 578 359 582
rect 363 578 447 582
rect 451 578 479 582
rect 483 578 543 582
rect 547 578 607 582
rect 611 578 639 582
rect 643 578 719 582
rect 723 578 775 582
rect 779 578 799 582
rect 91 577 799 578
rect 805 577 806 583
rect 96 521 97 527
rect 103 526 811 527
rect 103 522 111 526
rect 115 522 155 526
rect 159 522 203 526
rect 207 522 211 526
rect 215 522 267 526
rect 271 522 283 526
rect 287 522 331 526
rect 335 522 371 526
rect 375 522 403 526
rect 407 522 467 526
rect 471 522 483 526
rect 487 522 563 526
rect 567 522 571 526
rect 575 522 659 526
rect 663 522 667 526
rect 671 522 739 526
rect 743 522 775 526
rect 779 522 811 526
rect 103 521 811 522
rect 817 521 818 527
rect 84 465 85 471
rect 91 470 799 471
rect 91 466 111 470
rect 115 466 191 470
rect 195 466 247 470
rect 251 466 311 470
rect 315 466 351 470
rect 355 466 383 470
rect 387 466 399 470
rect 403 466 447 470
rect 451 466 463 470
rect 467 466 495 470
rect 499 466 543 470
rect 547 466 551 470
rect 555 466 599 470
rect 603 466 647 470
rect 651 466 663 470
rect 667 466 719 470
rect 723 466 775 470
rect 779 466 799 470
rect 91 465 799 466
rect 805 465 806 471
rect 96 405 97 411
rect 103 410 811 411
rect 103 406 111 410
rect 115 406 339 410
rect 343 406 371 410
rect 375 406 387 410
rect 391 406 419 410
rect 423 406 435 410
rect 439 406 467 410
rect 471 406 483 410
rect 487 406 515 410
rect 519 406 539 410
rect 543 406 563 410
rect 567 406 603 410
rect 607 406 619 410
rect 623 406 667 410
rect 671 406 683 410
rect 687 406 739 410
rect 743 406 775 410
rect 779 406 811 410
rect 103 405 811 406
rect 817 405 818 411
rect 84 341 85 347
rect 91 346 799 347
rect 91 342 111 346
rect 115 342 135 346
rect 139 342 199 346
rect 203 342 271 346
rect 275 342 319 346
rect 323 342 343 346
rect 347 342 367 346
rect 371 342 415 346
rect 419 342 423 346
rect 427 342 463 346
rect 467 342 511 346
rect 515 342 519 346
rect 523 342 583 346
rect 587 342 607 346
rect 611 342 647 346
rect 651 342 703 346
rect 707 342 719 346
rect 723 342 775 346
rect 779 342 799 346
rect 91 341 799 342
rect 805 341 806 347
rect 96 277 97 283
rect 103 282 811 283
rect 103 278 111 282
rect 115 278 155 282
rect 159 278 211 282
rect 215 278 219 282
rect 223 278 291 282
rect 295 278 299 282
rect 303 278 363 282
rect 367 278 387 282
rect 391 278 443 282
rect 447 278 475 282
rect 479 278 531 282
rect 535 278 563 282
rect 567 278 627 282
rect 631 278 659 282
rect 663 278 723 282
rect 727 278 739 282
rect 743 278 775 282
rect 779 278 811 282
rect 103 277 811 278
rect 817 277 818 283
rect 84 213 85 219
rect 91 218 799 219
rect 91 214 111 218
rect 115 214 135 218
rect 139 214 191 218
rect 195 214 279 218
rect 283 214 367 218
rect 371 214 455 218
rect 459 214 543 218
rect 547 214 551 218
rect 555 214 639 218
rect 643 214 647 218
rect 651 214 719 218
rect 723 214 775 218
rect 779 214 799 218
rect 91 213 799 214
rect 805 213 806 219
rect 96 149 97 155
rect 103 154 811 155
rect 103 150 111 154
rect 115 150 211 154
rect 215 150 259 154
rect 263 150 299 154
rect 303 150 307 154
rect 311 150 355 154
rect 359 150 387 154
rect 391 150 403 154
rect 407 150 451 154
rect 455 150 475 154
rect 479 150 499 154
rect 503 150 547 154
rect 551 150 571 154
rect 575 150 595 154
rect 599 150 643 154
rect 647 150 667 154
rect 671 150 691 154
rect 695 150 739 154
rect 743 150 775 154
rect 779 150 811 154
rect 103 149 811 150
rect 817 149 818 155
rect 84 93 85 99
rect 91 98 799 99
rect 91 94 111 98
rect 115 94 191 98
rect 195 94 239 98
rect 243 94 287 98
rect 291 94 335 98
rect 339 94 383 98
rect 387 94 431 98
rect 435 94 479 98
rect 483 94 527 98
rect 531 94 575 98
rect 579 94 623 98
rect 627 94 671 98
rect 675 94 719 98
rect 723 94 775 98
rect 779 94 799 98
rect 91 93 799 94
rect 805 93 806 99
<< m5c >>
rect 97 857 103 863
rect 811 857 817 863
rect 85 801 91 807
rect 799 801 805 807
rect 97 745 103 751
rect 811 745 817 751
rect 85 689 91 695
rect 799 689 805 695
rect 97 633 103 639
rect 811 633 817 639
rect 85 577 91 583
rect 799 577 805 583
rect 97 521 103 527
rect 811 521 817 527
rect 85 465 91 471
rect 799 465 805 471
rect 97 405 103 411
rect 811 405 817 411
rect 85 341 91 347
rect 799 341 805 347
rect 97 277 103 283
rect 811 277 817 283
rect 85 213 91 219
rect 799 213 805 219
rect 97 149 103 155
rect 811 149 817 155
rect 85 93 91 99
rect 799 93 805 99
<< m5 >>
rect 84 807 92 864
rect 84 801 85 807
rect 91 801 92 807
rect 84 695 92 801
rect 84 689 85 695
rect 91 689 92 695
rect 84 583 92 689
rect 84 577 85 583
rect 91 577 92 583
rect 84 471 92 577
rect 84 465 85 471
rect 91 465 92 471
rect 84 347 92 465
rect 84 341 85 347
rect 91 341 92 347
rect 84 219 92 341
rect 84 213 85 219
rect 91 213 92 219
rect 84 99 92 213
rect 84 93 85 99
rect 91 93 92 99
rect 84 72 92 93
rect 96 863 104 864
rect 96 857 97 863
rect 103 857 104 863
rect 96 751 104 857
rect 96 745 97 751
rect 103 745 104 751
rect 96 639 104 745
rect 96 633 97 639
rect 103 633 104 639
rect 96 527 104 633
rect 96 521 97 527
rect 103 521 104 527
rect 96 411 104 521
rect 96 405 97 411
rect 103 405 104 411
rect 96 283 104 405
rect 96 277 97 283
rect 103 277 104 283
rect 96 155 104 277
rect 96 149 97 155
rect 103 149 104 155
rect 96 72 104 149
rect 798 807 806 864
rect 798 801 799 807
rect 805 801 806 807
rect 798 695 806 801
rect 798 689 799 695
rect 805 689 806 695
rect 798 583 806 689
rect 798 577 799 583
rect 805 577 806 583
rect 798 471 806 577
rect 798 465 799 471
rect 805 465 806 471
rect 798 347 806 465
rect 798 341 799 347
rect 805 341 806 347
rect 798 219 806 341
rect 798 213 799 219
rect 805 213 806 219
rect 798 99 806 213
rect 798 93 799 99
rect 805 93 806 99
rect 798 72 806 93
rect 810 863 818 864
rect 810 857 811 863
rect 817 857 818 863
rect 810 751 818 857
rect 810 745 811 751
rect 817 745 818 751
rect 810 639 818 745
rect 810 633 811 639
rect 817 633 818 639
rect 810 527 818 633
rect 810 521 811 527
rect 817 521 818 527
rect 810 411 818 521
rect 810 405 811 411
rect 817 405 818 411
rect 810 283 818 405
rect 810 277 811 283
rect 817 277 818 283
rect 810 155 818 277
rect 810 149 811 155
rect 817 149 818 155
rect 810 72 818 149
use welltap_svt  __well_tap__0
timestamp 1730593976
transform 1 0 104 0 1 112
box 8 4 12 24
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__0
timestamp 1730593976
transform 1 0 104 0 1 112
box 8 4 12 24
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use _0_0std_0_0cells_0_0OR2X1  or_561_6
timestamp 1730593976
transform 1 0 184 0 1 96
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_561_6
timestamp 1730593976
transform 1 0 184 0 1 96
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_562_6
timestamp 1730593976
transform 1 0 232 0 1 96
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_562_6
timestamp 1730593976
transform 1 0 232 0 1 96
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_563_6
timestamp 1730593976
transform 1 0 280 0 1 96
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_563_6
timestamp 1730593976
transform 1 0 280 0 1 96
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_564_6
timestamp 1730593976
transform 1 0 328 0 1 96
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_564_6
timestamp 1730593976
transform 1 0 328 0 1 96
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_565_6
timestamp 1730593976
transform 1 0 376 0 1 96
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_565_6
timestamp 1730593976
transform 1 0 376 0 1 96
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_566_6
timestamp 1730593976
transform 1 0 424 0 1 96
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_566_6
timestamp 1730593976
transform 1 0 424 0 1 96
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_567_6
timestamp 1730593976
transform 1 0 472 0 1 96
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_567_6
timestamp 1730593976
transform 1 0 472 0 1 96
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_568_6
timestamp 1730593976
transform 1 0 520 0 1 96
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_568_6
timestamp 1730593976
transform 1 0 520 0 1 96
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_569_6
timestamp 1730593976
transform 1 0 568 0 1 96
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_569_6
timestamp 1730593976
transform 1 0 568 0 1 96
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_599_6
timestamp 1730593976
transform 1 0 616 0 1 96
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_599_6
timestamp 1730593976
transform 1 0 616 0 1 96
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_598_6
timestamp 1730593976
transform 1 0 664 0 1 96
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_598_6
timestamp 1730593976
transform 1 0 664 0 1 96
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_597_6
timestamp 1730593976
transform 1 0 712 0 1 96
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_597_6
timestamp 1730593976
transform 1 0 712 0 1 96
box 7 3 44 54
use welltap_svt  __well_tap__1
timestamp 1730593976
transform 1 0 768 0 1 112
box 8 4 12 24
use welltap_svt  __well_tap__1
timestamp 1730593976
transform 1 0 768 0 1 112
box 8 4 12 24
use _0_0std_0_0cells_0_0OR2X1  or_560_6
timestamp 1730593976
transform 1 0 184 0 -1 216
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_560_6
timestamp 1730593976
transform 1 0 184 0 -1 216
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_559_6
timestamp 1730593976
transform 1 0 272 0 -1 216
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_559_6
timestamp 1730593976
transform 1 0 272 0 -1 216
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_558_6
timestamp 1730593976
transform 1 0 360 0 -1 216
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_558_6
timestamp 1730593976
transform 1 0 360 0 -1 216
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_571_6
timestamp 1730593976
transform 1 0 448 0 -1 216
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_571_6
timestamp 1730593976
transform 1 0 448 0 -1 216
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_570_6
timestamp 1730593976
transform 1 0 544 0 -1 216
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_570_6
timestamp 1730593976
transform 1 0 544 0 -1 216
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_595_6
timestamp 1730593976
transform 1 0 640 0 -1 216
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_595_6
timestamp 1730593976
transform 1 0 640 0 -1 216
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_596_6
timestamp 1730593976
transform 1 0 712 0 -1 216
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_596_6
timestamp 1730593976
transform 1 0 712 0 -1 216
box 7 3 44 54
use welltap_svt  __well_tap__2
timestamp 1730593976
transform 1 0 104 0 -1 200
box 8 4 12 24
use welltap_svt  __well_tap__2
timestamp 1730593976
transform 1 0 104 0 -1 200
box 8 4 12 24
use _0_0std_0_0cells_0_0OR2X1  or_554_6
timestamp 1730593976
transform 1 0 128 0 1 224
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_554_6
timestamp 1730593976
transform 1 0 128 0 1 224
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_555_6
timestamp 1730593976
transform 1 0 184 0 1 224
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_555_6
timestamp 1730593976
transform 1 0 184 0 1 224
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_556_6
timestamp 1730593976
transform 1 0 272 0 1 224
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_556_6
timestamp 1730593976
transform 1 0 272 0 1 224
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_557_6
timestamp 1730593976
transform 1 0 360 0 1 224
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_557_6
timestamp 1730593976
transform 1 0 360 0 1 224
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_572_6
timestamp 1730593976
transform 1 0 448 0 1 224
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_572_6
timestamp 1730593976
transform 1 0 448 0 1 224
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_573_6
timestamp 1730593976
transform 1 0 536 0 1 224
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_573_6
timestamp 1730593976
transform 1 0 536 0 1 224
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_594_6
timestamp 1730593976
transform 1 0 632 0 1 224
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_594_6
timestamp 1730593976
transform 1 0 632 0 1 224
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_593_6
timestamp 1730593976
transform 1 0 712 0 1 224
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_593_6
timestamp 1730593976
transform 1 0 712 0 1 224
box 7 3 44 54
use welltap_svt  __well_tap__3
timestamp 1730593976
transform 1 0 768 0 -1 200
box 8 4 12 24
use welltap_svt  __well_tap__3
timestamp 1730593976
transform 1 0 768 0 -1 200
box 8 4 12 24
use welltap_svt  __well_tap__4
timestamp 1730593976
transform 1 0 104 0 1 240
box 8 4 12 24
use welltap_svt  __well_tap__4
timestamp 1730593976
transform 1 0 104 0 1 240
box 8 4 12 24
use welltap_svt  __well_tap__5
timestamp 1730593976
transform 1 0 768 0 1 240
box 8 4 12 24
use welltap_svt  __well_tap__5
timestamp 1730593976
transform 1 0 768 0 1 240
box 8 4 12 24
use welltap_svt  __well_tap__6
timestamp 1730593976
transform 1 0 104 0 -1 328
box 8 4 12 24
use welltap_svt  __well_tap__6
timestamp 1730593976
transform 1 0 104 0 -1 328
box 8 4 12 24
use _0_0std_0_0cells_0_0OR2X1  or_553_6
timestamp 1730593976
transform 1 0 128 0 -1 344
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_553_6
timestamp 1730593976
transform 1 0 128 0 -1 344
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_552_6
timestamp 1730593976
transform 1 0 192 0 -1 344
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_552_6
timestamp 1730593976
transform 1 0 192 0 -1 344
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_551_6
timestamp 1730593976
transform 1 0 264 0 -1 344
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_551_6
timestamp 1730593976
transform 1 0 264 0 -1 344
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_550_6
timestamp 1730593976
transform 1 0 336 0 -1 344
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_550_6
timestamp 1730593976
transform 1 0 336 0 -1 344
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_549_6
timestamp 1730593976
transform 1 0 416 0 -1 344
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_549_6
timestamp 1730593976
transform 1 0 416 0 -1 344
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_574_6
timestamp 1730593976
transform 1 0 504 0 -1 344
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_574_6
timestamp 1730593976
transform 1 0 504 0 -1 344
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_575_6
timestamp 1730593976
transform 1 0 600 0 -1 344
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_575_6
timestamp 1730593976
transform 1 0 600 0 -1 344
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_592_6
timestamp 1730593976
transform 1 0 696 0 -1 344
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_592_6
timestamp 1730593976
transform 1 0 696 0 -1 344
box 7 3 44 54
use welltap_svt  __well_tap__7
timestamp 1730593976
transform 1 0 768 0 -1 328
box 8 4 12 24
use welltap_svt  __well_tap__7
timestamp 1730593976
transform 1 0 768 0 -1 328
box 8 4 12 24
use welltap_svt  __well_tap__8
timestamp 1730593976
transform 1 0 104 0 1 368
box 8 4 12 24
use welltap_svt  __well_tap__8
timestamp 1730593976
transform 1 0 104 0 1 368
box 8 4 12 24
use _0_0std_0_0cells_0_0OR2X1  or_546_6
timestamp 1730593976
transform 1 0 312 0 1 352
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_546_6
timestamp 1730593976
transform 1 0 312 0 1 352
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_547_6
timestamp 1730593976
transform 1 0 360 0 1 352
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_547_6
timestamp 1730593976
transform 1 0 360 0 1 352
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_548_6
timestamp 1730593976
transform 1 0 408 0 1 352
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_548_6
timestamp 1730593976
transform 1 0 408 0 1 352
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_545_6
timestamp 1730593976
transform 1 0 456 0 1 352
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_545_6
timestamp 1730593976
transform 1 0 456 0 1 352
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_544_6
timestamp 1730593976
transform 1 0 512 0 1 352
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_544_6
timestamp 1730593976
transform 1 0 512 0 1 352
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_543_6
timestamp 1730593976
transform 1 0 576 0 1 352
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_543_6
timestamp 1730593976
transform 1 0 576 0 1 352
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_576_6
timestamp 1730593976
transform 1 0 640 0 1 352
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_576_6
timestamp 1730593976
transform 1 0 640 0 1 352
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_591_6
timestamp 1730593976
transform 1 0 712 0 1 352
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_591_6
timestamp 1730593976
transform 1 0 712 0 1 352
box 7 3 44 54
use welltap_svt  __well_tap__9
timestamp 1730593976
transform 1 0 768 0 1 368
box 8 4 12 24
use welltap_svt  __well_tap__9
timestamp 1730593976
transform 1 0 768 0 1 368
box 8 4 12 24
use welltap_svt  __well_tap__10
timestamp 1730593976
transform 1 0 104 0 -1 452
box 8 4 12 24
use welltap_svt  __well_tap__10
timestamp 1730593976
transform 1 0 104 0 -1 452
box 8 4 12 24
use _0_0std_0_0cells_0_0OR2X1  or_537_6
timestamp 1730593976
transform 1 0 344 0 -1 468
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_537_6
timestamp 1730593976
transform 1 0 344 0 -1 468
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_538_6
timestamp 1730593976
transform 1 0 392 0 -1 468
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_538_6
timestamp 1730593976
transform 1 0 392 0 -1 468
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_539_6
timestamp 1730593976
transform 1 0 440 0 -1 468
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_539_6
timestamp 1730593976
transform 1 0 440 0 -1 468
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_540_6
timestamp 1730593976
transform 1 0 488 0 -1 468
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_540_6
timestamp 1730593976
transform 1 0 488 0 -1 468
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_541_6
timestamp 1730593976
transform 1 0 536 0 -1 468
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_541_6
timestamp 1730593976
transform 1 0 536 0 -1 468
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_542_6
timestamp 1730593976
transform 1 0 592 0 -1 468
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_542_6
timestamp 1730593976
transform 1 0 592 0 -1 468
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_577_6
timestamp 1730593976
transform 1 0 656 0 -1 468
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_577_6
timestamp 1730593976
transform 1 0 656 0 -1 468
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_590_6
timestamp 1730593976
transform 1 0 712 0 -1 468
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_590_6
timestamp 1730593976
transform 1 0 712 0 -1 468
box 7 3 44 54
use welltap_svt  __well_tap__11
timestamp 1730593976
transform 1 0 768 0 -1 452
box 8 4 12 24
use welltap_svt  __well_tap__11
timestamp 1730593976
transform 1 0 768 0 -1 452
box 8 4 12 24
use _0_0std_0_0cells_0_0OR2X1  or_531_6
timestamp 1730593976
transform 1 0 184 0 1 468
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_531_6
timestamp 1730593976
transform 1 0 184 0 1 468
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_532_6
timestamp 1730593976
transform 1 0 240 0 1 468
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_532_6
timestamp 1730593976
transform 1 0 240 0 1 468
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_533_6
timestamp 1730593976
transform 1 0 304 0 1 468
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_533_6
timestamp 1730593976
transform 1 0 304 0 1 468
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_534_6
timestamp 1730593976
transform 1 0 376 0 1 468
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_534_6
timestamp 1730593976
transform 1 0 376 0 1 468
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_535_6
timestamp 1730593976
transform 1 0 456 0 1 468
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_535_6
timestamp 1730593976
transform 1 0 456 0 1 468
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_536_6
timestamp 1730593976
transform 1 0 544 0 1 468
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_536_6
timestamp 1730593976
transform 1 0 544 0 1 468
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_578_6
timestamp 1730593976
transform 1 0 640 0 1 468
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_578_6
timestamp 1730593976
transform 1 0 640 0 1 468
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_589_6
timestamp 1730593976
transform 1 0 712 0 1 468
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_589_6
timestamp 1730593976
transform 1 0 712 0 1 468
box 7 3 44 54
use welltap_svt  __well_tap__12
timestamp 1730593976
transform 1 0 104 0 1 484
box 8 4 12 24
use welltap_svt  __well_tap__12
timestamp 1730593976
transform 1 0 104 0 1 484
box 8 4 12 24
use _0_0std_0_0cells_0_0OR2X1  or_526_6
timestamp 1730593976
transform 1 0 128 0 -1 580
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_526_6
timestamp 1730593976
transform 1 0 128 0 -1 580
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_527_6
timestamp 1730593976
transform 1 0 176 0 -1 580
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_527_6
timestamp 1730593976
transform 1 0 176 0 -1 580
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_528_6
timestamp 1730593976
transform 1 0 256 0 -1 580
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_528_6
timestamp 1730593976
transform 1 0 256 0 -1 580
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_529_6
timestamp 1730593976
transform 1 0 344 0 -1 580
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_529_6
timestamp 1730593976
transform 1 0 344 0 -1 580
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_530_6
timestamp 1730593976
transform 1 0 440 0 -1 580
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_530_6
timestamp 1730593976
transform 1 0 440 0 -1 580
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_579_6
timestamp 1730593976
transform 1 0 536 0 -1 580
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_579_6
timestamp 1730593976
transform 1 0 536 0 -1 580
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_588_6
timestamp 1730593976
transform 1 0 632 0 -1 580
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_588_6
timestamp 1730593976
transform 1 0 632 0 -1 580
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_587_6
timestamp 1730593976
transform 1 0 712 0 -1 580
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_587_6
timestamp 1730593976
transform 1 0 712 0 -1 580
box 7 3 44 54
use welltap_svt  __well_tap__13
timestamp 1730593976
transform 1 0 768 0 1 484
box 8 4 12 24
use welltap_svt  __well_tap__13
timestamp 1730593976
transform 1 0 768 0 1 484
box 8 4 12 24
use welltap_svt  __well_tap__14
timestamp 1730593976
transform 1 0 104 0 -1 564
box 8 4 12 24
use welltap_svt  __well_tap__14
timestamp 1730593976
transform 1 0 104 0 -1 564
box 8 4 12 24
use _0_0std_0_0cells_0_0OR2X1  or_525_6
timestamp 1730593976
transform 1 0 128 0 1 580
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_525_6
timestamp 1730593976
transform 1 0 128 0 1 580
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_524_6
timestamp 1730593976
transform 1 0 176 0 1 580
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_524_6
timestamp 1730593976
transform 1 0 176 0 1 580
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_523_6
timestamp 1730593976
transform 1 0 248 0 1 580
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_523_6
timestamp 1730593976
transform 1 0 248 0 1 580
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_522_6
timestamp 1730593976
transform 1 0 352 0 1 580
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_522_6
timestamp 1730593976
transform 1 0 352 0 1 580
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_520_6
timestamp 1730593976
transform 1 0 472 0 1 580
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_520_6
timestamp 1730593976
transform 1 0 472 0 1 580
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_521_6
timestamp 1730593976
transform 1 0 600 0 1 580
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_521_6
timestamp 1730593976
transform 1 0 600 0 1 580
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_586_6
timestamp 1730593976
transform 1 0 712 0 1 580
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_586_6
timestamp 1730593976
transform 1 0 712 0 1 580
box 7 3 44 54
use welltap_svt  __well_tap__15
timestamp 1730593976
transform 1 0 768 0 -1 564
box 8 4 12 24
use welltap_svt  __well_tap__15
timestamp 1730593976
transform 1 0 768 0 -1 564
box 8 4 12 24
use welltap_svt  __well_tap__16
timestamp 1730593976
transform 1 0 104 0 1 596
box 8 4 12 24
use welltap_svt  __well_tap__16
timestamp 1730593976
transform 1 0 104 0 1 596
box 8 4 12 24
use _0_0std_0_0cells_0_0OR2X1  or_517_6
timestamp 1730593976
transform 1 0 328 0 -1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_517_6
timestamp 1730593976
transform 1 0 328 0 -1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_518_6
timestamp 1730593976
transform 1 0 376 0 -1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_518_6
timestamp 1730593976
transform 1 0 376 0 -1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_519_6
timestamp 1730593976
transform 1 0 424 0 -1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_519_6
timestamp 1730593976
transform 1 0 424 0 -1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_516_6
timestamp 1730593976
transform 1 0 472 0 -1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_516_6
timestamp 1730593976
transform 1 0 472 0 -1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_515_6
timestamp 1730593976
transform 1 0 520 0 -1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_515_6
timestamp 1730593976
transform 1 0 520 0 -1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_580_6
timestamp 1730593976
transform 1 0 568 0 -1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_580_6
timestamp 1730593976
transform 1 0 568 0 -1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_581_6
timestamp 1730593976
transform 1 0 616 0 -1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_581_6
timestamp 1730593976
transform 1 0 616 0 -1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_584_6
timestamp 1730593976
transform 1 0 664 0 -1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_584_6
timestamp 1730593976
transform 1 0 664 0 -1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_585_6
timestamp 1730593976
transform 1 0 712 0 -1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_585_6
timestamp 1730593976
transform 1 0 712 0 -1 692
box 7 3 44 54
use welltap_svt  __well_tap__17
timestamp 1730593976
transform 1 0 768 0 1 596
box 8 4 12 24
use welltap_svt  __well_tap__17
timestamp 1730593976
transform 1 0 768 0 1 596
box 8 4 12 24
use welltap_svt  __well_tap__18
timestamp 1730593976
transform 1 0 104 0 -1 676
box 8 4 12 24
use welltap_svt  __well_tap__18
timestamp 1730593976
transform 1 0 104 0 -1 676
box 8 4 12 24
use _0_0std_0_0cells_0_0OR2X1  or_59_6
timestamp 1730593976
transform 1 0 264 0 1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_59_6
timestamp 1730593976
transform 1 0 264 0 1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_510_6
timestamp 1730593976
transform 1 0 312 0 1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_510_6
timestamp 1730593976
transform 1 0 312 0 1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_511_6
timestamp 1730593976
transform 1 0 360 0 1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_511_6
timestamp 1730593976
transform 1 0 360 0 1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_512_6
timestamp 1730593976
transform 1 0 416 0 1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_512_6
timestamp 1730593976
transform 1 0 416 0 1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_513_6
timestamp 1730593976
transform 1 0 480 0 1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_513_6
timestamp 1730593976
transform 1 0 480 0 1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_514_6
timestamp 1730593976
transform 1 0 552 0 1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_514_6
timestamp 1730593976
transform 1 0 552 0 1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_582_6
timestamp 1730593976
transform 1 0 632 0 1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_582_6
timestamp 1730593976
transform 1 0 632 0 1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_583_6
timestamp 1730593976
transform 1 0 712 0 1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_583_6
timestamp 1730593976
transform 1 0 712 0 1 692
box 7 3 44 54
use welltap_svt  __well_tap__19
timestamp 1730593976
transform 1 0 768 0 -1 676
box 8 4 12 24
use welltap_svt  __well_tap__19
timestamp 1730593976
transform 1 0 768 0 -1 676
box 8 4 12 24
use welltap_svt  __well_tap__20
timestamp 1730593976
transform 1 0 104 0 1 708
box 8 4 12 24
use welltap_svt  __well_tap__20
timestamp 1730593976
transform 1 0 104 0 1 708
box 8 4 12 24
use welltap_svt  __well_tap__21
timestamp 1730593976
transform 1 0 768 0 1 708
box 8 4 12 24
use welltap_svt  __well_tap__21
timestamp 1730593976
transform 1 0 768 0 1 708
box 8 4 12 24
use welltap_svt  __well_tap__22
timestamp 1730593976
transform 1 0 104 0 -1 788
box 8 4 12 24
use welltap_svt  __well_tap__22
timestamp 1730593976
transform 1 0 104 0 -1 788
box 8 4 12 24
use _0_0std_0_0cells_0_0OR2X1  or_53_6
timestamp 1730593976
transform 1 0 128 0 -1 804
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_53_6
timestamp 1730593976
transform 1 0 128 0 -1 804
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_54_6
timestamp 1730593976
transform 1 0 176 0 -1 804
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_54_6
timestamp 1730593976
transform 1 0 176 0 -1 804
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_55_6
timestamp 1730593976
transform 1 0 224 0 -1 804
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_55_6
timestamp 1730593976
transform 1 0 224 0 -1 804
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_56_6
timestamp 1730593976
transform 1 0 272 0 -1 804
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_56_6
timestamp 1730593976
transform 1 0 272 0 -1 804
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_57_6
timestamp 1730593976
transform 1 0 320 0 -1 804
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_57_6
timestamp 1730593976
transform 1 0 320 0 -1 804
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_58_6
timestamp 1730593976
transform 1 0 368 0 -1 804
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_58_6
timestamp 1730593976
transform 1 0 368 0 -1 804
box 7 3 44 54
use welltap_svt  __well_tap__23
timestamp 1730593976
transform 1 0 768 0 -1 788
box 8 4 12 24
use welltap_svt  __well_tap__23
timestamp 1730593976
transform 1 0 768 0 -1 788
box 8 4 12 24
use welltap_svt  __well_tap__24
timestamp 1730593976
transform 1 0 104 0 1 820
box 8 4 12 24
use welltap_svt  __well_tap__24
timestamp 1730593976
transform 1 0 104 0 1 820
box 8 4 12 24
use _0_0std_0_0cells_0_0OR2X1  or_52_6
timestamp 1730593976
transform 1 0 128 0 1 804
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_52_6
timestamp 1730593976
transform 1 0 128 0 1 804
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_51_6
timestamp 1730593976
transform 1 0 176 0 1 804
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_51_6
timestamp 1730593976
transform 1 0 176 0 1 804
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_50_6
timestamp 1730593976
transform 1 0 224 0 1 804
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_50_6
timestamp 1730593976
transform 1 0 224 0 1 804
box 7 3 44 54
use welltap_svt  __well_tap__25
timestamp 1730593976
transform 1 0 768 0 1 820
box 8 4 12 24
use welltap_svt  __well_tap__25
timestamp 1730593976
transform 1 0 768 0 1 820
box 8 4 12 24
<< end >>
