magic
tech sky130l
timestamp 1731220645
<< m1 >>
rect 248 2315 252 2347
rect 992 2315 996 2347
rect 1392 2315 1396 2347
rect 1440 2315 1444 2347
rect 1504 2315 1508 2347
rect 1808 2315 1812 2347
rect 1888 2315 1892 2347
rect 1960 2315 1964 2347
rect 2104 2315 2108 2347
rect 2192 2315 2196 2399
rect 2336 2315 2340 2347
rect 1856 2263 1860 2295
rect 1928 2263 1932 2295
rect 600 2223 604 2255
rect 864 2223 868 2255
rect 944 2223 948 2255
rect 592 2183 596 2219
rect 1672 2167 1676 2199
rect 2216 2167 2220 2199
rect 1928 2119 1932 2151
rect 584 2079 588 2111
rect 640 2079 644 2111
rect 728 2031 732 2063
rect 1792 2027 1796 2059
rect 544 1935 548 1967
rect 664 1935 668 2027
rect 2344 2015 2348 2059
rect 248 1883 252 1915
rect 456 1891 460 1915
rect 672 1883 676 1915
rect 1336 1883 1340 1915
rect 1392 1883 1396 1915
rect 1608 1883 1612 1915
rect 2064 1883 2068 1967
rect 1528 1835 1532 1867
rect 1928 1843 1932 1867
rect 2008 1835 2012 1867
rect 248 1787 252 1819
rect 664 1787 668 1819
rect 760 1787 764 1819
rect 1064 1739 1068 1771
rect 1704 1651 1708 1727
rect 1840 1695 1844 1727
rect 1640 1559 1644 1591
rect 1816 1559 1820 1591
rect 1880 1515 1884 1591
rect 1872 1467 1876 1499
rect 304 1411 308 1443
rect 1568 1323 1572 1355
rect 1640 1323 1644 1355
rect 1800 1323 1804 1355
rect 1880 1323 1884 1355
rect 536 1275 540 1303
rect 1720 1275 1724 1307
rect 1944 1275 1948 1307
rect 264 1171 268 1211
rect 344 1179 348 1211
rect 432 1179 436 1211
rect 520 1179 524 1211
rect 776 1179 780 1211
rect 848 1179 852 1211
rect 912 1179 916 1211
rect 976 1179 980 1211
rect 1040 1179 1044 1211
rect 1336 1179 1340 1211
rect 1408 1179 1412 1211
rect 272 1131 276 1163
rect 1384 1131 1388 1163
rect 2216 1131 2220 1163
rect 568 1039 572 1071
rect 1856 1043 1860 1075
rect 1904 1043 1908 1075
rect 1952 1043 1956 1075
rect 2048 1043 2052 1075
rect 2096 1043 2100 1075
rect 1984 999 1988 1027
rect 392 903 396 935
rect 1104 903 1108 935
rect 1336 899 1340 931
rect 1384 899 1388 931
rect 1464 899 1468 931
rect 1656 899 1660 931
rect 1800 899 1804 931
rect 1888 899 1892 931
rect 1992 899 1996 991
rect 336 847 340 879
rect 1592 851 1596 883
rect 1688 855 1692 883
rect 1968 855 1972 883
rect 176 707 180 739
rect 320 707 324 739
rect 672 615 676 647
rect 744 615 748 647
rect 1656 611 1660 643
rect 2080 611 2084 643
rect 2144 611 2148 643
rect 2208 611 2212 643
rect 1824 571 1828 591
rect 1832 563 1836 591
rect 1952 559 1956 591
rect 176 463 180 495
rect 368 463 372 495
rect 448 463 452 495
rect 528 463 532 495
rect 768 463 772 495
rect 1408 471 1412 503
rect 1512 471 1516 503
rect 168 415 172 459
rect 648 415 652 447
rect 760 415 764 447
rect 1376 419 1380 451
rect 2336 427 2340 451
rect 376 327 380 359
rect 424 327 428 359
rect 2144 327 2148 359
rect 2208 327 2212 359
rect 2272 327 2276 359
rect 536 275 540 307
rect 1896 275 1900 307
rect 1528 183 1532 215
rect 1584 183 1588 215
rect 2104 183 2108 215
rect 2200 183 2204 215
rect 408 111 412 143
rect 664 115 668 143
rect 960 111 964 143
rect 1552 119 1556 151
rect 1616 123 1620 151
rect 1752 123 1756 151
rect 1800 119 1804 151
<< m2c >>
rect 172 2491 176 2495
rect 212 2491 216 2495
rect 252 2491 256 2495
rect 308 2491 312 2495
rect 388 2491 392 2495
rect 476 2491 480 2495
rect 564 2491 568 2495
rect 652 2491 656 2495
rect 740 2491 744 2495
rect 828 2491 832 2495
rect 924 2491 928 2495
rect 1560 2483 1564 2487
rect 1600 2483 1604 2487
rect 1640 2483 1644 2487
rect 1680 2483 1684 2487
rect 1720 2483 1724 2487
rect 1760 2483 1764 2487
rect 1800 2483 1804 2487
rect 1840 2483 1844 2487
rect 1880 2483 1884 2487
rect 1920 2483 1924 2487
rect 1960 2483 1964 2487
rect 2000 2483 2004 2487
rect 160 2455 164 2459
rect 200 2455 204 2459
rect 240 2455 244 2459
rect 280 2455 284 2459
rect 336 2455 340 2459
rect 416 2455 420 2459
rect 504 2455 508 2459
rect 592 2455 596 2459
rect 680 2455 684 2459
rect 768 2455 772 2459
rect 856 2455 860 2459
rect 952 2455 956 2459
rect 1532 2447 1536 2451
rect 1572 2447 1576 2451
rect 1612 2449 1616 2453
rect 1652 2447 1656 2451
rect 1692 2449 1696 2453
rect 1732 2447 1736 2451
rect 1772 2449 1776 2453
rect 1812 2447 1816 2451
rect 1852 2449 1856 2453
rect 1892 2447 1896 2451
rect 1932 2449 1936 2453
rect 1972 2447 1976 2451
rect 1356 2435 1360 2439
rect 1396 2435 1400 2439
rect 1452 2435 1456 2439
rect 1516 2435 1520 2439
rect 1596 2435 1600 2439
rect 1676 2435 1680 2439
rect 1756 2435 1760 2439
rect 1836 2435 1840 2439
rect 1916 2435 1920 2439
rect 1996 2435 2000 2439
rect 2076 2435 2080 2439
rect 2156 2435 2160 2439
rect 2244 2435 2248 2439
rect 2332 2435 2336 2439
rect 160 2403 164 2407
rect 208 2403 212 2407
rect 272 2403 276 2407
rect 344 2403 348 2407
rect 416 2403 420 2407
rect 496 2403 500 2407
rect 568 2403 572 2407
rect 640 2403 644 2407
rect 704 2403 708 2407
rect 760 2403 764 2407
rect 816 2403 820 2407
rect 864 2403 868 2407
rect 912 2403 916 2407
rect 960 2403 964 2407
rect 1016 2403 1020 2407
rect 1072 2403 1076 2407
rect 1384 2399 1388 2403
rect 1424 2399 1428 2403
rect 1480 2399 1484 2403
rect 1544 2399 1548 2403
rect 1624 2399 1628 2403
rect 1704 2399 1708 2403
rect 1784 2399 1788 2403
rect 1864 2399 1868 2403
rect 1944 2399 1948 2403
rect 2024 2399 2028 2403
rect 2104 2399 2108 2403
rect 2184 2399 2188 2403
rect 2192 2399 2196 2403
rect 2272 2399 2276 2403
rect 2360 2399 2364 2403
rect 132 2367 136 2371
rect 180 2367 184 2371
rect 244 2367 248 2371
rect 316 2367 320 2371
rect 388 2367 392 2371
rect 468 2367 472 2371
rect 540 2367 544 2371
rect 612 2367 616 2371
rect 676 2367 680 2371
rect 732 2367 736 2371
rect 788 2367 792 2371
rect 836 2367 840 2371
rect 884 2367 888 2371
rect 932 2367 936 2371
rect 988 2367 992 2371
rect 1044 2367 1048 2371
rect 132 2347 136 2351
rect 172 2347 176 2351
rect 212 2347 216 2351
rect 248 2347 252 2351
rect 268 2347 272 2351
rect 348 2347 352 2351
rect 428 2347 432 2351
rect 516 2347 520 2351
rect 596 2347 600 2351
rect 676 2347 680 2351
rect 748 2347 752 2351
rect 820 2349 824 2353
rect 884 2347 888 2351
rect 956 2347 960 2351
rect 992 2347 996 2351
rect 1028 2347 1032 2351
rect 1384 2347 1388 2351
rect 1392 2347 1396 2351
rect 1432 2347 1436 2351
rect 1440 2347 1444 2351
rect 1496 2347 1500 2351
rect 1504 2347 1508 2351
rect 1568 2347 1572 2351
rect 1640 2347 1644 2351
rect 1720 2347 1724 2351
rect 1800 2347 1804 2351
rect 1808 2347 1812 2351
rect 1880 2347 1884 2351
rect 1888 2347 1892 2351
rect 1952 2347 1956 2351
rect 1960 2347 1964 2351
rect 2024 2347 2028 2351
rect 2096 2347 2100 2351
rect 2104 2347 2108 2351
rect 2168 2347 2172 2351
rect 2248 2349 2252 2353
rect 2328 2347 2332 2351
rect 2336 2347 2340 2351
rect 2384 2347 2388 2351
rect 160 2311 164 2315
rect 200 2311 204 2315
rect 240 2311 244 2315
rect 248 2311 252 2315
rect 296 2311 300 2315
rect 376 2311 380 2315
rect 456 2311 460 2315
rect 544 2311 548 2315
rect 624 2311 628 2315
rect 704 2311 708 2315
rect 776 2311 780 2315
rect 848 2311 852 2315
rect 912 2311 916 2315
rect 984 2311 988 2315
rect 992 2311 996 2315
rect 1056 2311 1060 2315
rect 1356 2311 1360 2315
rect 1392 2311 1396 2315
rect 1404 2311 1408 2315
rect 1440 2311 1444 2315
rect 1468 2311 1472 2315
rect 1504 2311 1508 2315
rect 1540 2311 1544 2315
rect 1612 2311 1616 2315
rect 1692 2311 1696 2315
rect 1772 2311 1776 2315
rect 1808 2311 1812 2315
rect 1852 2311 1856 2315
rect 1888 2311 1892 2315
rect 1924 2311 1928 2315
rect 1960 2311 1964 2315
rect 1996 2311 2000 2315
rect 2068 2311 2072 2315
rect 2104 2311 2108 2315
rect 2140 2311 2144 2315
rect 2192 2311 2196 2315
rect 2220 2311 2224 2315
rect 2300 2311 2304 2315
rect 2336 2311 2340 2315
rect 2356 2311 2360 2315
rect 1500 2295 1504 2299
rect 1540 2295 1544 2299
rect 1580 2295 1584 2299
rect 1620 2295 1624 2299
rect 1660 2295 1664 2299
rect 1700 2295 1704 2299
rect 1756 2295 1760 2299
rect 1820 2295 1824 2299
rect 1856 2295 1860 2299
rect 1892 2295 1896 2299
rect 1928 2295 1932 2299
rect 1964 2295 1968 2299
rect 2044 2295 2048 2299
rect 2124 2295 2128 2299
rect 2204 2295 2208 2299
rect 2292 2295 2296 2299
rect 2356 2295 2360 2299
rect 1528 2259 1532 2263
rect 1568 2259 1572 2263
rect 1608 2259 1612 2263
rect 1648 2259 1652 2263
rect 1688 2259 1692 2263
rect 1728 2259 1732 2263
rect 1784 2259 1788 2263
rect 1848 2259 1852 2263
rect 1856 2259 1860 2263
rect 1920 2259 1924 2263
rect 1928 2259 1932 2263
rect 1992 2259 1996 2263
rect 2072 2259 2076 2263
rect 2152 2259 2156 2263
rect 2232 2259 2236 2263
rect 2320 2259 2324 2263
rect 2384 2259 2388 2263
rect 160 2255 164 2259
rect 200 2255 204 2259
rect 256 2255 260 2259
rect 328 2255 332 2259
rect 400 2255 404 2259
rect 480 2255 484 2259
rect 560 2255 564 2259
rect 600 2255 604 2259
rect 640 2255 644 2259
rect 712 2255 716 2259
rect 784 2255 788 2259
rect 856 2255 860 2259
rect 864 2255 868 2259
rect 936 2255 940 2259
rect 944 2255 948 2259
rect 1016 2255 1020 2259
rect 132 2219 136 2223
rect 172 2219 176 2223
rect 228 2219 232 2223
rect 300 2219 304 2223
rect 372 2219 376 2223
rect 452 2219 456 2223
rect 532 2219 536 2223
rect 592 2219 596 2223
rect 600 2219 604 2223
rect 612 2219 616 2223
rect 684 2219 688 2223
rect 756 2219 760 2223
rect 828 2219 832 2223
rect 864 2219 868 2223
rect 908 2219 912 2223
rect 944 2219 948 2223
rect 988 2219 992 2223
rect 244 2207 248 2211
rect 284 2207 288 2211
rect 324 2207 328 2211
rect 372 2207 376 2211
rect 428 2207 432 2211
rect 492 2207 496 2211
rect 548 2207 552 2211
rect 604 2207 608 2211
rect 660 2207 664 2211
rect 716 2207 720 2211
rect 780 2207 784 2211
rect 844 2207 848 2211
rect 908 2207 912 2211
rect 1328 2199 1332 2203
rect 1368 2199 1372 2203
rect 1408 2199 1412 2203
rect 1456 2199 1460 2203
rect 1520 2199 1524 2203
rect 1592 2199 1596 2203
rect 1664 2199 1668 2203
rect 1672 2199 1676 2203
rect 1736 2199 1740 2203
rect 1808 2199 1812 2203
rect 1880 2199 1884 2203
rect 1960 2199 1964 2203
rect 2040 2199 2044 2203
rect 2120 2199 2124 2203
rect 2208 2199 2212 2203
rect 2216 2199 2220 2203
rect 2304 2199 2308 2203
rect 2384 2199 2388 2203
rect 592 2179 596 2183
rect 272 2171 276 2175
rect 312 2171 316 2175
rect 352 2171 356 2175
rect 400 2171 404 2175
rect 456 2171 460 2175
rect 520 2171 524 2175
rect 576 2171 580 2175
rect 632 2171 636 2175
rect 688 2171 692 2175
rect 744 2171 748 2175
rect 808 2171 812 2175
rect 872 2171 876 2175
rect 936 2171 940 2175
rect 1300 2163 1304 2167
rect 1340 2163 1344 2167
rect 1380 2163 1384 2167
rect 1428 2163 1432 2167
rect 1492 2163 1496 2167
rect 1564 2163 1568 2167
rect 1636 2163 1640 2167
rect 1672 2163 1676 2167
rect 1708 2163 1712 2167
rect 1780 2163 1784 2167
rect 1852 2163 1856 2167
rect 1932 2163 1936 2167
rect 2012 2163 2016 2167
rect 2092 2163 2096 2167
rect 2180 2163 2184 2167
rect 2216 2163 2220 2167
rect 2276 2163 2280 2167
rect 2356 2163 2360 2167
rect 1300 2151 1304 2155
rect 1348 2151 1352 2155
rect 1436 2151 1440 2155
rect 1532 2151 1536 2155
rect 1628 2151 1632 2155
rect 1724 2151 1728 2155
rect 1812 2151 1816 2155
rect 1892 2151 1896 2155
rect 1928 2151 1932 2155
rect 1972 2151 1976 2155
rect 2044 2151 2048 2155
rect 2108 2151 2112 2155
rect 2172 2151 2176 2155
rect 2236 2151 2240 2155
rect 2308 2151 2312 2155
rect 2356 2151 2360 2155
rect 1328 2115 1332 2119
rect 1376 2115 1380 2119
rect 1464 2115 1468 2119
rect 1560 2115 1564 2119
rect 1656 2115 1660 2119
rect 1752 2115 1756 2119
rect 1840 2115 1844 2119
rect 1920 2115 1924 2119
rect 1928 2115 1932 2119
rect 2000 2115 2004 2119
rect 2072 2115 2076 2119
rect 2136 2115 2140 2119
rect 2200 2115 2204 2119
rect 2264 2115 2268 2119
rect 2336 2115 2340 2119
rect 2384 2115 2388 2119
rect 408 2111 412 2115
rect 448 2111 452 2115
rect 488 2111 492 2115
rect 528 2111 532 2115
rect 576 2111 580 2115
rect 584 2111 588 2115
rect 632 2111 636 2115
rect 640 2111 644 2115
rect 688 2111 692 2115
rect 752 2111 756 2115
rect 816 2111 820 2115
rect 880 2111 884 2115
rect 936 2111 940 2115
rect 992 2111 996 2115
rect 1048 2111 1052 2115
rect 1104 2111 1108 2115
rect 1168 2111 1172 2115
rect 380 2075 384 2079
rect 420 2075 424 2079
rect 460 2075 464 2079
rect 500 2075 504 2079
rect 548 2075 552 2079
rect 584 2075 588 2079
rect 604 2075 608 2079
rect 640 2075 644 2079
rect 660 2075 664 2079
rect 724 2075 728 2079
rect 788 2075 792 2079
rect 852 2075 856 2079
rect 908 2075 912 2079
rect 964 2075 968 2079
rect 1020 2075 1024 2079
rect 1076 2075 1080 2079
rect 1140 2075 1144 2079
rect 380 2063 384 2067
rect 420 2063 424 2067
rect 460 2063 464 2067
rect 500 2063 504 2067
rect 540 2063 544 2067
rect 580 2063 584 2067
rect 628 2063 632 2067
rect 684 2063 688 2067
rect 728 2063 732 2067
rect 740 2063 744 2067
rect 796 2063 800 2067
rect 844 2063 848 2067
rect 900 2063 904 2067
rect 956 2063 960 2067
rect 1012 2063 1016 2067
rect 1068 2063 1072 2067
rect 1328 2059 1332 2063
rect 1368 2059 1372 2063
rect 1424 2059 1428 2063
rect 1504 2059 1508 2063
rect 1592 2059 1596 2063
rect 1688 2059 1692 2063
rect 1784 2059 1788 2063
rect 1792 2059 1796 2063
rect 1872 2059 1876 2063
rect 1960 2059 1964 2063
rect 2040 2059 2044 2063
rect 2120 2059 2124 2063
rect 2192 2059 2196 2063
rect 2264 2059 2268 2063
rect 2336 2059 2340 2063
rect 2344 2059 2348 2063
rect 2384 2059 2388 2063
rect 408 2027 412 2031
rect 448 2027 452 2031
rect 488 2027 492 2031
rect 528 2027 532 2031
rect 568 2027 572 2031
rect 608 2027 612 2031
rect 656 2027 660 2031
rect 664 2027 668 2031
rect 712 2027 716 2031
rect 728 2027 732 2031
rect 768 2027 772 2031
rect 824 2027 828 2031
rect 872 2027 876 2031
rect 928 2027 932 2031
rect 984 2027 988 2031
rect 1040 2027 1044 2031
rect 1096 2027 1100 2031
rect 392 1967 396 1971
rect 432 1967 436 1971
rect 480 1967 484 1971
rect 536 1967 540 1971
rect 544 1967 548 1971
rect 592 1967 596 1971
rect 656 1967 660 1971
rect 1300 2023 1304 2027
rect 1340 2023 1344 2027
rect 1396 2023 1400 2027
rect 1476 2023 1480 2027
rect 1564 2023 1568 2027
rect 1660 2023 1664 2027
rect 1756 2023 1760 2027
rect 1792 2023 1796 2027
rect 1844 2023 1848 2027
rect 1932 2023 1936 2027
rect 2012 2023 2016 2027
rect 2092 2023 2096 2027
rect 2164 2023 2168 2027
rect 2236 2023 2240 2027
rect 2308 2023 2312 2027
rect 2356 2023 2360 2027
rect 2344 2011 2348 2015
rect 1300 2003 1304 2007
rect 1348 2003 1352 2007
rect 1420 2003 1424 2007
rect 1492 2003 1496 2007
rect 1572 2005 1576 2009
rect 1660 2003 1664 2007
rect 1748 2003 1752 2007
rect 1836 2003 1840 2007
rect 1916 2003 1920 2007
rect 1996 2003 2000 2007
rect 2068 2003 2072 2007
rect 2132 2003 2136 2007
rect 2188 2003 2192 2007
rect 2252 2005 2256 2009
rect 2316 2003 2320 2007
rect 2356 2003 2360 2007
rect 720 1967 724 1971
rect 784 1967 788 1971
rect 840 1967 844 1971
rect 896 1967 900 1971
rect 960 1967 964 1971
rect 1024 1967 1028 1971
rect 1088 1967 1092 1971
rect 1328 1967 1332 1971
rect 1376 1967 1380 1971
rect 1448 1967 1452 1971
rect 1520 1967 1524 1971
rect 1600 1967 1604 1971
rect 1688 1967 1692 1971
rect 1776 1967 1780 1971
rect 1864 1967 1868 1971
rect 1944 1967 1948 1971
rect 2024 1967 2028 1971
rect 2064 1967 2068 1971
rect 2096 1967 2100 1971
rect 2160 1967 2164 1971
rect 2216 1967 2220 1971
rect 2280 1967 2284 1971
rect 2344 1967 2348 1971
rect 2384 1967 2388 1971
rect 364 1931 368 1935
rect 404 1931 408 1935
rect 452 1931 456 1935
rect 508 1931 512 1935
rect 544 1931 548 1935
rect 564 1931 568 1935
rect 628 1931 632 1935
rect 664 1931 668 1935
rect 692 1931 696 1935
rect 756 1931 760 1935
rect 812 1931 816 1935
rect 868 1931 872 1935
rect 932 1931 936 1935
rect 996 1931 1000 1935
rect 1060 1931 1064 1935
rect 172 1915 176 1919
rect 212 1915 216 1919
rect 248 1915 252 1919
rect 260 1915 264 1919
rect 316 1915 320 1919
rect 388 1915 392 1919
rect 456 1915 460 1919
rect 468 1915 472 1919
rect 548 1915 552 1919
rect 636 1915 640 1919
rect 672 1915 676 1919
rect 716 1915 720 1919
rect 796 1915 800 1919
rect 876 1917 880 1921
rect 956 1915 960 1919
rect 1036 1915 1040 1919
rect 1116 1915 1120 1919
rect 1328 1915 1332 1919
rect 1336 1915 1340 1919
rect 1384 1915 1388 1919
rect 1392 1915 1396 1919
rect 1472 1915 1476 1919
rect 1560 1915 1564 1919
rect 1608 1915 1612 1919
rect 1648 1915 1652 1919
rect 1736 1915 1740 1919
rect 1816 1915 1820 1919
rect 1888 1915 1892 1919
rect 1960 1915 1964 1919
rect 2032 1915 2036 1919
rect 456 1887 460 1891
rect 2104 1915 2108 1919
rect 2176 1915 2180 1919
rect 2248 1915 2252 1919
rect 2328 1915 2332 1919
rect 2384 1915 2388 1919
rect 200 1879 204 1883
rect 240 1879 244 1883
rect 248 1879 252 1883
rect 288 1879 292 1883
rect 344 1879 348 1883
rect 416 1879 420 1883
rect 496 1879 500 1883
rect 576 1879 580 1883
rect 664 1879 668 1883
rect 672 1879 676 1883
rect 744 1879 748 1883
rect 824 1879 828 1883
rect 904 1879 908 1883
rect 984 1879 988 1883
rect 1064 1879 1068 1883
rect 1144 1879 1148 1883
rect 1300 1879 1304 1883
rect 1336 1879 1340 1883
rect 1356 1879 1360 1883
rect 1392 1879 1396 1883
rect 1444 1879 1448 1883
rect 1532 1879 1536 1883
rect 1608 1879 1612 1883
rect 1620 1879 1624 1883
rect 1708 1879 1712 1883
rect 1788 1879 1792 1883
rect 1860 1879 1864 1883
rect 1932 1879 1936 1883
rect 2004 1879 2008 1883
rect 2064 1879 2068 1883
rect 2076 1879 2080 1883
rect 2148 1879 2152 1883
rect 2220 1879 2224 1883
rect 2300 1879 2304 1883
rect 2356 1879 2360 1883
rect 1308 1867 1312 1871
rect 1356 1867 1360 1871
rect 1412 1867 1416 1871
rect 1476 1867 1480 1871
rect 1528 1867 1532 1871
rect 1540 1867 1544 1871
rect 1612 1867 1616 1871
rect 1684 1867 1688 1871
rect 1764 1867 1768 1871
rect 1860 1867 1864 1871
rect 1928 1867 1932 1871
rect 1972 1867 1976 1871
rect 2008 1867 2012 1871
rect 2092 1867 2096 1871
rect 2220 1867 2224 1871
rect 2356 1867 2360 1871
rect 1928 1839 1932 1843
rect 1336 1831 1340 1835
rect 1384 1831 1388 1835
rect 1440 1831 1444 1835
rect 1504 1831 1508 1835
rect 1528 1831 1532 1835
rect 1568 1831 1572 1835
rect 1640 1831 1644 1835
rect 1712 1831 1716 1835
rect 1792 1831 1796 1835
rect 1888 1831 1892 1835
rect 2000 1831 2004 1835
rect 2008 1831 2012 1835
rect 2120 1831 2124 1835
rect 2248 1831 2252 1835
rect 2384 1831 2388 1835
rect 160 1819 164 1823
rect 200 1819 204 1823
rect 240 1819 244 1823
rect 248 1819 252 1823
rect 296 1819 300 1823
rect 376 1819 380 1823
rect 464 1819 468 1823
rect 560 1819 564 1823
rect 656 1819 660 1823
rect 664 1819 668 1823
rect 752 1819 756 1823
rect 760 1819 764 1823
rect 848 1819 852 1823
rect 936 1819 940 1823
rect 1016 1819 1020 1823
rect 1088 1819 1092 1823
rect 1160 1819 1164 1823
rect 1216 1819 1220 1823
rect 132 1783 136 1787
rect 172 1783 176 1787
rect 212 1783 216 1787
rect 248 1783 252 1787
rect 268 1783 272 1787
rect 348 1783 352 1787
rect 436 1783 440 1787
rect 532 1783 536 1787
rect 628 1783 632 1787
rect 664 1783 668 1787
rect 724 1783 728 1787
rect 760 1783 764 1787
rect 820 1783 824 1787
rect 908 1783 912 1787
rect 988 1783 992 1787
rect 1060 1783 1064 1787
rect 1132 1783 1136 1787
rect 1188 1783 1192 1787
rect 1432 1775 1436 1779
rect 1496 1775 1500 1779
rect 1560 1775 1564 1779
rect 1624 1775 1628 1779
rect 1688 1775 1692 1779
rect 1752 1775 1756 1779
rect 1808 1775 1812 1779
rect 1864 1775 1868 1779
rect 1920 1775 1924 1779
rect 1984 1775 1988 1779
rect 132 1771 136 1775
rect 172 1771 176 1775
rect 212 1771 216 1775
rect 284 1771 288 1775
rect 372 1771 376 1775
rect 468 1771 472 1775
rect 564 1771 568 1775
rect 660 1771 664 1775
rect 748 1771 752 1775
rect 828 1771 832 1775
rect 900 1771 904 1775
rect 964 1771 968 1775
rect 1028 1771 1032 1775
rect 1064 1771 1068 1775
rect 1084 1771 1088 1775
rect 1148 1771 1152 1775
rect 1188 1771 1192 1775
rect 1404 1739 1408 1743
rect 1468 1739 1472 1743
rect 1532 1739 1536 1743
rect 1596 1739 1600 1743
rect 1660 1739 1664 1743
rect 1724 1739 1728 1743
rect 1780 1739 1784 1743
rect 1836 1739 1840 1743
rect 1892 1739 1896 1743
rect 1956 1739 1960 1743
rect 160 1735 164 1739
rect 200 1735 204 1739
rect 240 1735 244 1739
rect 312 1735 316 1739
rect 400 1735 404 1739
rect 496 1735 500 1739
rect 592 1735 596 1739
rect 688 1735 692 1739
rect 776 1735 780 1739
rect 856 1735 860 1739
rect 928 1735 932 1739
rect 992 1735 996 1739
rect 1056 1735 1060 1739
rect 1064 1735 1068 1739
rect 1112 1735 1116 1739
rect 1176 1735 1180 1739
rect 1216 1735 1220 1739
rect 1300 1729 1304 1733
rect 1348 1727 1352 1731
rect 1420 1727 1424 1731
rect 1500 1727 1504 1731
rect 1580 1727 1584 1731
rect 1660 1727 1664 1731
rect 1704 1727 1708 1731
rect 1732 1727 1736 1731
rect 1804 1727 1808 1731
rect 1840 1727 1844 1731
rect 1868 1727 1872 1731
rect 1932 1727 1936 1731
rect 1996 1727 2000 1731
rect 2060 1727 2064 1731
rect 1328 1691 1332 1695
rect 1376 1691 1380 1695
rect 1448 1691 1452 1695
rect 1528 1691 1532 1695
rect 1608 1691 1612 1695
rect 1688 1691 1692 1695
rect 160 1679 164 1683
rect 200 1679 204 1683
rect 264 1679 268 1683
rect 344 1679 348 1683
rect 440 1679 444 1683
rect 536 1679 540 1683
rect 640 1679 644 1683
rect 736 1679 740 1683
rect 824 1679 828 1683
rect 904 1679 908 1683
rect 976 1679 980 1683
rect 1040 1679 1044 1683
rect 1112 1679 1116 1683
rect 1184 1679 1188 1683
rect 1760 1691 1764 1695
rect 1832 1691 1836 1695
rect 1840 1691 1844 1695
rect 1896 1693 1900 1697
rect 1960 1691 1964 1695
rect 2024 1691 2028 1695
rect 2088 1691 2092 1695
rect 1704 1647 1708 1651
rect 132 1643 136 1647
rect 172 1643 176 1647
rect 236 1643 240 1647
rect 316 1643 320 1647
rect 412 1643 416 1647
rect 508 1643 512 1647
rect 612 1643 616 1647
rect 708 1643 712 1647
rect 796 1643 800 1647
rect 876 1643 880 1647
rect 948 1643 952 1647
rect 1012 1643 1016 1647
rect 1084 1643 1088 1647
rect 1156 1643 1160 1647
rect 1328 1639 1332 1643
rect 1384 1639 1388 1643
rect 1472 1639 1476 1643
rect 1568 1639 1572 1643
rect 1664 1639 1668 1643
rect 1752 1639 1756 1643
rect 1840 1639 1844 1643
rect 1920 1639 1924 1643
rect 1992 1639 1996 1643
rect 2056 1639 2060 1643
rect 2120 1639 2124 1643
rect 2184 1639 2188 1643
rect 2248 1639 2252 1643
rect 268 1627 272 1631
rect 308 1627 312 1631
rect 356 1627 360 1631
rect 412 1627 416 1631
rect 468 1627 472 1631
rect 532 1627 536 1631
rect 596 1627 600 1631
rect 660 1629 664 1633
rect 716 1627 720 1631
rect 772 1627 776 1631
rect 828 1627 832 1631
rect 884 1627 888 1631
rect 940 1627 944 1631
rect 996 1627 1000 1631
rect 1300 1603 1304 1607
rect 1356 1603 1360 1607
rect 1444 1603 1448 1607
rect 1540 1603 1544 1607
rect 1636 1603 1640 1607
rect 1724 1603 1728 1607
rect 1812 1603 1816 1607
rect 1892 1603 1896 1607
rect 1964 1603 1968 1607
rect 2028 1603 2032 1607
rect 2092 1603 2096 1607
rect 2156 1603 2160 1607
rect 2220 1603 2224 1607
rect 296 1591 300 1595
rect 336 1591 340 1595
rect 384 1591 388 1595
rect 440 1591 444 1595
rect 496 1591 500 1595
rect 560 1591 564 1595
rect 624 1591 628 1595
rect 688 1591 692 1595
rect 744 1591 748 1595
rect 800 1591 804 1595
rect 856 1591 860 1595
rect 912 1591 916 1595
rect 968 1591 972 1595
rect 1024 1591 1028 1595
rect 1324 1591 1328 1595
rect 1396 1591 1400 1595
rect 1476 1591 1480 1595
rect 1564 1591 1568 1595
rect 1640 1591 1644 1595
rect 1652 1591 1656 1595
rect 1740 1591 1744 1595
rect 1816 1591 1820 1595
rect 1828 1591 1832 1595
rect 1880 1591 1884 1595
rect 1908 1591 1912 1595
rect 1980 1591 1984 1595
rect 2044 1591 2048 1595
rect 2108 1591 2112 1595
rect 2164 1591 2168 1595
rect 2212 1591 2216 1595
rect 2268 1591 2272 1595
rect 2316 1591 2320 1595
rect 2356 1591 2360 1595
rect 1352 1555 1356 1559
rect 1424 1555 1428 1559
rect 1504 1555 1508 1559
rect 1592 1555 1596 1559
rect 1640 1555 1644 1559
rect 1680 1555 1684 1559
rect 1768 1555 1772 1559
rect 1816 1555 1820 1559
rect 1856 1555 1860 1559
rect 352 1531 356 1535
rect 392 1531 396 1535
rect 432 1531 436 1535
rect 472 1531 476 1535
rect 512 1531 516 1535
rect 552 1531 556 1535
rect 592 1531 596 1535
rect 632 1531 636 1535
rect 672 1531 676 1535
rect 712 1531 716 1535
rect 752 1531 756 1535
rect 792 1531 796 1535
rect 832 1531 836 1535
rect 872 1531 876 1535
rect 912 1531 916 1535
rect 952 1531 956 1535
rect 1936 1555 1940 1559
rect 2008 1555 2012 1559
rect 2072 1555 2076 1559
rect 2136 1555 2140 1559
rect 2192 1555 2196 1559
rect 2240 1555 2244 1559
rect 2296 1555 2300 1559
rect 2344 1555 2348 1559
rect 2384 1555 2388 1559
rect 1880 1511 1884 1515
rect 1360 1499 1364 1503
rect 1440 1499 1444 1503
rect 1528 1499 1532 1503
rect 1640 1499 1644 1503
rect 1768 1499 1772 1503
rect 1872 1499 1876 1503
rect 1912 1499 1916 1503
rect 2072 1499 2076 1503
rect 2240 1499 2244 1503
rect 2384 1499 2388 1503
rect 324 1495 328 1499
rect 364 1495 368 1499
rect 404 1495 408 1499
rect 444 1495 448 1499
rect 484 1495 488 1499
rect 524 1495 528 1499
rect 564 1495 568 1499
rect 604 1495 608 1499
rect 644 1495 648 1499
rect 684 1495 688 1499
rect 724 1495 728 1499
rect 764 1495 768 1499
rect 804 1495 808 1499
rect 844 1495 848 1499
rect 884 1495 888 1499
rect 924 1495 928 1499
rect 1332 1463 1336 1467
rect 1412 1463 1416 1467
rect 1500 1463 1504 1467
rect 1612 1463 1616 1467
rect 1740 1463 1744 1467
rect 1872 1463 1876 1467
rect 1884 1463 1888 1467
rect 2044 1463 2048 1467
rect 2212 1463 2216 1467
rect 2356 1463 2360 1467
rect 1372 1451 1376 1455
rect 1460 1451 1464 1455
rect 1548 1451 1552 1455
rect 1636 1451 1640 1455
rect 1724 1451 1728 1455
rect 1804 1451 1808 1455
rect 1876 1451 1880 1455
rect 1940 1451 1944 1455
rect 1996 1451 2000 1455
rect 2044 1451 2048 1455
rect 2092 1451 2096 1455
rect 2140 1451 2144 1455
rect 2188 1451 2192 1455
rect 2236 1451 2240 1455
rect 2276 1451 2280 1455
rect 2316 1451 2320 1455
rect 2356 1451 2360 1455
rect 140 1443 144 1447
rect 180 1443 184 1447
rect 220 1443 224 1447
rect 260 1443 264 1447
rect 304 1443 308 1447
rect 316 1443 320 1447
rect 388 1443 392 1447
rect 468 1443 472 1447
rect 556 1443 560 1447
rect 644 1443 648 1447
rect 724 1443 728 1447
rect 804 1443 808 1447
rect 876 1443 880 1447
rect 940 1443 944 1447
rect 996 1443 1000 1447
rect 1044 1443 1048 1447
rect 1100 1443 1104 1447
rect 1148 1443 1152 1447
rect 1188 1443 1192 1447
rect 1400 1415 1404 1419
rect 1488 1415 1492 1419
rect 1576 1415 1580 1419
rect 1664 1415 1668 1419
rect 1752 1415 1756 1419
rect 1832 1415 1836 1419
rect 1904 1415 1908 1419
rect 1968 1415 1972 1419
rect 2024 1415 2028 1419
rect 2072 1415 2076 1419
rect 2120 1415 2124 1419
rect 2168 1415 2172 1419
rect 2216 1415 2220 1419
rect 2264 1415 2268 1419
rect 2304 1415 2308 1419
rect 2344 1415 2348 1419
rect 2384 1415 2388 1419
rect 168 1407 172 1411
rect 208 1407 212 1411
rect 248 1407 252 1411
rect 288 1407 292 1411
rect 304 1407 308 1411
rect 344 1407 348 1411
rect 416 1407 420 1411
rect 496 1407 500 1411
rect 584 1407 588 1411
rect 672 1407 676 1411
rect 752 1407 756 1411
rect 832 1407 836 1411
rect 904 1407 908 1411
rect 968 1407 972 1411
rect 1024 1407 1028 1411
rect 1072 1407 1076 1411
rect 1128 1407 1132 1411
rect 1176 1407 1180 1411
rect 1216 1407 1220 1411
rect 192 1355 196 1359
rect 232 1355 236 1359
rect 272 1355 276 1359
rect 328 1355 332 1359
rect 392 1355 396 1359
rect 464 1355 468 1359
rect 544 1355 548 1359
rect 624 1355 628 1359
rect 704 1355 708 1359
rect 776 1355 780 1359
rect 848 1355 852 1359
rect 912 1355 916 1359
rect 976 1355 980 1359
rect 1040 1355 1044 1359
rect 1104 1355 1108 1359
rect 1168 1355 1172 1359
rect 1216 1355 1220 1359
rect 1328 1355 1332 1359
rect 1368 1355 1372 1359
rect 1424 1355 1428 1359
rect 1488 1355 1492 1359
rect 1560 1355 1564 1359
rect 1568 1355 1572 1359
rect 1632 1355 1636 1359
rect 1640 1355 1644 1359
rect 1712 1355 1716 1359
rect 1792 1355 1796 1359
rect 1800 1355 1804 1359
rect 1872 1355 1876 1359
rect 1880 1355 1884 1359
rect 1960 1355 1964 1359
rect 2048 1355 2052 1359
rect 2136 1355 2140 1359
rect 2224 1355 2228 1359
rect 2312 1355 2316 1359
rect 2384 1355 2388 1359
rect 164 1319 168 1323
rect 204 1319 208 1323
rect 244 1319 248 1323
rect 300 1319 304 1323
rect 364 1319 368 1323
rect 436 1319 440 1323
rect 516 1319 520 1323
rect 596 1319 600 1323
rect 676 1319 680 1323
rect 748 1319 752 1323
rect 820 1319 824 1323
rect 884 1319 888 1323
rect 948 1319 952 1323
rect 1012 1319 1016 1323
rect 1076 1319 1080 1323
rect 1140 1319 1144 1323
rect 1188 1319 1192 1323
rect 1300 1319 1304 1323
rect 1340 1319 1344 1323
rect 1396 1319 1400 1323
rect 1460 1319 1464 1323
rect 1532 1319 1536 1323
rect 1568 1319 1572 1323
rect 1604 1319 1608 1323
rect 1640 1319 1644 1323
rect 1684 1319 1688 1323
rect 1764 1319 1768 1323
rect 1800 1319 1804 1323
rect 1844 1319 1848 1323
rect 1880 1319 1884 1323
rect 1932 1319 1936 1323
rect 2020 1319 2024 1323
rect 2108 1319 2112 1323
rect 2196 1319 2200 1323
rect 2284 1319 2288 1323
rect 2356 1319 2360 1323
rect 1300 1307 1304 1311
rect 1340 1307 1344 1311
rect 1380 1307 1384 1311
rect 1420 1307 1424 1311
rect 1460 1307 1464 1311
rect 1500 1307 1504 1311
rect 1540 1307 1544 1311
rect 1580 1307 1584 1311
rect 1620 1307 1624 1311
rect 1676 1307 1680 1311
rect 1720 1307 1724 1311
rect 1732 1307 1736 1311
rect 1788 1307 1792 1311
rect 1844 1307 1848 1311
rect 1900 1307 1904 1311
rect 1944 1307 1948 1311
rect 1964 1307 1968 1311
rect 2036 1307 2040 1311
rect 2116 1307 2120 1311
rect 2196 1307 2200 1311
rect 2284 1307 2288 1311
rect 2356 1307 2360 1311
rect 180 1303 184 1307
rect 228 1303 232 1307
rect 284 1303 288 1307
rect 348 1303 352 1307
rect 420 1303 424 1307
rect 492 1303 496 1307
rect 536 1303 540 1307
rect 564 1303 568 1307
rect 636 1303 640 1307
rect 700 1303 704 1307
rect 764 1303 768 1307
rect 820 1303 824 1307
rect 876 1303 880 1307
rect 932 1303 936 1307
rect 996 1303 1000 1307
rect 208 1267 212 1271
rect 256 1267 260 1271
rect 312 1267 316 1271
rect 376 1267 380 1271
rect 448 1267 452 1271
rect 520 1269 524 1273
rect 536 1271 540 1275
rect 1328 1271 1332 1275
rect 1368 1271 1372 1275
rect 1408 1271 1412 1275
rect 1448 1271 1452 1275
rect 1488 1271 1492 1275
rect 1528 1271 1532 1275
rect 1568 1271 1572 1275
rect 1608 1271 1612 1275
rect 1648 1271 1652 1275
rect 1704 1271 1708 1275
rect 1720 1271 1724 1275
rect 1760 1271 1764 1275
rect 1816 1271 1820 1275
rect 1872 1271 1876 1275
rect 1928 1271 1932 1275
rect 1944 1271 1948 1275
rect 1992 1271 1996 1275
rect 2064 1271 2068 1275
rect 2144 1271 2148 1275
rect 2224 1271 2228 1275
rect 2312 1271 2316 1275
rect 2384 1271 2388 1275
rect 592 1267 596 1271
rect 664 1267 668 1271
rect 728 1267 732 1271
rect 792 1267 796 1271
rect 848 1267 852 1271
rect 904 1267 908 1271
rect 960 1267 964 1271
rect 1024 1267 1028 1271
rect 160 1211 164 1215
rect 200 1211 204 1215
rect 256 1211 260 1215
rect 264 1211 268 1215
rect 336 1211 340 1215
rect 344 1211 348 1215
rect 424 1211 428 1215
rect 432 1211 436 1215
rect 512 1211 516 1215
rect 520 1211 524 1215
rect 600 1211 604 1215
rect 688 1211 692 1215
rect 768 1211 772 1215
rect 776 1211 780 1215
rect 840 1211 844 1215
rect 848 1211 852 1215
rect 904 1211 908 1215
rect 912 1211 916 1215
rect 968 1211 972 1215
rect 976 1211 980 1215
rect 1032 1211 1036 1215
rect 1040 1211 1044 1215
rect 1096 1211 1100 1215
rect 1328 1211 1332 1215
rect 1336 1211 1340 1215
rect 1400 1211 1404 1215
rect 1408 1211 1412 1215
rect 1504 1211 1508 1215
rect 1608 1211 1612 1215
rect 1712 1211 1716 1215
rect 1816 1211 1820 1215
rect 1912 1211 1916 1215
rect 2008 1211 2012 1215
rect 2096 1211 2100 1215
rect 2176 1211 2180 1215
rect 2248 1211 2252 1215
rect 2328 1211 2332 1215
rect 2384 1211 2388 1215
rect 132 1175 136 1179
rect 172 1175 176 1179
rect 228 1175 232 1179
rect 308 1175 312 1179
rect 344 1175 348 1179
rect 396 1175 400 1179
rect 432 1175 436 1179
rect 484 1175 488 1179
rect 520 1175 524 1179
rect 572 1175 576 1179
rect 660 1175 664 1179
rect 740 1175 744 1179
rect 776 1175 780 1179
rect 812 1175 816 1179
rect 848 1175 852 1179
rect 876 1175 880 1179
rect 912 1175 916 1179
rect 940 1175 944 1179
rect 976 1175 980 1179
rect 1004 1175 1008 1179
rect 1040 1175 1044 1179
rect 1068 1175 1072 1179
rect 1300 1175 1304 1179
rect 1336 1175 1340 1179
rect 1372 1175 1376 1179
rect 1408 1175 1412 1179
rect 1476 1175 1480 1179
rect 1580 1175 1584 1179
rect 1684 1175 1688 1179
rect 1788 1175 1792 1179
rect 1884 1175 1888 1179
rect 1980 1175 1984 1179
rect 2068 1175 2072 1179
rect 2148 1175 2152 1179
rect 2220 1175 2224 1179
rect 2300 1175 2304 1179
rect 2356 1175 2360 1179
rect 132 1163 136 1167
rect 172 1163 176 1167
rect 236 1165 240 1169
rect 264 1167 268 1171
rect 272 1163 276 1167
rect 324 1163 328 1167
rect 428 1163 432 1167
rect 532 1163 536 1167
rect 636 1163 640 1167
rect 740 1163 744 1167
rect 836 1163 840 1167
rect 916 1163 920 1167
rect 996 1163 1000 1167
rect 1068 1163 1072 1167
rect 1140 1163 1144 1167
rect 1188 1163 1192 1167
rect 1300 1163 1304 1167
rect 1340 1163 1344 1167
rect 1384 1163 1388 1167
rect 1404 1163 1408 1167
rect 1484 1163 1488 1167
rect 1580 1163 1584 1167
rect 1684 1163 1688 1167
rect 1796 1163 1800 1167
rect 1900 1163 1904 1167
rect 1996 1163 2000 1167
rect 2076 1163 2080 1167
rect 2156 1163 2160 1167
rect 2216 1163 2220 1167
rect 2228 1163 2232 1167
rect 2300 1163 2304 1167
rect 2356 1163 2360 1167
rect 160 1127 164 1131
rect 200 1127 204 1131
rect 264 1127 268 1131
rect 272 1127 276 1131
rect 352 1127 356 1131
rect 456 1127 460 1131
rect 560 1127 564 1131
rect 664 1127 668 1131
rect 768 1127 772 1131
rect 864 1127 868 1131
rect 944 1127 948 1131
rect 1024 1127 1028 1131
rect 1096 1127 1100 1131
rect 1168 1127 1172 1131
rect 1216 1127 1220 1131
rect 1328 1127 1332 1131
rect 1368 1127 1372 1131
rect 1384 1127 1388 1131
rect 1432 1127 1436 1131
rect 1512 1127 1516 1131
rect 1608 1127 1612 1131
rect 1712 1127 1716 1131
rect 1824 1127 1828 1131
rect 1928 1127 1932 1131
rect 2024 1127 2028 1131
rect 2104 1127 2108 1131
rect 2184 1127 2188 1131
rect 2216 1127 2220 1131
rect 2256 1127 2260 1131
rect 2328 1127 2332 1131
rect 2384 1127 2388 1131
rect 1456 1075 1460 1079
rect 1496 1075 1500 1079
rect 1536 1075 1540 1079
rect 1584 1075 1588 1079
rect 1640 1075 1644 1079
rect 1696 1075 1700 1079
rect 1752 1075 1756 1079
rect 1800 1075 1804 1079
rect 1848 1075 1852 1079
rect 1856 1075 1860 1079
rect 1896 1075 1900 1079
rect 1904 1075 1908 1079
rect 1944 1075 1948 1079
rect 1952 1075 1956 1079
rect 1992 1075 1996 1079
rect 2040 1075 2044 1079
rect 2048 1075 2052 1079
rect 2088 1075 2092 1079
rect 2096 1075 2100 1079
rect 2144 1075 2148 1079
rect 2200 1075 2204 1079
rect 2256 1075 2260 1079
rect 160 1071 164 1075
rect 200 1071 204 1075
rect 272 1071 276 1075
rect 352 1071 356 1075
rect 440 1071 444 1075
rect 528 1071 532 1075
rect 568 1071 572 1075
rect 608 1071 612 1075
rect 688 1071 692 1075
rect 760 1071 764 1075
rect 824 1071 828 1075
rect 888 1071 892 1075
rect 944 1071 948 1075
rect 1008 1071 1012 1075
rect 1072 1071 1076 1075
rect 1428 1039 1432 1043
rect 1468 1039 1472 1043
rect 1508 1039 1512 1043
rect 1556 1039 1560 1043
rect 1612 1039 1616 1043
rect 1668 1039 1672 1043
rect 1724 1039 1728 1043
rect 1772 1039 1776 1043
rect 1820 1039 1824 1043
rect 1856 1039 1860 1043
rect 1868 1039 1872 1043
rect 1904 1039 1908 1043
rect 1916 1039 1920 1043
rect 1952 1039 1956 1043
rect 1964 1039 1968 1043
rect 2012 1039 2016 1043
rect 2048 1039 2052 1043
rect 2060 1039 2064 1043
rect 2096 1039 2100 1043
rect 2116 1039 2120 1043
rect 2172 1039 2176 1043
rect 2228 1039 2232 1043
rect 132 1035 136 1039
rect 172 1035 176 1039
rect 244 1035 248 1039
rect 324 1035 328 1039
rect 412 1035 416 1039
rect 500 1035 504 1039
rect 568 1035 572 1039
rect 580 1035 584 1039
rect 660 1035 664 1039
rect 732 1035 736 1039
rect 796 1035 800 1039
rect 860 1035 864 1039
rect 916 1035 920 1039
rect 980 1035 984 1039
rect 1044 1035 1048 1039
rect 1572 1027 1576 1031
rect 1612 1027 1616 1031
rect 1652 1027 1656 1031
rect 1692 1027 1696 1031
rect 1732 1027 1736 1031
rect 1772 1027 1776 1031
rect 1820 1027 1824 1031
rect 1876 1027 1880 1031
rect 1940 1027 1944 1031
rect 1984 1027 1988 1031
rect 2012 1027 2016 1031
rect 2092 1027 2096 1031
rect 2172 1027 2176 1031
rect 2252 1027 2256 1031
rect 172 1023 176 1027
rect 252 1023 256 1027
rect 324 1023 328 1027
rect 396 1023 400 1027
rect 460 1023 464 1027
rect 516 1023 520 1027
rect 572 1023 576 1027
rect 620 1023 624 1027
rect 668 1023 672 1027
rect 732 1023 736 1027
rect 804 1023 808 1027
rect 892 1023 896 1027
rect 996 1023 1000 1027
rect 1100 1023 1104 1027
rect 1188 1023 1192 1027
rect 1600 991 1604 995
rect 1640 991 1644 995
rect 1680 991 1684 995
rect 1720 991 1724 995
rect 1760 991 1764 995
rect 1800 991 1804 995
rect 1848 991 1852 995
rect 1904 991 1908 995
rect 1968 993 1972 997
rect 1984 995 1988 999
rect 1992 991 1996 995
rect 2040 991 2044 995
rect 2120 991 2124 995
rect 2200 991 2204 995
rect 2280 991 2284 995
rect 200 987 204 991
rect 280 987 284 991
rect 352 987 356 991
rect 424 987 428 991
rect 488 987 492 991
rect 544 987 548 991
rect 600 987 604 991
rect 648 987 652 991
rect 696 987 700 991
rect 760 987 764 991
rect 832 987 836 991
rect 920 987 924 991
rect 1024 987 1028 991
rect 1128 987 1132 991
rect 1216 987 1220 991
rect 240 935 244 939
rect 280 935 284 939
rect 328 935 332 939
rect 384 935 388 939
rect 392 935 396 939
rect 440 935 444 939
rect 488 935 492 939
rect 544 935 548 939
rect 600 935 604 939
rect 664 935 668 939
rect 736 935 740 939
rect 808 935 812 939
rect 880 935 884 939
rect 952 935 956 939
rect 1024 935 1028 939
rect 1096 935 1100 939
rect 1104 935 1108 939
rect 1168 935 1172 939
rect 1216 935 1220 939
rect 1328 931 1332 935
rect 1336 931 1340 935
rect 1376 931 1380 935
rect 1384 931 1388 935
rect 1456 931 1460 935
rect 1464 931 1468 935
rect 1536 931 1540 935
rect 1616 931 1620 935
rect 1656 931 1660 935
rect 1704 931 1708 935
rect 1792 931 1796 935
rect 1800 931 1804 935
rect 1880 931 1884 935
rect 1888 931 1892 935
rect 1968 931 1972 935
rect 212 899 216 903
rect 252 899 256 903
rect 300 899 304 903
rect 356 899 360 903
rect 392 899 396 903
rect 412 899 416 903
rect 460 899 464 903
rect 516 899 520 903
rect 572 899 576 903
rect 636 899 640 903
rect 708 899 712 903
rect 780 899 784 903
rect 852 899 856 903
rect 924 899 928 903
rect 996 899 1000 903
rect 1068 899 1072 903
rect 1104 899 1108 903
rect 1140 899 1144 903
rect 1188 899 1192 903
rect 2048 931 2052 935
rect 2128 931 2132 935
rect 2208 931 2212 935
rect 2296 931 2300 935
rect 1300 895 1304 899
rect 1336 895 1340 899
rect 1348 895 1352 899
rect 1384 895 1388 899
rect 1428 895 1432 899
rect 1464 895 1468 899
rect 1508 895 1512 899
rect 1588 895 1592 899
rect 1656 895 1660 899
rect 1676 895 1680 899
rect 1764 895 1768 899
rect 1800 895 1804 899
rect 1852 895 1856 899
rect 1888 895 1892 899
rect 1940 895 1944 899
rect 1992 895 1996 899
rect 2020 895 2024 899
rect 2100 895 2104 899
rect 2180 895 2184 899
rect 2268 895 2272 899
rect 188 881 192 885
rect 1436 883 1440 887
rect 1476 883 1480 887
rect 1516 883 1520 887
rect 1556 883 1560 887
rect 1592 883 1596 887
rect 1604 883 1608 887
rect 1652 883 1656 887
rect 1688 883 1692 887
rect 1708 883 1712 887
rect 1772 883 1776 887
rect 1844 883 1848 887
rect 1916 883 1920 887
rect 1968 883 1972 887
rect 1988 883 1992 887
rect 2060 883 2064 887
rect 2132 883 2136 887
rect 2212 883 2216 887
rect 2292 883 2296 887
rect 228 879 232 883
rect 284 879 288 883
rect 336 879 340 883
rect 356 879 360 883
rect 444 879 448 883
rect 540 879 544 883
rect 636 879 640 883
rect 724 879 728 883
rect 804 879 808 883
rect 884 879 888 883
rect 956 879 960 883
rect 1020 879 1024 883
rect 1084 879 1088 883
rect 1156 879 1160 883
rect 1464 847 1468 851
rect 1504 847 1508 851
rect 1544 847 1548 851
rect 1584 847 1588 851
rect 1592 847 1596 851
rect 1632 847 1636 851
rect 1680 849 1684 853
rect 1688 851 1692 855
rect 1736 847 1740 851
rect 1800 847 1804 851
rect 1872 847 1876 851
rect 1944 849 1948 853
rect 1968 851 1972 855
rect 2016 847 2020 851
rect 2088 847 2092 851
rect 2160 847 2164 851
rect 2240 847 2244 851
rect 2320 847 2324 851
rect 216 843 220 847
rect 256 843 260 847
rect 312 843 316 847
rect 336 843 340 847
rect 384 843 388 847
rect 472 843 476 847
rect 568 843 572 847
rect 664 843 668 847
rect 752 843 756 847
rect 832 843 836 847
rect 912 843 916 847
rect 984 843 988 847
rect 1048 843 1052 847
rect 1112 843 1116 847
rect 1184 843 1188 847
rect 160 791 164 795
rect 200 791 204 795
rect 264 791 268 795
rect 352 791 356 795
rect 440 791 444 795
rect 528 791 532 795
rect 616 791 620 795
rect 696 791 700 795
rect 768 791 772 795
rect 840 791 844 795
rect 904 791 908 795
rect 968 791 972 795
rect 1040 791 1044 795
rect 1384 783 1388 787
rect 1440 783 1444 787
rect 1496 783 1500 787
rect 1560 783 1564 787
rect 1616 783 1620 787
rect 1672 783 1676 787
rect 1728 783 1732 787
rect 1784 783 1788 787
rect 1840 783 1844 787
rect 1896 783 1900 787
rect 1960 783 1964 787
rect 2024 783 2028 787
rect 2096 783 2100 787
rect 2168 783 2172 787
rect 2248 783 2252 787
rect 2328 783 2332 787
rect 2384 783 2388 787
rect 132 755 136 759
rect 172 755 176 759
rect 236 755 240 759
rect 324 755 328 759
rect 412 755 416 759
rect 500 755 504 759
rect 588 755 592 759
rect 668 755 672 759
rect 740 755 744 759
rect 812 755 816 759
rect 876 755 880 759
rect 940 755 944 759
rect 1012 755 1016 759
rect 1356 747 1360 751
rect 1412 747 1416 751
rect 1468 747 1472 751
rect 1532 747 1536 751
rect 1588 747 1592 751
rect 1644 747 1648 751
rect 1700 747 1704 751
rect 1756 747 1760 751
rect 1812 747 1816 751
rect 1868 747 1872 751
rect 1932 747 1936 751
rect 1996 747 2000 751
rect 2068 747 2072 751
rect 2140 747 2144 751
rect 2220 747 2224 751
rect 2300 747 2304 751
rect 2356 747 2360 751
rect 132 739 136 743
rect 176 739 180 743
rect 188 739 192 743
rect 260 739 264 743
rect 320 739 324 743
rect 332 739 336 743
rect 396 739 400 743
rect 452 739 456 743
rect 500 739 504 743
rect 540 739 544 743
rect 580 739 584 743
rect 620 739 624 743
rect 668 739 672 743
rect 716 739 720 743
rect 764 739 768 743
rect 812 739 816 743
rect 860 739 864 743
rect 908 739 912 743
rect 1300 735 1304 739
rect 1340 735 1344 739
rect 1404 735 1408 739
rect 1484 735 1488 739
rect 1572 735 1576 739
rect 1660 735 1664 739
rect 1748 735 1752 739
rect 1828 735 1832 739
rect 1908 735 1912 739
rect 1988 735 1992 739
rect 2076 735 2080 739
rect 2172 735 2176 739
rect 2276 735 2280 739
rect 2356 735 2360 739
rect 160 703 164 707
rect 176 703 180 707
rect 216 703 220 707
rect 288 703 292 707
rect 320 703 324 707
rect 360 703 364 707
rect 424 703 428 707
rect 480 703 484 707
rect 528 703 532 707
rect 568 703 572 707
rect 608 703 612 707
rect 648 703 652 707
rect 696 703 700 707
rect 744 705 748 709
rect 792 703 796 707
rect 840 703 844 707
rect 888 703 892 707
rect 936 703 940 707
rect 1328 699 1332 703
rect 1368 699 1372 703
rect 1432 699 1436 703
rect 1512 699 1516 703
rect 1600 699 1604 703
rect 1688 699 1692 703
rect 1776 699 1780 703
rect 1856 699 1860 703
rect 1936 699 1940 703
rect 2016 699 2020 703
rect 2104 699 2108 703
rect 2200 699 2204 703
rect 2304 699 2308 703
rect 2384 699 2388 703
rect 160 647 164 651
rect 224 647 228 651
rect 304 647 308 651
rect 376 647 380 651
rect 440 647 444 651
rect 512 647 516 651
rect 584 647 588 651
rect 664 647 668 651
rect 672 647 676 651
rect 736 647 740 651
rect 744 647 748 651
rect 808 647 812 651
rect 880 647 884 651
rect 944 647 948 651
rect 1008 647 1012 651
rect 1064 647 1068 651
rect 1120 647 1124 651
rect 1176 647 1180 651
rect 1216 647 1220 651
rect 1328 643 1332 647
rect 1424 643 1428 647
rect 1536 643 1540 647
rect 1648 643 1652 647
rect 1656 643 1660 647
rect 1752 643 1756 647
rect 1840 643 1844 647
rect 1920 643 1924 647
rect 2000 643 2004 647
rect 2072 643 2076 647
rect 2080 643 2084 647
rect 2136 643 2140 647
rect 2144 643 2148 647
rect 2200 643 2204 647
rect 2208 643 2212 647
rect 2264 643 2268 647
rect 2336 643 2340 647
rect 2384 643 2388 647
rect 132 611 136 615
rect 196 611 200 615
rect 276 611 280 615
rect 348 611 352 615
rect 412 611 416 615
rect 484 611 488 615
rect 556 611 560 615
rect 636 611 640 615
rect 672 611 676 615
rect 708 611 712 615
rect 744 611 748 615
rect 780 611 784 615
rect 852 611 856 615
rect 916 611 920 615
rect 980 611 984 615
rect 1036 611 1040 615
rect 1092 611 1096 615
rect 1148 611 1152 615
rect 1188 611 1192 615
rect 1300 607 1304 611
rect 1396 607 1400 611
rect 1508 607 1512 611
rect 1620 607 1624 611
rect 1656 607 1660 611
rect 1724 607 1728 611
rect 1812 607 1816 611
rect 1892 607 1896 611
rect 1972 607 1976 611
rect 2044 607 2048 611
rect 2080 607 2084 611
rect 2108 607 2112 611
rect 2144 607 2148 611
rect 2172 607 2176 611
rect 2208 607 2212 611
rect 2236 607 2240 611
rect 2308 607 2312 611
rect 2356 607 2360 611
rect 132 591 136 595
rect 188 591 192 595
rect 268 591 272 595
rect 356 591 360 595
rect 444 591 448 595
rect 532 591 536 595
rect 620 591 624 595
rect 700 591 704 595
rect 780 591 784 595
rect 852 591 856 595
rect 916 591 920 595
rect 972 591 976 595
rect 1020 591 1024 595
rect 1076 591 1080 595
rect 1132 591 1136 595
rect 1188 591 1192 595
rect 1412 591 1416 595
rect 1452 591 1456 595
rect 1492 591 1496 595
rect 1540 591 1544 595
rect 1596 591 1600 595
rect 1660 591 1664 595
rect 1724 591 1728 595
rect 1788 591 1792 595
rect 1824 591 1828 595
rect 1824 567 1828 571
rect 1832 591 1836 595
rect 1844 591 1848 595
rect 1908 591 1912 595
rect 1952 591 1956 595
rect 1972 591 1976 595
rect 2044 591 2048 595
rect 2116 591 2120 595
rect 2196 591 2200 595
rect 2284 591 2288 595
rect 2356 591 2360 595
rect 160 555 164 559
rect 216 555 220 559
rect 296 555 300 559
rect 384 555 388 559
rect 472 555 476 559
rect 560 555 564 559
rect 648 555 652 559
rect 728 555 732 559
rect 808 555 812 559
rect 880 555 884 559
rect 944 555 948 559
rect 1000 555 1004 559
rect 1048 555 1052 559
rect 1104 555 1108 559
rect 1160 555 1164 559
rect 1216 555 1220 559
rect 1440 555 1444 559
rect 1480 555 1484 559
rect 1520 555 1524 559
rect 1568 555 1572 559
rect 1624 557 1628 561
rect 1688 555 1692 559
rect 1752 555 1756 559
rect 1816 557 1820 561
rect 1832 559 1836 563
rect 1872 555 1876 559
rect 1936 555 1940 559
rect 1952 555 1956 559
rect 2000 555 2004 559
rect 2072 555 2076 559
rect 2144 555 2148 559
rect 2224 555 2228 559
rect 2312 555 2316 559
rect 2384 555 2388 559
rect 1328 503 1332 507
rect 1400 503 1404 507
rect 1408 503 1412 507
rect 1504 503 1508 507
rect 1512 503 1516 507
rect 1608 503 1612 507
rect 1720 503 1724 507
rect 1824 503 1828 507
rect 1928 503 1932 507
rect 2032 503 2036 507
rect 2128 503 2132 507
rect 2216 503 2220 507
rect 2312 503 2316 507
rect 2384 503 2388 507
rect 160 495 164 499
rect 176 495 180 499
rect 216 495 220 499
rect 288 495 292 499
rect 360 495 364 499
rect 368 495 372 499
rect 440 495 444 499
rect 448 495 452 499
rect 520 495 524 499
rect 528 495 532 499
rect 600 495 604 499
rect 672 495 676 499
rect 744 495 748 499
rect 768 495 772 499
rect 808 495 812 499
rect 872 495 876 499
rect 928 495 932 499
rect 984 495 988 499
rect 1048 495 1052 499
rect 1112 495 1116 499
rect 1176 495 1180 499
rect 1216 495 1220 499
rect 132 459 136 463
rect 168 459 172 463
rect 176 459 180 463
rect 188 459 192 463
rect 260 459 264 463
rect 332 459 336 463
rect 368 459 372 463
rect 412 459 416 463
rect 448 459 452 463
rect 492 459 496 463
rect 528 459 532 463
rect 572 461 576 465
rect 1300 467 1304 471
rect 1372 467 1376 471
rect 1408 467 1412 471
rect 1476 467 1480 471
rect 1512 467 1516 471
rect 1580 467 1584 471
rect 1692 467 1696 471
rect 1796 467 1800 471
rect 1900 467 1904 471
rect 2004 467 2008 471
rect 2100 467 2104 471
rect 2188 467 2192 471
rect 2284 467 2288 471
rect 2356 467 2360 471
rect 644 459 648 463
rect 716 459 720 463
rect 768 459 772 463
rect 780 459 784 463
rect 844 459 848 463
rect 900 459 904 463
rect 956 459 960 463
rect 1020 459 1024 463
rect 1084 459 1088 463
rect 1148 459 1152 463
rect 1188 459 1192 463
rect 1300 451 1304 455
rect 1340 451 1344 455
rect 1376 451 1380 455
rect 1396 451 1400 455
rect 1460 451 1464 455
rect 1524 451 1528 455
rect 1588 451 1592 455
rect 1660 451 1664 455
rect 1732 451 1736 455
rect 1812 451 1816 455
rect 1892 451 1896 455
rect 1972 451 1976 455
rect 2052 451 2056 455
rect 2132 451 2136 455
rect 2212 451 2216 455
rect 2292 451 2296 455
rect 2336 451 2340 455
rect 2356 451 2360 455
rect 180 447 184 451
rect 220 447 224 451
rect 260 447 264 451
rect 308 447 312 451
rect 364 447 368 451
rect 428 447 432 451
rect 492 447 496 451
rect 556 447 560 451
rect 612 447 616 451
rect 648 447 652 451
rect 668 447 672 451
rect 716 447 720 451
rect 760 447 764 451
rect 772 447 776 451
rect 828 447 832 451
rect 884 447 888 451
rect 2336 423 2340 427
rect 1328 415 1332 419
rect 1368 415 1372 419
rect 1376 415 1380 419
rect 1424 415 1428 419
rect 1488 415 1492 419
rect 1552 415 1556 419
rect 1616 415 1620 419
rect 1688 415 1692 419
rect 1760 415 1764 419
rect 1840 415 1844 419
rect 1920 415 1924 419
rect 2000 415 2004 419
rect 2080 415 2084 419
rect 2160 415 2164 419
rect 2240 415 2244 419
rect 2320 415 2324 419
rect 2384 415 2388 419
rect 168 411 172 415
rect 208 411 212 415
rect 248 411 252 415
rect 288 411 292 415
rect 336 411 340 415
rect 392 411 396 415
rect 456 411 460 415
rect 520 411 524 415
rect 584 411 588 415
rect 640 411 644 415
rect 648 411 652 415
rect 696 411 700 415
rect 744 411 748 415
rect 760 411 764 415
rect 800 411 804 415
rect 856 411 860 415
rect 912 411 916 415
rect 160 359 164 363
rect 200 359 204 363
rect 256 359 260 363
rect 312 359 316 363
rect 368 359 372 363
rect 376 359 380 363
rect 416 359 420 363
rect 424 359 428 363
rect 464 359 468 363
rect 512 359 516 363
rect 560 359 564 363
rect 608 359 612 363
rect 656 359 660 363
rect 704 359 708 363
rect 752 359 756 363
rect 800 359 804 363
rect 1472 359 1476 363
rect 1512 359 1516 363
rect 1560 359 1564 363
rect 1616 359 1620 363
rect 1688 359 1692 363
rect 1760 359 1764 363
rect 1840 359 1844 363
rect 1920 359 1924 363
rect 1992 359 1996 363
rect 2064 359 2068 363
rect 2136 359 2140 363
rect 2144 359 2148 363
rect 2200 359 2204 363
rect 2208 359 2212 363
rect 2264 359 2268 363
rect 2272 359 2276 363
rect 2328 359 2332 363
rect 2384 359 2388 363
rect 132 323 136 327
rect 172 323 176 327
rect 228 323 232 327
rect 284 323 288 327
rect 340 323 344 327
rect 376 323 380 327
rect 388 323 392 327
rect 424 323 428 327
rect 436 323 440 327
rect 484 323 488 327
rect 532 323 536 327
rect 580 323 584 327
rect 628 323 632 327
rect 676 323 680 327
rect 724 323 728 327
rect 772 323 776 327
rect 1444 323 1448 327
rect 1484 323 1488 327
rect 1532 323 1536 327
rect 1588 323 1592 327
rect 1660 323 1664 327
rect 1732 323 1736 327
rect 1812 323 1816 327
rect 1892 323 1896 327
rect 1964 323 1968 327
rect 2036 323 2040 327
rect 2108 323 2112 327
rect 2144 323 2148 327
rect 2172 323 2176 327
rect 2208 323 2212 327
rect 2236 323 2240 327
rect 2272 323 2276 327
rect 2300 323 2304 327
rect 2356 323 2360 327
rect 132 307 136 311
rect 180 307 184 311
rect 252 307 256 311
rect 324 307 328 311
rect 388 307 392 311
rect 444 307 448 311
rect 500 307 504 311
rect 536 307 540 311
rect 548 307 552 311
rect 588 307 592 311
rect 628 307 632 311
rect 676 307 680 311
rect 724 307 728 311
rect 772 307 776 311
rect 820 307 824 311
rect 868 307 872 311
rect 916 307 920 311
rect 1492 309 1496 313
rect 1532 307 1536 311
rect 1572 307 1576 311
rect 1612 307 1616 311
rect 1652 307 1656 311
rect 1692 307 1696 311
rect 1740 307 1744 311
rect 1796 309 1800 313
rect 1860 307 1864 311
rect 1896 307 1900 311
rect 1932 307 1936 311
rect 2004 307 2008 311
rect 2068 307 2072 311
rect 2132 307 2136 311
rect 2188 307 2192 311
rect 2252 307 2256 311
rect 2316 307 2320 311
rect 2356 307 2360 311
rect 160 271 164 275
rect 208 271 212 275
rect 280 271 284 275
rect 352 271 356 275
rect 416 271 420 275
rect 472 271 476 275
rect 528 271 532 275
rect 536 271 540 275
rect 576 271 580 275
rect 616 271 620 275
rect 656 271 660 275
rect 704 271 708 275
rect 752 271 756 275
rect 800 271 804 275
rect 848 271 852 275
rect 896 271 900 275
rect 944 271 948 275
rect 1520 271 1524 275
rect 1560 271 1564 275
rect 1600 271 1604 275
rect 1640 271 1644 275
rect 1680 271 1684 275
rect 1720 271 1724 275
rect 1768 271 1772 275
rect 1824 271 1828 275
rect 1888 271 1892 275
rect 1896 271 1900 275
rect 1960 271 1964 275
rect 2032 271 2036 275
rect 2096 271 2100 275
rect 2160 271 2164 275
rect 2216 271 2220 275
rect 2280 271 2284 275
rect 2344 271 2348 275
rect 2384 271 2388 275
rect 1392 215 1396 219
rect 1432 215 1436 219
rect 1472 215 1476 219
rect 1520 215 1524 219
rect 1528 215 1532 219
rect 1576 215 1580 219
rect 1584 215 1588 219
rect 1632 215 1636 219
rect 1696 215 1700 219
rect 1760 215 1764 219
rect 1832 215 1836 219
rect 1912 215 1916 219
rect 2000 215 2004 219
rect 2096 215 2100 219
rect 2104 215 2108 219
rect 2192 215 2196 219
rect 2200 215 2204 219
rect 2296 215 2300 219
rect 2384 215 2388 219
rect 160 211 164 215
rect 200 211 204 215
rect 272 211 276 215
rect 352 211 356 215
rect 440 211 444 215
rect 520 211 524 215
rect 600 211 604 215
rect 680 211 684 215
rect 752 211 756 215
rect 816 211 820 215
rect 872 211 876 215
rect 928 211 932 215
rect 984 211 988 215
rect 1048 211 1052 215
rect 1364 179 1368 183
rect 1404 179 1408 183
rect 1444 179 1448 183
rect 1492 179 1496 183
rect 1528 179 1532 183
rect 1548 179 1552 183
rect 1584 179 1588 183
rect 1604 179 1608 183
rect 1668 179 1672 183
rect 1732 179 1736 183
rect 1804 179 1808 183
rect 1884 179 1888 183
rect 1972 179 1976 183
rect 2068 179 2072 183
rect 2104 179 2108 183
rect 2164 179 2168 183
rect 2200 179 2204 183
rect 2268 179 2272 183
rect 2356 179 2360 183
rect 132 175 136 179
rect 172 175 176 179
rect 244 175 248 179
rect 324 175 328 179
rect 412 175 416 179
rect 492 175 496 179
rect 572 175 576 179
rect 652 175 656 179
rect 724 175 728 179
rect 788 175 792 179
rect 844 175 848 179
rect 900 175 904 179
rect 956 175 960 179
rect 1020 175 1024 179
rect 1300 151 1304 155
rect 1340 151 1344 155
rect 1380 151 1384 155
rect 1420 151 1424 155
rect 1460 151 1464 155
rect 1516 151 1520 155
rect 1552 151 1556 155
rect 1580 151 1584 155
rect 1616 151 1620 155
rect 1644 151 1648 155
rect 1708 153 1712 157
rect 1752 151 1756 155
rect 1764 151 1768 155
rect 1800 151 1804 155
rect 1820 151 1824 155
rect 1868 151 1872 155
rect 1916 151 1920 155
rect 1964 151 1968 155
rect 2012 151 2016 155
rect 2060 151 2064 155
rect 2108 151 2112 155
rect 2156 151 2160 155
rect 2212 151 2216 155
rect 2268 151 2272 155
rect 2316 151 2320 155
rect 2356 151 2360 155
rect 132 143 136 147
rect 172 143 176 147
rect 212 143 216 147
rect 252 143 256 147
rect 292 143 296 147
rect 332 143 336 147
rect 372 143 376 147
rect 408 143 412 147
rect 420 143 424 147
rect 468 143 472 147
rect 524 143 528 147
rect 580 143 584 147
rect 628 143 632 147
rect 664 143 668 147
rect 676 143 680 147
rect 724 143 728 147
rect 764 143 768 147
rect 804 143 808 147
rect 844 143 848 147
rect 884 143 888 147
rect 924 143 928 147
rect 960 143 964 147
rect 972 143 976 147
rect 1020 143 1024 147
rect 1068 143 1072 147
rect 1108 143 1112 147
rect 1148 143 1152 147
rect 1188 143 1192 147
rect 160 107 164 111
rect 200 107 204 111
rect 240 107 244 111
rect 280 107 284 111
rect 320 107 324 111
rect 360 107 364 111
rect 400 107 404 111
rect 408 107 412 111
rect 448 107 452 111
rect 496 107 500 111
rect 552 107 556 111
rect 608 107 612 111
rect 656 109 660 113
rect 664 111 668 115
rect 1328 115 1332 119
rect 1368 115 1372 119
rect 1408 115 1412 119
rect 1448 115 1452 119
rect 1488 115 1492 119
rect 1544 115 1548 119
rect 1552 115 1556 119
rect 1608 117 1612 121
rect 1616 119 1620 123
rect 1672 115 1676 119
rect 1736 117 1740 121
rect 1752 119 1756 123
rect 1792 115 1796 119
rect 1800 115 1804 119
rect 1848 115 1852 119
rect 1896 115 1900 119
rect 1944 115 1948 119
rect 1992 115 1996 119
rect 2040 115 2044 119
rect 2088 115 2092 119
rect 2136 115 2140 119
rect 2184 115 2188 119
rect 2240 115 2244 119
rect 2344 115 2348 119
rect 2384 115 2388 119
rect 704 107 708 111
rect 752 107 756 111
rect 792 107 796 111
rect 832 107 836 111
rect 872 107 876 111
rect 912 107 916 111
rect 952 107 956 111
rect 960 107 964 111
rect 1000 107 1004 111
rect 1048 107 1052 111
rect 1096 107 1100 111
rect 1136 107 1140 111
rect 1176 107 1180 111
rect 1216 107 1220 111
<< m2 >>
rect 1534 2508 1540 2509
rect 1534 2504 1535 2508
rect 1539 2504 1540 2508
rect 1534 2503 1540 2504
rect 1574 2508 1580 2509
rect 1574 2504 1575 2508
rect 1579 2504 1580 2508
rect 1574 2503 1580 2504
rect 1614 2508 1620 2509
rect 1614 2504 1615 2508
rect 1619 2504 1620 2508
rect 1614 2503 1620 2504
rect 1654 2508 1660 2509
rect 1654 2504 1655 2508
rect 1659 2504 1660 2508
rect 1654 2503 1660 2504
rect 1694 2508 1700 2509
rect 1694 2504 1695 2508
rect 1699 2504 1700 2508
rect 1694 2503 1700 2504
rect 1734 2508 1740 2509
rect 1734 2504 1735 2508
rect 1739 2504 1740 2508
rect 1734 2503 1740 2504
rect 1774 2508 1780 2509
rect 1774 2504 1775 2508
rect 1779 2504 1780 2508
rect 1774 2503 1780 2504
rect 1814 2508 1820 2509
rect 1814 2504 1815 2508
rect 1819 2504 1820 2508
rect 1814 2503 1820 2504
rect 1854 2508 1860 2509
rect 1854 2504 1855 2508
rect 1859 2504 1860 2508
rect 1854 2503 1860 2504
rect 1894 2508 1900 2509
rect 1894 2504 1895 2508
rect 1899 2504 1900 2508
rect 1894 2503 1900 2504
rect 1934 2508 1940 2509
rect 1934 2504 1935 2508
rect 1939 2504 1940 2508
rect 1934 2503 1940 2504
rect 1974 2508 1980 2509
rect 1974 2504 1975 2508
rect 1979 2504 1980 2508
rect 1974 2503 1980 2504
rect 1278 2501 1284 2502
rect 1278 2497 1279 2501
rect 1283 2497 1284 2501
rect 1278 2496 1284 2497
rect 2406 2501 2412 2502
rect 2406 2497 2407 2501
rect 2411 2497 2412 2501
rect 2406 2496 2412 2497
rect 158 2495 164 2496
rect 158 2491 159 2495
rect 163 2494 164 2495
rect 171 2495 177 2496
rect 171 2494 172 2495
rect 163 2492 172 2494
rect 163 2491 164 2492
rect 158 2490 164 2491
rect 171 2491 172 2492
rect 176 2491 177 2495
rect 171 2490 177 2491
rect 202 2495 208 2496
rect 202 2491 203 2495
rect 207 2494 208 2495
rect 211 2495 217 2496
rect 211 2494 212 2495
rect 207 2492 212 2494
rect 207 2491 208 2492
rect 202 2490 208 2491
rect 211 2491 212 2492
rect 216 2491 217 2495
rect 211 2490 217 2491
rect 242 2495 248 2496
rect 242 2491 243 2495
rect 247 2494 248 2495
rect 251 2495 257 2496
rect 251 2494 252 2495
rect 247 2492 252 2494
rect 247 2491 248 2492
rect 242 2490 248 2491
rect 251 2491 252 2492
rect 256 2491 257 2495
rect 251 2490 257 2491
rect 282 2495 288 2496
rect 282 2491 283 2495
rect 287 2494 288 2495
rect 307 2495 313 2496
rect 307 2494 308 2495
rect 287 2492 308 2494
rect 287 2491 288 2492
rect 282 2490 288 2491
rect 307 2491 308 2492
rect 312 2491 313 2495
rect 307 2490 313 2491
rect 338 2495 344 2496
rect 338 2491 339 2495
rect 343 2494 344 2495
rect 387 2495 393 2496
rect 387 2494 388 2495
rect 343 2492 388 2494
rect 343 2491 344 2492
rect 338 2490 344 2491
rect 387 2491 388 2492
rect 392 2491 393 2495
rect 387 2490 393 2491
rect 418 2495 424 2496
rect 418 2491 419 2495
rect 423 2494 424 2495
rect 475 2495 481 2496
rect 475 2494 476 2495
rect 423 2492 476 2494
rect 423 2491 424 2492
rect 418 2490 424 2491
rect 475 2491 476 2492
rect 480 2491 481 2495
rect 475 2490 481 2491
rect 506 2495 512 2496
rect 506 2491 507 2495
rect 511 2494 512 2495
rect 563 2495 569 2496
rect 563 2494 564 2495
rect 511 2492 564 2494
rect 511 2491 512 2492
rect 506 2490 512 2491
rect 563 2491 564 2492
rect 568 2491 569 2495
rect 563 2490 569 2491
rect 651 2495 657 2496
rect 651 2491 652 2495
rect 656 2494 657 2495
rect 670 2495 676 2496
rect 670 2494 671 2495
rect 656 2492 671 2494
rect 656 2491 657 2492
rect 651 2490 657 2491
rect 670 2491 671 2492
rect 675 2491 676 2495
rect 670 2490 676 2491
rect 682 2495 688 2496
rect 682 2491 683 2495
rect 687 2494 688 2495
rect 739 2495 745 2496
rect 739 2494 740 2495
rect 687 2492 740 2494
rect 687 2491 688 2492
rect 682 2490 688 2491
rect 739 2491 740 2492
rect 744 2491 745 2495
rect 739 2490 745 2491
rect 798 2495 804 2496
rect 798 2491 799 2495
rect 803 2494 804 2495
rect 827 2495 833 2496
rect 827 2494 828 2495
rect 803 2492 828 2494
rect 803 2491 804 2492
rect 798 2490 804 2491
rect 827 2491 828 2492
rect 832 2491 833 2495
rect 827 2490 833 2491
rect 858 2495 864 2496
rect 858 2491 859 2495
rect 863 2494 864 2495
rect 923 2495 929 2496
rect 923 2494 924 2495
rect 863 2492 924 2494
rect 863 2491 864 2492
rect 858 2490 864 2491
rect 923 2491 924 2492
rect 928 2491 929 2495
rect 923 2490 929 2491
rect 134 2487 140 2488
rect 134 2483 135 2487
rect 139 2483 140 2487
rect 134 2482 140 2483
rect 174 2487 180 2488
rect 174 2483 175 2487
rect 179 2483 180 2487
rect 174 2482 180 2483
rect 214 2487 220 2488
rect 214 2483 215 2487
rect 219 2483 220 2487
rect 214 2482 220 2483
rect 254 2487 260 2488
rect 254 2483 255 2487
rect 259 2483 260 2487
rect 254 2482 260 2483
rect 310 2487 316 2488
rect 310 2483 311 2487
rect 315 2483 316 2487
rect 310 2482 316 2483
rect 390 2487 396 2488
rect 390 2483 391 2487
rect 395 2483 396 2487
rect 390 2482 396 2483
rect 478 2487 484 2488
rect 478 2483 479 2487
rect 483 2483 484 2487
rect 478 2482 484 2483
rect 566 2487 572 2488
rect 566 2483 567 2487
rect 571 2483 572 2487
rect 566 2482 572 2483
rect 654 2487 660 2488
rect 654 2483 655 2487
rect 659 2483 660 2487
rect 654 2482 660 2483
rect 742 2487 748 2488
rect 742 2483 743 2487
rect 747 2483 748 2487
rect 742 2482 748 2483
rect 830 2487 836 2488
rect 830 2483 831 2487
rect 835 2483 836 2487
rect 830 2482 836 2483
rect 926 2487 932 2488
rect 926 2483 927 2487
rect 931 2483 932 2487
rect 1559 2487 1568 2488
rect 926 2482 932 2483
rect 1278 2484 1284 2485
rect 1278 2480 1279 2484
rect 1283 2480 1284 2484
rect 1559 2483 1560 2487
rect 1567 2483 1568 2487
rect 1559 2482 1568 2483
rect 1599 2487 1608 2488
rect 1599 2483 1600 2487
rect 1607 2483 1608 2487
rect 1599 2482 1608 2483
rect 1639 2487 1648 2488
rect 1639 2483 1640 2487
rect 1647 2483 1648 2487
rect 1639 2482 1648 2483
rect 1679 2487 1688 2488
rect 1679 2483 1680 2487
rect 1687 2483 1688 2487
rect 1679 2482 1688 2483
rect 1719 2487 1728 2488
rect 1719 2483 1720 2487
rect 1727 2483 1728 2487
rect 1719 2482 1728 2483
rect 1759 2487 1768 2488
rect 1759 2483 1760 2487
rect 1767 2483 1768 2487
rect 1759 2482 1768 2483
rect 1799 2487 1808 2488
rect 1799 2483 1800 2487
rect 1807 2483 1808 2487
rect 1799 2482 1808 2483
rect 1839 2487 1848 2488
rect 1839 2483 1840 2487
rect 1847 2483 1848 2487
rect 1839 2482 1848 2483
rect 1879 2487 1888 2488
rect 1879 2483 1880 2487
rect 1887 2483 1888 2487
rect 1879 2482 1888 2483
rect 1919 2487 1928 2488
rect 1919 2483 1920 2487
rect 1927 2483 1928 2487
rect 1919 2482 1928 2483
rect 1959 2487 1968 2488
rect 1959 2483 1960 2487
rect 1967 2483 1968 2487
rect 1959 2482 1968 2483
rect 1999 2487 2005 2488
rect 1999 2483 2000 2487
rect 2004 2483 2005 2487
rect 1999 2482 2005 2483
rect 2406 2484 2412 2485
rect 1278 2479 1284 2480
rect 1830 2479 1836 2480
rect 1830 2475 1831 2479
rect 1835 2478 1836 2479
rect 1999 2478 2001 2482
rect 2406 2480 2407 2484
rect 2411 2480 2412 2484
rect 2406 2479 2412 2480
rect 1835 2476 2001 2478
rect 1835 2475 1836 2476
rect 1830 2474 1836 2475
rect 110 2464 116 2465
rect 110 2460 111 2464
rect 115 2460 116 2464
rect 1238 2464 1244 2465
rect 1238 2460 1239 2464
rect 1243 2460 1244 2464
rect 110 2459 116 2460
rect 158 2459 165 2460
rect 158 2455 159 2459
rect 164 2455 165 2459
rect 158 2454 165 2455
rect 199 2459 208 2460
rect 199 2455 200 2459
rect 207 2455 208 2459
rect 199 2454 208 2455
rect 239 2459 248 2460
rect 239 2455 240 2459
rect 247 2455 248 2459
rect 239 2454 248 2455
rect 279 2459 288 2460
rect 279 2455 280 2459
rect 287 2455 288 2459
rect 279 2454 288 2455
rect 335 2459 344 2460
rect 335 2455 336 2459
rect 343 2455 344 2459
rect 335 2454 344 2455
rect 415 2459 424 2460
rect 415 2455 416 2459
rect 423 2455 424 2459
rect 415 2454 424 2455
rect 503 2459 512 2460
rect 503 2455 504 2459
rect 511 2455 512 2459
rect 591 2459 597 2460
rect 591 2458 592 2459
rect 503 2454 512 2455
rect 516 2456 592 2458
rect 142 2451 148 2452
rect 110 2447 116 2448
rect 110 2443 111 2447
rect 115 2443 116 2447
rect 142 2447 143 2451
rect 147 2450 148 2451
rect 516 2450 518 2456
rect 591 2455 592 2456
rect 596 2455 597 2459
rect 591 2454 597 2455
rect 679 2459 688 2460
rect 679 2455 680 2459
rect 687 2455 688 2459
rect 679 2454 688 2455
rect 767 2459 773 2460
rect 767 2455 768 2459
rect 772 2458 773 2459
rect 798 2459 804 2460
rect 798 2458 799 2459
rect 772 2456 799 2458
rect 772 2455 773 2456
rect 767 2454 773 2455
rect 798 2455 799 2456
rect 803 2455 804 2459
rect 798 2454 804 2455
rect 855 2459 864 2460
rect 855 2455 856 2459
rect 863 2455 864 2459
rect 855 2454 864 2455
rect 866 2459 872 2460
rect 866 2455 867 2459
rect 871 2458 872 2459
rect 951 2459 957 2460
rect 1238 2459 1244 2460
rect 1534 2461 1540 2462
rect 951 2458 952 2459
rect 871 2456 952 2458
rect 871 2455 872 2456
rect 866 2454 872 2455
rect 951 2455 952 2456
rect 956 2455 957 2459
rect 1534 2457 1535 2461
rect 1539 2457 1540 2461
rect 1534 2456 1540 2457
rect 1574 2461 1580 2462
rect 1574 2457 1575 2461
rect 1579 2457 1580 2461
rect 1574 2456 1580 2457
rect 1614 2461 1620 2462
rect 1614 2457 1615 2461
rect 1619 2457 1620 2461
rect 1614 2456 1620 2457
rect 1654 2461 1660 2462
rect 1654 2457 1655 2461
rect 1659 2457 1660 2461
rect 1654 2456 1660 2457
rect 1694 2461 1700 2462
rect 1694 2457 1695 2461
rect 1699 2457 1700 2461
rect 1694 2456 1700 2457
rect 1734 2461 1740 2462
rect 1734 2457 1735 2461
rect 1739 2457 1740 2461
rect 1734 2456 1740 2457
rect 1774 2461 1780 2462
rect 1774 2457 1775 2461
rect 1779 2457 1780 2461
rect 1774 2456 1780 2457
rect 1814 2461 1820 2462
rect 1814 2457 1815 2461
rect 1819 2457 1820 2461
rect 1814 2456 1820 2457
rect 1854 2461 1860 2462
rect 1854 2457 1855 2461
rect 1859 2457 1860 2461
rect 1854 2456 1860 2457
rect 1894 2461 1900 2462
rect 1894 2457 1895 2461
rect 1899 2457 1900 2461
rect 1894 2456 1900 2457
rect 1934 2461 1940 2462
rect 1934 2457 1935 2461
rect 1939 2457 1940 2461
rect 1934 2456 1940 2457
rect 1974 2461 1980 2462
rect 1974 2457 1975 2461
rect 1979 2457 1980 2461
rect 1974 2456 1980 2457
rect 951 2454 957 2455
rect 1602 2455 1608 2456
rect 147 2448 518 2450
rect 1531 2451 1537 2452
rect 147 2447 148 2448
rect 142 2446 148 2447
rect 1238 2447 1244 2448
rect 110 2442 116 2443
rect 1238 2443 1239 2447
rect 1243 2443 1244 2447
rect 1531 2447 1532 2451
rect 1536 2450 1537 2451
rect 1554 2451 1560 2452
rect 1554 2450 1555 2451
rect 1536 2448 1555 2450
rect 1536 2447 1537 2448
rect 1531 2446 1537 2447
rect 1554 2447 1555 2448
rect 1559 2447 1560 2451
rect 1554 2446 1560 2447
rect 1562 2451 1568 2452
rect 1562 2447 1563 2451
rect 1567 2450 1568 2451
rect 1571 2451 1577 2452
rect 1571 2450 1572 2451
rect 1567 2448 1572 2450
rect 1567 2447 1568 2448
rect 1562 2446 1568 2447
rect 1571 2447 1572 2448
rect 1576 2447 1577 2451
rect 1602 2451 1603 2455
rect 1607 2454 1608 2455
rect 1682 2455 1688 2456
rect 1607 2453 1617 2454
rect 1607 2452 1612 2453
rect 1607 2451 1608 2452
rect 1602 2450 1608 2451
rect 1611 2449 1612 2452
rect 1616 2449 1617 2453
rect 1611 2448 1617 2449
rect 1642 2451 1648 2452
rect 1571 2446 1577 2447
rect 1642 2447 1643 2451
rect 1647 2450 1648 2451
rect 1651 2451 1657 2452
rect 1651 2450 1652 2451
rect 1647 2448 1652 2450
rect 1647 2447 1648 2448
rect 1642 2446 1648 2447
rect 1651 2447 1652 2448
rect 1656 2447 1657 2451
rect 1682 2451 1683 2455
rect 1687 2454 1688 2455
rect 1762 2455 1768 2456
rect 1687 2453 1697 2454
rect 1687 2452 1692 2453
rect 1687 2451 1688 2452
rect 1682 2450 1688 2451
rect 1691 2449 1692 2452
rect 1696 2449 1697 2453
rect 1691 2448 1697 2449
rect 1722 2451 1728 2452
rect 1651 2446 1657 2447
rect 1722 2447 1723 2451
rect 1727 2450 1728 2451
rect 1731 2451 1737 2452
rect 1731 2450 1732 2451
rect 1727 2448 1732 2450
rect 1727 2447 1728 2448
rect 1722 2446 1728 2447
rect 1731 2447 1732 2448
rect 1736 2447 1737 2451
rect 1762 2451 1763 2455
rect 1767 2454 1768 2455
rect 1842 2455 1848 2456
rect 1767 2453 1777 2454
rect 1767 2452 1772 2453
rect 1767 2451 1768 2452
rect 1762 2450 1768 2451
rect 1771 2449 1772 2452
rect 1776 2449 1777 2453
rect 1771 2448 1777 2449
rect 1802 2451 1808 2452
rect 1731 2446 1737 2447
rect 1802 2447 1803 2451
rect 1807 2450 1808 2451
rect 1811 2451 1817 2452
rect 1811 2450 1812 2451
rect 1807 2448 1812 2450
rect 1807 2447 1808 2448
rect 1802 2446 1808 2447
rect 1811 2447 1812 2448
rect 1816 2447 1817 2451
rect 1842 2451 1843 2455
rect 1847 2454 1848 2455
rect 1922 2455 1928 2456
rect 1847 2453 1857 2454
rect 1847 2452 1852 2453
rect 1847 2451 1848 2452
rect 1842 2450 1848 2451
rect 1851 2449 1852 2452
rect 1856 2449 1857 2453
rect 1851 2448 1857 2449
rect 1882 2451 1888 2452
rect 1811 2446 1817 2447
rect 1882 2447 1883 2451
rect 1887 2450 1888 2451
rect 1891 2451 1897 2452
rect 1891 2450 1892 2451
rect 1887 2448 1892 2450
rect 1887 2447 1888 2448
rect 1882 2446 1888 2447
rect 1891 2447 1892 2448
rect 1896 2447 1897 2451
rect 1922 2451 1923 2455
rect 1927 2454 1928 2455
rect 1927 2453 1937 2454
rect 1927 2452 1932 2453
rect 1927 2451 1928 2452
rect 1922 2450 1928 2451
rect 1931 2449 1932 2452
rect 1936 2449 1937 2453
rect 1931 2448 1937 2449
rect 1962 2451 1968 2452
rect 1891 2446 1897 2447
rect 1962 2447 1963 2451
rect 1967 2450 1968 2451
rect 1971 2451 1977 2452
rect 1971 2450 1972 2451
rect 1967 2448 1972 2450
rect 1967 2447 1968 2448
rect 1962 2446 1968 2447
rect 1971 2447 1972 2448
rect 1976 2447 1977 2451
rect 1971 2446 1977 2447
rect 1238 2442 1244 2443
rect 134 2440 140 2441
rect 134 2436 135 2440
rect 139 2436 140 2440
rect 134 2435 140 2436
rect 174 2440 180 2441
rect 174 2436 175 2440
rect 179 2436 180 2440
rect 174 2435 180 2436
rect 214 2440 220 2441
rect 214 2436 215 2440
rect 219 2436 220 2440
rect 214 2435 220 2436
rect 254 2440 260 2441
rect 254 2436 255 2440
rect 259 2436 260 2440
rect 254 2435 260 2436
rect 310 2440 316 2441
rect 310 2436 311 2440
rect 315 2436 316 2440
rect 310 2435 316 2436
rect 390 2440 396 2441
rect 390 2436 391 2440
rect 395 2436 396 2440
rect 390 2435 396 2436
rect 478 2440 484 2441
rect 478 2436 479 2440
rect 483 2436 484 2440
rect 478 2435 484 2436
rect 566 2440 572 2441
rect 566 2436 567 2440
rect 571 2436 572 2440
rect 566 2435 572 2436
rect 654 2440 660 2441
rect 654 2436 655 2440
rect 659 2436 660 2440
rect 654 2435 660 2436
rect 742 2440 748 2441
rect 742 2436 743 2440
rect 747 2436 748 2440
rect 742 2435 748 2436
rect 830 2440 836 2441
rect 830 2436 831 2440
rect 835 2436 836 2440
rect 830 2435 836 2436
rect 926 2440 932 2441
rect 926 2436 927 2440
rect 931 2436 932 2440
rect 926 2435 932 2436
rect 1355 2439 1361 2440
rect 1355 2435 1356 2439
rect 1360 2438 1361 2439
rect 1378 2439 1384 2440
rect 1378 2438 1379 2439
rect 1360 2436 1379 2438
rect 1360 2435 1361 2436
rect 1355 2434 1361 2435
rect 1378 2435 1379 2436
rect 1383 2435 1384 2439
rect 1378 2434 1384 2435
rect 1386 2439 1392 2440
rect 1386 2435 1387 2439
rect 1391 2438 1392 2439
rect 1395 2439 1401 2440
rect 1395 2438 1396 2439
rect 1391 2436 1396 2438
rect 1391 2435 1392 2436
rect 1386 2434 1392 2435
rect 1395 2435 1396 2436
rect 1400 2435 1401 2439
rect 1395 2434 1401 2435
rect 1426 2439 1432 2440
rect 1426 2435 1427 2439
rect 1431 2438 1432 2439
rect 1451 2439 1457 2440
rect 1451 2438 1452 2439
rect 1431 2436 1452 2438
rect 1431 2435 1432 2436
rect 1426 2434 1432 2435
rect 1451 2435 1452 2436
rect 1456 2435 1457 2439
rect 1451 2434 1457 2435
rect 1482 2439 1488 2440
rect 1482 2435 1483 2439
rect 1487 2438 1488 2439
rect 1515 2439 1521 2440
rect 1515 2438 1516 2439
rect 1487 2436 1516 2438
rect 1487 2435 1488 2436
rect 1482 2434 1488 2435
rect 1515 2435 1516 2436
rect 1520 2435 1521 2439
rect 1515 2434 1521 2435
rect 1546 2439 1552 2440
rect 1546 2435 1547 2439
rect 1551 2438 1552 2439
rect 1595 2439 1601 2440
rect 1595 2438 1596 2439
rect 1551 2436 1596 2438
rect 1551 2435 1552 2436
rect 1546 2434 1552 2435
rect 1595 2435 1596 2436
rect 1600 2435 1601 2439
rect 1595 2434 1601 2435
rect 1626 2439 1632 2440
rect 1626 2435 1627 2439
rect 1631 2438 1632 2439
rect 1675 2439 1681 2440
rect 1675 2438 1676 2439
rect 1631 2436 1676 2438
rect 1631 2435 1632 2436
rect 1626 2434 1632 2435
rect 1675 2435 1676 2436
rect 1680 2435 1681 2439
rect 1675 2434 1681 2435
rect 1706 2439 1712 2440
rect 1706 2435 1707 2439
rect 1711 2438 1712 2439
rect 1755 2439 1761 2440
rect 1755 2438 1756 2439
rect 1711 2436 1756 2438
rect 1711 2435 1712 2436
rect 1706 2434 1712 2435
rect 1755 2435 1756 2436
rect 1760 2435 1761 2439
rect 1755 2434 1761 2435
rect 1830 2439 1841 2440
rect 1830 2435 1831 2439
rect 1835 2435 1836 2439
rect 1840 2435 1841 2439
rect 1830 2434 1841 2435
rect 1866 2439 1872 2440
rect 1866 2435 1867 2439
rect 1871 2438 1872 2439
rect 1915 2439 1921 2440
rect 1915 2438 1916 2439
rect 1871 2436 1916 2438
rect 1871 2435 1872 2436
rect 1866 2434 1872 2435
rect 1915 2435 1916 2436
rect 1920 2435 1921 2439
rect 1915 2434 1921 2435
rect 1946 2439 1952 2440
rect 1946 2435 1947 2439
rect 1951 2438 1952 2439
rect 1995 2439 2001 2440
rect 1995 2438 1996 2439
rect 1951 2436 1996 2438
rect 1951 2435 1952 2436
rect 1946 2434 1952 2435
rect 1995 2435 1996 2436
rect 2000 2435 2001 2439
rect 1995 2434 2001 2435
rect 2026 2439 2032 2440
rect 2026 2435 2027 2439
rect 2031 2438 2032 2439
rect 2075 2439 2081 2440
rect 2075 2438 2076 2439
rect 2031 2436 2076 2438
rect 2031 2435 2032 2436
rect 2026 2434 2032 2435
rect 2075 2435 2076 2436
rect 2080 2435 2081 2439
rect 2075 2434 2081 2435
rect 2106 2439 2112 2440
rect 2106 2435 2107 2439
rect 2111 2438 2112 2439
rect 2155 2439 2161 2440
rect 2155 2438 2156 2439
rect 2111 2436 2156 2438
rect 2111 2435 2112 2436
rect 2106 2434 2112 2435
rect 2155 2435 2156 2436
rect 2160 2435 2161 2439
rect 2155 2434 2161 2435
rect 2182 2439 2188 2440
rect 2182 2435 2183 2439
rect 2187 2438 2188 2439
rect 2243 2439 2249 2440
rect 2243 2438 2244 2439
rect 2187 2436 2244 2438
rect 2187 2435 2188 2436
rect 2182 2434 2188 2435
rect 2243 2435 2244 2436
rect 2248 2435 2249 2439
rect 2243 2434 2249 2435
rect 2290 2439 2296 2440
rect 2290 2435 2291 2439
rect 2295 2438 2296 2439
rect 2331 2439 2337 2440
rect 2331 2438 2332 2439
rect 2295 2436 2332 2438
rect 2295 2435 2296 2436
rect 2290 2434 2296 2435
rect 2331 2435 2332 2436
rect 2336 2435 2337 2439
rect 2331 2434 2337 2435
rect 1358 2431 1364 2432
rect 134 2428 140 2429
rect 134 2424 135 2428
rect 139 2424 140 2428
rect 134 2423 140 2424
rect 182 2428 188 2429
rect 182 2424 183 2428
rect 187 2424 188 2428
rect 182 2423 188 2424
rect 246 2428 252 2429
rect 246 2424 247 2428
rect 251 2424 252 2428
rect 246 2423 252 2424
rect 318 2428 324 2429
rect 318 2424 319 2428
rect 323 2424 324 2428
rect 318 2423 324 2424
rect 390 2428 396 2429
rect 390 2424 391 2428
rect 395 2424 396 2428
rect 390 2423 396 2424
rect 470 2428 476 2429
rect 470 2424 471 2428
rect 475 2424 476 2428
rect 470 2423 476 2424
rect 542 2428 548 2429
rect 542 2424 543 2428
rect 547 2424 548 2428
rect 542 2423 548 2424
rect 614 2428 620 2429
rect 614 2424 615 2428
rect 619 2424 620 2428
rect 614 2423 620 2424
rect 678 2428 684 2429
rect 678 2424 679 2428
rect 683 2424 684 2428
rect 678 2423 684 2424
rect 734 2428 740 2429
rect 734 2424 735 2428
rect 739 2424 740 2428
rect 734 2423 740 2424
rect 790 2428 796 2429
rect 790 2424 791 2428
rect 795 2424 796 2428
rect 790 2423 796 2424
rect 838 2428 844 2429
rect 838 2424 839 2428
rect 843 2424 844 2428
rect 838 2423 844 2424
rect 886 2428 892 2429
rect 886 2424 887 2428
rect 891 2424 892 2428
rect 886 2423 892 2424
rect 934 2428 940 2429
rect 934 2424 935 2428
rect 939 2424 940 2428
rect 934 2423 940 2424
rect 990 2428 996 2429
rect 990 2424 991 2428
rect 995 2424 996 2428
rect 990 2423 996 2424
rect 1046 2428 1052 2429
rect 1046 2424 1047 2428
rect 1051 2424 1052 2428
rect 1358 2427 1359 2431
rect 1363 2427 1364 2431
rect 1358 2426 1364 2427
rect 1398 2431 1404 2432
rect 1398 2427 1399 2431
rect 1403 2427 1404 2431
rect 1398 2426 1404 2427
rect 1454 2431 1460 2432
rect 1454 2427 1455 2431
rect 1459 2427 1460 2431
rect 1454 2426 1460 2427
rect 1518 2431 1524 2432
rect 1518 2427 1519 2431
rect 1523 2427 1524 2431
rect 1518 2426 1524 2427
rect 1598 2431 1604 2432
rect 1598 2427 1599 2431
rect 1603 2427 1604 2431
rect 1598 2426 1604 2427
rect 1678 2431 1684 2432
rect 1678 2427 1679 2431
rect 1683 2427 1684 2431
rect 1678 2426 1684 2427
rect 1758 2431 1764 2432
rect 1758 2427 1759 2431
rect 1763 2427 1764 2431
rect 1758 2426 1764 2427
rect 1838 2431 1844 2432
rect 1838 2427 1839 2431
rect 1843 2427 1844 2431
rect 1838 2426 1844 2427
rect 1918 2431 1924 2432
rect 1918 2427 1919 2431
rect 1923 2427 1924 2431
rect 1918 2426 1924 2427
rect 1998 2431 2004 2432
rect 1998 2427 1999 2431
rect 2003 2427 2004 2431
rect 1998 2426 2004 2427
rect 2078 2431 2084 2432
rect 2078 2427 2079 2431
rect 2083 2427 2084 2431
rect 2078 2426 2084 2427
rect 2158 2431 2164 2432
rect 2158 2427 2159 2431
rect 2163 2427 2164 2431
rect 2158 2426 2164 2427
rect 2246 2431 2252 2432
rect 2246 2427 2247 2431
rect 2251 2427 2252 2431
rect 2246 2426 2252 2427
rect 2334 2431 2340 2432
rect 2334 2427 2335 2431
rect 2339 2427 2340 2431
rect 2334 2426 2340 2427
rect 1046 2423 1052 2424
rect 110 2421 116 2422
rect 110 2417 111 2421
rect 115 2417 116 2421
rect 110 2416 116 2417
rect 1238 2421 1244 2422
rect 1238 2417 1239 2421
rect 1243 2417 1244 2421
rect 1238 2416 1244 2417
rect 670 2415 676 2416
rect 670 2411 671 2415
rect 675 2414 676 2415
rect 675 2412 794 2414
rect 675 2411 676 2412
rect 670 2410 676 2411
rect 159 2407 165 2408
rect 110 2404 116 2405
rect 110 2400 111 2404
rect 115 2400 116 2404
rect 159 2403 160 2407
rect 164 2406 165 2407
rect 174 2407 180 2408
rect 174 2406 175 2407
rect 164 2404 175 2406
rect 164 2403 165 2404
rect 159 2402 165 2403
rect 174 2403 175 2404
rect 179 2403 180 2407
rect 174 2402 180 2403
rect 207 2407 213 2408
rect 207 2403 208 2407
rect 212 2406 213 2407
rect 238 2407 244 2408
rect 238 2406 239 2407
rect 212 2404 239 2406
rect 212 2403 213 2404
rect 207 2402 213 2403
rect 238 2403 239 2404
rect 243 2403 244 2407
rect 238 2402 244 2403
rect 271 2407 277 2408
rect 271 2403 272 2407
rect 276 2406 277 2407
rect 310 2407 316 2408
rect 310 2406 311 2407
rect 276 2404 311 2406
rect 276 2403 277 2404
rect 271 2402 277 2403
rect 310 2403 311 2404
rect 315 2403 316 2407
rect 310 2402 316 2403
rect 343 2407 349 2408
rect 343 2403 344 2407
rect 348 2406 349 2407
rect 382 2407 388 2408
rect 382 2406 383 2407
rect 348 2404 383 2406
rect 348 2403 349 2404
rect 343 2402 349 2403
rect 382 2403 383 2404
rect 387 2403 388 2407
rect 382 2402 388 2403
rect 415 2407 421 2408
rect 415 2403 416 2407
rect 420 2406 421 2407
rect 462 2407 468 2408
rect 462 2406 463 2407
rect 420 2404 463 2406
rect 420 2403 421 2404
rect 415 2402 421 2403
rect 462 2403 463 2404
rect 467 2403 468 2407
rect 462 2402 468 2403
rect 495 2407 501 2408
rect 495 2403 496 2407
rect 500 2406 501 2407
rect 510 2407 516 2408
rect 510 2406 511 2407
rect 500 2404 511 2406
rect 500 2403 501 2404
rect 495 2402 501 2403
rect 510 2403 511 2404
rect 515 2403 516 2407
rect 510 2402 516 2403
rect 567 2407 573 2408
rect 567 2403 568 2407
rect 572 2406 573 2407
rect 606 2407 612 2408
rect 606 2406 607 2407
rect 572 2404 607 2406
rect 572 2403 573 2404
rect 567 2402 573 2403
rect 606 2403 607 2404
rect 611 2403 612 2407
rect 606 2402 612 2403
rect 639 2407 645 2408
rect 639 2403 640 2407
rect 644 2406 645 2407
rect 670 2407 676 2408
rect 670 2406 671 2407
rect 644 2404 671 2406
rect 644 2403 645 2404
rect 639 2402 645 2403
rect 670 2403 671 2404
rect 675 2403 676 2407
rect 670 2402 676 2403
rect 703 2407 709 2408
rect 703 2403 704 2407
rect 708 2406 709 2407
rect 726 2407 732 2408
rect 726 2406 727 2407
rect 708 2404 727 2406
rect 708 2403 709 2404
rect 703 2402 709 2403
rect 726 2403 727 2404
rect 731 2403 732 2407
rect 726 2402 732 2403
rect 759 2407 765 2408
rect 759 2403 760 2407
rect 764 2406 765 2407
rect 782 2407 788 2408
rect 782 2406 783 2407
rect 764 2404 783 2406
rect 764 2403 765 2404
rect 759 2402 765 2403
rect 782 2403 783 2404
rect 787 2403 788 2407
rect 792 2406 794 2412
rect 1554 2411 1560 2412
rect 1278 2408 1284 2409
rect 815 2407 821 2408
rect 815 2406 816 2407
rect 792 2404 816 2406
rect 782 2402 788 2403
rect 815 2403 816 2404
rect 820 2403 821 2407
rect 815 2402 821 2403
rect 863 2407 869 2408
rect 863 2403 864 2407
rect 868 2406 869 2407
rect 878 2407 884 2408
rect 878 2406 879 2407
rect 868 2404 879 2406
rect 868 2403 869 2404
rect 863 2402 869 2403
rect 878 2403 879 2404
rect 883 2403 884 2407
rect 878 2402 884 2403
rect 911 2407 917 2408
rect 911 2403 912 2407
rect 916 2406 917 2407
rect 926 2407 932 2408
rect 926 2406 927 2407
rect 916 2404 927 2406
rect 916 2403 917 2404
rect 911 2402 917 2403
rect 926 2403 927 2404
rect 931 2403 932 2407
rect 926 2402 932 2403
rect 959 2407 965 2408
rect 959 2403 960 2407
rect 964 2406 965 2407
rect 974 2407 980 2408
rect 974 2406 975 2407
rect 964 2404 975 2406
rect 964 2403 965 2404
rect 959 2402 965 2403
rect 974 2403 975 2404
rect 979 2403 980 2407
rect 974 2402 980 2403
rect 1015 2407 1021 2408
rect 1015 2403 1016 2407
rect 1020 2406 1021 2407
rect 1038 2407 1044 2408
rect 1038 2406 1039 2407
rect 1020 2404 1039 2406
rect 1020 2403 1021 2404
rect 1015 2402 1021 2403
rect 1038 2403 1039 2404
rect 1043 2403 1044 2407
rect 1038 2402 1044 2403
rect 1054 2407 1060 2408
rect 1054 2403 1055 2407
rect 1059 2406 1060 2407
rect 1071 2407 1077 2408
rect 1071 2406 1072 2407
rect 1059 2404 1072 2406
rect 1059 2403 1060 2404
rect 1054 2402 1060 2403
rect 1071 2403 1072 2404
rect 1076 2403 1077 2407
rect 1071 2402 1077 2403
rect 1238 2404 1244 2405
rect 110 2399 116 2400
rect 1238 2400 1239 2404
rect 1243 2400 1244 2404
rect 1278 2404 1279 2408
rect 1283 2404 1284 2408
rect 1554 2407 1555 2411
rect 1559 2410 1560 2411
rect 1559 2408 1718 2410
rect 1559 2407 1560 2408
rect 1554 2406 1560 2407
rect 1278 2403 1284 2404
rect 1383 2403 1392 2404
rect 1238 2399 1244 2400
rect 1383 2399 1384 2403
rect 1391 2399 1392 2403
rect 1383 2398 1392 2399
rect 1423 2403 1432 2404
rect 1423 2399 1424 2403
rect 1431 2399 1432 2403
rect 1423 2398 1432 2399
rect 1479 2403 1488 2404
rect 1479 2399 1480 2403
rect 1487 2399 1488 2403
rect 1479 2398 1488 2399
rect 1543 2403 1552 2404
rect 1543 2399 1544 2403
rect 1551 2399 1552 2403
rect 1543 2398 1552 2399
rect 1623 2403 1632 2404
rect 1623 2399 1624 2403
rect 1631 2399 1632 2403
rect 1623 2398 1632 2399
rect 1703 2403 1712 2404
rect 1703 2399 1704 2403
rect 1711 2399 1712 2403
rect 1716 2402 1718 2408
rect 2406 2408 2412 2409
rect 2406 2404 2407 2408
rect 2411 2404 2412 2408
rect 1783 2403 1789 2404
rect 1783 2402 1784 2403
rect 1716 2400 1784 2402
rect 1703 2398 1712 2399
rect 1783 2399 1784 2400
rect 1788 2399 1789 2403
rect 1783 2398 1789 2399
rect 1863 2403 1872 2404
rect 1863 2399 1864 2403
rect 1871 2399 1872 2403
rect 1863 2398 1872 2399
rect 1943 2403 1952 2404
rect 1943 2399 1944 2403
rect 1951 2399 1952 2403
rect 1943 2398 1952 2399
rect 2023 2403 2032 2404
rect 2023 2399 2024 2403
rect 2031 2399 2032 2403
rect 2023 2398 2032 2399
rect 2103 2403 2112 2404
rect 2103 2399 2104 2403
rect 2111 2399 2112 2403
rect 2103 2398 2112 2399
rect 2182 2403 2189 2404
rect 2182 2399 2183 2403
rect 2188 2399 2189 2403
rect 2182 2398 2189 2399
rect 2191 2403 2197 2404
rect 2191 2399 2192 2403
rect 2196 2402 2197 2403
rect 2271 2403 2277 2404
rect 2271 2402 2272 2403
rect 2196 2400 2272 2402
rect 2196 2399 2197 2400
rect 2191 2398 2197 2399
rect 2271 2399 2272 2400
rect 2276 2399 2277 2403
rect 2271 2398 2277 2399
rect 2350 2403 2356 2404
rect 2350 2399 2351 2403
rect 2355 2402 2356 2403
rect 2359 2403 2365 2404
rect 2406 2403 2412 2404
rect 2359 2402 2360 2403
rect 2355 2400 2360 2402
rect 2355 2399 2356 2400
rect 2350 2398 2356 2399
rect 2359 2399 2360 2400
rect 2364 2399 2365 2403
rect 2359 2398 2365 2399
rect 1278 2391 1284 2392
rect 1278 2387 1279 2391
rect 1283 2387 1284 2391
rect 1278 2386 1284 2387
rect 2406 2391 2412 2392
rect 2406 2387 2407 2391
rect 2411 2387 2412 2391
rect 2406 2386 2412 2387
rect 1358 2384 1364 2385
rect 134 2381 140 2382
rect 134 2377 135 2381
rect 139 2377 140 2381
rect 134 2376 140 2377
rect 182 2381 188 2382
rect 182 2377 183 2381
rect 187 2377 188 2381
rect 182 2376 188 2377
rect 246 2381 252 2382
rect 246 2377 247 2381
rect 251 2377 252 2381
rect 246 2376 252 2377
rect 318 2381 324 2382
rect 318 2377 319 2381
rect 323 2377 324 2381
rect 318 2376 324 2377
rect 390 2381 396 2382
rect 390 2377 391 2381
rect 395 2377 396 2381
rect 390 2376 396 2377
rect 470 2381 476 2382
rect 470 2377 471 2381
rect 475 2377 476 2381
rect 470 2376 476 2377
rect 542 2381 548 2382
rect 542 2377 543 2381
rect 547 2377 548 2381
rect 542 2376 548 2377
rect 614 2381 620 2382
rect 614 2377 615 2381
rect 619 2377 620 2381
rect 614 2376 620 2377
rect 678 2381 684 2382
rect 678 2377 679 2381
rect 683 2377 684 2381
rect 678 2376 684 2377
rect 734 2381 740 2382
rect 734 2377 735 2381
rect 739 2377 740 2381
rect 734 2376 740 2377
rect 790 2381 796 2382
rect 790 2377 791 2381
rect 795 2377 796 2381
rect 790 2376 796 2377
rect 838 2381 844 2382
rect 838 2377 839 2381
rect 843 2377 844 2381
rect 838 2376 844 2377
rect 886 2381 892 2382
rect 886 2377 887 2381
rect 891 2377 892 2381
rect 886 2376 892 2377
rect 934 2381 940 2382
rect 934 2377 935 2381
rect 939 2377 940 2381
rect 934 2376 940 2377
rect 990 2381 996 2382
rect 990 2377 991 2381
rect 995 2377 996 2381
rect 990 2376 996 2377
rect 1046 2381 1052 2382
rect 1046 2377 1047 2381
rect 1051 2377 1052 2381
rect 1358 2380 1359 2384
rect 1363 2380 1364 2384
rect 1358 2379 1364 2380
rect 1398 2384 1404 2385
rect 1398 2380 1399 2384
rect 1403 2380 1404 2384
rect 1398 2379 1404 2380
rect 1454 2384 1460 2385
rect 1454 2380 1455 2384
rect 1459 2380 1460 2384
rect 1454 2379 1460 2380
rect 1518 2384 1524 2385
rect 1518 2380 1519 2384
rect 1523 2380 1524 2384
rect 1518 2379 1524 2380
rect 1598 2384 1604 2385
rect 1598 2380 1599 2384
rect 1603 2380 1604 2384
rect 1598 2379 1604 2380
rect 1678 2384 1684 2385
rect 1678 2380 1679 2384
rect 1683 2380 1684 2384
rect 1678 2379 1684 2380
rect 1758 2384 1764 2385
rect 1758 2380 1759 2384
rect 1763 2380 1764 2384
rect 1758 2379 1764 2380
rect 1838 2384 1844 2385
rect 1838 2380 1839 2384
rect 1843 2380 1844 2384
rect 1838 2379 1844 2380
rect 1918 2384 1924 2385
rect 1918 2380 1919 2384
rect 1923 2380 1924 2384
rect 1918 2379 1924 2380
rect 1998 2384 2004 2385
rect 1998 2380 1999 2384
rect 2003 2380 2004 2384
rect 1998 2379 2004 2380
rect 2078 2384 2084 2385
rect 2078 2380 2079 2384
rect 2083 2380 2084 2384
rect 2078 2379 2084 2380
rect 2158 2384 2164 2385
rect 2158 2380 2159 2384
rect 2163 2380 2164 2384
rect 2158 2379 2164 2380
rect 2246 2384 2252 2385
rect 2246 2380 2247 2384
rect 2251 2380 2252 2384
rect 2246 2379 2252 2380
rect 2334 2384 2340 2385
rect 2334 2380 2335 2384
rect 2339 2380 2340 2384
rect 2334 2379 2340 2380
rect 1046 2376 1052 2377
rect 1358 2372 1364 2373
rect 131 2371 137 2372
rect 131 2367 132 2371
rect 136 2370 137 2371
rect 142 2371 148 2372
rect 142 2370 143 2371
rect 136 2368 143 2370
rect 136 2367 137 2368
rect 131 2366 137 2367
rect 142 2367 143 2368
rect 147 2367 148 2371
rect 142 2366 148 2367
rect 174 2371 185 2372
rect 174 2367 175 2371
rect 179 2367 180 2371
rect 184 2367 185 2371
rect 174 2366 185 2367
rect 238 2371 249 2372
rect 238 2367 239 2371
rect 243 2367 244 2371
rect 248 2367 249 2371
rect 238 2366 249 2367
rect 310 2371 321 2372
rect 310 2367 311 2371
rect 315 2367 316 2371
rect 320 2367 321 2371
rect 310 2366 321 2367
rect 382 2371 393 2372
rect 382 2367 383 2371
rect 387 2367 388 2371
rect 392 2367 393 2371
rect 382 2366 393 2367
rect 462 2371 473 2372
rect 462 2367 463 2371
rect 467 2367 468 2371
rect 472 2367 473 2371
rect 462 2366 473 2367
rect 539 2371 545 2372
rect 539 2367 540 2371
rect 544 2370 545 2371
rect 590 2371 596 2372
rect 590 2370 591 2371
rect 544 2368 591 2370
rect 544 2367 545 2368
rect 539 2366 545 2367
rect 590 2367 591 2368
rect 595 2367 596 2371
rect 590 2366 596 2367
rect 606 2371 617 2372
rect 606 2367 607 2371
rect 611 2367 612 2371
rect 616 2367 617 2371
rect 606 2366 617 2367
rect 670 2371 681 2372
rect 670 2367 671 2371
rect 675 2367 676 2371
rect 680 2367 681 2371
rect 670 2366 681 2367
rect 726 2371 737 2372
rect 726 2367 727 2371
rect 731 2367 732 2371
rect 736 2367 737 2371
rect 726 2366 737 2367
rect 782 2371 793 2372
rect 782 2367 783 2371
rect 787 2367 788 2371
rect 792 2367 793 2371
rect 782 2366 793 2367
rect 835 2371 841 2372
rect 835 2367 836 2371
rect 840 2370 841 2371
rect 866 2371 872 2372
rect 866 2370 867 2371
rect 840 2368 867 2370
rect 840 2367 841 2368
rect 835 2366 841 2367
rect 866 2367 867 2368
rect 871 2367 872 2371
rect 866 2366 872 2367
rect 878 2371 889 2372
rect 878 2367 879 2371
rect 883 2367 884 2371
rect 888 2367 889 2371
rect 878 2366 889 2367
rect 926 2371 937 2372
rect 926 2367 927 2371
rect 931 2367 932 2371
rect 936 2367 937 2371
rect 926 2366 937 2367
rect 974 2371 980 2372
rect 974 2367 975 2371
rect 979 2370 980 2371
rect 987 2371 993 2372
rect 987 2370 988 2371
rect 979 2368 988 2370
rect 979 2367 980 2368
rect 974 2366 980 2367
rect 987 2367 988 2368
rect 992 2367 993 2371
rect 987 2366 993 2367
rect 1038 2371 1049 2372
rect 1038 2367 1039 2371
rect 1043 2367 1044 2371
rect 1048 2367 1049 2371
rect 1358 2368 1359 2372
rect 1363 2368 1364 2372
rect 1358 2367 1364 2368
rect 1406 2372 1412 2373
rect 1406 2368 1407 2372
rect 1411 2368 1412 2372
rect 1406 2367 1412 2368
rect 1470 2372 1476 2373
rect 1470 2368 1471 2372
rect 1475 2368 1476 2372
rect 1470 2367 1476 2368
rect 1542 2372 1548 2373
rect 1542 2368 1543 2372
rect 1547 2368 1548 2372
rect 1542 2367 1548 2368
rect 1614 2372 1620 2373
rect 1614 2368 1615 2372
rect 1619 2368 1620 2372
rect 1614 2367 1620 2368
rect 1694 2372 1700 2373
rect 1694 2368 1695 2372
rect 1699 2368 1700 2372
rect 1694 2367 1700 2368
rect 1774 2372 1780 2373
rect 1774 2368 1775 2372
rect 1779 2368 1780 2372
rect 1774 2367 1780 2368
rect 1854 2372 1860 2373
rect 1854 2368 1855 2372
rect 1859 2368 1860 2372
rect 1854 2367 1860 2368
rect 1926 2372 1932 2373
rect 1926 2368 1927 2372
rect 1931 2368 1932 2372
rect 1926 2367 1932 2368
rect 1998 2372 2004 2373
rect 1998 2368 1999 2372
rect 2003 2368 2004 2372
rect 1998 2367 2004 2368
rect 2070 2372 2076 2373
rect 2070 2368 2071 2372
rect 2075 2368 2076 2372
rect 2070 2367 2076 2368
rect 2142 2372 2148 2373
rect 2142 2368 2143 2372
rect 2147 2368 2148 2372
rect 2142 2367 2148 2368
rect 2222 2372 2228 2373
rect 2222 2368 2223 2372
rect 2227 2368 2228 2372
rect 2222 2367 2228 2368
rect 2302 2372 2308 2373
rect 2302 2368 2303 2372
rect 2307 2368 2308 2372
rect 2302 2367 2308 2368
rect 2358 2372 2364 2373
rect 2358 2368 2359 2372
rect 2363 2368 2364 2372
rect 2358 2367 2364 2368
rect 1038 2366 1049 2367
rect 1278 2365 1284 2366
rect 1278 2361 1279 2365
rect 1283 2361 1284 2365
rect 1278 2360 1284 2361
rect 2406 2365 2412 2366
rect 2406 2361 2407 2365
rect 2411 2361 2412 2365
rect 2406 2360 2412 2361
rect 1054 2359 1060 2360
rect 1054 2358 1055 2359
rect 820 2356 1055 2358
rect 820 2354 822 2356
rect 1054 2355 1055 2356
rect 1059 2355 1060 2359
rect 1054 2354 1060 2355
rect 2290 2355 2296 2356
rect 2290 2354 2291 2355
rect 819 2353 825 2354
rect 131 2351 137 2352
rect 131 2347 132 2351
rect 136 2350 137 2351
rect 154 2351 160 2352
rect 154 2350 155 2351
rect 136 2348 155 2350
rect 136 2347 137 2348
rect 131 2346 137 2347
rect 154 2347 155 2348
rect 159 2347 160 2351
rect 154 2346 160 2347
rect 162 2351 168 2352
rect 162 2347 163 2351
rect 167 2350 168 2351
rect 171 2351 177 2352
rect 171 2350 172 2351
rect 167 2348 172 2350
rect 167 2347 168 2348
rect 162 2346 168 2347
rect 171 2347 172 2348
rect 176 2347 177 2351
rect 171 2346 177 2347
rect 202 2351 208 2352
rect 202 2347 203 2351
rect 207 2350 208 2351
rect 211 2351 217 2352
rect 211 2350 212 2351
rect 207 2348 212 2350
rect 207 2347 208 2348
rect 202 2346 208 2347
rect 211 2347 212 2348
rect 216 2347 217 2351
rect 211 2346 217 2347
rect 247 2351 253 2352
rect 247 2347 248 2351
rect 252 2350 253 2351
rect 267 2351 273 2352
rect 267 2350 268 2351
rect 252 2348 268 2350
rect 252 2347 253 2348
rect 247 2346 253 2347
rect 267 2347 268 2348
rect 272 2347 273 2351
rect 267 2346 273 2347
rect 347 2351 353 2352
rect 347 2347 348 2351
rect 352 2350 353 2351
rect 418 2351 424 2352
rect 418 2350 419 2351
rect 352 2348 419 2350
rect 352 2347 353 2348
rect 347 2346 353 2347
rect 418 2347 419 2348
rect 423 2347 424 2351
rect 418 2346 424 2347
rect 427 2351 433 2352
rect 427 2347 428 2351
rect 432 2350 433 2351
rect 502 2351 508 2352
rect 502 2350 503 2351
rect 432 2348 503 2350
rect 432 2347 433 2348
rect 427 2346 433 2347
rect 502 2347 503 2348
rect 507 2347 508 2351
rect 502 2346 508 2347
rect 510 2351 521 2352
rect 510 2347 511 2351
rect 515 2347 516 2351
rect 520 2347 521 2351
rect 510 2346 521 2347
rect 595 2351 601 2352
rect 595 2347 596 2351
rect 600 2350 601 2351
rect 666 2351 672 2352
rect 666 2350 667 2351
rect 600 2348 667 2350
rect 600 2347 601 2348
rect 595 2346 601 2347
rect 666 2347 667 2348
rect 671 2347 672 2351
rect 666 2346 672 2347
rect 675 2351 681 2352
rect 675 2347 676 2351
rect 680 2350 681 2351
rect 726 2351 732 2352
rect 726 2350 727 2351
rect 680 2348 727 2350
rect 680 2347 681 2348
rect 675 2346 681 2347
rect 726 2347 727 2348
rect 731 2347 732 2351
rect 726 2346 732 2347
rect 747 2351 753 2352
rect 747 2347 748 2351
rect 752 2350 753 2351
rect 782 2351 788 2352
rect 782 2350 783 2351
rect 752 2348 783 2350
rect 752 2347 753 2348
rect 747 2346 753 2347
rect 782 2347 783 2348
rect 787 2347 788 2351
rect 819 2349 820 2353
rect 824 2349 825 2353
rect 2247 2353 2291 2354
rect 819 2348 825 2349
rect 850 2351 856 2352
rect 782 2346 788 2347
rect 850 2347 851 2351
rect 855 2350 856 2351
rect 883 2351 889 2352
rect 883 2350 884 2351
rect 855 2348 884 2350
rect 855 2347 856 2348
rect 850 2346 856 2347
rect 883 2347 884 2348
rect 888 2347 889 2351
rect 883 2346 889 2347
rect 914 2351 920 2352
rect 914 2347 915 2351
rect 919 2350 920 2351
rect 955 2351 961 2352
rect 955 2350 956 2351
rect 919 2348 956 2350
rect 919 2347 920 2348
rect 914 2346 920 2347
rect 955 2347 956 2348
rect 960 2347 961 2351
rect 955 2346 961 2347
rect 991 2351 997 2352
rect 991 2347 992 2351
rect 996 2350 997 2351
rect 1027 2351 1033 2352
rect 1027 2350 1028 2351
rect 996 2348 1028 2350
rect 996 2347 997 2348
rect 991 2346 997 2347
rect 1027 2347 1028 2348
rect 1032 2347 1033 2351
rect 1378 2351 1389 2352
rect 1027 2346 1033 2347
rect 1278 2348 1284 2349
rect 1278 2344 1279 2348
rect 1283 2344 1284 2348
rect 1378 2347 1379 2351
rect 1383 2347 1384 2351
rect 1388 2347 1389 2351
rect 1378 2346 1389 2347
rect 1391 2351 1397 2352
rect 1391 2347 1392 2351
rect 1396 2350 1397 2351
rect 1431 2351 1437 2352
rect 1431 2350 1432 2351
rect 1396 2348 1432 2350
rect 1396 2347 1397 2348
rect 1391 2346 1397 2347
rect 1431 2347 1432 2348
rect 1436 2347 1437 2351
rect 1431 2346 1437 2347
rect 1439 2351 1445 2352
rect 1439 2347 1440 2351
rect 1444 2350 1445 2351
rect 1495 2351 1501 2352
rect 1495 2350 1496 2351
rect 1444 2348 1496 2350
rect 1444 2347 1445 2348
rect 1439 2346 1445 2347
rect 1495 2347 1496 2348
rect 1500 2347 1501 2351
rect 1495 2346 1501 2347
rect 1503 2351 1509 2352
rect 1503 2347 1504 2351
rect 1508 2350 1509 2351
rect 1567 2351 1573 2352
rect 1567 2350 1568 2351
rect 1508 2348 1568 2350
rect 1508 2347 1509 2348
rect 1503 2346 1509 2347
rect 1567 2347 1568 2348
rect 1572 2347 1573 2351
rect 1567 2346 1573 2347
rect 1639 2351 1645 2352
rect 1639 2347 1640 2351
rect 1644 2350 1645 2351
rect 1686 2351 1692 2352
rect 1686 2350 1687 2351
rect 1644 2348 1687 2350
rect 1644 2347 1645 2348
rect 1639 2346 1645 2347
rect 1686 2347 1687 2348
rect 1691 2347 1692 2351
rect 1719 2351 1725 2352
rect 1719 2350 1720 2351
rect 1686 2346 1692 2347
rect 1696 2348 1720 2350
rect 134 2343 140 2344
rect 134 2339 135 2343
rect 139 2339 140 2343
rect 134 2338 140 2339
rect 174 2343 180 2344
rect 174 2339 175 2343
rect 179 2339 180 2343
rect 174 2338 180 2339
rect 214 2343 220 2344
rect 214 2339 215 2343
rect 219 2339 220 2343
rect 214 2338 220 2339
rect 270 2343 276 2344
rect 270 2339 271 2343
rect 275 2339 276 2343
rect 270 2338 276 2339
rect 350 2343 356 2344
rect 350 2339 351 2343
rect 355 2339 356 2343
rect 350 2338 356 2339
rect 430 2343 436 2344
rect 430 2339 431 2343
rect 435 2339 436 2343
rect 430 2338 436 2339
rect 518 2343 524 2344
rect 518 2339 519 2343
rect 523 2339 524 2343
rect 518 2338 524 2339
rect 598 2343 604 2344
rect 598 2339 599 2343
rect 603 2339 604 2343
rect 598 2338 604 2339
rect 678 2343 684 2344
rect 678 2339 679 2343
rect 683 2339 684 2343
rect 678 2338 684 2339
rect 750 2343 756 2344
rect 750 2339 751 2343
rect 755 2339 756 2343
rect 750 2338 756 2339
rect 822 2343 828 2344
rect 822 2339 823 2343
rect 827 2339 828 2343
rect 822 2338 828 2339
rect 886 2343 892 2344
rect 886 2339 887 2343
rect 891 2339 892 2343
rect 886 2338 892 2339
rect 958 2343 964 2344
rect 958 2339 959 2343
rect 963 2339 964 2343
rect 958 2338 964 2339
rect 1030 2343 1036 2344
rect 1278 2343 1284 2344
rect 1550 2343 1556 2344
rect 1030 2339 1031 2343
rect 1035 2339 1036 2343
rect 1030 2338 1036 2339
rect 1550 2339 1551 2343
rect 1555 2342 1556 2343
rect 1696 2342 1698 2348
rect 1719 2347 1720 2348
rect 1724 2347 1725 2351
rect 1719 2346 1725 2347
rect 1766 2351 1772 2352
rect 1766 2347 1767 2351
rect 1771 2350 1772 2351
rect 1799 2351 1805 2352
rect 1799 2350 1800 2351
rect 1771 2348 1800 2350
rect 1771 2347 1772 2348
rect 1766 2346 1772 2347
rect 1799 2347 1800 2348
rect 1804 2347 1805 2351
rect 1799 2346 1805 2347
rect 1807 2351 1813 2352
rect 1807 2347 1808 2351
rect 1812 2350 1813 2351
rect 1879 2351 1885 2352
rect 1879 2350 1880 2351
rect 1812 2348 1880 2350
rect 1812 2347 1813 2348
rect 1807 2346 1813 2347
rect 1879 2347 1880 2348
rect 1884 2347 1885 2351
rect 1879 2346 1885 2347
rect 1887 2351 1893 2352
rect 1887 2347 1888 2351
rect 1892 2350 1893 2351
rect 1951 2351 1957 2352
rect 1951 2350 1952 2351
rect 1892 2348 1952 2350
rect 1892 2347 1893 2348
rect 1887 2346 1893 2347
rect 1951 2347 1952 2348
rect 1956 2347 1957 2351
rect 1951 2346 1957 2347
rect 1959 2351 1965 2352
rect 1959 2347 1960 2351
rect 1964 2350 1965 2351
rect 2023 2351 2029 2352
rect 2023 2350 2024 2351
rect 1964 2348 2024 2350
rect 1964 2347 1965 2348
rect 1959 2346 1965 2347
rect 2023 2347 2024 2348
rect 2028 2347 2029 2351
rect 2023 2346 2029 2347
rect 2046 2351 2052 2352
rect 2046 2347 2047 2351
rect 2051 2350 2052 2351
rect 2095 2351 2101 2352
rect 2095 2350 2096 2351
rect 2051 2348 2096 2350
rect 2051 2347 2052 2348
rect 2046 2346 2052 2347
rect 2095 2347 2096 2348
rect 2100 2347 2101 2351
rect 2095 2346 2101 2347
rect 2103 2351 2109 2352
rect 2103 2347 2104 2351
rect 2108 2350 2109 2351
rect 2167 2351 2173 2352
rect 2167 2350 2168 2351
rect 2108 2348 2168 2350
rect 2108 2347 2109 2348
rect 2103 2346 2109 2347
rect 2167 2347 2168 2348
rect 2172 2347 2173 2351
rect 2247 2349 2248 2353
rect 2252 2352 2291 2353
rect 2252 2349 2253 2352
rect 2290 2351 2291 2352
rect 2295 2351 2296 2355
rect 2290 2350 2296 2351
rect 2310 2351 2316 2352
rect 2247 2348 2253 2349
rect 2167 2346 2173 2347
rect 2310 2347 2311 2351
rect 2315 2350 2316 2351
rect 2327 2351 2333 2352
rect 2327 2350 2328 2351
rect 2315 2348 2328 2350
rect 2315 2347 2316 2348
rect 2310 2346 2316 2347
rect 2327 2347 2328 2348
rect 2332 2347 2333 2351
rect 2327 2346 2333 2347
rect 2335 2351 2341 2352
rect 2335 2347 2336 2351
rect 2340 2350 2341 2351
rect 2383 2351 2389 2352
rect 2383 2350 2384 2351
rect 2340 2348 2384 2350
rect 2340 2347 2341 2348
rect 2335 2346 2341 2347
rect 2383 2347 2384 2348
rect 2388 2347 2389 2351
rect 2383 2346 2389 2347
rect 2406 2348 2412 2349
rect 2406 2344 2407 2348
rect 2411 2344 2412 2348
rect 2406 2343 2412 2344
rect 1555 2340 1698 2342
rect 1555 2339 1556 2340
rect 1550 2338 1556 2339
rect 1358 2325 1364 2326
rect 154 2323 160 2324
rect 110 2320 116 2321
rect 110 2316 111 2320
rect 115 2316 116 2320
rect 154 2319 155 2323
rect 159 2322 160 2323
rect 159 2320 321 2322
rect 1358 2321 1359 2325
rect 1363 2321 1364 2325
rect 159 2319 160 2320
rect 154 2318 160 2319
rect 110 2315 116 2316
rect 159 2315 168 2316
rect 159 2311 160 2315
rect 167 2311 168 2315
rect 159 2310 168 2311
rect 199 2315 208 2316
rect 199 2311 200 2315
rect 207 2311 208 2315
rect 199 2310 208 2311
rect 239 2315 245 2316
rect 239 2311 240 2315
rect 244 2314 245 2315
rect 247 2315 253 2316
rect 247 2314 248 2315
rect 244 2312 248 2314
rect 244 2311 245 2312
rect 239 2310 245 2311
rect 247 2311 248 2312
rect 252 2311 253 2315
rect 295 2315 301 2316
rect 295 2314 296 2315
rect 247 2310 253 2311
rect 256 2312 296 2314
rect 142 2307 148 2308
rect 110 2303 116 2304
rect 110 2299 111 2303
rect 115 2299 116 2303
rect 142 2303 143 2307
rect 147 2306 148 2307
rect 256 2306 258 2312
rect 295 2311 296 2312
rect 300 2311 301 2315
rect 319 2314 321 2320
rect 1238 2320 1244 2321
rect 1358 2320 1364 2321
rect 1406 2325 1412 2326
rect 1406 2321 1407 2325
rect 1411 2321 1412 2325
rect 1406 2320 1412 2321
rect 1470 2325 1476 2326
rect 1470 2321 1471 2325
rect 1475 2321 1476 2325
rect 1470 2320 1476 2321
rect 1542 2325 1548 2326
rect 1542 2321 1543 2325
rect 1547 2321 1548 2325
rect 1542 2320 1548 2321
rect 1614 2325 1620 2326
rect 1614 2321 1615 2325
rect 1619 2321 1620 2325
rect 1614 2320 1620 2321
rect 1694 2325 1700 2326
rect 1694 2321 1695 2325
rect 1699 2321 1700 2325
rect 1694 2320 1700 2321
rect 1774 2325 1780 2326
rect 1774 2321 1775 2325
rect 1779 2321 1780 2325
rect 1774 2320 1780 2321
rect 1854 2325 1860 2326
rect 1854 2321 1855 2325
rect 1859 2321 1860 2325
rect 1854 2320 1860 2321
rect 1926 2325 1932 2326
rect 1926 2321 1927 2325
rect 1931 2321 1932 2325
rect 1926 2320 1932 2321
rect 1998 2325 2004 2326
rect 1998 2321 1999 2325
rect 2003 2321 2004 2325
rect 1998 2320 2004 2321
rect 2070 2325 2076 2326
rect 2070 2321 2071 2325
rect 2075 2321 2076 2325
rect 2070 2320 2076 2321
rect 2142 2325 2148 2326
rect 2142 2321 2143 2325
rect 2147 2321 2148 2325
rect 2142 2320 2148 2321
rect 2222 2325 2228 2326
rect 2222 2321 2223 2325
rect 2227 2321 2228 2325
rect 2222 2320 2228 2321
rect 2302 2325 2308 2326
rect 2302 2321 2303 2325
rect 2307 2321 2308 2325
rect 2302 2320 2308 2321
rect 2358 2325 2364 2326
rect 2358 2321 2359 2325
rect 2363 2321 2364 2325
rect 2358 2320 2364 2321
rect 1238 2316 1239 2320
rect 1243 2316 1244 2320
rect 375 2315 381 2316
rect 375 2314 376 2315
rect 319 2312 376 2314
rect 295 2310 301 2311
rect 375 2311 376 2312
rect 380 2311 381 2315
rect 375 2310 381 2311
rect 418 2315 424 2316
rect 418 2311 419 2315
rect 423 2314 424 2315
rect 455 2315 461 2316
rect 455 2314 456 2315
rect 423 2312 456 2314
rect 423 2311 424 2312
rect 418 2310 424 2311
rect 455 2311 456 2312
rect 460 2311 461 2315
rect 455 2310 461 2311
rect 502 2315 508 2316
rect 502 2311 503 2315
rect 507 2314 508 2315
rect 543 2315 549 2316
rect 543 2314 544 2315
rect 507 2312 544 2314
rect 507 2311 508 2312
rect 502 2310 508 2311
rect 543 2311 544 2312
rect 548 2311 549 2315
rect 543 2310 549 2311
rect 590 2315 596 2316
rect 590 2311 591 2315
rect 595 2314 596 2315
rect 623 2315 629 2316
rect 623 2314 624 2315
rect 595 2312 624 2314
rect 595 2311 596 2312
rect 590 2310 596 2311
rect 623 2311 624 2312
rect 628 2311 629 2315
rect 623 2310 629 2311
rect 666 2315 672 2316
rect 666 2311 667 2315
rect 671 2314 672 2315
rect 703 2315 709 2316
rect 703 2314 704 2315
rect 671 2312 704 2314
rect 671 2311 672 2312
rect 666 2310 672 2311
rect 703 2311 704 2312
rect 708 2311 709 2315
rect 703 2310 709 2311
rect 726 2315 732 2316
rect 726 2311 727 2315
rect 731 2314 732 2315
rect 775 2315 781 2316
rect 775 2314 776 2315
rect 731 2312 776 2314
rect 731 2311 732 2312
rect 726 2310 732 2311
rect 775 2311 776 2312
rect 780 2311 781 2315
rect 775 2310 781 2311
rect 847 2315 856 2316
rect 847 2311 848 2315
rect 855 2311 856 2315
rect 847 2310 856 2311
rect 911 2315 920 2316
rect 911 2311 912 2315
rect 919 2311 920 2315
rect 911 2310 920 2311
rect 983 2315 989 2316
rect 983 2311 984 2315
rect 988 2314 989 2315
rect 991 2315 997 2316
rect 991 2314 992 2315
rect 988 2312 992 2314
rect 988 2311 989 2312
rect 983 2310 989 2311
rect 991 2311 992 2312
rect 996 2311 997 2315
rect 991 2310 997 2311
rect 1002 2315 1008 2316
rect 1002 2311 1003 2315
rect 1007 2314 1008 2315
rect 1055 2315 1061 2316
rect 1238 2315 1244 2316
rect 1355 2315 1361 2316
rect 1055 2314 1056 2315
rect 1007 2312 1056 2314
rect 1007 2311 1008 2312
rect 1002 2310 1008 2311
rect 1055 2311 1056 2312
rect 1060 2311 1061 2315
rect 1055 2310 1061 2311
rect 1355 2311 1356 2315
rect 1360 2314 1361 2315
rect 1391 2315 1397 2316
rect 1391 2314 1392 2315
rect 1360 2312 1392 2314
rect 1360 2311 1361 2312
rect 1355 2310 1361 2311
rect 1391 2311 1392 2312
rect 1396 2311 1397 2315
rect 1391 2310 1397 2311
rect 1403 2315 1409 2316
rect 1403 2311 1404 2315
rect 1408 2314 1409 2315
rect 1439 2315 1445 2316
rect 1439 2314 1440 2315
rect 1408 2312 1440 2314
rect 1408 2311 1409 2312
rect 1403 2310 1409 2311
rect 1439 2311 1440 2312
rect 1444 2311 1445 2315
rect 1439 2310 1445 2311
rect 1467 2315 1473 2316
rect 1467 2311 1468 2315
rect 1472 2314 1473 2315
rect 1503 2315 1509 2316
rect 1503 2314 1504 2315
rect 1472 2312 1504 2314
rect 1472 2311 1473 2312
rect 1467 2310 1473 2311
rect 1503 2311 1504 2312
rect 1508 2311 1509 2315
rect 1503 2310 1509 2311
rect 1539 2315 1545 2316
rect 1539 2311 1540 2315
rect 1544 2314 1545 2315
rect 1550 2315 1556 2316
rect 1550 2314 1551 2315
rect 1544 2312 1551 2314
rect 1544 2311 1545 2312
rect 1539 2310 1545 2311
rect 1550 2311 1551 2312
rect 1555 2311 1556 2315
rect 1550 2310 1556 2311
rect 1606 2315 1617 2316
rect 1606 2311 1607 2315
rect 1611 2311 1612 2315
rect 1616 2311 1617 2315
rect 1606 2310 1617 2311
rect 1686 2315 1697 2316
rect 1686 2311 1687 2315
rect 1691 2311 1692 2315
rect 1696 2311 1697 2315
rect 1686 2310 1697 2311
rect 1771 2315 1777 2316
rect 1771 2311 1772 2315
rect 1776 2314 1777 2315
rect 1807 2315 1813 2316
rect 1807 2314 1808 2315
rect 1776 2312 1808 2314
rect 1776 2311 1777 2312
rect 1771 2310 1777 2311
rect 1807 2311 1808 2312
rect 1812 2311 1813 2315
rect 1807 2310 1813 2311
rect 1851 2315 1857 2316
rect 1851 2311 1852 2315
rect 1856 2314 1857 2315
rect 1887 2315 1893 2316
rect 1887 2314 1888 2315
rect 1856 2312 1888 2314
rect 1856 2311 1857 2312
rect 1851 2310 1857 2311
rect 1887 2311 1888 2312
rect 1892 2311 1893 2315
rect 1887 2310 1893 2311
rect 1923 2315 1929 2316
rect 1923 2311 1924 2315
rect 1928 2314 1929 2315
rect 1959 2315 1965 2316
rect 1959 2314 1960 2315
rect 1928 2312 1960 2314
rect 1928 2311 1929 2312
rect 1923 2310 1929 2311
rect 1959 2311 1960 2312
rect 1964 2311 1965 2315
rect 1959 2310 1965 2311
rect 1995 2315 2001 2316
rect 1995 2311 1996 2315
rect 2000 2314 2001 2315
rect 2046 2315 2052 2316
rect 2046 2314 2047 2315
rect 2000 2312 2047 2314
rect 2000 2311 2001 2312
rect 1995 2310 2001 2311
rect 2046 2311 2047 2312
rect 2051 2311 2052 2315
rect 2046 2310 2052 2311
rect 2067 2315 2073 2316
rect 2067 2311 2068 2315
rect 2072 2314 2073 2315
rect 2103 2315 2109 2316
rect 2103 2314 2104 2315
rect 2072 2312 2104 2314
rect 2072 2311 2073 2312
rect 2067 2310 2073 2311
rect 2103 2311 2104 2312
rect 2108 2311 2109 2315
rect 2103 2310 2109 2311
rect 2139 2315 2145 2316
rect 2139 2311 2140 2315
rect 2144 2314 2145 2315
rect 2191 2315 2197 2316
rect 2191 2314 2192 2315
rect 2144 2312 2192 2314
rect 2144 2311 2145 2312
rect 2139 2310 2145 2311
rect 2191 2311 2192 2312
rect 2196 2311 2197 2315
rect 2191 2310 2197 2311
rect 2219 2315 2225 2316
rect 2219 2311 2220 2315
rect 2224 2314 2225 2315
rect 2230 2315 2236 2316
rect 2230 2314 2231 2315
rect 2224 2312 2231 2314
rect 2224 2311 2225 2312
rect 2219 2310 2225 2311
rect 2230 2311 2231 2312
rect 2235 2311 2236 2315
rect 2230 2310 2236 2311
rect 2299 2315 2305 2316
rect 2299 2311 2300 2315
rect 2304 2314 2305 2315
rect 2335 2315 2341 2316
rect 2335 2314 2336 2315
rect 2304 2312 2336 2314
rect 2304 2311 2305 2312
rect 2299 2310 2305 2311
rect 2335 2311 2336 2312
rect 2340 2311 2341 2315
rect 2335 2310 2341 2311
rect 2350 2315 2361 2316
rect 2350 2311 2351 2315
rect 2355 2311 2356 2315
rect 2360 2311 2361 2315
rect 2350 2310 2361 2311
rect 147 2304 258 2306
rect 147 2303 148 2304
rect 142 2302 148 2303
rect 1238 2303 1244 2304
rect 110 2298 116 2299
rect 1238 2299 1239 2303
rect 1243 2299 1244 2303
rect 1238 2298 1244 2299
rect 1499 2299 1505 2300
rect 134 2296 140 2297
rect 134 2292 135 2296
rect 139 2292 140 2296
rect 134 2291 140 2292
rect 174 2296 180 2297
rect 174 2292 175 2296
rect 179 2292 180 2296
rect 174 2291 180 2292
rect 214 2296 220 2297
rect 214 2292 215 2296
rect 219 2292 220 2296
rect 214 2291 220 2292
rect 270 2296 276 2297
rect 270 2292 271 2296
rect 275 2292 276 2296
rect 270 2291 276 2292
rect 350 2296 356 2297
rect 350 2292 351 2296
rect 355 2292 356 2296
rect 350 2291 356 2292
rect 430 2296 436 2297
rect 430 2292 431 2296
rect 435 2292 436 2296
rect 430 2291 436 2292
rect 518 2296 524 2297
rect 518 2292 519 2296
rect 523 2292 524 2296
rect 518 2291 524 2292
rect 598 2296 604 2297
rect 598 2292 599 2296
rect 603 2292 604 2296
rect 598 2291 604 2292
rect 678 2296 684 2297
rect 678 2292 679 2296
rect 683 2292 684 2296
rect 678 2291 684 2292
rect 750 2296 756 2297
rect 750 2292 751 2296
rect 755 2292 756 2296
rect 750 2291 756 2292
rect 822 2296 828 2297
rect 822 2292 823 2296
rect 827 2292 828 2296
rect 822 2291 828 2292
rect 886 2296 892 2297
rect 886 2292 887 2296
rect 891 2292 892 2296
rect 886 2291 892 2292
rect 958 2296 964 2297
rect 958 2292 959 2296
rect 963 2292 964 2296
rect 958 2291 964 2292
rect 1030 2296 1036 2297
rect 1030 2292 1031 2296
rect 1035 2292 1036 2296
rect 1499 2295 1500 2299
rect 1504 2298 1505 2299
rect 1522 2299 1528 2300
rect 1522 2298 1523 2299
rect 1504 2296 1523 2298
rect 1504 2295 1505 2296
rect 1499 2294 1505 2295
rect 1522 2295 1523 2296
rect 1527 2295 1528 2299
rect 1522 2294 1528 2295
rect 1530 2299 1536 2300
rect 1530 2295 1531 2299
rect 1535 2298 1536 2299
rect 1539 2299 1545 2300
rect 1539 2298 1540 2299
rect 1535 2296 1540 2298
rect 1535 2295 1536 2296
rect 1530 2294 1536 2295
rect 1539 2295 1540 2296
rect 1544 2295 1545 2299
rect 1539 2294 1545 2295
rect 1566 2299 1572 2300
rect 1566 2295 1567 2299
rect 1571 2298 1572 2299
rect 1579 2299 1585 2300
rect 1579 2298 1580 2299
rect 1571 2296 1580 2298
rect 1571 2295 1572 2296
rect 1566 2294 1572 2295
rect 1579 2295 1580 2296
rect 1584 2295 1585 2299
rect 1579 2294 1585 2295
rect 1619 2299 1625 2300
rect 1619 2295 1620 2299
rect 1624 2298 1625 2299
rect 1646 2299 1652 2300
rect 1646 2298 1647 2299
rect 1624 2296 1647 2298
rect 1624 2295 1625 2296
rect 1619 2294 1625 2295
rect 1646 2295 1647 2296
rect 1651 2295 1652 2299
rect 1646 2294 1652 2295
rect 1654 2299 1665 2300
rect 1654 2295 1655 2299
rect 1659 2295 1660 2299
rect 1664 2295 1665 2299
rect 1654 2294 1665 2295
rect 1686 2299 1692 2300
rect 1686 2295 1687 2299
rect 1691 2298 1692 2299
rect 1699 2299 1705 2300
rect 1699 2298 1700 2299
rect 1691 2296 1700 2298
rect 1691 2295 1692 2296
rect 1686 2294 1692 2295
rect 1699 2295 1700 2296
rect 1704 2295 1705 2299
rect 1699 2294 1705 2295
rect 1755 2299 1761 2300
rect 1755 2295 1756 2299
rect 1760 2298 1761 2299
rect 1766 2299 1772 2300
rect 1766 2298 1767 2299
rect 1760 2296 1767 2298
rect 1760 2295 1761 2296
rect 1755 2294 1761 2295
rect 1766 2295 1767 2296
rect 1771 2295 1772 2299
rect 1766 2294 1772 2295
rect 1786 2299 1792 2300
rect 1786 2295 1787 2299
rect 1791 2298 1792 2299
rect 1819 2299 1825 2300
rect 1819 2298 1820 2299
rect 1791 2296 1820 2298
rect 1791 2295 1792 2296
rect 1786 2294 1792 2295
rect 1819 2295 1820 2296
rect 1824 2295 1825 2299
rect 1819 2294 1825 2295
rect 1855 2299 1861 2300
rect 1855 2295 1856 2299
rect 1860 2298 1861 2299
rect 1891 2299 1897 2300
rect 1891 2298 1892 2299
rect 1860 2296 1892 2298
rect 1860 2295 1861 2296
rect 1855 2294 1861 2295
rect 1891 2295 1892 2296
rect 1896 2295 1897 2299
rect 1891 2294 1897 2295
rect 1927 2299 1933 2300
rect 1927 2295 1928 2299
rect 1932 2298 1933 2299
rect 1963 2299 1969 2300
rect 1963 2298 1964 2299
rect 1932 2296 1964 2298
rect 1932 2295 1933 2296
rect 1927 2294 1933 2295
rect 1963 2295 1964 2296
rect 1968 2295 1969 2299
rect 1963 2294 1969 2295
rect 2018 2299 2024 2300
rect 2018 2295 2019 2299
rect 2023 2298 2024 2299
rect 2043 2299 2049 2300
rect 2043 2298 2044 2299
rect 2023 2296 2044 2298
rect 2023 2295 2024 2296
rect 2018 2294 2024 2295
rect 2043 2295 2044 2296
rect 2048 2295 2049 2299
rect 2043 2294 2049 2295
rect 2123 2299 2129 2300
rect 2123 2295 2124 2299
rect 2128 2298 2129 2299
rect 2134 2299 2140 2300
rect 2134 2298 2135 2299
rect 2128 2296 2135 2298
rect 2128 2295 2129 2296
rect 2123 2294 2129 2295
rect 2134 2295 2135 2296
rect 2139 2295 2140 2299
rect 2134 2294 2140 2295
rect 2154 2299 2160 2300
rect 2154 2295 2155 2299
rect 2159 2298 2160 2299
rect 2203 2299 2209 2300
rect 2203 2298 2204 2299
rect 2159 2296 2204 2298
rect 2159 2295 2160 2296
rect 2154 2294 2160 2295
rect 2203 2295 2204 2296
rect 2208 2295 2209 2299
rect 2203 2294 2209 2295
rect 2291 2299 2297 2300
rect 2291 2295 2292 2299
rect 2296 2298 2297 2299
rect 2310 2299 2316 2300
rect 2310 2298 2311 2299
rect 2296 2296 2311 2298
rect 2296 2295 2297 2296
rect 2291 2294 2297 2295
rect 2310 2295 2311 2296
rect 2315 2295 2316 2299
rect 2310 2294 2316 2295
rect 2322 2299 2328 2300
rect 2322 2295 2323 2299
rect 2327 2298 2328 2299
rect 2355 2299 2361 2300
rect 2355 2298 2356 2299
rect 2327 2296 2356 2298
rect 2327 2295 2328 2296
rect 2322 2294 2328 2295
rect 2355 2295 2356 2296
rect 2360 2295 2361 2299
rect 2355 2294 2361 2295
rect 1030 2291 1036 2292
rect 1502 2291 1508 2292
rect 1502 2287 1503 2291
rect 1507 2287 1508 2291
rect 1502 2286 1508 2287
rect 1542 2291 1548 2292
rect 1542 2287 1543 2291
rect 1547 2287 1548 2291
rect 1542 2286 1548 2287
rect 1582 2291 1588 2292
rect 1582 2287 1583 2291
rect 1587 2287 1588 2291
rect 1582 2286 1588 2287
rect 1622 2291 1628 2292
rect 1622 2287 1623 2291
rect 1627 2287 1628 2291
rect 1622 2286 1628 2287
rect 1662 2291 1668 2292
rect 1662 2287 1663 2291
rect 1667 2287 1668 2291
rect 1662 2286 1668 2287
rect 1702 2291 1708 2292
rect 1702 2287 1703 2291
rect 1707 2287 1708 2291
rect 1702 2286 1708 2287
rect 1758 2291 1764 2292
rect 1758 2287 1759 2291
rect 1763 2287 1764 2291
rect 1758 2286 1764 2287
rect 1822 2291 1828 2292
rect 1822 2287 1823 2291
rect 1827 2287 1828 2291
rect 1822 2286 1828 2287
rect 1894 2291 1900 2292
rect 1894 2287 1895 2291
rect 1899 2287 1900 2291
rect 1894 2286 1900 2287
rect 1966 2291 1972 2292
rect 1966 2287 1967 2291
rect 1971 2287 1972 2291
rect 1966 2286 1972 2287
rect 2046 2291 2052 2292
rect 2046 2287 2047 2291
rect 2051 2287 2052 2291
rect 2046 2286 2052 2287
rect 2126 2291 2132 2292
rect 2126 2287 2127 2291
rect 2131 2287 2132 2291
rect 2126 2286 2132 2287
rect 2206 2291 2212 2292
rect 2206 2287 2207 2291
rect 2211 2287 2212 2291
rect 2206 2286 2212 2287
rect 2294 2291 2300 2292
rect 2294 2287 2295 2291
rect 2299 2287 2300 2291
rect 2294 2286 2300 2287
rect 2358 2291 2364 2292
rect 2358 2287 2359 2291
rect 2363 2287 2364 2291
rect 2358 2286 2364 2287
rect 134 2280 140 2281
rect 134 2276 135 2280
rect 139 2276 140 2280
rect 134 2275 140 2276
rect 174 2280 180 2281
rect 174 2276 175 2280
rect 179 2276 180 2280
rect 174 2275 180 2276
rect 230 2280 236 2281
rect 230 2276 231 2280
rect 235 2276 236 2280
rect 230 2275 236 2276
rect 302 2280 308 2281
rect 302 2276 303 2280
rect 307 2276 308 2280
rect 302 2275 308 2276
rect 374 2280 380 2281
rect 374 2276 375 2280
rect 379 2276 380 2280
rect 374 2275 380 2276
rect 454 2280 460 2281
rect 454 2276 455 2280
rect 459 2276 460 2280
rect 454 2275 460 2276
rect 534 2280 540 2281
rect 534 2276 535 2280
rect 539 2276 540 2280
rect 534 2275 540 2276
rect 614 2280 620 2281
rect 614 2276 615 2280
rect 619 2276 620 2280
rect 614 2275 620 2276
rect 686 2280 692 2281
rect 686 2276 687 2280
rect 691 2276 692 2280
rect 686 2275 692 2276
rect 758 2280 764 2281
rect 758 2276 759 2280
rect 763 2276 764 2280
rect 758 2275 764 2276
rect 830 2280 836 2281
rect 830 2276 831 2280
rect 835 2276 836 2280
rect 830 2275 836 2276
rect 910 2280 916 2281
rect 910 2276 911 2280
rect 915 2276 916 2280
rect 910 2275 916 2276
rect 990 2280 996 2281
rect 990 2276 991 2280
rect 995 2276 996 2280
rect 990 2275 996 2276
rect 110 2273 116 2274
rect 110 2269 111 2273
rect 115 2269 116 2273
rect 110 2268 116 2269
rect 1238 2273 1244 2274
rect 1238 2269 1239 2273
rect 1243 2269 1244 2273
rect 1522 2271 1528 2272
rect 1238 2268 1244 2269
rect 1278 2268 1284 2269
rect 1278 2264 1279 2268
rect 1283 2264 1284 2268
rect 1522 2267 1523 2271
rect 1527 2270 1528 2271
rect 1646 2271 1652 2272
rect 1527 2268 1618 2270
rect 1527 2267 1528 2268
rect 1522 2266 1528 2267
rect 1278 2263 1284 2264
rect 1527 2263 1536 2264
rect 159 2259 168 2260
rect 110 2256 116 2257
rect 110 2252 111 2256
rect 115 2252 116 2256
rect 159 2255 160 2259
rect 167 2255 168 2259
rect 159 2254 168 2255
rect 199 2259 205 2260
rect 199 2255 200 2259
rect 204 2258 205 2259
rect 214 2259 220 2260
rect 214 2258 215 2259
rect 204 2256 215 2258
rect 204 2255 205 2256
rect 199 2254 205 2255
rect 214 2255 215 2256
rect 219 2255 220 2259
rect 214 2254 220 2255
rect 255 2259 261 2260
rect 255 2255 256 2259
rect 260 2258 261 2259
rect 294 2259 300 2260
rect 294 2258 295 2259
rect 260 2256 295 2258
rect 260 2255 261 2256
rect 255 2254 261 2255
rect 294 2255 295 2256
rect 299 2255 300 2259
rect 294 2254 300 2255
rect 327 2259 333 2260
rect 327 2255 328 2259
rect 332 2258 333 2259
rect 366 2259 372 2260
rect 366 2258 367 2259
rect 332 2256 367 2258
rect 332 2255 333 2256
rect 327 2254 333 2255
rect 366 2255 367 2256
rect 371 2255 372 2259
rect 366 2254 372 2255
rect 399 2259 405 2260
rect 399 2255 400 2259
rect 404 2258 405 2259
rect 446 2259 452 2260
rect 446 2258 447 2259
rect 404 2256 447 2258
rect 404 2255 405 2256
rect 399 2254 405 2255
rect 446 2255 447 2256
rect 451 2255 452 2259
rect 479 2259 485 2260
rect 479 2258 480 2259
rect 446 2254 452 2255
rect 456 2256 480 2258
rect 110 2251 116 2252
rect 254 2251 260 2252
rect 254 2247 255 2251
rect 259 2250 260 2251
rect 456 2250 458 2256
rect 479 2255 480 2256
rect 484 2255 485 2259
rect 479 2254 485 2255
rect 559 2259 565 2260
rect 559 2255 560 2259
rect 564 2258 565 2259
rect 599 2259 605 2260
rect 599 2258 600 2259
rect 564 2256 600 2258
rect 564 2255 565 2256
rect 559 2254 565 2255
rect 599 2255 600 2256
rect 604 2255 605 2259
rect 599 2254 605 2255
rect 639 2259 645 2260
rect 639 2255 640 2259
rect 644 2258 645 2259
rect 678 2259 684 2260
rect 678 2258 679 2259
rect 644 2256 679 2258
rect 644 2255 645 2256
rect 639 2254 645 2255
rect 678 2255 679 2256
rect 683 2255 684 2259
rect 678 2254 684 2255
rect 711 2259 717 2260
rect 711 2255 712 2259
rect 716 2258 717 2259
rect 750 2259 756 2260
rect 750 2258 751 2259
rect 716 2256 751 2258
rect 716 2255 717 2256
rect 711 2254 717 2255
rect 750 2255 751 2256
rect 755 2255 756 2259
rect 750 2254 756 2255
rect 782 2259 789 2260
rect 782 2255 783 2259
rect 788 2255 789 2259
rect 782 2254 789 2255
rect 854 2259 861 2260
rect 854 2255 855 2259
rect 860 2255 861 2259
rect 854 2254 861 2255
rect 863 2259 869 2260
rect 863 2255 864 2259
rect 868 2258 869 2259
rect 935 2259 941 2260
rect 935 2258 936 2259
rect 868 2256 936 2258
rect 868 2255 869 2256
rect 863 2254 869 2255
rect 935 2255 936 2256
rect 940 2255 941 2259
rect 935 2254 941 2255
rect 943 2259 949 2260
rect 943 2255 944 2259
rect 948 2258 949 2259
rect 1015 2259 1021 2260
rect 1015 2258 1016 2259
rect 948 2256 1016 2258
rect 948 2255 949 2256
rect 943 2254 949 2255
rect 1015 2255 1016 2256
rect 1020 2255 1021 2259
rect 1527 2259 1528 2263
rect 1535 2259 1536 2263
rect 1527 2258 1536 2259
rect 1566 2263 1573 2264
rect 1566 2259 1567 2263
rect 1572 2259 1573 2263
rect 1566 2258 1573 2259
rect 1606 2263 1613 2264
rect 1606 2259 1607 2263
rect 1612 2259 1613 2263
rect 1616 2262 1618 2268
rect 1646 2267 1647 2271
rect 1651 2270 1652 2271
rect 1651 2268 1698 2270
rect 1651 2267 1652 2268
rect 1646 2266 1652 2267
rect 1647 2263 1653 2264
rect 1647 2262 1648 2263
rect 1616 2260 1648 2262
rect 1606 2258 1613 2259
rect 1647 2259 1648 2260
rect 1652 2259 1653 2263
rect 1647 2258 1653 2259
rect 1686 2263 1693 2264
rect 1686 2259 1687 2263
rect 1692 2259 1693 2263
rect 1696 2262 1698 2268
rect 2406 2268 2412 2269
rect 2406 2264 2407 2268
rect 2411 2264 2412 2268
rect 1727 2263 1733 2264
rect 1727 2262 1728 2263
rect 1696 2260 1728 2262
rect 1686 2258 1693 2259
rect 1727 2259 1728 2260
rect 1732 2259 1733 2263
rect 1727 2258 1733 2259
rect 1783 2263 1792 2264
rect 1783 2259 1784 2263
rect 1791 2259 1792 2263
rect 1783 2258 1792 2259
rect 1847 2263 1853 2264
rect 1847 2259 1848 2263
rect 1852 2262 1853 2263
rect 1855 2263 1861 2264
rect 1855 2262 1856 2263
rect 1852 2260 1856 2262
rect 1852 2259 1853 2260
rect 1847 2258 1853 2259
rect 1855 2259 1856 2260
rect 1860 2259 1861 2263
rect 1855 2258 1861 2259
rect 1919 2263 1925 2264
rect 1919 2259 1920 2263
rect 1924 2262 1925 2263
rect 1927 2263 1933 2264
rect 1927 2262 1928 2263
rect 1924 2260 1928 2262
rect 1924 2259 1925 2260
rect 1919 2258 1925 2259
rect 1927 2259 1928 2260
rect 1932 2259 1933 2263
rect 1927 2258 1933 2259
rect 1991 2263 1997 2264
rect 1991 2259 1992 2263
rect 1996 2262 1997 2263
rect 2018 2263 2024 2264
rect 2018 2262 2019 2263
rect 1996 2260 2019 2262
rect 1996 2259 1997 2260
rect 1991 2258 1997 2259
rect 2018 2259 2019 2260
rect 2023 2259 2024 2263
rect 2071 2263 2077 2264
rect 2071 2262 2072 2263
rect 2018 2258 2024 2259
rect 2036 2260 2072 2262
rect 1015 2254 1021 2255
rect 1238 2256 1244 2257
rect 1238 2252 1239 2256
rect 1243 2252 1244 2256
rect 1790 2255 1796 2256
rect 1238 2251 1244 2252
rect 1278 2251 1284 2252
rect 259 2248 458 2250
rect 259 2247 260 2248
rect 254 2246 260 2247
rect 1278 2247 1279 2251
rect 1283 2247 1284 2251
rect 1790 2251 1791 2255
rect 1795 2254 1796 2255
rect 2036 2254 2038 2260
rect 2071 2259 2072 2260
rect 2076 2259 2077 2263
rect 2071 2258 2077 2259
rect 2151 2263 2160 2264
rect 2151 2259 2152 2263
rect 2159 2259 2160 2263
rect 2151 2258 2160 2259
rect 2230 2263 2237 2264
rect 2230 2259 2231 2263
rect 2236 2259 2237 2263
rect 2230 2258 2237 2259
rect 2319 2263 2328 2264
rect 2319 2259 2320 2263
rect 2327 2259 2328 2263
rect 2319 2258 2328 2259
rect 2366 2263 2372 2264
rect 2366 2259 2367 2263
rect 2371 2262 2372 2263
rect 2383 2263 2389 2264
rect 2406 2263 2412 2264
rect 2383 2262 2384 2263
rect 2371 2260 2384 2262
rect 2371 2259 2372 2260
rect 2366 2258 2372 2259
rect 2383 2259 2384 2260
rect 2388 2259 2389 2263
rect 2383 2258 2389 2259
rect 1795 2252 2038 2254
rect 1795 2251 1796 2252
rect 1790 2250 1796 2251
rect 2406 2251 2412 2252
rect 1278 2246 1284 2247
rect 2406 2247 2407 2251
rect 2411 2247 2412 2251
rect 2406 2246 2412 2247
rect 1502 2244 1508 2245
rect 1502 2240 1503 2244
rect 1507 2240 1508 2244
rect 1502 2239 1508 2240
rect 1542 2244 1548 2245
rect 1542 2240 1543 2244
rect 1547 2240 1548 2244
rect 1542 2239 1548 2240
rect 1582 2244 1588 2245
rect 1582 2240 1583 2244
rect 1587 2240 1588 2244
rect 1582 2239 1588 2240
rect 1622 2244 1628 2245
rect 1622 2240 1623 2244
rect 1627 2240 1628 2244
rect 1622 2239 1628 2240
rect 1662 2244 1668 2245
rect 1662 2240 1663 2244
rect 1667 2240 1668 2244
rect 1662 2239 1668 2240
rect 1702 2244 1708 2245
rect 1702 2240 1703 2244
rect 1707 2240 1708 2244
rect 1702 2239 1708 2240
rect 1758 2244 1764 2245
rect 1758 2240 1759 2244
rect 1763 2240 1764 2244
rect 1758 2239 1764 2240
rect 1822 2244 1828 2245
rect 1822 2240 1823 2244
rect 1827 2240 1828 2244
rect 1822 2239 1828 2240
rect 1894 2244 1900 2245
rect 1894 2240 1895 2244
rect 1899 2240 1900 2244
rect 1894 2239 1900 2240
rect 1966 2244 1972 2245
rect 1966 2240 1967 2244
rect 1971 2240 1972 2244
rect 1966 2239 1972 2240
rect 2046 2244 2052 2245
rect 2046 2240 2047 2244
rect 2051 2240 2052 2244
rect 2046 2239 2052 2240
rect 2126 2244 2132 2245
rect 2126 2240 2127 2244
rect 2131 2240 2132 2244
rect 2126 2239 2132 2240
rect 2206 2244 2212 2245
rect 2206 2240 2207 2244
rect 2211 2240 2212 2244
rect 2206 2239 2212 2240
rect 2294 2244 2300 2245
rect 2294 2240 2295 2244
rect 2299 2240 2300 2244
rect 2294 2239 2300 2240
rect 2358 2244 2364 2245
rect 2358 2240 2359 2244
rect 2363 2240 2364 2244
rect 2358 2239 2364 2240
rect 134 2233 140 2234
rect 134 2229 135 2233
rect 139 2229 140 2233
rect 134 2228 140 2229
rect 174 2233 180 2234
rect 174 2229 175 2233
rect 179 2229 180 2233
rect 174 2228 180 2229
rect 230 2233 236 2234
rect 230 2229 231 2233
rect 235 2229 236 2233
rect 230 2228 236 2229
rect 302 2233 308 2234
rect 302 2229 303 2233
rect 307 2229 308 2233
rect 302 2228 308 2229
rect 374 2233 380 2234
rect 374 2229 375 2233
rect 379 2229 380 2233
rect 374 2228 380 2229
rect 454 2233 460 2234
rect 454 2229 455 2233
rect 459 2229 460 2233
rect 454 2228 460 2229
rect 534 2233 540 2234
rect 534 2229 535 2233
rect 539 2229 540 2233
rect 534 2228 540 2229
rect 614 2233 620 2234
rect 614 2229 615 2233
rect 619 2229 620 2233
rect 614 2228 620 2229
rect 686 2233 692 2234
rect 686 2229 687 2233
rect 691 2229 692 2233
rect 686 2228 692 2229
rect 758 2233 764 2234
rect 758 2229 759 2233
rect 763 2229 764 2233
rect 758 2228 764 2229
rect 830 2233 836 2234
rect 830 2229 831 2233
rect 835 2229 836 2233
rect 830 2228 836 2229
rect 910 2233 916 2234
rect 910 2229 911 2233
rect 915 2229 916 2233
rect 910 2228 916 2229
rect 990 2233 996 2234
rect 990 2229 991 2233
rect 995 2229 996 2233
rect 990 2228 996 2229
rect 1302 2224 1308 2225
rect 131 2223 137 2224
rect 131 2219 132 2223
rect 136 2222 137 2223
rect 142 2223 148 2224
rect 142 2222 143 2223
rect 136 2220 143 2222
rect 136 2219 137 2220
rect 131 2218 137 2219
rect 142 2219 143 2220
rect 147 2219 148 2223
rect 142 2218 148 2219
rect 162 2223 168 2224
rect 162 2219 163 2223
rect 167 2222 168 2223
rect 171 2223 177 2224
rect 171 2222 172 2223
rect 167 2220 172 2222
rect 167 2219 168 2220
rect 162 2218 168 2219
rect 171 2219 172 2220
rect 176 2219 177 2223
rect 171 2218 177 2219
rect 214 2223 220 2224
rect 214 2219 215 2223
rect 219 2222 220 2223
rect 227 2223 233 2224
rect 227 2222 228 2223
rect 219 2220 228 2222
rect 219 2219 220 2220
rect 214 2218 220 2219
rect 227 2219 228 2220
rect 232 2219 233 2223
rect 227 2218 233 2219
rect 294 2223 305 2224
rect 294 2219 295 2223
rect 299 2219 300 2223
rect 304 2219 305 2223
rect 294 2218 305 2219
rect 366 2223 377 2224
rect 366 2219 367 2223
rect 371 2219 372 2223
rect 376 2219 377 2223
rect 366 2218 377 2219
rect 446 2223 457 2224
rect 446 2219 447 2223
rect 451 2219 452 2223
rect 456 2219 457 2223
rect 446 2218 457 2219
rect 531 2223 537 2224
rect 531 2219 532 2223
rect 536 2222 537 2223
rect 591 2223 597 2224
rect 591 2222 592 2223
rect 536 2220 592 2222
rect 536 2219 537 2220
rect 531 2218 537 2219
rect 591 2219 592 2220
rect 596 2219 597 2223
rect 591 2218 597 2219
rect 599 2223 605 2224
rect 599 2219 600 2223
rect 604 2222 605 2223
rect 611 2223 617 2224
rect 611 2222 612 2223
rect 604 2220 612 2222
rect 604 2219 605 2220
rect 599 2218 605 2219
rect 611 2219 612 2220
rect 616 2219 617 2223
rect 611 2218 617 2219
rect 678 2223 689 2224
rect 678 2219 679 2223
rect 683 2219 684 2223
rect 688 2219 689 2223
rect 678 2218 689 2219
rect 750 2223 761 2224
rect 750 2219 751 2223
rect 755 2219 756 2223
rect 760 2219 761 2223
rect 750 2218 761 2219
rect 827 2223 833 2224
rect 827 2219 828 2223
rect 832 2222 833 2223
rect 863 2223 869 2224
rect 863 2222 864 2223
rect 832 2220 864 2222
rect 832 2219 833 2220
rect 827 2218 833 2219
rect 863 2219 864 2220
rect 868 2219 869 2223
rect 863 2218 869 2219
rect 907 2223 913 2224
rect 907 2219 908 2223
rect 912 2222 913 2223
rect 943 2223 949 2224
rect 943 2222 944 2223
rect 912 2220 944 2222
rect 912 2219 913 2220
rect 907 2218 913 2219
rect 943 2219 944 2220
rect 948 2219 949 2223
rect 943 2218 949 2219
rect 987 2223 993 2224
rect 987 2219 988 2223
rect 992 2222 993 2223
rect 1002 2223 1008 2224
rect 1002 2222 1003 2223
rect 992 2220 1003 2222
rect 992 2219 993 2220
rect 987 2218 993 2219
rect 1002 2219 1003 2220
rect 1007 2219 1008 2223
rect 1302 2220 1303 2224
rect 1307 2220 1308 2224
rect 1302 2219 1308 2220
rect 1342 2224 1348 2225
rect 1342 2220 1343 2224
rect 1347 2220 1348 2224
rect 1342 2219 1348 2220
rect 1382 2224 1388 2225
rect 1382 2220 1383 2224
rect 1387 2220 1388 2224
rect 1382 2219 1388 2220
rect 1430 2224 1436 2225
rect 1430 2220 1431 2224
rect 1435 2220 1436 2224
rect 1430 2219 1436 2220
rect 1494 2224 1500 2225
rect 1494 2220 1495 2224
rect 1499 2220 1500 2224
rect 1494 2219 1500 2220
rect 1566 2224 1572 2225
rect 1566 2220 1567 2224
rect 1571 2220 1572 2224
rect 1566 2219 1572 2220
rect 1638 2224 1644 2225
rect 1638 2220 1639 2224
rect 1643 2220 1644 2224
rect 1638 2219 1644 2220
rect 1710 2224 1716 2225
rect 1710 2220 1711 2224
rect 1715 2220 1716 2224
rect 1710 2219 1716 2220
rect 1782 2224 1788 2225
rect 1782 2220 1783 2224
rect 1787 2220 1788 2224
rect 1782 2219 1788 2220
rect 1854 2224 1860 2225
rect 1854 2220 1855 2224
rect 1859 2220 1860 2224
rect 1854 2219 1860 2220
rect 1934 2224 1940 2225
rect 1934 2220 1935 2224
rect 1939 2220 1940 2224
rect 1934 2219 1940 2220
rect 2014 2224 2020 2225
rect 2014 2220 2015 2224
rect 2019 2220 2020 2224
rect 2014 2219 2020 2220
rect 2094 2224 2100 2225
rect 2094 2220 2095 2224
rect 2099 2220 2100 2224
rect 2094 2219 2100 2220
rect 2182 2224 2188 2225
rect 2182 2220 2183 2224
rect 2187 2220 2188 2224
rect 2182 2219 2188 2220
rect 2278 2224 2284 2225
rect 2278 2220 2279 2224
rect 2283 2220 2284 2224
rect 2278 2219 2284 2220
rect 2358 2224 2364 2225
rect 2358 2220 2359 2224
rect 2363 2220 2364 2224
rect 2358 2219 2364 2220
rect 1002 2218 1008 2219
rect 1278 2217 1284 2218
rect 1278 2213 1279 2217
rect 1283 2213 1284 2217
rect 1278 2212 1284 2213
rect 2406 2217 2412 2218
rect 2406 2213 2407 2217
rect 2411 2213 2412 2217
rect 2406 2212 2412 2213
rect 243 2211 249 2212
rect 243 2207 244 2211
rect 248 2210 249 2211
rect 254 2211 260 2212
rect 254 2210 255 2211
rect 248 2208 255 2210
rect 248 2207 249 2208
rect 243 2206 249 2207
rect 254 2207 255 2208
rect 259 2207 260 2211
rect 254 2206 260 2207
rect 274 2211 280 2212
rect 274 2207 275 2211
rect 279 2210 280 2211
rect 283 2211 289 2212
rect 283 2210 284 2211
rect 279 2208 284 2210
rect 279 2207 280 2208
rect 274 2206 280 2207
rect 283 2207 284 2208
rect 288 2207 289 2211
rect 283 2206 289 2207
rect 314 2211 320 2212
rect 314 2207 315 2211
rect 319 2210 320 2211
rect 323 2211 329 2212
rect 323 2210 324 2211
rect 319 2208 324 2210
rect 319 2207 320 2208
rect 314 2206 320 2207
rect 323 2207 324 2208
rect 328 2207 329 2211
rect 323 2206 329 2207
rect 350 2211 356 2212
rect 350 2207 351 2211
rect 355 2210 356 2211
rect 371 2211 377 2212
rect 371 2210 372 2211
rect 355 2208 372 2210
rect 355 2207 356 2208
rect 350 2206 356 2207
rect 371 2207 372 2208
rect 376 2207 377 2211
rect 371 2206 377 2207
rect 402 2211 408 2212
rect 402 2207 403 2211
rect 407 2210 408 2211
rect 427 2211 433 2212
rect 427 2210 428 2211
rect 407 2208 428 2210
rect 407 2207 408 2208
rect 402 2206 408 2207
rect 427 2207 428 2208
rect 432 2207 433 2211
rect 427 2206 433 2207
rect 462 2211 468 2212
rect 462 2207 463 2211
rect 467 2210 468 2211
rect 491 2211 497 2212
rect 491 2210 492 2211
rect 467 2208 492 2210
rect 467 2207 468 2208
rect 462 2206 468 2207
rect 491 2207 492 2208
rect 496 2207 497 2211
rect 491 2206 497 2207
rect 547 2211 553 2212
rect 547 2207 548 2211
rect 552 2210 553 2211
rect 570 2211 576 2212
rect 570 2210 571 2211
rect 552 2208 571 2210
rect 552 2207 553 2208
rect 547 2206 553 2207
rect 570 2207 571 2208
rect 575 2207 576 2211
rect 570 2206 576 2207
rect 578 2211 584 2212
rect 578 2207 579 2211
rect 583 2210 584 2211
rect 603 2211 609 2212
rect 603 2210 604 2211
rect 583 2208 604 2210
rect 583 2207 584 2208
rect 578 2206 584 2207
rect 603 2207 604 2208
rect 608 2207 609 2211
rect 603 2206 609 2207
rect 634 2211 640 2212
rect 634 2207 635 2211
rect 639 2210 640 2211
rect 659 2211 665 2212
rect 659 2210 660 2211
rect 639 2208 660 2210
rect 639 2207 640 2208
rect 634 2206 640 2207
rect 659 2207 660 2208
rect 664 2207 665 2211
rect 659 2206 665 2207
rect 715 2211 721 2212
rect 715 2207 716 2211
rect 720 2210 721 2211
rect 738 2211 744 2212
rect 738 2210 739 2211
rect 720 2208 739 2210
rect 720 2207 721 2208
rect 715 2206 721 2207
rect 738 2207 739 2208
rect 743 2207 744 2211
rect 738 2206 744 2207
rect 746 2211 752 2212
rect 746 2207 747 2211
rect 751 2210 752 2211
rect 779 2211 785 2212
rect 779 2210 780 2211
rect 751 2208 780 2210
rect 751 2207 752 2208
rect 746 2206 752 2207
rect 779 2207 780 2208
rect 784 2207 785 2211
rect 779 2206 785 2207
rect 843 2211 849 2212
rect 843 2207 844 2211
rect 848 2210 849 2211
rect 854 2211 860 2212
rect 854 2210 855 2211
rect 848 2208 855 2210
rect 848 2207 849 2208
rect 843 2206 849 2207
rect 854 2207 855 2208
rect 859 2207 860 2211
rect 854 2206 860 2207
rect 874 2211 880 2212
rect 874 2207 875 2211
rect 879 2210 880 2211
rect 907 2211 913 2212
rect 907 2210 908 2211
rect 879 2208 908 2210
rect 879 2207 880 2208
rect 874 2206 880 2207
rect 907 2207 908 2208
rect 912 2207 913 2211
rect 907 2206 913 2207
rect 246 2203 252 2204
rect 246 2199 247 2203
rect 251 2199 252 2203
rect 246 2198 252 2199
rect 286 2203 292 2204
rect 286 2199 287 2203
rect 291 2199 292 2203
rect 286 2198 292 2199
rect 326 2203 332 2204
rect 326 2199 327 2203
rect 331 2199 332 2203
rect 326 2198 332 2199
rect 374 2203 380 2204
rect 374 2199 375 2203
rect 379 2199 380 2203
rect 374 2198 380 2199
rect 430 2203 436 2204
rect 430 2199 431 2203
rect 435 2199 436 2203
rect 430 2198 436 2199
rect 494 2203 500 2204
rect 494 2199 495 2203
rect 499 2199 500 2203
rect 494 2198 500 2199
rect 550 2203 556 2204
rect 550 2199 551 2203
rect 555 2199 556 2203
rect 550 2198 556 2199
rect 606 2203 612 2204
rect 606 2199 607 2203
rect 611 2199 612 2203
rect 606 2198 612 2199
rect 662 2203 668 2204
rect 662 2199 663 2203
rect 667 2199 668 2203
rect 662 2198 668 2199
rect 718 2203 724 2204
rect 718 2199 719 2203
rect 723 2199 724 2203
rect 718 2198 724 2199
rect 782 2203 788 2204
rect 782 2199 783 2203
rect 787 2199 788 2203
rect 782 2198 788 2199
rect 846 2203 852 2204
rect 846 2199 847 2203
rect 851 2199 852 2203
rect 846 2198 852 2199
rect 910 2203 916 2204
rect 910 2199 911 2203
rect 915 2199 916 2203
rect 1327 2203 1336 2204
rect 910 2198 916 2199
rect 1278 2200 1284 2201
rect 1278 2196 1279 2200
rect 1283 2196 1284 2200
rect 1327 2199 1328 2203
rect 1335 2199 1336 2203
rect 1327 2198 1336 2199
rect 1367 2203 1376 2204
rect 1367 2199 1368 2203
rect 1375 2199 1376 2203
rect 1367 2198 1376 2199
rect 1407 2203 1413 2204
rect 1407 2199 1408 2203
rect 1412 2202 1413 2203
rect 1422 2203 1428 2204
rect 1422 2202 1423 2203
rect 1412 2200 1423 2202
rect 1412 2199 1413 2200
rect 1407 2198 1413 2199
rect 1422 2199 1423 2200
rect 1427 2199 1428 2203
rect 1422 2198 1428 2199
rect 1455 2203 1461 2204
rect 1455 2199 1456 2203
rect 1460 2202 1461 2203
rect 1486 2203 1492 2204
rect 1486 2202 1487 2203
rect 1460 2200 1487 2202
rect 1460 2199 1461 2200
rect 1455 2198 1461 2199
rect 1486 2199 1487 2200
rect 1491 2199 1492 2203
rect 1486 2198 1492 2199
rect 1519 2203 1525 2204
rect 1519 2199 1520 2203
rect 1524 2202 1525 2203
rect 1558 2203 1564 2204
rect 1558 2202 1559 2203
rect 1524 2200 1559 2202
rect 1524 2199 1525 2200
rect 1519 2198 1525 2199
rect 1558 2199 1559 2200
rect 1563 2199 1564 2203
rect 1558 2198 1564 2199
rect 1591 2203 1597 2204
rect 1591 2199 1592 2203
rect 1596 2202 1597 2203
rect 1622 2203 1628 2204
rect 1622 2202 1623 2203
rect 1596 2200 1623 2202
rect 1596 2199 1597 2200
rect 1591 2198 1597 2199
rect 1622 2199 1623 2200
rect 1627 2199 1628 2203
rect 1622 2198 1628 2199
rect 1654 2203 1660 2204
rect 1654 2199 1655 2203
rect 1659 2202 1660 2203
rect 1663 2203 1669 2204
rect 1663 2202 1664 2203
rect 1659 2200 1664 2202
rect 1659 2199 1660 2200
rect 1654 2198 1660 2199
rect 1663 2199 1664 2200
rect 1668 2199 1669 2203
rect 1663 2198 1669 2199
rect 1671 2203 1677 2204
rect 1671 2199 1672 2203
rect 1676 2202 1677 2203
rect 1735 2203 1741 2204
rect 1735 2202 1736 2203
rect 1676 2200 1736 2202
rect 1676 2199 1677 2200
rect 1671 2198 1677 2199
rect 1735 2199 1736 2200
rect 1740 2199 1741 2203
rect 1735 2198 1741 2199
rect 1807 2203 1813 2204
rect 1807 2199 1808 2203
rect 1812 2202 1813 2203
rect 1846 2203 1852 2204
rect 1846 2202 1847 2203
rect 1812 2200 1847 2202
rect 1812 2199 1813 2200
rect 1807 2198 1813 2199
rect 1846 2199 1847 2200
rect 1851 2199 1852 2203
rect 1846 2198 1852 2199
rect 1879 2203 1885 2204
rect 1879 2199 1880 2203
rect 1884 2202 1885 2203
rect 1926 2203 1932 2204
rect 1926 2202 1927 2203
rect 1884 2200 1927 2202
rect 1884 2199 1885 2200
rect 1879 2198 1885 2199
rect 1926 2199 1927 2200
rect 1931 2199 1932 2203
rect 1926 2198 1932 2199
rect 1959 2203 1965 2204
rect 1959 2199 1960 2203
rect 1964 2202 1965 2203
rect 2006 2203 2012 2204
rect 2006 2202 2007 2203
rect 1964 2200 2007 2202
rect 1964 2199 1965 2200
rect 1959 2198 1965 2199
rect 2006 2199 2007 2200
rect 2011 2199 2012 2203
rect 2006 2198 2012 2199
rect 2039 2203 2045 2204
rect 2039 2199 2040 2203
rect 2044 2202 2045 2203
rect 2086 2203 2092 2204
rect 2086 2202 2087 2203
rect 2044 2200 2087 2202
rect 2044 2199 2045 2200
rect 2039 2198 2045 2199
rect 2086 2199 2087 2200
rect 2091 2199 2092 2203
rect 2119 2203 2125 2204
rect 2119 2202 2120 2203
rect 2086 2198 2092 2199
rect 2096 2200 2120 2202
rect 1278 2195 1284 2196
rect 1822 2195 1828 2196
rect 1822 2191 1823 2195
rect 1827 2194 1828 2195
rect 2096 2194 2098 2200
rect 2119 2199 2120 2200
rect 2124 2199 2125 2203
rect 2119 2198 2125 2199
rect 2134 2203 2140 2204
rect 2134 2199 2135 2203
rect 2139 2202 2140 2203
rect 2207 2203 2213 2204
rect 2207 2202 2208 2203
rect 2139 2200 2208 2202
rect 2139 2199 2140 2200
rect 2134 2198 2140 2199
rect 2207 2199 2208 2200
rect 2212 2199 2213 2203
rect 2207 2198 2213 2199
rect 2215 2203 2221 2204
rect 2215 2199 2216 2203
rect 2220 2202 2221 2203
rect 2303 2203 2309 2204
rect 2303 2202 2304 2203
rect 2220 2200 2304 2202
rect 2220 2199 2221 2200
rect 2215 2198 2221 2199
rect 2303 2199 2304 2200
rect 2308 2199 2309 2203
rect 2303 2198 2309 2199
rect 2318 2203 2324 2204
rect 2318 2199 2319 2203
rect 2323 2202 2324 2203
rect 2383 2203 2389 2204
rect 2383 2202 2384 2203
rect 2323 2200 2384 2202
rect 2323 2199 2324 2200
rect 2318 2198 2324 2199
rect 2383 2199 2384 2200
rect 2388 2199 2389 2203
rect 2383 2198 2389 2199
rect 2406 2200 2412 2201
rect 2406 2196 2407 2200
rect 2411 2196 2412 2200
rect 2406 2195 2412 2196
rect 1827 2192 2098 2194
rect 1827 2191 1828 2192
rect 1822 2190 1828 2191
rect 591 2183 597 2184
rect 110 2180 116 2181
rect 110 2176 111 2180
rect 115 2176 116 2180
rect 591 2179 592 2183
rect 596 2182 597 2183
rect 738 2183 744 2184
rect 596 2180 646 2182
rect 596 2179 597 2180
rect 591 2178 597 2179
rect 110 2175 116 2176
rect 271 2175 280 2176
rect 271 2171 272 2175
rect 279 2171 280 2175
rect 271 2170 280 2171
rect 311 2175 320 2176
rect 311 2171 312 2175
rect 319 2171 320 2175
rect 311 2170 320 2171
rect 350 2175 357 2176
rect 350 2171 351 2175
rect 356 2171 357 2175
rect 350 2170 357 2171
rect 399 2175 408 2176
rect 399 2171 400 2175
rect 407 2171 408 2175
rect 399 2170 408 2171
rect 455 2175 464 2176
rect 455 2171 456 2175
rect 463 2171 464 2175
rect 519 2175 525 2176
rect 519 2174 520 2175
rect 455 2170 464 2171
rect 472 2172 520 2174
rect 390 2167 396 2168
rect 110 2163 116 2164
rect 110 2159 111 2163
rect 115 2159 116 2163
rect 390 2163 391 2167
rect 395 2166 396 2167
rect 472 2166 474 2172
rect 519 2171 520 2172
rect 524 2171 525 2175
rect 519 2170 525 2171
rect 575 2175 584 2176
rect 575 2171 576 2175
rect 583 2171 584 2175
rect 575 2170 584 2171
rect 631 2175 640 2176
rect 631 2171 632 2175
rect 639 2171 640 2175
rect 644 2174 646 2180
rect 738 2179 739 2183
rect 743 2182 744 2183
rect 743 2180 886 2182
rect 743 2179 744 2180
rect 738 2178 744 2179
rect 687 2175 693 2176
rect 687 2174 688 2175
rect 644 2172 688 2174
rect 631 2170 640 2171
rect 687 2171 688 2172
rect 692 2171 693 2175
rect 687 2170 693 2171
rect 743 2175 752 2176
rect 743 2171 744 2175
rect 751 2171 752 2175
rect 743 2170 752 2171
rect 806 2175 813 2176
rect 806 2171 807 2175
rect 812 2171 813 2175
rect 806 2170 813 2171
rect 871 2175 880 2176
rect 871 2171 872 2175
rect 879 2171 880 2175
rect 884 2174 886 2180
rect 1238 2180 1244 2181
rect 1238 2176 1239 2180
rect 1243 2176 1244 2180
rect 935 2175 941 2176
rect 1238 2175 1244 2176
rect 1302 2177 1308 2178
rect 935 2174 936 2175
rect 884 2172 936 2174
rect 871 2170 880 2171
rect 935 2171 936 2172
rect 940 2171 941 2175
rect 1302 2173 1303 2177
rect 1307 2173 1308 2177
rect 1302 2172 1308 2173
rect 1342 2177 1348 2178
rect 1342 2173 1343 2177
rect 1347 2173 1348 2177
rect 1342 2172 1348 2173
rect 1382 2177 1388 2178
rect 1382 2173 1383 2177
rect 1387 2173 1388 2177
rect 1382 2172 1388 2173
rect 1430 2177 1436 2178
rect 1430 2173 1431 2177
rect 1435 2173 1436 2177
rect 1430 2172 1436 2173
rect 1494 2177 1500 2178
rect 1494 2173 1495 2177
rect 1499 2173 1500 2177
rect 1494 2172 1500 2173
rect 1566 2177 1572 2178
rect 1566 2173 1567 2177
rect 1571 2173 1572 2177
rect 1566 2172 1572 2173
rect 1638 2177 1644 2178
rect 1638 2173 1639 2177
rect 1643 2173 1644 2177
rect 1638 2172 1644 2173
rect 1710 2177 1716 2178
rect 1710 2173 1711 2177
rect 1715 2173 1716 2177
rect 1710 2172 1716 2173
rect 1782 2177 1788 2178
rect 1782 2173 1783 2177
rect 1787 2173 1788 2177
rect 1782 2172 1788 2173
rect 1854 2177 1860 2178
rect 1854 2173 1855 2177
rect 1859 2173 1860 2177
rect 1854 2172 1860 2173
rect 1934 2177 1940 2178
rect 1934 2173 1935 2177
rect 1939 2173 1940 2177
rect 1934 2172 1940 2173
rect 2014 2177 2020 2178
rect 2014 2173 2015 2177
rect 2019 2173 2020 2177
rect 2014 2172 2020 2173
rect 2094 2177 2100 2178
rect 2094 2173 2095 2177
rect 2099 2173 2100 2177
rect 2094 2172 2100 2173
rect 2182 2177 2188 2178
rect 2182 2173 2183 2177
rect 2187 2173 2188 2177
rect 2182 2172 2188 2173
rect 2278 2177 2284 2178
rect 2278 2173 2279 2177
rect 2283 2173 2284 2177
rect 2278 2172 2284 2173
rect 2358 2177 2364 2178
rect 2358 2173 2359 2177
rect 2363 2173 2364 2177
rect 2358 2172 2364 2173
rect 935 2170 941 2171
rect 395 2164 474 2166
rect 1299 2167 1305 2168
rect 395 2163 396 2164
rect 390 2162 396 2163
rect 1238 2163 1244 2164
rect 110 2158 116 2159
rect 1238 2159 1239 2163
rect 1243 2159 1244 2163
rect 1299 2163 1300 2167
rect 1304 2166 1305 2167
rect 1314 2167 1320 2168
rect 1314 2166 1315 2167
rect 1304 2164 1315 2166
rect 1304 2163 1305 2164
rect 1299 2162 1305 2163
rect 1314 2163 1315 2164
rect 1319 2163 1320 2167
rect 1314 2162 1320 2163
rect 1330 2167 1336 2168
rect 1330 2163 1331 2167
rect 1335 2166 1336 2167
rect 1339 2167 1345 2168
rect 1339 2166 1340 2167
rect 1335 2164 1340 2166
rect 1335 2163 1336 2164
rect 1330 2162 1336 2163
rect 1339 2163 1340 2164
rect 1344 2163 1345 2167
rect 1339 2162 1345 2163
rect 1370 2167 1376 2168
rect 1370 2163 1371 2167
rect 1375 2166 1376 2167
rect 1379 2167 1385 2168
rect 1379 2166 1380 2167
rect 1375 2164 1380 2166
rect 1375 2163 1376 2164
rect 1370 2162 1376 2163
rect 1379 2163 1380 2164
rect 1384 2163 1385 2167
rect 1379 2162 1385 2163
rect 1422 2167 1433 2168
rect 1422 2163 1423 2167
rect 1427 2163 1428 2167
rect 1432 2163 1433 2167
rect 1422 2162 1433 2163
rect 1486 2167 1497 2168
rect 1486 2163 1487 2167
rect 1491 2163 1492 2167
rect 1496 2163 1497 2167
rect 1486 2162 1497 2163
rect 1558 2167 1569 2168
rect 1558 2163 1559 2167
rect 1563 2163 1564 2167
rect 1568 2163 1569 2167
rect 1558 2162 1569 2163
rect 1635 2167 1641 2168
rect 1635 2163 1636 2167
rect 1640 2166 1641 2167
rect 1671 2167 1677 2168
rect 1671 2166 1672 2167
rect 1640 2164 1672 2166
rect 1640 2163 1641 2164
rect 1635 2162 1641 2163
rect 1671 2163 1672 2164
rect 1676 2163 1677 2167
rect 1671 2162 1677 2163
rect 1707 2167 1713 2168
rect 1707 2163 1708 2167
rect 1712 2166 1713 2167
rect 1750 2167 1756 2168
rect 1750 2166 1751 2167
rect 1712 2164 1751 2166
rect 1712 2163 1713 2164
rect 1707 2162 1713 2163
rect 1750 2163 1751 2164
rect 1755 2163 1756 2167
rect 1750 2162 1756 2163
rect 1779 2167 1785 2168
rect 1779 2163 1780 2167
rect 1784 2166 1785 2167
rect 1790 2167 1796 2168
rect 1790 2166 1791 2167
rect 1784 2164 1791 2166
rect 1784 2163 1785 2164
rect 1779 2162 1785 2163
rect 1790 2163 1791 2164
rect 1795 2163 1796 2167
rect 1790 2162 1796 2163
rect 1846 2167 1857 2168
rect 1846 2163 1847 2167
rect 1851 2163 1852 2167
rect 1856 2163 1857 2167
rect 1846 2162 1857 2163
rect 1926 2167 1937 2168
rect 1926 2163 1927 2167
rect 1931 2163 1932 2167
rect 1936 2163 1937 2167
rect 1926 2162 1937 2163
rect 2006 2167 2017 2168
rect 2006 2163 2007 2167
rect 2011 2163 2012 2167
rect 2016 2163 2017 2167
rect 2006 2162 2017 2163
rect 2086 2167 2097 2168
rect 2086 2163 2087 2167
rect 2091 2163 2092 2167
rect 2096 2163 2097 2167
rect 2086 2162 2097 2163
rect 2179 2167 2185 2168
rect 2179 2163 2180 2167
rect 2184 2166 2185 2167
rect 2215 2167 2221 2168
rect 2215 2166 2216 2167
rect 2184 2164 2216 2166
rect 2184 2163 2185 2164
rect 2179 2162 2185 2163
rect 2215 2163 2216 2164
rect 2220 2163 2221 2167
rect 2215 2162 2221 2163
rect 2266 2167 2272 2168
rect 2266 2163 2267 2167
rect 2271 2166 2272 2167
rect 2275 2167 2281 2168
rect 2275 2166 2276 2167
rect 2271 2164 2276 2166
rect 2271 2163 2272 2164
rect 2266 2162 2272 2163
rect 2275 2163 2276 2164
rect 2280 2163 2281 2167
rect 2275 2162 2281 2163
rect 2355 2167 2361 2168
rect 2355 2163 2356 2167
rect 2360 2166 2361 2167
rect 2366 2167 2372 2168
rect 2366 2166 2367 2167
rect 2360 2164 2367 2166
rect 2360 2163 2361 2164
rect 2355 2162 2361 2163
rect 2366 2163 2367 2164
rect 2371 2163 2372 2167
rect 2366 2162 2372 2163
rect 1238 2158 1244 2159
rect 246 2156 252 2157
rect 246 2152 247 2156
rect 251 2152 252 2156
rect 246 2151 252 2152
rect 286 2156 292 2157
rect 286 2152 287 2156
rect 291 2152 292 2156
rect 286 2151 292 2152
rect 326 2156 332 2157
rect 326 2152 327 2156
rect 331 2152 332 2156
rect 326 2151 332 2152
rect 374 2156 380 2157
rect 374 2152 375 2156
rect 379 2152 380 2156
rect 374 2151 380 2152
rect 430 2156 436 2157
rect 430 2152 431 2156
rect 435 2152 436 2156
rect 430 2151 436 2152
rect 494 2156 500 2157
rect 494 2152 495 2156
rect 499 2152 500 2156
rect 494 2151 500 2152
rect 550 2156 556 2157
rect 550 2152 551 2156
rect 555 2152 556 2156
rect 550 2151 556 2152
rect 606 2156 612 2157
rect 606 2152 607 2156
rect 611 2152 612 2156
rect 606 2151 612 2152
rect 662 2156 668 2157
rect 662 2152 663 2156
rect 667 2152 668 2156
rect 662 2151 668 2152
rect 718 2156 724 2157
rect 718 2152 719 2156
rect 723 2152 724 2156
rect 718 2151 724 2152
rect 782 2156 788 2157
rect 782 2152 783 2156
rect 787 2152 788 2156
rect 782 2151 788 2152
rect 846 2156 852 2157
rect 846 2152 847 2156
rect 851 2152 852 2156
rect 846 2151 852 2152
rect 910 2156 916 2157
rect 910 2152 911 2156
rect 915 2152 916 2156
rect 910 2151 916 2152
rect 1299 2155 1305 2156
rect 1299 2151 1300 2155
rect 1304 2154 1305 2155
rect 1322 2155 1328 2156
rect 1322 2154 1323 2155
rect 1304 2152 1323 2154
rect 1304 2151 1305 2152
rect 1299 2150 1305 2151
rect 1322 2151 1323 2152
rect 1327 2151 1328 2155
rect 1322 2150 1328 2151
rect 1330 2155 1336 2156
rect 1330 2151 1331 2155
rect 1335 2154 1336 2155
rect 1347 2155 1353 2156
rect 1347 2154 1348 2155
rect 1335 2152 1348 2154
rect 1335 2151 1336 2152
rect 1330 2150 1336 2151
rect 1347 2151 1348 2152
rect 1352 2151 1353 2155
rect 1347 2150 1353 2151
rect 1435 2155 1441 2156
rect 1435 2151 1436 2155
rect 1440 2154 1441 2155
rect 1522 2155 1528 2156
rect 1522 2154 1523 2155
rect 1440 2152 1523 2154
rect 1440 2151 1441 2152
rect 1435 2150 1441 2151
rect 1522 2151 1523 2152
rect 1527 2151 1528 2155
rect 1522 2150 1528 2151
rect 1531 2155 1537 2156
rect 1531 2151 1532 2155
rect 1536 2154 1537 2155
rect 1614 2155 1620 2156
rect 1614 2154 1615 2155
rect 1536 2152 1615 2154
rect 1536 2151 1537 2152
rect 1531 2150 1537 2151
rect 1614 2151 1615 2152
rect 1619 2151 1620 2155
rect 1614 2150 1620 2151
rect 1622 2155 1633 2156
rect 1622 2151 1623 2155
rect 1627 2151 1628 2155
rect 1632 2151 1633 2155
rect 1622 2150 1633 2151
rect 1723 2155 1729 2156
rect 1723 2151 1724 2155
rect 1728 2154 1729 2155
rect 1774 2155 1780 2156
rect 1774 2154 1775 2155
rect 1728 2152 1775 2154
rect 1728 2151 1729 2152
rect 1723 2150 1729 2151
rect 1774 2151 1775 2152
rect 1779 2151 1780 2155
rect 1774 2150 1780 2151
rect 1811 2155 1817 2156
rect 1811 2151 1812 2155
rect 1816 2154 1817 2155
rect 1822 2155 1828 2156
rect 1822 2154 1823 2155
rect 1816 2152 1823 2154
rect 1816 2151 1817 2152
rect 1811 2150 1817 2151
rect 1822 2151 1823 2152
rect 1827 2151 1828 2155
rect 1822 2150 1828 2151
rect 1842 2155 1848 2156
rect 1842 2151 1843 2155
rect 1847 2154 1848 2155
rect 1891 2155 1897 2156
rect 1891 2154 1892 2155
rect 1847 2152 1892 2154
rect 1847 2151 1848 2152
rect 1842 2150 1848 2151
rect 1891 2151 1892 2152
rect 1896 2151 1897 2155
rect 1891 2150 1897 2151
rect 1927 2155 1933 2156
rect 1927 2151 1928 2155
rect 1932 2154 1933 2155
rect 1971 2155 1977 2156
rect 1971 2154 1972 2155
rect 1932 2152 1972 2154
rect 1932 2151 1933 2152
rect 1927 2150 1933 2151
rect 1971 2151 1972 2152
rect 1976 2151 1977 2155
rect 1971 2150 1977 2151
rect 1998 2155 2004 2156
rect 1998 2151 1999 2155
rect 2003 2154 2004 2155
rect 2043 2155 2049 2156
rect 2043 2154 2044 2155
rect 2003 2152 2044 2154
rect 2003 2151 2004 2152
rect 1998 2150 2004 2151
rect 2043 2151 2044 2152
rect 2048 2151 2049 2155
rect 2043 2150 2049 2151
rect 2054 2155 2060 2156
rect 2054 2151 2055 2155
rect 2059 2154 2060 2155
rect 2107 2155 2113 2156
rect 2107 2154 2108 2155
rect 2059 2152 2108 2154
rect 2059 2151 2060 2152
rect 2054 2150 2060 2151
rect 2107 2151 2108 2152
rect 2112 2151 2113 2155
rect 2107 2150 2113 2151
rect 2138 2155 2144 2156
rect 2138 2151 2139 2155
rect 2143 2154 2144 2155
rect 2171 2155 2177 2156
rect 2171 2154 2172 2155
rect 2143 2152 2172 2154
rect 2143 2151 2144 2152
rect 2138 2150 2144 2151
rect 2171 2151 2172 2152
rect 2176 2151 2177 2155
rect 2171 2150 2177 2151
rect 2202 2155 2208 2156
rect 2202 2151 2203 2155
rect 2207 2154 2208 2155
rect 2235 2155 2241 2156
rect 2235 2154 2236 2155
rect 2207 2152 2236 2154
rect 2207 2151 2208 2152
rect 2202 2150 2208 2151
rect 2235 2151 2236 2152
rect 2240 2151 2241 2155
rect 2235 2150 2241 2151
rect 2307 2155 2313 2156
rect 2307 2151 2308 2155
rect 2312 2154 2313 2155
rect 2318 2155 2324 2156
rect 2318 2154 2319 2155
rect 2312 2152 2319 2154
rect 2312 2151 2313 2152
rect 2307 2150 2313 2151
rect 2318 2151 2319 2152
rect 2323 2151 2324 2155
rect 2318 2150 2324 2151
rect 2338 2155 2344 2156
rect 2338 2151 2339 2155
rect 2343 2154 2344 2155
rect 2355 2155 2361 2156
rect 2355 2154 2356 2155
rect 2343 2152 2356 2154
rect 2343 2151 2344 2152
rect 2338 2150 2344 2151
rect 2355 2151 2356 2152
rect 2360 2151 2361 2155
rect 2355 2150 2361 2151
rect 1302 2147 1308 2148
rect 1302 2143 1303 2147
rect 1307 2143 1308 2147
rect 1302 2142 1308 2143
rect 1350 2147 1356 2148
rect 1350 2143 1351 2147
rect 1355 2143 1356 2147
rect 1350 2142 1356 2143
rect 1438 2147 1444 2148
rect 1438 2143 1439 2147
rect 1443 2143 1444 2147
rect 1438 2142 1444 2143
rect 1534 2147 1540 2148
rect 1534 2143 1535 2147
rect 1539 2143 1540 2147
rect 1534 2142 1540 2143
rect 1630 2147 1636 2148
rect 1630 2143 1631 2147
rect 1635 2143 1636 2147
rect 1630 2142 1636 2143
rect 1726 2147 1732 2148
rect 1726 2143 1727 2147
rect 1731 2143 1732 2147
rect 1726 2142 1732 2143
rect 1814 2147 1820 2148
rect 1814 2143 1815 2147
rect 1819 2143 1820 2147
rect 1814 2142 1820 2143
rect 1894 2147 1900 2148
rect 1894 2143 1895 2147
rect 1899 2143 1900 2147
rect 1894 2142 1900 2143
rect 1974 2147 1980 2148
rect 1974 2143 1975 2147
rect 1979 2143 1980 2147
rect 1974 2142 1980 2143
rect 2046 2147 2052 2148
rect 2046 2143 2047 2147
rect 2051 2143 2052 2147
rect 2046 2142 2052 2143
rect 2110 2147 2116 2148
rect 2110 2143 2111 2147
rect 2115 2143 2116 2147
rect 2110 2142 2116 2143
rect 2174 2147 2180 2148
rect 2174 2143 2175 2147
rect 2179 2143 2180 2147
rect 2174 2142 2180 2143
rect 2238 2147 2244 2148
rect 2238 2143 2239 2147
rect 2243 2143 2244 2147
rect 2238 2142 2244 2143
rect 2310 2147 2316 2148
rect 2310 2143 2311 2147
rect 2315 2143 2316 2147
rect 2310 2142 2316 2143
rect 2358 2147 2364 2148
rect 2358 2143 2359 2147
rect 2363 2143 2364 2147
rect 2358 2142 2364 2143
rect 382 2136 388 2137
rect 382 2132 383 2136
rect 387 2132 388 2136
rect 382 2131 388 2132
rect 422 2136 428 2137
rect 422 2132 423 2136
rect 427 2132 428 2136
rect 422 2131 428 2132
rect 462 2136 468 2137
rect 462 2132 463 2136
rect 467 2132 468 2136
rect 462 2131 468 2132
rect 502 2136 508 2137
rect 502 2132 503 2136
rect 507 2132 508 2136
rect 502 2131 508 2132
rect 550 2136 556 2137
rect 550 2132 551 2136
rect 555 2132 556 2136
rect 550 2131 556 2132
rect 606 2136 612 2137
rect 606 2132 607 2136
rect 611 2132 612 2136
rect 606 2131 612 2132
rect 662 2136 668 2137
rect 662 2132 663 2136
rect 667 2132 668 2136
rect 662 2131 668 2132
rect 726 2136 732 2137
rect 726 2132 727 2136
rect 731 2132 732 2136
rect 726 2131 732 2132
rect 790 2136 796 2137
rect 790 2132 791 2136
rect 795 2132 796 2136
rect 790 2131 796 2132
rect 854 2136 860 2137
rect 854 2132 855 2136
rect 859 2132 860 2136
rect 854 2131 860 2132
rect 910 2136 916 2137
rect 910 2132 911 2136
rect 915 2132 916 2136
rect 910 2131 916 2132
rect 966 2136 972 2137
rect 966 2132 967 2136
rect 971 2132 972 2136
rect 966 2131 972 2132
rect 1022 2136 1028 2137
rect 1022 2132 1023 2136
rect 1027 2132 1028 2136
rect 1022 2131 1028 2132
rect 1078 2136 1084 2137
rect 1078 2132 1079 2136
rect 1083 2132 1084 2136
rect 1078 2131 1084 2132
rect 1142 2136 1148 2137
rect 1142 2132 1143 2136
rect 1147 2132 1148 2136
rect 1142 2131 1148 2132
rect 110 2129 116 2130
rect 110 2125 111 2129
rect 115 2125 116 2129
rect 110 2124 116 2125
rect 1238 2129 1244 2130
rect 1238 2125 1239 2129
rect 1243 2125 1244 2129
rect 1314 2127 1320 2128
rect 1238 2124 1244 2125
rect 1278 2124 1284 2125
rect 1278 2120 1279 2124
rect 1283 2120 1284 2124
rect 1314 2123 1315 2127
rect 1319 2126 1320 2127
rect 1319 2124 1342 2126
rect 1319 2123 1320 2124
rect 1314 2122 1320 2123
rect 1278 2119 1284 2120
rect 1327 2119 1336 2120
rect 407 2115 416 2116
rect 110 2112 116 2113
rect 110 2108 111 2112
rect 115 2108 116 2112
rect 407 2111 408 2115
rect 415 2111 416 2115
rect 407 2110 416 2111
rect 447 2115 456 2116
rect 447 2111 448 2115
rect 455 2111 456 2115
rect 447 2110 456 2111
rect 487 2115 496 2116
rect 487 2111 488 2115
rect 495 2111 496 2115
rect 527 2115 533 2116
rect 527 2114 528 2115
rect 487 2110 496 2111
rect 500 2112 528 2114
rect 110 2107 116 2108
rect 398 2107 404 2108
rect 398 2103 399 2107
rect 403 2106 404 2107
rect 500 2106 502 2112
rect 527 2111 528 2112
rect 532 2111 533 2115
rect 527 2110 533 2111
rect 570 2115 581 2116
rect 570 2111 571 2115
rect 575 2111 576 2115
rect 580 2111 581 2115
rect 570 2110 581 2111
rect 583 2115 589 2116
rect 583 2111 584 2115
rect 588 2114 589 2115
rect 631 2115 637 2116
rect 631 2114 632 2115
rect 588 2112 632 2114
rect 588 2111 589 2112
rect 583 2110 589 2111
rect 631 2111 632 2112
rect 636 2111 637 2115
rect 631 2110 637 2111
rect 639 2115 645 2116
rect 639 2111 640 2115
rect 644 2114 645 2115
rect 687 2115 693 2116
rect 687 2114 688 2115
rect 644 2112 688 2114
rect 644 2111 645 2112
rect 639 2110 645 2111
rect 687 2111 688 2112
rect 692 2111 693 2115
rect 687 2110 693 2111
rect 750 2115 757 2116
rect 750 2111 751 2115
rect 756 2111 757 2115
rect 750 2110 757 2111
rect 770 2115 776 2116
rect 770 2111 771 2115
rect 775 2114 776 2115
rect 815 2115 821 2116
rect 815 2114 816 2115
rect 775 2112 816 2114
rect 775 2111 776 2112
rect 770 2110 776 2111
rect 815 2111 816 2112
rect 820 2111 821 2115
rect 815 2110 821 2111
rect 879 2115 885 2116
rect 879 2111 880 2115
rect 884 2114 885 2115
rect 894 2115 900 2116
rect 894 2114 895 2115
rect 884 2112 895 2114
rect 884 2111 885 2112
rect 879 2110 885 2111
rect 894 2111 895 2112
rect 899 2111 900 2115
rect 894 2110 900 2111
rect 935 2115 941 2116
rect 935 2111 936 2115
rect 940 2114 941 2115
rect 950 2115 956 2116
rect 950 2114 951 2115
rect 940 2112 951 2114
rect 940 2111 941 2112
rect 935 2110 941 2111
rect 950 2111 951 2112
rect 955 2111 956 2115
rect 950 2110 956 2111
rect 991 2115 997 2116
rect 991 2111 992 2115
rect 996 2114 997 2115
rect 1006 2115 1012 2116
rect 1006 2114 1007 2115
rect 996 2112 1007 2114
rect 996 2111 997 2112
rect 991 2110 997 2111
rect 1006 2111 1007 2112
rect 1011 2111 1012 2115
rect 1006 2110 1012 2111
rect 1047 2115 1053 2116
rect 1047 2111 1048 2115
rect 1052 2114 1053 2115
rect 1062 2115 1068 2116
rect 1062 2114 1063 2115
rect 1052 2112 1063 2114
rect 1052 2111 1053 2112
rect 1047 2110 1053 2111
rect 1062 2111 1063 2112
rect 1067 2111 1068 2115
rect 1062 2110 1068 2111
rect 1103 2115 1109 2116
rect 1103 2111 1104 2115
rect 1108 2114 1109 2115
rect 1134 2115 1140 2116
rect 1134 2114 1135 2115
rect 1108 2112 1135 2114
rect 1108 2111 1109 2112
rect 1103 2110 1109 2111
rect 1134 2111 1135 2112
rect 1139 2111 1140 2115
rect 1134 2110 1140 2111
rect 1150 2115 1156 2116
rect 1150 2111 1151 2115
rect 1155 2114 1156 2115
rect 1167 2115 1173 2116
rect 1167 2114 1168 2115
rect 1155 2112 1168 2114
rect 1155 2111 1156 2112
rect 1150 2110 1156 2111
rect 1167 2111 1168 2112
rect 1172 2111 1173 2115
rect 1327 2115 1328 2119
rect 1335 2115 1336 2119
rect 1340 2118 1342 2124
rect 2406 2124 2412 2125
rect 2406 2120 2407 2124
rect 2411 2120 2412 2124
rect 1375 2119 1381 2120
rect 1375 2118 1376 2119
rect 1340 2116 1376 2118
rect 1327 2114 1336 2115
rect 1375 2115 1376 2116
rect 1380 2115 1381 2119
rect 1375 2114 1381 2115
rect 1406 2119 1412 2120
rect 1406 2115 1407 2119
rect 1411 2118 1412 2119
rect 1463 2119 1469 2120
rect 1463 2118 1464 2119
rect 1411 2116 1464 2118
rect 1411 2115 1412 2116
rect 1406 2114 1412 2115
rect 1463 2115 1464 2116
rect 1468 2115 1469 2119
rect 1463 2114 1469 2115
rect 1522 2119 1528 2120
rect 1522 2115 1523 2119
rect 1527 2118 1528 2119
rect 1559 2119 1565 2120
rect 1559 2118 1560 2119
rect 1527 2116 1560 2118
rect 1527 2115 1528 2116
rect 1522 2114 1528 2115
rect 1559 2115 1560 2116
rect 1564 2115 1565 2119
rect 1559 2114 1565 2115
rect 1614 2119 1620 2120
rect 1614 2115 1615 2119
rect 1619 2118 1620 2119
rect 1655 2119 1661 2120
rect 1655 2118 1656 2119
rect 1619 2116 1656 2118
rect 1619 2115 1620 2116
rect 1614 2114 1620 2115
rect 1655 2115 1656 2116
rect 1660 2115 1661 2119
rect 1655 2114 1661 2115
rect 1750 2119 1757 2120
rect 1750 2115 1751 2119
rect 1756 2115 1757 2119
rect 1750 2114 1757 2115
rect 1839 2119 1848 2120
rect 1839 2115 1840 2119
rect 1847 2115 1848 2119
rect 1839 2114 1848 2115
rect 1919 2119 1925 2120
rect 1919 2115 1920 2119
rect 1924 2118 1925 2119
rect 1927 2119 1933 2120
rect 1927 2118 1928 2119
rect 1924 2116 1928 2118
rect 1924 2115 1925 2116
rect 1919 2114 1925 2115
rect 1927 2115 1928 2116
rect 1932 2115 1933 2119
rect 1927 2114 1933 2115
rect 1998 2119 2005 2120
rect 1998 2115 1999 2119
rect 2004 2115 2005 2119
rect 2071 2119 2077 2120
rect 2071 2118 2072 2119
rect 1998 2114 2005 2115
rect 2036 2116 2072 2118
rect 1167 2110 1173 2111
rect 1238 2112 1244 2113
rect 1238 2108 1239 2112
rect 1243 2108 1244 2112
rect 1942 2111 1948 2112
rect 1238 2107 1244 2108
rect 1278 2107 1284 2108
rect 403 2104 502 2106
rect 403 2103 404 2104
rect 398 2102 404 2103
rect 1278 2103 1279 2107
rect 1283 2103 1284 2107
rect 1942 2107 1943 2111
rect 1947 2110 1948 2111
rect 2036 2110 2038 2116
rect 2071 2115 2072 2116
rect 2076 2115 2077 2119
rect 2071 2114 2077 2115
rect 2135 2119 2144 2120
rect 2135 2115 2136 2119
rect 2143 2115 2144 2119
rect 2135 2114 2144 2115
rect 2199 2119 2208 2120
rect 2199 2115 2200 2119
rect 2207 2115 2208 2119
rect 2199 2114 2208 2115
rect 2263 2119 2272 2120
rect 2263 2115 2264 2119
rect 2271 2115 2272 2119
rect 2263 2114 2272 2115
rect 2335 2119 2344 2120
rect 2335 2115 2336 2119
rect 2343 2115 2344 2119
rect 2335 2114 2344 2115
rect 2366 2119 2372 2120
rect 2366 2115 2367 2119
rect 2371 2118 2372 2119
rect 2383 2119 2389 2120
rect 2406 2119 2412 2120
rect 2383 2118 2384 2119
rect 2371 2116 2384 2118
rect 2371 2115 2372 2116
rect 2366 2114 2372 2115
rect 2383 2115 2384 2116
rect 2388 2115 2389 2119
rect 2383 2114 2389 2115
rect 1947 2108 2038 2110
rect 1947 2107 1948 2108
rect 1942 2106 1948 2107
rect 2406 2107 2412 2108
rect 1278 2102 1284 2103
rect 2406 2103 2407 2107
rect 2411 2103 2412 2107
rect 2406 2102 2412 2103
rect 1302 2100 1308 2101
rect 1302 2096 1303 2100
rect 1307 2096 1308 2100
rect 1302 2095 1308 2096
rect 1350 2100 1356 2101
rect 1350 2096 1351 2100
rect 1355 2096 1356 2100
rect 1350 2095 1356 2096
rect 1438 2100 1444 2101
rect 1438 2096 1439 2100
rect 1443 2096 1444 2100
rect 1438 2095 1444 2096
rect 1534 2100 1540 2101
rect 1534 2096 1535 2100
rect 1539 2096 1540 2100
rect 1534 2095 1540 2096
rect 1630 2100 1636 2101
rect 1630 2096 1631 2100
rect 1635 2096 1636 2100
rect 1630 2095 1636 2096
rect 1726 2100 1732 2101
rect 1726 2096 1727 2100
rect 1731 2096 1732 2100
rect 1726 2095 1732 2096
rect 1814 2100 1820 2101
rect 1814 2096 1815 2100
rect 1819 2096 1820 2100
rect 1814 2095 1820 2096
rect 1894 2100 1900 2101
rect 1894 2096 1895 2100
rect 1899 2096 1900 2100
rect 1894 2095 1900 2096
rect 1974 2100 1980 2101
rect 1974 2096 1975 2100
rect 1979 2096 1980 2100
rect 1974 2095 1980 2096
rect 2046 2100 2052 2101
rect 2046 2096 2047 2100
rect 2051 2096 2052 2100
rect 2046 2095 2052 2096
rect 2110 2100 2116 2101
rect 2110 2096 2111 2100
rect 2115 2096 2116 2100
rect 2110 2095 2116 2096
rect 2174 2100 2180 2101
rect 2174 2096 2175 2100
rect 2179 2096 2180 2100
rect 2174 2095 2180 2096
rect 2238 2100 2244 2101
rect 2238 2096 2239 2100
rect 2243 2096 2244 2100
rect 2238 2095 2244 2096
rect 2310 2100 2316 2101
rect 2310 2096 2311 2100
rect 2315 2096 2316 2100
rect 2310 2095 2316 2096
rect 2358 2100 2364 2101
rect 2358 2096 2359 2100
rect 2363 2096 2364 2100
rect 2358 2095 2364 2096
rect 382 2089 388 2090
rect 382 2085 383 2089
rect 387 2085 388 2089
rect 382 2084 388 2085
rect 422 2089 428 2090
rect 422 2085 423 2089
rect 427 2085 428 2089
rect 422 2084 428 2085
rect 462 2089 468 2090
rect 462 2085 463 2089
rect 467 2085 468 2089
rect 462 2084 468 2085
rect 502 2089 508 2090
rect 502 2085 503 2089
rect 507 2085 508 2089
rect 502 2084 508 2085
rect 550 2089 556 2090
rect 550 2085 551 2089
rect 555 2085 556 2089
rect 550 2084 556 2085
rect 606 2089 612 2090
rect 606 2085 607 2089
rect 611 2085 612 2089
rect 606 2084 612 2085
rect 662 2089 668 2090
rect 662 2085 663 2089
rect 667 2085 668 2089
rect 662 2084 668 2085
rect 726 2089 732 2090
rect 726 2085 727 2089
rect 731 2085 732 2089
rect 726 2084 732 2085
rect 790 2089 796 2090
rect 790 2085 791 2089
rect 795 2085 796 2089
rect 790 2084 796 2085
rect 854 2089 860 2090
rect 854 2085 855 2089
rect 859 2085 860 2089
rect 854 2084 860 2085
rect 910 2089 916 2090
rect 910 2085 911 2089
rect 915 2085 916 2089
rect 910 2084 916 2085
rect 966 2089 972 2090
rect 966 2085 967 2089
rect 971 2085 972 2089
rect 966 2084 972 2085
rect 1022 2089 1028 2090
rect 1022 2085 1023 2089
rect 1027 2085 1028 2089
rect 1022 2084 1028 2085
rect 1078 2089 1084 2090
rect 1078 2085 1079 2089
rect 1083 2085 1084 2089
rect 1078 2084 1084 2085
rect 1142 2089 1148 2090
rect 1142 2085 1143 2089
rect 1147 2085 1148 2089
rect 1142 2084 1148 2085
rect 1302 2084 1308 2085
rect 1302 2080 1303 2084
rect 1307 2080 1308 2084
rect 379 2079 385 2080
rect 379 2075 380 2079
rect 384 2078 385 2079
rect 390 2079 396 2080
rect 390 2078 391 2079
rect 384 2076 391 2078
rect 384 2075 385 2076
rect 379 2074 385 2075
rect 390 2075 391 2076
rect 395 2075 396 2079
rect 390 2074 396 2075
rect 410 2079 416 2080
rect 410 2075 411 2079
rect 415 2078 416 2079
rect 419 2079 425 2080
rect 419 2078 420 2079
rect 415 2076 420 2078
rect 415 2075 416 2076
rect 410 2074 416 2075
rect 419 2075 420 2076
rect 424 2075 425 2079
rect 419 2074 425 2075
rect 450 2079 456 2080
rect 450 2075 451 2079
rect 455 2078 456 2079
rect 459 2079 465 2080
rect 459 2078 460 2079
rect 455 2076 460 2078
rect 455 2075 456 2076
rect 450 2074 456 2075
rect 459 2075 460 2076
rect 464 2075 465 2079
rect 459 2074 465 2075
rect 490 2079 496 2080
rect 490 2075 491 2079
rect 495 2078 496 2079
rect 499 2079 505 2080
rect 499 2078 500 2079
rect 495 2076 500 2078
rect 495 2075 496 2076
rect 490 2074 496 2075
rect 499 2075 500 2076
rect 504 2075 505 2079
rect 499 2074 505 2075
rect 547 2079 553 2080
rect 547 2075 548 2079
rect 552 2078 553 2079
rect 583 2079 589 2080
rect 583 2078 584 2079
rect 552 2076 584 2078
rect 552 2075 553 2076
rect 547 2074 553 2075
rect 583 2075 584 2076
rect 588 2075 589 2079
rect 583 2074 589 2075
rect 603 2079 609 2080
rect 603 2075 604 2079
rect 608 2078 609 2079
rect 639 2079 645 2080
rect 639 2078 640 2079
rect 608 2076 640 2078
rect 608 2075 609 2076
rect 603 2074 609 2075
rect 639 2075 640 2076
rect 644 2075 645 2079
rect 639 2074 645 2075
rect 654 2079 665 2080
rect 654 2075 655 2079
rect 659 2075 660 2079
rect 664 2075 665 2079
rect 654 2074 665 2075
rect 723 2079 729 2080
rect 723 2075 724 2079
rect 728 2078 729 2079
rect 770 2079 776 2080
rect 770 2078 771 2079
rect 728 2076 771 2078
rect 728 2075 729 2076
rect 723 2074 729 2075
rect 770 2075 771 2076
rect 775 2075 776 2079
rect 770 2074 776 2075
rect 787 2079 793 2080
rect 787 2075 788 2079
rect 792 2078 793 2079
rect 806 2079 812 2080
rect 806 2078 807 2079
rect 792 2076 807 2078
rect 792 2075 793 2076
rect 787 2074 793 2075
rect 806 2075 807 2076
rect 811 2075 812 2079
rect 806 2074 812 2075
rect 851 2079 857 2080
rect 851 2075 852 2079
rect 856 2078 857 2079
rect 886 2079 892 2080
rect 886 2078 887 2079
rect 856 2076 887 2078
rect 856 2075 857 2076
rect 851 2074 857 2075
rect 886 2075 887 2076
rect 891 2075 892 2079
rect 886 2074 892 2075
rect 894 2079 900 2080
rect 894 2075 895 2079
rect 899 2078 900 2079
rect 907 2079 913 2080
rect 907 2078 908 2079
rect 899 2076 908 2078
rect 899 2075 900 2076
rect 894 2074 900 2075
rect 907 2075 908 2076
rect 912 2075 913 2079
rect 907 2074 913 2075
rect 950 2079 956 2080
rect 950 2075 951 2079
rect 955 2078 956 2079
rect 963 2079 969 2080
rect 963 2078 964 2079
rect 955 2076 964 2078
rect 955 2075 956 2076
rect 950 2074 956 2075
rect 963 2075 964 2076
rect 968 2075 969 2079
rect 963 2074 969 2075
rect 1006 2079 1012 2080
rect 1006 2075 1007 2079
rect 1011 2078 1012 2079
rect 1019 2079 1025 2080
rect 1019 2078 1020 2079
rect 1011 2076 1020 2078
rect 1011 2075 1012 2076
rect 1006 2074 1012 2075
rect 1019 2075 1020 2076
rect 1024 2075 1025 2079
rect 1019 2074 1025 2075
rect 1062 2079 1068 2080
rect 1062 2075 1063 2079
rect 1067 2078 1068 2079
rect 1075 2079 1081 2080
rect 1075 2078 1076 2079
rect 1067 2076 1076 2078
rect 1067 2075 1068 2076
rect 1062 2074 1068 2075
rect 1075 2075 1076 2076
rect 1080 2075 1081 2079
rect 1075 2074 1081 2075
rect 1134 2079 1145 2080
rect 1302 2079 1308 2080
rect 1342 2084 1348 2085
rect 1342 2080 1343 2084
rect 1347 2080 1348 2084
rect 1342 2079 1348 2080
rect 1398 2084 1404 2085
rect 1398 2080 1399 2084
rect 1403 2080 1404 2084
rect 1398 2079 1404 2080
rect 1478 2084 1484 2085
rect 1478 2080 1479 2084
rect 1483 2080 1484 2084
rect 1478 2079 1484 2080
rect 1566 2084 1572 2085
rect 1566 2080 1567 2084
rect 1571 2080 1572 2084
rect 1566 2079 1572 2080
rect 1662 2084 1668 2085
rect 1662 2080 1663 2084
rect 1667 2080 1668 2084
rect 1662 2079 1668 2080
rect 1758 2084 1764 2085
rect 1758 2080 1759 2084
rect 1763 2080 1764 2084
rect 1758 2079 1764 2080
rect 1846 2084 1852 2085
rect 1846 2080 1847 2084
rect 1851 2080 1852 2084
rect 1846 2079 1852 2080
rect 1934 2084 1940 2085
rect 1934 2080 1935 2084
rect 1939 2080 1940 2084
rect 1934 2079 1940 2080
rect 2014 2084 2020 2085
rect 2014 2080 2015 2084
rect 2019 2080 2020 2084
rect 2014 2079 2020 2080
rect 2094 2084 2100 2085
rect 2094 2080 2095 2084
rect 2099 2080 2100 2084
rect 2094 2079 2100 2080
rect 2166 2084 2172 2085
rect 2166 2080 2167 2084
rect 2171 2080 2172 2084
rect 2166 2079 2172 2080
rect 2238 2084 2244 2085
rect 2238 2080 2239 2084
rect 2243 2080 2244 2084
rect 2238 2079 2244 2080
rect 2310 2084 2316 2085
rect 2310 2080 2311 2084
rect 2315 2080 2316 2084
rect 2310 2079 2316 2080
rect 2358 2084 2364 2085
rect 2358 2080 2359 2084
rect 2363 2080 2364 2084
rect 2358 2079 2364 2080
rect 1134 2075 1135 2079
rect 1139 2075 1140 2079
rect 1144 2075 1145 2079
rect 1134 2074 1145 2075
rect 1278 2077 1284 2078
rect 1278 2073 1279 2077
rect 1283 2073 1284 2077
rect 1278 2072 1284 2073
rect 2406 2077 2412 2078
rect 2406 2073 2407 2077
rect 2411 2073 2412 2077
rect 2406 2072 2412 2073
rect 379 2067 385 2068
rect 379 2063 380 2067
rect 384 2066 385 2067
rect 398 2067 404 2068
rect 398 2066 399 2067
rect 384 2064 399 2066
rect 384 2063 385 2064
rect 379 2062 385 2063
rect 398 2063 399 2064
rect 403 2063 404 2067
rect 398 2062 404 2063
rect 410 2067 416 2068
rect 410 2063 411 2067
rect 415 2066 416 2067
rect 419 2067 425 2068
rect 419 2066 420 2067
rect 415 2064 420 2066
rect 415 2063 416 2064
rect 410 2062 416 2063
rect 419 2063 420 2064
rect 424 2063 425 2067
rect 419 2062 425 2063
rect 446 2067 452 2068
rect 446 2063 447 2067
rect 451 2066 452 2067
rect 459 2067 465 2068
rect 459 2066 460 2067
rect 451 2064 460 2066
rect 451 2063 452 2064
rect 446 2062 452 2063
rect 459 2063 460 2064
rect 464 2063 465 2067
rect 459 2062 465 2063
rect 490 2067 496 2068
rect 490 2063 491 2067
rect 495 2066 496 2067
rect 499 2067 505 2068
rect 499 2066 500 2067
rect 495 2064 500 2066
rect 495 2063 496 2064
rect 490 2062 496 2063
rect 499 2063 500 2064
rect 504 2063 505 2067
rect 499 2062 505 2063
rect 526 2067 532 2068
rect 526 2063 527 2067
rect 531 2066 532 2067
rect 539 2067 545 2068
rect 539 2066 540 2067
rect 531 2064 540 2066
rect 531 2063 532 2064
rect 526 2062 532 2063
rect 539 2063 540 2064
rect 544 2063 545 2067
rect 539 2062 545 2063
rect 570 2067 576 2068
rect 570 2063 571 2067
rect 575 2066 576 2067
rect 579 2067 585 2068
rect 579 2066 580 2067
rect 575 2064 580 2066
rect 575 2063 576 2064
rect 570 2062 576 2063
rect 579 2063 580 2064
rect 584 2063 585 2067
rect 579 2062 585 2063
rect 614 2067 620 2068
rect 614 2063 615 2067
rect 619 2066 620 2067
rect 627 2067 633 2068
rect 627 2066 628 2067
rect 619 2064 628 2066
rect 619 2063 620 2064
rect 614 2062 620 2063
rect 627 2063 628 2064
rect 632 2063 633 2067
rect 627 2062 633 2063
rect 683 2067 689 2068
rect 683 2063 684 2067
rect 688 2066 689 2067
rect 727 2067 733 2068
rect 727 2066 728 2067
rect 688 2064 728 2066
rect 688 2063 689 2064
rect 683 2062 689 2063
rect 727 2063 728 2064
rect 732 2063 733 2067
rect 727 2062 733 2063
rect 739 2067 745 2068
rect 739 2063 740 2067
rect 744 2066 745 2067
rect 750 2067 756 2068
rect 750 2066 751 2067
rect 744 2064 751 2066
rect 744 2063 745 2064
rect 739 2062 745 2063
rect 750 2063 751 2064
rect 755 2063 756 2067
rect 750 2062 756 2063
rect 782 2067 788 2068
rect 782 2063 783 2067
rect 787 2066 788 2067
rect 795 2067 801 2068
rect 795 2066 796 2067
rect 787 2064 796 2066
rect 787 2063 788 2064
rect 782 2062 788 2063
rect 795 2063 796 2064
rect 800 2063 801 2067
rect 795 2062 801 2063
rect 826 2067 832 2068
rect 826 2063 827 2067
rect 831 2066 832 2067
rect 843 2067 849 2068
rect 843 2066 844 2067
rect 831 2064 844 2066
rect 831 2063 832 2064
rect 826 2062 832 2063
rect 843 2063 844 2064
rect 848 2063 849 2067
rect 843 2062 849 2063
rect 874 2067 880 2068
rect 874 2063 875 2067
rect 879 2066 880 2067
rect 899 2067 905 2068
rect 899 2066 900 2067
rect 879 2064 900 2066
rect 879 2063 880 2064
rect 874 2062 880 2063
rect 899 2063 900 2064
rect 904 2063 905 2067
rect 899 2062 905 2063
rect 955 2067 961 2068
rect 955 2063 956 2067
rect 960 2066 961 2067
rect 1002 2067 1008 2068
rect 1002 2066 1003 2067
rect 960 2064 1003 2066
rect 960 2063 961 2064
rect 955 2062 961 2063
rect 1002 2063 1003 2064
rect 1007 2063 1008 2067
rect 1002 2062 1008 2063
rect 1011 2067 1017 2068
rect 1011 2063 1012 2067
rect 1016 2066 1017 2067
rect 1058 2067 1064 2068
rect 1058 2066 1059 2067
rect 1016 2064 1059 2066
rect 1016 2063 1017 2064
rect 1011 2062 1017 2063
rect 1058 2063 1059 2064
rect 1063 2063 1064 2067
rect 1058 2062 1064 2063
rect 1067 2067 1073 2068
rect 1067 2063 1068 2067
rect 1072 2066 1073 2067
rect 1150 2067 1156 2068
rect 1150 2066 1151 2067
rect 1072 2064 1151 2066
rect 1072 2063 1073 2064
rect 1067 2062 1073 2063
rect 1150 2063 1151 2064
rect 1155 2063 1156 2067
rect 1150 2062 1156 2063
rect 1322 2063 1333 2064
rect 1278 2060 1284 2061
rect 382 2059 388 2060
rect 382 2055 383 2059
rect 387 2055 388 2059
rect 382 2054 388 2055
rect 422 2059 428 2060
rect 422 2055 423 2059
rect 427 2055 428 2059
rect 422 2054 428 2055
rect 462 2059 468 2060
rect 462 2055 463 2059
rect 467 2055 468 2059
rect 462 2054 468 2055
rect 502 2059 508 2060
rect 502 2055 503 2059
rect 507 2055 508 2059
rect 502 2054 508 2055
rect 542 2059 548 2060
rect 542 2055 543 2059
rect 547 2055 548 2059
rect 542 2054 548 2055
rect 582 2059 588 2060
rect 582 2055 583 2059
rect 587 2055 588 2059
rect 582 2054 588 2055
rect 630 2059 636 2060
rect 630 2055 631 2059
rect 635 2055 636 2059
rect 630 2054 636 2055
rect 686 2059 692 2060
rect 686 2055 687 2059
rect 691 2055 692 2059
rect 686 2054 692 2055
rect 742 2059 748 2060
rect 742 2055 743 2059
rect 747 2055 748 2059
rect 742 2054 748 2055
rect 798 2059 804 2060
rect 798 2055 799 2059
rect 803 2055 804 2059
rect 798 2054 804 2055
rect 846 2059 852 2060
rect 846 2055 847 2059
rect 851 2055 852 2059
rect 846 2054 852 2055
rect 902 2059 908 2060
rect 902 2055 903 2059
rect 907 2055 908 2059
rect 902 2054 908 2055
rect 958 2059 964 2060
rect 958 2055 959 2059
rect 963 2055 964 2059
rect 958 2054 964 2055
rect 1014 2059 1020 2060
rect 1014 2055 1015 2059
rect 1019 2055 1020 2059
rect 1014 2054 1020 2055
rect 1070 2059 1076 2060
rect 1070 2055 1071 2059
rect 1075 2055 1076 2059
rect 1278 2056 1279 2060
rect 1283 2056 1284 2060
rect 1322 2059 1323 2063
rect 1327 2059 1328 2063
rect 1332 2059 1333 2063
rect 1322 2058 1333 2059
rect 1338 2063 1344 2064
rect 1338 2059 1339 2063
rect 1343 2062 1344 2063
rect 1367 2063 1373 2064
rect 1367 2062 1368 2063
rect 1343 2060 1368 2062
rect 1343 2059 1344 2060
rect 1338 2058 1344 2059
rect 1367 2059 1368 2060
rect 1372 2059 1373 2063
rect 1367 2058 1373 2059
rect 1423 2063 1429 2064
rect 1423 2059 1424 2063
rect 1428 2062 1429 2063
rect 1470 2063 1476 2064
rect 1470 2062 1471 2063
rect 1428 2060 1471 2062
rect 1428 2059 1429 2060
rect 1423 2058 1429 2059
rect 1470 2059 1471 2060
rect 1475 2059 1476 2063
rect 1470 2058 1476 2059
rect 1503 2063 1509 2064
rect 1503 2059 1504 2063
rect 1508 2062 1509 2063
rect 1546 2063 1552 2064
rect 1546 2062 1547 2063
rect 1508 2060 1547 2062
rect 1508 2059 1509 2060
rect 1503 2058 1509 2059
rect 1546 2059 1547 2060
rect 1551 2059 1552 2063
rect 1546 2058 1552 2059
rect 1591 2063 1597 2064
rect 1591 2059 1592 2063
rect 1596 2062 1597 2063
rect 1654 2063 1660 2064
rect 1654 2062 1655 2063
rect 1596 2060 1655 2062
rect 1596 2059 1597 2060
rect 1591 2058 1597 2059
rect 1654 2059 1655 2060
rect 1659 2059 1660 2063
rect 1654 2058 1660 2059
rect 1670 2063 1676 2064
rect 1670 2059 1671 2063
rect 1675 2062 1676 2063
rect 1687 2063 1693 2064
rect 1687 2062 1688 2063
rect 1675 2060 1688 2062
rect 1675 2059 1676 2060
rect 1670 2058 1676 2059
rect 1687 2059 1688 2060
rect 1692 2059 1693 2063
rect 1687 2058 1693 2059
rect 1774 2063 1780 2064
rect 1774 2059 1775 2063
rect 1779 2062 1780 2063
rect 1783 2063 1789 2064
rect 1783 2062 1784 2063
rect 1779 2060 1784 2062
rect 1779 2059 1780 2060
rect 1774 2058 1780 2059
rect 1783 2059 1784 2060
rect 1788 2059 1789 2063
rect 1783 2058 1789 2059
rect 1791 2063 1797 2064
rect 1791 2059 1792 2063
rect 1796 2062 1797 2063
rect 1871 2063 1877 2064
rect 1871 2062 1872 2063
rect 1796 2060 1872 2062
rect 1796 2059 1797 2060
rect 1791 2058 1797 2059
rect 1871 2059 1872 2060
rect 1876 2059 1877 2063
rect 1871 2058 1877 2059
rect 1959 2063 1965 2064
rect 1959 2059 1960 2063
rect 1964 2062 1965 2063
rect 2006 2063 2012 2064
rect 2006 2062 2007 2063
rect 1964 2060 2007 2062
rect 1964 2059 1965 2060
rect 1959 2058 1965 2059
rect 2006 2059 2007 2060
rect 2011 2059 2012 2063
rect 2006 2058 2012 2059
rect 2039 2063 2045 2064
rect 2039 2059 2040 2063
rect 2044 2062 2045 2063
rect 2054 2063 2060 2064
rect 2054 2062 2055 2063
rect 2044 2060 2055 2062
rect 2044 2059 2045 2060
rect 2039 2058 2045 2059
rect 2054 2059 2055 2060
rect 2059 2059 2060 2063
rect 2054 2058 2060 2059
rect 2119 2063 2125 2064
rect 2119 2059 2120 2063
rect 2124 2062 2125 2063
rect 2158 2063 2164 2064
rect 2158 2062 2159 2063
rect 2124 2060 2159 2062
rect 2124 2059 2125 2060
rect 2119 2058 2125 2059
rect 2158 2059 2159 2060
rect 2163 2059 2164 2063
rect 2158 2058 2164 2059
rect 2182 2063 2188 2064
rect 2182 2059 2183 2063
rect 2187 2062 2188 2063
rect 2191 2063 2197 2064
rect 2191 2062 2192 2063
rect 2187 2060 2192 2062
rect 2187 2059 2188 2060
rect 2182 2058 2188 2059
rect 2191 2059 2192 2060
rect 2196 2059 2197 2063
rect 2263 2063 2269 2064
rect 2263 2062 2264 2063
rect 2191 2058 2197 2059
rect 2200 2060 2264 2062
rect 1278 2055 1284 2056
rect 2102 2055 2108 2056
rect 1070 2054 1076 2055
rect 2102 2051 2103 2055
rect 2107 2054 2108 2055
rect 2200 2054 2202 2060
rect 2263 2059 2264 2060
rect 2268 2059 2269 2063
rect 2263 2058 2269 2059
rect 2274 2063 2280 2064
rect 2274 2059 2275 2063
rect 2279 2062 2280 2063
rect 2335 2063 2341 2064
rect 2335 2062 2336 2063
rect 2279 2060 2336 2062
rect 2279 2059 2280 2060
rect 2274 2058 2280 2059
rect 2335 2059 2336 2060
rect 2340 2059 2341 2063
rect 2335 2058 2341 2059
rect 2343 2063 2349 2064
rect 2343 2059 2344 2063
rect 2348 2062 2349 2063
rect 2383 2063 2389 2064
rect 2383 2062 2384 2063
rect 2348 2060 2384 2062
rect 2348 2059 2349 2060
rect 2343 2058 2349 2059
rect 2383 2059 2384 2060
rect 2388 2059 2389 2063
rect 2383 2058 2389 2059
rect 2406 2060 2412 2061
rect 2406 2056 2407 2060
rect 2411 2056 2412 2060
rect 2406 2055 2412 2056
rect 2107 2052 2202 2054
rect 2107 2051 2108 2052
rect 2102 2050 2108 2051
rect 1302 2037 1308 2038
rect 110 2036 116 2037
rect 110 2032 111 2036
rect 115 2032 116 2036
rect 1238 2036 1244 2037
rect 1238 2032 1239 2036
rect 1243 2032 1244 2036
rect 1302 2033 1303 2037
rect 1307 2033 1308 2037
rect 1302 2032 1308 2033
rect 1342 2037 1348 2038
rect 1342 2033 1343 2037
rect 1347 2033 1348 2037
rect 1342 2032 1348 2033
rect 1398 2037 1404 2038
rect 1398 2033 1399 2037
rect 1403 2033 1404 2037
rect 1398 2032 1404 2033
rect 1478 2037 1484 2038
rect 1478 2033 1479 2037
rect 1483 2033 1484 2037
rect 1478 2032 1484 2033
rect 1566 2037 1572 2038
rect 1566 2033 1567 2037
rect 1571 2033 1572 2037
rect 1566 2032 1572 2033
rect 1662 2037 1668 2038
rect 1662 2033 1663 2037
rect 1667 2033 1668 2037
rect 1662 2032 1668 2033
rect 1758 2037 1764 2038
rect 1758 2033 1759 2037
rect 1763 2033 1764 2037
rect 1758 2032 1764 2033
rect 1846 2037 1852 2038
rect 1846 2033 1847 2037
rect 1851 2033 1852 2037
rect 1846 2032 1852 2033
rect 1934 2037 1940 2038
rect 1934 2033 1935 2037
rect 1939 2033 1940 2037
rect 1934 2032 1940 2033
rect 2014 2037 2020 2038
rect 2014 2033 2015 2037
rect 2019 2033 2020 2037
rect 2014 2032 2020 2033
rect 2094 2037 2100 2038
rect 2094 2033 2095 2037
rect 2099 2033 2100 2037
rect 2094 2032 2100 2033
rect 2166 2037 2172 2038
rect 2166 2033 2167 2037
rect 2171 2033 2172 2037
rect 2166 2032 2172 2033
rect 2238 2037 2244 2038
rect 2238 2033 2239 2037
rect 2243 2033 2244 2037
rect 2238 2032 2244 2033
rect 2310 2037 2316 2038
rect 2310 2033 2311 2037
rect 2315 2033 2316 2037
rect 2310 2032 2316 2033
rect 2358 2037 2364 2038
rect 2358 2033 2359 2037
rect 2363 2033 2364 2037
rect 2358 2032 2364 2033
rect 110 2031 116 2032
rect 407 2031 416 2032
rect 407 2027 408 2031
rect 415 2027 416 2031
rect 407 2026 416 2027
rect 446 2031 453 2032
rect 446 2027 447 2031
rect 452 2027 453 2031
rect 446 2026 453 2027
rect 487 2031 496 2032
rect 487 2027 488 2031
rect 495 2027 496 2031
rect 487 2026 496 2027
rect 526 2031 533 2032
rect 526 2027 527 2031
rect 532 2027 533 2031
rect 526 2026 533 2027
rect 567 2031 576 2032
rect 567 2027 568 2031
rect 575 2027 576 2031
rect 567 2026 576 2027
rect 607 2031 616 2032
rect 607 2027 608 2031
rect 615 2027 616 2031
rect 607 2026 616 2027
rect 654 2031 661 2032
rect 654 2027 655 2031
rect 660 2027 661 2031
rect 654 2026 661 2027
rect 663 2031 669 2032
rect 663 2027 664 2031
rect 668 2030 669 2031
rect 711 2031 717 2032
rect 711 2030 712 2031
rect 668 2028 712 2030
rect 668 2027 669 2028
rect 663 2026 669 2027
rect 711 2027 712 2028
rect 716 2027 717 2031
rect 711 2026 717 2027
rect 727 2031 733 2032
rect 727 2027 728 2031
rect 732 2030 733 2031
rect 767 2031 773 2032
rect 767 2030 768 2031
rect 732 2028 768 2030
rect 732 2027 733 2028
rect 727 2026 733 2027
rect 767 2027 768 2028
rect 772 2027 773 2031
rect 767 2026 773 2027
rect 823 2031 832 2032
rect 823 2027 824 2031
rect 831 2027 832 2031
rect 823 2026 832 2027
rect 871 2031 880 2032
rect 871 2027 872 2031
rect 879 2027 880 2031
rect 871 2026 880 2027
rect 886 2031 892 2032
rect 886 2027 887 2031
rect 891 2030 892 2031
rect 927 2031 933 2032
rect 927 2030 928 2031
rect 891 2028 928 2030
rect 891 2027 892 2028
rect 886 2026 892 2027
rect 927 2027 928 2028
rect 932 2027 933 2031
rect 983 2031 989 2032
rect 983 2030 984 2031
rect 927 2026 933 2027
rect 936 2028 984 2030
rect 878 2023 884 2024
rect 110 2019 116 2020
rect 110 2015 111 2019
rect 115 2015 116 2019
rect 878 2019 879 2023
rect 883 2022 884 2023
rect 936 2022 938 2028
rect 983 2027 984 2028
rect 988 2027 989 2031
rect 983 2026 989 2027
rect 1002 2031 1008 2032
rect 1002 2027 1003 2031
rect 1007 2030 1008 2031
rect 1039 2031 1045 2032
rect 1039 2030 1040 2031
rect 1007 2028 1040 2030
rect 1007 2027 1008 2028
rect 1002 2026 1008 2027
rect 1039 2027 1040 2028
rect 1044 2027 1045 2031
rect 1039 2026 1045 2027
rect 1058 2031 1064 2032
rect 1058 2027 1059 2031
rect 1063 2030 1064 2031
rect 1095 2031 1101 2032
rect 1238 2031 1244 2032
rect 1095 2030 1096 2031
rect 1063 2028 1096 2030
rect 1063 2027 1064 2028
rect 1058 2026 1064 2027
rect 1095 2027 1096 2028
rect 1100 2027 1101 2031
rect 1095 2026 1101 2027
rect 1299 2027 1305 2028
rect 1299 2023 1300 2027
rect 1304 2026 1305 2027
rect 1330 2027 1336 2028
rect 1330 2026 1331 2027
rect 1304 2024 1331 2026
rect 1304 2023 1305 2024
rect 1299 2022 1305 2023
rect 1330 2023 1331 2024
rect 1335 2023 1336 2027
rect 1330 2022 1336 2023
rect 1339 2027 1345 2028
rect 1339 2023 1340 2027
rect 1344 2026 1345 2027
rect 1374 2027 1380 2028
rect 1374 2026 1375 2027
rect 1344 2024 1375 2026
rect 1344 2023 1345 2024
rect 1339 2022 1345 2023
rect 1374 2023 1375 2024
rect 1379 2023 1380 2027
rect 1374 2022 1380 2023
rect 1395 2027 1401 2028
rect 1395 2023 1396 2027
rect 1400 2026 1401 2027
rect 1406 2027 1412 2028
rect 1406 2026 1407 2027
rect 1400 2024 1407 2026
rect 1400 2023 1401 2024
rect 1395 2022 1401 2023
rect 1406 2023 1407 2024
rect 1411 2023 1412 2027
rect 1406 2022 1412 2023
rect 1470 2027 1481 2028
rect 1470 2023 1471 2027
rect 1475 2023 1476 2027
rect 1480 2023 1481 2027
rect 1470 2022 1481 2023
rect 1546 2027 1552 2028
rect 1546 2023 1547 2027
rect 1551 2026 1552 2027
rect 1563 2027 1569 2028
rect 1563 2026 1564 2027
rect 1551 2024 1564 2026
rect 1551 2023 1552 2024
rect 1546 2022 1552 2023
rect 1563 2023 1564 2024
rect 1568 2023 1569 2027
rect 1563 2022 1569 2023
rect 1654 2027 1665 2028
rect 1654 2023 1655 2027
rect 1659 2023 1660 2027
rect 1664 2023 1665 2027
rect 1654 2022 1665 2023
rect 1755 2027 1761 2028
rect 1755 2023 1756 2027
rect 1760 2026 1761 2027
rect 1791 2027 1797 2028
rect 1791 2026 1792 2027
rect 1760 2024 1792 2026
rect 1760 2023 1761 2024
rect 1755 2022 1761 2023
rect 1791 2023 1792 2024
rect 1796 2023 1797 2027
rect 1791 2022 1797 2023
rect 1843 2027 1849 2028
rect 1843 2023 1844 2027
rect 1848 2026 1849 2027
rect 1862 2027 1868 2028
rect 1862 2026 1863 2027
rect 1848 2024 1863 2026
rect 1848 2023 1849 2024
rect 1843 2022 1849 2023
rect 1862 2023 1863 2024
rect 1867 2023 1868 2027
rect 1862 2022 1868 2023
rect 1931 2027 1937 2028
rect 1931 2023 1932 2027
rect 1936 2026 1937 2027
rect 1942 2027 1948 2028
rect 1942 2026 1943 2027
rect 1936 2024 1943 2026
rect 1936 2023 1937 2024
rect 1931 2022 1937 2023
rect 1942 2023 1943 2024
rect 1947 2023 1948 2027
rect 1942 2022 1948 2023
rect 2006 2027 2017 2028
rect 2006 2023 2007 2027
rect 2011 2023 2012 2027
rect 2016 2023 2017 2027
rect 2006 2022 2017 2023
rect 2091 2027 2097 2028
rect 2091 2023 2092 2027
rect 2096 2026 2097 2027
rect 2102 2027 2108 2028
rect 2102 2026 2103 2027
rect 2096 2024 2103 2026
rect 2096 2023 2097 2024
rect 2091 2022 2097 2023
rect 2102 2023 2103 2024
rect 2107 2023 2108 2027
rect 2102 2022 2108 2023
rect 2158 2027 2169 2028
rect 2158 2023 2159 2027
rect 2163 2023 2164 2027
rect 2168 2023 2169 2027
rect 2158 2022 2169 2023
rect 2235 2027 2241 2028
rect 2235 2023 2236 2027
rect 2240 2026 2241 2027
rect 2274 2027 2280 2028
rect 2274 2026 2275 2027
rect 2240 2024 2275 2026
rect 2240 2023 2241 2024
rect 2235 2022 2241 2023
rect 2274 2023 2275 2024
rect 2279 2023 2280 2027
rect 2274 2022 2280 2023
rect 2307 2027 2313 2028
rect 2307 2023 2308 2027
rect 2312 2026 2313 2027
rect 2342 2027 2348 2028
rect 2342 2026 2343 2027
rect 2312 2024 2343 2026
rect 2312 2023 2313 2024
rect 2307 2022 2313 2023
rect 2342 2023 2343 2024
rect 2347 2023 2348 2027
rect 2342 2022 2348 2023
rect 2355 2027 2361 2028
rect 2355 2023 2356 2027
rect 2360 2026 2361 2027
rect 2366 2027 2372 2028
rect 2366 2026 2367 2027
rect 2360 2024 2367 2026
rect 2360 2023 2361 2024
rect 2355 2022 2361 2023
rect 2366 2023 2367 2024
rect 2371 2023 2372 2027
rect 2366 2022 2372 2023
rect 883 2020 938 2022
rect 883 2019 884 2020
rect 878 2018 884 2019
rect 1238 2019 1244 2020
rect 110 2014 116 2015
rect 1238 2015 1239 2019
rect 1243 2015 1244 2019
rect 1238 2014 1244 2015
rect 1670 2015 1676 2016
rect 1670 2014 1671 2015
rect 382 2012 388 2013
rect 382 2008 383 2012
rect 387 2008 388 2012
rect 382 2007 388 2008
rect 422 2012 428 2013
rect 422 2008 423 2012
rect 427 2008 428 2012
rect 422 2007 428 2008
rect 462 2012 468 2013
rect 462 2008 463 2012
rect 467 2008 468 2012
rect 462 2007 468 2008
rect 502 2012 508 2013
rect 502 2008 503 2012
rect 507 2008 508 2012
rect 502 2007 508 2008
rect 542 2012 548 2013
rect 542 2008 543 2012
rect 547 2008 548 2012
rect 542 2007 548 2008
rect 582 2012 588 2013
rect 582 2008 583 2012
rect 587 2008 588 2012
rect 582 2007 588 2008
rect 630 2012 636 2013
rect 630 2008 631 2012
rect 635 2008 636 2012
rect 630 2007 636 2008
rect 686 2012 692 2013
rect 686 2008 687 2012
rect 691 2008 692 2012
rect 686 2007 692 2008
rect 742 2012 748 2013
rect 742 2008 743 2012
rect 747 2008 748 2012
rect 742 2007 748 2008
rect 798 2012 804 2013
rect 798 2008 799 2012
rect 803 2008 804 2012
rect 798 2007 804 2008
rect 846 2012 852 2013
rect 846 2008 847 2012
rect 851 2008 852 2012
rect 846 2007 852 2008
rect 902 2012 908 2013
rect 902 2008 903 2012
rect 907 2008 908 2012
rect 902 2007 908 2008
rect 958 2012 964 2013
rect 958 2008 959 2012
rect 963 2008 964 2012
rect 958 2007 964 2008
rect 1014 2012 1020 2013
rect 1014 2008 1015 2012
rect 1019 2008 1020 2012
rect 1014 2007 1020 2008
rect 1070 2012 1076 2013
rect 1070 2008 1071 2012
rect 1075 2008 1076 2012
rect 1572 2012 1671 2014
rect 1572 2010 1574 2012
rect 1670 2011 1671 2012
rect 1675 2011 1676 2015
rect 2343 2015 2349 2016
rect 2343 2014 2344 2015
rect 1670 2010 1676 2011
rect 2252 2012 2344 2014
rect 2252 2010 2254 2012
rect 2343 2011 2344 2012
rect 2348 2011 2349 2015
rect 2343 2010 2349 2011
rect 1571 2009 1577 2010
rect 1070 2007 1076 2008
rect 1299 2007 1305 2008
rect 1299 2003 1300 2007
rect 1304 2006 1305 2007
rect 1322 2007 1328 2008
rect 1322 2006 1323 2007
rect 1304 2004 1323 2006
rect 1304 2003 1305 2004
rect 1299 2002 1305 2003
rect 1322 2003 1323 2004
rect 1327 2003 1328 2007
rect 1322 2002 1328 2003
rect 1330 2007 1336 2008
rect 1330 2003 1331 2007
rect 1335 2006 1336 2007
rect 1347 2007 1353 2008
rect 1347 2006 1348 2007
rect 1335 2004 1348 2006
rect 1335 2003 1336 2004
rect 1330 2002 1336 2003
rect 1347 2003 1348 2004
rect 1352 2003 1353 2007
rect 1347 2002 1353 2003
rect 1419 2007 1425 2008
rect 1419 2003 1420 2007
rect 1424 2006 1425 2007
rect 1442 2007 1448 2008
rect 1442 2006 1443 2007
rect 1424 2004 1443 2006
rect 1424 2003 1425 2004
rect 1419 2002 1425 2003
rect 1442 2003 1443 2004
rect 1447 2003 1448 2007
rect 1442 2002 1448 2003
rect 1450 2007 1456 2008
rect 1450 2003 1451 2007
rect 1455 2006 1456 2007
rect 1491 2007 1497 2008
rect 1491 2006 1492 2007
rect 1455 2004 1492 2006
rect 1455 2003 1456 2004
rect 1450 2002 1456 2003
rect 1491 2003 1492 2004
rect 1496 2003 1497 2007
rect 1571 2005 1572 2009
rect 1576 2005 1577 2009
rect 2251 2009 2257 2010
rect 1571 2004 1577 2005
rect 1659 2007 1665 2008
rect 1491 2002 1497 2003
rect 1659 2003 1660 2007
rect 1664 2006 1665 2007
rect 1690 2007 1696 2008
rect 1664 2004 1686 2006
rect 1664 2003 1665 2004
rect 1659 2002 1665 2003
rect 1302 1999 1308 2000
rect 1302 1995 1303 1999
rect 1307 1995 1308 1999
rect 1302 1994 1308 1995
rect 1350 1999 1356 2000
rect 1350 1995 1351 1999
rect 1355 1995 1356 1999
rect 1350 1994 1356 1995
rect 1422 1999 1428 2000
rect 1422 1995 1423 1999
rect 1427 1995 1428 1999
rect 1422 1994 1428 1995
rect 1494 1999 1500 2000
rect 1494 1995 1495 1999
rect 1499 1995 1500 1999
rect 1494 1994 1500 1995
rect 1574 1999 1580 2000
rect 1574 1995 1575 1999
rect 1579 1995 1580 1999
rect 1574 1994 1580 1995
rect 1662 1999 1668 2000
rect 1662 1995 1663 1999
rect 1667 1995 1668 1999
rect 1684 1998 1686 2004
rect 1690 2003 1691 2007
rect 1695 2006 1696 2007
rect 1747 2007 1753 2008
rect 1747 2006 1748 2007
rect 1695 2004 1748 2006
rect 1695 2003 1696 2004
rect 1690 2002 1696 2003
rect 1747 2003 1748 2004
rect 1752 2003 1753 2007
rect 1747 2002 1753 2003
rect 1778 2007 1784 2008
rect 1778 2003 1779 2007
rect 1783 2006 1784 2007
rect 1835 2007 1841 2008
rect 1835 2006 1836 2007
rect 1783 2004 1836 2006
rect 1783 2003 1784 2004
rect 1778 2002 1784 2003
rect 1835 2003 1836 2004
rect 1840 2003 1841 2007
rect 1835 2002 1841 2003
rect 1915 2007 1921 2008
rect 1915 2003 1916 2007
rect 1920 2006 1921 2007
rect 1926 2007 1932 2008
rect 1926 2006 1927 2007
rect 1920 2004 1927 2006
rect 1920 2003 1921 2004
rect 1915 2002 1921 2003
rect 1926 2003 1927 2004
rect 1931 2003 1932 2007
rect 1926 2002 1932 2003
rect 1946 2007 1952 2008
rect 1946 2003 1947 2007
rect 1951 2006 1952 2007
rect 1995 2007 2001 2008
rect 1995 2006 1996 2007
rect 1951 2004 1996 2006
rect 1951 2003 1952 2004
rect 1946 2002 1952 2003
rect 1995 2003 1996 2004
rect 2000 2003 2001 2007
rect 1995 2002 2001 2003
rect 2067 2007 2073 2008
rect 2067 2003 2068 2007
rect 2072 2006 2073 2007
rect 2122 2007 2128 2008
rect 2122 2006 2123 2007
rect 2072 2004 2123 2006
rect 2072 2003 2073 2004
rect 2067 2002 2073 2003
rect 2122 2003 2123 2004
rect 2127 2003 2128 2007
rect 2122 2002 2128 2003
rect 2131 2007 2137 2008
rect 2131 2003 2132 2007
rect 2136 2006 2137 2007
rect 2174 2007 2180 2008
rect 2174 2006 2175 2007
rect 2136 2004 2175 2006
rect 2136 2003 2137 2004
rect 2131 2002 2137 2003
rect 2174 2003 2175 2004
rect 2179 2003 2180 2007
rect 2174 2002 2180 2003
rect 2182 2007 2193 2008
rect 2182 2003 2183 2007
rect 2187 2003 2188 2007
rect 2192 2003 2193 2007
rect 2251 2005 2252 2009
rect 2256 2005 2257 2009
rect 2251 2004 2257 2005
rect 2315 2007 2321 2008
rect 2182 2002 2193 2003
rect 2315 2003 2316 2007
rect 2320 2006 2321 2007
rect 2334 2007 2340 2008
rect 2334 2006 2335 2007
rect 2320 2004 2335 2006
rect 2320 2003 2321 2004
rect 2315 2002 2321 2003
rect 2334 2003 2335 2004
rect 2339 2003 2340 2007
rect 2334 2002 2340 2003
rect 2355 2007 2361 2008
rect 2355 2003 2356 2007
rect 2360 2006 2361 2007
rect 2382 2007 2388 2008
rect 2382 2006 2383 2007
rect 2360 2004 2383 2006
rect 2360 2003 2361 2004
rect 2355 2002 2361 2003
rect 2382 2003 2383 2004
rect 2387 2003 2388 2007
rect 2382 2002 2388 2003
rect 1734 1999 1740 2000
rect 1734 1998 1735 1999
rect 1684 1996 1735 1998
rect 1662 1994 1668 1995
rect 1734 1995 1735 1996
rect 1739 1995 1740 1999
rect 1734 1994 1740 1995
rect 1750 1999 1756 2000
rect 1750 1995 1751 1999
rect 1755 1995 1756 1999
rect 1750 1994 1756 1995
rect 1838 1999 1844 2000
rect 1838 1995 1839 1999
rect 1843 1995 1844 1999
rect 1838 1994 1844 1995
rect 1918 1999 1924 2000
rect 1918 1995 1919 1999
rect 1923 1995 1924 1999
rect 1918 1994 1924 1995
rect 1998 1999 2004 2000
rect 1998 1995 1999 1999
rect 2003 1995 2004 1999
rect 1998 1994 2004 1995
rect 2070 1999 2076 2000
rect 2070 1995 2071 1999
rect 2075 1995 2076 1999
rect 2070 1994 2076 1995
rect 2134 1999 2140 2000
rect 2134 1995 2135 1999
rect 2139 1995 2140 1999
rect 2134 1994 2140 1995
rect 2190 1999 2196 2000
rect 2190 1995 2191 1999
rect 2195 1995 2196 1999
rect 2190 1994 2196 1995
rect 2254 1999 2260 2000
rect 2254 1995 2255 1999
rect 2259 1995 2260 1999
rect 2254 1994 2260 1995
rect 2318 1999 2324 2000
rect 2318 1995 2319 1999
rect 2323 1995 2324 1999
rect 2318 1994 2324 1995
rect 2358 1999 2364 2000
rect 2358 1995 2359 1999
rect 2363 1995 2364 1999
rect 2358 1994 2364 1995
rect 366 1992 372 1993
rect 366 1988 367 1992
rect 371 1988 372 1992
rect 366 1987 372 1988
rect 406 1992 412 1993
rect 406 1988 407 1992
rect 411 1988 412 1992
rect 406 1987 412 1988
rect 454 1992 460 1993
rect 454 1988 455 1992
rect 459 1988 460 1992
rect 454 1987 460 1988
rect 510 1992 516 1993
rect 510 1988 511 1992
rect 515 1988 516 1992
rect 510 1987 516 1988
rect 566 1992 572 1993
rect 566 1988 567 1992
rect 571 1988 572 1992
rect 566 1987 572 1988
rect 630 1992 636 1993
rect 630 1988 631 1992
rect 635 1988 636 1992
rect 630 1987 636 1988
rect 694 1992 700 1993
rect 694 1988 695 1992
rect 699 1988 700 1992
rect 694 1987 700 1988
rect 758 1992 764 1993
rect 758 1988 759 1992
rect 763 1988 764 1992
rect 758 1987 764 1988
rect 814 1992 820 1993
rect 814 1988 815 1992
rect 819 1988 820 1992
rect 814 1987 820 1988
rect 870 1992 876 1993
rect 870 1988 871 1992
rect 875 1988 876 1992
rect 870 1987 876 1988
rect 934 1992 940 1993
rect 934 1988 935 1992
rect 939 1988 940 1992
rect 934 1987 940 1988
rect 998 1992 1004 1993
rect 998 1988 999 1992
rect 1003 1988 1004 1992
rect 998 1987 1004 1988
rect 1062 1992 1068 1993
rect 1062 1988 1063 1992
rect 1067 1988 1068 1992
rect 1062 1987 1068 1988
rect 110 1985 116 1986
rect 110 1981 111 1985
rect 115 1981 116 1985
rect 110 1980 116 1981
rect 1238 1985 1244 1986
rect 1238 1981 1239 1985
rect 1243 1981 1244 1985
rect 1238 1980 1244 1981
rect 1442 1979 1448 1980
rect 1278 1976 1284 1977
rect 1278 1972 1279 1976
rect 1283 1972 1284 1976
rect 1442 1975 1443 1979
rect 1447 1978 1448 1979
rect 1926 1979 1932 1980
rect 1447 1976 1534 1978
rect 1447 1975 1448 1976
rect 1442 1974 1448 1975
rect 391 1971 400 1972
rect 110 1968 116 1969
rect 110 1964 111 1968
rect 115 1964 116 1968
rect 391 1967 392 1971
rect 399 1967 400 1971
rect 391 1966 400 1967
rect 431 1971 437 1972
rect 431 1967 432 1971
rect 436 1970 437 1971
rect 446 1971 452 1972
rect 446 1970 447 1971
rect 436 1968 447 1970
rect 436 1967 437 1968
rect 431 1966 437 1967
rect 446 1967 447 1968
rect 451 1967 452 1971
rect 446 1966 452 1967
rect 478 1971 485 1972
rect 478 1967 479 1971
rect 484 1967 485 1971
rect 535 1971 541 1972
rect 535 1970 536 1971
rect 478 1966 485 1967
rect 488 1968 536 1970
rect 110 1963 116 1964
rect 374 1963 380 1964
rect 374 1959 375 1963
rect 379 1962 380 1963
rect 488 1962 490 1968
rect 535 1967 536 1968
rect 540 1967 541 1971
rect 535 1966 541 1967
rect 543 1971 549 1972
rect 543 1967 544 1971
rect 548 1970 549 1971
rect 591 1971 597 1972
rect 591 1970 592 1971
rect 548 1968 592 1970
rect 548 1967 549 1968
rect 543 1966 549 1967
rect 591 1967 592 1968
rect 596 1967 597 1971
rect 591 1966 597 1967
rect 602 1971 608 1972
rect 602 1967 603 1971
rect 607 1970 608 1971
rect 655 1971 661 1972
rect 655 1970 656 1971
rect 607 1968 656 1970
rect 607 1967 608 1968
rect 602 1966 608 1967
rect 655 1967 656 1968
rect 660 1967 661 1971
rect 655 1966 661 1967
rect 719 1971 725 1972
rect 719 1967 720 1971
rect 724 1970 725 1971
rect 750 1971 756 1972
rect 750 1970 751 1971
rect 724 1968 751 1970
rect 724 1967 725 1968
rect 719 1966 725 1967
rect 750 1967 751 1968
rect 755 1967 756 1971
rect 750 1966 756 1967
rect 782 1971 789 1972
rect 782 1967 783 1971
rect 788 1967 789 1971
rect 839 1971 845 1972
rect 839 1970 840 1971
rect 782 1966 789 1967
rect 792 1968 840 1970
rect 379 1960 490 1962
rect 702 1963 708 1964
rect 379 1959 380 1960
rect 374 1958 380 1959
rect 702 1959 703 1963
rect 707 1962 708 1963
rect 792 1962 794 1968
rect 839 1967 840 1968
rect 844 1967 845 1971
rect 839 1966 845 1967
rect 895 1971 901 1972
rect 895 1967 896 1971
rect 900 1970 901 1971
rect 926 1971 932 1972
rect 926 1970 927 1971
rect 900 1968 927 1970
rect 900 1967 901 1968
rect 895 1966 901 1967
rect 926 1967 927 1968
rect 931 1967 932 1971
rect 926 1966 932 1967
rect 959 1971 965 1972
rect 959 1967 960 1971
rect 964 1970 965 1971
rect 990 1971 996 1972
rect 990 1970 991 1971
rect 964 1968 991 1970
rect 964 1967 965 1968
rect 959 1966 965 1967
rect 990 1967 991 1968
rect 995 1967 996 1971
rect 990 1966 996 1967
rect 1023 1971 1029 1972
rect 1023 1967 1024 1971
rect 1028 1970 1029 1971
rect 1054 1971 1060 1972
rect 1054 1970 1055 1971
rect 1028 1968 1055 1970
rect 1028 1967 1029 1968
rect 1023 1966 1029 1967
rect 1054 1967 1055 1968
rect 1059 1967 1060 1971
rect 1054 1966 1060 1967
rect 1070 1971 1076 1972
rect 1070 1967 1071 1971
rect 1075 1970 1076 1971
rect 1087 1971 1093 1972
rect 1278 1971 1284 1972
rect 1327 1971 1336 1972
rect 1087 1970 1088 1971
rect 1075 1968 1088 1970
rect 1075 1967 1076 1968
rect 1070 1966 1076 1967
rect 1087 1967 1088 1968
rect 1092 1967 1093 1971
rect 1087 1966 1093 1967
rect 1238 1968 1244 1969
rect 1238 1964 1239 1968
rect 1243 1964 1244 1968
rect 1327 1967 1328 1971
rect 1335 1967 1336 1971
rect 1327 1966 1336 1967
rect 1374 1971 1381 1972
rect 1374 1967 1375 1971
rect 1380 1967 1381 1971
rect 1374 1966 1381 1967
rect 1447 1971 1456 1972
rect 1447 1967 1448 1971
rect 1455 1967 1456 1971
rect 1447 1966 1456 1967
rect 1519 1971 1528 1972
rect 1519 1967 1520 1971
rect 1527 1967 1528 1971
rect 1532 1970 1534 1976
rect 1926 1975 1927 1979
rect 1931 1978 1932 1979
rect 2334 1979 2340 1980
rect 1931 1976 2074 1978
rect 1931 1975 1932 1976
rect 1926 1974 1932 1975
rect 1599 1971 1605 1972
rect 1599 1970 1600 1971
rect 1532 1968 1600 1970
rect 1519 1966 1528 1967
rect 1599 1967 1600 1968
rect 1604 1967 1605 1971
rect 1599 1966 1605 1967
rect 1687 1971 1696 1972
rect 1687 1967 1688 1971
rect 1695 1967 1696 1971
rect 1687 1966 1696 1967
rect 1775 1971 1784 1972
rect 1775 1967 1776 1971
rect 1783 1967 1784 1971
rect 1775 1966 1784 1967
rect 1862 1971 1869 1972
rect 1862 1967 1863 1971
rect 1868 1967 1869 1971
rect 1862 1966 1869 1967
rect 1943 1971 1952 1972
rect 1943 1967 1944 1971
rect 1951 1967 1952 1971
rect 1943 1966 1952 1967
rect 2023 1971 2029 1972
rect 2023 1967 2024 1971
rect 2028 1970 2029 1971
rect 2063 1971 2069 1972
rect 2063 1970 2064 1971
rect 2028 1968 2064 1970
rect 2028 1967 2029 1968
rect 2023 1966 2029 1967
rect 2063 1967 2064 1968
rect 2068 1967 2069 1971
rect 2072 1970 2074 1976
rect 2334 1975 2335 1979
rect 2339 1978 2340 1979
rect 2339 1976 2387 1978
rect 2339 1975 2340 1976
rect 2334 1974 2340 1975
rect 2385 1972 2387 1976
rect 2406 1976 2412 1977
rect 2406 1972 2407 1976
rect 2411 1972 2412 1976
rect 2095 1971 2101 1972
rect 2095 1970 2096 1971
rect 2072 1968 2096 1970
rect 2063 1966 2069 1967
rect 2095 1967 2096 1968
rect 2100 1967 2101 1971
rect 2095 1966 2101 1967
rect 2122 1971 2128 1972
rect 2122 1967 2123 1971
rect 2127 1970 2128 1971
rect 2159 1971 2165 1972
rect 2159 1970 2160 1971
rect 2127 1968 2160 1970
rect 2127 1967 2128 1968
rect 2122 1966 2128 1967
rect 2159 1967 2160 1968
rect 2164 1967 2165 1971
rect 2159 1966 2165 1967
rect 2174 1971 2180 1972
rect 2174 1967 2175 1971
rect 2179 1970 2180 1971
rect 2215 1971 2221 1972
rect 2215 1970 2216 1971
rect 2179 1968 2216 1970
rect 2179 1967 2180 1968
rect 2174 1966 2180 1967
rect 2215 1967 2216 1968
rect 2220 1967 2221 1971
rect 2215 1966 2221 1967
rect 2230 1971 2236 1972
rect 2230 1967 2231 1971
rect 2235 1970 2236 1971
rect 2279 1971 2285 1972
rect 2279 1970 2280 1971
rect 2235 1968 2280 1970
rect 2235 1967 2236 1968
rect 2230 1966 2236 1967
rect 2279 1967 2280 1968
rect 2284 1967 2285 1971
rect 2279 1966 2285 1967
rect 2342 1971 2349 1972
rect 2342 1967 2343 1971
rect 2348 1967 2349 1971
rect 2342 1966 2349 1967
rect 2383 1971 2389 1972
rect 2406 1971 2412 1972
rect 2383 1967 2384 1971
rect 2388 1967 2389 1971
rect 2383 1966 2389 1967
rect 1238 1963 1244 1964
rect 707 1960 794 1962
rect 707 1959 708 1960
rect 702 1958 708 1959
rect 1278 1959 1284 1960
rect 1278 1955 1279 1959
rect 1283 1955 1284 1959
rect 1278 1954 1284 1955
rect 2406 1959 2412 1960
rect 2406 1955 2407 1959
rect 2411 1955 2412 1959
rect 2406 1954 2412 1955
rect 1302 1952 1308 1953
rect 1302 1948 1303 1952
rect 1307 1948 1308 1952
rect 1302 1947 1308 1948
rect 1350 1952 1356 1953
rect 1350 1948 1351 1952
rect 1355 1948 1356 1952
rect 1350 1947 1356 1948
rect 1422 1952 1428 1953
rect 1422 1948 1423 1952
rect 1427 1948 1428 1952
rect 1422 1947 1428 1948
rect 1494 1952 1500 1953
rect 1494 1948 1495 1952
rect 1499 1948 1500 1952
rect 1494 1947 1500 1948
rect 1574 1952 1580 1953
rect 1574 1948 1575 1952
rect 1579 1948 1580 1952
rect 1574 1947 1580 1948
rect 1662 1952 1668 1953
rect 1662 1948 1663 1952
rect 1667 1948 1668 1952
rect 1662 1947 1668 1948
rect 1750 1952 1756 1953
rect 1750 1948 1751 1952
rect 1755 1948 1756 1952
rect 1750 1947 1756 1948
rect 1838 1952 1844 1953
rect 1838 1948 1839 1952
rect 1843 1948 1844 1952
rect 1838 1947 1844 1948
rect 1918 1952 1924 1953
rect 1918 1948 1919 1952
rect 1923 1948 1924 1952
rect 1918 1947 1924 1948
rect 1998 1952 2004 1953
rect 1998 1948 1999 1952
rect 2003 1948 2004 1952
rect 1998 1947 2004 1948
rect 2070 1952 2076 1953
rect 2070 1948 2071 1952
rect 2075 1948 2076 1952
rect 2070 1947 2076 1948
rect 2134 1952 2140 1953
rect 2134 1948 2135 1952
rect 2139 1948 2140 1952
rect 2134 1947 2140 1948
rect 2190 1952 2196 1953
rect 2190 1948 2191 1952
rect 2195 1948 2196 1952
rect 2190 1947 2196 1948
rect 2254 1952 2260 1953
rect 2254 1948 2255 1952
rect 2259 1948 2260 1952
rect 2254 1947 2260 1948
rect 2318 1952 2324 1953
rect 2318 1948 2319 1952
rect 2323 1948 2324 1952
rect 2318 1947 2324 1948
rect 2358 1952 2364 1953
rect 2358 1948 2359 1952
rect 2363 1948 2364 1952
rect 2358 1947 2364 1948
rect 366 1945 372 1946
rect 366 1941 367 1945
rect 371 1941 372 1945
rect 366 1940 372 1941
rect 406 1945 412 1946
rect 406 1941 407 1945
rect 411 1941 412 1945
rect 406 1940 412 1941
rect 454 1945 460 1946
rect 454 1941 455 1945
rect 459 1941 460 1945
rect 454 1940 460 1941
rect 510 1945 516 1946
rect 510 1941 511 1945
rect 515 1941 516 1945
rect 510 1940 516 1941
rect 566 1945 572 1946
rect 566 1941 567 1945
rect 571 1941 572 1945
rect 566 1940 572 1941
rect 630 1945 636 1946
rect 630 1941 631 1945
rect 635 1941 636 1945
rect 630 1940 636 1941
rect 694 1945 700 1946
rect 694 1941 695 1945
rect 699 1941 700 1945
rect 694 1940 700 1941
rect 758 1945 764 1946
rect 758 1941 759 1945
rect 763 1941 764 1945
rect 758 1940 764 1941
rect 814 1945 820 1946
rect 814 1941 815 1945
rect 819 1941 820 1945
rect 814 1940 820 1941
rect 870 1945 876 1946
rect 870 1941 871 1945
rect 875 1941 876 1945
rect 870 1940 876 1941
rect 934 1945 940 1946
rect 934 1941 935 1945
rect 939 1941 940 1945
rect 934 1940 940 1941
rect 998 1945 1004 1946
rect 998 1941 999 1945
rect 1003 1941 1004 1945
rect 998 1940 1004 1941
rect 1062 1945 1068 1946
rect 1062 1941 1063 1945
rect 1067 1941 1068 1945
rect 1062 1940 1068 1941
rect 1302 1940 1308 1941
rect 1302 1936 1303 1940
rect 1307 1936 1308 1940
rect 363 1935 369 1936
rect 363 1931 364 1935
rect 368 1934 369 1935
rect 374 1935 380 1936
rect 374 1934 375 1935
rect 368 1932 375 1934
rect 368 1931 369 1932
rect 363 1930 369 1931
rect 374 1931 375 1932
rect 379 1931 380 1935
rect 374 1930 380 1931
rect 394 1935 400 1936
rect 394 1931 395 1935
rect 399 1934 400 1935
rect 403 1935 409 1936
rect 403 1934 404 1935
rect 399 1932 404 1934
rect 399 1931 400 1932
rect 394 1930 400 1931
rect 403 1931 404 1932
rect 408 1931 409 1935
rect 403 1930 409 1931
rect 446 1935 457 1936
rect 446 1931 447 1935
rect 451 1931 452 1935
rect 456 1931 457 1935
rect 446 1930 457 1931
rect 507 1935 513 1936
rect 507 1931 508 1935
rect 512 1934 513 1935
rect 543 1935 549 1936
rect 543 1934 544 1935
rect 512 1932 544 1934
rect 512 1931 513 1932
rect 507 1930 513 1931
rect 543 1931 544 1932
rect 548 1931 549 1935
rect 543 1930 549 1931
rect 563 1935 569 1936
rect 563 1931 564 1935
rect 568 1934 569 1935
rect 602 1935 608 1936
rect 602 1934 603 1935
rect 568 1932 603 1934
rect 568 1931 569 1932
rect 563 1930 569 1931
rect 602 1931 603 1932
rect 607 1931 608 1935
rect 602 1930 608 1931
rect 627 1935 633 1936
rect 627 1931 628 1935
rect 632 1934 633 1935
rect 663 1935 669 1936
rect 663 1934 664 1935
rect 632 1932 664 1934
rect 632 1931 633 1932
rect 627 1930 633 1931
rect 663 1931 664 1932
rect 668 1931 669 1935
rect 663 1930 669 1931
rect 691 1935 697 1936
rect 691 1931 692 1935
rect 696 1934 697 1935
rect 702 1935 708 1936
rect 702 1934 703 1935
rect 696 1932 703 1934
rect 696 1931 697 1932
rect 691 1930 697 1931
rect 702 1931 703 1932
rect 707 1931 708 1935
rect 702 1930 708 1931
rect 750 1935 761 1936
rect 750 1931 751 1935
rect 755 1931 756 1935
rect 760 1931 761 1935
rect 750 1930 761 1931
rect 811 1935 817 1936
rect 811 1931 812 1935
rect 816 1934 817 1935
rect 822 1935 828 1936
rect 822 1934 823 1935
rect 816 1932 823 1934
rect 816 1931 817 1932
rect 811 1930 817 1931
rect 822 1931 823 1932
rect 827 1931 828 1935
rect 822 1930 828 1931
rect 867 1935 873 1936
rect 867 1931 868 1935
rect 872 1934 873 1935
rect 878 1935 884 1936
rect 878 1934 879 1935
rect 872 1932 879 1934
rect 872 1931 873 1932
rect 867 1930 873 1931
rect 878 1931 879 1932
rect 883 1931 884 1935
rect 878 1930 884 1931
rect 926 1935 937 1936
rect 926 1931 927 1935
rect 931 1931 932 1935
rect 936 1931 937 1935
rect 926 1930 937 1931
rect 990 1935 1001 1936
rect 990 1931 991 1935
rect 995 1931 996 1935
rect 1000 1931 1001 1935
rect 990 1930 1001 1931
rect 1054 1935 1065 1936
rect 1302 1935 1308 1936
rect 1358 1940 1364 1941
rect 1358 1936 1359 1940
rect 1363 1936 1364 1940
rect 1358 1935 1364 1936
rect 1446 1940 1452 1941
rect 1446 1936 1447 1940
rect 1451 1936 1452 1940
rect 1446 1935 1452 1936
rect 1534 1940 1540 1941
rect 1534 1936 1535 1940
rect 1539 1936 1540 1940
rect 1534 1935 1540 1936
rect 1622 1940 1628 1941
rect 1622 1936 1623 1940
rect 1627 1936 1628 1940
rect 1622 1935 1628 1936
rect 1710 1940 1716 1941
rect 1710 1936 1711 1940
rect 1715 1936 1716 1940
rect 1710 1935 1716 1936
rect 1790 1940 1796 1941
rect 1790 1936 1791 1940
rect 1795 1936 1796 1940
rect 1790 1935 1796 1936
rect 1862 1940 1868 1941
rect 1862 1936 1863 1940
rect 1867 1936 1868 1940
rect 1862 1935 1868 1936
rect 1934 1940 1940 1941
rect 1934 1936 1935 1940
rect 1939 1936 1940 1940
rect 1934 1935 1940 1936
rect 2006 1940 2012 1941
rect 2006 1936 2007 1940
rect 2011 1936 2012 1940
rect 2006 1935 2012 1936
rect 2078 1940 2084 1941
rect 2078 1936 2079 1940
rect 2083 1936 2084 1940
rect 2078 1935 2084 1936
rect 2150 1940 2156 1941
rect 2150 1936 2151 1940
rect 2155 1936 2156 1940
rect 2150 1935 2156 1936
rect 2222 1940 2228 1941
rect 2222 1936 2223 1940
rect 2227 1936 2228 1940
rect 2222 1935 2228 1936
rect 2302 1940 2308 1941
rect 2302 1936 2303 1940
rect 2307 1936 2308 1940
rect 2302 1935 2308 1936
rect 2358 1940 2364 1941
rect 2358 1936 2359 1940
rect 2363 1936 2364 1940
rect 2358 1935 2364 1936
rect 1054 1931 1055 1935
rect 1059 1931 1060 1935
rect 1064 1931 1065 1935
rect 1054 1930 1065 1931
rect 1278 1933 1284 1934
rect 1278 1929 1279 1933
rect 1283 1929 1284 1933
rect 1278 1928 1284 1929
rect 2406 1933 2412 1934
rect 2406 1929 2407 1933
rect 2411 1929 2412 1933
rect 2406 1928 2412 1929
rect 1070 1927 1076 1928
rect 1070 1926 1071 1927
rect 877 1924 1071 1926
rect 877 1922 879 1924
rect 1070 1923 1071 1924
rect 1075 1923 1076 1927
rect 1070 1922 1076 1923
rect 875 1921 881 1922
rect 171 1919 177 1920
rect 171 1915 172 1919
rect 176 1918 177 1919
rect 190 1919 196 1920
rect 190 1918 191 1919
rect 176 1916 191 1918
rect 176 1915 177 1916
rect 171 1914 177 1915
rect 190 1915 191 1916
rect 195 1915 196 1919
rect 190 1914 196 1915
rect 198 1919 204 1920
rect 198 1915 199 1919
rect 203 1918 204 1919
rect 211 1919 217 1920
rect 211 1918 212 1919
rect 203 1916 212 1918
rect 203 1915 204 1916
rect 198 1914 204 1915
rect 211 1915 212 1916
rect 216 1915 217 1919
rect 211 1914 217 1915
rect 247 1919 253 1920
rect 247 1915 248 1919
rect 252 1918 253 1919
rect 259 1919 265 1920
rect 259 1918 260 1919
rect 252 1916 260 1918
rect 252 1915 253 1916
rect 247 1914 253 1915
rect 259 1915 260 1916
rect 264 1915 265 1919
rect 259 1914 265 1915
rect 315 1919 321 1920
rect 315 1915 316 1919
rect 320 1918 321 1919
rect 378 1919 384 1920
rect 378 1918 379 1919
rect 320 1916 379 1918
rect 320 1915 321 1916
rect 315 1914 321 1915
rect 378 1915 379 1916
rect 383 1915 384 1919
rect 378 1914 384 1915
rect 387 1919 393 1920
rect 387 1915 388 1919
rect 392 1918 393 1919
rect 455 1919 461 1920
rect 455 1918 456 1919
rect 392 1916 456 1918
rect 392 1915 393 1916
rect 387 1914 393 1915
rect 455 1915 456 1916
rect 460 1915 461 1919
rect 455 1914 461 1915
rect 467 1919 473 1920
rect 467 1915 468 1919
rect 472 1918 473 1919
rect 478 1919 484 1920
rect 478 1918 479 1919
rect 472 1916 479 1918
rect 472 1915 473 1916
rect 467 1914 473 1915
rect 478 1915 479 1916
rect 483 1915 484 1919
rect 478 1914 484 1915
rect 498 1919 504 1920
rect 498 1915 499 1919
rect 503 1918 504 1919
rect 547 1919 553 1920
rect 547 1918 548 1919
rect 503 1916 548 1918
rect 503 1915 504 1916
rect 498 1914 504 1915
rect 547 1915 548 1916
rect 552 1915 553 1919
rect 547 1914 553 1915
rect 635 1919 641 1920
rect 635 1915 636 1919
rect 640 1918 641 1919
rect 654 1919 660 1920
rect 654 1918 655 1919
rect 640 1916 655 1918
rect 640 1915 641 1916
rect 635 1914 641 1915
rect 654 1915 655 1916
rect 659 1915 660 1919
rect 654 1914 660 1915
rect 671 1919 677 1920
rect 671 1915 672 1919
rect 676 1918 677 1919
rect 715 1919 721 1920
rect 715 1918 716 1919
rect 676 1916 716 1918
rect 676 1915 677 1916
rect 671 1914 677 1915
rect 715 1915 716 1916
rect 720 1915 721 1919
rect 715 1914 721 1915
rect 746 1919 752 1920
rect 746 1915 747 1919
rect 751 1918 752 1919
rect 795 1919 801 1920
rect 795 1918 796 1919
rect 751 1916 796 1918
rect 751 1915 752 1916
rect 746 1914 752 1915
rect 795 1915 796 1916
rect 800 1915 801 1919
rect 875 1917 876 1921
rect 880 1917 881 1921
rect 875 1916 881 1917
rect 902 1919 908 1920
rect 795 1914 801 1915
rect 902 1915 903 1919
rect 907 1918 908 1919
rect 955 1919 961 1920
rect 955 1918 956 1919
rect 907 1916 956 1918
rect 907 1915 908 1916
rect 902 1914 908 1915
rect 955 1915 956 1916
rect 960 1915 961 1919
rect 955 1914 961 1915
rect 986 1919 992 1920
rect 986 1915 987 1919
rect 991 1918 992 1919
rect 1035 1919 1041 1920
rect 1035 1918 1036 1919
rect 991 1916 1036 1918
rect 991 1915 992 1916
rect 986 1914 992 1915
rect 1035 1915 1036 1916
rect 1040 1915 1041 1919
rect 1035 1914 1041 1915
rect 1070 1919 1076 1920
rect 1070 1915 1071 1919
rect 1075 1918 1076 1919
rect 1115 1919 1121 1920
rect 1115 1918 1116 1919
rect 1075 1916 1116 1918
rect 1075 1915 1076 1916
rect 1070 1914 1076 1915
rect 1115 1915 1116 1916
rect 1120 1915 1121 1919
rect 1322 1919 1333 1920
rect 1115 1914 1121 1915
rect 1278 1916 1284 1917
rect 1278 1912 1279 1916
rect 1283 1912 1284 1916
rect 1322 1915 1323 1919
rect 1327 1915 1328 1919
rect 1332 1915 1333 1919
rect 1322 1914 1333 1915
rect 1335 1919 1341 1920
rect 1335 1915 1336 1919
rect 1340 1918 1341 1919
rect 1383 1919 1389 1920
rect 1383 1918 1384 1919
rect 1340 1916 1384 1918
rect 1340 1915 1341 1916
rect 1335 1914 1341 1915
rect 1383 1915 1384 1916
rect 1388 1915 1389 1919
rect 1383 1914 1389 1915
rect 1391 1919 1397 1920
rect 1391 1915 1392 1919
rect 1396 1918 1397 1919
rect 1471 1919 1477 1920
rect 1471 1918 1472 1919
rect 1396 1916 1472 1918
rect 1396 1915 1397 1916
rect 1391 1914 1397 1915
rect 1471 1915 1472 1916
rect 1476 1915 1477 1919
rect 1471 1914 1477 1915
rect 1559 1919 1565 1920
rect 1559 1915 1560 1919
rect 1564 1918 1565 1919
rect 1607 1919 1613 1920
rect 1607 1918 1608 1919
rect 1564 1916 1608 1918
rect 1564 1915 1565 1916
rect 1559 1914 1565 1915
rect 1607 1915 1608 1916
rect 1612 1915 1613 1919
rect 1607 1914 1613 1915
rect 1647 1919 1653 1920
rect 1647 1915 1648 1919
rect 1652 1918 1653 1919
rect 1702 1919 1708 1920
rect 1702 1918 1703 1919
rect 1652 1916 1703 1918
rect 1652 1915 1653 1916
rect 1647 1914 1653 1915
rect 1702 1915 1703 1916
rect 1707 1915 1708 1919
rect 1702 1914 1708 1915
rect 1734 1919 1741 1920
rect 1734 1915 1735 1919
rect 1740 1915 1741 1919
rect 1734 1914 1741 1915
rect 1815 1919 1821 1920
rect 1815 1915 1816 1919
rect 1820 1918 1821 1919
rect 1854 1919 1860 1920
rect 1854 1918 1855 1919
rect 1820 1916 1855 1918
rect 1820 1915 1821 1916
rect 1815 1914 1821 1915
rect 1854 1915 1855 1916
rect 1859 1915 1860 1919
rect 1854 1914 1860 1915
rect 1887 1919 1893 1920
rect 1887 1915 1888 1919
rect 1892 1918 1893 1919
rect 1926 1919 1932 1920
rect 1926 1918 1927 1919
rect 1892 1916 1927 1918
rect 1892 1915 1893 1916
rect 1887 1914 1893 1915
rect 1926 1915 1927 1916
rect 1931 1915 1932 1919
rect 1926 1914 1932 1915
rect 1959 1919 1968 1920
rect 1959 1915 1960 1919
rect 1967 1915 1968 1919
rect 2031 1919 2037 1920
rect 2031 1918 2032 1919
rect 1959 1914 1968 1915
rect 1999 1916 2032 1918
rect 174 1911 180 1912
rect 174 1907 175 1911
rect 179 1907 180 1911
rect 174 1906 180 1907
rect 214 1911 220 1912
rect 214 1907 215 1911
rect 219 1907 220 1911
rect 214 1906 220 1907
rect 262 1911 268 1912
rect 262 1907 263 1911
rect 267 1907 268 1911
rect 262 1906 268 1907
rect 318 1911 324 1912
rect 318 1907 319 1911
rect 323 1907 324 1911
rect 318 1906 324 1907
rect 390 1911 396 1912
rect 390 1907 391 1911
rect 395 1907 396 1911
rect 390 1906 396 1907
rect 470 1911 476 1912
rect 470 1907 471 1911
rect 475 1907 476 1911
rect 470 1906 476 1907
rect 550 1911 556 1912
rect 550 1907 551 1911
rect 555 1907 556 1911
rect 550 1906 556 1907
rect 638 1911 644 1912
rect 638 1907 639 1911
rect 643 1907 644 1911
rect 638 1906 644 1907
rect 718 1911 724 1912
rect 718 1907 719 1911
rect 723 1907 724 1911
rect 718 1906 724 1907
rect 798 1911 804 1912
rect 798 1907 799 1911
rect 803 1907 804 1911
rect 798 1906 804 1907
rect 878 1911 884 1912
rect 878 1907 879 1911
rect 883 1907 884 1911
rect 878 1906 884 1907
rect 958 1911 964 1912
rect 958 1907 959 1911
rect 963 1907 964 1911
rect 958 1906 964 1907
rect 1038 1911 1044 1912
rect 1038 1907 1039 1911
rect 1043 1907 1044 1911
rect 1038 1906 1044 1907
rect 1118 1911 1124 1912
rect 1278 1911 1284 1912
rect 1798 1911 1804 1912
rect 1118 1907 1119 1911
rect 1123 1907 1124 1911
rect 1118 1906 1124 1907
rect 1798 1907 1799 1911
rect 1803 1910 1804 1911
rect 1999 1910 2001 1916
rect 2031 1915 2032 1916
rect 2036 1915 2037 1919
rect 2031 1914 2037 1915
rect 2103 1919 2109 1920
rect 2103 1915 2104 1919
rect 2108 1918 2109 1919
rect 2142 1919 2148 1920
rect 2142 1918 2143 1919
rect 2108 1916 2143 1918
rect 2108 1915 2109 1916
rect 2103 1914 2109 1915
rect 2142 1915 2143 1916
rect 2147 1915 2148 1919
rect 2175 1919 2181 1920
rect 2175 1918 2176 1919
rect 2142 1914 2148 1915
rect 2152 1916 2176 1918
rect 1803 1908 2001 1910
rect 2014 1911 2020 1912
rect 1803 1907 1804 1908
rect 1798 1906 1804 1907
rect 2014 1907 2015 1911
rect 2019 1910 2020 1911
rect 2152 1910 2154 1916
rect 2175 1915 2176 1916
rect 2180 1915 2181 1919
rect 2175 1914 2181 1915
rect 2247 1919 2253 1920
rect 2247 1915 2248 1919
rect 2252 1918 2253 1919
rect 2294 1919 2300 1920
rect 2294 1918 2295 1919
rect 2252 1916 2295 1918
rect 2252 1915 2253 1916
rect 2247 1914 2253 1915
rect 2294 1915 2295 1916
rect 2299 1915 2300 1919
rect 2294 1914 2300 1915
rect 2327 1919 2333 1920
rect 2327 1915 2328 1919
rect 2332 1918 2333 1919
rect 2350 1919 2356 1920
rect 2350 1918 2351 1919
rect 2332 1916 2351 1918
rect 2332 1915 2333 1916
rect 2327 1914 2333 1915
rect 2350 1915 2351 1916
rect 2355 1915 2356 1919
rect 2350 1914 2356 1915
rect 2382 1919 2389 1920
rect 2382 1915 2383 1919
rect 2388 1915 2389 1919
rect 2382 1914 2389 1915
rect 2406 1916 2412 1917
rect 2406 1912 2407 1916
rect 2411 1912 2412 1916
rect 2406 1911 2412 1912
rect 2019 1908 2154 1910
rect 2019 1907 2020 1908
rect 2014 1906 2020 1907
rect 1302 1893 1308 1894
rect 190 1891 196 1892
rect 110 1888 116 1889
rect 110 1884 111 1888
rect 115 1884 116 1888
rect 190 1887 191 1891
rect 195 1890 196 1891
rect 455 1891 461 1892
rect 195 1888 346 1890
rect 195 1887 196 1888
rect 190 1886 196 1887
rect 344 1884 346 1888
rect 455 1887 456 1891
rect 460 1890 461 1891
rect 460 1888 510 1890
rect 1302 1889 1303 1893
rect 1307 1889 1308 1893
rect 460 1887 461 1888
rect 455 1886 461 1887
rect 110 1883 116 1884
rect 198 1883 205 1884
rect 198 1879 199 1883
rect 204 1879 205 1883
rect 198 1878 205 1879
rect 239 1883 245 1884
rect 239 1879 240 1883
rect 244 1882 245 1883
rect 247 1883 253 1884
rect 247 1882 248 1883
rect 244 1880 248 1882
rect 244 1879 245 1880
rect 239 1878 245 1879
rect 247 1879 248 1880
rect 252 1879 253 1883
rect 247 1878 253 1879
rect 287 1883 293 1884
rect 287 1879 288 1883
rect 292 1882 293 1883
rect 334 1883 340 1884
rect 334 1882 335 1883
rect 292 1880 335 1882
rect 292 1879 293 1880
rect 287 1878 293 1879
rect 334 1879 335 1880
rect 339 1879 340 1883
rect 334 1878 340 1879
rect 343 1883 349 1884
rect 343 1879 344 1883
rect 348 1879 349 1883
rect 343 1878 349 1879
rect 378 1883 384 1884
rect 378 1879 379 1883
rect 383 1882 384 1883
rect 415 1883 421 1884
rect 415 1882 416 1883
rect 383 1880 416 1882
rect 383 1879 384 1880
rect 378 1878 384 1879
rect 415 1879 416 1880
rect 420 1879 421 1883
rect 415 1878 421 1879
rect 495 1883 504 1884
rect 495 1879 496 1883
rect 503 1879 504 1883
rect 508 1882 510 1888
rect 1238 1888 1244 1889
rect 1302 1888 1308 1889
rect 1358 1893 1364 1894
rect 1358 1889 1359 1893
rect 1363 1889 1364 1893
rect 1358 1888 1364 1889
rect 1446 1893 1452 1894
rect 1446 1889 1447 1893
rect 1451 1889 1452 1893
rect 1446 1888 1452 1889
rect 1534 1893 1540 1894
rect 1534 1889 1535 1893
rect 1539 1889 1540 1893
rect 1534 1888 1540 1889
rect 1622 1893 1628 1894
rect 1622 1889 1623 1893
rect 1627 1889 1628 1893
rect 1622 1888 1628 1889
rect 1710 1893 1716 1894
rect 1710 1889 1711 1893
rect 1715 1889 1716 1893
rect 1710 1888 1716 1889
rect 1790 1893 1796 1894
rect 1790 1889 1791 1893
rect 1795 1889 1796 1893
rect 1790 1888 1796 1889
rect 1862 1893 1868 1894
rect 1862 1889 1863 1893
rect 1867 1889 1868 1893
rect 1862 1888 1868 1889
rect 1934 1893 1940 1894
rect 1934 1889 1935 1893
rect 1939 1889 1940 1893
rect 1934 1888 1940 1889
rect 2006 1893 2012 1894
rect 2006 1889 2007 1893
rect 2011 1889 2012 1893
rect 2006 1888 2012 1889
rect 2078 1893 2084 1894
rect 2078 1889 2079 1893
rect 2083 1889 2084 1893
rect 2078 1888 2084 1889
rect 2150 1893 2156 1894
rect 2150 1889 2151 1893
rect 2155 1889 2156 1893
rect 2150 1888 2156 1889
rect 2222 1893 2228 1894
rect 2222 1889 2223 1893
rect 2227 1889 2228 1893
rect 2222 1888 2228 1889
rect 2302 1893 2308 1894
rect 2302 1889 2303 1893
rect 2307 1889 2308 1893
rect 2302 1888 2308 1889
rect 2358 1893 2364 1894
rect 2358 1889 2359 1893
rect 2363 1889 2364 1893
rect 2358 1888 2364 1889
rect 1238 1884 1239 1888
rect 1243 1884 1244 1888
rect 575 1883 581 1884
rect 575 1882 576 1883
rect 508 1880 576 1882
rect 495 1878 504 1879
rect 575 1879 576 1880
rect 580 1879 581 1883
rect 575 1878 581 1879
rect 663 1883 669 1884
rect 663 1879 664 1883
rect 668 1882 669 1883
rect 671 1883 677 1884
rect 671 1882 672 1883
rect 668 1880 672 1882
rect 668 1879 669 1880
rect 663 1878 669 1879
rect 671 1879 672 1880
rect 676 1879 677 1883
rect 671 1878 677 1879
rect 743 1883 752 1884
rect 743 1879 744 1883
rect 751 1879 752 1883
rect 743 1878 752 1879
rect 822 1883 829 1884
rect 822 1879 823 1883
rect 828 1879 829 1883
rect 822 1878 829 1879
rect 902 1883 909 1884
rect 902 1879 903 1883
rect 908 1879 909 1883
rect 902 1878 909 1879
rect 983 1883 992 1884
rect 983 1879 984 1883
rect 991 1879 992 1883
rect 983 1878 992 1879
rect 1063 1883 1072 1884
rect 1063 1879 1064 1883
rect 1071 1879 1072 1883
rect 1143 1883 1149 1884
rect 1238 1883 1244 1884
rect 1299 1883 1305 1884
rect 1143 1882 1144 1883
rect 1063 1878 1072 1879
rect 1080 1880 1144 1882
rect 918 1875 924 1876
rect 110 1871 116 1872
rect 110 1867 111 1871
rect 115 1867 116 1871
rect 918 1871 919 1875
rect 923 1874 924 1875
rect 1080 1874 1082 1880
rect 1143 1879 1144 1880
rect 1148 1879 1149 1883
rect 1143 1878 1149 1879
rect 1299 1879 1300 1883
rect 1304 1882 1305 1883
rect 1335 1883 1341 1884
rect 1335 1882 1336 1883
rect 1304 1880 1336 1882
rect 1304 1879 1305 1880
rect 1299 1878 1305 1879
rect 1335 1879 1336 1880
rect 1340 1879 1341 1883
rect 1335 1878 1341 1879
rect 1355 1883 1361 1884
rect 1355 1879 1356 1883
rect 1360 1882 1361 1883
rect 1391 1883 1397 1884
rect 1391 1882 1392 1883
rect 1360 1880 1392 1882
rect 1360 1879 1361 1880
rect 1355 1878 1361 1879
rect 1391 1879 1392 1880
rect 1396 1879 1397 1883
rect 1391 1878 1397 1879
rect 1438 1883 1449 1884
rect 1438 1879 1439 1883
rect 1443 1879 1444 1883
rect 1448 1879 1449 1883
rect 1438 1878 1449 1879
rect 1522 1883 1528 1884
rect 1522 1879 1523 1883
rect 1527 1882 1528 1883
rect 1531 1883 1537 1884
rect 1531 1882 1532 1883
rect 1527 1880 1532 1882
rect 1527 1879 1528 1880
rect 1522 1878 1528 1879
rect 1531 1879 1532 1880
rect 1536 1879 1537 1883
rect 1531 1878 1537 1879
rect 1607 1883 1613 1884
rect 1607 1879 1608 1883
rect 1612 1882 1613 1883
rect 1619 1883 1625 1884
rect 1619 1882 1620 1883
rect 1612 1880 1620 1882
rect 1612 1879 1613 1880
rect 1607 1878 1613 1879
rect 1619 1879 1620 1880
rect 1624 1879 1625 1883
rect 1619 1878 1625 1879
rect 1702 1883 1713 1884
rect 1702 1879 1703 1883
rect 1707 1879 1708 1883
rect 1712 1879 1713 1883
rect 1702 1878 1713 1879
rect 1787 1883 1793 1884
rect 1787 1879 1788 1883
rect 1792 1882 1793 1883
rect 1798 1883 1804 1884
rect 1798 1882 1799 1883
rect 1792 1880 1799 1882
rect 1792 1879 1793 1880
rect 1787 1878 1793 1879
rect 1798 1879 1799 1880
rect 1803 1879 1804 1883
rect 1798 1878 1804 1879
rect 1854 1883 1865 1884
rect 1854 1879 1855 1883
rect 1859 1879 1860 1883
rect 1864 1879 1865 1883
rect 1854 1878 1865 1879
rect 1926 1883 1937 1884
rect 1926 1879 1927 1883
rect 1931 1879 1932 1883
rect 1936 1879 1937 1883
rect 1926 1878 1937 1879
rect 2003 1883 2009 1884
rect 2003 1879 2004 1883
rect 2008 1882 2009 1883
rect 2014 1883 2020 1884
rect 2014 1882 2015 1883
rect 2008 1880 2015 1882
rect 2008 1879 2009 1880
rect 2003 1878 2009 1879
rect 2014 1879 2015 1880
rect 2019 1879 2020 1883
rect 2014 1878 2020 1879
rect 2063 1883 2069 1884
rect 2063 1879 2064 1883
rect 2068 1882 2069 1883
rect 2075 1883 2081 1884
rect 2075 1882 2076 1883
rect 2068 1880 2076 1882
rect 2068 1879 2069 1880
rect 2063 1878 2069 1879
rect 2075 1879 2076 1880
rect 2080 1879 2081 1883
rect 2075 1878 2081 1879
rect 2142 1883 2153 1884
rect 2142 1879 2143 1883
rect 2147 1879 2148 1883
rect 2152 1879 2153 1883
rect 2142 1878 2153 1879
rect 2219 1883 2225 1884
rect 2219 1879 2220 1883
rect 2224 1882 2225 1883
rect 2230 1883 2236 1884
rect 2230 1882 2231 1883
rect 2224 1880 2231 1882
rect 2224 1879 2225 1880
rect 2219 1878 2225 1879
rect 2230 1879 2231 1880
rect 2235 1879 2236 1883
rect 2230 1878 2236 1879
rect 2294 1883 2305 1884
rect 2294 1879 2295 1883
rect 2299 1879 2300 1883
rect 2304 1879 2305 1883
rect 2294 1878 2305 1879
rect 2355 1883 2361 1884
rect 2355 1879 2356 1883
rect 2360 1882 2361 1883
rect 2382 1883 2388 1884
rect 2382 1882 2383 1883
rect 2360 1880 2383 1882
rect 2360 1879 2361 1880
rect 2355 1878 2361 1879
rect 2382 1879 2383 1880
rect 2387 1879 2388 1883
rect 2382 1878 2388 1879
rect 923 1872 1082 1874
rect 923 1871 924 1872
rect 918 1870 924 1871
rect 1238 1871 1244 1872
rect 110 1866 116 1867
rect 1238 1867 1239 1871
rect 1243 1867 1244 1871
rect 1238 1866 1244 1867
rect 1307 1871 1313 1872
rect 1307 1867 1308 1871
rect 1312 1870 1313 1871
rect 1330 1871 1336 1872
rect 1330 1870 1331 1871
rect 1312 1868 1331 1870
rect 1312 1867 1313 1868
rect 1307 1866 1313 1867
rect 1330 1867 1331 1868
rect 1335 1867 1336 1871
rect 1330 1866 1336 1867
rect 1338 1871 1344 1872
rect 1338 1867 1339 1871
rect 1343 1870 1344 1871
rect 1355 1871 1361 1872
rect 1355 1870 1356 1871
rect 1343 1868 1356 1870
rect 1343 1867 1344 1868
rect 1338 1866 1344 1867
rect 1355 1867 1356 1868
rect 1360 1867 1361 1871
rect 1355 1866 1361 1867
rect 1386 1871 1392 1872
rect 1386 1867 1387 1871
rect 1391 1870 1392 1871
rect 1411 1871 1417 1872
rect 1411 1870 1412 1871
rect 1391 1868 1412 1870
rect 1391 1867 1392 1868
rect 1386 1866 1392 1867
rect 1411 1867 1412 1868
rect 1416 1867 1417 1871
rect 1411 1866 1417 1867
rect 1475 1871 1481 1872
rect 1475 1867 1476 1871
rect 1480 1870 1481 1871
rect 1527 1871 1533 1872
rect 1527 1870 1528 1871
rect 1480 1868 1528 1870
rect 1480 1867 1481 1868
rect 1475 1866 1481 1867
rect 1527 1867 1528 1868
rect 1532 1867 1533 1871
rect 1527 1866 1533 1867
rect 1539 1871 1545 1872
rect 1539 1867 1540 1871
rect 1544 1870 1545 1871
rect 1598 1871 1604 1872
rect 1598 1870 1599 1871
rect 1544 1868 1599 1870
rect 1544 1867 1545 1868
rect 1539 1866 1545 1867
rect 1598 1867 1599 1868
rect 1603 1867 1604 1871
rect 1598 1866 1604 1867
rect 1606 1871 1617 1872
rect 1606 1867 1607 1871
rect 1611 1867 1612 1871
rect 1616 1867 1617 1871
rect 1606 1866 1617 1867
rect 1683 1871 1689 1872
rect 1683 1867 1684 1871
rect 1688 1870 1689 1871
rect 1754 1871 1760 1872
rect 1754 1870 1755 1871
rect 1688 1868 1755 1870
rect 1688 1867 1689 1868
rect 1683 1866 1689 1867
rect 1754 1867 1755 1868
rect 1759 1867 1760 1871
rect 1754 1866 1760 1867
rect 1763 1871 1769 1872
rect 1763 1867 1764 1871
rect 1768 1870 1769 1871
rect 1850 1871 1856 1872
rect 1850 1870 1851 1871
rect 1768 1868 1851 1870
rect 1768 1867 1769 1868
rect 1763 1866 1769 1867
rect 1850 1867 1851 1868
rect 1855 1867 1856 1871
rect 1850 1866 1856 1867
rect 1859 1871 1865 1872
rect 1859 1867 1860 1871
rect 1864 1870 1865 1871
rect 1927 1871 1933 1872
rect 1927 1870 1928 1871
rect 1864 1868 1928 1870
rect 1864 1867 1865 1868
rect 1859 1866 1865 1867
rect 1927 1867 1928 1868
rect 1932 1867 1933 1871
rect 1927 1866 1933 1867
rect 1962 1871 1968 1872
rect 1962 1867 1963 1871
rect 1967 1870 1968 1871
rect 1971 1871 1977 1872
rect 1971 1870 1972 1871
rect 1967 1868 1972 1870
rect 1967 1867 1968 1868
rect 1962 1866 1968 1867
rect 1971 1867 1972 1868
rect 1976 1867 1977 1871
rect 1971 1866 1977 1867
rect 2007 1871 2013 1872
rect 2007 1867 2008 1871
rect 2012 1870 2013 1871
rect 2091 1871 2097 1872
rect 2091 1870 2092 1871
rect 2012 1868 2092 1870
rect 2012 1867 2013 1868
rect 2007 1866 2013 1867
rect 2091 1867 2092 1868
rect 2096 1867 2097 1871
rect 2091 1866 2097 1867
rect 2122 1871 2128 1872
rect 2122 1867 2123 1871
rect 2127 1870 2128 1871
rect 2219 1871 2225 1872
rect 2219 1870 2220 1871
rect 2127 1868 2220 1870
rect 2127 1867 2128 1868
rect 2122 1866 2128 1867
rect 2219 1867 2220 1868
rect 2224 1867 2225 1871
rect 2219 1866 2225 1867
rect 2350 1871 2361 1872
rect 2350 1867 2351 1871
rect 2355 1867 2356 1871
rect 2360 1867 2361 1871
rect 2350 1866 2361 1867
rect 174 1864 180 1865
rect 174 1860 175 1864
rect 179 1860 180 1864
rect 174 1859 180 1860
rect 214 1864 220 1865
rect 214 1860 215 1864
rect 219 1860 220 1864
rect 214 1859 220 1860
rect 262 1864 268 1865
rect 262 1860 263 1864
rect 267 1860 268 1864
rect 262 1859 268 1860
rect 318 1864 324 1865
rect 318 1860 319 1864
rect 323 1860 324 1864
rect 318 1859 324 1860
rect 390 1864 396 1865
rect 390 1860 391 1864
rect 395 1860 396 1864
rect 390 1859 396 1860
rect 470 1864 476 1865
rect 470 1860 471 1864
rect 475 1860 476 1864
rect 470 1859 476 1860
rect 550 1864 556 1865
rect 550 1860 551 1864
rect 555 1860 556 1864
rect 550 1859 556 1860
rect 638 1864 644 1865
rect 638 1860 639 1864
rect 643 1860 644 1864
rect 638 1859 644 1860
rect 718 1864 724 1865
rect 718 1860 719 1864
rect 723 1860 724 1864
rect 718 1859 724 1860
rect 798 1864 804 1865
rect 798 1860 799 1864
rect 803 1860 804 1864
rect 798 1859 804 1860
rect 878 1864 884 1865
rect 878 1860 879 1864
rect 883 1860 884 1864
rect 878 1859 884 1860
rect 958 1864 964 1865
rect 958 1860 959 1864
rect 963 1860 964 1864
rect 958 1859 964 1860
rect 1038 1864 1044 1865
rect 1038 1860 1039 1864
rect 1043 1860 1044 1864
rect 1038 1859 1044 1860
rect 1118 1864 1124 1865
rect 1118 1860 1119 1864
rect 1123 1860 1124 1864
rect 1118 1859 1124 1860
rect 1310 1863 1316 1864
rect 1310 1859 1311 1863
rect 1315 1859 1316 1863
rect 1310 1858 1316 1859
rect 1358 1863 1364 1864
rect 1358 1859 1359 1863
rect 1363 1859 1364 1863
rect 1358 1858 1364 1859
rect 1414 1863 1420 1864
rect 1414 1859 1415 1863
rect 1419 1859 1420 1863
rect 1414 1858 1420 1859
rect 1478 1863 1484 1864
rect 1478 1859 1479 1863
rect 1483 1859 1484 1863
rect 1478 1858 1484 1859
rect 1542 1863 1548 1864
rect 1542 1859 1543 1863
rect 1547 1859 1548 1863
rect 1542 1858 1548 1859
rect 1614 1863 1620 1864
rect 1614 1859 1615 1863
rect 1619 1859 1620 1863
rect 1614 1858 1620 1859
rect 1686 1863 1692 1864
rect 1686 1859 1687 1863
rect 1691 1859 1692 1863
rect 1686 1858 1692 1859
rect 1766 1863 1772 1864
rect 1766 1859 1767 1863
rect 1771 1859 1772 1863
rect 1766 1858 1772 1859
rect 1862 1863 1868 1864
rect 1862 1859 1863 1863
rect 1867 1859 1868 1863
rect 1862 1858 1868 1859
rect 1974 1863 1980 1864
rect 1974 1859 1975 1863
rect 1979 1859 1980 1863
rect 1974 1858 1980 1859
rect 2094 1863 2100 1864
rect 2094 1859 2095 1863
rect 2099 1859 2100 1863
rect 2094 1858 2100 1859
rect 2222 1863 2228 1864
rect 2222 1859 2223 1863
rect 2227 1859 2228 1863
rect 2222 1858 2228 1859
rect 2358 1863 2364 1864
rect 2358 1859 2359 1863
rect 2363 1859 2364 1863
rect 2358 1858 2364 1859
rect 134 1844 140 1845
rect 134 1840 135 1844
rect 139 1840 140 1844
rect 134 1839 140 1840
rect 174 1844 180 1845
rect 174 1840 175 1844
rect 179 1840 180 1844
rect 174 1839 180 1840
rect 214 1844 220 1845
rect 214 1840 215 1844
rect 219 1840 220 1844
rect 214 1839 220 1840
rect 270 1844 276 1845
rect 270 1840 271 1844
rect 275 1840 276 1844
rect 270 1839 276 1840
rect 350 1844 356 1845
rect 350 1840 351 1844
rect 355 1840 356 1844
rect 350 1839 356 1840
rect 438 1844 444 1845
rect 438 1840 439 1844
rect 443 1840 444 1844
rect 438 1839 444 1840
rect 534 1844 540 1845
rect 534 1840 535 1844
rect 539 1840 540 1844
rect 534 1839 540 1840
rect 630 1844 636 1845
rect 630 1840 631 1844
rect 635 1840 636 1844
rect 630 1839 636 1840
rect 726 1844 732 1845
rect 726 1840 727 1844
rect 731 1840 732 1844
rect 726 1839 732 1840
rect 822 1844 828 1845
rect 822 1840 823 1844
rect 827 1840 828 1844
rect 822 1839 828 1840
rect 910 1844 916 1845
rect 910 1840 911 1844
rect 915 1840 916 1844
rect 910 1839 916 1840
rect 990 1844 996 1845
rect 990 1840 991 1844
rect 995 1840 996 1844
rect 990 1839 996 1840
rect 1062 1844 1068 1845
rect 1062 1840 1063 1844
rect 1067 1840 1068 1844
rect 1062 1839 1068 1840
rect 1134 1844 1140 1845
rect 1134 1840 1135 1844
rect 1139 1840 1140 1844
rect 1134 1839 1140 1840
rect 1190 1844 1196 1845
rect 1190 1840 1191 1844
rect 1195 1840 1196 1844
rect 1330 1843 1336 1844
rect 1190 1839 1196 1840
rect 1278 1840 1284 1841
rect 110 1837 116 1838
rect 110 1833 111 1837
rect 115 1833 116 1837
rect 110 1832 116 1833
rect 1238 1837 1244 1838
rect 1238 1833 1239 1837
rect 1243 1833 1244 1837
rect 1278 1836 1279 1840
rect 1283 1836 1284 1840
rect 1330 1839 1331 1843
rect 1335 1842 1336 1843
rect 1927 1843 1933 1844
rect 1335 1840 1450 1842
rect 1335 1839 1336 1840
rect 1330 1838 1336 1839
rect 1278 1835 1284 1836
rect 1335 1835 1344 1836
rect 1238 1832 1244 1833
rect 1335 1831 1336 1835
rect 1343 1831 1344 1835
rect 1335 1830 1344 1831
rect 1383 1835 1392 1836
rect 1383 1831 1384 1835
rect 1391 1831 1392 1835
rect 1383 1830 1392 1831
rect 1438 1835 1445 1836
rect 1438 1831 1439 1835
rect 1444 1831 1445 1835
rect 1448 1834 1450 1840
rect 1927 1839 1928 1843
rect 1932 1842 1933 1843
rect 1932 1840 2134 1842
rect 1932 1839 1933 1840
rect 1927 1838 1933 1839
rect 1503 1835 1509 1836
rect 1503 1834 1504 1835
rect 1448 1832 1504 1834
rect 1438 1830 1445 1831
rect 1503 1831 1504 1832
rect 1508 1831 1509 1835
rect 1503 1830 1509 1831
rect 1527 1835 1533 1836
rect 1527 1831 1528 1835
rect 1532 1834 1533 1835
rect 1567 1835 1573 1836
rect 1567 1834 1568 1835
rect 1532 1832 1568 1834
rect 1532 1831 1533 1832
rect 1527 1830 1533 1831
rect 1567 1831 1568 1832
rect 1572 1831 1573 1835
rect 1567 1830 1573 1831
rect 1598 1835 1604 1836
rect 1598 1831 1599 1835
rect 1603 1834 1604 1835
rect 1639 1835 1645 1836
rect 1639 1834 1640 1835
rect 1603 1832 1640 1834
rect 1603 1831 1604 1832
rect 1598 1830 1604 1831
rect 1639 1831 1640 1832
rect 1644 1831 1645 1835
rect 1639 1830 1645 1831
rect 1670 1835 1676 1836
rect 1670 1831 1671 1835
rect 1675 1834 1676 1835
rect 1711 1835 1717 1836
rect 1711 1834 1712 1835
rect 1675 1832 1712 1834
rect 1675 1831 1676 1832
rect 1670 1830 1676 1831
rect 1711 1831 1712 1832
rect 1716 1831 1717 1835
rect 1711 1830 1717 1831
rect 1754 1835 1760 1836
rect 1754 1831 1755 1835
rect 1759 1834 1760 1835
rect 1791 1835 1797 1836
rect 1791 1834 1792 1835
rect 1759 1832 1792 1834
rect 1759 1831 1760 1832
rect 1754 1830 1760 1831
rect 1791 1831 1792 1832
rect 1796 1831 1797 1835
rect 1791 1830 1797 1831
rect 1850 1835 1856 1836
rect 1850 1831 1851 1835
rect 1855 1834 1856 1835
rect 1887 1835 1893 1836
rect 1887 1834 1888 1835
rect 1855 1832 1888 1834
rect 1855 1831 1856 1832
rect 1850 1830 1856 1831
rect 1887 1831 1888 1832
rect 1892 1831 1893 1835
rect 1887 1830 1893 1831
rect 1999 1835 2005 1836
rect 1999 1831 2000 1835
rect 2004 1834 2005 1835
rect 2007 1835 2013 1836
rect 2007 1834 2008 1835
rect 2004 1832 2008 1834
rect 2004 1831 2005 1832
rect 1999 1830 2005 1831
rect 2007 1831 2008 1832
rect 2012 1831 2013 1835
rect 2007 1830 2013 1831
rect 2119 1835 2128 1836
rect 2119 1831 2120 1835
rect 2127 1831 2128 1835
rect 2132 1834 2134 1840
rect 2406 1840 2412 1841
rect 2406 1836 2407 1840
rect 2411 1836 2412 1840
rect 2247 1835 2253 1836
rect 2247 1834 2248 1835
rect 2132 1832 2248 1834
rect 2119 1830 2128 1831
rect 2247 1831 2248 1832
rect 2252 1831 2253 1835
rect 2247 1830 2253 1831
rect 2382 1835 2389 1836
rect 2406 1835 2412 1836
rect 2382 1831 2383 1835
rect 2388 1831 2389 1835
rect 2382 1830 2389 1831
rect 142 1823 148 1824
rect 110 1820 116 1821
rect 110 1816 111 1820
rect 115 1816 116 1820
rect 142 1819 143 1823
rect 147 1822 148 1823
rect 159 1823 165 1824
rect 159 1822 160 1823
rect 147 1820 160 1822
rect 147 1819 148 1820
rect 142 1818 148 1819
rect 159 1819 160 1820
rect 164 1819 165 1823
rect 199 1823 205 1824
rect 199 1822 200 1823
rect 159 1818 165 1819
rect 168 1820 200 1822
rect 110 1815 116 1816
rect 150 1815 156 1816
rect 150 1811 151 1815
rect 155 1814 156 1815
rect 168 1814 170 1820
rect 199 1819 200 1820
rect 204 1819 205 1823
rect 239 1823 245 1824
rect 239 1822 240 1823
rect 199 1818 205 1819
rect 208 1820 240 1822
rect 155 1812 170 1814
rect 182 1815 188 1816
rect 155 1811 156 1812
rect 150 1810 156 1811
rect 182 1811 183 1815
rect 187 1814 188 1815
rect 208 1814 210 1820
rect 239 1819 240 1820
rect 244 1819 245 1823
rect 239 1818 245 1819
rect 247 1823 253 1824
rect 247 1819 248 1823
rect 252 1822 253 1823
rect 295 1823 301 1824
rect 295 1822 296 1823
rect 252 1820 296 1822
rect 252 1819 253 1820
rect 247 1818 253 1819
rect 295 1819 296 1820
rect 300 1819 301 1823
rect 295 1818 301 1819
rect 375 1823 381 1824
rect 375 1819 376 1823
rect 380 1822 381 1823
rect 430 1823 436 1824
rect 430 1822 431 1823
rect 380 1820 431 1822
rect 380 1819 381 1820
rect 375 1818 381 1819
rect 430 1819 431 1820
rect 435 1819 436 1823
rect 430 1818 436 1819
rect 463 1823 469 1824
rect 463 1819 464 1823
rect 468 1822 469 1823
rect 526 1823 532 1824
rect 526 1822 527 1823
rect 468 1820 527 1822
rect 468 1819 469 1820
rect 463 1818 469 1819
rect 526 1819 527 1820
rect 531 1819 532 1823
rect 559 1823 565 1824
rect 559 1822 560 1823
rect 526 1818 532 1819
rect 536 1820 560 1822
rect 187 1812 210 1814
rect 294 1815 300 1816
rect 187 1811 188 1812
rect 182 1810 188 1811
rect 294 1811 295 1815
rect 299 1814 300 1815
rect 536 1814 538 1820
rect 559 1819 560 1820
rect 564 1819 565 1823
rect 559 1818 565 1819
rect 654 1823 661 1824
rect 654 1819 655 1823
rect 660 1819 661 1823
rect 654 1818 661 1819
rect 663 1823 669 1824
rect 663 1819 664 1823
rect 668 1822 669 1823
rect 751 1823 757 1824
rect 751 1822 752 1823
rect 668 1820 752 1822
rect 668 1819 669 1820
rect 663 1818 669 1819
rect 751 1819 752 1820
rect 756 1819 757 1823
rect 751 1818 757 1819
rect 759 1823 765 1824
rect 759 1819 760 1823
rect 764 1822 765 1823
rect 847 1823 853 1824
rect 847 1822 848 1823
rect 764 1820 848 1822
rect 764 1819 765 1820
rect 759 1818 765 1819
rect 847 1819 848 1820
rect 852 1819 853 1823
rect 847 1818 853 1819
rect 935 1823 941 1824
rect 935 1819 936 1823
rect 940 1822 941 1823
rect 982 1823 988 1824
rect 982 1822 983 1823
rect 940 1820 983 1822
rect 940 1819 941 1820
rect 935 1818 941 1819
rect 982 1819 983 1820
rect 987 1819 988 1823
rect 982 1818 988 1819
rect 1015 1823 1021 1824
rect 1015 1819 1016 1823
rect 1020 1822 1021 1823
rect 1054 1823 1060 1824
rect 1054 1822 1055 1823
rect 1020 1820 1055 1822
rect 1020 1819 1021 1820
rect 1015 1818 1021 1819
rect 1054 1819 1055 1820
rect 1059 1819 1060 1823
rect 1054 1818 1060 1819
rect 1087 1823 1093 1824
rect 1087 1819 1088 1823
rect 1092 1822 1093 1823
rect 1126 1823 1132 1824
rect 1126 1822 1127 1823
rect 1092 1820 1127 1822
rect 1092 1819 1093 1820
rect 1087 1818 1093 1819
rect 1126 1819 1127 1820
rect 1131 1819 1132 1823
rect 1126 1818 1132 1819
rect 1159 1823 1165 1824
rect 1159 1819 1160 1823
rect 1164 1822 1165 1823
rect 1182 1823 1188 1824
rect 1182 1822 1183 1823
rect 1164 1820 1183 1822
rect 1164 1819 1165 1820
rect 1159 1818 1165 1819
rect 1182 1819 1183 1820
rect 1187 1819 1188 1823
rect 1215 1823 1221 1824
rect 1215 1822 1216 1823
rect 1182 1818 1188 1819
rect 1192 1820 1216 1822
rect 299 1812 538 1814
rect 1038 1815 1044 1816
rect 299 1811 300 1812
rect 294 1810 300 1811
rect 1038 1811 1039 1815
rect 1043 1814 1044 1815
rect 1192 1814 1194 1820
rect 1215 1819 1216 1820
rect 1220 1819 1221 1823
rect 1278 1823 1284 1824
rect 1215 1818 1221 1819
rect 1238 1820 1244 1821
rect 1238 1816 1239 1820
rect 1243 1816 1244 1820
rect 1278 1819 1279 1823
rect 1283 1819 1284 1823
rect 1278 1818 1284 1819
rect 2406 1823 2412 1824
rect 2406 1819 2407 1823
rect 2411 1819 2412 1823
rect 2406 1818 2412 1819
rect 1238 1815 1244 1816
rect 1310 1816 1316 1817
rect 1043 1812 1194 1814
rect 1310 1812 1311 1816
rect 1315 1812 1316 1816
rect 1043 1811 1044 1812
rect 1310 1811 1316 1812
rect 1358 1816 1364 1817
rect 1358 1812 1359 1816
rect 1363 1812 1364 1816
rect 1358 1811 1364 1812
rect 1414 1816 1420 1817
rect 1414 1812 1415 1816
rect 1419 1812 1420 1816
rect 1414 1811 1420 1812
rect 1478 1816 1484 1817
rect 1478 1812 1479 1816
rect 1483 1812 1484 1816
rect 1478 1811 1484 1812
rect 1542 1816 1548 1817
rect 1542 1812 1543 1816
rect 1547 1812 1548 1816
rect 1542 1811 1548 1812
rect 1614 1816 1620 1817
rect 1614 1812 1615 1816
rect 1619 1812 1620 1816
rect 1614 1811 1620 1812
rect 1686 1816 1692 1817
rect 1686 1812 1687 1816
rect 1691 1812 1692 1816
rect 1686 1811 1692 1812
rect 1766 1816 1772 1817
rect 1766 1812 1767 1816
rect 1771 1812 1772 1816
rect 1766 1811 1772 1812
rect 1862 1816 1868 1817
rect 1862 1812 1863 1816
rect 1867 1812 1868 1816
rect 1862 1811 1868 1812
rect 1974 1816 1980 1817
rect 1974 1812 1975 1816
rect 1979 1812 1980 1816
rect 1974 1811 1980 1812
rect 2094 1816 2100 1817
rect 2094 1812 2095 1816
rect 2099 1812 2100 1816
rect 2094 1811 2100 1812
rect 2222 1816 2228 1817
rect 2222 1812 2223 1816
rect 2227 1812 2228 1816
rect 2222 1811 2228 1812
rect 2358 1816 2364 1817
rect 2358 1812 2359 1816
rect 2363 1812 2364 1816
rect 2358 1811 2364 1812
rect 1038 1810 1044 1811
rect 1406 1800 1412 1801
rect 134 1797 140 1798
rect 134 1793 135 1797
rect 139 1793 140 1797
rect 134 1792 140 1793
rect 174 1797 180 1798
rect 174 1793 175 1797
rect 179 1793 180 1797
rect 174 1792 180 1793
rect 214 1797 220 1798
rect 214 1793 215 1797
rect 219 1793 220 1797
rect 214 1792 220 1793
rect 270 1797 276 1798
rect 270 1793 271 1797
rect 275 1793 276 1797
rect 270 1792 276 1793
rect 350 1797 356 1798
rect 350 1793 351 1797
rect 355 1793 356 1797
rect 350 1792 356 1793
rect 438 1797 444 1798
rect 438 1793 439 1797
rect 443 1793 444 1797
rect 438 1792 444 1793
rect 534 1797 540 1798
rect 534 1793 535 1797
rect 539 1793 540 1797
rect 534 1792 540 1793
rect 630 1797 636 1798
rect 630 1793 631 1797
rect 635 1793 636 1797
rect 630 1792 636 1793
rect 726 1797 732 1798
rect 726 1793 727 1797
rect 731 1793 732 1797
rect 726 1792 732 1793
rect 822 1797 828 1798
rect 822 1793 823 1797
rect 827 1793 828 1797
rect 822 1792 828 1793
rect 910 1797 916 1798
rect 910 1793 911 1797
rect 915 1793 916 1797
rect 910 1792 916 1793
rect 990 1797 996 1798
rect 990 1793 991 1797
rect 995 1793 996 1797
rect 990 1792 996 1793
rect 1062 1797 1068 1798
rect 1062 1793 1063 1797
rect 1067 1793 1068 1797
rect 1062 1792 1068 1793
rect 1134 1797 1140 1798
rect 1134 1793 1135 1797
rect 1139 1793 1140 1797
rect 1134 1792 1140 1793
rect 1190 1797 1196 1798
rect 1190 1793 1191 1797
rect 1195 1793 1196 1797
rect 1406 1796 1407 1800
rect 1411 1796 1412 1800
rect 1406 1795 1412 1796
rect 1470 1800 1476 1801
rect 1470 1796 1471 1800
rect 1475 1796 1476 1800
rect 1470 1795 1476 1796
rect 1534 1800 1540 1801
rect 1534 1796 1535 1800
rect 1539 1796 1540 1800
rect 1534 1795 1540 1796
rect 1598 1800 1604 1801
rect 1598 1796 1599 1800
rect 1603 1796 1604 1800
rect 1598 1795 1604 1796
rect 1662 1800 1668 1801
rect 1662 1796 1663 1800
rect 1667 1796 1668 1800
rect 1662 1795 1668 1796
rect 1726 1800 1732 1801
rect 1726 1796 1727 1800
rect 1731 1796 1732 1800
rect 1726 1795 1732 1796
rect 1782 1800 1788 1801
rect 1782 1796 1783 1800
rect 1787 1796 1788 1800
rect 1782 1795 1788 1796
rect 1838 1800 1844 1801
rect 1838 1796 1839 1800
rect 1843 1796 1844 1800
rect 1838 1795 1844 1796
rect 1894 1800 1900 1801
rect 1894 1796 1895 1800
rect 1899 1796 1900 1800
rect 1894 1795 1900 1796
rect 1958 1800 1964 1801
rect 1958 1796 1959 1800
rect 1963 1796 1964 1800
rect 1958 1795 1964 1796
rect 1190 1792 1196 1793
rect 1278 1793 1284 1794
rect 1278 1789 1279 1793
rect 1283 1789 1284 1793
rect 1278 1788 1284 1789
rect 2406 1793 2412 1794
rect 2406 1789 2407 1793
rect 2411 1789 2412 1793
rect 2406 1788 2412 1789
rect 131 1787 137 1788
rect 131 1783 132 1787
rect 136 1786 137 1787
rect 150 1787 156 1788
rect 150 1786 151 1787
rect 136 1784 151 1786
rect 136 1783 137 1784
rect 131 1782 137 1783
rect 150 1783 151 1784
rect 155 1783 156 1787
rect 150 1782 156 1783
rect 171 1787 177 1788
rect 171 1783 172 1787
rect 176 1786 177 1787
rect 182 1787 188 1788
rect 182 1786 183 1787
rect 176 1784 183 1786
rect 176 1783 177 1784
rect 171 1782 177 1783
rect 182 1783 183 1784
rect 187 1783 188 1787
rect 182 1782 188 1783
rect 211 1787 217 1788
rect 211 1783 212 1787
rect 216 1786 217 1787
rect 247 1787 253 1788
rect 247 1786 248 1787
rect 216 1784 248 1786
rect 216 1783 217 1784
rect 211 1782 217 1783
rect 247 1783 248 1784
rect 252 1783 253 1787
rect 247 1782 253 1783
rect 267 1787 273 1788
rect 267 1783 268 1787
rect 272 1786 273 1787
rect 294 1787 300 1788
rect 294 1786 295 1787
rect 272 1784 295 1786
rect 272 1783 273 1784
rect 267 1782 273 1783
rect 294 1783 295 1784
rect 299 1783 300 1787
rect 294 1782 300 1783
rect 334 1787 340 1788
rect 334 1783 335 1787
rect 339 1786 340 1787
rect 347 1787 353 1788
rect 347 1786 348 1787
rect 339 1784 348 1786
rect 339 1783 340 1784
rect 334 1782 340 1783
rect 347 1783 348 1784
rect 352 1783 353 1787
rect 347 1782 353 1783
rect 430 1787 441 1788
rect 430 1783 431 1787
rect 435 1783 436 1787
rect 440 1783 441 1787
rect 430 1782 441 1783
rect 526 1787 537 1788
rect 526 1783 527 1787
rect 531 1783 532 1787
rect 536 1783 537 1787
rect 526 1782 537 1783
rect 627 1787 633 1788
rect 627 1783 628 1787
rect 632 1786 633 1787
rect 663 1787 669 1788
rect 663 1786 664 1787
rect 632 1784 664 1786
rect 632 1783 633 1784
rect 627 1782 633 1783
rect 663 1783 664 1784
rect 668 1783 669 1787
rect 663 1782 669 1783
rect 723 1787 729 1788
rect 723 1783 724 1787
rect 728 1786 729 1787
rect 759 1787 765 1788
rect 759 1786 760 1787
rect 728 1784 760 1786
rect 728 1783 729 1784
rect 723 1782 729 1783
rect 759 1783 760 1784
rect 764 1783 765 1787
rect 759 1782 765 1783
rect 778 1787 784 1788
rect 778 1783 779 1787
rect 783 1786 784 1787
rect 819 1787 825 1788
rect 819 1786 820 1787
rect 783 1784 820 1786
rect 783 1783 784 1784
rect 778 1782 784 1783
rect 819 1783 820 1784
rect 824 1783 825 1787
rect 819 1782 825 1783
rect 907 1787 913 1788
rect 907 1783 908 1787
rect 912 1786 913 1787
rect 918 1787 924 1788
rect 918 1786 919 1787
rect 912 1784 919 1786
rect 912 1783 913 1784
rect 907 1782 913 1783
rect 918 1783 919 1784
rect 923 1783 924 1787
rect 918 1782 924 1783
rect 982 1787 993 1788
rect 982 1783 983 1787
rect 987 1783 988 1787
rect 992 1783 993 1787
rect 982 1782 993 1783
rect 1054 1787 1065 1788
rect 1054 1783 1055 1787
rect 1059 1783 1060 1787
rect 1064 1783 1065 1787
rect 1054 1782 1065 1783
rect 1126 1787 1137 1788
rect 1126 1783 1127 1787
rect 1131 1783 1132 1787
rect 1136 1783 1137 1787
rect 1126 1782 1137 1783
rect 1182 1787 1193 1788
rect 1182 1783 1183 1787
rect 1187 1783 1188 1787
rect 1192 1783 1193 1787
rect 1182 1782 1193 1783
rect 1431 1779 1437 1780
rect 1278 1776 1284 1777
rect 131 1775 137 1776
rect 131 1771 132 1775
rect 136 1774 137 1775
rect 142 1775 148 1776
rect 142 1774 143 1775
rect 136 1772 143 1774
rect 136 1771 137 1772
rect 131 1770 137 1771
rect 142 1771 143 1772
rect 147 1771 148 1775
rect 142 1770 148 1771
rect 158 1775 164 1776
rect 158 1771 159 1775
rect 163 1774 164 1775
rect 171 1775 177 1776
rect 171 1774 172 1775
rect 163 1772 172 1774
rect 163 1771 164 1772
rect 158 1770 164 1771
rect 171 1771 172 1772
rect 176 1771 177 1775
rect 171 1770 177 1771
rect 198 1775 204 1776
rect 198 1771 199 1775
rect 203 1774 204 1775
rect 211 1775 217 1776
rect 211 1774 212 1775
rect 203 1772 212 1774
rect 203 1771 204 1772
rect 198 1770 204 1771
rect 211 1771 212 1772
rect 216 1771 217 1775
rect 211 1770 217 1771
rect 242 1775 248 1776
rect 242 1771 243 1775
rect 247 1774 248 1775
rect 283 1775 289 1776
rect 283 1774 284 1775
rect 247 1772 284 1774
rect 247 1771 248 1772
rect 242 1770 248 1771
rect 283 1771 284 1772
rect 288 1771 289 1775
rect 283 1770 289 1771
rect 314 1775 320 1776
rect 314 1771 315 1775
rect 319 1774 320 1775
rect 371 1775 377 1776
rect 371 1774 372 1775
rect 319 1772 372 1774
rect 319 1771 320 1772
rect 314 1770 320 1771
rect 371 1771 372 1772
rect 376 1771 377 1775
rect 371 1770 377 1771
rect 402 1775 408 1776
rect 402 1771 403 1775
rect 407 1774 408 1775
rect 467 1775 473 1776
rect 467 1774 468 1775
rect 407 1772 468 1774
rect 407 1771 408 1772
rect 402 1770 408 1771
rect 467 1771 468 1772
rect 472 1771 473 1775
rect 467 1770 473 1771
rect 498 1775 504 1776
rect 498 1771 499 1775
rect 503 1774 504 1775
rect 563 1775 569 1776
rect 563 1774 564 1775
rect 503 1772 564 1774
rect 503 1771 504 1772
rect 498 1770 504 1771
rect 563 1771 564 1772
rect 568 1771 569 1775
rect 563 1770 569 1771
rect 659 1775 665 1776
rect 659 1771 660 1775
rect 664 1774 665 1775
rect 682 1775 688 1776
rect 682 1774 683 1775
rect 664 1772 683 1774
rect 664 1771 665 1772
rect 659 1770 665 1771
rect 682 1771 683 1772
rect 687 1771 688 1775
rect 682 1770 688 1771
rect 690 1775 696 1776
rect 690 1771 691 1775
rect 695 1774 696 1775
rect 747 1775 753 1776
rect 747 1774 748 1775
rect 695 1772 748 1774
rect 695 1771 696 1772
rect 690 1770 696 1771
rect 747 1771 748 1772
rect 752 1771 753 1775
rect 747 1770 753 1771
rect 827 1775 833 1776
rect 827 1771 828 1775
rect 832 1774 833 1775
rect 890 1775 896 1776
rect 890 1774 891 1775
rect 832 1772 891 1774
rect 832 1771 833 1772
rect 827 1770 833 1771
rect 890 1771 891 1772
rect 895 1771 896 1775
rect 890 1770 896 1771
rect 899 1775 905 1776
rect 899 1771 900 1775
rect 904 1774 905 1775
rect 954 1775 960 1776
rect 954 1774 955 1775
rect 904 1772 955 1774
rect 904 1771 905 1772
rect 899 1770 905 1771
rect 954 1771 955 1772
rect 959 1771 960 1775
rect 954 1770 960 1771
rect 963 1775 969 1776
rect 963 1771 964 1775
rect 968 1774 969 1775
rect 1006 1775 1012 1776
rect 1006 1774 1007 1775
rect 968 1772 1007 1774
rect 968 1771 969 1772
rect 963 1770 969 1771
rect 1006 1771 1007 1772
rect 1011 1771 1012 1775
rect 1006 1770 1012 1771
rect 1027 1775 1033 1776
rect 1027 1771 1028 1775
rect 1032 1774 1033 1775
rect 1038 1775 1044 1776
rect 1038 1774 1039 1775
rect 1032 1772 1039 1774
rect 1032 1771 1033 1772
rect 1027 1770 1033 1771
rect 1038 1771 1039 1772
rect 1043 1771 1044 1775
rect 1038 1770 1044 1771
rect 1063 1775 1069 1776
rect 1063 1771 1064 1775
rect 1068 1774 1069 1775
rect 1083 1775 1089 1776
rect 1083 1774 1084 1775
rect 1068 1772 1084 1774
rect 1068 1771 1069 1772
rect 1063 1770 1069 1771
rect 1083 1771 1084 1772
rect 1088 1771 1089 1775
rect 1083 1770 1089 1771
rect 1114 1775 1120 1776
rect 1114 1771 1115 1775
rect 1119 1774 1120 1775
rect 1147 1775 1153 1776
rect 1147 1774 1148 1775
rect 1119 1772 1148 1774
rect 1119 1771 1120 1772
rect 1114 1770 1120 1771
rect 1147 1771 1148 1772
rect 1152 1771 1153 1775
rect 1147 1770 1153 1771
rect 1174 1775 1180 1776
rect 1174 1771 1175 1775
rect 1179 1774 1180 1775
rect 1187 1775 1193 1776
rect 1187 1774 1188 1775
rect 1179 1772 1188 1774
rect 1179 1771 1180 1772
rect 1174 1770 1180 1771
rect 1187 1771 1188 1772
rect 1192 1771 1193 1775
rect 1278 1772 1279 1776
rect 1283 1772 1284 1776
rect 1431 1775 1432 1779
rect 1436 1778 1437 1779
rect 1462 1779 1468 1780
rect 1462 1778 1463 1779
rect 1436 1776 1463 1778
rect 1436 1775 1437 1776
rect 1431 1774 1437 1775
rect 1462 1775 1463 1776
rect 1467 1775 1468 1779
rect 1462 1774 1468 1775
rect 1495 1779 1501 1780
rect 1495 1775 1496 1779
rect 1500 1778 1501 1779
rect 1526 1779 1532 1780
rect 1526 1778 1527 1779
rect 1500 1776 1527 1778
rect 1500 1775 1501 1776
rect 1495 1774 1501 1775
rect 1526 1775 1527 1776
rect 1531 1775 1532 1779
rect 1526 1774 1532 1775
rect 1559 1779 1565 1780
rect 1559 1775 1560 1779
rect 1564 1778 1565 1779
rect 1590 1779 1596 1780
rect 1590 1778 1591 1779
rect 1564 1776 1591 1778
rect 1564 1775 1565 1776
rect 1559 1774 1565 1775
rect 1590 1775 1591 1776
rect 1595 1775 1596 1779
rect 1590 1774 1596 1775
rect 1606 1779 1612 1780
rect 1606 1775 1607 1779
rect 1611 1778 1612 1779
rect 1623 1779 1629 1780
rect 1623 1778 1624 1779
rect 1611 1776 1624 1778
rect 1611 1775 1612 1776
rect 1606 1774 1612 1775
rect 1623 1775 1624 1776
rect 1628 1775 1629 1779
rect 1623 1774 1629 1775
rect 1687 1779 1693 1780
rect 1687 1775 1688 1779
rect 1692 1778 1693 1779
rect 1718 1779 1724 1780
rect 1718 1778 1719 1779
rect 1692 1776 1719 1778
rect 1692 1775 1693 1776
rect 1687 1774 1693 1775
rect 1718 1775 1719 1776
rect 1723 1775 1724 1779
rect 1718 1774 1724 1775
rect 1751 1779 1757 1780
rect 1751 1775 1752 1779
rect 1756 1778 1757 1779
rect 1774 1779 1780 1780
rect 1774 1778 1775 1779
rect 1756 1776 1775 1778
rect 1756 1775 1757 1776
rect 1751 1774 1757 1775
rect 1774 1775 1775 1776
rect 1779 1775 1780 1779
rect 1774 1774 1780 1775
rect 1807 1779 1813 1780
rect 1807 1775 1808 1779
rect 1812 1778 1813 1779
rect 1830 1779 1836 1780
rect 1830 1778 1831 1779
rect 1812 1776 1831 1778
rect 1812 1775 1813 1776
rect 1807 1774 1813 1775
rect 1830 1775 1831 1776
rect 1835 1775 1836 1779
rect 1830 1774 1836 1775
rect 1863 1779 1869 1780
rect 1863 1775 1864 1779
rect 1868 1778 1869 1779
rect 1886 1779 1892 1780
rect 1886 1778 1887 1779
rect 1868 1776 1887 1778
rect 1868 1775 1869 1776
rect 1863 1774 1869 1775
rect 1886 1775 1887 1776
rect 1891 1775 1892 1779
rect 1886 1774 1892 1775
rect 1919 1779 1925 1780
rect 1919 1775 1920 1779
rect 1924 1778 1925 1779
rect 1950 1779 1956 1780
rect 1950 1778 1951 1779
rect 1924 1776 1951 1778
rect 1924 1775 1925 1776
rect 1919 1774 1925 1775
rect 1950 1775 1951 1776
rect 1955 1775 1956 1779
rect 1983 1779 1989 1780
rect 1983 1778 1984 1779
rect 1950 1774 1956 1775
rect 1960 1776 1984 1778
rect 1278 1771 1284 1772
rect 1742 1771 1748 1772
rect 1187 1770 1193 1771
rect 134 1767 140 1768
rect 134 1763 135 1767
rect 139 1763 140 1767
rect 134 1762 140 1763
rect 174 1767 180 1768
rect 174 1763 175 1767
rect 179 1763 180 1767
rect 174 1762 180 1763
rect 214 1767 220 1768
rect 214 1763 215 1767
rect 219 1763 220 1767
rect 214 1762 220 1763
rect 286 1767 292 1768
rect 286 1763 287 1767
rect 291 1763 292 1767
rect 286 1762 292 1763
rect 374 1767 380 1768
rect 374 1763 375 1767
rect 379 1763 380 1767
rect 374 1762 380 1763
rect 470 1767 476 1768
rect 470 1763 471 1767
rect 475 1763 476 1767
rect 470 1762 476 1763
rect 566 1767 572 1768
rect 566 1763 567 1767
rect 571 1763 572 1767
rect 566 1762 572 1763
rect 662 1767 668 1768
rect 662 1763 663 1767
rect 667 1763 668 1767
rect 662 1762 668 1763
rect 750 1767 756 1768
rect 750 1763 751 1767
rect 755 1763 756 1767
rect 750 1762 756 1763
rect 830 1767 836 1768
rect 830 1763 831 1767
rect 835 1763 836 1767
rect 830 1762 836 1763
rect 902 1767 908 1768
rect 902 1763 903 1767
rect 907 1763 908 1767
rect 902 1762 908 1763
rect 966 1767 972 1768
rect 966 1763 967 1767
rect 971 1763 972 1767
rect 966 1762 972 1763
rect 1030 1767 1036 1768
rect 1030 1763 1031 1767
rect 1035 1763 1036 1767
rect 1030 1762 1036 1763
rect 1086 1767 1092 1768
rect 1086 1763 1087 1767
rect 1091 1763 1092 1767
rect 1086 1762 1092 1763
rect 1150 1767 1156 1768
rect 1150 1763 1151 1767
rect 1155 1763 1156 1767
rect 1150 1762 1156 1763
rect 1190 1767 1196 1768
rect 1190 1763 1191 1767
rect 1195 1763 1196 1767
rect 1742 1767 1743 1771
rect 1747 1770 1748 1771
rect 1960 1770 1962 1776
rect 1983 1775 1984 1776
rect 1988 1775 1989 1779
rect 1983 1774 1989 1775
rect 2406 1776 2412 1777
rect 2406 1772 2407 1776
rect 2411 1772 2412 1776
rect 2406 1771 2412 1772
rect 1747 1768 1962 1770
rect 1747 1767 1748 1768
rect 1742 1766 1748 1767
rect 1190 1762 1196 1763
rect 1406 1753 1412 1754
rect 1406 1749 1407 1753
rect 1411 1749 1412 1753
rect 1406 1748 1412 1749
rect 1470 1753 1476 1754
rect 1470 1749 1471 1753
rect 1475 1749 1476 1753
rect 1470 1748 1476 1749
rect 1534 1753 1540 1754
rect 1534 1749 1535 1753
rect 1539 1749 1540 1753
rect 1534 1748 1540 1749
rect 1598 1753 1604 1754
rect 1598 1749 1599 1753
rect 1603 1749 1604 1753
rect 1598 1748 1604 1749
rect 1662 1753 1668 1754
rect 1662 1749 1663 1753
rect 1667 1749 1668 1753
rect 1662 1748 1668 1749
rect 1726 1753 1732 1754
rect 1726 1749 1727 1753
rect 1731 1749 1732 1753
rect 1726 1748 1732 1749
rect 1782 1753 1788 1754
rect 1782 1749 1783 1753
rect 1787 1749 1788 1753
rect 1782 1748 1788 1749
rect 1838 1753 1844 1754
rect 1838 1749 1839 1753
rect 1843 1749 1844 1753
rect 1838 1748 1844 1749
rect 1894 1753 1900 1754
rect 1894 1749 1895 1753
rect 1899 1749 1900 1753
rect 1894 1748 1900 1749
rect 1958 1753 1964 1754
rect 1958 1749 1959 1753
rect 1963 1749 1964 1753
rect 1958 1748 1964 1749
rect 682 1747 688 1748
rect 110 1744 116 1745
rect 110 1740 111 1744
rect 115 1740 116 1744
rect 682 1743 683 1747
rect 687 1746 688 1747
rect 687 1744 790 1746
rect 687 1743 688 1744
rect 682 1742 688 1743
rect 110 1739 116 1740
rect 158 1739 165 1740
rect 158 1735 159 1739
rect 164 1735 165 1739
rect 158 1734 165 1735
rect 198 1739 205 1740
rect 198 1735 199 1739
rect 204 1735 205 1739
rect 198 1734 205 1735
rect 239 1739 248 1740
rect 239 1735 240 1739
rect 247 1735 248 1739
rect 239 1734 248 1735
rect 311 1739 320 1740
rect 311 1735 312 1739
rect 319 1735 320 1739
rect 311 1734 320 1735
rect 399 1739 408 1740
rect 399 1735 400 1739
rect 407 1735 408 1739
rect 399 1734 408 1735
rect 495 1739 504 1740
rect 495 1735 496 1739
rect 503 1735 504 1739
rect 591 1739 597 1740
rect 591 1738 592 1739
rect 495 1734 504 1735
rect 508 1736 592 1738
rect 142 1731 148 1732
rect 110 1727 116 1728
rect 110 1723 111 1727
rect 115 1723 116 1727
rect 142 1727 143 1731
rect 147 1730 148 1731
rect 508 1730 510 1736
rect 591 1735 592 1736
rect 596 1735 597 1739
rect 591 1734 597 1735
rect 687 1739 696 1740
rect 687 1735 688 1739
rect 695 1735 696 1739
rect 687 1734 696 1735
rect 775 1739 784 1740
rect 775 1735 776 1739
rect 783 1735 784 1739
rect 788 1738 790 1744
rect 1238 1744 1244 1745
rect 1238 1740 1239 1744
rect 1243 1740 1244 1744
rect 855 1739 861 1740
rect 855 1738 856 1739
rect 788 1736 856 1738
rect 775 1734 784 1735
rect 855 1735 856 1736
rect 860 1735 861 1739
rect 855 1734 861 1735
rect 890 1739 896 1740
rect 890 1735 891 1739
rect 895 1738 896 1739
rect 927 1739 933 1740
rect 927 1738 928 1739
rect 895 1736 928 1738
rect 895 1735 896 1736
rect 890 1734 896 1735
rect 927 1735 928 1736
rect 932 1735 933 1739
rect 927 1734 933 1735
rect 954 1739 960 1740
rect 954 1735 955 1739
rect 959 1738 960 1739
rect 991 1739 997 1740
rect 991 1738 992 1739
rect 959 1736 992 1738
rect 959 1735 960 1736
rect 954 1734 960 1735
rect 991 1735 992 1736
rect 996 1735 997 1739
rect 991 1734 997 1735
rect 1055 1739 1061 1740
rect 1055 1735 1056 1739
rect 1060 1738 1061 1739
rect 1063 1739 1069 1740
rect 1063 1738 1064 1739
rect 1060 1736 1064 1738
rect 1060 1735 1061 1736
rect 1055 1734 1061 1735
rect 1063 1735 1064 1736
rect 1068 1735 1069 1739
rect 1063 1734 1069 1735
rect 1111 1739 1120 1740
rect 1111 1735 1112 1739
rect 1119 1735 1120 1739
rect 1111 1734 1120 1735
rect 1174 1739 1181 1740
rect 1174 1735 1175 1739
rect 1180 1735 1181 1739
rect 1174 1734 1181 1735
rect 1215 1739 1221 1740
rect 1238 1739 1244 1740
rect 1403 1743 1409 1744
rect 1403 1739 1404 1743
rect 1408 1742 1409 1743
rect 1446 1743 1452 1744
rect 1446 1742 1447 1743
rect 1408 1740 1447 1742
rect 1408 1739 1409 1740
rect 1215 1735 1216 1739
rect 1220 1738 1221 1739
rect 1403 1738 1409 1739
rect 1446 1739 1447 1740
rect 1451 1739 1452 1743
rect 1446 1738 1452 1739
rect 1462 1743 1473 1744
rect 1462 1739 1463 1743
rect 1467 1739 1468 1743
rect 1472 1739 1473 1743
rect 1462 1738 1473 1739
rect 1526 1743 1537 1744
rect 1526 1739 1527 1743
rect 1531 1739 1532 1743
rect 1536 1739 1537 1743
rect 1526 1738 1537 1739
rect 1590 1743 1601 1744
rect 1590 1739 1591 1743
rect 1595 1739 1596 1743
rect 1600 1739 1601 1743
rect 1590 1738 1601 1739
rect 1659 1743 1665 1744
rect 1659 1739 1660 1743
rect 1664 1742 1665 1743
rect 1670 1743 1676 1744
rect 1670 1742 1671 1743
rect 1664 1740 1671 1742
rect 1664 1739 1665 1740
rect 1659 1738 1665 1739
rect 1670 1739 1671 1740
rect 1675 1739 1676 1743
rect 1670 1738 1676 1739
rect 1718 1743 1729 1744
rect 1718 1739 1719 1743
rect 1723 1739 1724 1743
rect 1728 1739 1729 1743
rect 1718 1738 1729 1739
rect 1774 1743 1785 1744
rect 1774 1739 1775 1743
rect 1779 1739 1780 1743
rect 1784 1739 1785 1743
rect 1774 1738 1785 1739
rect 1830 1743 1841 1744
rect 1830 1739 1831 1743
rect 1835 1739 1836 1743
rect 1840 1739 1841 1743
rect 1830 1738 1841 1739
rect 1886 1743 1897 1744
rect 1886 1739 1887 1743
rect 1891 1739 1892 1743
rect 1896 1739 1897 1743
rect 1886 1738 1897 1739
rect 1950 1743 1961 1744
rect 1950 1739 1951 1743
rect 1955 1739 1956 1743
rect 1960 1739 1961 1743
rect 1950 1738 1961 1739
rect 1220 1736 1234 1738
rect 1220 1735 1221 1736
rect 1215 1734 1221 1735
rect 1232 1734 1234 1736
rect 1232 1733 1305 1734
rect 1232 1732 1300 1733
rect 147 1728 510 1730
rect 1299 1729 1300 1732
rect 1304 1729 1305 1733
rect 1299 1728 1305 1729
rect 1330 1731 1336 1732
rect 147 1727 148 1728
rect 142 1726 148 1727
rect 1238 1727 1244 1728
rect 110 1722 116 1723
rect 1238 1723 1239 1727
rect 1243 1723 1244 1727
rect 1330 1727 1331 1731
rect 1335 1730 1336 1731
rect 1347 1731 1353 1732
rect 1347 1730 1348 1731
rect 1335 1728 1348 1730
rect 1335 1727 1336 1728
rect 1330 1726 1336 1727
rect 1347 1727 1348 1728
rect 1352 1727 1353 1731
rect 1347 1726 1353 1727
rect 1419 1731 1425 1732
rect 1419 1727 1420 1731
rect 1424 1730 1425 1731
rect 1486 1731 1492 1732
rect 1486 1730 1487 1731
rect 1424 1728 1487 1730
rect 1424 1727 1425 1728
rect 1419 1726 1425 1727
rect 1486 1727 1487 1728
rect 1491 1727 1492 1731
rect 1486 1726 1492 1727
rect 1499 1731 1505 1732
rect 1499 1727 1500 1731
rect 1504 1730 1505 1731
rect 1570 1731 1576 1732
rect 1570 1730 1571 1731
rect 1504 1728 1571 1730
rect 1504 1727 1505 1728
rect 1499 1726 1505 1727
rect 1570 1727 1571 1728
rect 1575 1727 1576 1731
rect 1570 1726 1576 1727
rect 1579 1731 1585 1732
rect 1579 1727 1580 1731
rect 1584 1730 1585 1731
rect 1650 1731 1656 1732
rect 1650 1730 1651 1731
rect 1584 1728 1651 1730
rect 1584 1727 1585 1728
rect 1579 1726 1585 1727
rect 1650 1727 1651 1728
rect 1655 1727 1656 1731
rect 1650 1726 1656 1727
rect 1659 1731 1665 1732
rect 1659 1727 1660 1731
rect 1664 1730 1665 1731
rect 1703 1731 1709 1732
rect 1703 1730 1704 1731
rect 1664 1728 1704 1730
rect 1664 1727 1665 1728
rect 1659 1726 1665 1727
rect 1703 1727 1704 1728
rect 1708 1727 1709 1731
rect 1703 1726 1709 1727
rect 1731 1731 1737 1732
rect 1731 1727 1732 1731
rect 1736 1730 1737 1731
rect 1742 1731 1748 1732
rect 1742 1730 1743 1731
rect 1736 1728 1743 1730
rect 1736 1727 1737 1728
rect 1731 1726 1737 1727
rect 1742 1727 1743 1728
rect 1747 1727 1748 1731
rect 1742 1726 1748 1727
rect 1762 1731 1768 1732
rect 1762 1727 1763 1731
rect 1767 1730 1768 1731
rect 1803 1731 1809 1732
rect 1803 1730 1804 1731
rect 1767 1728 1804 1730
rect 1767 1727 1768 1728
rect 1762 1726 1768 1727
rect 1803 1727 1804 1728
rect 1808 1727 1809 1731
rect 1803 1726 1809 1727
rect 1839 1731 1845 1732
rect 1839 1727 1840 1731
rect 1844 1730 1845 1731
rect 1867 1731 1873 1732
rect 1867 1730 1868 1731
rect 1844 1728 1868 1730
rect 1844 1727 1845 1728
rect 1839 1726 1845 1727
rect 1867 1727 1868 1728
rect 1872 1727 1873 1731
rect 1867 1726 1873 1727
rect 1918 1731 1924 1732
rect 1918 1727 1919 1731
rect 1923 1730 1924 1731
rect 1931 1731 1937 1732
rect 1931 1730 1932 1731
rect 1923 1728 1932 1730
rect 1923 1727 1924 1728
rect 1918 1726 1924 1727
rect 1931 1727 1932 1728
rect 1936 1727 1937 1731
rect 1931 1726 1937 1727
rect 1966 1731 1972 1732
rect 1966 1727 1967 1731
rect 1971 1730 1972 1731
rect 1995 1731 2001 1732
rect 1995 1730 1996 1731
rect 1971 1728 1996 1730
rect 1971 1727 1972 1728
rect 1966 1726 1972 1727
rect 1995 1727 1996 1728
rect 2000 1727 2001 1731
rect 1995 1726 2001 1727
rect 2026 1731 2032 1732
rect 2026 1727 2027 1731
rect 2031 1730 2032 1731
rect 2059 1731 2065 1732
rect 2059 1730 2060 1731
rect 2031 1728 2060 1730
rect 2031 1727 2032 1728
rect 2026 1726 2032 1727
rect 2059 1727 2060 1728
rect 2064 1727 2065 1731
rect 2059 1726 2065 1727
rect 1238 1722 1244 1723
rect 1302 1723 1308 1724
rect 134 1720 140 1721
rect 134 1716 135 1720
rect 139 1716 140 1720
rect 134 1715 140 1716
rect 174 1720 180 1721
rect 174 1716 175 1720
rect 179 1716 180 1720
rect 174 1715 180 1716
rect 214 1720 220 1721
rect 214 1716 215 1720
rect 219 1716 220 1720
rect 214 1715 220 1716
rect 286 1720 292 1721
rect 286 1716 287 1720
rect 291 1716 292 1720
rect 286 1715 292 1716
rect 374 1720 380 1721
rect 374 1716 375 1720
rect 379 1716 380 1720
rect 374 1715 380 1716
rect 470 1720 476 1721
rect 470 1716 471 1720
rect 475 1716 476 1720
rect 470 1715 476 1716
rect 566 1720 572 1721
rect 566 1716 567 1720
rect 571 1716 572 1720
rect 566 1715 572 1716
rect 662 1720 668 1721
rect 662 1716 663 1720
rect 667 1716 668 1720
rect 662 1715 668 1716
rect 750 1720 756 1721
rect 750 1716 751 1720
rect 755 1716 756 1720
rect 750 1715 756 1716
rect 830 1720 836 1721
rect 830 1716 831 1720
rect 835 1716 836 1720
rect 830 1715 836 1716
rect 902 1720 908 1721
rect 902 1716 903 1720
rect 907 1716 908 1720
rect 902 1715 908 1716
rect 966 1720 972 1721
rect 966 1716 967 1720
rect 971 1716 972 1720
rect 966 1715 972 1716
rect 1030 1720 1036 1721
rect 1030 1716 1031 1720
rect 1035 1716 1036 1720
rect 1030 1715 1036 1716
rect 1086 1720 1092 1721
rect 1086 1716 1087 1720
rect 1091 1716 1092 1720
rect 1086 1715 1092 1716
rect 1150 1720 1156 1721
rect 1150 1716 1151 1720
rect 1155 1716 1156 1720
rect 1150 1715 1156 1716
rect 1190 1720 1196 1721
rect 1190 1716 1191 1720
rect 1195 1716 1196 1720
rect 1302 1719 1303 1723
rect 1307 1719 1308 1723
rect 1302 1718 1308 1719
rect 1350 1723 1356 1724
rect 1350 1719 1351 1723
rect 1355 1719 1356 1723
rect 1350 1718 1356 1719
rect 1422 1723 1428 1724
rect 1422 1719 1423 1723
rect 1427 1719 1428 1723
rect 1422 1718 1428 1719
rect 1502 1723 1508 1724
rect 1502 1719 1503 1723
rect 1507 1719 1508 1723
rect 1502 1718 1508 1719
rect 1582 1723 1588 1724
rect 1582 1719 1583 1723
rect 1587 1719 1588 1723
rect 1582 1718 1588 1719
rect 1662 1723 1668 1724
rect 1662 1719 1663 1723
rect 1667 1719 1668 1723
rect 1662 1718 1668 1719
rect 1734 1723 1740 1724
rect 1734 1719 1735 1723
rect 1739 1719 1740 1723
rect 1734 1718 1740 1719
rect 1806 1723 1812 1724
rect 1806 1719 1807 1723
rect 1811 1719 1812 1723
rect 1806 1718 1812 1719
rect 1870 1723 1876 1724
rect 1870 1719 1871 1723
rect 1875 1719 1876 1723
rect 1870 1718 1876 1719
rect 1934 1723 1940 1724
rect 1934 1719 1935 1723
rect 1939 1719 1940 1723
rect 1934 1718 1940 1719
rect 1998 1723 2004 1724
rect 1998 1719 1999 1723
rect 2003 1719 2004 1723
rect 1998 1718 2004 1719
rect 2062 1723 2068 1724
rect 2062 1719 2063 1723
rect 2067 1719 2068 1723
rect 2062 1718 2068 1719
rect 1190 1715 1196 1716
rect 134 1704 140 1705
rect 134 1700 135 1704
rect 139 1700 140 1704
rect 134 1699 140 1700
rect 174 1704 180 1705
rect 174 1700 175 1704
rect 179 1700 180 1704
rect 174 1699 180 1700
rect 238 1704 244 1705
rect 238 1700 239 1704
rect 243 1700 244 1704
rect 238 1699 244 1700
rect 318 1704 324 1705
rect 318 1700 319 1704
rect 323 1700 324 1704
rect 318 1699 324 1700
rect 414 1704 420 1705
rect 414 1700 415 1704
rect 419 1700 420 1704
rect 414 1699 420 1700
rect 510 1704 516 1705
rect 510 1700 511 1704
rect 515 1700 516 1704
rect 510 1699 516 1700
rect 614 1704 620 1705
rect 614 1700 615 1704
rect 619 1700 620 1704
rect 614 1699 620 1700
rect 710 1704 716 1705
rect 710 1700 711 1704
rect 715 1700 716 1704
rect 710 1699 716 1700
rect 798 1704 804 1705
rect 798 1700 799 1704
rect 803 1700 804 1704
rect 798 1699 804 1700
rect 878 1704 884 1705
rect 878 1700 879 1704
rect 883 1700 884 1704
rect 878 1699 884 1700
rect 950 1704 956 1705
rect 950 1700 951 1704
rect 955 1700 956 1704
rect 950 1699 956 1700
rect 1014 1704 1020 1705
rect 1014 1700 1015 1704
rect 1019 1700 1020 1704
rect 1014 1699 1020 1700
rect 1086 1704 1092 1705
rect 1086 1700 1087 1704
rect 1091 1700 1092 1704
rect 1086 1699 1092 1700
rect 1158 1704 1164 1705
rect 1158 1700 1159 1704
rect 1163 1700 1164 1704
rect 1158 1699 1164 1700
rect 1278 1700 1284 1701
rect 2406 1700 2412 1701
rect 110 1697 116 1698
rect 110 1693 111 1697
rect 115 1693 116 1697
rect 110 1692 116 1693
rect 1238 1697 1244 1698
rect 1238 1693 1239 1697
rect 1243 1693 1244 1697
rect 1278 1696 1279 1700
rect 1283 1696 1284 1700
rect 1918 1699 1924 1700
rect 1918 1698 1919 1699
rect 1895 1697 1919 1698
rect 1278 1695 1284 1696
rect 1327 1695 1336 1696
rect 1238 1692 1244 1693
rect 1006 1691 1012 1692
rect 1006 1687 1007 1691
rect 1011 1690 1012 1691
rect 1327 1691 1328 1695
rect 1335 1691 1336 1695
rect 1327 1690 1336 1691
rect 1338 1695 1344 1696
rect 1338 1691 1339 1695
rect 1343 1694 1344 1695
rect 1375 1695 1381 1696
rect 1375 1694 1376 1695
rect 1343 1692 1376 1694
rect 1343 1691 1344 1692
rect 1338 1690 1344 1691
rect 1375 1691 1376 1692
rect 1380 1691 1381 1695
rect 1375 1690 1381 1691
rect 1446 1695 1453 1696
rect 1446 1691 1447 1695
rect 1452 1691 1453 1695
rect 1446 1690 1453 1691
rect 1486 1695 1492 1696
rect 1486 1691 1487 1695
rect 1491 1694 1492 1695
rect 1527 1695 1533 1696
rect 1527 1694 1528 1695
rect 1491 1692 1528 1694
rect 1491 1691 1492 1692
rect 1486 1690 1492 1691
rect 1527 1691 1528 1692
rect 1532 1691 1533 1695
rect 1527 1690 1533 1691
rect 1570 1695 1576 1696
rect 1570 1691 1571 1695
rect 1575 1694 1576 1695
rect 1607 1695 1613 1696
rect 1607 1694 1608 1695
rect 1575 1692 1608 1694
rect 1575 1691 1576 1692
rect 1570 1690 1576 1691
rect 1607 1691 1608 1692
rect 1612 1691 1613 1695
rect 1607 1690 1613 1691
rect 1650 1695 1656 1696
rect 1650 1691 1651 1695
rect 1655 1694 1656 1695
rect 1687 1695 1693 1696
rect 1687 1694 1688 1695
rect 1655 1692 1688 1694
rect 1655 1691 1656 1692
rect 1650 1690 1656 1691
rect 1687 1691 1688 1692
rect 1692 1691 1693 1695
rect 1687 1690 1693 1691
rect 1759 1695 1768 1696
rect 1759 1691 1760 1695
rect 1767 1691 1768 1695
rect 1759 1690 1768 1691
rect 1831 1695 1837 1696
rect 1831 1691 1832 1695
rect 1836 1694 1837 1695
rect 1839 1695 1845 1696
rect 1839 1694 1840 1695
rect 1836 1692 1840 1694
rect 1836 1691 1837 1692
rect 1831 1690 1837 1691
rect 1839 1691 1840 1692
rect 1844 1691 1845 1695
rect 1895 1693 1896 1697
rect 1900 1696 1919 1697
rect 1900 1693 1901 1696
rect 1918 1695 1919 1696
rect 1923 1695 1924 1699
rect 2406 1696 2407 1700
rect 2411 1696 2412 1700
rect 1918 1694 1924 1695
rect 1959 1695 1968 1696
rect 1895 1692 1901 1693
rect 1839 1690 1845 1691
rect 1959 1691 1960 1695
rect 1967 1691 1968 1695
rect 1959 1690 1968 1691
rect 2023 1695 2032 1696
rect 2023 1691 2024 1695
rect 2031 1691 2032 1695
rect 2023 1690 2032 1691
rect 2087 1695 2093 1696
rect 2406 1695 2412 1696
rect 2087 1691 2088 1695
rect 2092 1691 2093 1695
rect 2087 1690 2093 1691
rect 1011 1688 1161 1690
rect 1011 1687 1012 1688
rect 1006 1686 1012 1687
rect 159 1683 168 1684
rect 110 1680 116 1681
rect 110 1676 111 1680
rect 115 1676 116 1680
rect 159 1679 160 1683
rect 167 1679 168 1683
rect 159 1678 168 1679
rect 199 1683 205 1684
rect 199 1679 200 1683
rect 204 1682 205 1683
rect 230 1683 236 1684
rect 230 1682 231 1683
rect 204 1680 231 1682
rect 204 1679 205 1680
rect 199 1678 205 1679
rect 230 1679 231 1680
rect 235 1679 236 1683
rect 230 1678 236 1679
rect 263 1683 269 1684
rect 263 1679 264 1683
rect 268 1682 269 1683
rect 310 1683 316 1684
rect 310 1682 311 1683
rect 268 1680 311 1682
rect 268 1679 269 1680
rect 263 1678 269 1679
rect 310 1679 311 1680
rect 315 1679 316 1683
rect 310 1678 316 1679
rect 343 1683 349 1684
rect 343 1679 344 1683
rect 348 1682 349 1683
rect 406 1683 412 1684
rect 406 1682 407 1683
rect 348 1680 407 1682
rect 348 1679 349 1680
rect 343 1678 349 1679
rect 406 1679 407 1680
rect 411 1679 412 1683
rect 406 1678 412 1679
rect 439 1683 445 1684
rect 439 1679 440 1683
rect 444 1682 445 1683
rect 502 1683 508 1684
rect 502 1682 503 1683
rect 444 1680 503 1682
rect 444 1679 445 1680
rect 439 1678 445 1679
rect 502 1679 503 1680
rect 507 1679 508 1683
rect 502 1678 508 1679
rect 535 1683 541 1684
rect 535 1679 536 1683
rect 540 1682 541 1683
rect 606 1683 612 1684
rect 606 1682 607 1683
rect 540 1680 607 1682
rect 540 1679 541 1680
rect 535 1678 541 1679
rect 606 1679 607 1680
rect 611 1679 612 1683
rect 606 1678 612 1679
rect 622 1683 628 1684
rect 622 1679 623 1683
rect 627 1682 628 1683
rect 639 1683 645 1684
rect 639 1682 640 1683
rect 627 1680 640 1682
rect 627 1679 628 1680
rect 622 1678 628 1679
rect 639 1679 640 1680
rect 644 1679 645 1683
rect 639 1678 645 1679
rect 735 1683 741 1684
rect 735 1679 736 1683
rect 740 1682 741 1683
rect 790 1683 796 1684
rect 790 1682 791 1683
rect 740 1680 791 1682
rect 740 1679 741 1680
rect 735 1678 741 1679
rect 790 1679 791 1680
rect 795 1679 796 1683
rect 790 1678 796 1679
rect 823 1683 829 1684
rect 823 1679 824 1683
rect 828 1682 829 1683
rect 870 1683 876 1684
rect 870 1682 871 1683
rect 828 1680 871 1682
rect 828 1679 829 1680
rect 823 1678 829 1679
rect 870 1679 871 1680
rect 875 1679 876 1683
rect 870 1678 876 1679
rect 903 1683 909 1684
rect 903 1679 904 1683
rect 908 1682 909 1683
rect 942 1683 948 1684
rect 942 1682 943 1683
rect 908 1680 943 1682
rect 908 1679 909 1680
rect 903 1678 909 1679
rect 942 1679 943 1680
rect 947 1679 948 1683
rect 942 1678 948 1679
rect 975 1683 981 1684
rect 975 1679 976 1683
rect 980 1682 981 1683
rect 1006 1683 1012 1684
rect 1006 1682 1007 1683
rect 980 1680 1007 1682
rect 980 1679 981 1680
rect 975 1678 981 1679
rect 1006 1679 1007 1680
rect 1011 1679 1012 1683
rect 1006 1678 1012 1679
rect 1039 1683 1045 1684
rect 1039 1679 1040 1683
rect 1044 1682 1045 1683
rect 1078 1683 1084 1684
rect 1078 1682 1079 1683
rect 1044 1680 1079 1682
rect 1044 1679 1045 1680
rect 1039 1678 1045 1679
rect 1078 1679 1079 1680
rect 1083 1679 1084 1683
rect 1078 1678 1084 1679
rect 1111 1683 1117 1684
rect 1111 1679 1112 1683
rect 1116 1682 1117 1683
rect 1150 1683 1156 1684
rect 1150 1682 1151 1683
rect 1116 1680 1151 1682
rect 1116 1679 1117 1680
rect 1111 1678 1117 1679
rect 1150 1679 1151 1680
rect 1155 1679 1156 1683
rect 1159 1682 1161 1688
rect 1822 1687 1828 1688
rect 1183 1683 1189 1684
rect 1183 1682 1184 1683
rect 1159 1680 1184 1682
rect 1150 1678 1156 1679
rect 1183 1679 1184 1680
rect 1188 1679 1189 1683
rect 1278 1683 1284 1684
rect 1183 1678 1189 1679
rect 1238 1680 1244 1681
rect 110 1675 116 1676
rect 1238 1676 1239 1680
rect 1243 1676 1244 1680
rect 1278 1679 1279 1683
rect 1283 1679 1284 1683
rect 1822 1683 1823 1687
rect 1827 1686 1828 1687
rect 2089 1686 2091 1690
rect 1827 1684 2091 1686
rect 1827 1683 1828 1684
rect 1822 1682 1828 1683
rect 2406 1683 2412 1684
rect 1278 1678 1284 1679
rect 2406 1679 2407 1683
rect 2411 1679 2412 1683
rect 2406 1678 2412 1679
rect 1238 1675 1244 1676
rect 1302 1676 1308 1677
rect 1302 1672 1303 1676
rect 1307 1672 1308 1676
rect 1302 1671 1308 1672
rect 1350 1676 1356 1677
rect 1350 1672 1351 1676
rect 1355 1672 1356 1676
rect 1350 1671 1356 1672
rect 1422 1676 1428 1677
rect 1422 1672 1423 1676
rect 1427 1672 1428 1676
rect 1422 1671 1428 1672
rect 1502 1676 1508 1677
rect 1502 1672 1503 1676
rect 1507 1672 1508 1676
rect 1502 1671 1508 1672
rect 1582 1676 1588 1677
rect 1582 1672 1583 1676
rect 1587 1672 1588 1676
rect 1582 1671 1588 1672
rect 1662 1676 1668 1677
rect 1662 1672 1663 1676
rect 1667 1672 1668 1676
rect 1662 1671 1668 1672
rect 1734 1676 1740 1677
rect 1734 1672 1735 1676
rect 1739 1672 1740 1676
rect 1734 1671 1740 1672
rect 1806 1676 1812 1677
rect 1806 1672 1807 1676
rect 1811 1672 1812 1676
rect 1806 1671 1812 1672
rect 1870 1676 1876 1677
rect 1870 1672 1871 1676
rect 1875 1672 1876 1676
rect 1870 1671 1876 1672
rect 1934 1676 1940 1677
rect 1934 1672 1935 1676
rect 1939 1672 1940 1676
rect 1934 1671 1940 1672
rect 1998 1676 2004 1677
rect 1998 1672 1999 1676
rect 2003 1672 2004 1676
rect 1998 1671 2004 1672
rect 2062 1676 2068 1677
rect 2062 1672 2063 1676
rect 2067 1672 2068 1676
rect 2062 1671 2068 1672
rect 1302 1664 1308 1665
rect 1302 1660 1303 1664
rect 1307 1660 1308 1664
rect 1302 1659 1308 1660
rect 1358 1664 1364 1665
rect 1358 1660 1359 1664
rect 1363 1660 1364 1664
rect 1358 1659 1364 1660
rect 1446 1664 1452 1665
rect 1446 1660 1447 1664
rect 1451 1660 1452 1664
rect 1446 1659 1452 1660
rect 1542 1664 1548 1665
rect 1542 1660 1543 1664
rect 1547 1660 1548 1664
rect 1542 1659 1548 1660
rect 1638 1664 1644 1665
rect 1638 1660 1639 1664
rect 1643 1660 1644 1664
rect 1638 1659 1644 1660
rect 1726 1664 1732 1665
rect 1726 1660 1727 1664
rect 1731 1660 1732 1664
rect 1726 1659 1732 1660
rect 1814 1664 1820 1665
rect 1814 1660 1815 1664
rect 1819 1660 1820 1664
rect 1814 1659 1820 1660
rect 1894 1664 1900 1665
rect 1894 1660 1895 1664
rect 1899 1660 1900 1664
rect 1894 1659 1900 1660
rect 1966 1664 1972 1665
rect 1966 1660 1967 1664
rect 1971 1660 1972 1664
rect 1966 1659 1972 1660
rect 2030 1664 2036 1665
rect 2030 1660 2031 1664
rect 2035 1660 2036 1664
rect 2030 1659 2036 1660
rect 2094 1664 2100 1665
rect 2094 1660 2095 1664
rect 2099 1660 2100 1664
rect 2094 1659 2100 1660
rect 2158 1664 2164 1665
rect 2158 1660 2159 1664
rect 2163 1660 2164 1664
rect 2158 1659 2164 1660
rect 2222 1664 2228 1665
rect 2222 1660 2223 1664
rect 2227 1660 2228 1664
rect 2222 1659 2228 1660
rect 134 1657 140 1658
rect 134 1653 135 1657
rect 139 1653 140 1657
rect 134 1652 140 1653
rect 174 1657 180 1658
rect 174 1653 175 1657
rect 179 1653 180 1657
rect 174 1652 180 1653
rect 238 1657 244 1658
rect 238 1653 239 1657
rect 243 1653 244 1657
rect 238 1652 244 1653
rect 318 1657 324 1658
rect 318 1653 319 1657
rect 323 1653 324 1657
rect 318 1652 324 1653
rect 414 1657 420 1658
rect 414 1653 415 1657
rect 419 1653 420 1657
rect 414 1652 420 1653
rect 510 1657 516 1658
rect 510 1653 511 1657
rect 515 1653 516 1657
rect 510 1652 516 1653
rect 614 1657 620 1658
rect 614 1653 615 1657
rect 619 1653 620 1657
rect 614 1652 620 1653
rect 710 1657 716 1658
rect 710 1653 711 1657
rect 715 1653 716 1657
rect 710 1652 716 1653
rect 798 1657 804 1658
rect 798 1653 799 1657
rect 803 1653 804 1657
rect 798 1652 804 1653
rect 878 1657 884 1658
rect 878 1653 879 1657
rect 883 1653 884 1657
rect 878 1652 884 1653
rect 950 1657 956 1658
rect 950 1653 951 1657
rect 955 1653 956 1657
rect 950 1652 956 1653
rect 1014 1657 1020 1658
rect 1014 1653 1015 1657
rect 1019 1653 1020 1657
rect 1014 1652 1020 1653
rect 1086 1657 1092 1658
rect 1086 1653 1087 1657
rect 1091 1653 1092 1657
rect 1086 1652 1092 1653
rect 1158 1657 1164 1658
rect 1158 1653 1159 1657
rect 1163 1653 1164 1657
rect 1158 1652 1164 1653
rect 1278 1657 1284 1658
rect 1278 1653 1279 1657
rect 1283 1653 1284 1657
rect 1278 1652 1284 1653
rect 2406 1657 2412 1658
rect 2406 1653 2407 1657
rect 2411 1653 2412 1657
rect 2406 1652 2412 1653
rect 1703 1651 1709 1652
rect 131 1647 137 1648
rect 131 1643 132 1647
rect 136 1646 137 1647
rect 142 1647 148 1648
rect 142 1646 143 1647
rect 136 1644 143 1646
rect 136 1643 137 1644
rect 131 1642 137 1643
rect 142 1643 143 1644
rect 147 1643 148 1647
rect 142 1642 148 1643
rect 162 1647 168 1648
rect 162 1643 163 1647
rect 167 1646 168 1647
rect 171 1647 177 1648
rect 171 1646 172 1647
rect 167 1644 172 1646
rect 167 1643 168 1644
rect 162 1642 168 1643
rect 171 1643 172 1644
rect 176 1643 177 1647
rect 171 1642 177 1643
rect 230 1647 241 1648
rect 230 1643 231 1647
rect 235 1643 236 1647
rect 240 1643 241 1647
rect 230 1642 241 1643
rect 310 1647 321 1648
rect 310 1643 311 1647
rect 315 1643 316 1647
rect 320 1643 321 1647
rect 310 1642 321 1643
rect 406 1647 417 1648
rect 406 1643 407 1647
rect 411 1643 412 1647
rect 416 1643 417 1647
rect 406 1642 417 1643
rect 502 1647 513 1648
rect 502 1643 503 1647
rect 507 1643 508 1647
rect 512 1643 513 1647
rect 502 1642 513 1643
rect 606 1647 617 1648
rect 606 1643 607 1647
rect 611 1643 612 1647
rect 616 1643 617 1647
rect 606 1642 617 1643
rect 707 1647 713 1648
rect 707 1643 708 1647
rect 712 1646 713 1647
rect 790 1647 801 1648
rect 712 1644 786 1646
rect 712 1643 713 1644
rect 707 1642 713 1643
rect 766 1639 772 1640
rect 766 1638 767 1639
rect 660 1636 767 1638
rect 660 1634 662 1636
rect 766 1635 767 1636
rect 771 1635 772 1639
rect 784 1638 786 1644
rect 790 1643 791 1647
rect 795 1643 796 1647
rect 800 1643 801 1647
rect 790 1642 801 1643
rect 870 1647 881 1648
rect 870 1643 871 1647
rect 875 1643 876 1647
rect 880 1643 881 1647
rect 870 1642 881 1643
rect 942 1647 953 1648
rect 942 1643 943 1647
rect 947 1643 948 1647
rect 952 1643 953 1647
rect 942 1642 953 1643
rect 1006 1647 1017 1648
rect 1006 1643 1007 1647
rect 1011 1643 1012 1647
rect 1016 1643 1017 1647
rect 1006 1642 1017 1643
rect 1078 1647 1089 1648
rect 1078 1643 1079 1647
rect 1083 1643 1084 1647
rect 1088 1643 1089 1647
rect 1078 1642 1089 1643
rect 1150 1647 1161 1648
rect 1150 1643 1151 1647
rect 1155 1643 1156 1647
rect 1160 1643 1161 1647
rect 1703 1647 1704 1651
rect 1708 1650 1709 1651
rect 1708 1648 1755 1650
rect 1708 1647 1709 1648
rect 1703 1646 1709 1647
rect 1753 1644 1755 1648
rect 1150 1642 1161 1643
rect 1327 1643 1333 1644
rect 1278 1640 1284 1641
rect 1022 1639 1028 1640
rect 1022 1638 1023 1639
rect 784 1636 1023 1638
rect 766 1634 772 1635
rect 1022 1635 1023 1636
rect 1027 1635 1028 1639
rect 1278 1636 1279 1640
rect 1283 1636 1284 1640
rect 1327 1639 1328 1643
rect 1332 1642 1333 1643
rect 1350 1643 1356 1644
rect 1350 1642 1351 1643
rect 1332 1640 1351 1642
rect 1332 1639 1333 1640
rect 1327 1638 1333 1639
rect 1350 1639 1351 1640
rect 1355 1639 1356 1643
rect 1350 1638 1356 1639
rect 1383 1643 1389 1644
rect 1383 1639 1384 1643
rect 1388 1642 1389 1643
rect 1438 1643 1444 1644
rect 1438 1642 1439 1643
rect 1388 1640 1439 1642
rect 1388 1639 1389 1640
rect 1383 1638 1389 1639
rect 1438 1639 1439 1640
rect 1443 1639 1444 1643
rect 1438 1638 1444 1639
rect 1454 1643 1460 1644
rect 1454 1639 1455 1643
rect 1459 1642 1460 1643
rect 1471 1643 1477 1644
rect 1471 1642 1472 1643
rect 1459 1640 1472 1642
rect 1459 1639 1460 1640
rect 1454 1638 1460 1639
rect 1471 1639 1472 1640
rect 1476 1639 1477 1643
rect 1471 1638 1477 1639
rect 1567 1643 1573 1644
rect 1567 1639 1568 1643
rect 1572 1642 1573 1643
rect 1630 1643 1636 1644
rect 1630 1642 1631 1643
rect 1572 1640 1631 1642
rect 1572 1639 1573 1640
rect 1567 1638 1573 1639
rect 1630 1639 1631 1640
rect 1635 1639 1636 1643
rect 1630 1638 1636 1639
rect 1663 1643 1669 1644
rect 1663 1639 1664 1643
rect 1668 1642 1669 1643
rect 1718 1643 1724 1644
rect 1718 1642 1719 1643
rect 1668 1640 1719 1642
rect 1668 1639 1669 1640
rect 1663 1638 1669 1639
rect 1718 1639 1719 1640
rect 1723 1639 1724 1643
rect 1718 1638 1724 1639
rect 1751 1643 1757 1644
rect 1751 1639 1752 1643
rect 1756 1639 1757 1643
rect 1751 1638 1757 1639
rect 1839 1643 1845 1644
rect 1839 1639 1840 1643
rect 1844 1642 1845 1643
rect 1886 1643 1892 1644
rect 1886 1642 1887 1643
rect 1844 1640 1887 1642
rect 1844 1639 1845 1640
rect 1839 1638 1845 1639
rect 1886 1639 1887 1640
rect 1891 1639 1892 1643
rect 1886 1638 1892 1639
rect 1919 1643 1925 1644
rect 1919 1639 1920 1643
rect 1924 1642 1925 1643
rect 1958 1643 1964 1644
rect 1958 1642 1959 1643
rect 1924 1640 1959 1642
rect 1924 1639 1925 1640
rect 1919 1638 1925 1639
rect 1958 1639 1959 1640
rect 1963 1639 1964 1643
rect 1958 1638 1964 1639
rect 1991 1643 1997 1644
rect 1991 1639 1992 1643
rect 1996 1642 1997 1643
rect 2022 1643 2028 1644
rect 2022 1642 2023 1643
rect 1996 1640 2023 1642
rect 1996 1639 1997 1640
rect 1991 1638 1997 1639
rect 2022 1639 2023 1640
rect 2027 1639 2028 1643
rect 2022 1638 2028 1639
rect 2055 1643 2061 1644
rect 2055 1639 2056 1643
rect 2060 1642 2061 1643
rect 2086 1643 2092 1644
rect 2086 1642 2087 1643
rect 2060 1640 2087 1642
rect 2060 1639 2061 1640
rect 2055 1638 2061 1639
rect 2086 1639 2087 1640
rect 2091 1639 2092 1643
rect 2086 1638 2092 1639
rect 2119 1643 2125 1644
rect 2119 1639 2120 1643
rect 2124 1642 2125 1643
rect 2150 1643 2156 1644
rect 2150 1642 2151 1643
rect 2124 1640 2151 1642
rect 2124 1639 2125 1640
rect 2119 1638 2125 1639
rect 2150 1639 2151 1640
rect 2155 1639 2156 1643
rect 2150 1638 2156 1639
rect 2183 1643 2189 1644
rect 2183 1639 2184 1643
rect 2188 1642 2189 1643
rect 2206 1643 2212 1644
rect 2206 1642 2207 1643
rect 2188 1640 2207 1642
rect 2188 1639 2189 1640
rect 2183 1638 2189 1639
rect 2206 1639 2207 1640
rect 2211 1639 2212 1643
rect 2247 1643 2253 1644
rect 2247 1642 2248 1643
rect 2206 1638 2212 1639
rect 2216 1640 2248 1642
rect 1278 1635 1284 1636
rect 1918 1635 1924 1636
rect 1022 1634 1028 1635
rect 659 1633 665 1634
rect 267 1631 273 1632
rect 267 1627 268 1631
rect 272 1630 273 1631
rect 278 1631 284 1632
rect 278 1630 279 1631
rect 272 1628 279 1630
rect 272 1627 273 1628
rect 267 1626 273 1627
rect 278 1627 279 1628
rect 283 1627 284 1631
rect 278 1626 284 1627
rect 298 1631 304 1632
rect 298 1627 299 1631
rect 303 1630 304 1631
rect 307 1631 313 1632
rect 307 1630 308 1631
rect 303 1628 308 1630
rect 303 1627 304 1628
rect 298 1626 304 1627
rect 307 1627 308 1628
rect 312 1627 313 1631
rect 307 1626 313 1627
rect 338 1631 344 1632
rect 338 1627 339 1631
rect 343 1630 344 1631
rect 355 1631 361 1632
rect 355 1630 356 1631
rect 343 1628 356 1630
rect 343 1627 344 1628
rect 338 1626 344 1627
rect 355 1627 356 1628
rect 360 1627 361 1631
rect 355 1626 361 1627
rect 394 1631 400 1632
rect 394 1627 395 1631
rect 399 1630 400 1631
rect 411 1631 417 1632
rect 411 1630 412 1631
rect 399 1628 412 1630
rect 399 1627 400 1628
rect 394 1626 400 1627
rect 411 1627 412 1628
rect 416 1627 417 1631
rect 411 1626 417 1627
rect 442 1631 448 1632
rect 442 1627 443 1631
rect 447 1630 448 1631
rect 467 1631 473 1632
rect 467 1630 468 1631
rect 447 1628 468 1630
rect 447 1627 448 1628
rect 442 1626 448 1627
rect 467 1627 468 1628
rect 472 1627 473 1631
rect 467 1626 473 1627
rect 498 1631 504 1632
rect 498 1627 499 1631
rect 503 1630 504 1631
rect 531 1631 537 1632
rect 531 1630 532 1631
rect 503 1628 532 1630
rect 503 1627 504 1628
rect 498 1626 504 1627
rect 531 1627 532 1628
rect 536 1627 537 1631
rect 531 1626 537 1627
rect 562 1631 568 1632
rect 562 1627 563 1631
rect 567 1630 568 1631
rect 595 1631 601 1632
rect 595 1630 596 1631
rect 567 1628 596 1630
rect 567 1627 568 1628
rect 562 1626 568 1627
rect 595 1627 596 1628
rect 600 1627 601 1631
rect 659 1629 660 1633
rect 664 1629 665 1633
rect 659 1628 665 1629
rect 690 1631 696 1632
rect 595 1626 601 1627
rect 690 1627 691 1631
rect 695 1630 696 1631
rect 715 1631 721 1632
rect 715 1630 716 1631
rect 695 1628 716 1630
rect 695 1627 696 1628
rect 690 1626 696 1627
rect 715 1627 716 1628
rect 720 1627 721 1631
rect 715 1626 721 1627
rect 746 1631 752 1632
rect 746 1627 747 1631
rect 751 1630 752 1631
rect 771 1631 777 1632
rect 771 1630 772 1631
rect 751 1628 772 1630
rect 751 1627 752 1628
rect 746 1626 752 1627
rect 771 1627 772 1628
rect 776 1627 777 1631
rect 771 1626 777 1627
rect 810 1631 816 1632
rect 810 1627 811 1631
rect 815 1630 816 1631
rect 827 1631 833 1632
rect 827 1630 828 1631
rect 815 1628 828 1630
rect 815 1627 816 1628
rect 810 1626 816 1627
rect 827 1627 828 1628
rect 832 1627 833 1631
rect 827 1626 833 1627
rect 858 1631 864 1632
rect 858 1627 859 1631
rect 863 1630 864 1631
rect 883 1631 889 1632
rect 883 1630 884 1631
rect 863 1628 884 1630
rect 863 1627 864 1628
rect 858 1626 864 1627
rect 883 1627 884 1628
rect 888 1627 889 1631
rect 883 1626 889 1627
rect 914 1631 920 1632
rect 914 1627 915 1631
rect 919 1630 920 1631
rect 939 1631 945 1632
rect 939 1630 940 1631
rect 919 1628 940 1630
rect 919 1627 920 1628
rect 914 1626 920 1627
rect 939 1627 940 1628
rect 944 1627 945 1631
rect 939 1626 945 1627
rect 970 1631 976 1632
rect 970 1627 971 1631
rect 975 1630 976 1631
rect 995 1631 1001 1632
rect 995 1630 996 1631
rect 975 1628 996 1630
rect 975 1627 976 1628
rect 970 1626 976 1627
rect 995 1627 996 1628
rect 1000 1627 1001 1631
rect 1918 1631 1919 1635
rect 1923 1634 1924 1635
rect 2216 1634 2218 1640
rect 2247 1639 2248 1640
rect 2252 1639 2253 1643
rect 2247 1638 2253 1639
rect 2406 1640 2412 1641
rect 2406 1636 2407 1640
rect 2411 1636 2412 1640
rect 2406 1635 2412 1636
rect 1923 1632 2218 1634
rect 1923 1631 1924 1632
rect 1918 1630 1924 1631
rect 995 1626 1001 1627
rect 270 1623 276 1624
rect 270 1619 271 1623
rect 275 1619 276 1623
rect 270 1618 276 1619
rect 310 1623 316 1624
rect 310 1619 311 1623
rect 315 1619 316 1623
rect 310 1618 316 1619
rect 358 1623 364 1624
rect 358 1619 359 1623
rect 363 1619 364 1623
rect 358 1618 364 1619
rect 414 1623 420 1624
rect 414 1619 415 1623
rect 419 1619 420 1623
rect 414 1618 420 1619
rect 470 1623 476 1624
rect 470 1619 471 1623
rect 475 1619 476 1623
rect 470 1618 476 1619
rect 534 1623 540 1624
rect 534 1619 535 1623
rect 539 1619 540 1623
rect 534 1618 540 1619
rect 598 1623 604 1624
rect 598 1619 599 1623
rect 603 1619 604 1623
rect 598 1618 604 1619
rect 662 1623 668 1624
rect 662 1619 663 1623
rect 667 1619 668 1623
rect 662 1618 668 1619
rect 718 1623 724 1624
rect 718 1619 719 1623
rect 723 1619 724 1623
rect 718 1618 724 1619
rect 774 1623 780 1624
rect 774 1619 775 1623
rect 779 1619 780 1623
rect 774 1618 780 1619
rect 830 1623 836 1624
rect 830 1619 831 1623
rect 835 1619 836 1623
rect 830 1618 836 1619
rect 886 1623 892 1624
rect 886 1619 887 1623
rect 891 1619 892 1623
rect 886 1618 892 1619
rect 942 1623 948 1624
rect 942 1619 943 1623
rect 947 1619 948 1623
rect 942 1618 948 1619
rect 998 1623 1004 1624
rect 998 1619 999 1623
rect 1003 1619 1004 1623
rect 998 1618 1004 1619
rect 1302 1617 1308 1618
rect 1302 1613 1303 1617
rect 1307 1613 1308 1617
rect 1302 1612 1308 1613
rect 1358 1617 1364 1618
rect 1358 1613 1359 1617
rect 1363 1613 1364 1617
rect 1358 1612 1364 1613
rect 1446 1617 1452 1618
rect 1446 1613 1447 1617
rect 1451 1613 1452 1617
rect 1446 1612 1452 1613
rect 1542 1617 1548 1618
rect 1542 1613 1543 1617
rect 1547 1613 1548 1617
rect 1542 1612 1548 1613
rect 1638 1617 1644 1618
rect 1638 1613 1639 1617
rect 1643 1613 1644 1617
rect 1638 1612 1644 1613
rect 1726 1617 1732 1618
rect 1726 1613 1727 1617
rect 1731 1613 1732 1617
rect 1726 1612 1732 1613
rect 1814 1617 1820 1618
rect 1814 1613 1815 1617
rect 1819 1613 1820 1617
rect 1814 1612 1820 1613
rect 1894 1617 1900 1618
rect 1894 1613 1895 1617
rect 1899 1613 1900 1617
rect 1894 1612 1900 1613
rect 1966 1617 1972 1618
rect 1966 1613 1967 1617
rect 1971 1613 1972 1617
rect 1966 1612 1972 1613
rect 2030 1617 2036 1618
rect 2030 1613 2031 1617
rect 2035 1613 2036 1617
rect 2030 1612 2036 1613
rect 2094 1617 2100 1618
rect 2094 1613 2095 1617
rect 2099 1613 2100 1617
rect 2094 1612 2100 1613
rect 2158 1617 2164 1618
rect 2158 1613 2159 1617
rect 2163 1613 2164 1617
rect 2158 1612 2164 1613
rect 2222 1617 2228 1618
rect 2222 1613 2223 1617
rect 2227 1613 2228 1617
rect 2222 1612 2228 1613
rect 1299 1607 1305 1608
rect 1299 1603 1300 1607
rect 1304 1606 1305 1607
rect 1338 1607 1344 1608
rect 1338 1606 1339 1607
rect 1304 1604 1339 1606
rect 1304 1603 1305 1604
rect 1299 1602 1305 1603
rect 1338 1603 1339 1604
rect 1343 1603 1344 1607
rect 1338 1602 1344 1603
rect 1350 1607 1361 1608
rect 1350 1603 1351 1607
rect 1355 1603 1356 1607
rect 1360 1603 1361 1607
rect 1350 1602 1361 1603
rect 1438 1607 1449 1608
rect 1438 1603 1439 1607
rect 1443 1603 1444 1607
rect 1448 1603 1449 1607
rect 1438 1602 1449 1603
rect 1506 1607 1512 1608
rect 1506 1603 1507 1607
rect 1511 1606 1512 1607
rect 1539 1607 1545 1608
rect 1539 1606 1540 1607
rect 1511 1604 1540 1606
rect 1511 1603 1512 1604
rect 1506 1602 1512 1603
rect 1539 1603 1540 1604
rect 1544 1603 1545 1607
rect 1539 1602 1545 1603
rect 1630 1607 1641 1608
rect 1630 1603 1631 1607
rect 1635 1603 1636 1607
rect 1640 1603 1641 1607
rect 1630 1602 1641 1603
rect 1718 1607 1729 1608
rect 1718 1603 1719 1607
rect 1723 1603 1724 1607
rect 1728 1603 1729 1607
rect 1718 1602 1729 1603
rect 1811 1607 1817 1608
rect 1811 1603 1812 1607
rect 1816 1606 1817 1607
rect 1822 1607 1828 1608
rect 1822 1606 1823 1607
rect 1816 1604 1823 1606
rect 1816 1603 1817 1604
rect 1811 1602 1817 1603
rect 1822 1603 1823 1604
rect 1827 1603 1828 1607
rect 1822 1602 1828 1603
rect 1886 1607 1897 1608
rect 1886 1603 1887 1607
rect 1891 1603 1892 1607
rect 1896 1603 1897 1607
rect 1886 1602 1897 1603
rect 1958 1607 1969 1608
rect 1958 1603 1959 1607
rect 1963 1603 1964 1607
rect 1968 1603 1969 1607
rect 1958 1602 1969 1603
rect 2022 1607 2033 1608
rect 2022 1603 2023 1607
rect 2027 1603 2028 1607
rect 2032 1603 2033 1607
rect 2022 1602 2033 1603
rect 2086 1607 2097 1608
rect 2086 1603 2087 1607
rect 2091 1603 2092 1607
rect 2096 1603 2097 1607
rect 2086 1602 2097 1603
rect 2150 1607 2161 1608
rect 2150 1603 2151 1607
rect 2155 1603 2156 1607
rect 2160 1603 2161 1607
rect 2150 1602 2161 1603
rect 2206 1607 2212 1608
rect 2206 1603 2207 1607
rect 2211 1606 2212 1607
rect 2219 1607 2225 1608
rect 2219 1606 2220 1607
rect 2211 1604 2220 1606
rect 2211 1603 2212 1604
rect 2206 1602 2212 1603
rect 2219 1603 2220 1604
rect 2224 1603 2225 1607
rect 2219 1602 2225 1603
rect 110 1600 116 1601
rect 110 1596 111 1600
rect 115 1596 116 1600
rect 1238 1600 1244 1601
rect 1238 1596 1239 1600
rect 1243 1596 1244 1600
rect 110 1595 116 1596
rect 295 1595 304 1596
rect 295 1591 296 1595
rect 303 1591 304 1595
rect 295 1590 304 1591
rect 335 1595 344 1596
rect 335 1591 336 1595
rect 343 1591 344 1595
rect 335 1590 344 1591
rect 383 1595 389 1596
rect 383 1591 384 1595
rect 388 1594 389 1595
rect 394 1595 400 1596
rect 394 1594 395 1595
rect 388 1592 395 1594
rect 388 1591 389 1592
rect 383 1590 389 1591
rect 394 1591 395 1592
rect 399 1591 400 1595
rect 394 1590 400 1591
rect 439 1595 448 1596
rect 439 1591 440 1595
rect 447 1591 448 1595
rect 439 1590 448 1591
rect 495 1595 504 1596
rect 495 1591 496 1595
rect 503 1591 504 1595
rect 495 1590 504 1591
rect 559 1595 568 1596
rect 559 1591 560 1595
rect 567 1591 568 1595
rect 559 1590 568 1591
rect 623 1595 629 1596
rect 623 1591 624 1595
rect 628 1591 629 1595
rect 623 1590 629 1591
rect 687 1595 696 1596
rect 687 1591 688 1595
rect 695 1591 696 1595
rect 687 1590 696 1591
rect 743 1595 752 1596
rect 743 1591 744 1595
rect 751 1591 752 1595
rect 743 1590 752 1591
rect 799 1595 805 1596
rect 799 1591 800 1595
rect 804 1594 805 1595
rect 810 1595 816 1596
rect 810 1594 811 1595
rect 804 1592 811 1594
rect 804 1591 805 1592
rect 799 1590 805 1591
rect 810 1591 811 1592
rect 815 1591 816 1595
rect 810 1590 816 1591
rect 855 1595 864 1596
rect 855 1591 856 1595
rect 863 1591 864 1595
rect 855 1590 864 1591
rect 911 1595 920 1596
rect 911 1591 912 1595
rect 919 1591 920 1595
rect 911 1590 920 1591
rect 967 1595 976 1596
rect 967 1591 968 1595
rect 975 1591 976 1595
rect 967 1590 976 1591
rect 1022 1595 1029 1596
rect 1238 1595 1244 1596
rect 1323 1595 1329 1596
rect 1022 1591 1023 1595
rect 1028 1591 1029 1595
rect 1022 1590 1029 1591
rect 1323 1591 1324 1595
rect 1328 1594 1329 1595
rect 1382 1595 1388 1596
rect 1382 1594 1383 1595
rect 1328 1592 1383 1594
rect 1328 1591 1329 1592
rect 1323 1590 1329 1591
rect 1382 1591 1383 1592
rect 1387 1591 1388 1595
rect 1382 1590 1388 1591
rect 1395 1595 1401 1596
rect 1395 1591 1396 1595
rect 1400 1594 1401 1595
rect 1454 1595 1460 1596
rect 1454 1594 1455 1595
rect 1400 1592 1455 1594
rect 1400 1591 1401 1592
rect 1395 1590 1401 1591
rect 1454 1591 1455 1592
rect 1459 1591 1460 1595
rect 1454 1590 1460 1591
rect 1475 1595 1481 1596
rect 1475 1591 1476 1595
rect 1480 1594 1481 1595
rect 1554 1595 1560 1596
rect 1554 1594 1555 1595
rect 1480 1592 1555 1594
rect 1480 1591 1481 1592
rect 1475 1590 1481 1591
rect 1554 1591 1555 1592
rect 1559 1591 1560 1595
rect 1554 1590 1560 1591
rect 1563 1595 1569 1596
rect 1563 1591 1564 1595
rect 1568 1594 1569 1595
rect 1639 1595 1645 1596
rect 1639 1594 1640 1595
rect 1568 1592 1640 1594
rect 1568 1591 1569 1592
rect 1563 1590 1569 1591
rect 1639 1591 1640 1592
rect 1644 1591 1645 1595
rect 1639 1590 1645 1591
rect 1651 1595 1657 1596
rect 1651 1591 1652 1595
rect 1656 1594 1657 1595
rect 1718 1595 1724 1596
rect 1718 1594 1719 1595
rect 1656 1592 1719 1594
rect 1656 1591 1657 1592
rect 1651 1590 1657 1591
rect 1718 1591 1719 1592
rect 1723 1591 1724 1595
rect 1718 1590 1724 1591
rect 1739 1595 1745 1596
rect 1739 1591 1740 1595
rect 1744 1594 1745 1595
rect 1815 1595 1821 1596
rect 1815 1594 1816 1595
rect 1744 1592 1816 1594
rect 1744 1591 1745 1592
rect 1739 1590 1745 1591
rect 1815 1591 1816 1592
rect 1820 1591 1821 1595
rect 1815 1590 1821 1591
rect 1827 1595 1833 1596
rect 1827 1591 1828 1595
rect 1832 1594 1833 1595
rect 1879 1595 1885 1596
rect 1879 1594 1880 1595
rect 1832 1592 1880 1594
rect 1832 1591 1833 1592
rect 1827 1590 1833 1591
rect 1879 1591 1880 1592
rect 1884 1591 1885 1595
rect 1879 1590 1885 1591
rect 1907 1595 1913 1596
rect 1907 1591 1908 1595
rect 1912 1594 1913 1595
rect 1918 1595 1924 1596
rect 1918 1594 1919 1595
rect 1912 1592 1919 1594
rect 1912 1591 1913 1592
rect 1907 1590 1913 1591
rect 1918 1591 1919 1592
rect 1923 1591 1924 1595
rect 1918 1590 1924 1591
rect 1938 1595 1944 1596
rect 1938 1591 1939 1595
rect 1943 1594 1944 1595
rect 1979 1595 1985 1596
rect 1979 1594 1980 1595
rect 1943 1592 1980 1594
rect 1943 1591 1944 1592
rect 1938 1590 1944 1591
rect 1979 1591 1980 1592
rect 1984 1591 1985 1595
rect 1979 1590 1985 1591
rect 2010 1595 2016 1596
rect 2010 1591 2011 1595
rect 2015 1594 2016 1595
rect 2043 1595 2049 1596
rect 2043 1594 2044 1595
rect 2015 1592 2044 1594
rect 2015 1591 2016 1592
rect 2010 1590 2016 1591
rect 2043 1591 2044 1592
rect 2048 1591 2049 1595
rect 2043 1590 2049 1591
rect 2074 1595 2080 1596
rect 2074 1591 2075 1595
rect 2079 1594 2080 1595
rect 2107 1595 2113 1596
rect 2107 1594 2108 1595
rect 2079 1592 2108 1594
rect 2079 1591 2080 1592
rect 2074 1590 2080 1591
rect 2107 1591 2108 1592
rect 2112 1591 2113 1595
rect 2107 1590 2113 1591
rect 2150 1595 2156 1596
rect 2150 1591 2151 1595
rect 2155 1594 2156 1595
rect 2163 1595 2169 1596
rect 2163 1594 2164 1595
rect 2155 1592 2164 1594
rect 2155 1591 2156 1592
rect 2150 1590 2156 1591
rect 2163 1591 2164 1592
rect 2168 1591 2169 1595
rect 2163 1590 2169 1591
rect 2194 1595 2200 1596
rect 2194 1591 2195 1595
rect 2199 1594 2200 1595
rect 2211 1595 2217 1596
rect 2211 1594 2212 1595
rect 2199 1592 2212 1594
rect 2199 1591 2200 1592
rect 2194 1590 2200 1591
rect 2211 1591 2212 1592
rect 2216 1591 2217 1595
rect 2211 1590 2217 1591
rect 2242 1595 2248 1596
rect 2242 1591 2243 1595
rect 2247 1594 2248 1595
rect 2267 1595 2273 1596
rect 2267 1594 2268 1595
rect 2247 1592 2268 1594
rect 2247 1591 2248 1592
rect 2242 1590 2248 1591
rect 2267 1591 2268 1592
rect 2272 1591 2273 1595
rect 2267 1590 2273 1591
rect 2298 1595 2304 1596
rect 2298 1591 2299 1595
rect 2303 1594 2304 1595
rect 2315 1595 2321 1596
rect 2315 1594 2316 1595
rect 2303 1592 2316 1594
rect 2303 1591 2304 1592
rect 2298 1590 2304 1591
rect 2315 1591 2316 1592
rect 2320 1591 2321 1595
rect 2315 1590 2321 1591
rect 2346 1595 2352 1596
rect 2346 1591 2347 1595
rect 2351 1594 2352 1595
rect 2355 1595 2361 1596
rect 2355 1594 2356 1595
rect 2351 1592 2356 1594
rect 2351 1591 2352 1592
rect 2346 1590 2352 1591
rect 2355 1591 2356 1592
rect 2360 1591 2361 1595
rect 2355 1590 2361 1591
rect 346 1587 352 1588
rect 110 1583 116 1584
rect 110 1579 111 1583
rect 115 1579 116 1583
rect 346 1583 347 1587
rect 351 1586 352 1587
rect 625 1586 627 1590
rect 351 1584 627 1586
rect 766 1587 772 1588
rect 351 1583 352 1584
rect 346 1582 352 1583
rect 766 1583 767 1587
rect 771 1586 772 1587
rect 950 1587 956 1588
rect 950 1586 951 1587
rect 771 1584 951 1586
rect 771 1583 772 1584
rect 766 1582 772 1583
rect 950 1583 951 1584
rect 955 1583 956 1587
rect 1326 1587 1332 1588
rect 950 1582 956 1583
rect 1238 1583 1244 1584
rect 110 1578 116 1579
rect 1238 1579 1239 1583
rect 1243 1579 1244 1583
rect 1326 1583 1327 1587
rect 1331 1583 1332 1587
rect 1326 1582 1332 1583
rect 1398 1587 1404 1588
rect 1398 1583 1399 1587
rect 1403 1583 1404 1587
rect 1398 1582 1404 1583
rect 1478 1587 1484 1588
rect 1478 1583 1479 1587
rect 1483 1583 1484 1587
rect 1478 1582 1484 1583
rect 1566 1587 1572 1588
rect 1566 1583 1567 1587
rect 1571 1583 1572 1587
rect 1566 1582 1572 1583
rect 1654 1587 1660 1588
rect 1654 1583 1655 1587
rect 1659 1583 1660 1587
rect 1654 1582 1660 1583
rect 1742 1587 1748 1588
rect 1742 1583 1743 1587
rect 1747 1583 1748 1587
rect 1742 1582 1748 1583
rect 1830 1587 1836 1588
rect 1830 1583 1831 1587
rect 1835 1583 1836 1587
rect 1830 1582 1836 1583
rect 1910 1587 1916 1588
rect 1910 1583 1911 1587
rect 1915 1583 1916 1587
rect 1910 1582 1916 1583
rect 1982 1587 1988 1588
rect 1982 1583 1983 1587
rect 1987 1583 1988 1587
rect 1982 1582 1988 1583
rect 2046 1587 2052 1588
rect 2046 1583 2047 1587
rect 2051 1583 2052 1587
rect 2046 1582 2052 1583
rect 2110 1587 2116 1588
rect 2110 1583 2111 1587
rect 2115 1583 2116 1587
rect 2110 1582 2116 1583
rect 2166 1587 2172 1588
rect 2166 1583 2167 1587
rect 2171 1583 2172 1587
rect 2166 1582 2172 1583
rect 2214 1587 2220 1588
rect 2214 1583 2215 1587
rect 2219 1583 2220 1587
rect 2214 1582 2220 1583
rect 2270 1587 2276 1588
rect 2270 1583 2271 1587
rect 2275 1583 2276 1587
rect 2270 1582 2276 1583
rect 2318 1587 2324 1588
rect 2318 1583 2319 1587
rect 2323 1583 2324 1587
rect 2318 1582 2324 1583
rect 2358 1587 2364 1588
rect 2358 1583 2359 1587
rect 2363 1583 2364 1587
rect 2358 1582 2364 1583
rect 1238 1578 1244 1579
rect 270 1576 276 1577
rect 270 1572 271 1576
rect 275 1572 276 1576
rect 270 1571 276 1572
rect 310 1576 316 1577
rect 310 1572 311 1576
rect 315 1572 316 1576
rect 310 1571 316 1572
rect 358 1576 364 1577
rect 358 1572 359 1576
rect 363 1572 364 1576
rect 358 1571 364 1572
rect 414 1576 420 1577
rect 414 1572 415 1576
rect 419 1572 420 1576
rect 414 1571 420 1572
rect 470 1576 476 1577
rect 470 1572 471 1576
rect 475 1572 476 1576
rect 470 1571 476 1572
rect 534 1576 540 1577
rect 534 1572 535 1576
rect 539 1572 540 1576
rect 534 1571 540 1572
rect 598 1576 604 1577
rect 598 1572 599 1576
rect 603 1572 604 1576
rect 598 1571 604 1572
rect 662 1576 668 1577
rect 662 1572 663 1576
rect 667 1572 668 1576
rect 662 1571 668 1572
rect 718 1576 724 1577
rect 718 1572 719 1576
rect 723 1572 724 1576
rect 718 1571 724 1572
rect 774 1576 780 1577
rect 774 1572 775 1576
rect 779 1572 780 1576
rect 774 1571 780 1572
rect 830 1576 836 1577
rect 830 1572 831 1576
rect 835 1572 836 1576
rect 830 1571 836 1572
rect 886 1576 892 1577
rect 886 1572 887 1576
rect 891 1572 892 1576
rect 886 1571 892 1572
rect 942 1576 948 1577
rect 942 1572 943 1576
rect 947 1572 948 1576
rect 942 1571 948 1572
rect 998 1576 1004 1577
rect 998 1572 999 1576
rect 1003 1572 1004 1576
rect 998 1571 1004 1572
rect 1278 1564 1284 1565
rect 1278 1560 1279 1564
rect 1283 1560 1284 1564
rect 2406 1564 2412 1565
rect 2406 1560 2407 1564
rect 2411 1560 2412 1564
rect 1278 1559 1284 1560
rect 1342 1559 1348 1560
rect 326 1556 332 1557
rect 326 1552 327 1556
rect 331 1552 332 1556
rect 326 1551 332 1552
rect 366 1556 372 1557
rect 366 1552 367 1556
rect 371 1552 372 1556
rect 366 1551 372 1552
rect 406 1556 412 1557
rect 406 1552 407 1556
rect 411 1552 412 1556
rect 406 1551 412 1552
rect 446 1556 452 1557
rect 446 1552 447 1556
rect 451 1552 452 1556
rect 446 1551 452 1552
rect 486 1556 492 1557
rect 486 1552 487 1556
rect 491 1552 492 1556
rect 486 1551 492 1552
rect 526 1556 532 1557
rect 526 1552 527 1556
rect 531 1552 532 1556
rect 526 1551 532 1552
rect 566 1556 572 1557
rect 566 1552 567 1556
rect 571 1552 572 1556
rect 566 1551 572 1552
rect 606 1556 612 1557
rect 606 1552 607 1556
rect 611 1552 612 1556
rect 606 1551 612 1552
rect 646 1556 652 1557
rect 646 1552 647 1556
rect 651 1552 652 1556
rect 646 1551 652 1552
rect 686 1556 692 1557
rect 686 1552 687 1556
rect 691 1552 692 1556
rect 686 1551 692 1552
rect 726 1556 732 1557
rect 726 1552 727 1556
rect 731 1552 732 1556
rect 726 1551 732 1552
rect 766 1556 772 1557
rect 766 1552 767 1556
rect 771 1552 772 1556
rect 766 1551 772 1552
rect 806 1556 812 1557
rect 806 1552 807 1556
rect 811 1552 812 1556
rect 806 1551 812 1552
rect 846 1556 852 1557
rect 846 1552 847 1556
rect 851 1552 852 1556
rect 846 1551 852 1552
rect 886 1556 892 1557
rect 886 1552 887 1556
rect 891 1552 892 1556
rect 886 1551 892 1552
rect 926 1556 932 1557
rect 926 1552 927 1556
rect 931 1552 932 1556
rect 1342 1555 1343 1559
rect 1347 1558 1348 1559
rect 1351 1559 1357 1560
rect 1351 1558 1352 1559
rect 1347 1556 1352 1558
rect 1347 1555 1348 1556
rect 1342 1554 1348 1555
rect 1351 1555 1352 1556
rect 1356 1555 1357 1559
rect 1351 1554 1357 1555
rect 1382 1559 1388 1560
rect 1382 1555 1383 1559
rect 1387 1558 1388 1559
rect 1423 1559 1429 1560
rect 1423 1558 1424 1559
rect 1387 1556 1424 1558
rect 1387 1555 1388 1556
rect 1382 1554 1388 1555
rect 1423 1555 1424 1556
rect 1428 1555 1429 1559
rect 1423 1554 1429 1555
rect 1503 1559 1512 1560
rect 1503 1555 1504 1559
rect 1511 1555 1512 1559
rect 1503 1554 1512 1555
rect 1554 1559 1560 1560
rect 1554 1555 1555 1559
rect 1559 1558 1560 1559
rect 1591 1559 1597 1560
rect 1591 1558 1592 1559
rect 1559 1556 1592 1558
rect 1559 1555 1560 1556
rect 1554 1554 1560 1555
rect 1591 1555 1592 1556
rect 1596 1555 1597 1559
rect 1591 1554 1597 1555
rect 1639 1559 1645 1560
rect 1639 1555 1640 1559
rect 1644 1558 1645 1559
rect 1679 1559 1685 1560
rect 1679 1558 1680 1559
rect 1644 1556 1680 1558
rect 1644 1555 1645 1556
rect 1639 1554 1645 1555
rect 1679 1555 1680 1556
rect 1684 1555 1685 1559
rect 1679 1554 1685 1555
rect 1718 1559 1724 1560
rect 1718 1555 1719 1559
rect 1723 1558 1724 1559
rect 1767 1559 1773 1560
rect 1767 1558 1768 1559
rect 1723 1556 1768 1558
rect 1723 1555 1724 1556
rect 1718 1554 1724 1555
rect 1767 1555 1768 1556
rect 1772 1555 1773 1559
rect 1767 1554 1773 1555
rect 1815 1559 1821 1560
rect 1815 1555 1816 1559
rect 1820 1558 1821 1559
rect 1855 1559 1861 1560
rect 1855 1558 1856 1559
rect 1820 1556 1856 1558
rect 1820 1555 1821 1556
rect 1815 1554 1821 1555
rect 1855 1555 1856 1556
rect 1860 1555 1861 1559
rect 1855 1554 1861 1555
rect 1935 1559 1944 1560
rect 1935 1555 1936 1559
rect 1943 1555 1944 1559
rect 1935 1554 1944 1555
rect 2007 1559 2016 1560
rect 2007 1555 2008 1559
rect 2015 1555 2016 1559
rect 2007 1554 2016 1555
rect 2071 1559 2080 1560
rect 2071 1555 2072 1559
rect 2079 1555 2080 1559
rect 2071 1554 2080 1555
rect 2135 1559 2141 1560
rect 2135 1555 2136 1559
rect 2140 1558 2141 1559
rect 2150 1559 2156 1560
rect 2150 1558 2151 1559
rect 2140 1556 2151 1558
rect 2140 1555 2141 1556
rect 2135 1554 2141 1555
rect 2150 1555 2151 1556
rect 2155 1555 2156 1559
rect 2150 1554 2156 1555
rect 2191 1559 2200 1560
rect 2191 1555 2192 1559
rect 2199 1555 2200 1559
rect 2191 1554 2200 1555
rect 2239 1559 2248 1560
rect 2239 1555 2240 1559
rect 2247 1555 2248 1559
rect 2239 1554 2248 1555
rect 2295 1559 2304 1560
rect 2295 1555 2296 1559
rect 2303 1555 2304 1559
rect 2295 1554 2304 1555
rect 2343 1559 2352 1560
rect 2343 1555 2344 1559
rect 2351 1555 2352 1559
rect 2383 1559 2389 1560
rect 2406 1559 2412 1560
rect 2383 1558 2384 1559
rect 2343 1554 2352 1555
rect 2356 1556 2384 1558
rect 926 1551 932 1552
rect 2222 1551 2228 1552
rect 110 1549 116 1550
rect 110 1545 111 1549
rect 115 1545 116 1549
rect 110 1544 116 1545
rect 1238 1549 1244 1550
rect 1238 1545 1239 1549
rect 1243 1545 1244 1549
rect 1238 1544 1244 1545
rect 1278 1547 1284 1548
rect 1278 1543 1279 1547
rect 1283 1543 1284 1547
rect 2222 1547 2223 1551
rect 2227 1550 2228 1551
rect 2356 1550 2358 1556
rect 2383 1555 2384 1556
rect 2388 1555 2389 1559
rect 2383 1554 2389 1555
rect 2227 1548 2358 1550
rect 2227 1547 2228 1548
rect 2222 1546 2228 1547
rect 2406 1547 2412 1548
rect 1278 1542 1284 1543
rect 2406 1543 2407 1547
rect 2411 1543 2412 1547
rect 2406 1542 2412 1543
rect 1326 1540 1332 1541
rect 1326 1536 1327 1540
rect 1331 1536 1332 1540
rect 351 1535 360 1536
rect 110 1532 116 1533
rect 110 1528 111 1532
rect 115 1528 116 1532
rect 351 1531 352 1535
rect 359 1531 360 1535
rect 351 1530 360 1531
rect 391 1535 400 1536
rect 391 1531 392 1535
rect 399 1531 400 1535
rect 391 1530 400 1531
rect 431 1535 440 1536
rect 431 1531 432 1535
rect 439 1531 440 1535
rect 431 1530 440 1531
rect 471 1535 480 1536
rect 471 1531 472 1535
rect 479 1531 480 1535
rect 471 1530 480 1531
rect 511 1535 520 1536
rect 511 1531 512 1535
rect 519 1531 520 1535
rect 511 1530 520 1531
rect 551 1535 560 1536
rect 551 1531 552 1535
rect 559 1531 560 1535
rect 551 1530 560 1531
rect 591 1535 600 1536
rect 591 1531 592 1535
rect 599 1531 600 1535
rect 591 1530 600 1531
rect 631 1535 640 1536
rect 631 1531 632 1535
rect 639 1531 640 1535
rect 631 1530 640 1531
rect 671 1535 680 1536
rect 671 1531 672 1535
rect 679 1531 680 1535
rect 671 1530 680 1531
rect 711 1535 720 1536
rect 711 1531 712 1535
rect 719 1531 720 1535
rect 711 1530 720 1531
rect 751 1535 760 1536
rect 751 1531 752 1535
rect 759 1531 760 1535
rect 751 1530 760 1531
rect 791 1535 800 1536
rect 791 1531 792 1535
rect 799 1531 800 1535
rect 791 1530 800 1531
rect 831 1535 840 1536
rect 831 1531 832 1535
rect 839 1531 840 1535
rect 831 1530 840 1531
rect 871 1535 880 1536
rect 871 1531 872 1535
rect 879 1531 880 1535
rect 871 1530 880 1531
rect 911 1535 920 1536
rect 911 1531 912 1535
rect 919 1531 920 1535
rect 911 1530 920 1531
rect 950 1535 957 1536
rect 1326 1535 1332 1536
rect 1398 1540 1404 1541
rect 1398 1536 1399 1540
rect 1403 1536 1404 1540
rect 1398 1535 1404 1536
rect 1478 1540 1484 1541
rect 1478 1536 1479 1540
rect 1483 1536 1484 1540
rect 1478 1535 1484 1536
rect 1566 1540 1572 1541
rect 1566 1536 1567 1540
rect 1571 1536 1572 1540
rect 1566 1535 1572 1536
rect 1654 1540 1660 1541
rect 1654 1536 1655 1540
rect 1659 1536 1660 1540
rect 1654 1535 1660 1536
rect 1742 1540 1748 1541
rect 1742 1536 1743 1540
rect 1747 1536 1748 1540
rect 1742 1535 1748 1536
rect 1830 1540 1836 1541
rect 1830 1536 1831 1540
rect 1835 1536 1836 1540
rect 1830 1535 1836 1536
rect 1910 1540 1916 1541
rect 1910 1536 1911 1540
rect 1915 1536 1916 1540
rect 1910 1535 1916 1536
rect 1982 1540 1988 1541
rect 1982 1536 1983 1540
rect 1987 1536 1988 1540
rect 1982 1535 1988 1536
rect 2046 1540 2052 1541
rect 2046 1536 2047 1540
rect 2051 1536 2052 1540
rect 2046 1535 2052 1536
rect 2110 1540 2116 1541
rect 2110 1536 2111 1540
rect 2115 1536 2116 1540
rect 2110 1535 2116 1536
rect 2166 1540 2172 1541
rect 2166 1536 2167 1540
rect 2171 1536 2172 1540
rect 2166 1535 2172 1536
rect 2214 1540 2220 1541
rect 2214 1536 2215 1540
rect 2219 1536 2220 1540
rect 2214 1535 2220 1536
rect 2270 1540 2276 1541
rect 2270 1536 2271 1540
rect 2275 1536 2276 1540
rect 2270 1535 2276 1536
rect 2318 1540 2324 1541
rect 2318 1536 2319 1540
rect 2323 1536 2324 1540
rect 2318 1535 2324 1536
rect 2358 1540 2364 1541
rect 2358 1536 2359 1540
rect 2363 1536 2364 1540
rect 2358 1535 2364 1536
rect 950 1531 951 1535
rect 956 1531 957 1535
rect 950 1530 957 1531
rect 1238 1532 1244 1533
rect 110 1527 116 1528
rect 1238 1528 1239 1532
rect 1243 1528 1244 1532
rect 1238 1527 1244 1528
rect 1334 1524 1340 1525
rect 1334 1520 1335 1524
rect 1339 1520 1340 1524
rect 1334 1519 1340 1520
rect 1414 1524 1420 1525
rect 1414 1520 1415 1524
rect 1419 1520 1420 1524
rect 1414 1519 1420 1520
rect 1502 1524 1508 1525
rect 1502 1520 1503 1524
rect 1507 1520 1508 1524
rect 1502 1519 1508 1520
rect 1614 1524 1620 1525
rect 1614 1520 1615 1524
rect 1619 1520 1620 1524
rect 1614 1519 1620 1520
rect 1742 1524 1748 1525
rect 1742 1520 1743 1524
rect 1747 1520 1748 1524
rect 1742 1519 1748 1520
rect 1886 1524 1892 1525
rect 1886 1520 1887 1524
rect 1891 1520 1892 1524
rect 1886 1519 1892 1520
rect 2046 1524 2052 1525
rect 2046 1520 2047 1524
rect 2051 1520 2052 1524
rect 2046 1519 2052 1520
rect 2214 1524 2220 1525
rect 2214 1520 2215 1524
rect 2219 1520 2220 1524
rect 2214 1519 2220 1520
rect 2358 1524 2364 1525
rect 2358 1520 2359 1524
rect 2363 1520 2364 1524
rect 2358 1519 2364 1520
rect 1278 1517 1284 1518
rect 1278 1513 1279 1517
rect 1283 1513 1284 1517
rect 2406 1517 2412 1518
rect 1278 1512 1284 1513
rect 1879 1515 1885 1516
rect 1879 1511 1880 1515
rect 1884 1514 1885 1515
rect 1884 1512 2001 1514
rect 2406 1513 2407 1517
rect 2411 1513 2412 1517
rect 2406 1512 2412 1513
rect 1884 1511 1885 1512
rect 1879 1510 1885 1511
rect 1999 1510 2001 1512
rect 326 1509 332 1510
rect 326 1505 327 1509
rect 331 1505 332 1509
rect 326 1504 332 1505
rect 366 1509 372 1510
rect 366 1505 367 1509
rect 371 1505 372 1509
rect 366 1504 372 1505
rect 406 1509 412 1510
rect 406 1505 407 1509
rect 411 1505 412 1509
rect 406 1504 412 1505
rect 446 1509 452 1510
rect 446 1505 447 1509
rect 451 1505 452 1509
rect 446 1504 452 1505
rect 486 1509 492 1510
rect 486 1505 487 1509
rect 491 1505 492 1509
rect 486 1504 492 1505
rect 526 1509 532 1510
rect 526 1505 527 1509
rect 531 1505 532 1509
rect 526 1504 532 1505
rect 566 1509 572 1510
rect 566 1505 567 1509
rect 571 1505 572 1509
rect 566 1504 572 1505
rect 606 1509 612 1510
rect 606 1505 607 1509
rect 611 1505 612 1509
rect 606 1504 612 1505
rect 646 1509 652 1510
rect 646 1505 647 1509
rect 651 1505 652 1509
rect 646 1504 652 1505
rect 686 1509 692 1510
rect 686 1505 687 1509
rect 691 1505 692 1509
rect 686 1504 692 1505
rect 726 1509 732 1510
rect 726 1505 727 1509
rect 731 1505 732 1509
rect 726 1504 732 1505
rect 766 1509 772 1510
rect 766 1505 767 1509
rect 771 1505 772 1509
rect 766 1504 772 1505
rect 806 1509 812 1510
rect 806 1505 807 1509
rect 811 1505 812 1509
rect 806 1504 812 1505
rect 846 1509 852 1510
rect 846 1505 847 1509
rect 851 1505 852 1509
rect 846 1504 852 1505
rect 886 1509 892 1510
rect 886 1505 887 1509
rect 891 1505 892 1509
rect 886 1504 892 1505
rect 926 1509 932 1510
rect 926 1505 927 1509
rect 931 1505 932 1509
rect 1999 1508 2050 1510
rect 926 1504 932 1505
rect 1359 1503 1365 1504
rect 1278 1500 1284 1501
rect 323 1499 329 1500
rect 323 1495 324 1499
rect 328 1498 329 1499
rect 346 1499 352 1500
rect 346 1498 347 1499
rect 328 1496 347 1498
rect 328 1495 329 1496
rect 323 1494 329 1495
rect 346 1495 347 1496
rect 351 1495 352 1499
rect 346 1494 352 1495
rect 354 1499 360 1500
rect 354 1495 355 1499
rect 359 1498 360 1499
rect 363 1499 369 1500
rect 363 1498 364 1499
rect 359 1496 364 1498
rect 359 1495 360 1496
rect 354 1494 360 1495
rect 363 1495 364 1496
rect 368 1495 369 1499
rect 363 1494 369 1495
rect 394 1499 400 1500
rect 394 1495 395 1499
rect 399 1498 400 1499
rect 403 1499 409 1500
rect 403 1498 404 1499
rect 399 1496 404 1498
rect 399 1495 400 1496
rect 394 1494 400 1495
rect 403 1495 404 1496
rect 408 1495 409 1499
rect 403 1494 409 1495
rect 434 1499 440 1500
rect 434 1495 435 1499
rect 439 1498 440 1499
rect 443 1499 449 1500
rect 443 1498 444 1499
rect 439 1496 444 1498
rect 439 1495 440 1496
rect 434 1494 440 1495
rect 443 1495 444 1496
rect 448 1495 449 1499
rect 443 1494 449 1495
rect 474 1499 480 1500
rect 474 1495 475 1499
rect 479 1498 480 1499
rect 483 1499 489 1500
rect 483 1498 484 1499
rect 479 1496 484 1498
rect 479 1495 480 1496
rect 474 1494 480 1495
rect 483 1495 484 1496
rect 488 1495 489 1499
rect 483 1494 489 1495
rect 514 1499 520 1500
rect 514 1495 515 1499
rect 519 1498 520 1499
rect 523 1499 529 1500
rect 523 1498 524 1499
rect 519 1496 524 1498
rect 519 1495 520 1496
rect 514 1494 520 1495
rect 523 1495 524 1496
rect 528 1495 529 1499
rect 523 1494 529 1495
rect 554 1499 560 1500
rect 554 1495 555 1499
rect 559 1498 560 1499
rect 563 1499 569 1500
rect 563 1498 564 1499
rect 559 1496 564 1498
rect 559 1495 560 1496
rect 554 1494 560 1495
rect 563 1495 564 1496
rect 568 1495 569 1499
rect 563 1494 569 1495
rect 594 1499 600 1500
rect 594 1495 595 1499
rect 599 1498 600 1499
rect 603 1499 609 1500
rect 603 1498 604 1499
rect 599 1496 604 1498
rect 599 1495 600 1496
rect 594 1494 600 1495
rect 603 1495 604 1496
rect 608 1495 609 1499
rect 603 1494 609 1495
rect 634 1499 640 1500
rect 634 1495 635 1499
rect 639 1498 640 1499
rect 643 1499 649 1500
rect 643 1498 644 1499
rect 639 1496 644 1498
rect 639 1495 640 1496
rect 634 1494 640 1495
rect 643 1495 644 1496
rect 648 1495 649 1499
rect 643 1494 649 1495
rect 674 1499 680 1500
rect 674 1495 675 1499
rect 679 1498 680 1499
rect 683 1499 689 1500
rect 683 1498 684 1499
rect 679 1496 684 1498
rect 679 1495 680 1496
rect 674 1494 680 1495
rect 683 1495 684 1496
rect 688 1495 689 1499
rect 683 1494 689 1495
rect 714 1499 720 1500
rect 714 1495 715 1499
rect 719 1498 720 1499
rect 723 1499 729 1500
rect 723 1498 724 1499
rect 719 1496 724 1498
rect 719 1495 720 1496
rect 714 1494 720 1495
rect 723 1495 724 1496
rect 728 1495 729 1499
rect 723 1494 729 1495
rect 754 1499 760 1500
rect 754 1495 755 1499
rect 759 1498 760 1499
rect 763 1499 769 1500
rect 763 1498 764 1499
rect 759 1496 764 1498
rect 759 1495 760 1496
rect 754 1494 760 1495
rect 763 1495 764 1496
rect 768 1495 769 1499
rect 763 1494 769 1495
rect 794 1499 800 1500
rect 794 1495 795 1499
rect 799 1498 800 1499
rect 803 1499 809 1500
rect 803 1498 804 1499
rect 799 1496 804 1498
rect 799 1495 800 1496
rect 794 1494 800 1495
rect 803 1495 804 1496
rect 808 1495 809 1499
rect 803 1494 809 1495
rect 834 1499 840 1500
rect 834 1495 835 1499
rect 839 1498 840 1499
rect 843 1499 849 1500
rect 843 1498 844 1499
rect 839 1496 844 1498
rect 839 1495 840 1496
rect 834 1494 840 1495
rect 843 1495 844 1496
rect 848 1495 849 1499
rect 843 1494 849 1495
rect 874 1499 880 1500
rect 874 1495 875 1499
rect 879 1498 880 1499
rect 883 1499 889 1500
rect 883 1498 884 1499
rect 879 1496 884 1498
rect 879 1495 880 1496
rect 874 1494 880 1495
rect 883 1495 884 1496
rect 888 1495 889 1499
rect 883 1494 889 1495
rect 914 1499 920 1500
rect 914 1495 915 1499
rect 919 1498 920 1499
rect 923 1499 929 1500
rect 923 1498 924 1499
rect 919 1496 924 1498
rect 919 1495 920 1496
rect 914 1494 920 1495
rect 923 1495 924 1496
rect 928 1495 929 1499
rect 1278 1496 1279 1500
rect 1283 1496 1284 1500
rect 1359 1499 1360 1503
rect 1364 1502 1365 1503
rect 1406 1503 1412 1504
rect 1406 1502 1407 1503
rect 1364 1500 1407 1502
rect 1364 1499 1365 1500
rect 1359 1498 1365 1499
rect 1406 1499 1407 1500
rect 1411 1499 1412 1503
rect 1406 1498 1412 1499
rect 1439 1503 1445 1504
rect 1439 1499 1440 1503
rect 1444 1502 1445 1503
rect 1486 1503 1492 1504
rect 1486 1502 1487 1503
rect 1444 1500 1487 1502
rect 1444 1499 1445 1500
rect 1439 1498 1445 1499
rect 1486 1499 1487 1500
rect 1491 1499 1492 1503
rect 1486 1498 1492 1499
rect 1494 1503 1500 1504
rect 1494 1499 1495 1503
rect 1499 1502 1500 1503
rect 1527 1503 1533 1504
rect 1527 1502 1528 1503
rect 1499 1500 1528 1502
rect 1499 1499 1500 1500
rect 1494 1498 1500 1499
rect 1527 1499 1528 1500
rect 1532 1499 1533 1503
rect 1527 1498 1533 1499
rect 1639 1503 1645 1504
rect 1639 1499 1640 1503
rect 1644 1502 1645 1503
rect 1734 1503 1740 1504
rect 1734 1502 1735 1503
rect 1644 1500 1735 1502
rect 1644 1499 1645 1500
rect 1639 1498 1645 1499
rect 1734 1499 1735 1500
rect 1739 1499 1740 1503
rect 1734 1498 1740 1499
rect 1767 1503 1773 1504
rect 1767 1499 1768 1503
rect 1772 1502 1773 1503
rect 1871 1503 1877 1504
rect 1871 1502 1872 1503
rect 1772 1500 1872 1502
rect 1772 1499 1773 1500
rect 1767 1498 1773 1499
rect 1871 1499 1872 1500
rect 1876 1499 1877 1503
rect 1871 1498 1877 1499
rect 1911 1503 1917 1504
rect 1911 1499 1912 1503
rect 1916 1502 1917 1503
rect 2038 1503 2044 1504
rect 2038 1502 2039 1503
rect 1916 1500 2039 1502
rect 1916 1499 1917 1500
rect 1911 1498 1917 1499
rect 2038 1499 2039 1500
rect 2043 1499 2044 1503
rect 2048 1502 2050 1508
rect 2071 1503 2077 1504
rect 2071 1502 2072 1503
rect 2048 1500 2072 1502
rect 2038 1498 2044 1499
rect 2071 1499 2072 1500
rect 2076 1499 2077 1503
rect 2071 1498 2077 1499
rect 2239 1503 2245 1504
rect 2239 1499 2240 1503
rect 2244 1502 2245 1503
rect 2350 1503 2356 1504
rect 2350 1502 2351 1503
rect 2244 1500 2351 1502
rect 2244 1499 2245 1500
rect 2239 1498 2245 1499
rect 2350 1499 2351 1500
rect 2355 1499 2356 1503
rect 2350 1498 2356 1499
rect 2366 1503 2372 1504
rect 2366 1499 2367 1503
rect 2371 1502 2372 1503
rect 2383 1503 2389 1504
rect 2383 1502 2384 1503
rect 2371 1500 2384 1502
rect 2371 1499 2372 1500
rect 2366 1498 2372 1499
rect 2383 1499 2384 1500
rect 2388 1499 2389 1503
rect 2383 1498 2389 1499
rect 2406 1500 2412 1501
rect 1278 1495 1284 1496
rect 2406 1496 2407 1500
rect 2411 1496 2412 1500
rect 2406 1495 2412 1496
rect 923 1494 929 1495
rect 1334 1477 1340 1478
rect 1334 1473 1335 1477
rect 1339 1473 1340 1477
rect 1334 1472 1340 1473
rect 1414 1477 1420 1478
rect 1414 1473 1415 1477
rect 1419 1473 1420 1477
rect 1414 1472 1420 1473
rect 1502 1477 1508 1478
rect 1502 1473 1503 1477
rect 1507 1473 1508 1477
rect 1502 1472 1508 1473
rect 1614 1477 1620 1478
rect 1614 1473 1615 1477
rect 1619 1473 1620 1477
rect 1614 1472 1620 1473
rect 1742 1477 1748 1478
rect 1742 1473 1743 1477
rect 1747 1473 1748 1477
rect 1742 1472 1748 1473
rect 1886 1477 1892 1478
rect 1886 1473 1887 1477
rect 1891 1473 1892 1477
rect 1886 1472 1892 1473
rect 2046 1477 2052 1478
rect 2046 1473 2047 1477
rect 2051 1473 2052 1477
rect 2046 1472 2052 1473
rect 2214 1477 2220 1478
rect 2214 1473 2215 1477
rect 2219 1473 2220 1477
rect 2214 1472 2220 1473
rect 2358 1477 2364 1478
rect 2358 1473 2359 1477
rect 2363 1473 2364 1477
rect 2358 1472 2364 1473
rect 1331 1467 1337 1468
rect 1331 1463 1332 1467
rect 1336 1466 1337 1467
rect 1342 1467 1348 1468
rect 1342 1466 1343 1467
rect 1336 1464 1343 1466
rect 1336 1463 1337 1464
rect 1331 1462 1337 1463
rect 1342 1463 1343 1464
rect 1347 1463 1348 1467
rect 1342 1462 1348 1463
rect 1406 1467 1417 1468
rect 1406 1463 1407 1467
rect 1411 1463 1412 1467
rect 1416 1463 1417 1467
rect 1406 1462 1417 1463
rect 1486 1467 1492 1468
rect 1486 1463 1487 1467
rect 1491 1466 1492 1467
rect 1499 1467 1505 1468
rect 1499 1466 1500 1467
rect 1491 1464 1500 1466
rect 1491 1463 1492 1464
rect 1486 1462 1492 1463
rect 1499 1463 1500 1464
rect 1504 1463 1505 1467
rect 1499 1462 1505 1463
rect 1611 1467 1617 1468
rect 1611 1463 1612 1467
rect 1616 1466 1617 1467
rect 1718 1467 1724 1468
rect 1718 1466 1719 1467
rect 1616 1464 1719 1466
rect 1616 1463 1617 1464
rect 1611 1462 1617 1463
rect 1718 1463 1719 1464
rect 1723 1463 1724 1467
rect 1718 1462 1724 1463
rect 1734 1467 1745 1468
rect 1734 1463 1735 1467
rect 1739 1463 1740 1467
rect 1744 1463 1745 1467
rect 1734 1462 1745 1463
rect 1871 1467 1877 1468
rect 1871 1463 1872 1467
rect 1876 1466 1877 1467
rect 1883 1467 1889 1468
rect 1883 1466 1884 1467
rect 1876 1464 1884 1466
rect 1876 1463 1877 1464
rect 1871 1462 1877 1463
rect 1883 1463 1884 1464
rect 1888 1463 1889 1467
rect 1883 1462 1889 1463
rect 2038 1467 2049 1468
rect 2038 1463 2039 1467
rect 2043 1463 2044 1467
rect 2048 1463 2049 1467
rect 2038 1462 2049 1463
rect 2211 1467 2217 1468
rect 2211 1463 2212 1467
rect 2216 1466 2217 1467
rect 2222 1467 2228 1468
rect 2222 1466 2223 1467
rect 2216 1464 2223 1466
rect 2216 1463 2217 1464
rect 2211 1462 2217 1463
rect 2222 1463 2223 1464
rect 2227 1463 2228 1467
rect 2222 1462 2228 1463
rect 2350 1467 2361 1468
rect 2350 1463 2351 1467
rect 2355 1463 2356 1467
rect 2360 1463 2361 1467
rect 2350 1462 2361 1463
rect 1371 1455 1377 1456
rect 1371 1451 1372 1455
rect 1376 1454 1377 1455
rect 1450 1455 1456 1456
rect 1450 1454 1451 1455
rect 1376 1452 1451 1454
rect 1376 1451 1377 1452
rect 1371 1450 1377 1451
rect 1450 1451 1451 1452
rect 1455 1451 1456 1455
rect 1450 1450 1456 1451
rect 1459 1455 1465 1456
rect 1459 1451 1460 1455
rect 1464 1454 1465 1455
rect 1494 1455 1500 1456
rect 1494 1454 1495 1455
rect 1464 1452 1495 1454
rect 1464 1451 1465 1452
rect 1459 1450 1465 1451
rect 1494 1451 1495 1452
rect 1499 1451 1500 1455
rect 1494 1450 1500 1451
rect 1547 1455 1553 1456
rect 1547 1451 1548 1455
rect 1552 1454 1553 1455
rect 1558 1455 1564 1456
rect 1558 1454 1559 1455
rect 1552 1452 1559 1454
rect 1552 1451 1553 1452
rect 1547 1450 1553 1451
rect 1558 1451 1559 1452
rect 1563 1451 1564 1455
rect 1558 1450 1564 1451
rect 1578 1455 1584 1456
rect 1578 1451 1579 1455
rect 1583 1454 1584 1455
rect 1635 1455 1641 1456
rect 1635 1454 1636 1455
rect 1583 1452 1636 1454
rect 1583 1451 1584 1452
rect 1578 1450 1584 1451
rect 1635 1451 1636 1452
rect 1640 1451 1641 1455
rect 1635 1450 1641 1451
rect 1666 1455 1672 1456
rect 1666 1451 1667 1455
rect 1671 1454 1672 1455
rect 1723 1455 1729 1456
rect 1723 1454 1724 1455
rect 1671 1452 1724 1454
rect 1671 1451 1672 1452
rect 1666 1450 1672 1451
rect 1723 1451 1724 1452
rect 1728 1451 1729 1455
rect 1723 1450 1729 1451
rect 1803 1455 1809 1456
rect 1803 1451 1804 1455
rect 1808 1454 1809 1455
rect 1826 1455 1832 1456
rect 1826 1454 1827 1455
rect 1808 1452 1827 1454
rect 1808 1451 1809 1452
rect 1803 1450 1809 1451
rect 1826 1451 1827 1452
rect 1831 1451 1832 1455
rect 1826 1450 1832 1451
rect 1834 1455 1840 1456
rect 1834 1451 1835 1455
rect 1839 1454 1840 1455
rect 1875 1455 1881 1456
rect 1875 1454 1876 1455
rect 1839 1452 1876 1454
rect 1839 1451 1840 1452
rect 1834 1450 1840 1451
rect 1875 1451 1876 1452
rect 1880 1451 1881 1455
rect 1875 1450 1881 1451
rect 1906 1455 1912 1456
rect 1906 1451 1907 1455
rect 1911 1454 1912 1455
rect 1939 1455 1945 1456
rect 1939 1454 1940 1455
rect 1911 1452 1940 1454
rect 1911 1451 1912 1452
rect 1906 1450 1912 1451
rect 1939 1451 1940 1452
rect 1944 1451 1945 1455
rect 1939 1450 1945 1451
rect 1995 1455 2001 1456
rect 1995 1451 1996 1455
rect 2000 1454 2001 1455
rect 2034 1455 2040 1456
rect 2034 1454 2035 1455
rect 2000 1452 2035 1454
rect 2000 1451 2001 1452
rect 1995 1450 2001 1451
rect 2034 1451 2035 1452
rect 2039 1451 2040 1455
rect 2034 1450 2040 1451
rect 2043 1455 2049 1456
rect 2043 1451 2044 1455
rect 2048 1454 2049 1455
rect 2082 1455 2088 1456
rect 2082 1454 2083 1455
rect 2048 1452 2083 1454
rect 2048 1451 2049 1452
rect 2043 1450 2049 1451
rect 2082 1451 2083 1452
rect 2087 1451 2088 1455
rect 2082 1450 2088 1451
rect 2091 1455 2097 1456
rect 2091 1451 2092 1455
rect 2096 1454 2097 1455
rect 2130 1455 2136 1456
rect 2130 1454 2131 1455
rect 2096 1452 2131 1454
rect 2096 1451 2097 1452
rect 2091 1450 2097 1451
rect 2130 1451 2131 1452
rect 2135 1451 2136 1455
rect 2130 1450 2136 1451
rect 2139 1455 2145 1456
rect 2139 1451 2140 1455
rect 2144 1454 2145 1455
rect 2178 1455 2184 1456
rect 2178 1454 2179 1455
rect 2144 1452 2179 1454
rect 2144 1451 2145 1452
rect 2139 1450 2145 1451
rect 2178 1451 2179 1452
rect 2183 1451 2184 1455
rect 2178 1450 2184 1451
rect 2187 1455 2193 1456
rect 2187 1451 2188 1455
rect 2192 1454 2193 1455
rect 2226 1455 2232 1456
rect 2226 1454 2227 1455
rect 2192 1452 2227 1454
rect 2192 1451 2193 1452
rect 2187 1450 2193 1451
rect 2226 1451 2227 1452
rect 2231 1451 2232 1455
rect 2226 1450 2232 1451
rect 2235 1455 2241 1456
rect 2235 1451 2236 1455
rect 2240 1454 2241 1455
rect 2266 1455 2272 1456
rect 2266 1454 2267 1455
rect 2240 1452 2267 1454
rect 2240 1451 2241 1452
rect 2235 1450 2241 1451
rect 2266 1451 2267 1452
rect 2271 1451 2272 1455
rect 2266 1450 2272 1451
rect 2275 1455 2281 1456
rect 2275 1451 2276 1455
rect 2280 1454 2281 1455
rect 2302 1455 2308 1456
rect 2302 1454 2303 1455
rect 2280 1452 2303 1454
rect 2280 1451 2281 1452
rect 2275 1450 2281 1451
rect 2302 1451 2303 1452
rect 2307 1451 2308 1455
rect 2302 1450 2308 1451
rect 2310 1455 2321 1456
rect 2310 1451 2311 1455
rect 2315 1451 2316 1455
rect 2320 1451 2321 1455
rect 2310 1450 2321 1451
rect 2355 1455 2361 1456
rect 2355 1451 2356 1455
rect 2360 1454 2361 1455
rect 2366 1455 2372 1456
rect 2366 1454 2367 1455
rect 2360 1452 2367 1454
rect 2360 1451 2361 1452
rect 2355 1450 2361 1451
rect 2366 1451 2367 1452
rect 2371 1451 2372 1455
rect 2366 1450 2372 1451
rect 139 1447 145 1448
rect 139 1443 140 1447
rect 144 1446 145 1447
rect 158 1447 164 1448
rect 158 1446 159 1447
rect 144 1444 159 1446
rect 144 1443 145 1444
rect 139 1442 145 1443
rect 158 1443 159 1444
rect 163 1443 164 1447
rect 158 1442 164 1443
rect 166 1447 172 1448
rect 166 1443 167 1447
rect 171 1446 172 1447
rect 179 1447 185 1448
rect 179 1446 180 1447
rect 171 1444 180 1446
rect 171 1443 172 1444
rect 166 1442 172 1443
rect 179 1443 180 1444
rect 184 1443 185 1447
rect 179 1442 185 1443
rect 206 1447 212 1448
rect 206 1443 207 1447
rect 211 1446 212 1447
rect 219 1447 225 1448
rect 219 1446 220 1447
rect 211 1444 220 1446
rect 211 1443 212 1444
rect 206 1442 212 1443
rect 219 1443 220 1444
rect 224 1443 225 1447
rect 219 1442 225 1443
rect 250 1447 256 1448
rect 250 1443 251 1447
rect 255 1446 256 1447
rect 259 1447 265 1448
rect 259 1446 260 1447
rect 255 1444 260 1446
rect 255 1443 256 1444
rect 250 1442 256 1443
rect 259 1443 260 1444
rect 264 1443 265 1447
rect 259 1442 265 1443
rect 303 1447 309 1448
rect 303 1443 304 1447
rect 308 1446 309 1447
rect 315 1447 321 1448
rect 315 1446 316 1447
rect 308 1444 316 1446
rect 308 1443 309 1444
rect 303 1442 309 1443
rect 315 1443 316 1444
rect 320 1443 321 1447
rect 315 1442 321 1443
rect 346 1447 352 1448
rect 346 1443 347 1447
rect 351 1446 352 1447
rect 387 1447 393 1448
rect 387 1446 388 1447
rect 351 1444 388 1446
rect 351 1443 352 1444
rect 346 1442 352 1443
rect 387 1443 388 1444
rect 392 1443 393 1447
rect 387 1442 393 1443
rect 418 1447 424 1448
rect 418 1443 419 1447
rect 423 1446 424 1447
rect 467 1447 473 1448
rect 467 1446 468 1447
rect 423 1444 468 1446
rect 423 1443 424 1444
rect 418 1442 424 1443
rect 467 1443 468 1444
rect 472 1443 473 1447
rect 467 1442 473 1443
rect 498 1447 504 1448
rect 498 1443 499 1447
rect 503 1446 504 1447
rect 555 1447 561 1448
rect 555 1446 556 1447
rect 503 1444 556 1446
rect 503 1443 504 1444
rect 498 1442 504 1443
rect 555 1443 556 1444
rect 560 1443 561 1447
rect 555 1442 561 1443
rect 586 1447 592 1448
rect 586 1443 587 1447
rect 591 1446 592 1447
rect 643 1447 649 1448
rect 643 1446 644 1447
rect 591 1444 644 1446
rect 591 1443 592 1444
rect 586 1442 592 1443
rect 643 1443 644 1444
rect 648 1443 649 1447
rect 643 1442 649 1443
rect 723 1447 729 1448
rect 723 1443 724 1447
rect 728 1446 729 1447
rect 742 1447 748 1448
rect 742 1446 743 1447
rect 728 1444 743 1446
rect 728 1443 729 1444
rect 723 1442 729 1443
rect 742 1443 743 1444
rect 747 1443 748 1447
rect 742 1442 748 1443
rect 754 1447 760 1448
rect 754 1443 755 1447
rect 759 1446 760 1447
rect 803 1447 809 1448
rect 803 1446 804 1447
rect 759 1444 804 1446
rect 759 1443 760 1444
rect 754 1442 760 1443
rect 803 1443 804 1444
rect 808 1443 809 1447
rect 803 1442 809 1443
rect 834 1447 840 1448
rect 834 1443 835 1447
rect 839 1446 840 1447
rect 875 1447 881 1448
rect 875 1446 876 1447
rect 839 1444 876 1446
rect 839 1443 840 1444
rect 834 1442 840 1443
rect 875 1443 876 1444
rect 880 1443 881 1447
rect 875 1442 881 1443
rect 906 1447 912 1448
rect 906 1443 907 1447
rect 911 1446 912 1447
rect 939 1447 945 1448
rect 939 1446 940 1447
rect 911 1444 940 1446
rect 911 1443 912 1444
rect 906 1442 912 1443
rect 939 1443 940 1444
rect 944 1443 945 1447
rect 939 1442 945 1443
rect 970 1447 976 1448
rect 970 1443 971 1447
rect 975 1446 976 1447
rect 995 1447 1001 1448
rect 995 1446 996 1447
rect 975 1444 996 1446
rect 975 1443 976 1444
rect 970 1442 976 1443
rect 995 1443 996 1444
rect 1000 1443 1001 1447
rect 995 1442 1001 1443
rect 1026 1447 1032 1448
rect 1026 1443 1027 1447
rect 1031 1446 1032 1447
rect 1043 1447 1049 1448
rect 1043 1446 1044 1447
rect 1031 1444 1044 1446
rect 1031 1443 1032 1444
rect 1026 1442 1032 1443
rect 1043 1443 1044 1444
rect 1048 1443 1049 1447
rect 1043 1442 1049 1443
rect 1074 1447 1080 1448
rect 1074 1443 1075 1447
rect 1079 1446 1080 1447
rect 1099 1447 1105 1448
rect 1099 1446 1100 1447
rect 1079 1444 1100 1446
rect 1079 1443 1080 1444
rect 1074 1442 1080 1443
rect 1099 1443 1100 1444
rect 1104 1443 1105 1447
rect 1099 1442 1105 1443
rect 1138 1447 1144 1448
rect 1138 1443 1139 1447
rect 1143 1446 1144 1447
rect 1147 1447 1153 1448
rect 1147 1446 1148 1447
rect 1143 1444 1148 1446
rect 1143 1443 1144 1444
rect 1138 1442 1144 1443
rect 1147 1443 1148 1444
rect 1152 1443 1153 1447
rect 1147 1442 1153 1443
rect 1174 1447 1180 1448
rect 1174 1443 1175 1447
rect 1179 1446 1180 1447
rect 1187 1447 1193 1448
rect 1187 1446 1188 1447
rect 1179 1444 1188 1446
rect 1179 1443 1180 1444
rect 1174 1442 1180 1443
rect 1187 1443 1188 1444
rect 1192 1443 1193 1447
rect 1187 1442 1193 1443
rect 1374 1447 1380 1448
rect 1374 1443 1375 1447
rect 1379 1443 1380 1447
rect 1374 1442 1380 1443
rect 1462 1447 1468 1448
rect 1462 1443 1463 1447
rect 1467 1443 1468 1447
rect 1462 1442 1468 1443
rect 1550 1447 1556 1448
rect 1550 1443 1551 1447
rect 1555 1443 1556 1447
rect 1550 1442 1556 1443
rect 1638 1447 1644 1448
rect 1638 1443 1639 1447
rect 1643 1443 1644 1447
rect 1638 1442 1644 1443
rect 1726 1447 1732 1448
rect 1726 1443 1727 1447
rect 1731 1443 1732 1447
rect 1726 1442 1732 1443
rect 1806 1447 1812 1448
rect 1806 1443 1807 1447
rect 1811 1443 1812 1447
rect 1806 1442 1812 1443
rect 1878 1447 1884 1448
rect 1878 1443 1879 1447
rect 1883 1443 1884 1447
rect 1878 1442 1884 1443
rect 1942 1447 1948 1448
rect 1942 1443 1943 1447
rect 1947 1443 1948 1447
rect 1942 1442 1948 1443
rect 1998 1447 2004 1448
rect 1998 1443 1999 1447
rect 2003 1443 2004 1447
rect 1998 1442 2004 1443
rect 2046 1447 2052 1448
rect 2046 1443 2047 1447
rect 2051 1443 2052 1447
rect 2046 1442 2052 1443
rect 2094 1447 2100 1448
rect 2094 1443 2095 1447
rect 2099 1443 2100 1447
rect 2094 1442 2100 1443
rect 2142 1447 2148 1448
rect 2142 1443 2143 1447
rect 2147 1443 2148 1447
rect 2142 1442 2148 1443
rect 2190 1447 2196 1448
rect 2190 1443 2191 1447
rect 2195 1443 2196 1447
rect 2190 1442 2196 1443
rect 2238 1447 2244 1448
rect 2238 1443 2239 1447
rect 2243 1443 2244 1447
rect 2238 1442 2244 1443
rect 2278 1447 2284 1448
rect 2278 1443 2279 1447
rect 2283 1443 2284 1447
rect 2278 1442 2284 1443
rect 2318 1447 2324 1448
rect 2318 1443 2319 1447
rect 2323 1443 2324 1447
rect 2318 1442 2324 1443
rect 2358 1447 2364 1448
rect 2358 1443 2359 1447
rect 2363 1443 2364 1447
rect 2358 1442 2364 1443
rect 142 1439 148 1440
rect 142 1435 143 1439
rect 147 1435 148 1439
rect 142 1434 148 1435
rect 182 1439 188 1440
rect 182 1435 183 1439
rect 187 1435 188 1439
rect 182 1434 188 1435
rect 222 1439 228 1440
rect 222 1435 223 1439
rect 227 1435 228 1439
rect 222 1434 228 1435
rect 262 1439 268 1440
rect 262 1435 263 1439
rect 267 1435 268 1439
rect 262 1434 268 1435
rect 318 1439 324 1440
rect 318 1435 319 1439
rect 323 1435 324 1439
rect 318 1434 324 1435
rect 390 1439 396 1440
rect 390 1435 391 1439
rect 395 1435 396 1439
rect 390 1434 396 1435
rect 470 1439 476 1440
rect 470 1435 471 1439
rect 475 1435 476 1439
rect 470 1434 476 1435
rect 558 1439 564 1440
rect 558 1435 559 1439
rect 563 1435 564 1439
rect 558 1434 564 1435
rect 646 1439 652 1440
rect 646 1435 647 1439
rect 651 1435 652 1439
rect 646 1434 652 1435
rect 726 1439 732 1440
rect 726 1435 727 1439
rect 731 1435 732 1439
rect 726 1434 732 1435
rect 806 1439 812 1440
rect 806 1435 807 1439
rect 811 1435 812 1439
rect 806 1434 812 1435
rect 878 1439 884 1440
rect 878 1435 879 1439
rect 883 1435 884 1439
rect 878 1434 884 1435
rect 942 1439 948 1440
rect 942 1435 943 1439
rect 947 1435 948 1439
rect 942 1434 948 1435
rect 998 1439 1004 1440
rect 998 1435 999 1439
rect 1003 1435 1004 1439
rect 998 1434 1004 1435
rect 1046 1439 1052 1440
rect 1046 1435 1047 1439
rect 1051 1435 1052 1439
rect 1046 1434 1052 1435
rect 1102 1439 1108 1440
rect 1102 1435 1103 1439
rect 1107 1435 1108 1439
rect 1102 1434 1108 1435
rect 1150 1439 1156 1440
rect 1150 1435 1151 1439
rect 1155 1435 1156 1439
rect 1150 1434 1156 1435
rect 1190 1439 1196 1440
rect 1190 1435 1191 1439
rect 1195 1435 1196 1439
rect 1190 1434 1196 1435
rect 1826 1427 1832 1428
rect 1278 1424 1284 1425
rect 1278 1420 1279 1424
rect 1283 1420 1284 1424
rect 1826 1423 1827 1427
rect 1831 1426 1832 1427
rect 2266 1427 2272 1428
rect 1831 1424 2001 1426
rect 1831 1423 1832 1424
rect 1826 1422 1832 1423
rect 1999 1422 2001 1424
rect 2266 1423 2267 1427
rect 2271 1426 2272 1427
rect 2302 1427 2308 1428
rect 2271 1423 2274 1426
rect 2266 1422 2274 1423
rect 2302 1423 2303 1427
rect 2307 1426 2308 1427
rect 2307 1424 2314 1426
rect 2307 1423 2308 1424
rect 2302 1422 2308 1423
rect 1999 1420 2014 1422
rect 1278 1419 1284 1420
rect 1350 1419 1356 1420
rect 110 1416 116 1417
rect 110 1412 111 1416
rect 115 1412 116 1416
rect 1238 1416 1244 1417
rect 1238 1412 1239 1416
rect 1243 1412 1244 1416
rect 1350 1415 1351 1419
rect 1355 1418 1356 1419
rect 1399 1419 1405 1420
rect 1399 1418 1400 1419
rect 1355 1416 1400 1418
rect 1355 1415 1356 1416
rect 1350 1414 1356 1415
rect 1399 1415 1400 1416
rect 1404 1415 1405 1419
rect 1399 1414 1405 1415
rect 1450 1419 1456 1420
rect 1450 1415 1451 1419
rect 1455 1418 1456 1419
rect 1487 1419 1493 1420
rect 1487 1418 1488 1419
rect 1455 1416 1488 1418
rect 1455 1415 1456 1416
rect 1450 1414 1456 1415
rect 1487 1415 1488 1416
rect 1492 1415 1493 1419
rect 1487 1414 1493 1415
rect 1575 1419 1584 1420
rect 1575 1415 1576 1419
rect 1583 1415 1584 1419
rect 1575 1414 1584 1415
rect 1663 1419 1672 1420
rect 1663 1415 1664 1419
rect 1671 1415 1672 1419
rect 1663 1414 1672 1415
rect 1718 1419 1724 1420
rect 1718 1415 1719 1419
rect 1723 1418 1724 1419
rect 1751 1419 1757 1420
rect 1751 1418 1752 1419
rect 1723 1416 1752 1418
rect 1723 1415 1724 1416
rect 1718 1414 1724 1415
rect 1751 1415 1752 1416
rect 1756 1415 1757 1419
rect 1751 1414 1757 1415
rect 1831 1419 1840 1420
rect 1831 1415 1832 1419
rect 1839 1415 1840 1419
rect 1831 1414 1840 1415
rect 1903 1419 1912 1420
rect 1903 1415 1904 1419
rect 1911 1415 1912 1419
rect 1903 1414 1912 1415
rect 1967 1419 1973 1420
rect 1967 1415 1968 1419
rect 1972 1418 1973 1419
rect 2012 1418 2014 1420
rect 2023 1419 2029 1420
rect 2023 1418 2024 1419
rect 1972 1416 2001 1418
rect 2012 1416 2024 1418
rect 1972 1415 1973 1416
rect 1967 1414 1973 1415
rect 110 1411 116 1412
rect 166 1411 173 1412
rect 166 1407 167 1411
rect 172 1407 173 1411
rect 166 1406 173 1407
rect 206 1411 213 1412
rect 206 1407 207 1411
rect 212 1407 213 1411
rect 206 1406 213 1407
rect 247 1411 256 1412
rect 247 1407 248 1411
rect 255 1407 256 1411
rect 247 1406 256 1407
rect 287 1411 293 1412
rect 287 1407 288 1411
rect 292 1410 293 1411
rect 303 1411 309 1412
rect 303 1410 304 1411
rect 292 1408 304 1410
rect 292 1407 293 1408
rect 287 1406 293 1407
rect 303 1407 304 1408
rect 308 1407 309 1411
rect 303 1406 309 1407
rect 343 1411 352 1412
rect 343 1407 344 1411
rect 351 1407 352 1411
rect 343 1406 352 1407
rect 415 1411 424 1412
rect 415 1407 416 1411
rect 423 1407 424 1411
rect 415 1406 424 1407
rect 495 1411 504 1412
rect 495 1407 496 1411
rect 503 1407 504 1411
rect 495 1406 504 1407
rect 583 1411 592 1412
rect 583 1407 584 1411
rect 591 1407 592 1411
rect 671 1411 677 1412
rect 671 1410 672 1411
rect 583 1406 592 1407
rect 596 1408 672 1410
rect 374 1403 380 1404
rect 110 1399 116 1400
rect 110 1395 111 1399
rect 115 1395 116 1399
rect 374 1399 375 1403
rect 379 1402 380 1403
rect 596 1402 598 1408
rect 671 1407 672 1408
rect 676 1407 677 1411
rect 671 1406 677 1407
rect 751 1411 760 1412
rect 751 1407 752 1411
rect 759 1407 760 1411
rect 751 1406 760 1407
rect 831 1411 840 1412
rect 831 1407 832 1411
rect 839 1407 840 1411
rect 831 1406 840 1407
rect 903 1411 912 1412
rect 903 1407 904 1411
rect 911 1407 912 1411
rect 903 1406 912 1407
rect 967 1411 976 1412
rect 967 1407 968 1411
rect 975 1407 976 1411
rect 967 1406 976 1407
rect 1023 1411 1032 1412
rect 1023 1407 1024 1411
rect 1031 1407 1032 1411
rect 1023 1406 1032 1407
rect 1071 1411 1080 1412
rect 1071 1407 1072 1411
rect 1079 1407 1080 1411
rect 1071 1406 1080 1407
rect 1127 1411 1133 1412
rect 1127 1407 1128 1411
rect 1132 1410 1133 1411
rect 1138 1411 1144 1412
rect 1138 1410 1139 1411
rect 1132 1408 1139 1410
rect 1132 1407 1133 1408
rect 1127 1406 1133 1407
rect 1138 1407 1139 1408
rect 1143 1407 1144 1411
rect 1138 1406 1144 1407
rect 1174 1411 1181 1412
rect 1174 1407 1175 1411
rect 1180 1407 1181 1411
rect 1215 1411 1221 1412
rect 1238 1411 1244 1412
rect 1215 1410 1216 1411
rect 1174 1406 1181 1407
rect 1188 1408 1216 1410
rect 379 1400 598 1402
rect 1086 1403 1092 1404
rect 379 1399 380 1400
rect 374 1398 380 1399
rect 1086 1399 1087 1403
rect 1091 1402 1092 1403
rect 1188 1402 1190 1408
rect 1215 1407 1216 1408
rect 1220 1407 1221 1411
rect 1999 1410 2001 1416
rect 2023 1415 2024 1416
rect 2028 1415 2029 1419
rect 2023 1414 2029 1415
rect 2034 1419 2040 1420
rect 2034 1415 2035 1419
rect 2039 1418 2040 1419
rect 2071 1419 2077 1420
rect 2071 1418 2072 1419
rect 2039 1416 2072 1418
rect 2039 1415 2040 1416
rect 2034 1414 2040 1415
rect 2071 1415 2072 1416
rect 2076 1415 2077 1419
rect 2071 1414 2077 1415
rect 2082 1419 2088 1420
rect 2082 1415 2083 1419
rect 2087 1418 2088 1419
rect 2119 1419 2125 1420
rect 2119 1418 2120 1419
rect 2087 1416 2120 1418
rect 2087 1415 2088 1416
rect 2082 1414 2088 1415
rect 2119 1415 2120 1416
rect 2124 1415 2125 1419
rect 2119 1414 2125 1415
rect 2130 1419 2136 1420
rect 2130 1415 2131 1419
rect 2135 1418 2136 1419
rect 2167 1419 2173 1420
rect 2167 1418 2168 1419
rect 2135 1416 2168 1418
rect 2135 1415 2136 1416
rect 2130 1414 2136 1415
rect 2167 1415 2168 1416
rect 2172 1415 2173 1419
rect 2167 1414 2173 1415
rect 2178 1419 2184 1420
rect 2178 1415 2179 1419
rect 2183 1418 2184 1419
rect 2215 1419 2221 1420
rect 2215 1418 2216 1419
rect 2183 1416 2216 1418
rect 2183 1415 2184 1416
rect 2178 1414 2184 1415
rect 2215 1415 2216 1416
rect 2220 1415 2221 1419
rect 2215 1414 2221 1415
rect 2226 1419 2232 1420
rect 2226 1415 2227 1419
rect 2231 1418 2232 1419
rect 2263 1419 2269 1420
rect 2263 1418 2264 1419
rect 2231 1416 2264 1418
rect 2231 1415 2232 1416
rect 2226 1414 2232 1415
rect 2263 1415 2264 1416
rect 2268 1415 2269 1419
rect 2272 1418 2274 1422
rect 2303 1419 2309 1420
rect 2303 1418 2304 1419
rect 2272 1416 2304 1418
rect 2263 1414 2269 1415
rect 2303 1415 2304 1416
rect 2308 1415 2309 1419
rect 2312 1418 2314 1424
rect 2406 1424 2412 1425
rect 2406 1420 2407 1424
rect 2411 1420 2412 1424
rect 2343 1419 2349 1420
rect 2343 1418 2344 1419
rect 2312 1416 2344 1418
rect 2303 1414 2309 1415
rect 2343 1415 2344 1416
rect 2348 1415 2349 1419
rect 2343 1414 2349 1415
rect 2374 1419 2380 1420
rect 2374 1415 2375 1419
rect 2379 1418 2380 1419
rect 2383 1419 2389 1420
rect 2406 1419 2412 1420
rect 2383 1418 2384 1419
rect 2379 1416 2384 1418
rect 2379 1415 2380 1416
rect 2374 1414 2380 1415
rect 2383 1415 2384 1416
rect 2388 1415 2389 1419
rect 2383 1414 2389 1415
rect 2014 1411 2020 1412
rect 2014 1410 2015 1411
rect 1999 1408 2015 1410
rect 1215 1406 1221 1407
rect 1278 1407 1284 1408
rect 1278 1403 1279 1407
rect 1283 1403 1284 1407
rect 2014 1407 2015 1408
rect 2019 1407 2020 1411
rect 2014 1406 2020 1407
rect 2406 1407 2412 1408
rect 1278 1402 1284 1403
rect 2406 1403 2407 1407
rect 2411 1403 2412 1407
rect 2406 1402 2412 1403
rect 1091 1400 1190 1402
rect 1374 1400 1380 1401
rect 1091 1399 1092 1400
rect 1086 1398 1092 1399
rect 1238 1399 1244 1400
rect 110 1394 116 1395
rect 1238 1395 1239 1399
rect 1243 1395 1244 1399
rect 1374 1396 1375 1400
rect 1379 1396 1380 1400
rect 1374 1395 1380 1396
rect 1462 1400 1468 1401
rect 1462 1396 1463 1400
rect 1467 1396 1468 1400
rect 1462 1395 1468 1396
rect 1550 1400 1556 1401
rect 1550 1396 1551 1400
rect 1555 1396 1556 1400
rect 1550 1395 1556 1396
rect 1638 1400 1644 1401
rect 1638 1396 1639 1400
rect 1643 1396 1644 1400
rect 1638 1395 1644 1396
rect 1726 1400 1732 1401
rect 1726 1396 1727 1400
rect 1731 1396 1732 1400
rect 1726 1395 1732 1396
rect 1806 1400 1812 1401
rect 1806 1396 1807 1400
rect 1811 1396 1812 1400
rect 1806 1395 1812 1396
rect 1878 1400 1884 1401
rect 1878 1396 1879 1400
rect 1883 1396 1884 1400
rect 1878 1395 1884 1396
rect 1942 1400 1948 1401
rect 1942 1396 1943 1400
rect 1947 1396 1948 1400
rect 1942 1395 1948 1396
rect 1998 1400 2004 1401
rect 1998 1396 1999 1400
rect 2003 1396 2004 1400
rect 1998 1395 2004 1396
rect 2046 1400 2052 1401
rect 2046 1396 2047 1400
rect 2051 1396 2052 1400
rect 2046 1395 2052 1396
rect 2094 1400 2100 1401
rect 2094 1396 2095 1400
rect 2099 1396 2100 1400
rect 2094 1395 2100 1396
rect 2142 1400 2148 1401
rect 2142 1396 2143 1400
rect 2147 1396 2148 1400
rect 2142 1395 2148 1396
rect 2190 1400 2196 1401
rect 2190 1396 2191 1400
rect 2195 1396 2196 1400
rect 2190 1395 2196 1396
rect 2238 1400 2244 1401
rect 2238 1396 2239 1400
rect 2243 1396 2244 1400
rect 2238 1395 2244 1396
rect 2278 1400 2284 1401
rect 2278 1396 2279 1400
rect 2283 1396 2284 1400
rect 2278 1395 2284 1396
rect 2318 1400 2324 1401
rect 2318 1396 2319 1400
rect 2323 1396 2324 1400
rect 2318 1395 2324 1396
rect 2358 1400 2364 1401
rect 2358 1396 2359 1400
rect 2363 1396 2364 1400
rect 2358 1395 2364 1396
rect 1238 1394 1244 1395
rect 142 1392 148 1393
rect 142 1388 143 1392
rect 147 1388 148 1392
rect 142 1387 148 1388
rect 182 1392 188 1393
rect 182 1388 183 1392
rect 187 1388 188 1392
rect 182 1387 188 1388
rect 222 1392 228 1393
rect 222 1388 223 1392
rect 227 1388 228 1392
rect 222 1387 228 1388
rect 262 1392 268 1393
rect 262 1388 263 1392
rect 267 1388 268 1392
rect 262 1387 268 1388
rect 318 1392 324 1393
rect 318 1388 319 1392
rect 323 1388 324 1392
rect 318 1387 324 1388
rect 390 1392 396 1393
rect 390 1388 391 1392
rect 395 1388 396 1392
rect 390 1387 396 1388
rect 470 1392 476 1393
rect 470 1388 471 1392
rect 475 1388 476 1392
rect 470 1387 476 1388
rect 558 1392 564 1393
rect 558 1388 559 1392
rect 563 1388 564 1392
rect 558 1387 564 1388
rect 646 1392 652 1393
rect 646 1388 647 1392
rect 651 1388 652 1392
rect 646 1387 652 1388
rect 726 1392 732 1393
rect 726 1388 727 1392
rect 731 1388 732 1392
rect 726 1387 732 1388
rect 806 1392 812 1393
rect 806 1388 807 1392
rect 811 1388 812 1392
rect 806 1387 812 1388
rect 878 1392 884 1393
rect 878 1388 879 1392
rect 883 1388 884 1392
rect 878 1387 884 1388
rect 942 1392 948 1393
rect 942 1388 943 1392
rect 947 1388 948 1392
rect 942 1387 948 1388
rect 998 1392 1004 1393
rect 998 1388 999 1392
rect 1003 1388 1004 1392
rect 998 1387 1004 1388
rect 1046 1392 1052 1393
rect 1046 1388 1047 1392
rect 1051 1388 1052 1392
rect 1046 1387 1052 1388
rect 1102 1392 1108 1393
rect 1102 1388 1103 1392
rect 1107 1388 1108 1392
rect 1102 1387 1108 1388
rect 1150 1392 1156 1393
rect 1150 1388 1151 1392
rect 1155 1388 1156 1392
rect 1150 1387 1156 1388
rect 1190 1392 1196 1393
rect 1190 1388 1191 1392
rect 1195 1388 1196 1392
rect 1190 1387 1196 1388
rect 166 1380 172 1381
rect 166 1376 167 1380
rect 171 1376 172 1380
rect 166 1375 172 1376
rect 206 1380 212 1381
rect 206 1376 207 1380
rect 211 1376 212 1380
rect 206 1375 212 1376
rect 246 1380 252 1381
rect 246 1376 247 1380
rect 251 1376 252 1380
rect 246 1375 252 1376
rect 302 1380 308 1381
rect 302 1376 303 1380
rect 307 1376 308 1380
rect 302 1375 308 1376
rect 366 1380 372 1381
rect 366 1376 367 1380
rect 371 1376 372 1380
rect 366 1375 372 1376
rect 438 1380 444 1381
rect 438 1376 439 1380
rect 443 1376 444 1380
rect 438 1375 444 1376
rect 518 1380 524 1381
rect 518 1376 519 1380
rect 523 1376 524 1380
rect 518 1375 524 1376
rect 598 1380 604 1381
rect 598 1376 599 1380
rect 603 1376 604 1380
rect 598 1375 604 1376
rect 678 1380 684 1381
rect 678 1376 679 1380
rect 683 1376 684 1380
rect 678 1375 684 1376
rect 750 1380 756 1381
rect 750 1376 751 1380
rect 755 1376 756 1380
rect 750 1375 756 1376
rect 822 1380 828 1381
rect 822 1376 823 1380
rect 827 1376 828 1380
rect 822 1375 828 1376
rect 886 1380 892 1381
rect 886 1376 887 1380
rect 891 1376 892 1380
rect 886 1375 892 1376
rect 950 1380 956 1381
rect 950 1376 951 1380
rect 955 1376 956 1380
rect 950 1375 956 1376
rect 1014 1380 1020 1381
rect 1014 1376 1015 1380
rect 1019 1376 1020 1380
rect 1014 1375 1020 1376
rect 1078 1380 1084 1381
rect 1078 1376 1079 1380
rect 1083 1376 1084 1380
rect 1078 1375 1084 1376
rect 1142 1380 1148 1381
rect 1142 1376 1143 1380
rect 1147 1376 1148 1380
rect 1142 1375 1148 1376
rect 1190 1380 1196 1381
rect 1190 1376 1191 1380
rect 1195 1376 1196 1380
rect 1190 1375 1196 1376
rect 1302 1380 1308 1381
rect 1302 1376 1303 1380
rect 1307 1376 1308 1380
rect 1302 1375 1308 1376
rect 1342 1380 1348 1381
rect 1342 1376 1343 1380
rect 1347 1376 1348 1380
rect 1342 1375 1348 1376
rect 1398 1380 1404 1381
rect 1398 1376 1399 1380
rect 1403 1376 1404 1380
rect 1398 1375 1404 1376
rect 1462 1380 1468 1381
rect 1462 1376 1463 1380
rect 1467 1376 1468 1380
rect 1462 1375 1468 1376
rect 1534 1380 1540 1381
rect 1534 1376 1535 1380
rect 1539 1376 1540 1380
rect 1534 1375 1540 1376
rect 1606 1380 1612 1381
rect 1606 1376 1607 1380
rect 1611 1376 1612 1380
rect 1606 1375 1612 1376
rect 1686 1380 1692 1381
rect 1686 1376 1687 1380
rect 1691 1376 1692 1380
rect 1686 1375 1692 1376
rect 1766 1380 1772 1381
rect 1766 1376 1767 1380
rect 1771 1376 1772 1380
rect 1766 1375 1772 1376
rect 1846 1380 1852 1381
rect 1846 1376 1847 1380
rect 1851 1376 1852 1380
rect 1846 1375 1852 1376
rect 1934 1380 1940 1381
rect 1934 1376 1935 1380
rect 1939 1376 1940 1380
rect 1934 1375 1940 1376
rect 2022 1380 2028 1381
rect 2022 1376 2023 1380
rect 2027 1376 2028 1380
rect 2022 1375 2028 1376
rect 2110 1380 2116 1381
rect 2110 1376 2111 1380
rect 2115 1376 2116 1380
rect 2110 1375 2116 1376
rect 2198 1380 2204 1381
rect 2198 1376 2199 1380
rect 2203 1376 2204 1380
rect 2198 1375 2204 1376
rect 2286 1380 2292 1381
rect 2286 1376 2287 1380
rect 2291 1376 2292 1380
rect 2286 1375 2292 1376
rect 2358 1380 2364 1381
rect 2358 1376 2359 1380
rect 2363 1376 2364 1380
rect 2358 1375 2364 1376
rect 110 1373 116 1374
rect 110 1369 111 1373
rect 115 1369 116 1373
rect 110 1368 116 1369
rect 1238 1373 1244 1374
rect 1238 1369 1239 1373
rect 1243 1369 1244 1373
rect 1238 1368 1244 1369
rect 1278 1373 1284 1374
rect 1278 1369 1279 1373
rect 1283 1369 1284 1373
rect 1278 1368 1284 1369
rect 2406 1373 2412 1374
rect 2406 1369 2407 1373
rect 2411 1369 2412 1373
rect 2406 1368 2412 1369
rect 158 1367 164 1368
rect 158 1363 159 1367
rect 163 1366 164 1367
rect 742 1367 748 1368
rect 163 1364 321 1366
rect 163 1363 164 1364
rect 158 1362 164 1363
rect 191 1359 200 1360
rect 110 1356 116 1357
rect 110 1352 111 1356
rect 115 1352 116 1356
rect 191 1355 192 1359
rect 199 1355 200 1359
rect 191 1354 200 1355
rect 231 1359 240 1360
rect 231 1355 232 1359
rect 239 1355 240 1359
rect 231 1354 240 1355
rect 271 1359 277 1360
rect 271 1355 272 1359
rect 276 1358 277 1359
rect 294 1359 300 1360
rect 294 1358 295 1359
rect 276 1356 295 1358
rect 276 1355 277 1356
rect 271 1354 277 1355
rect 294 1355 295 1356
rect 299 1355 300 1359
rect 319 1358 321 1364
rect 742 1363 743 1367
rect 747 1366 748 1367
rect 747 1364 1018 1366
rect 747 1363 748 1364
rect 742 1362 748 1363
rect 327 1359 333 1360
rect 327 1358 328 1359
rect 319 1356 328 1358
rect 294 1354 300 1355
rect 327 1355 328 1356
rect 332 1355 333 1359
rect 327 1354 333 1355
rect 391 1359 397 1360
rect 391 1355 392 1359
rect 396 1358 397 1359
rect 430 1359 436 1360
rect 430 1358 431 1359
rect 396 1356 431 1358
rect 396 1355 397 1356
rect 391 1354 397 1355
rect 430 1355 431 1356
rect 435 1355 436 1359
rect 430 1354 436 1355
rect 463 1359 469 1360
rect 463 1355 464 1359
rect 468 1358 469 1359
rect 510 1359 516 1360
rect 510 1358 511 1359
rect 468 1356 511 1358
rect 468 1355 469 1356
rect 463 1354 469 1355
rect 510 1355 511 1356
rect 515 1355 516 1359
rect 510 1354 516 1355
rect 543 1359 549 1360
rect 543 1355 544 1359
rect 548 1358 549 1359
rect 590 1359 596 1360
rect 590 1358 591 1359
rect 548 1356 591 1358
rect 548 1355 549 1356
rect 543 1354 549 1355
rect 590 1355 591 1356
rect 595 1355 596 1359
rect 590 1354 596 1355
rect 606 1359 612 1360
rect 606 1355 607 1359
rect 611 1358 612 1359
rect 623 1359 629 1360
rect 623 1358 624 1359
rect 611 1356 624 1358
rect 611 1355 612 1356
rect 606 1354 612 1355
rect 623 1355 624 1356
rect 628 1355 629 1359
rect 623 1354 629 1355
rect 703 1359 709 1360
rect 703 1355 704 1359
rect 708 1358 709 1359
rect 742 1359 748 1360
rect 742 1358 743 1359
rect 708 1356 743 1358
rect 708 1355 709 1356
rect 703 1354 709 1355
rect 742 1355 743 1356
rect 747 1355 748 1359
rect 742 1354 748 1355
rect 775 1359 781 1360
rect 775 1355 776 1359
rect 780 1358 781 1359
rect 814 1359 820 1360
rect 814 1358 815 1359
rect 780 1356 815 1358
rect 780 1355 781 1356
rect 775 1354 781 1355
rect 814 1355 815 1356
rect 819 1355 820 1359
rect 814 1354 820 1355
rect 847 1359 853 1360
rect 847 1355 848 1359
rect 852 1358 853 1359
rect 878 1359 884 1360
rect 878 1358 879 1359
rect 852 1356 879 1358
rect 852 1355 853 1356
rect 847 1354 853 1355
rect 878 1355 879 1356
rect 883 1355 884 1359
rect 878 1354 884 1355
rect 911 1359 917 1360
rect 911 1355 912 1359
rect 916 1358 917 1359
rect 942 1359 948 1360
rect 942 1358 943 1359
rect 916 1356 943 1358
rect 916 1355 917 1356
rect 911 1354 917 1355
rect 942 1355 943 1356
rect 947 1355 948 1359
rect 942 1354 948 1355
rect 975 1359 981 1360
rect 975 1355 976 1359
rect 980 1358 981 1359
rect 1006 1359 1012 1360
rect 1006 1358 1007 1359
rect 980 1356 1007 1358
rect 980 1355 981 1356
rect 975 1354 981 1355
rect 1006 1355 1007 1356
rect 1011 1355 1012 1359
rect 1016 1358 1018 1364
rect 1039 1359 1045 1360
rect 1039 1358 1040 1359
rect 1016 1356 1040 1358
rect 1006 1354 1012 1355
rect 1039 1355 1040 1356
rect 1044 1355 1045 1359
rect 1039 1354 1045 1355
rect 1103 1359 1109 1360
rect 1103 1355 1104 1359
rect 1108 1358 1109 1359
rect 1134 1359 1140 1360
rect 1134 1358 1135 1359
rect 1108 1356 1135 1358
rect 1108 1355 1109 1356
rect 1103 1354 1109 1355
rect 1134 1355 1135 1356
rect 1139 1355 1140 1359
rect 1134 1354 1140 1355
rect 1167 1359 1173 1360
rect 1167 1355 1168 1359
rect 1172 1358 1173 1359
rect 1182 1359 1188 1360
rect 1182 1358 1183 1359
rect 1172 1356 1183 1358
rect 1172 1355 1173 1356
rect 1167 1354 1173 1355
rect 1182 1355 1183 1356
rect 1187 1355 1188 1359
rect 1182 1354 1188 1355
rect 1215 1359 1221 1360
rect 1215 1355 1216 1359
rect 1220 1358 1221 1359
rect 1230 1359 1236 1360
rect 1230 1358 1231 1359
rect 1220 1356 1231 1358
rect 1220 1355 1221 1356
rect 1215 1354 1221 1355
rect 1230 1355 1231 1356
rect 1235 1355 1236 1359
rect 1310 1359 1316 1360
rect 1230 1354 1236 1355
rect 1238 1356 1244 1357
rect 110 1351 116 1352
rect 1238 1352 1239 1356
rect 1243 1352 1244 1356
rect 1238 1351 1244 1352
rect 1278 1356 1284 1357
rect 1278 1352 1279 1356
rect 1283 1352 1284 1356
rect 1310 1355 1311 1359
rect 1315 1358 1316 1359
rect 1327 1359 1333 1360
rect 1327 1358 1328 1359
rect 1315 1356 1328 1358
rect 1315 1355 1316 1356
rect 1310 1354 1316 1355
rect 1327 1355 1328 1356
rect 1332 1355 1333 1359
rect 1327 1354 1333 1355
rect 1367 1359 1373 1360
rect 1367 1355 1368 1359
rect 1372 1358 1373 1359
rect 1390 1359 1396 1360
rect 1390 1358 1391 1359
rect 1372 1356 1391 1358
rect 1372 1355 1373 1356
rect 1367 1354 1373 1355
rect 1390 1355 1391 1356
rect 1395 1355 1396 1359
rect 1390 1354 1396 1355
rect 1423 1359 1429 1360
rect 1423 1355 1424 1359
rect 1428 1358 1429 1359
rect 1454 1359 1460 1360
rect 1454 1358 1455 1359
rect 1428 1356 1455 1358
rect 1428 1355 1429 1356
rect 1423 1354 1429 1355
rect 1454 1355 1455 1356
rect 1459 1355 1460 1359
rect 1454 1354 1460 1355
rect 1487 1359 1496 1360
rect 1487 1355 1488 1359
rect 1495 1355 1496 1359
rect 1487 1354 1496 1355
rect 1558 1359 1565 1360
rect 1558 1355 1559 1359
rect 1564 1355 1565 1359
rect 1558 1354 1565 1355
rect 1567 1359 1573 1360
rect 1567 1355 1568 1359
rect 1572 1358 1573 1359
rect 1631 1359 1637 1360
rect 1631 1358 1632 1359
rect 1572 1356 1632 1358
rect 1572 1355 1573 1356
rect 1567 1354 1573 1355
rect 1631 1355 1632 1356
rect 1636 1355 1637 1359
rect 1631 1354 1637 1355
rect 1639 1359 1645 1360
rect 1639 1355 1640 1359
rect 1644 1358 1645 1359
rect 1711 1359 1717 1360
rect 1711 1358 1712 1359
rect 1644 1356 1712 1358
rect 1644 1355 1645 1356
rect 1639 1354 1645 1355
rect 1711 1355 1712 1356
rect 1716 1355 1717 1359
rect 1711 1354 1717 1355
rect 1782 1359 1788 1360
rect 1782 1355 1783 1359
rect 1787 1358 1788 1359
rect 1791 1359 1797 1360
rect 1791 1358 1792 1359
rect 1787 1356 1792 1358
rect 1787 1355 1788 1356
rect 1782 1354 1788 1355
rect 1791 1355 1792 1356
rect 1796 1355 1797 1359
rect 1791 1354 1797 1355
rect 1799 1359 1805 1360
rect 1799 1355 1800 1359
rect 1804 1358 1805 1359
rect 1871 1359 1877 1360
rect 1871 1358 1872 1359
rect 1804 1356 1872 1358
rect 1804 1355 1805 1356
rect 1799 1354 1805 1355
rect 1871 1355 1872 1356
rect 1876 1355 1877 1359
rect 1871 1354 1877 1355
rect 1879 1359 1885 1360
rect 1879 1355 1880 1359
rect 1884 1358 1885 1359
rect 1959 1359 1965 1360
rect 1959 1358 1960 1359
rect 1884 1356 1960 1358
rect 1884 1355 1885 1356
rect 1879 1354 1885 1355
rect 1959 1355 1960 1356
rect 1964 1355 1965 1359
rect 1959 1354 1965 1355
rect 2047 1359 2053 1360
rect 2047 1355 2048 1359
rect 2052 1358 2053 1359
rect 2102 1359 2108 1360
rect 2102 1358 2103 1359
rect 2052 1356 2103 1358
rect 2052 1355 2053 1356
rect 2047 1354 2053 1355
rect 2102 1355 2103 1356
rect 2107 1355 2108 1359
rect 2135 1359 2141 1360
rect 2135 1358 2136 1359
rect 2102 1354 2108 1355
rect 2112 1356 2136 1358
rect 1278 1351 1284 1352
rect 1942 1351 1948 1352
rect 1942 1347 1943 1351
rect 1947 1350 1948 1351
rect 2112 1350 2114 1356
rect 2135 1355 2136 1356
rect 2140 1355 2141 1359
rect 2135 1354 2141 1355
rect 2223 1359 2229 1360
rect 2223 1355 2224 1359
rect 2228 1358 2229 1359
rect 2270 1359 2276 1360
rect 2270 1358 2271 1359
rect 2228 1356 2271 1358
rect 2228 1355 2229 1356
rect 2223 1354 2229 1355
rect 2270 1355 2271 1356
rect 2275 1355 2276 1359
rect 2270 1354 2276 1355
rect 2310 1359 2317 1360
rect 2310 1355 2311 1359
rect 2316 1355 2317 1359
rect 2310 1354 2317 1355
rect 2366 1359 2372 1360
rect 2366 1355 2367 1359
rect 2371 1358 2372 1359
rect 2383 1359 2389 1360
rect 2383 1358 2384 1359
rect 2371 1356 2384 1358
rect 2371 1355 2372 1356
rect 2366 1354 2372 1355
rect 2383 1355 2384 1356
rect 2388 1355 2389 1359
rect 2383 1354 2389 1355
rect 2406 1356 2412 1357
rect 2406 1352 2407 1356
rect 2411 1352 2412 1356
rect 2406 1351 2412 1352
rect 1947 1348 2114 1350
rect 1947 1347 1948 1348
rect 1942 1346 1948 1347
rect 166 1333 172 1334
rect 166 1329 167 1333
rect 171 1329 172 1333
rect 166 1328 172 1329
rect 206 1333 212 1334
rect 206 1329 207 1333
rect 211 1329 212 1333
rect 206 1328 212 1329
rect 246 1333 252 1334
rect 246 1329 247 1333
rect 251 1329 252 1333
rect 246 1328 252 1329
rect 302 1333 308 1334
rect 302 1329 303 1333
rect 307 1329 308 1333
rect 302 1328 308 1329
rect 366 1333 372 1334
rect 366 1329 367 1333
rect 371 1329 372 1333
rect 366 1328 372 1329
rect 438 1333 444 1334
rect 438 1329 439 1333
rect 443 1329 444 1333
rect 438 1328 444 1329
rect 518 1333 524 1334
rect 518 1329 519 1333
rect 523 1329 524 1333
rect 518 1328 524 1329
rect 598 1333 604 1334
rect 598 1329 599 1333
rect 603 1329 604 1333
rect 598 1328 604 1329
rect 678 1333 684 1334
rect 678 1329 679 1333
rect 683 1329 684 1333
rect 678 1328 684 1329
rect 750 1333 756 1334
rect 750 1329 751 1333
rect 755 1329 756 1333
rect 750 1328 756 1329
rect 822 1333 828 1334
rect 822 1329 823 1333
rect 827 1329 828 1333
rect 822 1328 828 1329
rect 886 1333 892 1334
rect 886 1329 887 1333
rect 891 1329 892 1333
rect 886 1328 892 1329
rect 950 1333 956 1334
rect 950 1329 951 1333
rect 955 1329 956 1333
rect 950 1328 956 1329
rect 1014 1333 1020 1334
rect 1014 1329 1015 1333
rect 1019 1329 1020 1333
rect 1014 1328 1020 1329
rect 1078 1333 1084 1334
rect 1078 1329 1079 1333
rect 1083 1329 1084 1333
rect 1078 1328 1084 1329
rect 1142 1333 1148 1334
rect 1142 1329 1143 1333
rect 1147 1329 1148 1333
rect 1142 1328 1148 1329
rect 1190 1333 1196 1334
rect 1190 1329 1191 1333
rect 1195 1329 1196 1333
rect 1190 1328 1196 1329
rect 1302 1333 1308 1334
rect 1302 1329 1303 1333
rect 1307 1329 1308 1333
rect 1302 1328 1308 1329
rect 1342 1333 1348 1334
rect 1342 1329 1343 1333
rect 1347 1329 1348 1333
rect 1342 1328 1348 1329
rect 1398 1333 1404 1334
rect 1398 1329 1399 1333
rect 1403 1329 1404 1333
rect 1398 1328 1404 1329
rect 1462 1333 1468 1334
rect 1462 1329 1463 1333
rect 1467 1329 1468 1333
rect 1462 1328 1468 1329
rect 1534 1333 1540 1334
rect 1534 1329 1535 1333
rect 1539 1329 1540 1333
rect 1534 1328 1540 1329
rect 1606 1333 1612 1334
rect 1606 1329 1607 1333
rect 1611 1329 1612 1333
rect 1606 1328 1612 1329
rect 1686 1333 1692 1334
rect 1686 1329 1687 1333
rect 1691 1329 1692 1333
rect 1686 1328 1692 1329
rect 1766 1333 1772 1334
rect 1766 1329 1767 1333
rect 1771 1329 1772 1333
rect 1766 1328 1772 1329
rect 1846 1333 1852 1334
rect 1846 1329 1847 1333
rect 1851 1329 1852 1333
rect 1846 1328 1852 1329
rect 1934 1333 1940 1334
rect 1934 1329 1935 1333
rect 1939 1329 1940 1333
rect 1934 1328 1940 1329
rect 2022 1333 2028 1334
rect 2022 1329 2023 1333
rect 2027 1329 2028 1333
rect 2022 1328 2028 1329
rect 2110 1333 2116 1334
rect 2110 1329 2111 1333
rect 2115 1329 2116 1333
rect 2110 1328 2116 1329
rect 2198 1333 2204 1334
rect 2198 1329 2199 1333
rect 2203 1329 2204 1333
rect 2198 1328 2204 1329
rect 2286 1333 2292 1334
rect 2286 1329 2287 1333
rect 2291 1329 2292 1333
rect 2286 1328 2292 1329
rect 2358 1333 2364 1334
rect 2358 1329 2359 1333
rect 2363 1329 2364 1333
rect 2358 1328 2364 1329
rect 163 1323 169 1324
rect 163 1319 164 1323
rect 168 1322 169 1323
rect 174 1323 180 1324
rect 174 1322 175 1323
rect 168 1320 175 1322
rect 168 1319 169 1320
rect 163 1318 169 1319
rect 174 1319 175 1320
rect 179 1319 180 1323
rect 174 1318 180 1319
rect 194 1323 200 1324
rect 194 1319 195 1323
rect 199 1322 200 1323
rect 203 1323 209 1324
rect 203 1322 204 1323
rect 199 1320 204 1322
rect 199 1319 200 1320
rect 194 1318 200 1319
rect 203 1319 204 1320
rect 208 1319 209 1323
rect 203 1318 209 1319
rect 234 1323 240 1324
rect 234 1319 235 1323
rect 239 1322 240 1323
rect 243 1323 249 1324
rect 243 1322 244 1323
rect 239 1320 244 1322
rect 239 1319 240 1320
rect 234 1318 240 1319
rect 243 1319 244 1320
rect 248 1319 249 1323
rect 243 1318 249 1319
rect 294 1323 305 1324
rect 294 1319 295 1323
rect 299 1319 300 1323
rect 304 1319 305 1323
rect 294 1318 305 1319
rect 363 1323 369 1324
rect 363 1319 364 1323
rect 368 1322 369 1323
rect 374 1323 380 1324
rect 374 1322 375 1323
rect 368 1320 375 1322
rect 368 1319 369 1320
rect 363 1318 369 1319
rect 374 1319 375 1320
rect 379 1319 380 1323
rect 374 1318 380 1319
rect 430 1323 441 1324
rect 430 1319 431 1323
rect 435 1319 436 1323
rect 440 1319 441 1323
rect 430 1318 441 1319
rect 510 1323 521 1324
rect 510 1319 511 1323
rect 515 1319 516 1323
rect 520 1319 521 1323
rect 510 1318 521 1319
rect 590 1323 601 1324
rect 590 1319 591 1323
rect 595 1319 596 1323
rect 600 1319 601 1323
rect 590 1318 601 1319
rect 675 1323 681 1324
rect 675 1319 676 1323
rect 680 1319 681 1323
rect 675 1318 681 1319
rect 742 1323 753 1324
rect 742 1319 743 1323
rect 747 1319 748 1323
rect 752 1319 753 1323
rect 742 1318 753 1319
rect 814 1323 825 1324
rect 814 1319 815 1323
rect 819 1319 820 1323
rect 824 1319 825 1323
rect 814 1318 825 1319
rect 878 1323 889 1324
rect 878 1319 879 1323
rect 883 1319 884 1323
rect 888 1319 889 1323
rect 878 1318 889 1319
rect 942 1323 953 1324
rect 942 1319 943 1323
rect 947 1319 948 1323
rect 952 1319 953 1323
rect 942 1318 953 1319
rect 1006 1323 1017 1324
rect 1006 1319 1007 1323
rect 1011 1319 1012 1323
rect 1016 1319 1017 1323
rect 1006 1318 1017 1319
rect 1075 1323 1081 1324
rect 1075 1319 1076 1323
rect 1080 1322 1081 1323
rect 1086 1323 1092 1324
rect 1086 1322 1087 1323
rect 1080 1320 1087 1322
rect 1080 1319 1081 1320
rect 1075 1318 1081 1319
rect 1086 1319 1087 1320
rect 1091 1319 1092 1323
rect 1086 1318 1092 1319
rect 1134 1323 1145 1324
rect 1134 1319 1135 1323
rect 1139 1319 1140 1323
rect 1144 1319 1145 1323
rect 1134 1318 1145 1319
rect 1182 1323 1193 1324
rect 1182 1319 1183 1323
rect 1187 1319 1188 1323
rect 1192 1319 1193 1323
rect 1182 1318 1193 1319
rect 1230 1323 1236 1324
rect 1230 1319 1231 1323
rect 1235 1322 1236 1323
rect 1299 1323 1305 1324
rect 1299 1322 1300 1323
rect 1235 1320 1300 1322
rect 1235 1319 1236 1320
rect 1230 1318 1236 1319
rect 1299 1319 1300 1320
rect 1304 1319 1305 1323
rect 1299 1318 1305 1319
rect 1339 1323 1345 1324
rect 1339 1319 1340 1323
rect 1344 1322 1345 1323
rect 1350 1323 1356 1324
rect 1350 1322 1351 1323
rect 1344 1320 1351 1322
rect 1344 1319 1345 1320
rect 1339 1318 1345 1319
rect 1350 1319 1351 1320
rect 1355 1319 1356 1323
rect 1350 1318 1356 1319
rect 1390 1323 1401 1324
rect 1390 1319 1391 1323
rect 1395 1319 1396 1323
rect 1400 1319 1401 1323
rect 1390 1318 1401 1319
rect 1454 1323 1465 1324
rect 1454 1319 1455 1323
rect 1459 1319 1460 1323
rect 1464 1319 1465 1323
rect 1454 1318 1465 1319
rect 1531 1323 1537 1324
rect 1531 1319 1532 1323
rect 1536 1322 1537 1323
rect 1567 1323 1573 1324
rect 1567 1322 1568 1323
rect 1536 1320 1568 1322
rect 1536 1319 1537 1320
rect 1531 1318 1537 1319
rect 1567 1319 1568 1320
rect 1572 1319 1573 1323
rect 1567 1318 1573 1319
rect 1603 1323 1609 1324
rect 1603 1319 1604 1323
rect 1608 1322 1609 1323
rect 1639 1323 1645 1324
rect 1639 1322 1640 1323
rect 1608 1320 1640 1322
rect 1608 1319 1609 1320
rect 1603 1318 1609 1319
rect 1639 1319 1640 1320
rect 1644 1319 1645 1323
rect 1639 1318 1645 1319
rect 1683 1323 1689 1324
rect 1683 1319 1684 1323
rect 1688 1322 1689 1323
rect 1754 1323 1760 1324
rect 1754 1322 1755 1323
rect 1688 1320 1755 1322
rect 1688 1319 1689 1320
rect 1683 1318 1689 1319
rect 1754 1319 1755 1320
rect 1759 1319 1760 1323
rect 1754 1318 1760 1319
rect 1763 1323 1769 1324
rect 1763 1319 1764 1323
rect 1768 1322 1769 1323
rect 1799 1323 1805 1324
rect 1799 1322 1800 1323
rect 1768 1320 1800 1322
rect 1768 1319 1769 1320
rect 1763 1318 1769 1319
rect 1799 1319 1800 1320
rect 1804 1319 1805 1323
rect 1799 1318 1805 1319
rect 1843 1323 1849 1324
rect 1843 1319 1844 1323
rect 1848 1322 1849 1323
rect 1879 1323 1885 1324
rect 1879 1322 1880 1323
rect 1848 1320 1880 1322
rect 1848 1319 1849 1320
rect 1843 1318 1849 1319
rect 1879 1319 1880 1320
rect 1884 1319 1885 1323
rect 1879 1318 1885 1319
rect 1931 1323 1937 1324
rect 1931 1319 1932 1323
rect 1936 1322 1937 1323
rect 1942 1323 1948 1324
rect 1942 1322 1943 1323
rect 1936 1320 1943 1322
rect 1936 1319 1937 1320
rect 1931 1318 1937 1319
rect 1942 1319 1943 1320
rect 1947 1319 1948 1323
rect 1942 1318 1948 1319
rect 2014 1323 2025 1324
rect 2014 1319 2015 1323
rect 2019 1319 2020 1323
rect 2024 1319 2025 1323
rect 2014 1318 2025 1319
rect 2102 1323 2113 1324
rect 2102 1319 2103 1323
rect 2107 1319 2108 1323
rect 2112 1319 2113 1323
rect 2102 1318 2113 1319
rect 2195 1323 2201 1324
rect 2195 1319 2196 1323
rect 2200 1322 2201 1323
rect 2262 1323 2268 1324
rect 2262 1322 2263 1323
rect 2200 1320 2263 1322
rect 2200 1319 2201 1320
rect 2195 1318 2201 1319
rect 2262 1319 2263 1320
rect 2267 1319 2268 1323
rect 2262 1318 2268 1319
rect 2270 1323 2276 1324
rect 2270 1319 2271 1323
rect 2275 1322 2276 1323
rect 2283 1323 2289 1324
rect 2283 1322 2284 1323
rect 2275 1320 2284 1322
rect 2275 1319 2276 1320
rect 2270 1318 2276 1319
rect 2283 1319 2284 1320
rect 2288 1319 2289 1323
rect 2283 1318 2289 1319
rect 2355 1323 2361 1324
rect 2355 1319 2356 1323
rect 2360 1322 2361 1323
rect 2374 1323 2380 1324
rect 2374 1322 2375 1323
rect 2360 1320 2375 1322
rect 2360 1319 2361 1320
rect 2355 1318 2361 1319
rect 2374 1319 2375 1320
rect 2379 1319 2380 1323
rect 2374 1318 2380 1319
rect 679 1314 681 1318
rect 1022 1315 1028 1316
rect 1022 1314 1023 1315
rect 679 1312 1023 1314
rect 1022 1311 1023 1312
rect 1027 1311 1028 1315
rect 1022 1310 1028 1311
rect 1299 1311 1305 1312
rect 179 1307 185 1308
rect 179 1303 180 1307
rect 184 1306 185 1307
rect 218 1307 224 1308
rect 218 1306 219 1307
rect 184 1304 219 1306
rect 184 1303 185 1304
rect 179 1302 185 1303
rect 218 1303 219 1304
rect 223 1303 224 1307
rect 218 1302 224 1303
rect 227 1307 233 1308
rect 227 1303 228 1307
rect 232 1306 233 1307
rect 254 1307 260 1308
rect 254 1306 255 1307
rect 232 1304 255 1306
rect 232 1303 233 1304
rect 227 1302 233 1303
rect 254 1303 255 1304
rect 259 1303 260 1307
rect 254 1302 260 1303
rect 278 1307 289 1308
rect 278 1303 279 1307
rect 283 1303 284 1307
rect 288 1303 289 1307
rect 278 1302 289 1303
rect 314 1307 320 1308
rect 314 1303 315 1307
rect 319 1306 320 1307
rect 347 1307 353 1308
rect 347 1306 348 1307
rect 319 1304 348 1306
rect 319 1303 320 1304
rect 314 1302 320 1303
rect 347 1303 348 1304
rect 352 1303 353 1307
rect 347 1302 353 1303
rect 378 1307 384 1308
rect 378 1303 379 1307
rect 383 1306 384 1307
rect 419 1307 425 1308
rect 419 1306 420 1307
rect 383 1304 420 1306
rect 383 1303 384 1304
rect 378 1302 384 1303
rect 419 1303 420 1304
rect 424 1303 425 1307
rect 419 1302 425 1303
rect 450 1307 456 1308
rect 450 1303 451 1307
rect 455 1306 456 1307
rect 491 1307 497 1308
rect 491 1306 492 1307
rect 455 1304 492 1306
rect 455 1303 456 1304
rect 450 1302 456 1303
rect 491 1303 492 1304
rect 496 1303 497 1307
rect 491 1302 497 1303
rect 535 1307 541 1308
rect 535 1303 536 1307
rect 540 1306 541 1307
rect 563 1307 569 1308
rect 563 1306 564 1307
rect 540 1304 564 1306
rect 540 1303 541 1304
rect 535 1302 541 1303
rect 563 1303 564 1304
rect 568 1303 569 1307
rect 563 1302 569 1303
rect 635 1307 641 1308
rect 635 1303 636 1307
rect 640 1306 641 1307
rect 654 1307 660 1308
rect 654 1306 655 1307
rect 640 1304 655 1306
rect 640 1303 641 1304
rect 635 1302 641 1303
rect 654 1303 655 1304
rect 659 1303 660 1307
rect 654 1302 660 1303
rect 666 1307 672 1308
rect 666 1303 667 1307
rect 671 1306 672 1307
rect 699 1307 705 1308
rect 699 1306 700 1307
rect 671 1304 700 1306
rect 671 1303 672 1304
rect 666 1302 672 1303
rect 699 1303 700 1304
rect 704 1303 705 1307
rect 699 1302 705 1303
rect 730 1307 736 1308
rect 730 1303 731 1307
rect 735 1306 736 1307
rect 763 1307 769 1308
rect 763 1306 764 1307
rect 735 1304 764 1306
rect 735 1303 736 1304
rect 730 1302 736 1303
rect 763 1303 764 1304
rect 768 1303 769 1307
rect 763 1302 769 1303
rect 794 1307 800 1308
rect 794 1303 795 1307
rect 799 1306 800 1307
rect 819 1307 825 1308
rect 819 1306 820 1307
rect 799 1304 820 1306
rect 799 1303 800 1304
rect 794 1302 800 1303
rect 819 1303 820 1304
rect 824 1303 825 1307
rect 819 1302 825 1303
rect 850 1307 856 1308
rect 850 1303 851 1307
rect 855 1306 856 1307
rect 875 1307 881 1308
rect 875 1306 876 1307
rect 855 1304 876 1306
rect 855 1303 856 1304
rect 850 1302 856 1303
rect 875 1303 876 1304
rect 880 1303 881 1307
rect 875 1302 881 1303
rect 906 1307 912 1308
rect 906 1303 907 1307
rect 911 1306 912 1307
rect 931 1307 937 1308
rect 931 1306 932 1307
rect 911 1304 932 1306
rect 911 1303 912 1304
rect 906 1302 912 1303
rect 931 1303 932 1304
rect 936 1303 937 1307
rect 931 1302 937 1303
rect 962 1307 968 1308
rect 962 1303 963 1307
rect 967 1306 968 1307
rect 995 1307 1001 1308
rect 995 1306 996 1307
rect 967 1304 996 1306
rect 967 1303 968 1304
rect 962 1302 968 1303
rect 995 1303 996 1304
rect 1000 1303 1001 1307
rect 1299 1307 1300 1311
rect 1304 1310 1305 1311
rect 1310 1311 1316 1312
rect 1310 1310 1311 1311
rect 1304 1308 1311 1310
rect 1304 1307 1305 1308
rect 1299 1306 1305 1307
rect 1310 1307 1311 1308
rect 1315 1307 1316 1311
rect 1310 1306 1316 1307
rect 1330 1311 1336 1312
rect 1330 1307 1331 1311
rect 1335 1310 1336 1311
rect 1339 1311 1345 1312
rect 1339 1310 1340 1311
rect 1335 1308 1340 1310
rect 1335 1307 1336 1308
rect 1330 1306 1336 1307
rect 1339 1307 1340 1308
rect 1344 1307 1345 1311
rect 1339 1306 1345 1307
rect 1370 1311 1376 1312
rect 1370 1307 1371 1311
rect 1375 1310 1376 1311
rect 1379 1311 1385 1312
rect 1379 1310 1380 1311
rect 1375 1308 1380 1310
rect 1375 1307 1376 1308
rect 1370 1306 1376 1307
rect 1379 1307 1380 1308
rect 1384 1307 1385 1311
rect 1379 1306 1385 1307
rect 1410 1311 1416 1312
rect 1410 1307 1411 1311
rect 1415 1310 1416 1311
rect 1419 1311 1425 1312
rect 1419 1310 1420 1311
rect 1415 1308 1420 1310
rect 1415 1307 1416 1308
rect 1410 1306 1416 1307
rect 1419 1307 1420 1308
rect 1424 1307 1425 1311
rect 1419 1306 1425 1307
rect 1446 1311 1452 1312
rect 1446 1307 1447 1311
rect 1451 1310 1452 1311
rect 1459 1311 1465 1312
rect 1459 1310 1460 1311
rect 1451 1308 1460 1310
rect 1451 1307 1452 1308
rect 1446 1306 1452 1307
rect 1459 1307 1460 1308
rect 1464 1307 1465 1311
rect 1459 1306 1465 1307
rect 1490 1311 1496 1312
rect 1490 1307 1491 1311
rect 1495 1310 1496 1311
rect 1499 1311 1505 1312
rect 1499 1310 1500 1311
rect 1495 1308 1500 1310
rect 1495 1307 1496 1308
rect 1490 1306 1496 1307
rect 1499 1307 1500 1308
rect 1504 1307 1505 1311
rect 1499 1306 1505 1307
rect 1526 1311 1532 1312
rect 1526 1307 1527 1311
rect 1531 1310 1532 1311
rect 1539 1311 1545 1312
rect 1539 1310 1540 1311
rect 1531 1308 1540 1310
rect 1531 1307 1532 1308
rect 1526 1306 1532 1307
rect 1539 1307 1540 1308
rect 1544 1307 1545 1311
rect 1539 1306 1545 1307
rect 1550 1311 1556 1312
rect 1550 1307 1551 1311
rect 1555 1310 1556 1311
rect 1579 1311 1585 1312
rect 1579 1310 1580 1311
rect 1555 1308 1580 1310
rect 1555 1307 1556 1308
rect 1550 1306 1556 1307
rect 1579 1307 1580 1308
rect 1584 1307 1585 1311
rect 1579 1306 1585 1307
rect 1614 1311 1625 1312
rect 1614 1307 1615 1311
rect 1619 1307 1620 1311
rect 1624 1307 1625 1311
rect 1614 1306 1625 1307
rect 1650 1311 1656 1312
rect 1650 1307 1651 1311
rect 1655 1310 1656 1311
rect 1675 1311 1681 1312
rect 1675 1310 1676 1311
rect 1655 1308 1676 1310
rect 1655 1307 1656 1308
rect 1650 1306 1656 1307
rect 1675 1307 1676 1308
rect 1680 1307 1681 1311
rect 1675 1306 1681 1307
rect 1719 1311 1725 1312
rect 1719 1307 1720 1311
rect 1724 1310 1725 1311
rect 1731 1311 1737 1312
rect 1731 1310 1732 1311
rect 1724 1308 1732 1310
rect 1724 1307 1725 1308
rect 1719 1306 1725 1307
rect 1731 1307 1732 1308
rect 1736 1307 1737 1311
rect 1731 1306 1737 1307
rect 1782 1311 1793 1312
rect 1782 1307 1783 1311
rect 1787 1307 1788 1311
rect 1792 1307 1793 1311
rect 1782 1306 1793 1307
rect 1818 1311 1824 1312
rect 1818 1307 1819 1311
rect 1823 1310 1824 1311
rect 1843 1311 1849 1312
rect 1843 1310 1844 1311
rect 1823 1308 1844 1310
rect 1823 1307 1824 1308
rect 1818 1306 1824 1307
rect 1843 1307 1844 1308
rect 1848 1307 1849 1311
rect 1843 1306 1849 1307
rect 1874 1311 1880 1312
rect 1874 1307 1875 1311
rect 1879 1310 1880 1311
rect 1899 1311 1905 1312
rect 1899 1310 1900 1311
rect 1879 1308 1900 1310
rect 1879 1307 1880 1308
rect 1874 1306 1880 1307
rect 1899 1307 1900 1308
rect 1904 1307 1905 1311
rect 1899 1306 1905 1307
rect 1943 1311 1949 1312
rect 1943 1307 1944 1311
rect 1948 1310 1949 1311
rect 1963 1311 1969 1312
rect 1963 1310 1964 1311
rect 1948 1308 1964 1310
rect 1948 1307 1949 1308
rect 1943 1306 1949 1307
rect 1963 1307 1964 1308
rect 1968 1307 1969 1311
rect 1963 1306 1969 1307
rect 1994 1311 2000 1312
rect 1994 1307 1995 1311
rect 1999 1310 2000 1311
rect 2035 1311 2041 1312
rect 2035 1310 2036 1311
rect 1999 1308 2036 1310
rect 1999 1307 2000 1308
rect 1994 1306 2000 1307
rect 2035 1307 2036 1308
rect 2040 1307 2041 1311
rect 2035 1306 2041 1307
rect 2066 1311 2072 1312
rect 2066 1307 2067 1311
rect 2071 1310 2072 1311
rect 2115 1311 2121 1312
rect 2115 1310 2116 1311
rect 2071 1308 2116 1310
rect 2071 1307 2072 1308
rect 2066 1306 2072 1307
rect 2115 1307 2116 1308
rect 2120 1307 2121 1311
rect 2115 1306 2121 1307
rect 2146 1311 2152 1312
rect 2146 1307 2147 1311
rect 2151 1310 2152 1311
rect 2195 1311 2201 1312
rect 2195 1310 2196 1311
rect 2151 1308 2196 1310
rect 2151 1307 2152 1308
rect 2146 1306 2152 1307
rect 2195 1307 2196 1308
rect 2200 1307 2201 1311
rect 2195 1306 2201 1307
rect 2250 1311 2256 1312
rect 2250 1307 2251 1311
rect 2255 1310 2256 1311
rect 2283 1311 2289 1312
rect 2283 1310 2284 1311
rect 2255 1308 2284 1310
rect 2255 1307 2256 1308
rect 2250 1306 2256 1307
rect 2283 1307 2284 1308
rect 2288 1307 2289 1311
rect 2283 1306 2289 1307
rect 2355 1311 2361 1312
rect 2355 1307 2356 1311
rect 2360 1310 2361 1311
rect 2366 1311 2372 1312
rect 2366 1310 2367 1311
rect 2360 1308 2367 1310
rect 2360 1307 2361 1308
rect 2355 1306 2361 1307
rect 2366 1307 2367 1308
rect 2371 1307 2372 1311
rect 2366 1306 2372 1307
rect 995 1302 1001 1303
rect 1302 1303 1308 1304
rect 182 1299 188 1300
rect 182 1295 183 1299
rect 187 1295 188 1299
rect 182 1294 188 1295
rect 230 1299 236 1300
rect 230 1295 231 1299
rect 235 1295 236 1299
rect 230 1294 236 1295
rect 286 1299 292 1300
rect 286 1295 287 1299
rect 291 1295 292 1299
rect 286 1294 292 1295
rect 350 1299 356 1300
rect 350 1295 351 1299
rect 355 1295 356 1299
rect 350 1294 356 1295
rect 422 1299 428 1300
rect 422 1295 423 1299
rect 427 1295 428 1299
rect 422 1294 428 1295
rect 494 1299 500 1300
rect 494 1295 495 1299
rect 499 1295 500 1299
rect 494 1294 500 1295
rect 566 1299 572 1300
rect 566 1295 567 1299
rect 571 1295 572 1299
rect 566 1294 572 1295
rect 638 1299 644 1300
rect 638 1295 639 1299
rect 643 1295 644 1299
rect 638 1294 644 1295
rect 702 1299 708 1300
rect 702 1295 703 1299
rect 707 1295 708 1299
rect 702 1294 708 1295
rect 766 1299 772 1300
rect 766 1295 767 1299
rect 771 1295 772 1299
rect 766 1294 772 1295
rect 822 1299 828 1300
rect 822 1295 823 1299
rect 827 1295 828 1299
rect 822 1294 828 1295
rect 878 1299 884 1300
rect 878 1295 879 1299
rect 883 1295 884 1299
rect 878 1294 884 1295
rect 934 1299 940 1300
rect 934 1295 935 1299
rect 939 1295 940 1299
rect 934 1294 940 1295
rect 998 1299 1004 1300
rect 998 1295 999 1299
rect 1003 1295 1004 1299
rect 1302 1299 1303 1303
rect 1307 1299 1308 1303
rect 1302 1298 1308 1299
rect 1342 1303 1348 1304
rect 1342 1299 1343 1303
rect 1347 1299 1348 1303
rect 1342 1298 1348 1299
rect 1382 1303 1388 1304
rect 1382 1299 1383 1303
rect 1387 1299 1388 1303
rect 1382 1298 1388 1299
rect 1422 1303 1428 1304
rect 1422 1299 1423 1303
rect 1427 1299 1428 1303
rect 1422 1298 1428 1299
rect 1462 1303 1468 1304
rect 1462 1299 1463 1303
rect 1467 1299 1468 1303
rect 1462 1298 1468 1299
rect 1502 1303 1508 1304
rect 1502 1299 1503 1303
rect 1507 1299 1508 1303
rect 1502 1298 1508 1299
rect 1542 1303 1548 1304
rect 1542 1299 1543 1303
rect 1547 1299 1548 1303
rect 1542 1298 1548 1299
rect 1582 1303 1588 1304
rect 1582 1299 1583 1303
rect 1587 1299 1588 1303
rect 1582 1298 1588 1299
rect 1622 1303 1628 1304
rect 1622 1299 1623 1303
rect 1627 1299 1628 1303
rect 1622 1298 1628 1299
rect 1678 1303 1684 1304
rect 1678 1299 1679 1303
rect 1683 1299 1684 1303
rect 1678 1298 1684 1299
rect 1734 1303 1740 1304
rect 1734 1299 1735 1303
rect 1739 1299 1740 1303
rect 1734 1298 1740 1299
rect 1790 1303 1796 1304
rect 1790 1299 1791 1303
rect 1795 1299 1796 1303
rect 1790 1298 1796 1299
rect 1846 1303 1852 1304
rect 1846 1299 1847 1303
rect 1851 1299 1852 1303
rect 1846 1298 1852 1299
rect 1902 1303 1908 1304
rect 1902 1299 1903 1303
rect 1907 1299 1908 1303
rect 1902 1298 1908 1299
rect 1966 1303 1972 1304
rect 1966 1299 1967 1303
rect 1971 1299 1972 1303
rect 1966 1298 1972 1299
rect 2038 1303 2044 1304
rect 2038 1299 2039 1303
rect 2043 1299 2044 1303
rect 2038 1298 2044 1299
rect 2118 1303 2124 1304
rect 2118 1299 2119 1303
rect 2123 1299 2124 1303
rect 2118 1298 2124 1299
rect 2198 1303 2204 1304
rect 2198 1299 2199 1303
rect 2203 1299 2204 1303
rect 2198 1298 2204 1299
rect 2286 1303 2292 1304
rect 2286 1299 2287 1303
rect 2291 1299 2292 1303
rect 2286 1298 2292 1299
rect 2358 1303 2364 1304
rect 2358 1299 2359 1303
rect 2363 1299 2364 1303
rect 2358 1298 2364 1299
rect 998 1294 1004 1295
rect 1550 1283 1556 1284
rect 1550 1282 1551 1283
rect 1278 1280 1284 1281
rect 110 1276 116 1277
rect 1238 1276 1244 1277
rect 110 1272 111 1276
rect 115 1272 116 1276
rect 535 1275 541 1276
rect 535 1274 536 1275
rect 519 1273 536 1274
rect 110 1271 116 1272
rect 174 1271 180 1272
rect 174 1267 175 1271
rect 179 1270 180 1271
rect 207 1271 213 1272
rect 207 1270 208 1271
rect 179 1268 208 1270
rect 179 1267 180 1268
rect 174 1266 180 1267
rect 207 1267 208 1268
rect 212 1267 213 1271
rect 207 1266 213 1267
rect 218 1271 224 1272
rect 218 1267 219 1271
rect 223 1270 224 1271
rect 255 1271 261 1272
rect 255 1270 256 1271
rect 223 1268 256 1270
rect 223 1267 224 1268
rect 218 1266 224 1267
rect 255 1267 256 1268
rect 260 1267 261 1271
rect 255 1266 261 1267
rect 311 1271 320 1272
rect 311 1267 312 1271
rect 319 1267 320 1271
rect 311 1266 320 1267
rect 375 1271 384 1272
rect 375 1267 376 1271
rect 383 1267 384 1271
rect 375 1266 384 1267
rect 447 1271 456 1272
rect 447 1267 448 1271
rect 455 1267 456 1271
rect 519 1269 520 1273
rect 524 1272 536 1273
rect 524 1269 525 1272
rect 535 1271 536 1272
rect 540 1271 541 1275
rect 1238 1272 1239 1276
rect 1243 1272 1244 1276
rect 1278 1276 1279 1280
rect 1283 1276 1284 1280
rect 1520 1280 1551 1282
rect 1278 1275 1284 1276
rect 1327 1275 1336 1276
rect 535 1270 541 1271
rect 582 1271 588 1272
rect 519 1268 525 1269
rect 447 1266 456 1267
rect 582 1267 583 1271
rect 587 1270 588 1271
rect 591 1271 597 1272
rect 591 1270 592 1271
rect 587 1268 592 1270
rect 587 1267 588 1268
rect 582 1266 588 1267
rect 591 1267 592 1268
rect 596 1267 597 1271
rect 591 1266 597 1267
rect 663 1271 672 1272
rect 663 1267 664 1271
rect 671 1267 672 1271
rect 663 1266 672 1267
rect 727 1271 736 1272
rect 727 1267 728 1271
rect 735 1267 736 1271
rect 727 1266 736 1267
rect 791 1271 800 1272
rect 791 1267 792 1271
rect 799 1267 800 1271
rect 791 1266 800 1267
rect 847 1271 856 1272
rect 847 1267 848 1271
rect 855 1267 856 1271
rect 847 1266 856 1267
rect 903 1271 912 1272
rect 903 1267 904 1271
rect 911 1267 912 1271
rect 903 1266 912 1267
rect 959 1271 968 1272
rect 959 1267 960 1271
rect 967 1267 968 1271
rect 959 1266 968 1267
rect 1022 1271 1029 1272
rect 1238 1271 1244 1272
rect 1327 1271 1328 1275
rect 1335 1271 1336 1275
rect 1022 1267 1023 1271
rect 1028 1267 1029 1271
rect 1327 1270 1336 1271
rect 1367 1275 1376 1276
rect 1367 1271 1368 1275
rect 1375 1271 1376 1275
rect 1367 1270 1376 1271
rect 1407 1275 1416 1276
rect 1407 1271 1408 1275
rect 1415 1271 1416 1275
rect 1407 1270 1416 1271
rect 1446 1275 1453 1276
rect 1446 1271 1447 1275
rect 1452 1271 1453 1275
rect 1446 1270 1453 1271
rect 1487 1275 1493 1276
rect 1487 1271 1488 1275
rect 1492 1274 1493 1275
rect 1520 1274 1522 1280
rect 1550 1279 1551 1280
rect 1555 1279 1556 1283
rect 1550 1278 1556 1279
rect 2406 1280 2412 1281
rect 2406 1276 2407 1280
rect 2411 1276 2412 1280
rect 1492 1272 1522 1274
rect 1526 1275 1533 1276
rect 1492 1271 1493 1272
rect 1487 1270 1493 1271
rect 1526 1271 1527 1275
rect 1532 1271 1533 1275
rect 1526 1270 1533 1271
rect 1567 1275 1576 1276
rect 1567 1271 1568 1275
rect 1575 1271 1576 1275
rect 1567 1270 1576 1271
rect 1607 1275 1616 1276
rect 1607 1271 1608 1275
rect 1615 1271 1616 1275
rect 1607 1270 1616 1271
rect 1647 1275 1656 1276
rect 1647 1271 1648 1275
rect 1655 1271 1656 1275
rect 1647 1270 1656 1271
rect 1703 1275 1709 1276
rect 1703 1271 1704 1275
rect 1708 1274 1709 1275
rect 1719 1275 1725 1276
rect 1719 1274 1720 1275
rect 1708 1272 1720 1274
rect 1708 1271 1709 1272
rect 1703 1270 1709 1271
rect 1719 1271 1720 1272
rect 1724 1271 1725 1275
rect 1719 1270 1725 1271
rect 1754 1275 1765 1276
rect 1754 1271 1755 1275
rect 1759 1271 1760 1275
rect 1764 1271 1765 1275
rect 1754 1270 1765 1271
rect 1815 1275 1824 1276
rect 1815 1271 1816 1275
rect 1823 1271 1824 1275
rect 1815 1270 1824 1271
rect 1871 1275 1880 1276
rect 1871 1271 1872 1275
rect 1879 1271 1880 1275
rect 1871 1270 1880 1271
rect 1927 1275 1933 1276
rect 1927 1271 1928 1275
rect 1932 1274 1933 1275
rect 1943 1275 1949 1276
rect 1943 1274 1944 1275
rect 1932 1272 1944 1274
rect 1932 1271 1933 1272
rect 1927 1270 1933 1271
rect 1943 1271 1944 1272
rect 1948 1271 1949 1275
rect 1943 1270 1949 1271
rect 1991 1275 2000 1276
rect 1991 1271 1992 1275
rect 1999 1271 2000 1275
rect 1991 1270 2000 1271
rect 2063 1275 2072 1276
rect 2063 1271 2064 1275
rect 2071 1271 2072 1275
rect 2063 1270 2072 1271
rect 2143 1275 2152 1276
rect 2143 1271 2144 1275
rect 2151 1271 2152 1275
rect 2223 1275 2229 1276
rect 2223 1274 2224 1275
rect 2143 1270 2152 1271
rect 2156 1272 2224 1274
rect 1022 1266 1029 1267
rect 1806 1267 1812 1268
rect 1278 1263 1284 1264
rect 110 1259 116 1260
rect 110 1255 111 1259
rect 115 1255 116 1259
rect 110 1254 116 1255
rect 1238 1259 1244 1260
rect 1238 1255 1239 1259
rect 1243 1255 1244 1259
rect 1278 1259 1279 1263
rect 1283 1259 1284 1263
rect 1806 1263 1807 1267
rect 1811 1266 1812 1267
rect 2156 1266 2158 1272
rect 2223 1271 2224 1272
rect 2228 1271 2229 1275
rect 2223 1270 2229 1271
rect 2262 1275 2268 1276
rect 2262 1271 2263 1275
rect 2267 1274 2268 1275
rect 2311 1275 2317 1276
rect 2311 1274 2312 1275
rect 2267 1272 2312 1274
rect 2267 1271 2268 1272
rect 2262 1270 2268 1271
rect 2311 1271 2312 1272
rect 2316 1271 2317 1275
rect 2311 1270 2317 1271
rect 2366 1275 2372 1276
rect 2366 1271 2367 1275
rect 2371 1274 2372 1275
rect 2383 1275 2389 1276
rect 2406 1275 2412 1276
rect 2383 1274 2384 1275
rect 2371 1272 2384 1274
rect 2371 1271 2372 1272
rect 2366 1270 2372 1271
rect 2383 1271 2384 1272
rect 2388 1271 2389 1275
rect 2383 1270 2389 1271
rect 1811 1264 2158 1266
rect 1811 1263 1812 1264
rect 1806 1262 1812 1263
rect 2406 1263 2412 1264
rect 1278 1258 1284 1259
rect 2406 1259 2407 1263
rect 2411 1259 2412 1263
rect 2406 1258 2412 1259
rect 1238 1254 1244 1255
rect 1302 1256 1308 1257
rect 182 1252 188 1253
rect 182 1248 183 1252
rect 187 1248 188 1252
rect 182 1247 188 1248
rect 230 1252 236 1253
rect 230 1248 231 1252
rect 235 1248 236 1252
rect 230 1247 236 1248
rect 286 1252 292 1253
rect 286 1248 287 1252
rect 291 1248 292 1252
rect 286 1247 292 1248
rect 350 1252 356 1253
rect 350 1248 351 1252
rect 355 1248 356 1252
rect 350 1247 356 1248
rect 422 1252 428 1253
rect 422 1248 423 1252
rect 427 1248 428 1252
rect 422 1247 428 1248
rect 494 1252 500 1253
rect 494 1248 495 1252
rect 499 1248 500 1252
rect 494 1247 500 1248
rect 566 1252 572 1253
rect 566 1248 567 1252
rect 571 1248 572 1252
rect 566 1247 572 1248
rect 638 1252 644 1253
rect 638 1248 639 1252
rect 643 1248 644 1252
rect 638 1247 644 1248
rect 702 1252 708 1253
rect 702 1248 703 1252
rect 707 1248 708 1252
rect 702 1247 708 1248
rect 766 1252 772 1253
rect 766 1248 767 1252
rect 771 1248 772 1252
rect 766 1247 772 1248
rect 822 1252 828 1253
rect 822 1248 823 1252
rect 827 1248 828 1252
rect 822 1247 828 1248
rect 878 1252 884 1253
rect 878 1248 879 1252
rect 883 1248 884 1252
rect 878 1247 884 1248
rect 934 1252 940 1253
rect 934 1248 935 1252
rect 939 1248 940 1252
rect 934 1247 940 1248
rect 998 1252 1004 1253
rect 998 1248 999 1252
rect 1003 1248 1004 1252
rect 1302 1252 1303 1256
rect 1307 1252 1308 1256
rect 1302 1251 1308 1252
rect 1342 1256 1348 1257
rect 1342 1252 1343 1256
rect 1347 1252 1348 1256
rect 1342 1251 1348 1252
rect 1382 1256 1388 1257
rect 1382 1252 1383 1256
rect 1387 1252 1388 1256
rect 1382 1251 1388 1252
rect 1422 1256 1428 1257
rect 1422 1252 1423 1256
rect 1427 1252 1428 1256
rect 1422 1251 1428 1252
rect 1462 1256 1468 1257
rect 1462 1252 1463 1256
rect 1467 1252 1468 1256
rect 1462 1251 1468 1252
rect 1502 1256 1508 1257
rect 1502 1252 1503 1256
rect 1507 1252 1508 1256
rect 1502 1251 1508 1252
rect 1542 1256 1548 1257
rect 1542 1252 1543 1256
rect 1547 1252 1548 1256
rect 1542 1251 1548 1252
rect 1582 1256 1588 1257
rect 1582 1252 1583 1256
rect 1587 1252 1588 1256
rect 1582 1251 1588 1252
rect 1622 1256 1628 1257
rect 1622 1252 1623 1256
rect 1627 1252 1628 1256
rect 1622 1251 1628 1252
rect 1678 1256 1684 1257
rect 1678 1252 1679 1256
rect 1683 1252 1684 1256
rect 1678 1251 1684 1252
rect 1734 1256 1740 1257
rect 1734 1252 1735 1256
rect 1739 1252 1740 1256
rect 1734 1251 1740 1252
rect 1790 1256 1796 1257
rect 1790 1252 1791 1256
rect 1795 1252 1796 1256
rect 1790 1251 1796 1252
rect 1846 1256 1852 1257
rect 1846 1252 1847 1256
rect 1851 1252 1852 1256
rect 1846 1251 1852 1252
rect 1902 1256 1908 1257
rect 1902 1252 1903 1256
rect 1907 1252 1908 1256
rect 1902 1251 1908 1252
rect 1966 1256 1972 1257
rect 1966 1252 1967 1256
rect 1971 1252 1972 1256
rect 1966 1251 1972 1252
rect 2038 1256 2044 1257
rect 2038 1252 2039 1256
rect 2043 1252 2044 1256
rect 2038 1251 2044 1252
rect 2118 1256 2124 1257
rect 2118 1252 2119 1256
rect 2123 1252 2124 1256
rect 2118 1251 2124 1252
rect 2198 1256 2204 1257
rect 2198 1252 2199 1256
rect 2203 1252 2204 1256
rect 2198 1251 2204 1252
rect 2286 1256 2292 1257
rect 2286 1252 2287 1256
rect 2291 1252 2292 1256
rect 2286 1251 2292 1252
rect 2358 1256 2364 1257
rect 2358 1252 2359 1256
rect 2363 1252 2364 1256
rect 2358 1251 2364 1252
rect 998 1247 1004 1248
rect 134 1236 140 1237
rect 134 1232 135 1236
rect 139 1232 140 1236
rect 134 1231 140 1232
rect 174 1236 180 1237
rect 174 1232 175 1236
rect 179 1232 180 1236
rect 174 1231 180 1232
rect 230 1236 236 1237
rect 230 1232 231 1236
rect 235 1232 236 1236
rect 230 1231 236 1232
rect 310 1236 316 1237
rect 310 1232 311 1236
rect 315 1232 316 1236
rect 310 1231 316 1232
rect 398 1236 404 1237
rect 398 1232 399 1236
rect 403 1232 404 1236
rect 398 1231 404 1232
rect 486 1236 492 1237
rect 486 1232 487 1236
rect 491 1232 492 1236
rect 486 1231 492 1232
rect 574 1236 580 1237
rect 574 1232 575 1236
rect 579 1232 580 1236
rect 574 1231 580 1232
rect 662 1236 668 1237
rect 662 1232 663 1236
rect 667 1232 668 1236
rect 662 1231 668 1232
rect 742 1236 748 1237
rect 742 1232 743 1236
rect 747 1232 748 1236
rect 742 1231 748 1232
rect 814 1236 820 1237
rect 814 1232 815 1236
rect 819 1232 820 1236
rect 814 1231 820 1232
rect 878 1236 884 1237
rect 878 1232 879 1236
rect 883 1232 884 1236
rect 878 1231 884 1232
rect 942 1236 948 1237
rect 942 1232 943 1236
rect 947 1232 948 1236
rect 942 1231 948 1232
rect 1006 1236 1012 1237
rect 1006 1232 1007 1236
rect 1011 1232 1012 1236
rect 1006 1231 1012 1232
rect 1070 1236 1076 1237
rect 1070 1232 1071 1236
rect 1075 1232 1076 1236
rect 1070 1231 1076 1232
rect 1302 1236 1308 1237
rect 1302 1232 1303 1236
rect 1307 1232 1308 1236
rect 1302 1231 1308 1232
rect 1374 1236 1380 1237
rect 1374 1232 1375 1236
rect 1379 1232 1380 1236
rect 1374 1231 1380 1232
rect 1478 1236 1484 1237
rect 1478 1232 1479 1236
rect 1483 1232 1484 1236
rect 1478 1231 1484 1232
rect 1582 1236 1588 1237
rect 1582 1232 1583 1236
rect 1587 1232 1588 1236
rect 1582 1231 1588 1232
rect 1686 1236 1692 1237
rect 1686 1232 1687 1236
rect 1691 1232 1692 1236
rect 1686 1231 1692 1232
rect 1790 1236 1796 1237
rect 1790 1232 1791 1236
rect 1795 1232 1796 1236
rect 1790 1231 1796 1232
rect 1886 1236 1892 1237
rect 1886 1232 1887 1236
rect 1891 1232 1892 1236
rect 1886 1231 1892 1232
rect 1982 1236 1988 1237
rect 1982 1232 1983 1236
rect 1987 1232 1988 1236
rect 1982 1231 1988 1232
rect 2070 1236 2076 1237
rect 2070 1232 2071 1236
rect 2075 1232 2076 1236
rect 2070 1231 2076 1232
rect 2150 1236 2156 1237
rect 2150 1232 2151 1236
rect 2155 1232 2156 1236
rect 2150 1231 2156 1232
rect 2222 1236 2228 1237
rect 2222 1232 2223 1236
rect 2227 1232 2228 1236
rect 2222 1231 2228 1232
rect 2302 1236 2308 1237
rect 2302 1232 2303 1236
rect 2307 1232 2308 1236
rect 2302 1231 2308 1232
rect 2358 1236 2364 1237
rect 2358 1232 2359 1236
rect 2363 1232 2364 1236
rect 2358 1231 2364 1232
rect 110 1229 116 1230
rect 110 1225 111 1229
rect 115 1225 116 1229
rect 110 1224 116 1225
rect 1238 1229 1244 1230
rect 1238 1225 1239 1229
rect 1243 1225 1244 1229
rect 1238 1224 1244 1225
rect 1278 1229 1284 1230
rect 1278 1225 1279 1229
rect 1283 1225 1284 1229
rect 1278 1224 1284 1225
rect 2406 1229 2412 1230
rect 2406 1225 2407 1229
rect 2411 1225 2412 1229
rect 2406 1224 2412 1225
rect 159 1215 168 1216
rect 110 1212 116 1213
rect 110 1208 111 1212
rect 115 1208 116 1212
rect 159 1211 160 1215
rect 167 1211 168 1215
rect 159 1210 168 1211
rect 199 1215 205 1216
rect 199 1211 200 1215
rect 204 1214 205 1215
rect 222 1215 228 1216
rect 222 1214 223 1215
rect 204 1212 223 1214
rect 204 1211 205 1212
rect 199 1210 205 1211
rect 222 1211 223 1212
rect 227 1211 228 1215
rect 222 1210 228 1211
rect 254 1215 261 1216
rect 254 1211 255 1215
rect 260 1211 261 1215
rect 254 1210 261 1211
rect 263 1215 269 1216
rect 263 1211 264 1215
rect 268 1214 269 1215
rect 335 1215 341 1216
rect 335 1214 336 1215
rect 268 1212 336 1214
rect 268 1211 269 1212
rect 263 1210 269 1211
rect 335 1211 336 1212
rect 340 1211 341 1215
rect 335 1210 341 1211
rect 343 1215 349 1216
rect 343 1211 344 1215
rect 348 1214 349 1215
rect 423 1215 429 1216
rect 423 1214 424 1215
rect 348 1212 424 1214
rect 348 1211 349 1212
rect 343 1210 349 1211
rect 423 1211 424 1212
rect 428 1211 429 1215
rect 423 1210 429 1211
rect 431 1215 437 1216
rect 431 1211 432 1215
rect 436 1214 437 1215
rect 511 1215 517 1216
rect 511 1214 512 1215
rect 436 1212 512 1214
rect 436 1211 437 1212
rect 431 1210 437 1211
rect 511 1211 512 1212
rect 516 1211 517 1215
rect 511 1210 517 1211
rect 519 1215 525 1216
rect 519 1211 520 1215
rect 524 1214 525 1215
rect 599 1215 605 1216
rect 599 1214 600 1215
rect 524 1212 600 1214
rect 524 1211 525 1212
rect 519 1210 525 1211
rect 599 1211 600 1212
rect 604 1211 605 1215
rect 599 1210 605 1211
rect 654 1215 660 1216
rect 654 1211 655 1215
rect 659 1214 660 1215
rect 687 1215 693 1216
rect 687 1214 688 1215
rect 659 1212 688 1214
rect 659 1211 660 1212
rect 654 1210 660 1211
rect 687 1211 688 1212
rect 692 1211 693 1215
rect 687 1210 693 1211
rect 710 1215 716 1216
rect 710 1211 711 1215
rect 715 1214 716 1215
rect 767 1215 773 1216
rect 767 1214 768 1215
rect 715 1212 768 1214
rect 715 1211 716 1212
rect 710 1210 716 1211
rect 767 1211 768 1212
rect 772 1211 773 1215
rect 767 1210 773 1211
rect 775 1215 781 1216
rect 775 1211 776 1215
rect 780 1214 781 1215
rect 839 1215 845 1216
rect 839 1214 840 1215
rect 780 1212 840 1214
rect 780 1211 781 1212
rect 775 1210 781 1211
rect 839 1211 840 1212
rect 844 1211 845 1215
rect 839 1210 845 1211
rect 847 1215 853 1216
rect 847 1211 848 1215
rect 852 1214 853 1215
rect 903 1215 909 1216
rect 903 1214 904 1215
rect 852 1212 904 1214
rect 852 1211 853 1212
rect 847 1210 853 1211
rect 903 1211 904 1212
rect 908 1211 909 1215
rect 903 1210 909 1211
rect 911 1215 917 1216
rect 911 1211 912 1215
rect 916 1214 917 1215
rect 967 1215 973 1216
rect 967 1214 968 1215
rect 916 1212 968 1214
rect 916 1211 917 1212
rect 911 1210 917 1211
rect 967 1211 968 1212
rect 972 1211 973 1215
rect 967 1210 973 1211
rect 975 1215 981 1216
rect 975 1211 976 1215
rect 980 1214 981 1215
rect 1031 1215 1037 1216
rect 1031 1214 1032 1215
rect 980 1212 1032 1214
rect 980 1211 981 1212
rect 975 1210 981 1211
rect 1031 1211 1032 1212
rect 1036 1211 1037 1215
rect 1031 1210 1037 1211
rect 1039 1215 1045 1216
rect 1039 1211 1040 1215
rect 1044 1214 1045 1215
rect 1095 1215 1101 1216
rect 1095 1214 1096 1215
rect 1044 1212 1096 1214
rect 1044 1211 1045 1212
rect 1039 1210 1045 1211
rect 1095 1211 1096 1212
rect 1100 1211 1101 1215
rect 1310 1215 1316 1216
rect 1095 1210 1101 1211
rect 1238 1212 1244 1213
rect 110 1207 116 1208
rect 1238 1208 1239 1212
rect 1243 1208 1244 1212
rect 1238 1207 1244 1208
rect 1278 1212 1284 1213
rect 1278 1208 1279 1212
rect 1283 1208 1284 1212
rect 1310 1211 1311 1215
rect 1315 1214 1316 1215
rect 1327 1215 1333 1216
rect 1327 1214 1328 1215
rect 1315 1212 1328 1214
rect 1315 1211 1316 1212
rect 1310 1210 1316 1211
rect 1327 1211 1328 1212
rect 1332 1211 1333 1215
rect 1327 1210 1333 1211
rect 1335 1215 1341 1216
rect 1335 1211 1336 1215
rect 1340 1214 1341 1215
rect 1399 1215 1405 1216
rect 1399 1214 1400 1215
rect 1340 1212 1400 1214
rect 1340 1211 1341 1212
rect 1335 1210 1341 1211
rect 1399 1211 1400 1212
rect 1404 1211 1405 1215
rect 1399 1210 1405 1211
rect 1407 1215 1413 1216
rect 1407 1211 1408 1215
rect 1412 1214 1413 1215
rect 1503 1215 1509 1216
rect 1503 1214 1504 1215
rect 1412 1212 1504 1214
rect 1412 1211 1413 1212
rect 1407 1210 1413 1211
rect 1503 1211 1504 1212
rect 1508 1211 1509 1215
rect 1503 1210 1509 1211
rect 1607 1215 1613 1216
rect 1607 1211 1608 1215
rect 1612 1214 1613 1215
rect 1678 1215 1684 1216
rect 1678 1214 1679 1215
rect 1612 1212 1679 1214
rect 1612 1211 1613 1212
rect 1607 1210 1613 1211
rect 1678 1211 1679 1212
rect 1683 1211 1684 1215
rect 1711 1215 1717 1216
rect 1711 1214 1712 1215
rect 1678 1210 1684 1211
rect 1688 1212 1712 1214
rect 1278 1207 1284 1208
rect 1494 1207 1500 1208
rect 1494 1203 1495 1207
rect 1499 1206 1500 1207
rect 1688 1206 1690 1212
rect 1711 1211 1712 1212
rect 1716 1211 1717 1215
rect 1711 1210 1717 1211
rect 1815 1215 1821 1216
rect 1815 1211 1816 1215
rect 1820 1214 1821 1215
rect 1878 1215 1884 1216
rect 1878 1214 1879 1215
rect 1820 1212 1879 1214
rect 1820 1211 1821 1212
rect 1815 1210 1821 1211
rect 1878 1211 1879 1212
rect 1883 1211 1884 1215
rect 1878 1210 1884 1211
rect 1911 1215 1917 1216
rect 1911 1211 1912 1215
rect 1916 1214 1917 1215
rect 1974 1215 1980 1216
rect 1974 1214 1975 1215
rect 1916 1212 1975 1214
rect 1916 1211 1917 1212
rect 1911 1210 1917 1211
rect 1974 1211 1975 1212
rect 1979 1211 1980 1215
rect 1974 1210 1980 1211
rect 2007 1215 2013 1216
rect 2007 1211 2008 1215
rect 2012 1214 2013 1215
rect 2062 1215 2068 1216
rect 2062 1214 2063 1215
rect 2012 1212 2063 1214
rect 2012 1211 2013 1212
rect 2007 1210 2013 1211
rect 2062 1211 2063 1212
rect 2067 1211 2068 1215
rect 2062 1210 2068 1211
rect 2095 1215 2101 1216
rect 2095 1211 2096 1215
rect 2100 1214 2101 1215
rect 2142 1215 2148 1216
rect 2142 1214 2143 1215
rect 2100 1212 2143 1214
rect 2100 1211 2101 1212
rect 2095 1210 2101 1211
rect 2142 1211 2143 1212
rect 2147 1211 2148 1215
rect 2175 1215 2181 1216
rect 2175 1214 2176 1215
rect 2142 1210 2148 1211
rect 2152 1212 2176 1214
rect 1499 1204 1690 1206
rect 1910 1207 1916 1208
rect 1499 1203 1500 1204
rect 1494 1202 1500 1203
rect 1910 1203 1911 1207
rect 1915 1206 1916 1207
rect 2152 1206 2154 1212
rect 2175 1211 2176 1212
rect 2180 1211 2181 1215
rect 2175 1210 2181 1211
rect 2247 1215 2256 1216
rect 2247 1211 2248 1215
rect 2255 1211 2256 1215
rect 2247 1210 2256 1211
rect 2327 1215 2333 1216
rect 2327 1211 2328 1215
rect 2332 1214 2333 1215
rect 2350 1215 2356 1216
rect 2350 1214 2351 1215
rect 2332 1212 2351 1214
rect 2332 1211 2333 1212
rect 2327 1210 2333 1211
rect 2350 1211 2351 1212
rect 2355 1211 2356 1215
rect 2383 1215 2389 1216
rect 2383 1214 2384 1215
rect 2350 1210 2356 1211
rect 2360 1212 2384 1214
rect 1915 1204 2154 1206
rect 2310 1207 2316 1208
rect 1915 1203 1916 1204
rect 1910 1202 1916 1203
rect 2310 1203 2311 1207
rect 2315 1206 2316 1207
rect 2360 1206 2362 1212
rect 2383 1211 2384 1212
rect 2388 1211 2389 1215
rect 2383 1210 2389 1211
rect 2406 1212 2412 1213
rect 2406 1208 2407 1212
rect 2411 1208 2412 1212
rect 2406 1207 2412 1208
rect 2315 1204 2362 1206
rect 2315 1203 2316 1204
rect 2310 1202 2316 1203
rect 134 1189 140 1190
rect 134 1185 135 1189
rect 139 1185 140 1189
rect 134 1184 140 1185
rect 174 1189 180 1190
rect 174 1185 175 1189
rect 179 1185 180 1189
rect 174 1184 180 1185
rect 230 1189 236 1190
rect 230 1185 231 1189
rect 235 1185 236 1189
rect 230 1184 236 1185
rect 310 1189 316 1190
rect 310 1185 311 1189
rect 315 1185 316 1189
rect 310 1184 316 1185
rect 398 1189 404 1190
rect 398 1185 399 1189
rect 403 1185 404 1189
rect 398 1184 404 1185
rect 486 1189 492 1190
rect 486 1185 487 1189
rect 491 1185 492 1189
rect 486 1184 492 1185
rect 574 1189 580 1190
rect 574 1185 575 1189
rect 579 1185 580 1189
rect 574 1184 580 1185
rect 662 1189 668 1190
rect 662 1185 663 1189
rect 667 1185 668 1189
rect 662 1184 668 1185
rect 742 1189 748 1190
rect 742 1185 743 1189
rect 747 1185 748 1189
rect 742 1184 748 1185
rect 814 1189 820 1190
rect 814 1185 815 1189
rect 819 1185 820 1189
rect 814 1184 820 1185
rect 878 1189 884 1190
rect 878 1185 879 1189
rect 883 1185 884 1189
rect 878 1184 884 1185
rect 942 1189 948 1190
rect 942 1185 943 1189
rect 947 1185 948 1189
rect 942 1184 948 1185
rect 1006 1189 1012 1190
rect 1006 1185 1007 1189
rect 1011 1185 1012 1189
rect 1006 1184 1012 1185
rect 1070 1189 1076 1190
rect 1070 1185 1071 1189
rect 1075 1185 1076 1189
rect 1070 1184 1076 1185
rect 1302 1189 1308 1190
rect 1302 1185 1303 1189
rect 1307 1185 1308 1189
rect 1302 1184 1308 1185
rect 1374 1189 1380 1190
rect 1374 1185 1375 1189
rect 1379 1185 1380 1189
rect 1374 1184 1380 1185
rect 1478 1189 1484 1190
rect 1478 1185 1479 1189
rect 1483 1185 1484 1189
rect 1478 1184 1484 1185
rect 1582 1189 1588 1190
rect 1582 1185 1583 1189
rect 1587 1185 1588 1189
rect 1582 1184 1588 1185
rect 1686 1189 1692 1190
rect 1686 1185 1687 1189
rect 1691 1185 1692 1189
rect 1686 1184 1692 1185
rect 1790 1189 1796 1190
rect 1790 1185 1791 1189
rect 1795 1185 1796 1189
rect 1790 1184 1796 1185
rect 1886 1189 1892 1190
rect 1886 1185 1887 1189
rect 1891 1185 1892 1189
rect 1886 1184 1892 1185
rect 1982 1189 1988 1190
rect 1982 1185 1983 1189
rect 1987 1185 1988 1189
rect 1982 1184 1988 1185
rect 2070 1189 2076 1190
rect 2070 1185 2071 1189
rect 2075 1185 2076 1189
rect 2070 1184 2076 1185
rect 2150 1189 2156 1190
rect 2150 1185 2151 1189
rect 2155 1185 2156 1189
rect 2150 1184 2156 1185
rect 2222 1189 2228 1190
rect 2222 1185 2223 1189
rect 2227 1185 2228 1189
rect 2222 1184 2228 1185
rect 2302 1189 2308 1190
rect 2302 1185 2303 1189
rect 2307 1185 2308 1189
rect 2302 1184 2308 1185
rect 2358 1189 2364 1190
rect 2358 1185 2359 1189
rect 2363 1185 2364 1189
rect 2358 1184 2364 1185
rect 131 1179 137 1180
rect 131 1175 132 1179
rect 136 1178 137 1179
rect 154 1179 160 1180
rect 154 1178 155 1179
rect 136 1176 155 1178
rect 136 1175 137 1176
rect 131 1174 137 1175
rect 154 1175 155 1176
rect 159 1175 160 1179
rect 154 1174 160 1175
rect 162 1179 168 1180
rect 162 1175 163 1179
rect 167 1178 168 1179
rect 171 1179 177 1180
rect 171 1178 172 1179
rect 167 1176 172 1178
rect 167 1175 168 1176
rect 162 1174 168 1175
rect 171 1175 172 1176
rect 176 1175 177 1179
rect 171 1174 177 1175
rect 222 1179 233 1180
rect 222 1175 223 1179
rect 227 1175 228 1179
rect 232 1175 233 1179
rect 222 1174 233 1175
rect 307 1179 313 1180
rect 307 1175 308 1179
rect 312 1178 313 1179
rect 343 1179 349 1180
rect 343 1178 344 1179
rect 312 1176 344 1178
rect 312 1175 313 1176
rect 307 1174 313 1175
rect 343 1175 344 1176
rect 348 1175 349 1179
rect 343 1174 349 1175
rect 395 1179 401 1180
rect 395 1175 396 1179
rect 400 1178 401 1179
rect 431 1179 437 1180
rect 431 1178 432 1179
rect 400 1176 432 1178
rect 400 1175 401 1176
rect 395 1174 401 1175
rect 431 1175 432 1176
rect 436 1175 437 1179
rect 431 1174 437 1175
rect 483 1179 489 1180
rect 483 1175 484 1179
rect 488 1178 489 1179
rect 519 1179 525 1180
rect 519 1178 520 1179
rect 488 1176 520 1178
rect 488 1175 489 1176
rect 483 1174 489 1175
rect 519 1175 520 1176
rect 524 1175 525 1179
rect 519 1174 525 1175
rect 571 1179 577 1180
rect 571 1175 572 1179
rect 576 1178 577 1179
rect 582 1179 588 1180
rect 582 1178 583 1179
rect 576 1176 583 1178
rect 576 1175 577 1176
rect 571 1174 577 1175
rect 582 1175 583 1176
rect 587 1175 588 1179
rect 582 1174 588 1175
rect 659 1179 665 1180
rect 659 1175 660 1179
rect 664 1178 665 1179
rect 710 1179 716 1180
rect 710 1178 711 1179
rect 664 1176 711 1178
rect 664 1175 665 1176
rect 659 1174 665 1175
rect 710 1175 711 1176
rect 715 1175 716 1179
rect 710 1174 716 1175
rect 739 1179 745 1180
rect 739 1175 740 1179
rect 744 1178 745 1179
rect 775 1179 781 1180
rect 775 1178 776 1179
rect 744 1176 776 1178
rect 744 1175 745 1176
rect 739 1174 745 1175
rect 775 1175 776 1176
rect 780 1175 781 1179
rect 775 1174 781 1175
rect 811 1179 817 1180
rect 811 1175 812 1179
rect 816 1178 817 1179
rect 847 1179 853 1180
rect 847 1178 848 1179
rect 816 1176 848 1178
rect 816 1175 817 1176
rect 811 1174 817 1175
rect 847 1175 848 1176
rect 852 1175 853 1179
rect 847 1174 853 1175
rect 875 1179 881 1180
rect 875 1175 876 1179
rect 880 1178 881 1179
rect 911 1179 917 1180
rect 911 1178 912 1179
rect 880 1176 912 1178
rect 880 1175 881 1176
rect 875 1174 881 1175
rect 911 1175 912 1176
rect 916 1175 917 1179
rect 911 1174 917 1175
rect 939 1179 945 1180
rect 939 1175 940 1179
rect 944 1178 945 1179
rect 975 1179 981 1180
rect 975 1178 976 1179
rect 944 1176 976 1178
rect 944 1175 945 1176
rect 939 1174 945 1175
rect 975 1175 976 1176
rect 980 1175 981 1179
rect 975 1174 981 1175
rect 1003 1179 1009 1180
rect 1003 1175 1004 1179
rect 1008 1178 1009 1179
rect 1039 1179 1045 1180
rect 1039 1178 1040 1179
rect 1008 1176 1040 1178
rect 1008 1175 1009 1176
rect 1003 1174 1009 1175
rect 1039 1175 1040 1176
rect 1044 1175 1045 1179
rect 1039 1174 1045 1175
rect 1067 1179 1073 1180
rect 1067 1175 1068 1179
rect 1072 1178 1073 1179
rect 1214 1179 1220 1180
rect 1214 1178 1215 1179
rect 1072 1176 1215 1178
rect 1072 1175 1073 1176
rect 1067 1174 1073 1175
rect 1214 1175 1215 1176
rect 1219 1175 1220 1179
rect 1214 1174 1220 1175
rect 1299 1179 1305 1180
rect 1299 1175 1300 1179
rect 1304 1178 1305 1179
rect 1335 1179 1341 1180
rect 1335 1178 1336 1179
rect 1304 1176 1336 1178
rect 1304 1175 1305 1176
rect 1299 1174 1305 1175
rect 1335 1175 1336 1176
rect 1340 1175 1341 1179
rect 1335 1174 1341 1175
rect 1371 1179 1377 1180
rect 1371 1175 1372 1179
rect 1376 1178 1377 1179
rect 1407 1179 1413 1180
rect 1407 1178 1408 1179
rect 1376 1176 1408 1178
rect 1376 1175 1377 1176
rect 1371 1174 1377 1175
rect 1407 1175 1408 1176
rect 1412 1175 1413 1179
rect 1407 1174 1413 1175
rect 1475 1179 1481 1180
rect 1475 1175 1476 1179
rect 1480 1178 1481 1179
rect 1494 1179 1500 1180
rect 1494 1178 1495 1179
rect 1480 1176 1495 1178
rect 1480 1175 1481 1176
rect 1475 1174 1481 1175
rect 1494 1175 1495 1176
rect 1499 1175 1500 1179
rect 1494 1174 1500 1175
rect 1570 1179 1576 1180
rect 1570 1175 1571 1179
rect 1575 1178 1576 1179
rect 1579 1179 1585 1180
rect 1579 1178 1580 1179
rect 1575 1176 1580 1178
rect 1575 1175 1576 1176
rect 1570 1174 1576 1175
rect 1579 1175 1580 1176
rect 1584 1175 1585 1179
rect 1579 1174 1585 1175
rect 1678 1179 1689 1180
rect 1678 1175 1679 1179
rect 1683 1175 1684 1179
rect 1688 1175 1689 1179
rect 1678 1174 1689 1175
rect 1787 1179 1793 1180
rect 1787 1175 1788 1179
rect 1792 1178 1793 1179
rect 1806 1179 1812 1180
rect 1806 1178 1807 1179
rect 1792 1176 1807 1178
rect 1792 1175 1793 1176
rect 1787 1174 1793 1175
rect 1806 1175 1807 1176
rect 1811 1175 1812 1179
rect 1806 1174 1812 1175
rect 1878 1179 1889 1180
rect 1878 1175 1879 1179
rect 1883 1175 1884 1179
rect 1888 1175 1889 1179
rect 1878 1174 1889 1175
rect 1974 1179 1985 1180
rect 1974 1175 1975 1179
rect 1979 1175 1980 1179
rect 1984 1175 1985 1179
rect 1974 1174 1985 1175
rect 2062 1179 2073 1180
rect 2062 1175 2063 1179
rect 2067 1175 2068 1179
rect 2072 1175 2073 1179
rect 2062 1174 2073 1175
rect 2142 1179 2153 1180
rect 2142 1175 2143 1179
rect 2147 1175 2148 1179
rect 2152 1175 2153 1179
rect 2142 1174 2153 1175
rect 2186 1179 2192 1180
rect 2186 1175 2187 1179
rect 2191 1178 2192 1179
rect 2219 1179 2225 1180
rect 2219 1178 2220 1179
rect 2191 1176 2220 1178
rect 2191 1175 2192 1176
rect 2186 1174 2192 1175
rect 2219 1175 2220 1176
rect 2224 1175 2225 1179
rect 2219 1174 2225 1175
rect 2299 1179 2305 1180
rect 2299 1175 2300 1179
rect 2304 1178 2305 1179
rect 2310 1179 2316 1180
rect 2310 1178 2311 1179
rect 2304 1176 2311 1178
rect 2304 1175 2305 1176
rect 2299 1174 2305 1175
rect 2310 1175 2311 1176
rect 2315 1175 2316 1179
rect 2310 1174 2316 1175
rect 2355 1179 2361 1180
rect 2355 1175 2356 1179
rect 2360 1178 2361 1179
rect 2366 1179 2372 1180
rect 2366 1178 2367 1179
rect 2360 1176 2367 1178
rect 2360 1175 2361 1176
rect 2355 1174 2361 1175
rect 2366 1175 2367 1176
rect 2371 1175 2372 1179
rect 2366 1174 2372 1175
rect 263 1171 269 1172
rect 263 1170 264 1171
rect 235 1169 264 1170
rect 131 1167 137 1168
rect 131 1163 132 1167
rect 136 1166 137 1167
rect 146 1167 152 1168
rect 146 1166 147 1167
rect 136 1164 147 1166
rect 136 1163 137 1164
rect 131 1162 137 1163
rect 146 1163 147 1164
rect 151 1163 152 1167
rect 146 1162 152 1163
rect 162 1167 168 1168
rect 162 1163 163 1167
rect 167 1166 168 1167
rect 171 1167 177 1168
rect 171 1166 172 1167
rect 167 1164 172 1166
rect 167 1163 168 1164
rect 162 1162 168 1163
rect 171 1163 172 1164
rect 176 1163 177 1167
rect 235 1165 236 1169
rect 240 1168 264 1169
rect 240 1165 241 1168
rect 263 1167 264 1168
rect 268 1167 269 1171
rect 263 1166 269 1167
rect 271 1167 277 1168
rect 235 1164 241 1165
rect 171 1162 177 1163
rect 271 1163 272 1167
rect 276 1166 277 1167
rect 323 1167 329 1168
rect 323 1166 324 1167
rect 276 1164 324 1166
rect 276 1163 277 1164
rect 271 1162 277 1163
rect 323 1163 324 1164
rect 328 1163 329 1167
rect 323 1162 329 1163
rect 354 1167 360 1168
rect 354 1163 355 1167
rect 359 1166 360 1167
rect 427 1167 433 1168
rect 427 1166 428 1167
rect 359 1164 428 1166
rect 359 1163 360 1164
rect 354 1162 360 1163
rect 427 1163 428 1164
rect 432 1163 433 1167
rect 427 1162 433 1163
rect 458 1167 464 1168
rect 458 1163 459 1167
rect 463 1166 464 1167
rect 531 1167 537 1168
rect 531 1166 532 1167
rect 463 1164 532 1166
rect 463 1163 464 1164
rect 458 1162 464 1163
rect 531 1163 532 1164
rect 536 1163 537 1167
rect 531 1162 537 1163
rect 562 1167 568 1168
rect 562 1163 563 1167
rect 567 1166 568 1167
rect 635 1167 641 1168
rect 635 1166 636 1167
rect 567 1164 636 1166
rect 567 1163 568 1164
rect 562 1162 568 1163
rect 635 1163 636 1164
rect 640 1163 641 1167
rect 635 1162 641 1163
rect 739 1167 745 1168
rect 739 1163 740 1167
rect 744 1166 745 1167
rect 762 1167 768 1168
rect 762 1166 763 1167
rect 744 1164 763 1166
rect 744 1163 745 1164
rect 739 1162 745 1163
rect 762 1163 763 1164
rect 767 1163 768 1167
rect 762 1162 768 1163
rect 770 1167 776 1168
rect 770 1163 771 1167
rect 775 1166 776 1167
rect 835 1167 841 1168
rect 835 1166 836 1167
rect 775 1164 836 1166
rect 775 1163 776 1164
rect 770 1162 776 1163
rect 835 1163 836 1164
rect 840 1163 841 1167
rect 835 1162 841 1163
rect 866 1167 872 1168
rect 866 1163 867 1167
rect 871 1166 872 1167
rect 915 1167 921 1168
rect 915 1166 916 1167
rect 871 1164 916 1166
rect 871 1163 872 1164
rect 866 1162 872 1163
rect 915 1163 916 1164
rect 920 1163 921 1167
rect 915 1162 921 1163
rect 970 1167 976 1168
rect 970 1163 971 1167
rect 975 1166 976 1167
rect 995 1167 1001 1168
rect 995 1166 996 1167
rect 975 1164 996 1166
rect 975 1163 976 1164
rect 970 1162 976 1163
rect 995 1163 996 1164
rect 1000 1163 1001 1167
rect 995 1162 1001 1163
rect 1026 1167 1032 1168
rect 1026 1163 1027 1167
rect 1031 1166 1032 1167
rect 1067 1167 1073 1168
rect 1067 1166 1068 1167
rect 1031 1164 1068 1166
rect 1031 1163 1032 1164
rect 1026 1162 1032 1163
rect 1067 1163 1068 1164
rect 1072 1163 1073 1167
rect 1067 1162 1073 1163
rect 1098 1167 1104 1168
rect 1098 1163 1099 1167
rect 1103 1166 1104 1167
rect 1139 1167 1145 1168
rect 1139 1166 1140 1167
rect 1103 1164 1140 1166
rect 1103 1163 1104 1164
rect 1098 1162 1104 1163
rect 1139 1163 1140 1164
rect 1144 1163 1145 1167
rect 1139 1162 1145 1163
rect 1170 1167 1176 1168
rect 1170 1163 1171 1167
rect 1175 1166 1176 1167
rect 1187 1167 1193 1168
rect 1187 1166 1188 1167
rect 1175 1164 1188 1166
rect 1175 1163 1176 1164
rect 1170 1162 1176 1163
rect 1187 1163 1188 1164
rect 1192 1163 1193 1167
rect 1187 1162 1193 1163
rect 1299 1167 1305 1168
rect 1299 1163 1300 1167
rect 1304 1166 1305 1167
rect 1310 1167 1316 1168
rect 1310 1166 1311 1167
rect 1304 1164 1311 1166
rect 1304 1163 1305 1164
rect 1299 1162 1305 1163
rect 1310 1163 1311 1164
rect 1315 1163 1316 1167
rect 1310 1162 1316 1163
rect 1330 1167 1336 1168
rect 1330 1163 1331 1167
rect 1335 1166 1336 1167
rect 1339 1167 1345 1168
rect 1339 1166 1340 1167
rect 1335 1164 1340 1166
rect 1335 1163 1336 1164
rect 1330 1162 1336 1163
rect 1339 1163 1340 1164
rect 1344 1163 1345 1167
rect 1339 1162 1345 1163
rect 1383 1167 1389 1168
rect 1383 1163 1384 1167
rect 1388 1166 1389 1167
rect 1403 1167 1409 1168
rect 1403 1166 1404 1167
rect 1388 1164 1404 1166
rect 1388 1163 1389 1164
rect 1383 1162 1389 1163
rect 1403 1163 1404 1164
rect 1408 1163 1409 1167
rect 1403 1162 1409 1163
rect 1434 1167 1440 1168
rect 1434 1163 1435 1167
rect 1439 1166 1440 1167
rect 1483 1167 1489 1168
rect 1483 1166 1484 1167
rect 1439 1164 1484 1166
rect 1439 1163 1440 1164
rect 1434 1162 1440 1163
rect 1483 1163 1484 1164
rect 1488 1163 1489 1167
rect 1483 1162 1489 1163
rect 1514 1167 1520 1168
rect 1514 1163 1515 1167
rect 1519 1166 1520 1167
rect 1579 1167 1585 1168
rect 1579 1166 1580 1167
rect 1519 1164 1580 1166
rect 1519 1163 1520 1164
rect 1514 1162 1520 1163
rect 1579 1163 1580 1164
rect 1584 1163 1585 1167
rect 1579 1162 1585 1163
rect 1610 1167 1616 1168
rect 1610 1163 1611 1167
rect 1615 1166 1616 1167
rect 1683 1167 1689 1168
rect 1683 1166 1684 1167
rect 1615 1164 1684 1166
rect 1615 1163 1616 1164
rect 1610 1162 1616 1163
rect 1683 1163 1684 1164
rect 1688 1163 1689 1167
rect 1683 1162 1689 1163
rect 1714 1167 1720 1168
rect 1714 1163 1715 1167
rect 1719 1166 1720 1167
rect 1795 1167 1801 1168
rect 1795 1166 1796 1167
rect 1719 1164 1796 1166
rect 1719 1163 1720 1164
rect 1714 1162 1720 1163
rect 1795 1163 1796 1164
rect 1800 1163 1801 1167
rect 1795 1162 1801 1163
rect 1899 1167 1905 1168
rect 1899 1163 1900 1167
rect 1904 1166 1905 1167
rect 1910 1167 1916 1168
rect 1910 1166 1911 1167
rect 1904 1164 1911 1166
rect 1904 1163 1905 1164
rect 1899 1162 1905 1163
rect 1910 1163 1911 1164
rect 1915 1163 1916 1167
rect 1910 1162 1916 1163
rect 1930 1167 1936 1168
rect 1930 1163 1931 1167
rect 1935 1166 1936 1167
rect 1995 1167 2001 1168
rect 1995 1166 1996 1167
rect 1935 1164 1996 1166
rect 1935 1163 1936 1164
rect 1930 1162 1936 1163
rect 1995 1163 1996 1164
rect 2000 1163 2001 1167
rect 1995 1162 2001 1163
rect 2026 1167 2032 1168
rect 2026 1163 2027 1167
rect 2031 1166 2032 1167
rect 2075 1167 2081 1168
rect 2075 1166 2076 1167
rect 2031 1164 2076 1166
rect 2031 1163 2032 1164
rect 2026 1162 2032 1163
rect 2075 1163 2076 1164
rect 2080 1163 2081 1167
rect 2075 1162 2081 1163
rect 2155 1167 2161 1168
rect 2155 1163 2156 1167
rect 2160 1166 2161 1167
rect 2215 1167 2221 1168
rect 2215 1166 2216 1167
rect 2160 1164 2216 1166
rect 2160 1163 2161 1164
rect 2155 1162 2161 1163
rect 2215 1163 2216 1164
rect 2220 1163 2221 1167
rect 2215 1162 2221 1163
rect 2227 1167 2233 1168
rect 2227 1163 2228 1167
rect 2232 1166 2233 1167
rect 2290 1167 2296 1168
rect 2290 1166 2291 1167
rect 2232 1164 2291 1166
rect 2232 1163 2233 1164
rect 2227 1162 2233 1163
rect 2290 1163 2291 1164
rect 2295 1163 2296 1167
rect 2290 1162 2296 1163
rect 2299 1167 2305 1168
rect 2299 1163 2300 1167
rect 2304 1166 2305 1167
rect 2342 1167 2348 1168
rect 2342 1166 2343 1167
rect 2304 1164 2343 1166
rect 2304 1163 2305 1164
rect 2299 1162 2305 1163
rect 2342 1163 2343 1164
rect 2347 1163 2348 1167
rect 2342 1162 2348 1163
rect 2350 1167 2361 1168
rect 2350 1163 2351 1167
rect 2355 1163 2356 1167
rect 2360 1163 2361 1167
rect 2350 1162 2361 1163
rect 134 1159 140 1160
rect 134 1155 135 1159
rect 139 1155 140 1159
rect 134 1154 140 1155
rect 174 1159 180 1160
rect 174 1155 175 1159
rect 179 1155 180 1159
rect 174 1154 180 1155
rect 238 1159 244 1160
rect 238 1155 239 1159
rect 243 1155 244 1159
rect 238 1154 244 1155
rect 326 1159 332 1160
rect 326 1155 327 1159
rect 331 1155 332 1159
rect 326 1154 332 1155
rect 430 1159 436 1160
rect 430 1155 431 1159
rect 435 1155 436 1159
rect 430 1154 436 1155
rect 534 1159 540 1160
rect 534 1155 535 1159
rect 539 1155 540 1159
rect 534 1154 540 1155
rect 638 1159 644 1160
rect 638 1155 639 1159
rect 643 1155 644 1159
rect 638 1154 644 1155
rect 742 1159 748 1160
rect 742 1155 743 1159
rect 747 1155 748 1159
rect 742 1154 748 1155
rect 838 1159 844 1160
rect 838 1155 839 1159
rect 843 1155 844 1159
rect 838 1154 844 1155
rect 918 1159 924 1160
rect 918 1155 919 1159
rect 923 1155 924 1159
rect 918 1154 924 1155
rect 998 1159 1004 1160
rect 998 1155 999 1159
rect 1003 1155 1004 1159
rect 998 1154 1004 1155
rect 1070 1159 1076 1160
rect 1070 1155 1071 1159
rect 1075 1155 1076 1159
rect 1070 1154 1076 1155
rect 1142 1159 1148 1160
rect 1142 1155 1143 1159
rect 1147 1155 1148 1159
rect 1142 1154 1148 1155
rect 1190 1159 1196 1160
rect 1190 1155 1191 1159
rect 1195 1155 1196 1159
rect 1190 1154 1196 1155
rect 1302 1159 1308 1160
rect 1302 1155 1303 1159
rect 1307 1155 1308 1159
rect 1302 1154 1308 1155
rect 1342 1159 1348 1160
rect 1342 1155 1343 1159
rect 1347 1155 1348 1159
rect 1342 1154 1348 1155
rect 1406 1159 1412 1160
rect 1406 1155 1407 1159
rect 1411 1155 1412 1159
rect 1406 1154 1412 1155
rect 1486 1159 1492 1160
rect 1486 1155 1487 1159
rect 1491 1155 1492 1159
rect 1486 1154 1492 1155
rect 1582 1159 1588 1160
rect 1582 1155 1583 1159
rect 1587 1155 1588 1159
rect 1582 1154 1588 1155
rect 1686 1159 1692 1160
rect 1686 1155 1687 1159
rect 1691 1155 1692 1159
rect 1686 1154 1692 1155
rect 1798 1159 1804 1160
rect 1798 1155 1799 1159
rect 1803 1155 1804 1159
rect 1798 1154 1804 1155
rect 1902 1159 1908 1160
rect 1902 1155 1903 1159
rect 1907 1155 1908 1159
rect 1902 1154 1908 1155
rect 1998 1159 2004 1160
rect 1998 1155 1999 1159
rect 2003 1155 2004 1159
rect 1998 1154 2004 1155
rect 2078 1159 2084 1160
rect 2078 1155 2079 1159
rect 2083 1155 2084 1159
rect 2078 1154 2084 1155
rect 2158 1159 2164 1160
rect 2158 1155 2159 1159
rect 2163 1155 2164 1159
rect 2158 1154 2164 1155
rect 2230 1159 2236 1160
rect 2230 1155 2231 1159
rect 2235 1155 2236 1159
rect 2230 1154 2236 1155
rect 2302 1159 2308 1160
rect 2302 1155 2303 1159
rect 2307 1155 2308 1159
rect 2302 1154 2308 1155
rect 2358 1159 2364 1160
rect 2358 1155 2359 1159
rect 2363 1155 2364 1159
rect 2358 1154 2364 1155
rect 146 1139 152 1140
rect 110 1136 116 1137
rect 110 1132 111 1136
rect 115 1132 116 1136
rect 146 1135 147 1139
rect 151 1138 152 1139
rect 151 1136 203 1138
rect 151 1135 152 1136
rect 146 1134 152 1135
rect 201 1132 203 1136
rect 1238 1136 1244 1137
rect 1238 1132 1239 1136
rect 1243 1132 1244 1136
rect 110 1131 116 1132
rect 154 1131 165 1132
rect 154 1127 155 1131
rect 159 1127 160 1131
rect 164 1127 165 1131
rect 154 1126 165 1127
rect 199 1131 205 1132
rect 199 1127 200 1131
rect 204 1127 205 1131
rect 199 1126 205 1127
rect 263 1131 269 1132
rect 263 1127 264 1131
rect 268 1130 269 1131
rect 271 1131 277 1132
rect 271 1130 272 1131
rect 268 1128 272 1130
rect 268 1127 269 1128
rect 263 1126 269 1127
rect 271 1127 272 1128
rect 276 1127 277 1131
rect 271 1126 277 1127
rect 351 1131 360 1132
rect 351 1127 352 1131
rect 359 1127 360 1131
rect 351 1126 360 1127
rect 455 1131 464 1132
rect 455 1127 456 1131
rect 463 1127 464 1131
rect 455 1126 464 1127
rect 559 1131 568 1132
rect 559 1127 560 1131
rect 567 1127 568 1131
rect 559 1126 568 1127
rect 663 1131 669 1132
rect 663 1127 664 1131
rect 668 1127 669 1131
rect 663 1126 669 1127
rect 767 1131 776 1132
rect 767 1127 768 1131
rect 775 1127 776 1131
rect 767 1126 776 1127
rect 863 1131 872 1132
rect 863 1127 864 1131
rect 871 1127 872 1131
rect 863 1126 872 1127
rect 943 1131 949 1132
rect 943 1127 944 1131
rect 948 1130 949 1131
rect 970 1131 976 1132
rect 970 1130 971 1131
rect 948 1128 971 1130
rect 948 1127 949 1128
rect 943 1126 949 1127
rect 970 1127 971 1128
rect 975 1127 976 1131
rect 970 1126 976 1127
rect 1023 1131 1032 1132
rect 1023 1127 1024 1131
rect 1031 1127 1032 1131
rect 1023 1126 1032 1127
rect 1095 1131 1104 1132
rect 1095 1127 1096 1131
rect 1103 1127 1104 1131
rect 1095 1126 1104 1127
rect 1167 1131 1176 1132
rect 1167 1127 1168 1131
rect 1175 1127 1176 1131
rect 1167 1126 1176 1127
rect 1214 1131 1221 1132
rect 1238 1131 1244 1132
rect 1278 1136 1284 1137
rect 1278 1132 1279 1136
rect 1283 1132 1284 1136
rect 2406 1136 2412 1137
rect 2406 1132 2407 1136
rect 2411 1132 2412 1136
rect 1278 1131 1284 1132
rect 1327 1131 1336 1132
rect 1214 1127 1215 1131
rect 1220 1127 1221 1131
rect 1214 1126 1221 1127
rect 1327 1127 1328 1131
rect 1335 1127 1336 1131
rect 1327 1126 1336 1127
rect 1367 1131 1373 1132
rect 1367 1127 1368 1131
rect 1372 1130 1373 1131
rect 1383 1131 1389 1132
rect 1383 1130 1384 1131
rect 1372 1128 1384 1130
rect 1372 1127 1373 1128
rect 1367 1126 1373 1127
rect 1383 1127 1384 1128
rect 1388 1127 1389 1131
rect 1383 1126 1389 1127
rect 1431 1131 1440 1132
rect 1431 1127 1432 1131
rect 1439 1127 1440 1131
rect 1431 1126 1440 1127
rect 1511 1131 1520 1132
rect 1511 1127 1512 1131
rect 1519 1127 1520 1131
rect 1511 1126 1520 1127
rect 1607 1131 1616 1132
rect 1607 1127 1608 1131
rect 1615 1127 1616 1131
rect 1607 1126 1616 1127
rect 1711 1131 1720 1132
rect 1711 1127 1712 1131
rect 1719 1127 1720 1131
rect 1711 1126 1720 1127
rect 1734 1131 1740 1132
rect 1734 1127 1735 1131
rect 1739 1130 1740 1131
rect 1823 1131 1829 1132
rect 1823 1130 1824 1131
rect 1739 1128 1824 1130
rect 1739 1127 1740 1128
rect 1734 1126 1740 1127
rect 1823 1127 1824 1128
rect 1828 1127 1829 1131
rect 1823 1126 1829 1127
rect 1927 1131 1936 1132
rect 1927 1127 1928 1131
rect 1935 1127 1936 1131
rect 1927 1126 1936 1127
rect 2023 1131 2032 1132
rect 2023 1127 2024 1131
rect 2031 1127 2032 1131
rect 2023 1126 2032 1127
rect 2103 1131 2109 1132
rect 2103 1127 2104 1131
rect 2108 1130 2109 1131
rect 2166 1131 2172 1132
rect 2166 1130 2167 1131
rect 2108 1128 2167 1130
rect 2108 1127 2109 1128
rect 2103 1126 2109 1127
rect 2166 1127 2167 1128
rect 2171 1127 2172 1131
rect 2166 1126 2172 1127
rect 2183 1131 2192 1132
rect 2183 1127 2184 1131
rect 2191 1127 2192 1131
rect 2183 1126 2192 1127
rect 2215 1131 2221 1132
rect 2215 1127 2216 1131
rect 2220 1130 2221 1131
rect 2255 1131 2261 1132
rect 2255 1130 2256 1131
rect 2220 1128 2256 1130
rect 2220 1127 2221 1128
rect 2215 1126 2221 1127
rect 2255 1127 2256 1128
rect 2260 1127 2261 1131
rect 2255 1126 2261 1127
rect 2290 1131 2296 1132
rect 2290 1127 2291 1131
rect 2295 1130 2296 1131
rect 2327 1131 2333 1132
rect 2327 1130 2328 1131
rect 2295 1128 2328 1130
rect 2295 1127 2296 1128
rect 2290 1126 2296 1127
rect 2327 1127 2328 1128
rect 2332 1127 2333 1131
rect 2327 1126 2333 1127
rect 2342 1131 2348 1132
rect 2342 1127 2343 1131
rect 2347 1130 2348 1131
rect 2383 1131 2389 1132
rect 2406 1131 2412 1132
rect 2383 1130 2384 1131
rect 2347 1128 2384 1130
rect 2347 1127 2348 1128
rect 2342 1126 2348 1127
rect 2383 1127 2384 1128
rect 2388 1127 2389 1131
rect 2383 1126 2389 1127
rect 346 1123 352 1124
rect 110 1119 116 1120
rect 110 1115 111 1119
rect 115 1115 116 1119
rect 346 1119 347 1123
rect 351 1122 352 1123
rect 665 1122 667 1126
rect 351 1120 667 1122
rect 351 1119 352 1120
rect 346 1118 352 1119
rect 1238 1119 1244 1120
rect 110 1114 116 1115
rect 1238 1115 1239 1119
rect 1243 1115 1244 1119
rect 1238 1114 1244 1115
rect 1278 1119 1284 1120
rect 1278 1115 1279 1119
rect 1283 1115 1284 1119
rect 1278 1114 1284 1115
rect 2406 1119 2412 1120
rect 2406 1115 2407 1119
rect 2411 1115 2412 1119
rect 2406 1114 2412 1115
rect 134 1112 140 1113
rect 134 1108 135 1112
rect 139 1108 140 1112
rect 134 1107 140 1108
rect 174 1112 180 1113
rect 174 1108 175 1112
rect 179 1108 180 1112
rect 174 1107 180 1108
rect 238 1112 244 1113
rect 238 1108 239 1112
rect 243 1108 244 1112
rect 238 1107 244 1108
rect 326 1112 332 1113
rect 326 1108 327 1112
rect 331 1108 332 1112
rect 326 1107 332 1108
rect 430 1112 436 1113
rect 430 1108 431 1112
rect 435 1108 436 1112
rect 430 1107 436 1108
rect 534 1112 540 1113
rect 534 1108 535 1112
rect 539 1108 540 1112
rect 534 1107 540 1108
rect 638 1112 644 1113
rect 638 1108 639 1112
rect 643 1108 644 1112
rect 638 1107 644 1108
rect 742 1112 748 1113
rect 742 1108 743 1112
rect 747 1108 748 1112
rect 742 1107 748 1108
rect 838 1112 844 1113
rect 838 1108 839 1112
rect 843 1108 844 1112
rect 838 1107 844 1108
rect 918 1112 924 1113
rect 918 1108 919 1112
rect 923 1108 924 1112
rect 918 1107 924 1108
rect 998 1112 1004 1113
rect 998 1108 999 1112
rect 1003 1108 1004 1112
rect 998 1107 1004 1108
rect 1070 1112 1076 1113
rect 1070 1108 1071 1112
rect 1075 1108 1076 1112
rect 1070 1107 1076 1108
rect 1142 1112 1148 1113
rect 1142 1108 1143 1112
rect 1147 1108 1148 1112
rect 1142 1107 1148 1108
rect 1190 1112 1196 1113
rect 1190 1108 1191 1112
rect 1195 1108 1196 1112
rect 1190 1107 1196 1108
rect 1302 1112 1308 1113
rect 1302 1108 1303 1112
rect 1307 1108 1308 1112
rect 1302 1107 1308 1108
rect 1342 1112 1348 1113
rect 1342 1108 1343 1112
rect 1347 1108 1348 1112
rect 1342 1107 1348 1108
rect 1406 1112 1412 1113
rect 1406 1108 1407 1112
rect 1411 1108 1412 1112
rect 1406 1107 1412 1108
rect 1486 1112 1492 1113
rect 1486 1108 1487 1112
rect 1491 1108 1492 1112
rect 1486 1107 1492 1108
rect 1582 1112 1588 1113
rect 1582 1108 1583 1112
rect 1587 1108 1588 1112
rect 1582 1107 1588 1108
rect 1686 1112 1692 1113
rect 1686 1108 1687 1112
rect 1691 1108 1692 1112
rect 1686 1107 1692 1108
rect 1798 1112 1804 1113
rect 1798 1108 1799 1112
rect 1803 1108 1804 1112
rect 1798 1107 1804 1108
rect 1902 1112 1908 1113
rect 1902 1108 1903 1112
rect 1907 1108 1908 1112
rect 1902 1107 1908 1108
rect 1998 1112 2004 1113
rect 1998 1108 1999 1112
rect 2003 1108 2004 1112
rect 1998 1107 2004 1108
rect 2078 1112 2084 1113
rect 2078 1108 2079 1112
rect 2083 1108 2084 1112
rect 2078 1107 2084 1108
rect 2158 1112 2164 1113
rect 2158 1108 2159 1112
rect 2163 1108 2164 1112
rect 2158 1107 2164 1108
rect 2230 1112 2236 1113
rect 2230 1108 2231 1112
rect 2235 1108 2236 1112
rect 2230 1107 2236 1108
rect 2302 1112 2308 1113
rect 2302 1108 2303 1112
rect 2307 1108 2308 1112
rect 2302 1107 2308 1108
rect 2358 1112 2364 1113
rect 2358 1108 2359 1112
rect 2363 1108 2364 1112
rect 2358 1107 2364 1108
rect 1430 1100 1436 1101
rect 134 1096 140 1097
rect 134 1092 135 1096
rect 139 1092 140 1096
rect 134 1091 140 1092
rect 174 1096 180 1097
rect 174 1092 175 1096
rect 179 1092 180 1096
rect 174 1091 180 1092
rect 246 1096 252 1097
rect 246 1092 247 1096
rect 251 1092 252 1096
rect 246 1091 252 1092
rect 326 1096 332 1097
rect 326 1092 327 1096
rect 331 1092 332 1096
rect 326 1091 332 1092
rect 414 1096 420 1097
rect 414 1092 415 1096
rect 419 1092 420 1096
rect 414 1091 420 1092
rect 502 1096 508 1097
rect 502 1092 503 1096
rect 507 1092 508 1096
rect 502 1091 508 1092
rect 582 1096 588 1097
rect 582 1092 583 1096
rect 587 1092 588 1096
rect 582 1091 588 1092
rect 662 1096 668 1097
rect 662 1092 663 1096
rect 667 1092 668 1096
rect 662 1091 668 1092
rect 734 1096 740 1097
rect 734 1092 735 1096
rect 739 1092 740 1096
rect 734 1091 740 1092
rect 798 1096 804 1097
rect 798 1092 799 1096
rect 803 1092 804 1096
rect 798 1091 804 1092
rect 862 1096 868 1097
rect 862 1092 863 1096
rect 867 1092 868 1096
rect 862 1091 868 1092
rect 918 1096 924 1097
rect 918 1092 919 1096
rect 923 1092 924 1096
rect 918 1091 924 1092
rect 982 1096 988 1097
rect 982 1092 983 1096
rect 987 1092 988 1096
rect 982 1091 988 1092
rect 1046 1096 1052 1097
rect 1046 1092 1047 1096
rect 1051 1092 1052 1096
rect 1430 1096 1431 1100
rect 1435 1096 1436 1100
rect 1430 1095 1436 1096
rect 1470 1100 1476 1101
rect 1470 1096 1471 1100
rect 1475 1096 1476 1100
rect 1470 1095 1476 1096
rect 1510 1100 1516 1101
rect 1510 1096 1511 1100
rect 1515 1096 1516 1100
rect 1510 1095 1516 1096
rect 1558 1100 1564 1101
rect 1558 1096 1559 1100
rect 1563 1096 1564 1100
rect 1558 1095 1564 1096
rect 1614 1100 1620 1101
rect 1614 1096 1615 1100
rect 1619 1096 1620 1100
rect 1614 1095 1620 1096
rect 1670 1100 1676 1101
rect 1670 1096 1671 1100
rect 1675 1096 1676 1100
rect 1670 1095 1676 1096
rect 1726 1100 1732 1101
rect 1726 1096 1727 1100
rect 1731 1096 1732 1100
rect 1726 1095 1732 1096
rect 1774 1100 1780 1101
rect 1774 1096 1775 1100
rect 1779 1096 1780 1100
rect 1774 1095 1780 1096
rect 1822 1100 1828 1101
rect 1822 1096 1823 1100
rect 1827 1096 1828 1100
rect 1822 1095 1828 1096
rect 1870 1100 1876 1101
rect 1870 1096 1871 1100
rect 1875 1096 1876 1100
rect 1870 1095 1876 1096
rect 1918 1100 1924 1101
rect 1918 1096 1919 1100
rect 1923 1096 1924 1100
rect 1918 1095 1924 1096
rect 1966 1100 1972 1101
rect 1966 1096 1967 1100
rect 1971 1096 1972 1100
rect 1966 1095 1972 1096
rect 2014 1100 2020 1101
rect 2014 1096 2015 1100
rect 2019 1096 2020 1100
rect 2014 1095 2020 1096
rect 2062 1100 2068 1101
rect 2062 1096 2063 1100
rect 2067 1096 2068 1100
rect 2062 1095 2068 1096
rect 2118 1100 2124 1101
rect 2118 1096 2119 1100
rect 2123 1096 2124 1100
rect 2118 1095 2124 1096
rect 2174 1100 2180 1101
rect 2174 1096 2175 1100
rect 2179 1096 2180 1100
rect 2174 1095 2180 1096
rect 2230 1100 2236 1101
rect 2230 1096 2231 1100
rect 2235 1096 2236 1100
rect 2230 1095 2236 1096
rect 1046 1091 1052 1092
rect 1278 1093 1284 1094
rect 110 1089 116 1090
rect 110 1085 111 1089
rect 115 1085 116 1089
rect 110 1084 116 1085
rect 1238 1089 1244 1090
rect 1238 1085 1239 1089
rect 1243 1085 1244 1089
rect 1278 1089 1279 1093
rect 1283 1089 1284 1093
rect 1278 1088 1284 1089
rect 2406 1093 2412 1094
rect 2406 1089 2407 1093
rect 2411 1089 2412 1093
rect 2406 1088 2412 1089
rect 1238 1084 1244 1085
rect 1455 1079 1464 1080
rect 1278 1076 1284 1077
rect 159 1075 168 1076
rect 110 1072 116 1073
rect 110 1068 111 1072
rect 115 1068 116 1072
rect 159 1071 160 1075
rect 167 1071 168 1075
rect 159 1070 168 1071
rect 199 1075 205 1076
rect 199 1071 200 1075
rect 204 1074 205 1075
rect 238 1075 244 1076
rect 238 1074 239 1075
rect 204 1072 239 1074
rect 204 1071 205 1072
rect 199 1070 205 1071
rect 238 1071 239 1072
rect 243 1071 244 1075
rect 271 1075 277 1076
rect 271 1074 272 1075
rect 238 1070 244 1071
rect 248 1072 272 1074
rect 110 1067 116 1068
rect 142 1067 148 1068
rect 142 1063 143 1067
rect 147 1066 148 1067
rect 248 1066 250 1072
rect 271 1071 272 1072
rect 276 1071 277 1075
rect 271 1070 277 1071
rect 351 1075 357 1076
rect 351 1071 352 1075
rect 356 1074 357 1075
rect 406 1075 412 1076
rect 406 1074 407 1075
rect 356 1072 407 1074
rect 356 1071 357 1072
rect 351 1070 357 1071
rect 406 1071 407 1072
rect 411 1071 412 1075
rect 406 1070 412 1071
rect 439 1075 445 1076
rect 439 1071 440 1075
rect 444 1074 445 1075
rect 494 1075 500 1076
rect 494 1074 495 1075
rect 444 1072 495 1074
rect 444 1071 445 1072
rect 439 1070 445 1071
rect 494 1071 495 1072
rect 499 1071 500 1075
rect 494 1070 500 1071
rect 527 1075 533 1076
rect 527 1071 528 1075
rect 532 1074 533 1075
rect 567 1075 573 1076
rect 567 1074 568 1075
rect 532 1072 568 1074
rect 532 1071 533 1072
rect 527 1070 533 1071
rect 567 1071 568 1072
rect 572 1071 573 1075
rect 607 1075 613 1076
rect 607 1074 608 1075
rect 567 1070 573 1071
rect 576 1072 608 1074
rect 147 1064 250 1066
rect 334 1067 340 1068
rect 147 1063 148 1064
rect 142 1062 148 1063
rect 334 1063 335 1067
rect 339 1066 340 1067
rect 576 1066 578 1072
rect 607 1071 608 1072
rect 612 1071 613 1075
rect 607 1070 613 1071
rect 687 1075 693 1076
rect 687 1071 688 1075
rect 692 1074 693 1075
rect 726 1075 732 1076
rect 726 1074 727 1075
rect 692 1072 727 1074
rect 692 1071 693 1072
rect 687 1070 693 1071
rect 726 1071 727 1072
rect 731 1071 732 1075
rect 726 1070 732 1071
rect 759 1075 765 1076
rect 759 1071 760 1075
rect 764 1074 765 1075
rect 790 1075 796 1076
rect 790 1074 791 1075
rect 764 1072 791 1074
rect 764 1071 765 1072
rect 759 1070 765 1071
rect 790 1071 791 1072
rect 795 1071 796 1075
rect 790 1070 796 1071
rect 823 1075 829 1076
rect 823 1071 824 1075
rect 828 1074 829 1075
rect 854 1075 860 1076
rect 854 1074 855 1075
rect 828 1072 855 1074
rect 828 1071 829 1072
rect 823 1070 829 1071
rect 854 1071 855 1072
rect 859 1071 860 1075
rect 854 1070 860 1071
rect 887 1075 893 1076
rect 887 1071 888 1075
rect 892 1074 893 1075
rect 910 1075 916 1076
rect 910 1074 911 1075
rect 892 1072 911 1074
rect 892 1071 893 1072
rect 887 1070 893 1071
rect 910 1071 911 1072
rect 915 1071 916 1075
rect 910 1070 916 1071
rect 943 1075 949 1076
rect 943 1071 944 1075
rect 948 1074 949 1075
rect 974 1075 980 1076
rect 974 1074 975 1075
rect 948 1072 975 1074
rect 948 1071 949 1072
rect 943 1070 949 1071
rect 974 1071 975 1072
rect 979 1071 980 1075
rect 974 1070 980 1071
rect 1007 1075 1013 1076
rect 1007 1071 1008 1075
rect 1012 1074 1013 1075
rect 1038 1075 1044 1076
rect 1038 1074 1039 1075
rect 1012 1072 1039 1074
rect 1012 1071 1013 1072
rect 1007 1070 1013 1071
rect 1038 1071 1039 1072
rect 1043 1071 1044 1075
rect 1038 1070 1044 1071
rect 1070 1075 1077 1076
rect 1070 1071 1071 1075
rect 1076 1071 1077 1075
rect 1070 1070 1077 1071
rect 1238 1072 1244 1073
rect 1238 1068 1239 1072
rect 1243 1068 1244 1072
rect 1278 1072 1279 1076
rect 1283 1072 1284 1076
rect 1455 1075 1456 1079
rect 1463 1075 1464 1079
rect 1455 1074 1464 1075
rect 1495 1079 1504 1080
rect 1495 1075 1496 1079
rect 1503 1075 1504 1079
rect 1495 1074 1504 1075
rect 1535 1079 1541 1080
rect 1535 1075 1536 1079
rect 1540 1078 1541 1079
rect 1550 1079 1556 1080
rect 1550 1078 1551 1079
rect 1540 1076 1551 1078
rect 1540 1075 1541 1076
rect 1535 1074 1541 1075
rect 1550 1075 1551 1076
rect 1555 1075 1556 1079
rect 1550 1074 1556 1075
rect 1583 1079 1589 1080
rect 1583 1075 1584 1079
rect 1588 1078 1589 1079
rect 1606 1079 1612 1080
rect 1606 1078 1607 1079
rect 1588 1076 1607 1078
rect 1588 1075 1589 1076
rect 1583 1074 1589 1075
rect 1606 1075 1607 1076
rect 1611 1075 1612 1079
rect 1606 1074 1612 1075
rect 1639 1079 1645 1080
rect 1639 1075 1640 1079
rect 1644 1078 1645 1079
rect 1662 1079 1668 1080
rect 1662 1078 1663 1079
rect 1644 1076 1663 1078
rect 1644 1075 1645 1076
rect 1639 1074 1645 1075
rect 1662 1075 1663 1076
rect 1667 1075 1668 1079
rect 1662 1074 1668 1075
rect 1695 1079 1701 1080
rect 1695 1075 1696 1079
rect 1700 1078 1701 1079
rect 1714 1079 1720 1080
rect 1714 1078 1715 1079
rect 1700 1076 1715 1078
rect 1700 1075 1701 1076
rect 1695 1074 1701 1075
rect 1714 1075 1715 1076
rect 1719 1075 1720 1079
rect 1751 1079 1757 1080
rect 1751 1078 1752 1079
rect 1714 1074 1720 1075
rect 1724 1076 1752 1078
rect 1278 1071 1284 1072
rect 1582 1071 1588 1072
rect 1238 1067 1244 1068
rect 1582 1067 1583 1071
rect 1587 1070 1588 1071
rect 1724 1070 1726 1076
rect 1751 1075 1752 1076
rect 1756 1075 1757 1079
rect 1751 1074 1757 1075
rect 1799 1079 1805 1080
rect 1799 1075 1800 1079
rect 1804 1078 1805 1079
rect 1814 1079 1820 1080
rect 1814 1078 1815 1079
rect 1804 1076 1815 1078
rect 1804 1075 1805 1076
rect 1799 1074 1805 1075
rect 1814 1075 1815 1076
rect 1819 1075 1820 1079
rect 1847 1079 1853 1080
rect 1847 1078 1848 1079
rect 1814 1074 1820 1075
rect 1824 1076 1848 1078
rect 1587 1068 1726 1070
rect 1782 1071 1788 1072
rect 1587 1067 1588 1068
rect 1582 1066 1588 1067
rect 1782 1067 1783 1071
rect 1787 1070 1788 1071
rect 1824 1070 1826 1076
rect 1847 1075 1848 1076
rect 1852 1075 1853 1079
rect 1847 1074 1853 1075
rect 1855 1079 1861 1080
rect 1855 1075 1856 1079
rect 1860 1078 1861 1079
rect 1895 1079 1901 1080
rect 1895 1078 1896 1079
rect 1860 1076 1896 1078
rect 1860 1075 1861 1076
rect 1855 1074 1861 1075
rect 1895 1075 1896 1076
rect 1900 1075 1901 1079
rect 1895 1074 1901 1075
rect 1903 1079 1909 1080
rect 1903 1075 1904 1079
rect 1908 1078 1909 1079
rect 1943 1079 1949 1080
rect 1943 1078 1944 1079
rect 1908 1076 1944 1078
rect 1908 1075 1909 1076
rect 1903 1074 1909 1075
rect 1943 1075 1944 1076
rect 1948 1075 1949 1079
rect 1943 1074 1949 1075
rect 1951 1079 1957 1080
rect 1951 1075 1952 1079
rect 1956 1078 1957 1079
rect 1991 1079 1997 1080
rect 1991 1078 1992 1079
rect 1956 1076 1992 1078
rect 1956 1075 1957 1076
rect 1951 1074 1957 1075
rect 1991 1075 1992 1076
rect 1996 1075 1997 1079
rect 1991 1074 1997 1075
rect 2002 1079 2008 1080
rect 2002 1075 2003 1079
rect 2007 1078 2008 1079
rect 2039 1079 2045 1080
rect 2039 1078 2040 1079
rect 2007 1076 2040 1078
rect 2007 1075 2008 1076
rect 2002 1074 2008 1075
rect 2039 1075 2040 1076
rect 2044 1075 2045 1079
rect 2039 1074 2045 1075
rect 2047 1079 2053 1080
rect 2047 1075 2048 1079
rect 2052 1078 2053 1079
rect 2087 1079 2093 1080
rect 2087 1078 2088 1079
rect 2052 1076 2088 1078
rect 2052 1075 2053 1076
rect 2047 1074 2053 1075
rect 2087 1075 2088 1076
rect 2092 1075 2093 1079
rect 2087 1074 2093 1075
rect 2095 1079 2101 1080
rect 2095 1075 2096 1079
rect 2100 1078 2101 1079
rect 2143 1079 2149 1080
rect 2143 1078 2144 1079
rect 2100 1076 2144 1078
rect 2100 1075 2101 1076
rect 2095 1074 2101 1075
rect 2143 1075 2144 1076
rect 2148 1075 2149 1079
rect 2143 1074 2149 1075
rect 2199 1079 2205 1080
rect 2199 1075 2200 1079
rect 2204 1078 2205 1079
rect 2222 1079 2228 1080
rect 2222 1078 2223 1079
rect 2204 1076 2223 1078
rect 2204 1075 2205 1076
rect 2199 1074 2205 1075
rect 2222 1075 2223 1076
rect 2227 1075 2228 1079
rect 2222 1074 2228 1075
rect 2246 1079 2252 1080
rect 2246 1075 2247 1079
rect 2251 1078 2252 1079
rect 2255 1079 2261 1080
rect 2255 1078 2256 1079
rect 2251 1076 2256 1078
rect 2251 1075 2252 1076
rect 2246 1074 2252 1075
rect 2255 1075 2256 1076
rect 2260 1075 2261 1079
rect 2255 1074 2261 1075
rect 2406 1076 2412 1077
rect 2406 1072 2407 1076
rect 2411 1072 2412 1076
rect 2406 1071 2412 1072
rect 1787 1068 1826 1070
rect 1787 1067 1788 1068
rect 1782 1066 1788 1067
rect 339 1064 578 1066
rect 339 1063 340 1064
rect 334 1062 340 1063
rect 1430 1053 1436 1054
rect 134 1049 140 1050
rect 134 1045 135 1049
rect 139 1045 140 1049
rect 134 1044 140 1045
rect 174 1049 180 1050
rect 174 1045 175 1049
rect 179 1045 180 1049
rect 174 1044 180 1045
rect 246 1049 252 1050
rect 246 1045 247 1049
rect 251 1045 252 1049
rect 246 1044 252 1045
rect 326 1049 332 1050
rect 326 1045 327 1049
rect 331 1045 332 1049
rect 326 1044 332 1045
rect 414 1049 420 1050
rect 414 1045 415 1049
rect 419 1045 420 1049
rect 414 1044 420 1045
rect 502 1049 508 1050
rect 502 1045 503 1049
rect 507 1045 508 1049
rect 502 1044 508 1045
rect 582 1049 588 1050
rect 582 1045 583 1049
rect 587 1045 588 1049
rect 582 1044 588 1045
rect 662 1049 668 1050
rect 662 1045 663 1049
rect 667 1045 668 1049
rect 662 1044 668 1045
rect 734 1049 740 1050
rect 734 1045 735 1049
rect 739 1045 740 1049
rect 734 1044 740 1045
rect 798 1049 804 1050
rect 798 1045 799 1049
rect 803 1045 804 1049
rect 798 1044 804 1045
rect 862 1049 868 1050
rect 862 1045 863 1049
rect 867 1045 868 1049
rect 862 1044 868 1045
rect 918 1049 924 1050
rect 918 1045 919 1049
rect 923 1045 924 1049
rect 918 1044 924 1045
rect 982 1049 988 1050
rect 982 1045 983 1049
rect 987 1045 988 1049
rect 982 1044 988 1045
rect 1046 1049 1052 1050
rect 1046 1045 1047 1049
rect 1051 1045 1052 1049
rect 1430 1049 1431 1053
rect 1435 1049 1436 1053
rect 1430 1048 1436 1049
rect 1470 1053 1476 1054
rect 1470 1049 1471 1053
rect 1475 1049 1476 1053
rect 1470 1048 1476 1049
rect 1510 1053 1516 1054
rect 1510 1049 1511 1053
rect 1515 1049 1516 1053
rect 1510 1048 1516 1049
rect 1558 1053 1564 1054
rect 1558 1049 1559 1053
rect 1563 1049 1564 1053
rect 1558 1048 1564 1049
rect 1614 1053 1620 1054
rect 1614 1049 1615 1053
rect 1619 1049 1620 1053
rect 1614 1048 1620 1049
rect 1670 1053 1676 1054
rect 1670 1049 1671 1053
rect 1675 1049 1676 1053
rect 1670 1048 1676 1049
rect 1726 1053 1732 1054
rect 1726 1049 1727 1053
rect 1731 1049 1732 1053
rect 1726 1048 1732 1049
rect 1774 1053 1780 1054
rect 1774 1049 1775 1053
rect 1779 1049 1780 1053
rect 1774 1048 1780 1049
rect 1822 1053 1828 1054
rect 1822 1049 1823 1053
rect 1827 1049 1828 1053
rect 1822 1048 1828 1049
rect 1870 1053 1876 1054
rect 1870 1049 1871 1053
rect 1875 1049 1876 1053
rect 1870 1048 1876 1049
rect 1918 1053 1924 1054
rect 1918 1049 1919 1053
rect 1923 1049 1924 1053
rect 1918 1048 1924 1049
rect 1966 1053 1972 1054
rect 1966 1049 1967 1053
rect 1971 1049 1972 1053
rect 1966 1048 1972 1049
rect 2014 1053 2020 1054
rect 2014 1049 2015 1053
rect 2019 1049 2020 1053
rect 2014 1048 2020 1049
rect 2062 1053 2068 1054
rect 2062 1049 2063 1053
rect 2067 1049 2068 1053
rect 2062 1048 2068 1049
rect 2118 1053 2124 1054
rect 2118 1049 2119 1053
rect 2123 1049 2124 1053
rect 2118 1048 2124 1049
rect 2174 1053 2180 1054
rect 2174 1049 2175 1053
rect 2179 1049 2180 1053
rect 2174 1048 2180 1049
rect 2230 1053 2236 1054
rect 2230 1049 2231 1053
rect 2235 1049 2236 1053
rect 2230 1048 2236 1049
rect 1046 1044 1052 1045
rect 1427 1043 1433 1044
rect 131 1039 137 1040
rect 131 1035 132 1039
rect 136 1038 137 1039
rect 142 1039 148 1040
rect 142 1038 143 1039
rect 136 1036 143 1038
rect 136 1035 137 1036
rect 131 1034 137 1035
rect 142 1035 143 1036
rect 147 1035 148 1039
rect 142 1034 148 1035
rect 171 1039 177 1040
rect 171 1035 172 1039
rect 176 1038 177 1039
rect 198 1039 204 1040
rect 198 1038 199 1039
rect 176 1036 199 1038
rect 176 1035 177 1036
rect 171 1034 177 1035
rect 198 1035 199 1036
rect 203 1035 204 1039
rect 198 1034 204 1035
rect 238 1039 249 1040
rect 238 1035 239 1039
rect 243 1035 244 1039
rect 248 1035 249 1039
rect 238 1034 249 1035
rect 323 1039 329 1040
rect 323 1035 324 1039
rect 328 1038 329 1039
rect 346 1039 352 1040
rect 346 1038 347 1039
rect 328 1036 347 1038
rect 328 1035 329 1036
rect 323 1034 329 1035
rect 346 1035 347 1036
rect 351 1035 352 1039
rect 346 1034 352 1035
rect 406 1039 417 1040
rect 406 1035 407 1039
rect 411 1035 412 1039
rect 416 1035 417 1039
rect 406 1034 417 1035
rect 494 1039 505 1040
rect 494 1035 495 1039
rect 499 1035 500 1039
rect 504 1035 505 1039
rect 494 1034 505 1035
rect 567 1039 573 1040
rect 567 1035 568 1039
rect 572 1038 573 1039
rect 579 1039 585 1040
rect 579 1038 580 1039
rect 572 1036 580 1038
rect 572 1035 573 1036
rect 567 1034 573 1035
rect 579 1035 580 1036
rect 584 1035 585 1039
rect 579 1034 585 1035
rect 659 1039 665 1040
rect 659 1035 660 1039
rect 664 1038 665 1039
rect 718 1039 724 1040
rect 718 1038 719 1039
rect 664 1036 719 1038
rect 664 1035 665 1036
rect 659 1034 665 1035
rect 718 1035 719 1036
rect 723 1035 724 1039
rect 718 1034 724 1035
rect 726 1039 737 1040
rect 726 1035 727 1039
rect 731 1035 732 1039
rect 736 1035 737 1039
rect 726 1034 737 1035
rect 790 1039 801 1040
rect 790 1035 791 1039
rect 795 1035 796 1039
rect 800 1035 801 1039
rect 790 1034 801 1035
rect 854 1039 865 1040
rect 854 1035 855 1039
rect 859 1035 860 1039
rect 864 1035 865 1039
rect 854 1034 865 1035
rect 910 1039 921 1040
rect 910 1035 911 1039
rect 915 1035 916 1039
rect 920 1035 921 1039
rect 910 1034 921 1035
rect 974 1039 985 1040
rect 974 1035 975 1039
rect 979 1035 980 1039
rect 984 1035 985 1039
rect 974 1034 985 1035
rect 1038 1039 1049 1040
rect 1038 1035 1039 1039
rect 1043 1035 1044 1039
rect 1048 1035 1049 1039
rect 1427 1039 1428 1043
rect 1432 1042 1433 1043
rect 1438 1043 1444 1044
rect 1438 1042 1439 1043
rect 1432 1040 1439 1042
rect 1432 1039 1433 1040
rect 1427 1038 1433 1039
rect 1438 1039 1439 1040
rect 1443 1039 1444 1043
rect 1438 1038 1444 1039
rect 1458 1043 1464 1044
rect 1458 1039 1459 1043
rect 1463 1042 1464 1043
rect 1467 1043 1473 1044
rect 1467 1042 1468 1043
rect 1463 1040 1468 1042
rect 1463 1039 1464 1040
rect 1458 1038 1464 1039
rect 1467 1039 1468 1040
rect 1472 1039 1473 1043
rect 1467 1038 1473 1039
rect 1498 1043 1504 1044
rect 1498 1039 1499 1043
rect 1503 1042 1504 1043
rect 1507 1043 1513 1044
rect 1507 1042 1508 1043
rect 1503 1040 1508 1042
rect 1503 1039 1504 1040
rect 1498 1038 1504 1039
rect 1507 1039 1508 1040
rect 1512 1039 1513 1043
rect 1507 1038 1513 1039
rect 1550 1043 1561 1044
rect 1550 1039 1551 1043
rect 1555 1039 1556 1043
rect 1560 1039 1561 1043
rect 1550 1038 1561 1039
rect 1606 1043 1617 1044
rect 1606 1039 1607 1043
rect 1611 1039 1612 1043
rect 1616 1039 1617 1043
rect 1606 1038 1617 1039
rect 1662 1043 1673 1044
rect 1662 1039 1663 1043
rect 1667 1039 1668 1043
rect 1672 1039 1673 1043
rect 1662 1038 1673 1039
rect 1714 1043 1720 1044
rect 1714 1039 1715 1043
rect 1719 1042 1720 1043
rect 1723 1043 1729 1044
rect 1723 1042 1724 1043
rect 1719 1040 1724 1042
rect 1719 1039 1720 1040
rect 1714 1038 1720 1039
rect 1723 1039 1724 1040
rect 1728 1039 1729 1043
rect 1723 1038 1729 1039
rect 1771 1043 1777 1044
rect 1771 1039 1772 1043
rect 1776 1042 1777 1043
rect 1782 1043 1788 1044
rect 1782 1042 1783 1043
rect 1776 1040 1783 1042
rect 1776 1039 1777 1040
rect 1771 1038 1777 1039
rect 1782 1039 1783 1040
rect 1787 1039 1788 1043
rect 1782 1038 1788 1039
rect 1819 1043 1825 1044
rect 1819 1039 1820 1043
rect 1824 1042 1825 1043
rect 1855 1043 1861 1044
rect 1855 1042 1856 1043
rect 1824 1040 1856 1042
rect 1824 1039 1825 1040
rect 1819 1038 1825 1039
rect 1855 1039 1856 1040
rect 1860 1039 1861 1043
rect 1855 1038 1861 1039
rect 1867 1043 1873 1044
rect 1867 1039 1868 1043
rect 1872 1042 1873 1043
rect 1903 1043 1909 1044
rect 1903 1042 1904 1043
rect 1872 1040 1904 1042
rect 1872 1039 1873 1040
rect 1867 1038 1873 1039
rect 1903 1039 1904 1040
rect 1908 1039 1909 1043
rect 1903 1038 1909 1039
rect 1915 1043 1921 1044
rect 1915 1039 1916 1043
rect 1920 1042 1921 1043
rect 1951 1043 1957 1044
rect 1951 1042 1952 1043
rect 1920 1040 1952 1042
rect 1920 1039 1921 1040
rect 1915 1038 1921 1039
rect 1951 1039 1952 1040
rect 1956 1039 1957 1043
rect 1951 1038 1957 1039
rect 1963 1043 1969 1044
rect 1963 1039 1964 1043
rect 1968 1042 1969 1043
rect 2002 1043 2008 1044
rect 2002 1042 2003 1043
rect 1968 1040 2003 1042
rect 1968 1039 1969 1040
rect 1963 1038 1969 1039
rect 2002 1039 2003 1040
rect 2007 1039 2008 1043
rect 2002 1038 2008 1039
rect 2011 1043 2017 1044
rect 2011 1039 2012 1043
rect 2016 1042 2017 1043
rect 2047 1043 2053 1044
rect 2047 1042 2048 1043
rect 2016 1040 2048 1042
rect 2016 1039 2017 1040
rect 2011 1038 2017 1039
rect 2047 1039 2048 1040
rect 2052 1039 2053 1043
rect 2047 1038 2053 1039
rect 2059 1043 2065 1044
rect 2059 1039 2060 1043
rect 2064 1042 2065 1043
rect 2095 1043 2101 1044
rect 2095 1042 2096 1043
rect 2064 1040 2096 1042
rect 2064 1039 2065 1040
rect 2059 1038 2065 1039
rect 2095 1039 2096 1040
rect 2100 1039 2101 1043
rect 2095 1038 2101 1039
rect 2110 1043 2121 1044
rect 2110 1039 2111 1043
rect 2115 1039 2116 1043
rect 2120 1039 2121 1043
rect 2110 1038 2121 1039
rect 2166 1043 2177 1044
rect 2166 1039 2167 1043
rect 2171 1039 2172 1043
rect 2176 1039 2177 1043
rect 2166 1038 2177 1039
rect 2222 1043 2233 1044
rect 2222 1039 2223 1043
rect 2227 1039 2228 1043
rect 2232 1039 2233 1043
rect 2222 1038 2233 1039
rect 1038 1034 1049 1035
rect 1571 1031 1577 1032
rect 171 1027 177 1028
rect 171 1023 172 1027
rect 176 1026 177 1027
rect 238 1027 244 1028
rect 238 1026 239 1027
rect 176 1024 239 1026
rect 176 1023 177 1024
rect 171 1022 177 1023
rect 238 1023 239 1024
rect 243 1023 244 1027
rect 238 1022 244 1023
rect 251 1027 257 1028
rect 251 1023 252 1027
rect 256 1026 257 1027
rect 278 1027 284 1028
rect 278 1026 279 1027
rect 256 1024 279 1026
rect 256 1023 257 1024
rect 251 1022 257 1023
rect 278 1023 279 1024
rect 283 1023 284 1027
rect 278 1022 284 1023
rect 323 1027 329 1028
rect 323 1023 324 1027
rect 328 1026 329 1027
rect 334 1027 340 1028
rect 334 1026 335 1027
rect 328 1024 335 1026
rect 328 1023 329 1024
rect 323 1022 329 1023
rect 334 1023 335 1024
rect 339 1023 340 1027
rect 334 1022 340 1023
rect 354 1027 360 1028
rect 354 1023 355 1027
rect 359 1026 360 1027
rect 395 1027 401 1028
rect 395 1026 396 1027
rect 359 1024 396 1026
rect 359 1023 360 1024
rect 354 1022 360 1023
rect 395 1023 396 1024
rect 400 1023 401 1027
rect 395 1022 401 1023
rect 426 1027 432 1028
rect 426 1023 427 1027
rect 431 1026 432 1027
rect 459 1027 465 1028
rect 459 1026 460 1027
rect 431 1024 460 1026
rect 431 1023 432 1024
rect 426 1022 432 1023
rect 459 1023 460 1024
rect 464 1023 465 1027
rect 459 1022 465 1023
rect 490 1027 496 1028
rect 490 1023 491 1027
rect 495 1026 496 1027
rect 515 1027 521 1028
rect 515 1026 516 1027
rect 495 1024 516 1026
rect 495 1023 496 1024
rect 490 1022 496 1023
rect 515 1023 516 1024
rect 520 1023 521 1027
rect 515 1022 521 1023
rect 546 1027 552 1028
rect 546 1023 547 1027
rect 551 1026 552 1027
rect 571 1027 577 1028
rect 571 1026 572 1027
rect 551 1024 572 1026
rect 551 1023 552 1024
rect 546 1022 552 1023
rect 571 1023 572 1024
rect 576 1023 577 1027
rect 571 1022 577 1023
rect 619 1027 625 1028
rect 619 1023 620 1027
rect 624 1026 625 1027
rect 630 1027 636 1028
rect 630 1026 631 1027
rect 624 1024 631 1026
rect 624 1023 625 1024
rect 619 1022 625 1023
rect 630 1023 631 1024
rect 635 1023 636 1027
rect 630 1022 636 1023
rect 650 1027 656 1028
rect 650 1023 651 1027
rect 655 1026 656 1027
rect 667 1027 673 1028
rect 667 1026 668 1027
rect 655 1024 668 1026
rect 655 1023 656 1024
rect 650 1022 656 1023
rect 667 1023 668 1024
rect 672 1023 673 1027
rect 667 1022 673 1023
rect 698 1027 704 1028
rect 698 1023 699 1027
rect 703 1026 704 1027
rect 731 1027 737 1028
rect 731 1026 732 1027
rect 703 1024 732 1026
rect 703 1023 704 1024
rect 698 1022 704 1023
rect 731 1023 732 1024
rect 736 1023 737 1027
rect 731 1022 737 1023
rect 762 1027 768 1028
rect 762 1023 763 1027
rect 767 1026 768 1027
rect 803 1027 809 1028
rect 803 1026 804 1027
rect 767 1024 804 1026
rect 767 1023 768 1024
rect 762 1022 768 1023
rect 803 1023 804 1024
rect 808 1023 809 1027
rect 803 1022 809 1023
rect 834 1027 840 1028
rect 834 1023 835 1027
rect 839 1026 840 1027
rect 891 1027 897 1028
rect 891 1026 892 1027
rect 839 1024 892 1026
rect 839 1023 840 1024
rect 834 1022 840 1023
rect 891 1023 892 1024
rect 896 1023 897 1027
rect 891 1022 897 1023
rect 926 1027 932 1028
rect 926 1023 927 1027
rect 931 1026 932 1027
rect 995 1027 1001 1028
rect 995 1026 996 1027
rect 931 1024 996 1026
rect 931 1023 932 1024
rect 926 1022 932 1023
rect 995 1023 996 1024
rect 1000 1023 1001 1027
rect 995 1022 1001 1023
rect 1026 1027 1032 1028
rect 1026 1023 1027 1027
rect 1031 1026 1032 1027
rect 1099 1027 1105 1028
rect 1099 1026 1100 1027
rect 1031 1024 1100 1026
rect 1031 1023 1032 1024
rect 1026 1022 1032 1023
rect 1099 1023 1100 1024
rect 1104 1023 1105 1027
rect 1099 1022 1105 1023
rect 1187 1027 1193 1028
rect 1187 1023 1188 1027
rect 1192 1026 1193 1027
rect 1214 1027 1220 1028
rect 1214 1026 1215 1027
rect 1192 1024 1215 1026
rect 1192 1023 1193 1024
rect 1187 1022 1193 1023
rect 1214 1023 1215 1024
rect 1219 1023 1220 1027
rect 1571 1027 1572 1031
rect 1576 1030 1577 1031
rect 1582 1031 1588 1032
rect 1582 1030 1583 1031
rect 1576 1028 1583 1030
rect 1576 1027 1577 1028
rect 1571 1026 1577 1027
rect 1582 1027 1583 1028
rect 1587 1027 1588 1031
rect 1582 1026 1588 1027
rect 1602 1031 1608 1032
rect 1602 1027 1603 1031
rect 1607 1030 1608 1031
rect 1611 1031 1617 1032
rect 1611 1030 1612 1031
rect 1607 1028 1612 1030
rect 1607 1027 1608 1028
rect 1602 1026 1608 1027
rect 1611 1027 1612 1028
rect 1616 1027 1617 1031
rect 1611 1026 1617 1027
rect 1642 1031 1648 1032
rect 1642 1027 1643 1031
rect 1647 1030 1648 1031
rect 1651 1031 1657 1032
rect 1651 1030 1652 1031
rect 1647 1028 1652 1030
rect 1647 1027 1648 1028
rect 1642 1026 1648 1027
rect 1651 1027 1652 1028
rect 1656 1027 1657 1031
rect 1651 1026 1657 1027
rect 1682 1031 1688 1032
rect 1682 1027 1683 1031
rect 1687 1030 1688 1031
rect 1691 1031 1697 1032
rect 1691 1030 1692 1031
rect 1687 1028 1692 1030
rect 1687 1027 1688 1028
rect 1682 1026 1688 1027
rect 1691 1027 1692 1028
rect 1696 1027 1697 1031
rect 1691 1026 1697 1027
rect 1718 1031 1724 1032
rect 1718 1027 1719 1031
rect 1723 1030 1724 1031
rect 1731 1031 1737 1032
rect 1731 1030 1732 1031
rect 1723 1028 1732 1030
rect 1723 1027 1724 1028
rect 1718 1026 1724 1027
rect 1731 1027 1732 1028
rect 1736 1027 1737 1031
rect 1731 1026 1737 1027
rect 1762 1031 1768 1032
rect 1762 1027 1763 1031
rect 1767 1030 1768 1031
rect 1771 1031 1777 1032
rect 1771 1030 1772 1031
rect 1767 1028 1772 1030
rect 1767 1027 1768 1028
rect 1762 1026 1768 1027
rect 1771 1027 1772 1028
rect 1776 1027 1777 1031
rect 1771 1026 1777 1027
rect 1814 1031 1825 1032
rect 1814 1027 1815 1031
rect 1819 1027 1820 1031
rect 1824 1027 1825 1031
rect 1814 1026 1825 1027
rect 1850 1031 1856 1032
rect 1850 1027 1851 1031
rect 1855 1030 1856 1031
rect 1875 1031 1881 1032
rect 1875 1030 1876 1031
rect 1855 1028 1876 1030
rect 1855 1027 1856 1028
rect 1850 1026 1856 1027
rect 1875 1027 1876 1028
rect 1880 1027 1881 1031
rect 1875 1026 1881 1027
rect 1906 1031 1912 1032
rect 1906 1027 1907 1031
rect 1911 1030 1912 1031
rect 1939 1031 1945 1032
rect 1939 1030 1940 1031
rect 1911 1028 1940 1030
rect 1911 1027 1912 1028
rect 1906 1026 1912 1027
rect 1939 1027 1940 1028
rect 1944 1027 1945 1031
rect 1939 1026 1945 1027
rect 1983 1031 1989 1032
rect 1983 1027 1984 1031
rect 1988 1030 1989 1031
rect 2011 1031 2017 1032
rect 2011 1030 2012 1031
rect 1988 1028 2012 1030
rect 1988 1027 1989 1028
rect 1983 1026 1989 1027
rect 2011 1027 2012 1028
rect 2016 1027 2017 1031
rect 2011 1026 2017 1027
rect 2091 1031 2097 1032
rect 2091 1027 2092 1031
rect 2096 1030 2097 1031
rect 2126 1031 2132 1032
rect 2126 1030 2127 1031
rect 2096 1028 2127 1030
rect 2096 1027 2097 1028
rect 2091 1026 2097 1027
rect 2126 1027 2127 1028
rect 2131 1027 2132 1031
rect 2126 1026 2132 1027
rect 2171 1031 2177 1032
rect 2171 1027 2172 1031
rect 2176 1030 2177 1031
rect 2238 1031 2244 1032
rect 2238 1030 2239 1031
rect 2176 1028 2239 1030
rect 2176 1027 2177 1028
rect 2171 1026 2177 1027
rect 2238 1027 2239 1028
rect 2243 1027 2244 1031
rect 2238 1026 2244 1027
rect 2246 1031 2257 1032
rect 2246 1027 2247 1031
rect 2251 1027 2252 1031
rect 2256 1027 2257 1031
rect 2246 1026 2257 1027
rect 1214 1022 1220 1023
rect 1574 1023 1580 1024
rect 174 1019 180 1020
rect 174 1015 175 1019
rect 179 1015 180 1019
rect 174 1014 180 1015
rect 254 1019 260 1020
rect 254 1015 255 1019
rect 259 1015 260 1019
rect 254 1014 260 1015
rect 326 1019 332 1020
rect 326 1015 327 1019
rect 331 1015 332 1019
rect 326 1014 332 1015
rect 398 1019 404 1020
rect 398 1015 399 1019
rect 403 1015 404 1019
rect 398 1014 404 1015
rect 462 1019 468 1020
rect 462 1015 463 1019
rect 467 1015 468 1019
rect 462 1014 468 1015
rect 518 1019 524 1020
rect 518 1015 519 1019
rect 523 1015 524 1019
rect 518 1014 524 1015
rect 574 1019 580 1020
rect 574 1015 575 1019
rect 579 1015 580 1019
rect 574 1014 580 1015
rect 622 1019 628 1020
rect 622 1015 623 1019
rect 627 1015 628 1019
rect 622 1014 628 1015
rect 670 1019 676 1020
rect 670 1015 671 1019
rect 675 1015 676 1019
rect 670 1014 676 1015
rect 734 1019 740 1020
rect 734 1015 735 1019
rect 739 1015 740 1019
rect 734 1014 740 1015
rect 806 1019 812 1020
rect 806 1015 807 1019
rect 811 1015 812 1019
rect 806 1014 812 1015
rect 894 1019 900 1020
rect 894 1015 895 1019
rect 899 1015 900 1019
rect 894 1014 900 1015
rect 998 1019 1004 1020
rect 998 1015 999 1019
rect 1003 1015 1004 1019
rect 998 1014 1004 1015
rect 1102 1019 1108 1020
rect 1102 1015 1103 1019
rect 1107 1015 1108 1019
rect 1102 1014 1108 1015
rect 1190 1019 1196 1020
rect 1190 1015 1191 1019
rect 1195 1015 1196 1019
rect 1574 1019 1575 1023
rect 1579 1019 1580 1023
rect 1574 1018 1580 1019
rect 1614 1023 1620 1024
rect 1614 1019 1615 1023
rect 1619 1019 1620 1023
rect 1614 1018 1620 1019
rect 1654 1023 1660 1024
rect 1654 1019 1655 1023
rect 1659 1019 1660 1023
rect 1654 1018 1660 1019
rect 1694 1023 1700 1024
rect 1694 1019 1695 1023
rect 1699 1019 1700 1023
rect 1694 1018 1700 1019
rect 1734 1023 1740 1024
rect 1734 1019 1735 1023
rect 1739 1019 1740 1023
rect 1734 1018 1740 1019
rect 1774 1023 1780 1024
rect 1774 1019 1775 1023
rect 1779 1019 1780 1023
rect 1774 1018 1780 1019
rect 1822 1023 1828 1024
rect 1822 1019 1823 1023
rect 1827 1019 1828 1023
rect 1822 1018 1828 1019
rect 1878 1023 1884 1024
rect 1878 1019 1879 1023
rect 1883 1019 1884 1023
rect 1878 1018 1884 1019
rect 1942 1023 1948 1024
rect 1942 1019 1943 1023
rect 1947 1019 1948 1023
rect 1942 1018 1948 1019
rect 2014 1023 2020 1024
rect 2014 1019 2015 1023
rect 2019 1019 2020 1023
rect 2014 1018 2020 1019
rect 2094 1023 2100 1024
rect 2094 1019 2095 1023
rect 2099 1019 2100 1023
rect 2094 1018 2100 1019
rect 2174 1023 2180 1024
rect 2174 1019 2175 1023
rect 2179 1019 2180 1023
rect 2174 1018 2180 1019
rect 2254 1023 2260 1024
rect 2254 1019 2255 1023
rect 2259 1019 2260 1023
rect 2254 1018 2260 1019
rect 1190 1014 1196 1015
rect 1278 1000 1284 1001
rect 2406 1000 2412 1001
rect 110 996 116 997
rect 110 992 111 996
rect 115 992 116 996
rect 1238 996 1244 997
rect 1238 992 1239 996
rect 1243 992 1244 996
rect 1278 996 1279 1000
rect 1283 996 1284 1000
rect 1983 999 1989 1000
rect 1983 998 1984 999
rect 1967 997 1984 998
rect 1278 995 1284 996
rect 1599 995 1608 996
rect 110 991 116 992
rect 198 991 205 992
rect 198 987 199 991
rect 204 987 205 991
rect 198 986 205 987
rect 238 991 244 992
rect 238 987 239 991
rect 243 990 244 991
rect 279 991 285 992
rect 279 990 280 991
rect 243 988 280 990
rect 243 987 244 988
rect 238 986 244 987
rect 279 987 280 988
rect 284 987 285 991
rect 279 986 285 987
rect 351 991 360 992
rect 351 987 352 991
rect 359 987 360 991
rect 351 986 360 987
rect 423 991 432 992
rect 423 987 424 991
rect 431 987 432 991
rect 423 986 432 987
rect 487 991 496 992
rect 487 987 488 991
rect 495 987 496 991
rect 487 986 496 987
rect 543 991 552 992
rect 543 987 544 991
rect 551 987 552 991
rect 599 991 605 992
rect 599 990 600 991
rect 543 986 552 987
rect 556 988 600 990
rect 470 983 476 984
rect 110 979 116 980
rect 110 975 111 979
rect 115 975 116 979
rect 470 979 471 983
rect 475 982 476 983
rect 556 982 558 988
rect 599 987 600 988
rect 604 987 605 991
rect 599 986 605 987
rect 647 991 656 992
rect 647 987 648 991
rect 655 987 656 991
rect 647 986 656 987
rect 695 991 704 992
rect 695 987 696 991
rect 703 987 704 991
rect 695 986 704 987
rect 759 991 768 992
rect 759 987 760 991
rect 767 987 768 991
rect 759 986 768 987
rect 831 991 840 992
rect 831 987 832 991
rect 839 987 840 991
rect 831 986 840 987
rect 919 991 928 992
rect 919 987 920 991
rect 927 987 928 991
rect 919 986 928 987
rect 1023 991 1032 992
rect 1023 987 1024 991
rect 1031 987 1032 991
rect 1023 986 1032 987
rect 1126 991 1133 992
rect 1126 987 1127 991
rect 1132 987 1133 991
rect 1126 986 1133 987
rect 1150 991 1156 992
rect 1150 987 1151 991
rect 1155 990 1156 991
rect 1215 991 1221 992
rect 1238 991 1244 992
rect 1599 991 1600 995
rect 1607 991 1608 995
rect 1215 990 1216 991
rect 1155 988 1216 990
rect 1155 987 1156 988
rect 1150 986 1156 987
rect 1215 987 1216 988
rect 1220 987 1221 991
rect 1599 990 1608 991
rect 1639 995 1648 996
rect 1639 991 1640 995
rect 1647 991 1648 995
rect 1639 990 1648 991
rect 1679 995 1688 996
rect 1679 991 1680 995
rect 1687 991 1688 995
rect 1679 990 1688 991
rect 1718 995 1725 996
rect 1718 991 1719 995
rect 1724 991 1725 995
rect 1718 990 1725 991
rect 1759 995 1768 996
rect 1759 991 1760 995
rect 1767 991 1768 995
rect 1799 995 1805 996
rect 1799 994 1800 995
rect 1759 990 1768 991
rect 1772 992 1800 994
rect 1215 986 1221 987
rect 1686 987 1692 988
rect 475 980 558 982
rect 1278 983 1284 984
rect 475 979 476 980
rect 470 978 476 979
rect 1238 979 1244 980
rect 110 974 116 975
rect 1238 975 1239 979
rect 1243 975 1244 979
rect 1278 979 1279 983
rect 1283 979 1284 983
rect 1686 983 1687 987
rect 1691 986 1692 987
rect 1772 986 1774 992
rect 1799 991 1800 992
rect 1804 991 1805 995
rect 1799 990 1805 991
rect 1847 995 1856 996
rect 1847 991 1848 995
rect 1855 991 1856 995
rect 1847 990 1856 991
rect 1903 995 1912 996
rect 1903 991 1904 995
rect 1911 991 1912 995
rect 1967 993 1968 997
rect 1972 996 1984 997
rect 1972 993 1973 996
rect 1983 995 1984 996
rect 1988 995 1989 999
rect 2406 996 2407 1000
rect 2411 996 2412 1000
rect 1983 994 1989 995
rect 1991 995 1997 996
rect 1967 992 1973 993
rect 1903 990 1912 991
rect 1991 991 1992 995
rect 1996 994 1997 995
rect 2039 995 2045 996
rect 2039 994 2040 995
rect 1996 992 2040 994
rect 1996 991 1997 992
rect 1991 990 1997 991
rect 2039 991 2040 992
rect 2044 991 2045 995
rect 2039 990 2045 991
rect 2110 995 2116 996
rect 2110 991 2111 995
rect 2115 994 2116 995
rect 2119 995 2125 996
rect 2119 994 2120 995
rect 2115 992 2120 994
rect 2115 991 2116 992
rect 2110 990 2116 991
rect 2119 991 2120 992
rect 2124 991 2125 995
rect 2119 990 2125 991
rect 2190 995 2196 996
rect 2190 991 2191 995
rect 2195 994 2196 995
rect 2199 995 2205 996
rect 2199 994 2200 995
rect 2195 992 2200 994
rect 2195 991 2196 992
rect 2190 990 2196 991
rect 2199 991 2200 992
rect 2204 991 2205 995
rect 2199 990 2205 991
rect 2238 995 2244 996
rect 2238 991 2239 995
rect 2243 994 2244 995
rect 2279 995 2285 996
rect 2406 995 2412 996
rect 2279 994 2280 995
rect 2243 992 2280 994
rect 2243 991 2244 992
rect 2238 990 2244 991
rect 2279 991 2280 992
rect 2284 991 2285 995
rect 2279 990 2285 991
rect 1691 984 1774 986
rect 1691 983 1692 984
rect 1686 982 1692 983
rect 2406 983 2412 984
rect 1278 978 1284 979
rect 2406 979 2407 983
rect 2411 979 2412 983
rect 2406 978 2412 979
rect 1238 974 1244 975
rect 1574 976 1580 977
rect 174 972 180 973
rect 174 968 175 972
rect 179 968 180 972
rect 174 967 180 968
rect 254 972 260 973
rect 254 968 255 972
rect 259 968 260 972
rect 254 967 260 968
rect 326 972 332 973
rect 326 968 327 972
rect 331 968 332 972
rect 326 967 332 968
rect 398 972 404 973
rect 398 968 399 972
rect 403 968 404 972
rect 398 967 404 968
rect 462 972 468 973
rect 462 968 463 972
rect 467 968 468 972
rect 462 967 468 968
rect 518 972 524 973
rect 518 968 519 972
rect 523 968 524 972
rect 518 967 524 968
rect 574 972 580 973
rect 574 968 575 972
rect 579 968 580 972
rect 574 967 580 968
rect 622 972 628 973
rect 622 968 623 972
rect 627 968 628 972
rect 622 967 628 968
rect 670 972 676 973
rect 670 968 671 972
rect 675 968 676 972
rect 670 967 676 968
rect 734 972 740 973
rect 734 968 735 972
rect 739 968 740 972
rect 734 967 740 968
rect 806 972 812 973
rect 806 968 807 972
rect 811 968 812 972
rect 806 967 812 968
rect 894 972 900 973
rect 894 968 895 972
rect 899 968 900 972
rect 894 967 900 968
rect 998 972 1004 973
rect 998 968 999 972
rect 1003 968 1004 972
rect 998 967 1004 968
rect 1102 972 1108 973
rect 1102 968 1103 972
rect 1107 968 1108 972
rect 1102 967 1108 968
rect 1190 972 1196 973
rect 1190 968 1191 972
rect 1195 968 1196 972
rect 1574 972 1575 976
rect 1579 972 1580 976
rect 1574 971 1580 972
rect 1614 976 1620 977
rect 1614 972 1615 976
rect 1619 972 1620 976
rect 1614 971 1620 972
rect 1654 976 1660 977
rect 1654 972 1655 976
rect 1659 972 1660 976
rect 1654 971 1660 972
rect 1694 976 1700 977
rect 1694 972 1695 976
rect 1699 972 1700 976
rect 1694 971 1700 972
rect 1734 976 1740 977
rect 1734 972 1735 976
rect 1739 972 1740 976
rect 1734 971 1740 972
rect 1774 976 1780 977
rect 1774 972 1775 976
rect 1779 972 1780 976
rect 1774 971 1780 972
rect 1822 976 1828 977
rect 1822 972 1823 976
rect 1827 972 1828 976
rect 1822 971 1828 972
rect 1878 976 1884 977
rect 1878 972 1879 976
rect 1883 972 1884 976
rect 1878 971 1884 972
rect 1942 976 1948 977
rect 1942 972 1943 976
rect 1947 972 1948 976
rect 1942 971 1948 972
rect 2014 976 2020 977
rect 2014 972 2015 976
rect 2019 972 2020 976
rect 2014 971 2020 972
rect 2094 976 2100 977
rect 2094 972 2095 976
rect 2099 972 2100 976
rect 2094 971 2100 972
rect 2174 976 2180 977
rect 2174 972 2175 976
rect 2179 972 2180 976
rect 2174 971 2180 972
rect 2254 976 2260 977
rect 2254 972 2255 976
rect 2259 972 2260 976
rect 2254 971 2260 972
rect 1190 967 1196 968
rect 214 960 220 961
rect 214 956 215 960
rect 219 956 220 960
rect 214 955 220 956
rect 254 960 260 961
rect 254 956 255 960
rect 259 956 260 960
rect 254 955 260 956
rect 302 960 308 961
rect 302 956 303 960
rect 307 956 308 960
rect 302 955 308 956
rect 358 960 364 961
rect 358 956 359 960
rect 363 956 364 960
rect 358 955 364 956
rect 414 960 420 961
rect 414 956 415 960
rect 419 956 420 960
rect 414 955 420 956
rect 462 960 468 961
rect 462 956 463 960
rect 467 956 468 960
rect 462 955 468 956
rect 518 960 524 961
rect 518 956 519 960
rect 523 956 524 960
rect 518 955 524 956
rect 574 960 580 961
rect 574 956 575 960
rect 579 956 580 960
rect 574 955 580 956
rect 638 960 644 961
rect 638 956 639 960
rect 643 956 644 960
rect 638 955 644 956
rect 710 960 716 961
rect 710 956 711 960
rect 715 956 716 960
rect 710 955 716 956
rect 782 960 788 961
rect 782 956 783 960
rect 787 956 788 960
rect 782 955 788 956
rect 854 960 860 961
rect 854 956 855 960
rect 859 956 860 960
rect 854 955 860 956
rect 926 960 932 961
rect 926 956 927 960
rect 931 956 932 960
rect 926 955 932 956
rect 998 960 1004 961
rect 998 956 999 960
rect 1003 956 1004 960
rect 998 955 1004 956
rect 1070 960 1076 961
rect 1070 956 1071 960
rect 1075 956 1076 960
rect 1070 955 1076 956
rect 1142 960 1148 961
rect 1142 956 1143 960
rect 1147 956 1148 960
rect 1142 955 1148 956
rect 1190 960 1196 961
rect 1190 956 1191 960
rect 1195 956 1196 960
rect 1190 955 1196 956
rect 1302 956 1308 957
rect 110 953 116 954
rect 110 949 111 953
rect 115 949 116 953
rect 110 948 116 949
rect 1238 953 1244 954
rect 1238 949 1239 953
rect 1243 949 1244 953
rect 1302 952 1303 956
rect 1307 952 1308 956
rect 1302 951 1308 952
rect 1350 956 1356 957
rect 1350 952 1351 956
rect 1355 952 1356 956
rect 1350 951 1356 952
rect 1430 956 1436 957
rect 1430 952 1431 956
rect 1435 952 1436 956
rect 1430 951 1436 952
rect 1510 956 1516 957
rect 1510 952 1511 956
rect 1515 952 1516 956
rect 1510 951 1516 952
rect 1590 956 1596 957
rect 1590 952 1591 956
rect 1595 952 1596 956
rect 1590 951 1596 952
rect 1678 956 1684 957
rect 1678 952 1679 956
rect 1683 952 1684 956
rect 1678 951 1684 952
rect 1766 956 1772 957
rect 1766 952 1767 956
rect 1771 952 1772 956
rect 1766 951 1772 952
rect 1854 956 1860 957
rect 1854 952 1855 956
rect 1859 952 1860 956
rect 1854 951 1860 952
rect 1942 956 1948 957
rect 1942 952 1943 956
rect 1947 952 1948 956
rect 1942 951 1948 952
rect 2022 956 2028 957
rect 2022 952 2023 956
rect 2027 952 2028 956
rect 2022 951 2028 952
rect 2102 956 2108 957
rect 2102 952 2103 956
rect 2107 952 2108 956
rect 2102 951 2108 952
rect 2182 956 2188 957
rect 2182 952 2183 956
rect 2187 952 2188 956
rect 2182 951 2188 952
rect 2270 956 2276 957
rect 2270 952 2271 956
rect 2275 952 2276 956
rect 2270 951 2276 952
rect 1238 948 1244 949
rect 1278 949 1284 950
rect 630 947 636 948
rect 630 943 631 947
rect 635 946 636 947
rect 635 944 858 946
rect 1278 945 1279 949
rect 1283 945 1284 949
rect 1278 944 1284 945
rect 2406 949 2412 950
rect 2406 945 2407 949
rect 2411 945 2412 949
rect 2406 944 2412 945
rect 635 943 636 944
rect 630 942 636 943
rect 239 939 248 940
rect 110 936 116 937
rect 110 932 111 936
rect 115 932 116 936
rect 239 935 240 939
rect 247 935 248 939
rect 239 934 248 935
rect 278 939 285 940
rect 278 935 279 939
rect 284 935 285 939
rect 327 939 333 940
rect 327 938 328 939
rect 278 934 285 935
rect 288 936 328 938
rect 110 931 116 932
rect 222 931 228 932
rect 222 927 223 931
rect 227 930 228 931
rect 288 930 290 936
rect 327 935 328 936
rect 332 935 333 939
rect 327 934 333 935
rect 346 939 352 940
rect 346 935 347 939
rect 351 938 352 939
rect 383 939 389 940
rect 383 938 384 939
rect 351 936 384 938
rect 351 935 352 936
rect 346 934 352 935
rect 383 935 384 936
rect 388 935 389 939
rect 383 934 389 935
rect 391 939 397 940
rect 391 935 392 939
rect 396 938 397 939
rect 439 939 445 940
rect 439 938 440 939
rect 396 936 440 938
rect 396 935 397 936
rect 391 934 397 935
rect 439 935 440 936
rect 444 935 445 939
rect 439 934 445 935
rect 487 939 493 940
rect 487 935 488 939
rect 492 938 493 939
rect 502 939 508 940
rect 502 938 503 939
rect 492 936 503 938
rect 492 935 493 936
rect 487 934 493 935
rect 502 935 503 936
rect 507 935 508 939
rect 502 934 508 935
rect 543 939 549 940
rect 543 935 544 939
rect 548 938 549 939
rect 558 939 564 940
rect 558 938 559 939
rect 548 936 559 938
rect 548 935 549 936
rect 543 934 549 935
rect 558 935 559 936
rect 563 935 564 939
rect 558 934 564 935
rect 599 939 605 940
rect 599 935 600 939
rect 604 938 605 939
rect 630 939 636 940
rect 630 938 631 939
rect 604 936 631 938
rect 604 935 605 936
rect 599 934 605 935
rect 630 935 631 936
rect 635 935 636 939
rect 630 934 636 935
rect 663 939 669 940
rect 663 935 664 939
rect 668 938 669 939
rect 702 939 708 940
rect 702 938 703 939
rect 668 936 703 938
rect 668 935 669 936
rect 663 934 669 935
rect 702 935 703 936
rect 707 935 708 939
rect 702 934 708 935
rect 735 939 741 940
rect 735 935 736 939
rect 740 938 741 939
rect 774 939 780 940
rect 774 938 775 939
rect 740 936 775 938
rect 740 935 741 936
rect 735 934 741 935
rect 774 935 775 936
rect 779 935 780 939
rect 774 934 780 935
rect 807 939 813 940
rect 807 935 808 939
rect 812 938 813 939
rect 846 939 852 940
rect 846 938 847 939
rect 812 936 847 938
rect 812 935 813 936
rect 807 934 813 935
rect 846 935 847 936
rect 851 935 852 939
rect 856 938 858 944
rect 879 939 885 940
rect 879 938 880 939
rect 856 936 880 938
rect 846 934 852 935
rect 879 935 880 936
rect 884 935 885 939
rect 879 934 885 935
rect 951 939 957 940
rect 951 935 952 939
rect 956 938 957 939
rect 990 939 996 940
rect 990 938 991 939
rect 956 936 991 938
rect 956 935 957 936
rect 951 934 957 935
rect 990 935 991 936
rect 995 935 996 939
rect 990 934 996 935
rect 1014 939 1020 940
rect 1014 935 1015 939
rect 1019 938 1020 939
rect 1023 939 1029 940
rect 1023 938 1024 939
rect 1019 936 1024 938
rect 1019 935 1020 936
rect 1014 934 1020 935
rect 1023 935 1024 936
rect 1028 935 1029 939
rect 1095 939 1101 940
rect 1095 938 1096 939
rect 1023 934 1029 935
rect 1032 936 1096 938
rect 227 928 290 930
rect 938 931 944 932
rect 227 927 228 928
rect 222 926 228 927
rect 938 927 939 931
rect 943 930 944 931
rect 1032 930 1034 936
rect 1095 935 1096 936
rect 1100 935 1101 939
rect 1095 934 1101 935
rect 1103 939 1109 940
rect 1103 935 1104 939
rect 1108 938 1109 939
rect 1167 939 1173 940
rect 1167 938 1168 939
rect 1108 936 1168 938
rect 1108 935 1109 936
rect 1103 934 1109 935
rect 1167 935 1168 936
rect 1172 935 1173 939
rect 1167 934 1173 935
rect 1214 939 1221 940
rect 1214 935 1215 939
rect 1220 935 1221 939
rect 1214 934 1221 935
rect 1238 936 1244 937
rect 1238 932 1239 936
rect 1243 932 1244 936
rect 1286 935 1292 936
rect 1238 931 1244 932
rect 1278 932 1284 933
rect 943 928 1034 930
rect 1278 928 1279 932
rect 1283 928 1284 932
rect 1286 931 1287 935
rect 1291 934 1292 935
rect 1327 935 1333 936
rect 1327 934 1328 935
rect 1291 932 1328 934
rect 1291 931 1292 932
rect 1286 930 1292 931
rect 1327 931 1328 932
rect 1332 931 1333 935
rect 1327 930 1333 931
rect 1335 935 1341 936
rect 1335 931 1336 935
rect 1340 934 1341 935
rect 1375 935 1381 936
rect 1375 934 1376 935
rect 1340 932 1376 934
rect 1340 931 1341 932
rect 1335 930 1341 931
rect 1375 931 1376 932
rect 1380 931 1381 935
rect 1375 930 1381 931
rect 1383 935 1389 936
rect 1383 931 1384 935
rect 1388 934 1389 935
rect 1455 935 1461 936
rect 1455 934 1456 935
rect 1388 932 1456 934
rect 1388 931 1389 932
rect 1383 930 1389 931
rect 1455 931 1456 932
rect 1460 931 1461 935
rect 1455 930 1461 931
rect 1463 935 1469 936
rect 1463 931 1464 935
rect 1468 934 1469 935
rect 1535 935 1541 936
rect 1535 934 1536 935
rect 1468 932 1536 934
rect 1468 931 1469 932
rect 1463 930 1469 931
rect 1535 931 1536 932
rect 1540 931 1541 935
rect 1535 930 1541 931
rect 1615 935 1621 936
rect 1615 931 1616 935
rect 1620 934 1621 935
rect 1646 935 1652 936
rect 1646 934 1647 935
rect 1620 932 1647 934
rect 1620 931 1621 932
rect 1615 930 1621 931
rect 1646 931 1647 932
rect 1651 931 1652 935
rect 1646 930 1652 931
rect 1655 935 1661 936
rect 1655 931 1656 935
rect 1660 934 1661 935
rect 1703 935 1709 936
rect 1703 934 1704 935
rect 1660 932 1704 934
rect 1660 931 1661 932
rect 1655 930 1661 931
rect 1703 931 1704 932
rect 1708 931 1709 935
rect 1703 930 1709 931
rect 1782 935 1788 936
rect 1782 931 1783 935
rect 1787 934 1788 935
rect 1791 935 1797 936
rect 1791 934 1792 935
rect 1787 932 1792 934
rect 1787 931 1788 932
rect 1782 930 1788 931
rect 1791 931 1792 932
rect 1796 931 1797 935
rect 1791 930 1797 931
rect 1799 935 1805 936
rect 1799 931 1800 935
rect 1804 934 1805 935
rect 1879 935 1885 936
rect 1879 934 1880 935
rect 1804 932 1880 934
rect 1804 931 1805 932
rect 1799 930 1805 931
rect 1879 931 1880 932
rect 1884 931 1885 935
rect 1879 930 1885 931
rect 1887 935 1893 936
rect 1887 931 1888 935
rect 1892 934 1893 935
rect 1967 935 1973 936
rect 1967 934 1968 935
rect 1892 932 1968 934
rect 1892 931 1893 932
rect 1887 930 1893 931
rect 1967 931 1968 932
rect 1972 931 1973 935
rect 1967 930 1973 931
rect 2047 935 2053 936
rect 2047 931 2048 935
rect 2052 934 2053 935
rect 2094 935 2100 936
rect 2094 934 2095 935
rect 2052 932 2095 934
rect 2052 931 2053 932
rect 2047 930 2053 931
rect 2094 931 2095 932
rect 2099 931 2100 935
rect 2094 930 2100 931
rect 2126 935 2133 936
rect 2126 931 2127 935
rect 2132 931 2133 935
rect 2126 930 2133 931
rect 2207 935 2213 936
rect 2207 931 2208 935
rect 2212 934 2213 935
rect 2262 935 2268 936
rect 2262 934 2263 935
rect 2212 932 2263 934
rect 2212 931 2213 932
rect 2207 930 2213 931
rect 2262 931 2263 932
rect 2267 931 2268 935
rect 2262 930 2268 931
rect 2286 935 2292 936
rect 2286 931 2287 935
rect 2291 934 2292 935
rect 2295 935 2301 936
rect 2295 934 2296 935
rect 2291 932 2296 934
rect 2291 931 2292 932
rect 2286 930 2292 931
rect 2295 931 2296 932
rect 2300 931 2301 935
rect 2295 930 2301 931
rect 2406 932 2412 933
rect 943 927 944 928
rect 1278 927 1284 928
rect 2406 928 2407 932
rect 2411 928 2412 932
rect 2406 927 2412 928
rect 938 926 944 927
rect 214 913 220 914
rect 214 909 215 913
rect 219 909 220 913
rect 214 908 220 909
rect 254 913 260 914
rect 254 909 255 913
rect 259 909 260 913
rect 254 908 260 909
rect 302 913 308 914
rect 302 909 303 913
rect 307 909 308 913
rect 302 908 308 909
rect 358 913 364 914
rect 358 909 359 913
rect 363 909 364 913
rect 358 908 364 909
rect 414 913 420 914
rect 414 909 415 913
rect 419 909 420 913
rect 414 908 420 909
rect 462 913 468 914
rect 462 909 463 913
rect 467 909 468 913
rect 462 908 468 909
rect 518 913 524 914
rect 518 909 519 913
rect 523 909 524 913
rect 518 908 524 909
rect 574 913 580 914
rect 574 909 575 913
rect 579 909 580 913
rect 574 908 580 909
rect 638 913 644 914
rect 638 909 639 913
rect 643 909 644 913
rect 638 908 644 909
rect 710 913 716 914
rect 710 909 711 913
rect 715 909 716 913
rect 710 908 716 909
rect 782 913 788 914
rect 782 909 783 913
rect 787 909 788 913
rect 782 908 788 909
rect 854 913 860 914
rect 854 909 855 913
rect 859 909 860 913
rect 854 908 860 909
rect 926 913 932 914
rect 926 909 927 913
rect 931 909 932 913
rect 926 908 932 909
rect 998 913 1004 914
rect 998 909 999 913
rect 1003 909 1004 913
rect 998 908 1004 909
rect 1070 913 1076 914
rect 1070 909 1071 913
rect 1075 909 1076 913
rect 1070 908 1076 909
rect 1142 913 1148 914
rect 1142 909 1143 913
rect 1147 909 1148 913
rect 1142 908 1148 909
rect 1190 913 1196 914
rect 1190 909 1191 913
rect 1195 909 1196 913
rect 1190 908 1196 909
rect 1302 909 1308 910
rect 1302 905 1303 909
rect 1307 905 1308 909
rect 1302 904 1308 905
rect 1350 909 1356 910
rect 1350 905 1351 909
rect 1355 905 1356 909
rect 1350 904 1356 905
rect 1430 909 1436 910
rect 1430 905 1431 909
rect 1435 905 1436 909
rect 1430 904 1436 905
rect 1510 909 1516 910
rect 1510 905 1511 909
rect 1515 905 1516 909
rect 1510 904 1516 905
rect 1590 909 1596 910
rect 1590 905 1591 909
rect 1595 905 1596 909
rect 1590 904 1596 905
rect 1678 909 1684 910
rect 1678 905 1679 909
rect 1683 905 1684 909
rect 1678 904 1684 905
rect 1766 909 1772 910
rect 1766 905 1767 909
rect 1771 905 1772 909
rect 1766 904 1772 905
rect 1854 909 1860 910
rect 1854 905 1855 909
rect 1859 905 1860 909
rect 1854 904 1860 905
rect 1942 909 1948 910
rect 1942 905 1943 909
rect 1947 905 1948 909
rect 1942 904 1948 905
rect 2022 909 2028 910
rect 2022 905 2023 909
rect 2027 905 2028 909
rect 2022 904 2028 905
rect 2102 909 2108 910
rect 2102 905 2103 909
rect 2107 905 2108 909
rect 2102 904 2108 905
rect 2182 909 2188 910
rect 2182 905 2183 909
rect 2187 905 2188 909
rect 2182 904 2188 905
rect 2270 909 2276 910
rect 2270 905 2271 909
rect 2275 905 2276 909
rect 2270 904 2276 905
rect 211 903 217 904
rect 211 899 212 903
rect 216 902 217 903
rect 222 903 228 904
rect 222 902 223 903
rect 216 900 223 902
rect 216 899 217 900
rect 211 898 217 899
rect 222 899 223 900
rect 227 899 228 903
rect 222 898 228 899
rect 242 903 248 904
rect 242 899 243 903
rect 247 902 248 903
rect 251 903 257 904
rect 251 902 252 903
rect 247 900 252 902
rect 247 899 248 900
rect 242 898 248 899
rect 251 899 252 900
rect 256 899 257 903
rect 251 898 257 899
rect 299 903 305 904
rect 299 899 300 903
rect 304 902 305 903
rect 346 903 352 904
rect 346 902 347 903
rect 304 900 347 902
rect 304 899 305 900
rect 299 898 305 899
rect 346 899 347 900
rect 351 899 352 903
rect 346 898 352 899
rect 355 903 361 904
rect 355 899 356 903
rect 360 902 361 903
rect 391 903 397 904
rect 391 902 392 903
rect 360 900 392 902
rect 360 899 361 900
rect 355 898 361 899
rect 391 899 392 900
rect 396 899 397 903
rect 391 898 397 899
rect 411 903 417 904
rect 411 899 412 903
rect 416 902 417 903
rect 459 903 465 904
rect 416 900 454 902
rect 416 899 417 900
rect 411 898 417 899
rect 452 894 454 900
rect 459 899 460 903
rect 464 902 465 903
rect 470 903 476 904
rect 470 902 471 903
rect 464 900 471 902
rect 464 899 465 900
rect 459 898 465 899
rect 470 899 471 900
rect 475 899 476 903
rect 470 898 476 899
rect 502 903 508 904
rect 502 899 503 903
rect 507 902 508 903
rect 515 903 521 904
rect 515 902 516 903
rect 507 900 516 902
rect 507 899 508 900
rect 502 898 508 899
rect 515 899 516 900
rect 520 899 521 903
rect 515 898 521 899
rect 558 903 564 904
rect 558 899 559 903
rect 563 902 564 903
rect 571 903 577 904
rect 571 902 572 903
rect 563 900 572 902
rect 563 899 564 900
rect 558 898 564 899
rect 571 899 572 900
rect 576 899 577 903
rect 571 898 577 899
rect 630 903 641 904
rect 630 899 631 903
rect 635 899 636 903
rect 640 899 641 903
rect 630 898 641 899
rect 702 903 713 904
rect 702 899 703 903
rect 707 899 708 903
rect 712 899 713 903
rect 702 898 713 899
rect 774 903 785 904
rect 774 899 775 903
rect 779 899 780 903
rect 784 899 785 903
rect 774 898 785 899
rect 846 903 857 904
rect 846 899 847 903
rect 851 899 852 903
rect 856 899 857 903
rect 846 898 857 899
rect 923 903 929 904
rect 923 899 924 903
rect 928 902 929 903
rect 938 903 944 904
rect 938 902 939 903
rect 928 900 939 902
rect 928 899 929 900
rect 923 898 929 899
rect 938 899 939 900
rect 943 899 944 903
rect 938 898 944 899
rect 990 903 1001 904
rect 990 899 991 903
rect 995 899 996 903
rect 1000 899 1001 903
rect 990 898 1001 899
rect 1067 903 1073 904
rect 1067 899 1068 903
rect 1072 902 1073 903
rect 1103 903 1109 904
rect 1103 902 1104 903
rect 1072 900 1104 902
rect 1072 899 1073 900
rect 1067 898 1073 899
rect 1103 899 1104 900
rect 1108 899 1109 903
rect 1103 898 1109 899
rect 1139 903 1145 904
rect 1139 899 1140 903
rect 1144 902 1145 903
rect 1150 903 1156 904
rect 1150 902 1151 903
rect 1144 900 1151 902
rect 1144 899 1145 900
rect 1139 898 1145 899
rect 1150 899 1151 900
rect 1155 899 1156 903
rect 1150 898 1156 899
rect 1187 903 1193 904
rect 1187 899 1188 903
rect 1192 902 1193 903
rect 1286 903 1292 904
rect 1286 902 1287 903
rect 1192 900 1287 902
rect 1192 899 1193 900
rect 1187 898 1193 899
rect 1286 899 1287 900
rect 1291 899 1292 903
rect 1286 898 1292 899
rect 1299 899 1305 900
rect 662 895 668 896
rect 662 894 663 895
rect 452 892 663 894
rect 274 891 280 892
rect 274 890 275 891
rect 188 888 275 890
rect 188 886 190 888
rect 274 887 275 888
rect 279 887 280 891
rect 662 891 663 892
rect 667 891 668 895
rect 1299 895 1300 899
rect 1304 898 1305 899
rect 1335 899 1341 900
rect 1335 898 1336 899
rect 1304 896 1336 898
rect 1304 895 1305 896
rect 1299 894 1305 895
rect 1335 895 1336 896
rect 1340 895 1341 899
rect 1335 894 1341 895
rect 1347 899 1353 900
rect 1347 895 1348 899
rect 1352 898 1353 899
rect 1383 899 1389 900
rect 1383 898 1384 899
rect 1352 896 1384 898
rect 1352 895 1353 896
rect 1347 894 1353 895
rect 1383 895 1384 896
rect 1388 895 1389 899
rect 1383 894 1389 895
rect 1427 899 1433 900
rect 1427 895 1428 899
rect 1432 898 1433 899
rect 1463 899 1469 900
rect 1463 898 1464 899
rect 1432 896 1464 898
rect 1432 895 1433 896
rect 1427 894 1433 895
rect 1463 895 1464 896
rect 1468 895 1469 899
rect 1463 894 1469 895
rect 1507 899 1513 900
rect 1507 895 1508 899
rect 1512 898 1513 899
rect 1570 899 1576 900
rect 1570 898 1571 899
rect 1512 896 1571 898
rect 1512 895 1513 896
rect 1507 894 1513 895
rect 1570 895 1571 896
rect 1575 895 1576 899
rect 1570 894 1576 895
rect 1587 899 1593 900
rect 1587 895 1588 899
rect 1592 898 1593 899
rect 1655 899 1661 900
rect 1655 898 1656 899
rect 1592 896 1656 898
rect 1592 895 1593 896
rect 1587 894 1593 895
rect 1655 895 1656 896
rect 1660 895 1661 899
rect 1655 894 1661 895
rect 1675 899 1681 900
rect 1675 895 1676 899
rect 1680 898 1681 899
rect 1686 899 1692 900
rect 1686 898 1687 899
rect 1680 896 1687 898
rect 1680 895 1681 896
rect 1675 894 1681 895
rect 1686 895 1687 896
rect 1691 895 1692 899
rect 1686 894 1692 895
rect 1763 899 1769 900
rect 1763 895 1764 899
rect 1768 898 1769 899
rect 1799 899 1805 900
rect 1799 898 1800 899
rect 1768 896 1800 898
rect 1768 895 1769 896
rect 1763 894 1769 895
rect 1799 895 1800 896
rect 1804 895 1805 899
rect 1799 894 1805 895
rect 1851 899 1857 900
rect 1851 895 1852 899
rect 1856 898 1857 899
rect 1887 899 1893 900
rect 1887 898 1888 899
rect 1856 896 1888 898
rect 1856 895 1857 896
rect 1851 894 1857 895
rect 1887 895 1888 896
rect 1892 895 1893 899
rect 1887 894 1893 895
rect 1939 899 1945 900
rect 1939 895 1940 899
rect 1944 898 1945 899
rect 1991 899 1997 900
rect 1991 898 1992 899
rect 1944 896 1992 898
rect 1944 895 1945 896
rect 1939 894 1945 895
rect 1991 895 1992 896
rect 1996 895 1997 899
rect 1991 894 1997 895
rect 2019 899 2025 900
rect 2019 895 2020 899
rect 2024 898 2025 899
rect 2086 899 2092 900
rect 2086 898 2087 899
rect 2024 896 2087 898
rect 2024 895 2025 896
rect 2019 894 2025 895
rect 2086 895 2087 896
rect 2091 895 2092 899
rect 2086 894 2092 895
rect 2094 899 2105 900
rect 2094 895 2095 899
rect 2099 895 2100 899
rect 2104 895 2105 899
rect 2094 894 2105 895
rect 2179 899 2185 900
rect 2179 895 2180 899
rect 2184 898 2185 899
rect 2190 899 2196 900
rect 2190 898 2191 899
rect 2184 896 2191 898
rect 2184 895 2185 896
rect 2179 894 2185 895
rect 2190 895 2191 896
rect 2195 895 2196 899
rect 2190 894 2196 895
rect 2262 899 2273 900
rect 2262 895 2263 899
rect 2267 895 2268 899
rect 2272 895 2273 899
rect 2262 894 2273 895
rect 662 890 668 891
rect 274 886 280 887
rect 1435 887 1441 888
rect 187 885 193 886
rect 187 881 188 885
rect 192 881 193 885
rect 227 883 233 884
rect 227 882 228 883
rect 187 880 193 881
rect 216 880 228 882
rect 214 879 220 880
rect 190 875 196 876
rect 190 871 191 875
rect 195 871 196 875
rect 214 875 215 879
rect 219 875 220 879
rect 227 879 228 880
rect 232 879 233 883
rect 283 883 289 884
rect 283 882 284 883
rect 256 880 284 882
rect 227 878 233 879
rect 254 879 260 880
rect 214 874 220 875
rect 230 875 236 876
rect 190 870 196 871
rect 230 871 231 875
rect 235 871 236 875
rect 254 875 255 879
rect 259 875 260 879
rect 283 879 284 880
rect 288 879 289 883
rect 283 878 289 879
rect 335 883 341 884
rect 335 879 336 883
rect 340 882 341 883
rect 355 883 361 884
rect 355 882 356 883
rect 340 880 356 882
rect 340 879 341 880
rect 335 878 341 879
rect 355 879 356 880
rect 360 879 361 883
rect 355 878 361 879
rect 386 883 392 884
rect 386 879 387 883
rect 391 882 392 883
rect 443 883 449 884
rect 443 882 444 883
rect 391 880 444 882
rect 391 879 392 880
rect 386 878 392 879
rect 443 879 444 880
rect 448 879 449 883
rect 443 878 449 879
rect 498 883 504 884
rect 498 879 499 883
rect 503 882 504 883
rect 539 883 545 884
rect 539 882 540 883
rect 503 880 540 882
rect 503 879 504 880
rect 498 878 504 879
rect 539 879 540 880
rect 544 879 545 883
rect 539 878 545 879
rect 602 883 608 884
rect 602 879 603 883
rect 607 882 608 883
rect 635 883 641 884
rect 635 882 636 883
rect 607 880 636 882
rect 607 879 608 880
rect 602 878 608 879
rect 635 879 636 880
rect 640 879 641 883
rect 635 878 641 879
rect 723 883 729 884
rect 723 879 724 883
rect 728 882 729 883
rect 746 883 752 884
rect 746 882 747 883
rect 728 880 747 882
rect 728 879 729 880
rect 723 878 729 879
rect 746 879 747 880
rect 751 879 752 883
rect 746 878 752 879
rect 754 883 760 884
rect 754 879 755 883
rect 759 882 760 883
rect 803 883 809 884
rect 803 882 804 883
rect 759 880 804 882
rect 759 879 760 880
rect 754 878 760 879
rect 803 879 804 880
rect 808 879 809 883
rect 803 878 809 879
rect 883 883 889 884
rect 883 879 884 883
rect 888 882 889 883
rect 946 883 952 884
rect 946 882 947 883
rect 888 880 947 882
rect 888 879 889 880
rect 883 878 889 879
rect 946 879 947 880
rect 951 879 952 883
rect 946 878 952 879
rect 955 883 961 884
rect 955 879 956 883
rect 960 882 961 883
rect 1006 883 1012 884
rect 1006 882 1007 883
rect 960 880 1007 882
rect 960 879 961 880
rect 955 878 961 879
rect 1006 879 1007 880
rect 1011 879 1012 883
rect 1006 878 1012 879
rect 1014 883 1025 884
rect 1014 879 1015 883
rect 1019 879 1020 883
rect 1024 879 1025 883
rect 1014 878 1025 879
rect 1050 883 1056 884
rect 1050 879 1051 883
rect 1055 882 1056 883
rect 1083 883 1089 884
rect 1083 882 1084 883
rect 1055 880 1084 882
rect 1055 879 1056 880
rect 1050 878 1056 879
rect 1083 879 1084 880
rect 1088 879 1089 883
rect 1083 878 1089 879
rect 1114 883 1120 884
rect 1114 879 1115 883
rect 1119 882 1120 883
rect 1155 883 1161 884
rect 1155 882 1156 883
rect 1119 880 1156 882
rect 1119 879 1120 880
rect 1114 878 1120 879
rect 1155 879 1156 880
rect 1160 879 1161 883
rect 1435 883 1436 887
rect 1440 886 1441 887
rect 1454 887 1460 888
rect 1454 886 1455 887
rect 1440 884 1455 886
rect 1440 883 1441 884
rect 1435 882 1441 883
rect 1454 883 1455 884
rect 1459 883 1460 887
rect 1454 882 1460 883
rect 1462 887 1468 888
rect 1462 883 1463 887
rect 1467 886 1468 887
rect 1475 887 1481 888
rect 1475 886 1476 887
rect 1467 884 1476 886
rect 1467 883 1468 884
rect 1462 882 1468 883
rect 1475 883 1476 884
rect 1480 883 1481 887
rect 1475 882 1481 883
rect 1502 887 1508 888
rect 1502 883 1503 887
rect 1507 886 1508 887
rect 1515 887 1521 888
rect 1515 886 1516 887
rect 1507 884 1516 886
rect 1507 883 1508 884
rect 1502 882 1508 883
rect 1515 883 1516 884
rect 1520 883 1521 887
rect 1515 882 1521 883
rect 1546 887 1552 888
rect 1546 883 1547 887
rect 1551 886 1552 887
rect 1555 887 1561 888
rect 1555 886 1556 887
rect 1551 884 1556 886
rect 1551 883 1552 884
rect 1546 882 1552 883
rect 1555 883 1556 884
rect 1560 883 1561 887
rect 1555 882 1561 883
rect 1591 887 1597 888
rect 1591 883 1592 887
rect 1596 886 1597 887
rect 1603 887 1609 888
rect 1603 886 1604 887
rect 1596 884 1604 886
rect 1596 883 1597 884
rect 1591 882 1597 883
rect 1603 883 1604 884
rect 1608 883 1609 887
rect 1603 882 1609 883
rect 1646 887 1657 888
rect 1646 883 1647 887
rect 1651 883 1652 887
rect 1656 883 1657 887
rect 1646 882 1657 883
rect 1687 887 1693 888
rect 1687 883 1688 887
rect 1692 886 1693 887
rect 1707 887 1713 888
rect 1707 886 1708 887
rect 1692 884 1708 886
rect 1692 883 1693 884
rect 1687 882 1693 883
rect 1707 883 1708 884
rect 1712 883 1713 887
rect 1707 882 1713 883
rect 1771 887 1777 888
rect 1771 883 1772 887
rect 1776 886 1777 887
rect 1782 887 1788 888
rect 1782 886 1783 887
rect 1776 884 1783 886
rect 1776 883 1777 884
rect 1771 882 1777 883
rect 1782 883 1783 884
rect 1787 883 1788 887
rect 1782 882 1788 883
rect 1802 887 1808 888
rect 1802 883 1803 887
rect 1807 886 1808 887
rect 1843 887 1849 888
rect 1843 886 1844 887
rect 1807 884 1844 886
rect 1807 883 1808 884
rect 1802 882 1808 883
rect 1843 883 1844 884
rect 1848 883 1849 887
rect 1843 882 1849 883
rect 1874 887 1880 888
rect 1874 883 1875 887
rect 1879 886 1880 887
rect 1915 887 1921 888
rect 1915 886 1916 887
rect 1879 884 1916 886
rect 1879 883 1880 884
rect 1874 882 1880 883
rect 1915 883 1916 884
rect 1920 883 1921 887
rect 1915 882 1921 883
rect 1967 887 1973 888
rect 1967 883 1968 887
rect 1972 886 1973 887
rect 1987 887 1993 888
rect 1987 886 1988 887
rect 1972 884 1988 886
rect 1972 883 1973 884
rect 1967 882 1973 883
rect 1987 883 1988 884
rect 1992 883 1993 887
rect 1987 882 1993 883
rect 2059 887 2065 888
rect 2059 883 2060 887
rect 2064 886 2065 887
rect 2110 887 2116 888
rect 2110 886 2111 887
rect 2064 884 2111 886
rect 2064 883 2065 884
rect 2059 882 2065 883
rect 2110 883 2111 884
rect 2115 883 2116 887
rect 2110 882 2116 883
rect 2131 887 2137 888
rect 2131 883 2132 887
rect 2136 886 2137 887
rect 2202 887 2208 888
rect 2202 886 2203 887
rect 2136 884 2203 886
rect 2136 883 2137 884
rect 2131 882 2137 883
rect 2202 883 2203 884
rect 2207 883 2208 887
rect 2202 882 2208 883
rect 2211 887 2217 888
rect 2211 883 2212 887
rect 2216 886 2217 887
rect 2278 887 2284 888
rect 2278 886 2279 887
rect 2216 884 2279 886
rect 2216 883 2217 884
rect 2211 882 2217 883
rect 2278 883 2279 884
rect 2283 883 2284 887
rect 2278 882 2284 883
rect 2286 887 2297 888
rect 2286 883 2287 887
rect 2291 883 2292 887
rect 2296 883 2297 887
rect 2286 882 2297 883
rect 1155 878 1161 879
rect 1438 879 1444 880
rect 254 874 260 875
rect 286 875 292 876
rect 230 870 236 871
rect 286 871 287 875
rect 291 871 292 875
rect 286 870 292 871
rect 358 875 364 876
rect 358 871 359 875
rect 363 871 364 875
rect 358 870 364 871
rect 446 875 452 876
rect 446 871 447 875
rect 451 871 452 875
rect 446 870 452 871
rect 542 875 548 876
rect 542 871 543 875
rect 547 871 548 875
rect 542 870 548 871
rect 638 875 644 876
rect 638 871 639 875
rect 643 871 644 875
rect 638 870 644 871
rect 726 875 732 876
rect 726 871 727 875
rect 731 871 732 875
rect 726 870 732 871
rect 806 875 812 876
rect 806 871 807 875
rect 811 871 812 875
rect 806 870 812 871
rect 886 875 892 876
rect 886 871 887 875
rect 891 871 892 875
rect 886 870 892 871
rect 958 875 964 876
rect 958 871 959 875
rect 963 871 964 875
rect 958 870 964 871
rect 1022 875 1028 876
rect 1022 871 1023 875
rect 1027 871 1028 875
rect 1022 870 1028 871
rect 1086 875 1092 876
rect 1086 871 1087 875
rect 1091 871 1092 875
rect 1086 870 1092 871
rect 1158 875 1164 876
rect 1158 871 1159 875
rect 1163 871 1164 875
rect 1438 875 1439 879
rect 1443 875 1444 879
rect 1438 874 1444 875
rect 1478 879 1484 880
rect 1478 875 1479 879
rect 1483 875 1484 879
rect 1478 874 1484 875
rect 1518 879 1524 880
rect 1518 875 1519 879
rect 1523 875 1524 879
rect 1518 874 1524 875
rect 1558 879 1564 880
rect 1558 875 1559 879
rect 1563 875 1564 879
rect 1558 874 1564 875
rect 1606 879 1612 880
rect 1606 875 1607 879
rect 1611 875 1612 879
rect 1606 874 1612 875
rect 1654 879 1660 880
rect 1654 875 1655 879
rect 1659 875 1660 879
rect 1654 874 1660 875
rect 1710 879 1716 880
rect 1710 875 1711 879
rect 1715 875 1716 879
rect 1710 874 1716 875
rect 1774 879 1780 880
rect 1774 875 1775 879
rect 1779 875 1780 879
rect 1774 874 1780 875
rect 1846 879 1852 880
rect 1846 875 1847 879
rect 1851 875 1852 879
rect 1846 874 1852 875
rect 1918 879 1924 880
rect 1918 875 1919 879
rect 1923 875 1924 879
rect 1918 874 1924 875
rect 1990 879 1996 880
rect 1990 875 1991 879
rect 1995 875 1996 879
rect 1990 874 1996 875
rect 2062 879 2068 880
rect 2062 875 2063 879
rect 2067 875 2068 879
rect 2062 874 2068 875
rect 2134 879 2140 880
rect 2134 875 2135 879
rect 2139 875 2140 879
rect 2134 874 2140 875
rect 2214 879 2220 880
rect 2214 875 2215 879
rect 2219 875 2220 879
rect 2214 874 2220 875
rect 2294 879 2300 880
rect 2294 875 2295 879
rect 2299 875 2300 879
rect 2294 874 2300 875
rect 1158 870 1164 871
rect 1570 859 1576 860
rect 1278 856 1284 857
rect 746 855 752 856
rect 110 852 116 853
rect 110 848 111 852
rect 115 848 116 852
rect 746 851 747 855
rect 751 854 752 855
rect 1006 855 1012 856
rect 751 852 882 854
rect 751 851 752 852
rect 746 850 752 851
rect 110 847 116 848
rect 214 847 221 848
rect 214 843 215 847
rect 220 843 221 847
rect 214 842 221 843
rect 254 847 261 848
rect 254 843 255 847
rect 260 843 261 847
rect 254 842 261 843
rect 311 847 317 848
rect 311 843 312 847
rect 316 846 317 847
rect 335 847 341 848
rect 335 846 336 847
rect 316 844 336 846
rect 316 843 317 844
rect 311 842 317 843
rect 335 843 336 844
rect 340 843 341 847
rect 335 842 341 843
rect 383 847 392 848
rect 383 843 384 847
rect 391 843 392 847
rect 383 842 392 843
rect 471 847 477 848
rect 471 843 472 847
rect 476 846 477 847
rect 498 847 504 848
rect 498 846 499 847
rect 476 844 499 846
rect 476 843 477 844
rect 471 842 477 843
rect 498 843 499 844
rect 503 843 504 847
rect 498 842 504 843
rect 567 847 573 848
rect 567 843 568 847
rect 572 846 573 847
rect 602 847 608 848
rect 602 846 603 847
rect 572 844 603 846
rect 572 843 573 844
rect 567 842 573 843
rect 602 843 603 844
rect 607 843 608 847
rect 602 842 608 843
rect 662 847 669 848
rect 662 843 663 847
rect 668 843 669 847
rect 662 842 669 843
rect 751 847 760 848
rect 751 843 752 847
rect 759 843 760 847
rect 751 842 760 843
rect 831 847 837 848
rect 831 843 832 847
rect 836 846 837 847
rect 870 847 876 848
rect 870 846 871 847
rect 836 844 871 846
rect 836 843 837 844
rect 831 842 837 843
rect 870 843 871 844
rect 875 843 876 847
rect 880 846 882 852
rect 1006 851 1007 855
rect 1011 854 1012 855
rect 1011 852 1161 854
rect 1011 851 1012 852
rect 1006 850 1012 851
rect 911 847 917 848
rect 911 846 912 847
rect 880 844 912 846
rect 870 842 876 843
rect 911 843 912 844
rect 916 843 917 847
rect 911 842 917 843
rect 946 847 952 848
rect 946 843 947 847
rect 951 846 952 847
rect 983 847 989 848
rect 983 846 984 847
rect 951 844 984 846
rect 951 843 952 844
rect 946 842 952 843
rect 983 843 984 844
rect 988 843 989 847
rect 983 842 989 843
rect 1047 847 1056 848
rect 1047 843 1048 847
rect 1055 843 1056 847
rect 1047 842 1056 843
rect 1111 847 1120 848
rect 1111 843 1112 847
rect 1119 843 1120 847
rect 1159 846 1161 852
rect 1238 852 1244 853
rect 1238 848 1239 852
rect 1243 848 1244 852
rect 1278 852 1279 856
rect 1283 852 1284 856
rect 1570 855 1571 859
rect 1575 858 1576 859
rect 1575 856 1602 858
rect 2406 856 2412 857
rect 1575 855 1576 856
rect 1570 854 1576 855
rect 1278 851 1284 852
rect 1462 851 1469 852
rect 1183 847 1189 848
rect 1238 847 1244 848
rect 1462 847 1463 851
rect 1468 847 1469 851
rect 1183 846 1184 847
rect 1159 844 1184 846
rect 1111 842 1120 843
rect 1183 843 1184 844
rect 1188 843 1189 847
rect 1462 846 1469 847
rect 1502 851 1509 852
rect 1502 847 1503 851
rect 1508 847 1509 851
rect 1502 846 1509 847
rect 1543 851 1552 852
rect 1543 847 1544 851
rect 1551 847 1552 851
rect 1543 846 1552 847
rect 1583 851 1589 852
rect 1583 847 1584 851
rect 1588 850 1589 851
rect 1591 851 1597 852
rect 1591 850 1592 851
rect 1588 848 1592 850
rect 1588 847 1589 848
rect 1583 846 1589 847
rect 1591 847 1592 848
rect 1596 847 1597 851
rect 1600 850 1602 856
rect 1687 855 1693 856
rect 1687 854 1688 855
rect 1679 853 1688 854
rect 1631 851 1637 852
rect 1631 850 1632 851
rect 1600 848 1632 850
rect 1591 846 1597 847
rect 1631 847 1632 848
rect 1636 847 1637 851
rect 1679 849 1680 853
rect 1684 852 1688 853
rect 1684 849 1685 852
rect 1687 851 1688 852
rect 1692 851 1693 855
rect 1967 855 1973 856
rect 1967 854 1968 855
rect 1943 853 1968 854
rect 1687 850 1693 851
rect 1718 851 1724 852
rect 1679 848 1685 849
rect 1631 846 1637 847
rect 1718 847 1719 851
rect 1723 850 1724 851
rect 1735 851 1741 852
rect 1735 850 1736 851
rect 1723 848 1736 850
rect 1723 847 1724 848
rect 1718 846 1724 847
rect 1735 847 1736 848
rect 1740 847 1741 851
rect 1735 846 1741 847
rect 1799 851 1808 852
rect 1799 847 1800 851
rect 1807 847 1808 851
rect 1799 846 1808 847
rect 1871 851 1880 852
rect 1871 847 1872 851
rect 1879 847 1880 851
rect 1943 849 1944 853
rect 1948 852 1968 853
rect 1948 849 1949 852
rect 1967 851 1968 852
rect 1972 851 1973 855
rect 2406 852 2407 856
rect 2411 852 2412 856
rect 1967 850 1973 851
rect 2015 851 2021 852
rect 2015 850 2016 851
rect 1943 848 1949 849
rect 1999 848 2016 850
rect 1871 846 1880 847
rect 1183 842 1189 843
rect 1766 843 1772 844
rect 1278 839 1284 840
rect 110 835 116 836
rect 110 831 111 835
rect 115 831 116 835
rect 110 830 116 831
rect 1238 835 1244 836
rect 1238 831 1239 835
rect 1243 831 1244 835
rect 1278 835 1279 839
rect 1283 835 1284 839
rect 1766 839 1767 843
rect 1771 842 1772 843
rect 1999 842 2001 848
rect 2015 847 2016 848
rect 2020 847 2021 851
rect 2015 846 2021 847
rect 2086 851 2093 852
rect 2086 847 2087 851
rect 2092 847 2093 851
rect 2086 846 2093 847
rect 2110 851 2116 852
rect 2110 847 2111 851
rect 2115 850 2116 851
rect 2159 851 2165 852
rect 2159 850 2160 851
rect 2115 848 2160 850
rect 2115 847 2116 848
rect 2110 846 2116 847
rect 2159 847 2160 848
rect 2164 847 2165 851
rect 2159 846 2165 847
rect 2202 851 2208 852
rect 2202 847 2203 851
rect 2207 850 2208 851
rect 2239 851 2245 852
rect 2239 850 2240 851
rect 2207 848 2240 850
rect 2207 847 2208 848
rect 2202 846 2208 847
rect 2239 847 2240 848
rect 2244 847 2245 851
rect 2239 846 2245 847
rect 2278 851 2284 852
rect 2278 847 2279 851
rect 2283 850 2284 851
rect 2319 851 2325 852
rect 2406 851 2412 852
rect 2319 850 2320 851
rect 2283 848 2320 850
rect 2283 847 2284 848
rect 2278 846 2284 847
rect 2319 847 2320 848
rect 2324 847 2325 851
rect 2319 846 2325 847
rect 1771 840 2001 842
rect 1771 839 1772 840
rect 1766 838 1772 839
rect 2406 839 2412 840
rect 1278 834 1284 835
rect 2406 835 2407 839
rect 2411 835 2412 839
rect 2406 834 2412 835
rect 1238 830 1244 831
rect 1438 832 1444 833
rect 190 828 196 829
rect 190 824 191 828
rect 195 824 196 828
rect 190 823 196 824
rect 230 828 236 829
rect 230 824 231 828
rect 235 824 236 828
rect 230 823 236 824
rect 286 828 292 829
rect 286 824 287 828
rect 291 824 292 828
rect 286 823 292 824
rect 358 828 364 829
rect 358 824 359 828
rect 363 824 364 828
rect 358 823 364 824
rect 446 828 452 829
rect 446 824 447 828
rect 451 824 452 828
rect 446 823 452 824
rect 542 828 548 829
rect 542 824 543 828
rect 547 824 548 828
rect 542 823 548 824
rect 638 828 644 829
rect 638 824 639 828
rect 643 824 644 828
rect 638 823 644 824
rect 726 828 732 829
rect 726 824 727 828
rect 731 824 732 828
rect 726 823 732 824
rect 806 828 812 829
rect 806 824 807 828
rect 811 824 812 828
rect 806 823 812 824
rect 886 828 892 829
rect 886 824 887 828
rect 891 824 892 828
rect 886 823 892 824
rect 958 828 964 829
rect 958 824 959 828
rect 963 824 964 828
rect 958 823 964 824
rect 1022 828 1028 829
rect 1022 824 1023 828
rect 1027 824 1028 828
rect 1022 823 1028 824
rect 1086 828 1092 829
rect 1086 824 1087 828
rect 1091 824 1092 828
rect 1086 823 1092 824
rect 1158 828 1164 829
rect 1158 824 1159 828
rect 1163 824 1164 828
rect 1438 828 1439 832
rect 1443 828 1444 832
rect 1438 827 1444 828
rect 1478 832 1484 833
rect 1478 828 1479 832
rect 1483 828 1484 832
rect 1478 827 1484 828
rect 1518 832 1524 833
rect 1518 828 1519 832
rect 1523 828 1524 832
rect 1518 827 1524 828
rect 1558 832 1564 833
rect 1558 828 1559 832
rect 1563 828 1564 832
rect 1558 827 1564 828
rect 1606 832 1612 833
rect 1606 828 1607 832
rect 1611 828 1612 832
rect 1606 827 1612 828
rect 1654 832 1660 833
rect 1654 828 1655 832
rect 1659 828 1660 832
rect 1654 827 1660 828
rect 1710 832 1716 833
rect 1710 828 1711 832
rect 1715 828 1716 832
rect 1710 827 1716 828
rect 1774 832 1780 833
rect 1774 828 1775 832
rect 1779 828 1780 832
rect 1774 827 1780 828
rect 1846 832 1852 833
rect 1846 828 1847 832
rect 1851 828 1852 832
rect 1846 827 1852 828
rect 1918 832 1924 833
rect 1918 828 1919 832
rect 1923 828 1924 832
rect 1918 827 1924 828
rect 1990 832 1996 833
rect 1990 828 1991 832
rect 1995 828 1996 832
rect 1990 827 1996 828
rect 2062 832 2068 833
rect 2062 828 2063 832
rect 2067 828 2068 832
rect 2062 827 2068 828
rect 2134 832 2140 833
rect 2134 828 2135 832
rect 2139 828 2140 832
rect 2134 827 2140 828
rect 2214 832 2220 833
rect 2214 828 2215 832
rect 2219 828 2220 832
rect 2214 827 2220 828
rect 2294 832 2300 833
rect 2294 828 2295 832
rect 2299 828 2300 832
rect 2294 827 2300 828
rect 1158 823 1164 824
rect 134 816 140 817
rect 134 812 135 816
rect 139 812 140 816
rect 134 811 140 812
rect 174 816 180 817
rect 174 812 175 816
rect 179 812 180 816
rect 174 811 180 812
rect 238 816 244 817
rect 238 812 239 816
rect 243 812 244 816
rect 238 811 244 812
rect 326 816 332 817
rect 326 812 327 816
rect 331 812 332 816
rect 326 811 332 812
rect 414 816 420 817
rect 414 812 415 816
rect 419 812 420 816
rect 414 811 420 812
rect 502 816 508 817
rect 502 812 503 816
rect 507 812 508 816
rect 502 811 508 812
rect 590 816 596 817
rect 590 812 591 816
rect 595 812 596 816
rect 590 811 596 812
rect 670 816 676 817
rect 670 812 671 816
rect 675 812 676 816
rect 670 811 676 812
rect 742 816 748 817
rect 742 812 743 816
rect 747 812 748 816
rect 742 811 748 812
rect 814 816 820 817
rect 814 812 815 816
rect 819 812 820 816
rect 814 811 820 812
rect 878 816 884 817
rect 878 812 879 816
rect 883 812 884 816
rect 878 811 884 812
rect 942 816 948 817
rect 942 812 943 816
rect 947 812 948 816
rect 942 811 948 812
rect 1014 816 1020 817
rect 1014 812 1015 816
rect 1019 812 1020 816
rect 1014 811 1020 812
rect 110 809 116 810
rect 110 805 111 809
rect 115 805 116 809
rect 110 804 116 805
rect 1238 809 1244 810
rect 1238 805 1239 809
rect 1243 805 1244 809
rect 1238 804 1244 805
rect 1358 808 1364 809
rect 1358 804 1359 808
rect 1363 804 1364 808
rect 274 803 280 804
rect 1358 803 1364 804
rect 1414 808 1420 809
rect 1414 804 1415 808
rect 1419 804 1420 808
rect 1414 803 1420 804
rect 1470 808 1476 809
rect 1470 804 1471 808
rect 1475 804 1476 808
rect 1470 803 1476 804
rect 1534 808 1540 809
rect 1534 804 1535 808
rect 1539 804 1540 808
rect 1534 803 1540 804
rect 1590 808 1596 809
rect 1590 804 1591 808
rect 1595 804 1596 808
rect 1590 803 1596 804
rect 1646 808 1652 809
rect 1646 804 1647 808
rect 1651 804 1652 808
rect 1646 803 1652 804
rect 1702 808 1708 809
rect 1702 804 1703 808
rect 1707 804 1708 808
rect 1702 803 1708 804
rect 1758 808 1764 809
rect 1758 804 1759 808
rect 1763 804 1764 808
rect 1758 803 1764 804
rect 1814 808 1820 809
rect 1814 804 1815 808
rect 1819 804 1820 808
rect 1814 803 1820 804
rect 1870 808 1876 809
rect 1870 804 1871 808
rect 1875 804 1876 808
rect 1870 803 1876 804
rect 1934 808 1940 809
rect 1934 804 1935 808
rect 1939 804 1940 808
rect 1934 803 1940 804
rect 1998 808 2004 809
rect 1998 804 1999 808
rect 2003 804 2004 808
rect 1998 803 2004 804
rect 2070 808 2076 809
rect 2070 804 2071 808
rect 2075 804 2076 808
rect 2070 803 2076 804
rect 2142 808 2148 809
rect 2142 804 2143 808
rect 2147 804 2148 808
rect 2142 803 2148 804
rect 2222 808 2228 809
rect 2222 804 2223 808
rect 2227 804 2228 808
rect 2222 803 2228 804
rect 2302 808 2308 809
rect 2302 804 2303 808
rect 2307 804 2308 808
rect 2302 803 2308 804
rect 2358 808 2364 809
rect 2358 804 2359 808
rect 2363 804 2364 808
rect 2358 803 2364 804
rect 274 799 275 803
rect 279 802 280 803
rect 279 800 506 802
rect 279 799 280 800
rect 274 798 280 799
rect 159 795 168 796
rect 110 792 116 793
rect 110 788 111 792
rect 115 788 116 792
rect 159 791 160 795
rect 167 791 168 795
rect 159 790 168 791
rect 199 795 205 796
rect 199 791 200 795
rect 204 794 205 795
rect 230 795 236 796
rect 230 794 231 795
rect 204 792 231 794
rect 204 791 205 792
rect 199 790 205 791
rect 230 791 231 792
rect 235 791 236 795
rect 230 790 236 791
rect 263 795 269 796
rect 263 791 264 795
rect 268 794 269 795
rect 318 795 324 796
rect 318 794 319 795
rect 268 792 319 794
rect 268 791 269 792
rect 263 790 269 791
rect 318 791 319 792
rect 323 791 324 795
rect 318 790 324 791
rect 351 795 357 796
rect 351 791 352 795
rect 356 794 357 795
rect 406 795 412 796
rect 406 794 407 795
rect 356 792 407 794
rect 356 791 357 792
rect 351 790 357 791
rect 406 791 407 792
rect 411 791 412 795
rect 406 790 412 791
rect 439 795 445 796
rect 439 791 440 795
rect 444 794 445 795
rect 494 795 500 796
rect 494 794 495 795
rect 444 792 495 794
rect 444 791 445 792
rect 439 790 445 791
rect 494 791 495 792
rect 499 791 500 795
rect 504 794 506 800
rect 1278 801 1284 802
rect 1278 797 1279 801
rect 1283 797 1284 801
rect 1278 796 1284 797
rect 2406 801 2412 802
rect 2406 797 2407 801
rect 2411 797 2412 801
rect 2406 796 2412 797
rect 527 795 533 796
rect 527 794 528 795
rect 504 792 528 794
rect 494 790 500 791
rect 527 791 528 792
rect 532 791 533 795
rect 527 790 533 791
rect 615 795 621 796
rect 615 791 616 795
rect 620 794 621 795
rect 662 795 668 796
rect 662 794 663 795
rect 620 792 663 794
rect 620 791 621 792
rect 615 790 621 791
rect 662 791 663 792
rect 667 791 668 795
rect 662 790 668 791
rect 695 795 701 796
rect 695 791 696 795
rect 700 794 701 795
rect 734 795 740 796
rect 734 794 735 795
rect 700 792 735 794
rect 700 791 701 792
rect 695 790 701 791
rect 734 791 735 792
rect 739 791 740 795
rect 734 790 740 791
rect 767 795 773 796
rect 767 791 768 795
rect 772 794 773 795
rect 806 795 812 796
rect 806 794 807 795
rect 772 792 807 794
rect 772 791 773 792
rect 767 790 773 791
rect 806 791 807 792
rect 811 791 812 795
rect 839 795 845 796
rect 839 794 840 795
rect 806 790 812 791
rect 816 792 840 794
rect 110 787 116 788
rect 606 787 612 788
rect 606 783 607 787
rect 611 786 612 787
rect 816 786 818 792
rect 839 791 840 792
rect 844 791 845 795
rect 839 790 845 791
rect 903 795 909 796
rect 903 791 904 795
rect 908 794 909 795
rect 934 795 940 796
rect 934 794 935 795
rect 908 792 935 794
rect 908 791 909 792
rect 903 790 909 791
rect 934 791 935 792
rect 939 791 940 795
rect 934 790 940 791
rect 967 795 973 796
rect 967 791 968 795
rect 972 794 973 795
rect 1006 795 1012 796
rect 1006 794 1007 795
rect 972 792 1007 794
rect 972 791 973 792
rect 967 790 973 791
rect 1006 791 1007 792
rect 1011 791 1012 795
rect 1039 795 1045 796
rect 1039 794 1040 795
rect 1006 790 1012 791
rect 1016 792 1040 794
rect 611 784 818 786
rect 822 787 828 788
rect 611 783 612 784
rect 606 782 612 783
rect 822 783 823 787
rect 827 786 828 787
rect 1016 786 1018 792
rect 1039 791 1040 792
rect 1044 791 1045 795
rect 1454 795 1460 796
rect 1039 790 1045 791
rect 1238 792 1244 793
rect 1238 788 1239 792
rect 1243 788 1244 792
rect 1454 791 1455 795
rect 1459 794 1460 795
rect 1459 792 1538 794
rect 1459 791 1460 792
rect 1454 790 1460 791
rect 1238 787 1244 788
rect 1383 787 1389 788
rect 827 784 1018 786
rect 1278 784 1284 785
rect 827 783 828 784
rect 822 782 828 783
rect 1278 780 1279 784
rect 1283 780 1284 784
rect 1383 783 1384 787
rect 1388 786 1389 787
rect 1398 787 1404 788
rect 1398 786 1399 787
rect 1388 784 1399 786
rect 1388 783 1389 784
rect 1383 782 1389 783
rect 1398 783 1399 784
rect 1403 783 1404 787
rect 1398 782 1404 783
rect 1439 787 1445 788
rect 1439 783 1440 787
rect 1444 786 1445 787
rect 1462 787 1468 788
rect 1462 786 1463 787
rect 1444 784 1463 786
rect 1444 783 1445 784
rect 1439 782 1445 783
rect 1462 783 1463 784
rect 1467 783 1468 787
rect 1462 782 1468 783
rect 1495 787 1501 788
rect 1495 783 1496 787
rect 1500 786 1501 787
rect 1526 787 1532 788
rect 1526 786 1527 787
rect 1500 784 1527 786
rect 1500 783 1501 784
rect 1495 782 1501 783
rect 1526 783 1527 784
rect 1531 783 1532 787
rect 1536 786 1538 792
rect 1559 787 1565 788
rect 1559 786 1560 787
rect 1536 784 1560 786
rect 1526 782 1532 783
rect 1559 783 1560 784
rect 1564 783 1565 787
rect 1559 782 1565 783
rect 1615 787 1621 788
rect 1615 783 1616 787
rect 1620 786 1621 787
rect 1638 787 1644 788
rect 1638 786 1639 787
rect 1620 784 1639 786
rect 1620 783 1621 784
rect 1615 782 1621 783
rect 1638 783 1639 784
rect 1643 783 1644 787
rect 1638 782 1644 783
rect 1670 787 1677 788
rect 1670 783 1671 787
rect 1676 783 1677 787
rect 1727 787 1733 788
rect 1727 786 1728 787
rect 1670 782 1677 783
rect 1680 784 1728 786
rect 1278 779 1284 780
rect 1598 779 1604 780
rect 1598 775 1599 779
rect 1603 778 1604 779
rect 1680 778 1682 784
rect 1727 783 1728 784
rect 1732 783 1733 787
rect 1727 782 1733 783
rect 1783 787 1789 788
rect 1783 783 1784 787
rect 1788 786 1789 787
rect 1798 787 1804 788
rect 1798 786 1799 787
rect 1788 784 1799 786
rect 1788 783 1789 784
rect 1783 782 1789 783
rect 1798 783 1799 784
rect 1803 783 1804 787
rect 1798 782 1804 783
rect 1839 787 1845 788
rect 1839 783 1840 787
rect 1844 786 1845 787
rect 1862 787 1868 788
rect 1862 786 1863 787
rect 1844 784 1863 786
rect 1844 783 1845 784
rect 1839 782 1845 783
rect 1862 783 1863 784
rect 1867 783 1868 787
rect 1862 782 1868 783
rect 1895 787 1901 788
rect 1895 783 1896 787
rect 1900 786 1901 787
rect 1926 787 1932 788
rect 1926 786 1927 787
rect 1900 784 1927 786
rect 1900 783 1901 784
rect 1895 782 1901 783
rect 1926 783 1927 784
rect 1931 783 1932 787
rect 1926 782 1932 783
rect 1959 787 1965 788
rect 1959 783 1960 787
rect 1964 786 1965 787
rect 1982 787 1988 788
rect 1982 786 1983 787
rect 1964 784 1983 786
rect 1964 783 1965 784
rect 1959 782 1965 783
rect 1982 783 1983 784
rect 1987 783 1988 787
rect 1982 782 1988 783
rect 2023 787 2029 788
rect 2023 783 2024 787
rect 2028 786 2029 787
rect 2062 787 2068 788
rect 2062 786 2063 787
rect 2028 784 2063 786
rect 2028 783 2029 784
rect 2023 782 2029 783
rect 2062 783 2063 784
rect 2067 783 2068 787
rect 2062 782 2068 783
rect 2095 787 2101 788
rect 2095 783 2096 787
rect 2100 786 2101 787
rect 2134 787 2140 788
rect 2134 786 2135 787
rect 2100 784 2135 786
rect 2100 783 2101 784
rect 2095 782 2101 783
rect 2134 783 2135 784
rect 2139 783 2140 787
rect 2134 782 2140 783
rect 2150 787 2156 788
rect 2150 783 2151 787
rect 2155 786 2156 787
rect 2167 787 2173 788
rect 2167 786 2168 787
rect 2155 784 2168 786
rect 2155 783 2156 784
rect 2150 782 2156 783
rect 2167 783 2168 784
rect 2172 783 2173 787
rect 2167 782 2173 783
rect 2247 787 2253 788
rect 2247 783 2248 787
rect 2252 786 2253 787
rect 2294 787 2300 788
rect 2294 786 2295 787
rect 2252 784 2295 786
rect 2252 783 2253 784
rect 2247 782 2253 783
rect 2294 783 2295 784
rect 2299 783 2300 787
rect 2294 782 2300 783
rect 2327 787 2333 788
rect 2327 783 2328 787
rect 2332 786 2333 787
rect 2350 787 2356 788
rect 2350 786 2351 787
rect 2332 784 2351 786
rect 2332 783 2333 784
rect 2327 782 2333 783
rect 2350 783 2351 784
rect 2355 783 2356 787
rect 2350 782 2356 783
rect 2370 787 2376 788
rect 2370 783 2371 787
rect 2375 786 2376 787
rect 2383 787 2389 788
rect 2383 786 2384 787
rect 2375 784 2384 786
rect 2375 783 2376 784
rect 2370 782 2376 783
rect 2383 783 2384 784
rect 2388 783 2389 787
rect 2383 782 2389 783
rect 2406 784 2412 785
rect 2406 780 2407 784
rect 2411 780 2412 784
rect 2406 779 2412 780
rect 1603 776 1682 778
rect 1603 775 1604 776
rect 1598 774 1604 775
rect 134 769 140 770
rect 134 765 135 769
rect 139 765 140 769
rect 134 764 140 765
rect 174 769 180 770
rect 174 765 175 769
rect 179 765 180 769
rect 174 764 180 765
rect 238 769 244 770
rect 238 765 239 769
rect 243 765 244 769
rect 238 764 244 765
rect 326 769 332 770
rect 326 765 327 769
rect 331 765 332 769
rect 326 764 332 765
rect 414 769 420 770
rect 414 765 415 769
rect 419 765 420 769
rect 414 764 420 765
rect 502 769 508 770
rect 502 765 503 769
rect 507 765 508 769
rect 502 764 508 765
rect 590 769 596 770
rect 590 765 591 769
rect 595 765 596 769
rect 590 764 596 765
rect 670 769 676 770
rect 670 765 671 769
rect 675 765 676 769
rect 670 764 676 765
rect 742 769 748 770
rect 742 765 743 769
rect 747 765 748 769
rect 742 764 748 765
rect 814 769 820 770
rect 814 765 815 769
rect 819 765 820 769
rect 814 764 820 765
rect 878 769 884 770
rect 878 765 879 769
rect 883 765 884 769
rect 878 764 884 765
rect 942 769 948 770
rect 942 765 943 769
rect 947 765 948 769
rect 942 764 948 765
rect 1014 769 1020 770
rect 1014 765 1015 769
rect 1019 765 1020 769
rect 1014 764 1020 765
rect 1358 761 1364 762
rect 131 759 137 760
rect 131 755 132 759
rect 136 758 137 759
rect 154 759 160 760
rect 154 758 155 759
rect 136 756 155 758
rect 136 755 137 756
rect 131 754 137 755
rect 154 755 155 756
rect 159 755 160 759
rect 154 754 160 755
rect 162 759 168 760
rect 162 755 163 759
rect 167 758 168 759
rect 171 759 177 760
rect 171 758 172 759
rect 167 756 172 758
rect 167 755 168 756
rect 162 754 168 755
rect 171 755 172 756
rect 176 755 177 759
rect 171 754 177 755
rect 230 759 241 760
rect 230 755 231 759
rect 235 755 236 759
rect 240 755 241 759
rect 230 754 241 755
rect 318 759 329 760
rect 318 755 319 759
rect 323 755 324 759
rect 328 755 329 759
rect 318 754 329 755
rect 406 759 417 760
rect 406 755 407 759
rect 411 755 412 759
rect 416 755 417 759
rect 406 754 417 755
rect 494 759 505 760
rect 494 755 495 759
rect 499 755 500 759
rect 504 755 505 759
rect 494 754 505 755
rect 587 759 593 760
rect 587 755 588 759
rect 592 758 593 759
rect 606 759 612 760
rect 606 758 607 759
rect 592 756 607 758
rect 592 755 593 756
rect 587 754 593 755
rect 606 755 607 756
rect 611 755 612 759
rect 606 754 612 755
rect 662 759 673 760
rect 662 755 663 759
rect 667 755 668 759
rect 672 755 673 759
rect 662 754 673 755
rect 734 759 745 760
rect 734 755 735 759
rect 739 755 740 759
rect 744 755 745 759
rect 734 754 745 755
rect 811 759 817 760
rect 811 755 812 759
rect 816 758 817 759
rect 822 759 828 760
rect 822 758 823 759
rect 816 756 823 758
rect 816 755 817 756
rect 811 754 817 755
rect 822 755 823 756
rect 827 755 828 759
rect 822 754 828 755
rect 870 759 881 760
rect 870 755 871 759
rect 875 755 876 759
rect 880 755 881 759
rect 870 754 881 755
rect 934 759 945 760
rect 934 755 935 759
rect 939 755 940 759
rect 944 755 945 759
rect 934 754 945 755
rect 1006 759 1017 760
rect 1006 755 1007 759
rect 1011 755 1012 759
rect 1016 755 1017 759
rect 1358 757 1359 761
rect 1363 757 1364 761
rect 1358 756 1364 757
rect 1414 761 1420 762
rect 1414 757 1415 761
rect 1419 757 1420 761
rect 1414 756 1420 757
rect 1470 761 1476 762
rect 1470 757 1471 761
rect 1475 757 1476 761
rect 1470 756 1476 757
rect 1534 761 1540 762
rect 1534 757 1535 761
rect 1539 757 1540 761
rect 1534 756 1540 757
rect 1590 761 1596 762
rect 1590 757 1591 761
rect 1595 757 1596 761
rect 1590 756 1596 757
rect 1646 761 1652 762
rect 1646 757 1647 761
rect 1651 757 1652 761
rect 1646 756 1652 757
rect 1702 761 1708 762
rect 1702 757 1703 761
rect 1707 757 1708 761
rect 1702 756 1708 757
rect 1758 761 1764 762
rect 1758 757 1759 761
rect 1763 757 1764 761
rect 1758 756 1764 757
rect 1814 761 1820 762
rect 1814 757 1815 761
rect 1819 757 1820 761
rect 1814 756 1820 757
rect 1870 761 1876 762
rect 1870 757 1871 761
rect 1875 757 1876 761
rect 1870 756 1876 757
rect 1934 761 1940 762
rect 1934 757 1935 761
rect 1939 757 1940 761
rect 1934 756 1940 757
rect 1998 761 2004 762
rect 1998 757 1999 761
rect 2003 757 2004 761
rect 1998 756 2004 757
rect 2070 761 2076 762
rect 2070 757 2071 761
rect 2075 757 2076 761
rect 2070 756 2076 757
rect 2142 761 2148 762
rect 2142 757 2143 761
rect 2147 757 2148 761
rect 2142 756 2148 757
rect 2222 761 2228 762
rect 2222 757 2223 761
rect 2227 757 2228 761
rect 2222 756 2228 757
rect 2302 761 2308 762
rect 2302 757 2303 761
rect 2307 757 2308 761
rect 2302 756 2308 757
rect 2358 761 2364 762
rect 2358 757 2359 761
rect 2363 757 2364 761
rect 2358 756 2364 757
rect 1006 754 1017 755
rect 1355 751 1361 752
rect 1355 747 1356 751
rect 1360 750 1361 751
rect 1390 751 1396 752
rect 1390 750 1391 751
rect 1360 748 1391 750
rect 1360 747 1361 748
rect 1355 746 1361 747
rect 1390 747 1391 748
rect 1395 747 1396 751
rect 1390 746 1396 747
rect 1398 751 1404 752
rect 1398 747 1399 751
rect 1403 750 1404 751
rect 1411 751 1417 752
rect 1411 750 1412 751
rect 1403 748 1412 750
rect 1403 747 1404 748
rect 1398 746 1404 747
rect 1411 747 1412 748
rect 1416 747 1417 751
rect 1411 746 1417 747
rect 1462 751 1473 752
rect 1462 747 1463 751
rect 1467 747 1468 751
rect 1472 747 1473 751
rect 1462 746 1473 747
rect 1526 751 1537 752
rect 1526 747 1527 751
rect 1531 747 1532 751
rect 1536 747 1537 751
rect 1526 746 1537 747
rect 1587 751 1593 752
rect 1587 747 1588 751
rect 1592 750 1593 751
rect 1598 751 1604 752
rect 1598 750 1599 751
rect 1592 748 1599 750
rect 1592 747 1593 748
rect 1587 746 1593 747
rect 1598 747 1599 748
rect 1603 747 1604 751
rect 1598 746 1604 747
rect 1638 751 1649 752
rect 1638 747 1639 751
rect 1643 747 1644 751
rect 1648 747 1649 751
rect 1638 746 1649 747
rect 1699 751 1705 752
rect 1699 747 1700 751
rect 1704 750 1705 751
rect 1718 751 1724 752
rect 1718 750 1719 751
rect 1704 748 1719 750
rect 1704 747 1705 748
rect 1699 746 1705 747
rect 1718 747 1719 748
rect 1723 747 1724 751
rect 1718 746 1724 747
rect 1755 751 1761 752
rect 1755 747 1756 751
rect 1760 750 1761 751
rect 1766 751 1772 752
rect 1766 750 1767 751
rect 1760 748 1767 750
rect 1760 747 1761 748
rect 1755 746 1761 747
rect 1766 747 1767 748
rect 1771 747 1772 751
rect 1766 746 1772 747
rect 1798 751 1804 752
rect 1798 747 1799 751
rect 1803 750 1804 751
rect 1811 751 1817 752
rect 1811 750 1812 751
rect 1803 748 1812 750
rect 1803 747 1804 748
rect 1798 746 1804 747
rect 1811 747 1812 748
rect 1816 747 1817 751
rect 1811 746 1817 747
rect 1862 751 1873 752
rect 1862 747 1863 751
rect 1867 747 1868 751
rect 1872 747 1873 751
rect 1862 746 1873 747
rect 1926 751 1937 752
rect 1926 747 1927 751
rect 1931 747 1932 751
rect 1936 747 1937 751
rect 1926 746 1937 747
rect 1982 751 1988 752
rect 1982 747 1983 751
rect 1987 750 1988 751
rect 1995 751 2001 752
rect 1995 750 1996 751
rect 1987 748 1996 750
rect 1987 747 1988 748
rect 1982 746 1988 747
rect 1995 747 1996 748
rect 2000 747 2001 751
rect 1995 746 2001 747
rect 2062 751 2073 752
rect 2062 747 2063 751
rect 2067 747 2068 751
rect 2072 747 2073 751
rect 2062 746 2073 747
rect 2134 751 2145 752
rect 2134 747 2135 751
rect 2139 747 2140 751
rect 2144 747 2145 751
rect 2134 746 2145 747
rect 2219 751 2225 752
rect 2219 747 2220 751
rect 2224 750 2225 751
rect 2286 751 2292 752
rect 2286 750 2287 751
rect 2224 748 2287 750
rect 2224 747 2225 748
rect 2219 746 2225 747
rect 2286 747 2287 748
rect 2291 747 2292 751
rect 2286 746 2292 747
rect 2294 751 2305 752
rect 2294 747 2295 751
rect 2299 747 2300 751
rect 2304 747 2305 751
rect 2294 746 2305 747
rect 2350 751 2361 752
rect 2350 747 2351 751
rect 2355 747 2356 751
rect 2360 747 2361 751
rect 2350 746 2361 747
rect 131 743 137 744
rect 131 739 132 743
rect 136 742 137 743
rect 175 743 181 744
rect 175 742 176 743
rect 136 740 176 742
rect 136 739 137 740
rect 131 738 137 739
rect 175 739 176 740
rect 180 739 181 743
rect 175 738 181 739
rect 187 743 193 744
rect 187 739 188 743
rect 192 742 193 743
rect 222 743 228 744
rect 222 742 223 743
rect 192 740 223 742
rect 192 739 193 740
rect 187 738 193 739
rect 222 739 223 740
rect 227 739 228 743
rect 222 738 228 739
rect 259 743 265 744
rect 259 739 260 743
rect 264 742 265 743
rect 319 743 325 744
rect 319 742 320 743
rect 264 740 320 742
rect 264 739 265 740
rect 259 738 265 739
rect 319 739 320 740
rect 324 739 325 743
rect 319 738 325 739
rect 331 743 337 744
rect 331 739 332 743
rect 336 742 337 743
rect 386 743 392 744
rect 386 742 387 743
rect 336 740 387 742
rect 336 739 337 740
rect 331 738 337 739
rect 386 739 387 740
rect 391 739 392 743
rect 386 738 392 739
rect 395 743 401 744
rect 395 739 396 743
rect 400 742 401 743
rect 442 743 448 744
rect 442 742 443 743
rect 400 740 443 742
rect 400 739 401 740
rect 395 738 401 739
rect 442 739 443 740
rect 447 739 448 743
rect 442 738 448 739
rect 451 743 457 744
rect 451 739 452 743
rect 456 742 457 743
rect 490 743 496 744
rect 490 742 491 743
rect 456 740 491 742
rect 456 739 457 740
rect 451 738 457 739
rect 490 739 491 740
rect 495 739 496 743
rect 490 738 496 739
rect 499 743 505 744
rect 499 739 500 743
rect 504 742 505 743
rect 530 743 536 744
rect 530 742 531 743
rect 504 740 531 742
rect 504 739 505 740
rect 499 738 505 739
rect 530 739 531 740
rect 535 739 536 743
rect 530 738 536 739
rect 539 743 545 744
rect 539 739 540 743
rect 544 742 545 743
rect 570 743 576 744
rect 570 742 571 743
rect 544 740 571 742
rect 544 739 545 740
rect 539 738 545 739
rect 570 739 571 740
rect 575 739 576 743
rect 570 738 576 739
rect 579 743 585 744
rect 579 739 580 743
rect 584 742 585 743
rect 610 743 616 744
rect 610 742 611 743
rect 584 740 611 742
rect 584 739 585 740
rect 579 738 585 739
rect 610 739 611 740
rect 615 739 616 743
rect 610 738 616 739
rect 619 743 625 744
rect 619 739 620 743
rect 624 742 625 743
rect 658 743 664 744
rect 658 742 659 743
rect 624 740 659 742
rect 624 739 625 740
rect 619 738 625 739
rect 658 739 659 740
rect 663 739 664 743
rect 658 738 664 739
rect 667 743 673 744
rect 667 739 668 743
rect 672 742 673 743
rect 698 743 704 744
rect 698 742 699 743
rect 672 740 699 742
rect 672 739 673 740
rect 667 738 673 739
rect 698 739 699 740
rect 703 739 704 743
rect 698 738 704 739
rect 706 743 712 744
rect 706 739 707 743
rect 711 742 712 743
rect 715 743 721 744
rect 715 742 716 743
rect 711 740 716 742
rect 711 739 712 740
rect 706 738 712 739
rect 715 739 716 740
rect 720 739 721 743
rect 715 738 721 739
rect 754 743 760 744
rect 754 739 755 743
rect 759 742 760 743
rect 763 743 769 744
rect 763 742 764 743
rect 759 740 764 742
rect 759 739 760 740
rect 754 738 760 739
rect 763 739 764 740
rect 768 739 769 743
rect 763 738 769 739
rect 806 743 817 744
rect 806 739 807 743
rect 811 739 812 743
rect 816 739 817 743
rect 806 738 817 739
rect 850 743 856 744
rect 850 739 851 743
rect 855 742 856 743
rect 859 743 865 744
rect 859 742 860 743
rect 855 740 860 742
rect 855 739 856 740
rect 850 738 856 739
rect 859 739 860 740
rect 864 739 865 743
rect 859 738 865 739
rect 898 743 904 744
rect 898 739 899 743
rect 903 742 904 743
rect 907 743 913 744
rect 907 742 908 743
rect 903 740 908 742
rect 903 739 904 740
rect 898 738 904 739
rect 907 739 908 740
rect 912 739 913 743
rect 907 738 913 739
rect 1299 739 1305 740
rect 134 735 140 736
rect 134 731 135 735
rect 139 731 140 735
rect 134 730 140 731
rect 190 735 196 736
rect 190 731 191 735
rect 195 731 196 735
rect 190 730 196 731
rect 262 735 268 736
rect 262 731 263 735
rect 267 731 268 735
rect 262 730 268 731
rect 334 735 340 736
rect 334 731 335 735
rect 339 731 340 735
rect 334 730 340 731
rect 398 735 404 736
rect 398 731 399 735
rect 403 731 404 735
rect 398 730 404 731
rect 454 735 460 736
rect 454 731 455 735
rect 459 731 460 735
rect 454 730 460 731
rect 502 735 508 736
rect 502 731 503 735
rect 507 731 508 735
rect 502 730 508 731
rect 542 735 548 736
rect 542 731 543 735
rect 547 731 548 735
rect 542 730 548 731
rect 582 735 588 736
rect 582 731 583 735
rect 587 731 588 735
rect 582 730 588 731
rect 622 735 628 736
rect 622 731 623 735
rect 627 731 628 735
rect 622 730 628 731
rect 670 735 676 736
rect 670 731 671 735
rect 675 731 676 735
rect 670 730 676 731
rect 718 735 724 736
rect 718 731 719 735
rect 723 731 724 735
rect 718 730 724 731
rect 766 735 772 736
rect 766 731 767 735
rect 771 731 772 735
rect 766 730 772 731
rect 814 735 820 736
rect 814 731 815 735
rect 819 731 820 735
rect 814 730 820 731
rect 862 735 868 736
rect 862 731 863 735
rect 867 731 868 735
rect 862 730 868 731
rect 910 735 916 736
rect 910 731 911 735
rect 915 731 916 735
rect 1299 735 1300 739
rect 1304 738 1305 739
rect 1322 739 1328 740
rect 1322 738 1323 739
rect 1304 736 1323 738
rect 1304 735 1305 736
rect 1299 734 1305 735
rect 1322 735 1323 736
rect 1327 735 1328 739
rect 1322 734 1328 735
rect 1330 739 1336 740
rect 1330 735 1331 739
rect 1335 738 1336 739
rect 1339 739 1345 740
rect 1339 738 1340 739
rect 1335 736 1340 738
rect 1335 735 1336 736
rect 1330 734 1336 735
rect 1339 735 1340 736
rect 1344 735 1345 739
rect 1339 734 1345 735
rect 1370 739 1376 740
rect 1370 735 1371 739
rect 1375 738 1376 739
rect 1403 739 1409 740
rect 1403 738 1404 739
rect 1375 736 1404 738
rect 1375 735 1376 736
rect 1370 734 1376 735
rect 1403 735 1404 736
rect 1408 735 1409 739
rect 1403 734 1409 735
rect 1434 739 1440 740
rect 1434 735 1435 739
rect 1439 738 1440 739
rect 1483 739 1489 740
rect 1483 738 1484 739
rect 1439 736 1484 738
rect 1439 735 1440 736
rect 1434 734 1440 735
rect 1483 735 1484 736
rect 1488 735 1489 739
rect 1483 734 1489 735
rect 1514 739 1520 740
rect 1514 735 1515 739
rect 1519 738 1520 739
rect 1571 739 1577 740
rect 1571 738 1572 739
rect 1519 736 1572 738
rect 1519 735 1520 736
rect 1514 734 1520 735
rect 1571 735 1572 736
rect 1576 735 1577 739
rect 1571 734 1577 735
rect 1659 739 1665 740
rect 1659 735 1660 739
rect 1664 738 1665 739
rect 1670 739 1676 740
rect 1670 738 1671 739
rect 1664 736 1671 738
rect 1664 735 1665 736
rect 1659 734 1665 735
rect 1670 735 1671 736
rect 1675 735 1676 739
rect 1670 734 1676 735
rect 1690 739 1696 740
rect 1690 735 1691 739
rect 1695 738 1696 739
rect 1747 739 1753 740
rect 1747 738 1748 739
rect 1695 736 1748 738
rect 1695 735 1696 736
rect 1690 734 1696 735
rect 1747 735 1748 736
rect 1752 735 1753 739
rect 1747 734 1753 735
rect 1827 739 1833 740
rect 1827 735 1828 739
rect 1832 738 1833 739
rect 1838 739 1844 740
rect 1838 738 1839 739
rect 1832 736 1839 738
rect 1832 735 1833 736
rect 1827 734 1833 735
rect 1838 735 1839 736
rect 1843 735 1844 739
rect 1838 734 1844 735
rect 1858 739 1864 740
rect 1858 735 1859 739
rect 1863 738 1864 739
rect 1907 739 1913 740
rect 1907 738 1908 739
rect 1863 736 1908 738
rect 1863 735 1864 736
rect 1858 734 1864 735
rect 1907 735 1908 736
rect 1912 735 1913 739
rect 1987 739 1993 740
rect 1987 738 1988 739
rect 1936 736 1988 738
rect 1907 734 1913 735
rect 1934 735 1940 736
rect 910 730 916 731
rect 1302 731 1308 732
rect 1302 727 1303 731
rect 1307 727 1308 731
rect 1302 726 1308 727
rect 1342 731 1348 732
rect 1342 727 1343 731
rect 1347 727 1348 731
rect 1342 726 1348 727
rect 1406 731 1412 732
rect 1406 727 1407 731
rect 1411 727 1412 731
rect 1406 726 1412 727
rect 1486 731 1492 732
rect 1486 727 1487 731
rect 1491 727 1492 731
rect 1486 726 1492 727
rect 1574 731 1580 732
rect 1574 727 1575 731
rect 1579 727 1580 731
rect 1574 726 1580 727
rect 1662 731 1668 732
rect 1662 727 1663 731
rect 1667 727 1668 731
rect 1662 726 1668 727
rect 1750 731 1756 732
rect 1750 727 1751 731
rect 1755 727 1756 731
rect 1750 726 1756 727
rect 1830 731 1836 732
rect 1830 727 1831 731
rect 1835 727 1836 731
rect 1830 726 1836 727
rect 1910 731 1916 732
rect 1910 727 1911 731
rect 1915 727 1916 731
rect 1934 731 1935 735
rect 1939 731 1940 735
rect 1987 735 1988 736
rect 1992 735 1993 739
rect 1987 734 1993 735
rect 2018 739 2024 740
rect 2018 735 2019 739
rect 2023 738 2024 739
rect 2075 739 2081 740
rect 2075 738 2076 739
rect 2023 736 2076 738
rect 2023 735 2024 736
rect 2018 734 2024 735
rect 2075 735 2076 736
rect 2080 735 2081 739
rect 2075 734 2081 735
rect 2106 739 2112 740
rect 2106 735 2107 739
rect 2111 738 2112 739
rect 2171 739 2177 740
rect 2171 738 2172 739
rect 2111 736 2172 738
rect 2111 735 2112 736
rect 2106 734 2112 735
rect 2171 735 2172 736
rect 2176 735 2177 739
rect 2171 734 2177 735
rect 2202 739 2208 740
rect 2202 735 2203 739
rect 2207 738 2208 739
rect 2275 739 2281 740
rect 2275 738 2276 739
rect 2207 736 2276 738
rect 2207 735 2208 736
rect 2202 734 2208 735
rect 2275 735 2276 736
rect 2280 735 2281 739
rect 2275 734 2281 735
rect 2355 739 2361 740
rect 2355 735 2356 739
rect 2360 738 2361 739
rect 2370 739 2376 740
rect 2370 738 2371 739
rect 2360 736 2371 738
rect 2360 735 2361 736
rect 2355 734 2361 735
rect 2370 735 2371 736
rect 2375 735 2376 739
rect 2370 734 2376 735
rect 1934 730 1940 731
rect 1990 731 1996 732
rect 1910 726 1916 727
rect 1990 727 1991 731
rect 1995 727 1996 731
rect 1990 726 1996 727
rect 2078 731 2084 732
rect 2078 727 2079 731
rect 2083 727 2084 731
rect 2078 726 2084 727
rect 2174 731 2180 732
rect 2174 727 2175 731
rect 2179 727 2180 731
rect 2174 726 2180 727
rect 2278 731 2284 732
rect 2278 727 2279 731
rect 2283 727 2284 731
rect 2278 726 2284 727
rect 2358 731 2364 732
rect 2358 727 2359 731
rect 2363 727 2364 731
rect 2358 726 2364 727
rect 698 719 704 720
rect 698 715 699 719
rect 703 718 704 719
rect 703 716 910 718
rect 703 715 704 716
rect 698 714 704 715
rect 110 712 116 713
rect 110 708 111 712
rect 115 708 116 712
rect 754 711 760 712
rect 754 710 755 711
rect 743 709 755 710
rect 110 707 116 708
rect 154 707 165 708
rect 154 703 155 707
rect 159 703 160 707
rect 164 703 165 707
rect 154 702 165 703
rect 175 707 181 708
rect 175 703 176 707
rect 180 706 181 707
rect 215 707 221 708
rect 215 706 216 707
rect 180 704 216 706
rect 180 703 181 704
rect 175 702 181 703
rect 215 703 216 704
rect 220 703 221 707
rect 215 702 221 703
rect 286 707 293 708
rect 286 703 287 707
rect 292 703 293 707
rect 286 702 293 703
rect 319 707 325 708
rect 319 703 320 707
rect 324 706 325 707
rect 359 707 365 708
rect 359 706 360 707
rect 324 704 360 706
rect 324 703 325 704
rect 319 702 325 703
rect 359 703 360 704
rect 364 703 365 707
rect 359 702 365 703
rect 386 707 392 708
rect 386 703 387 707
rect 391 706 392 707
rect 423 707 429 708
rect 423 706 424 707
rect 391 704 424 706
rect 391 703 392 704
rect 386 702 392 703
rect 423 703 424 704
rect 428 703 429 707
rect 423 702 429 703
rect 442 707 448 708
rect 442 703 443 707
rect 447 706 448 707
rect 479 707 485 708
rect 479 706 480 707
rect 447 704 480 706
rect 447 703 448 704
rect 442 702 448 703
rect 479 703 480 704
rect 484 703 485 707
rect 479 702 485 703
rect 490 707 496 708
rect 490 703 491 707
rect 495 706 496 707
rect 527 707 533 708
rect 527 706 528 707
rect 495 704 528 706
rect 495 703 496 704
rect 490 702 496 703
rect 527 703 528 704
rect 532 703 533 707
rect 527 702 533 703
rect 538 707 544 708
rect 538 703 539 707
rect 543 706 544 707
rect 567 707 573 708
rect 567 706 568 707
rect 543 704 568 706
rect 543 703 544 704
rect 538 702 544 703
rect 567 703 568 704
rect 572 703 573 707
rect 567 702 573 703
rect 578 707 584 708
rect 578 703 579 707
rect 583 706 584 707
rect 607 707 613 708
rect 607 706 608 707
rect 583 704 608 706
rect 583 703 584 704
rect 578 702 584 703
rect 607 703 608 704
rect 612 703 613 707
rect 607 702 613 703
rect 618 707 624 708
rect 618 703 619 707
rect 623 706 624 707
rect 647 707 653 708
rect 647 706 648 707
rect 623 704 648 706
rect 623 703 624 704
rect 618 702 624 703
rect 647 703 648 704
rect 652 703 653 707
rect 647 702 653 703
rect 695 707 701 708
rect 695 703 696 707
rect 700 706 701 707
rect 706 707 712 708
rect 706 706 707 707
rect 700 704 707 706
rect 700 703 701 704
rect 695 702 701 703
rect 706 703 707 704
rect 711 703 712 707
rect 743 705 744 709
rect 748 708 755 709
rect 748 705 749 708
rect 754 707 755 708
rect 759 707 760 711
rect 754 706 760 707
rect 790 707 797 708
rect 743 704 749 705
rect 706 702 712 703
rect 790 703 791 707
rect 796 703 797 707
rect 790 702 797 703
rect 839 707 845 708
rect 839 703 840 707
rect 844 706 845 707
rect 850 707 856 708
rect 850 706 851 707
rect 844 704 851 706
rect 844 703 845 704
rect 839 702 845 703
rect 850 703 851 704
rect 855 703 856 707
rect 850 702 856 703
rect 887 707 893 708
rect 887 703 888 707
rect 892 706 893 707
rect 898 707 904 708
rect 898 706 899 707
rect 892 704 899 706
rect 892 703 893 704
rect 887 702 893 703
rect 898 703 899 704
rect 903 703 904 707
rect 908 706 910 716
rect 1238 712 1244 713
rect 1238 708 1239 712
rect 1243 708 1244 712
rect 1390 711 1396 712
rect 935 707 941 708
rect 1238 707 1244 708
rect 1278 708 1284 709
rect 935 706 936 707
rect 908 704 936 706
rect 898 702 904 703
rect 935 703 936 704
rect 940 703 941 707
rect 1278 704 1279 708
rect 1283 704 1284 708
rect 1390 707 1391 711
rect 1395 710 1396 711
rect 1395 708 1526 710
rect 1395 707 1396 708
rect 1390 706 1396 707
rect 1278 703 1284 704
rect 1327 703 1336 704
rect 935 702 941 703
rect 1327 699 1328 703
rect 1335 699 1336 703
rect 1327 698 1336 699
rect 1367 703 1376 704
rect 1367 699 1368 703
rect 1375 699 1376 703
rect 1367 698 1376 699
rect 1431 703 1440 704
rect 1431 699 1432 703
rect 1439 699 1440 703
rect 1431 698 1440 699
rect 1511 703 1520 704
rect 1511 699 1512 703
rect 1519 699 1520 703
rect 1524 702 1526 708
rect 2406 708 2412 709
rect 2406 704 2407 708
rect 2411 704 2412 708
rect 1599 703 1605 704
rect 1599 702 1600 703
rect 1524 700 1600 702
rect 1511 698 1520 699
rect 1599 699 1600 700
rect 1604 699 1605 703
rect 1599 698 1605 699
rect 1687 703 1696 704
rect 1687 699 1688 703
rect 1695 699 1696 703
rect 1687 698 1696 699
rect 1734 703 1740 704
rect 1734 699 1735 703
rect 1739 702 1740 703
rect 1775 703 1781 704
rect 1775 702 1776 703
rect 1739 700 1776 702
rect 1739 699 1740 700
rect 1734 698 1740 699
rect 1775 699 1776 700
rect 1780 699 1781 703
rect 1775 698 1781 699
rect 1855 703 1864 704
rect 1855 699 1856 703
rect 1863 699 1864 703
rect 1855 698 1864 699
rect 1934 703 1941 704
rect 1934 699 1935 703
rect 1940 699 1941 703
rect 1934 698 1941 699
rect 2015 703 2024 704
rect 2015 699 2016 703
rect 2023 699 2024 703
rect 2015 698 2024 699
rect 2103 703 2112 704
rect 2103 699 2104 703
rect 2111 699 2112 703
rect 2103 698 2112 699
rect 2199 703 2208 704
rect 2199 699 2200 703
rect 2207 699 2208 703
rect 2199 698 2208 699
rect 2246 703 2252 704
rect 2246 699 2247 703
rect 2251 702 2252 703
rect 2303 703 2309 704
rect 2303 702 2304 703
rect 2251 700 2304 702
rect 2251 699 2252 700
rect 2246 698 2252 699
rect 2303 699 2304 700
rect 2308 699 2309 703
rect 2303 698 2309 699
rect 2378 703 2389 704
rect 2406 703 2412 704
rect 2378 699 2379 703
rect 2383 699 2384 703
rect 2388 699 2389 703
rect 2378 698 2389 699
rect 110 695 116 696
rect 110 691 111 695
rect 115 691 116 695
rect 110 690 116 691
rect 1238 695 1244 696
rect 1238 691 1239 695
rect 1243 691 1244 695
rect 1238 690 1244 691
rect 1278 691 1284 692
rect 134 688 140 689
rect 134 684 135 688
rect 139 684 140 688
rect 134 683 140 684
rect 190 688 196 689
rect 190 684 191 688
rect 195 684 196 688
rect 190 683 196 684
rect 262 688 268 689
rect 262 684 263 688
rect 267 684 268 688
rect 262 683 268 684
rect 334 688 340 689
rect 334 684 335 688
rect 339 684 340 688
rect 334 683 340 684
rect 398 688 404 689
rect 398 684 399 688
rect 403 684 404 688
rect 398 683 404 684
rect 454 688 460 689
rect 454 684 455 688
rect 459 684 460 688
rect 454 683 460 684
rect 502 688 508 689
rect 502 684 503 688
rect 507 684 508 688
rect 502 683 508 684
rect 542 688 548 689
rect 542 684 543 688
rect 547 684 548 688
rect 542 683 548 684
rect 582 688 588 689
rect 582 684 583 688
rect 587 684 588 688
rect 582 683 588 684
rect 622 688 628 689
rect 622 684 623 688
rect 627 684 628 688
rect 622 683 628 684
rect 670 688 676 689
rect 670 684 671 688
rect 675 684 676 688
rect 670 683 676 684
rect 718 688 724 689
rect 718 684 719 688
rect 723 684 724 688
rect 718 683 724 684
rect 766 688 772 689
rect 766 684 767 688
rect 771 684 772 688
rect 766 683 772 684
rect 814 688 820 689
rect 814 684 815 688
rect 819 684 820 688
rect 814 683 820 684
rect 862 688 868 689
rect 862 684 863 688
rect 867 684 868 688
rect 862 683 868 684
rect 910 688 916 689
rect 910 684 911 688
rect 915 684 916 688
rect 1278 687 1279 691
rect 1283 687 1284 691
rect 1278 686 1284 687
rect 2406 691 2412 692
rect 2406 687 2407 691
rect 2411 687 2412 691
rect 2406 686 2412 687
rect 910 683 916 684
rect 1302 684 1308 685
rect 1302 680 1303 684
rect 1307 680 1308 684
rect 1302 679 1308 680
rect 1342 684 1348 685
rect 1342 680 1343 684
rect 1347 680 1348 684
rect 1342 679 1348 680
rect 1406 684 1412 685
rect 1406 680 1407 684
rect 1411 680 1412 684
rect 1406 679 1412 680
rect 1486 684 1492 685
rect 1486 680 1487 684
rect 1491 680 1492 684
rect 1486 679 1492 680
rect 1574 684 1580 685
rect 1574 680 1575 684
rect 1579 680 1580 684
rect 1574 679 1580 680
rect 1662 684 1668 685
rect 1662 680 1663 684
rect 1667 680 1668 684
rect 1662 679 1668 680
rect 1750 684 1756 685
rect 1750 680 1751 684
rect 1755 680 1756 684
rect 1750 679 1756 680
rect 1830 684 1836 685
rect 1830 680 1831 684
rect 1835 680 1836 684
rect 1830 679 1836 680
rect 1910 684 1916 685
rect 1910 680 1911 684
rect 1915 680 1916 684
rect 1910 679 1916 680
rect 1990 684 1996 685
rect 1990 680 1991 684
rect 1995 680 1996 684
rect 1990 679 1996 680
rect 2078 684 2084 685
rect 2078 680 2079 684
rect 2083 680 2084 684
rect 2078 679 2084 680
rect 2174 684 2180 685
rect 2174 680 2175 684
rect 2179 680 2180 684
rect 2174 679 2180 680
rect 2278 684 2284 685
rect 2278 680 2279 684
rect 2283 680 2284 684
rect 2278 679 2284 680
rect 2358 684 2364 685
rect 2358 680 2359 684
rect 2363 680 2364 684
rect 2358 679 2364 680
rect 134 672 140 673
rect 134 668 135 672
rect 139 668 140 672
rect 134 667 140 668
rect 198 672 204 673
rect 198 668 199 672
rect 203 668 204 672
rect 198 667 204 668
rect 278 672 284 673
rect 278 668 279 672
rect 283 668 284 672
rect 278 667 284 668
rect 350 672 356 673
rect 350 668 351 672
rect 355 668 356 672
rect 350 667 356 668
rect 414 672 420 673
rect 414 668 415 672
rect 419 668 420 672
rect 414 667 420 668
rect 486 672 492 673
rect 486 668 487 672
rect 491 668 492 672
rect 486 667 492 668
rect 558 672 564 673
rect 558 668 559 672
rect 563 668 564 672
rect 558 667 564 668
rect 638 672 644 673
rect 638 668 639 672
rect 643 668 644 672
rect 638 667 644 668
rect 710 672 716 673
rect 710 668 711 672
rect 715 668 716 672
rect 710 667 716 668
rect 782 672 788 673
rect 782 668 783 672
rect 787 668 788 672
rect 782 667 788 668
rect 854 672 860 673
rect 854 668 855 672
rect 859 668 860 672
rect 854 667 860 668
rect 918 672 924 673
rect 918 668 919 672
rect 923 668 924 672
rect 918 667 924 668
rect 982 672 988 673
rect 982 668 983 672
rect 987 668 988 672
rect 982 667 988 668
rect 1038 672 1044 673
rect 1038 668 1039 672
rect 1043 668 1044 672
rect 1038 667 1044 668
rect 1094 672 1100 673
rect 1094 668 1095 672
rect 1099 668 1100 672
rect 1094 667 1100 668
rect 1150 672 1156 673
rect 1150 668 1151 672
rect 1155 668 1156 672
rect 1150 667 1156 668
rect 1190 672 1196 673
rect 1190 668 1191 672
rect 1195 668 1196 672
rect 1190 667 1196 668
rect 1302 668 1308 669
rect 110 665 116 666
rect 110 661 111 665
rect 115 661 116 665
rect 110 660 116 661
rect 1238 665 1244 666
rect 1238 661 1239 665
rect 1243 661 1244 665
rect 1302 664 1303 668
rect 1307 664 1308 668
rect 1302 663 1308 664
rect 1398 668 1404 669
rect 1398 664 1399 668
rect 1403 664 1404 668
rect 1398 663 1404 664
rect 1510 668 1516 669
rect 1510 664 1511 668
rect 1515 664 1516 668
rect 1510 663 1516 664
rect 1622 668 1628 669
rect 1622 664 1623 668
rect 1627 664 1628 668
rect 1622 663 1628 664
rect 1726 668 1732 669
rect 1726 664 1727 668
rect 1731 664 1732 668
rect 1726 663 1732 664
rect 1814 668 1820 669
rect 1814 664 1815 668
rect 1819 664 1820 668
rect 1814 663 1820 664
rect 1894 668 1900 669
rect 1894 664 1895 668
rect 1899 664 1900 668
rect 1894 663 1900 664
rect 1974 668 1980 669
rect 1974 664 1975 668
rect 1979 664 1980 668
rect 1974 663 1980 664
rect 2046 668 2052 669
rect 2046 664 2047 668
rect 2051 664 2052 668
rect 2046 663 2052 664
rect 2110 668 2116 669
rect 2110 664 2111 668
rect 2115 664 2116 668
rect 2110 663 2116 664
rect 2174 668 2180 669
rect 2174 664 2175 668
rect 2179 664 2180 668
rect 2174 663 2180 664
rect 2238 668 2244 669
rect 2238 664 2239 668
rect 2243 664 2244 668
rect 2238 663 2244 664
rect 2310 668 2316 669
rect 2310 664 2311 668
rect 2315 664 2316 668
rect 2310 663 2316 664
rect 2358 668 2364 669
rect 2358 664 2359 668
rect 2363 664 2364 668
rect 2358 663 2364 664
rect 1238 660 1244 661
rect 1278 661 1284 662
rect 1278 657 1279 661
rect 1283 657 1284 661
rect 1278 656 1284 657
rect 2406 661 2412 662
rect 2406 657 2407 661
rect 2411 657 2412 661
rect 2406 656 2412 657
rect 159 651 165 652
rect 110 648 116 649
rect 110 644 111 648
rect 115 644 116 648
rect 159 647 160 651
rect 164 650 165 651
rect 190 651 196 652
rect 190 650 191 651
rect 164 648 191 650
rect 164 647 165 648
rect 159 646 165 647
rect 190 647 191 648
rect 195 647 196 651
rect 190 646 196 647
rect 222 651 229 652
rect 222 647 223 651
rect 228 647 229 651
rect 222 646 229 647
rect 303 651 309 652
rect 303 647 304 651
rect 308 650 309 651
rect 342 651 348 652
rect 342 650 343 651
rect 308 648 343 650
rect 308 647 309 648
rect 303 646 309 647
rect 342 647 343 648
rect 347 647 348 651
rect 342 646 348 647
rect 375 651 381 652
rect 375 647 376 651
rect 380 650 381 651
rect 406 651 412 652
rect 406 650 407 651
rect 380 648 407 650
rect 380 647 381 648
rect 375 646 381 647
rect 406 647 407 648
rect 411 647 412 651
rect 406 646 412 647
rect 439 651 445 652
rect 439 647 440 651
rect 444 650 445 651
rect 478 651 484 652
rect 478 650 479 651
rect 444 648 479 650
rect 444 647 445 648
rect 439 646 445 647
rect 478 647 479 648
rect 483 647 484 651
rect 478 646 484 647
rect 511 651 517 652
rect 511 647 512 651
rect 516 650 517 651
rect 550 651 556 652
rect 550 650 551 651
rect 516 648 551 650
rect 516 647 517 648
rect 511 646 517 647
rect 550 647 551 648
rect 555 647 556 651
rect 550 646 556 647
rect 583 651 589 652
rect 583 647 584 651
rect 588 650 589 651
rect 614 651 620 652
rect 614 650 615 651
rect 588 648 615 650
rect 588 647 589 648
rect 583 646 589 647
rect 614 647 615 648
rect 619 647 620 651
rect 614 646 620 647
rect 658 651 669 652
rect 658 647 659 651
rect 663 647 664 651
rect 668 647 669 651
rect 658 646 669 647
rect 671 651 677 652
rect 671 647 672 651
rect 676 650 677 651
rect 735 651 741 652
rect 735 650 736 651
rect 676 648 736 650
rect 676 647 677 648
rect 671 646 677 647
rect 735 647 736 648
rect 740 647 741 651
rect 735 646 741 647
rect 743 651 749 652
rect 743 647 744 651
rect 748 650 749 651
rect 807 651 813 652
rect 807 650 808 651
rect 748 648 808 650
rect 748 647 749 648
rect 743 646 749 647
rect 807 647 808 648
rect 812 647 813 651
rect 807 646 813 647
rect 879 651 885 652
rect 879 647 880 651
rect 884 650 885 651
rect 910 651 916 652
rect 910 650 911 651
rect 884 648 911 650
rect 884 647 885 648
rect 879 646 885 647
rect 910 647 911 648
rect 915 647 916 651
rect 910 646 916 647
rect 943 651 949 652
rect 943 647 944 651
rect 948 650 949 651
rect 974 651 980 652
rect 974 650 975 651
rect 948 648 975 650
rect 948 647 949 648
rect 943 646 949 647
rect 974 647 975 648
rect 979 647 980 651
rect 974 646 980 647
rect 1007 651 1013 652
rect 1007 647 1008 651
rect 1012 650 1013 651
rect 1022 651 1028 652
rect 1022 650 1023 651
rect 1012 648 1023 650
rect 1012 647 1013 648
rect 1007 646 1013 647
rect 1022 647 1023 648
rect 1027 647 1028 651
rect 1022 646 1028 647
rect 1063 651 1069 652
rect 1063 647 1064 651
rect 1068 650 1069 651
rect 1086 651 1092 652
rect 1086 650 1087 651
rect 1068 648 1087 650
rect 1068 647 1069 648
rect 1063 646 1069 647
rect 1086 647 1087 648
rect 1091 647 1092 651
rect 1086 646 1092 647
rect 1119 651 1125 652
rect 1119 647 1120 651
rect 1124 650 1125 651
rect 1142 651 1148 652
rect 1142 650 1143 651
rect 1124 648 1143 650
rect 1124 647 1125 648
rect 1119 646 1125 647
rect 1142 647 1143 648
rect 1147 647 1148 651
rect 1142 646 1148 647
rect 1175 651 1184 652
rect 1175 647 1176 651
rect 1183 647 1184 651
rect 1175 646 1184 647
rect 1215 651 1221 652
rect 1215 647 1216 651
rect 1220 650 1221 651
rect 1230 651 1236 652
rect 1230 650 1231 651
rect 1220 648 1231 650
rect 1220 647 1221 648
rect 1215 646 1221 647
rect 1230 647 1231 648
rect 1235 647 1236 651
rect 1230 646 1236 647
rect 1238 648 1244 649
rect 110 643 116 644
rect 1238 644 1239 648
rect 1243 644 1244 648
rect 1322 647 1333 648
rect 1238 643 1244 644
rect 1278 644 1284 645
rect 1278 640 1279 644
rect 1283 640 1284 644
rect 1322 643 1323 647
rect 1327 643 1328 647
rect 1332 643 1333 647
rect 1322 642 1333 643
rect 1423 647 1429 648
rect 1423 643 1424 647
rect 1428 646 1429 647
rect 1502 647 1508 648
rect 1502 646 1503 647
rect 1428 644 1503 646
rect 1428 643 1429 644
rect 1423 642 1429 643
rect 1502 643 1503 644
rect 1507 643 1508 647
rect 1502 642 1508 643
rect 1535 647 1541 648
rect 1535 643 1536 647
rect 1540 646 1541 647
rect 1590 647 1596 648
rect 1590 646 1591 647
rect 1540 644 1591 646
rect 1540 643 1541 644
rect 1535 642 1541 643
rect 1590 643 1591 644
rect 1595 643 1596 647
rect 1647 647 1653 648
rect 1647 646 1648 647
rect 1590 642 1596 643
rect 1600 644 1648 646
rect 1278 639 1284 640
rect 1406 639 1412 640
rect 1406 635 1407 639
rect 1411 638 1412 639
rect 1600 638 1602 644
rect 1647 643 1648 644
rect 1652 643 1653 647
rect 1647 642 1653 643
rect 1655 647 1661 648
rect 1655 643 1656 647
rect 1660 646 1661 647
rect 1751 647 1757 648
rect 1751 646 1752 647
rect 1660 644 1752 646
rect 1660 643 1661 644
rect 1655 642 1661 643
rect 1751 643 1752 644
rect 1756 643 1757 647
rect 1751 642 1757 643
rect 1839 647 1845 648
rect 1839 643 1840 647
rect 1844 646 1845 647
rect 1886 647 1892 648
rect 1886 646 1887 647
rect 1844 644 1887 646
rect 1844 643 1845 644
rect 1839 642 1845 643
rect 1886 643 1887 644
rect 1891 643 1892 647
rect 1886 642 1892 643
rect 1919 647 1925 648
rect 1919 643 1920 647
rect 1924 646 1925 647
rect 1966 647 1972 648
rect 1966 646 1967 647
rect 1924 644 1967 646
rect 1924 643 1925 644
rect 1919 642 1925 643
rect 1966 643 1967 644
rect 1971 643 1972 647
rect 1966 642 1972 643
rect 1999 647 2005 648
rect 1999 643 2000 647
rect 2004 646 2005 647
rect 2022 647 2028 648
rect 2022 646 2023 647
rect 2004 644 2023 646
rect 2004 643 2005 644
rect 1999 642 2005 643
rect 2022 643 2023 644
rect 2027 643 2028 647
rect 2071 647 2077 648
rect 2071 646 2072 647
rect 2022 642 2028 643
rect 2036 644 2072 646
rect 1411 636 1602 638
rect 1822 639 1828 640
rect 1411 635 1412 636
rect 1406 634 1412 635
rect 1822 635 1823 639
rect 1827 638 1828 639
rect 2036 638 2038 644
rect 2071 643 2072 644
rect 2076 643 2077 647
rect 2071 642 2077 643
rect 2079 647 2085 648
rect 2079 643 2080 647
rect 2084 646 2085 647
rect 2135 647 2141 648
rect 2135 646 2136 647
rect 2084 644 2136 646
rect 2084 643 2085 644
rect 2079 642 2085 643
rect 2135 643 2136 644
rect 2140 643 2141 647
rect 2135 642 2141 643
rect 2143 647 2149 648
rect 2143 643 2144 647
rect 2148 646 2149 647
rect 2199 647 2205 648
rect 2199 646 2200 647
rect 2148 644 2200 646
rect 2148 643 2149 644
rect 2143 642 2149 643
rect 2199 643 2200 644
rect 2204 643 2205 647
rect 2199 642 2205 643
rect 2207 647 2213 648
rect 2207 643 2208 647
rect 2212 646 2213 647
rect 2263 647 2269 648
rect 2263 646 2264 647
rect 2212 644 2264 646
rect 2212 643 2213 644
rect 2207 642 2213 643
rect 2263 643 2264 644
rect 2268 643 2269 647
rect 2263 642 2269 643
rect 2286 647 2292 648
rect 2286 643 2287 647
rect 2291 646 2292 647
rect 2335 647 2341 648
rect 2335 646 2336 647
rect 2291 644 2336 646
rect 2291 643 2292 644
rect 2286 642 2292 643
rect 2335 643 2336 644
rect 2340 643 2341 647
rect 2335 642 2341 643
rect 2370 647 2376 648
rect 2370 643 2371 647
rect 2375 646 2376 647
rect 2383 647 2389 648
rect 2383 646 2384 647
rect 2375 644 2384 646
rect 2375 643 2376 644
rect 2370 642 2376 643
rect 2383 643 2384 644
rect 2388 643 2389 647
rect 2383 642 2389 643
rect 2406 644 2412 645
rect 2406 640 2407 644
rect 2411 640 2412 644
rect 2406 639 2412 640
rect 1827 636 2038 638
rect 1827 635 1828 636
rect 1822 634 1828 635
rect 134 625 140 626
rect 134 621 135 625
rect 139 621 140 625
rect 134 620 140 621
rect 198 625 204 626
rect 198 621 199 625
rect 203 621 204 625
rect 198 620 204 621
rect 278 625 284 626
rect 278 621 279 625
rect 283 621 284 625
rect 278 620 284 621
rect 350 625 356 626
rect 350 621 351 625
rect 355 621 356 625
rect 350 620 356 621
rect 414 625 420 626
rect 414 621 415 625
rect 419 621 420 625
rect 414 620 420 621
rect 486 625 492 626
rect 486 621 487 625
rect 491 621 492 625
rect 486 620 492 621
rect 558 625 564 626
rect 558 621 559 625
rect 563 621 564 625
rect 558 620 564 621
rect 638 625 644 626
rect 638 621 639 625
rect 643 621 644 625
rect 638 620 644 621
rect 710 625 716 626
rect 710 621 711 625
rect 715 621 716 625
rect 710 620 716 621
rect 782 625 788 626
rect 782 621 783 625
rect 787 621 788 625
rect 782 620 788 621
rect 854 625 860 626
rect 854 621 855 625
rect 859 621 860 625
rect 854 620 860 621
rect 918 625 924 626
rect 918 621 919 625
rect 923 621 924 625
rect 918 620 924 621
rect 982 625 988 626
rect 982 621 983 625
rect 987 621 988 625
rect 982 620 988 621
rect 1038 625 1044 626
rect 1038 621 1039 625
rect 1043 621 1044 625
rect 1038 620 1044 621
rect 1094 625 1100 626
rect 1094 621 1095 625
rect 1099 621 1100 625
rect 1094 620 1100 621
rect 1150 625 1156 626
rect 1150 621 1151 625
rect 1155 621 1156 625
rect 1150 620 1156 621
rect 1190 625 1196 626
rect 1190 621 1191 625
rect 1195 621 1196 625
rect 1190 620 1196 621
rect 1302 621 1308 622
rect 1302 617 1303 621
rect 1307 617 1308 621
rect 1302 616 1308 617
rect 1398 621 1404 622
rect 1398 617 1399 621
rect 1403 617 1404 621
rect 1398 616 1404 617
rect 1510 621 1516 622
rect 1510 617 1511 621
rect 1515 617 1516 621
rect 1510 616 1516 617
rect 1622 621 1628 622
rect 1622 617 1623 621
rect 1627 617 1628 621
rect 1622 616 1628 617
rect 1726 621 1732 622
rect 1726 617 1727 621
rect 1731 617 1732 621
rect 1726 616 1732 617
rect 1814 621 1820 622
rect 1814 617 1815 621
rect 1819 617 1820 621
rect 1814 616 1820 617
rect 1894 621 1900 622
rect 1894 617 1895 621
rect 1899 617 1900 621
rect 1894 616 1900 617
rect 1974 621 1980 622
rect 1974 617 1975 621
rect 1979 617 1980 621
rect 1974 616 1980 617
rect 2046 621 2052 622
rect 2046 617 2047 621
rect 2051 617 2052 621
rect 2046 616 2052 617
rect 2110 621 2116 622
rect 2110 617 2111 621
rect 2115 617 2116 621
rect 2110 616 2116 617
rect 2174 621 2180 622
rect 2174 617 2175 621
rect 2179 617 2180 621
rect 2174 616 2180 617
rect 2238 621 2244 622
rect 2238 617 2239 621
rect 2243 617 2244 621
rect 2238 616 2244 617
rect 2310 621 2316 622
rect 2310 617 2311 621
rect 2315 617 2316 621
rect 2310 616 2316 617
rect 2358 621 2364 622
rect 2358 617 2359 621
rect 2363 617 2364 621
rect 2358 616 2364 617
rect 131 615 137 616
rect 131 611 132 615
rect 136 614 137 615
rect 158 615 164 616
rect 158 614 159 615
rect 136 612 159 614
rect 136 611 137 612
rect 131 610 137 611
rect 158 611 159 612
rect 163 611 164 615
rect 158 610 164 611
rect 190 615 201 616
rect 190 611 191 615
rect 195 611 196 615
rect 200 611 201 615
rect 190 610 201 611
rect 275 615 281 616
rect 275 611 276 615
rect 280 614 281 615
rect 286 615 292 616
rect 286 614 287 615
rect 280 612 287 614
rect 280 611 281 612
rect 275 610 281 611
rect 286 611 287 612
rect 291 611 292 615
rect 286 610 292 611
rect 342 615 353 616
rect 342 611 343 615
rect 347 611 348 615
rect 352 611 353 615
rect 342 610 353 611
rect 406 615 417 616
rect 406 611 407 615
rect 411 611 412 615
rect 416 611 417 615
rect 406 610 417 611
rect 478 615 489 616
rect 478 611 479 615
rect 483 611 484 615
rect 488 611 489 615
rect 478 610 489 611
rect 550 615 561 616
rect 550 611 551 615
rect 555 611 556 615
rect 560 611 561 615
rect 550 610 561 611
rect 635 615 641 616
rect 635 611 636 615
rect 640 614 641 615
rect 671 615 677 616
rect 671 614 672 615
rect 640 612 672 614
rect 640 611 641 612
rect 635 610 641 611
rect 671 611 672 612
rect 676 611 677 615
rect 671 610 677 611
rect 707 615 713 616
rect 707 611 708 615
rect 712 614 713 615
rect 743 615 749 616
rect 743 614 744 615
rect 712 612 744 614
rect 712 611 713 612
rect 707 610 713 611
rect 743 611 744 612
rect 748 611 749 615
rect 743 610 749 611
rect 779 615 785 616
rect 779 611 780 615
rect 784 614 785 615
rect 790 615 796 616
rect 790 614 791 615
rect 784 612 791 614
rect 784 611 785 612
rect 779 610 785 611
rect 790 611 791 612
rect 795 611 796 615
rect 790 610 796 611
rect 851 615 857 616
rect 851 611 852 615
rect 856 614 857 615
rect 902 615 908 616
rect 902 614 903 615
rect 856 612 903 614
rect 856 611 857 612
rect 851 610 857 611
rect 902 611 903 612
rect 907 611 908 615
rect 902 610 908 611
rect 910 615 921 616
rect 910 611 911 615
rect 915 611 916 615
rect 920 611 921 615
rect 910 610 921 611
rect 974 615 985 616
rect 974 611 975 615
rect 979 611 980 615
rect 984 611 985 615
rect 974 610 985 611
rect 1022 615 1028 616
rect 1022 611 1023 615
rect 1027 614 1028 615
rect 1035 615 1041 616
rect 1035 614 1036 615
rect 1027 612 1036 614
rect 1027 611 1028 612
rect 1022 610 1028 611
rect 1035 611 1036 612
rect 1040 611 1041 615
rect 1035 610 1041 611
rect 1086 615 1097 616
rect 1086 611 1087 615
rect 1091 611 1092 615
rect 1096 611 1097 615
rect 1086 610 1097 611
rect 1142 615 1153 616
rect 1142 611 1143 615
rect 1147 611 1148 615
rect 1152 611 1153 615
rect 1142 610 1153 611
rect 1178 615 1184 616
rect 1178 611 1179 615
rect 1183 614 1184 615
rect 1187 615 1193 616
rect 1187 614 1188 615
rect 1183 612 1188 614
rect 1183 611 1184 612
rect 1178 610 1184 611
rect 1187 611 1188 612
rect 1192 611 1193 615
rect 1187 610 1193 611
rect 1230 611 1236 612
rect 1230 607 1231 611
rect 1235 610 1236 611
rect 1299 611 1305 612
rect 1299 610 1300 611
rect 1235 608 1300 610
rect 1235 607 1236 608
rect 1230 606 1236 607
rect 1299 607 1300 608
rect 1304 607 1305 611
rect 1299 606 1305 607
rect 1395 611 1401 612
rect 1395 607 1396 611
rect 1400 610 1401 611
rect 1406 611 1412 612
rect 1406 610 1407 611
rect 1400 608 1407 610
rect 1400 607 1401 608
rect 1395 606 1401 607
rect 1406 607 1407 608
rect 1411 607 1412 611
rect 1406 606 1412 607
rect 1502 611 1513 612
rect 1502 607 1503 611
rect 1507 607 1508 611
rect 1512 607 1513 611
rect 1502 606 1513 607
rect 1619 611 1625 612
rect 1619 607 1620 611
rect 1624 610 1625 611
rect 1655 611 1661 612
rect 1655 610 1656 611
rect 1624 608 1656 610
rect 1624 607 1625 608
rect 1619 606 1625 607
rect 1655 607 1656 608
rect 1660 607 1661 611
rect 1655 606 1661 607
rect 1723 611 1729 612
rect 1723 607 1724 611
rect 1728 610 1729 611
rect 1734 611 1740 612
rect 1734 610 1735 611
rect 1728 608 1735 610
rect 1728 607 1729 608
rect 1723 606 1729 607
rect 1734 607 1735 608
rect 1739 607 1740 611
rect 1734 606 1740 607
rect 1811 611 1817 612
rect 1811 607 1812 611
rect 1816 610 1817 611
rect 1822 611 1828 612
rect 1822 610 1823 611
rect 1816 608 1823 610
rect 1816 607 1817 608
rect 1811 606 1817 607
rect 1822 607 1823 608
rect 1827 607 1828 611
rect 1822 606 1828 607
rect 1886 611 1897 612
rect 1886 607 1887 611
rect 1891 607 1892 611
rect 1896 607 1897 611
rect 1886 606 1897 607
rect 1966 611 1977 612
rect 1966 607 1967 611
rect 1971 607 1972 611
rect 1976 607 1977 611
rect 1966 606 1977 607
rect 2043 611 2049 612
rect 2043 607 2044 611
rect 2048 610 2049 611
rect 2079 611 2085 612
rect 2079 610 2080 611
rect 2048 608 2080 610
rect 2048 607 2049 608
rect 2043 606 2049 607
rect 2079 607 2080 608
rect 2084 607 2085 611
rect 2079 606 2085 607
rect 2107 611 2113 612
rect 2107 607 2108 611
rect 2112 610 2113 611
rect 2143 611 2149 612
rect 2143 610 2144 611
rect 2112 608 2144 610
rect 2112 607 2113 608
rect 2107 606 2113 607
rect 2143 607 2144 608
rect 2148 607 2149 611
rect 2143 606 2149 607
rect 2171 611 2177 612
rect 2171 607 2172 611
rect 2176 610 2177 611
rect 2207 611 2213 612
rect 2207 610 2208 611
rect 2176 608 2208 610
rect 2176 607 2177 608
rect 2171 606 2177 607
rect 2207 607 2208 608
rect 2212 607 2213 611
rect 2207 606 2213 607
rect 2235 611 2241 612
rect 2235 607 2236 611
rect 2240 610 2241 611
rect 2246 611 2252 612
rect 2246 610 2247 611
rect 2240 608 2247 610
rect 2240 607 2241 608
rect 2235 606 2241 607
rect 2246 607 2247 608
rect 2251 607 2252 611
rect 2246 606 2252 607
rect 2302 611 2313 612
rect 2302 607 2303 611
rect 2307 607 2308 611
rect 2312 607 2313 611
rect 2302 606 2313 607
rect 2355 611 2361 612
rect 2355 607 2356 611
rect 2360 610 2361 611
rect 2378 611 2384 612
rect 2378 610 2379 611
rect 2360 608 2379 610
rect 2360 607 2361 608
rect 2355 606 2361 607
rect 2378 607 2379 608
rect 2383 607 2384 611
rect 2378 606 2384 607
rect 131 595 137 596
rect 131 591 132 595
rect 136 594 137 595
rect 178 595 184 596
rect 178 594 179 595
rect 136 592 179 594
rect 136 591 137 592
rect 131 590 137 591
rect 178 591 179 592
rect 183 591 184 595
rect 178 590 184 591
rect 187 595 193 596
rect 187 591 188 595
rect 192 594 193 595
rect 258 595 264 596
rect 258 594 259 595
rect 192 592 259 594
rect 192 591 193 592
rect 187 590 193 591
rect 258 591 259 592
rect 263 591 264 595
rect 258 590 264 591
rect 267 595 273 596
rect 267 591 268 595
rect 272 594 273 595
rect 286 595 292 596
rect 286 594 287 595
rect 272 592 287 594
rect 272 591 273 592
rect 267 590 273 591
rect 286 591 287 592
rect 291 591 292 595
rect 286 590 292 591
rect 355 595 361 596
rect 355 591 356 595
rect 360 594 361 595
rect 378 595 384 596
rect 378 594 379 595
rect 360 592 379 594
rect 360 591 361 592
rect 355 590 361 591
rect 378 591 379 592
rect 383 591 384 595
rect 378 590 384 591
rect 386 595 392 596
rect 386 591 387 595
rect 391 594 392 595
rect 443 595 449 596
rect 443 594 444 595
rect 391 592 444 594
rect 391 591 392 592
rect 386 590 392 591
rect 443 591 444 592
rect 448 591 449 595
rect 443 590 449 591
rect 474 595 480 596
rect 474 591 475 595
rect 479 594 480 595
rect 531 595 537 596
rect 531 594 532 595
rect 479 592 532 594
rect 479 591 480 592
rect 474 590 480 591
rect 531 591 532 592
rect 536 591 537 595
rect 531 590 537 591
rect 614 595 625 596
rect 614 591 615 595
rect 619 591 620 595
rect 624 591 625 595
rect 614 590 625 591
rect 650 595 656 596
rect 650 591 651 595
rect 655 594 656 595
rect 699 595 705 596
rect 699 594 700 595
rect 655 592 700 594
rect 655 591 656 592
rect 650 590 656 591
rect 699 591 700 592
rect 704 591 705 595
rect 699 590 705 591
rect 779 595 785 596
rect 779 591 780 595
rect 784 594 785 595
rect 802 595 808 596
rect 802 594 803 595
rect 784 592 803 594
rect 784 591 785 592
rect 779 590 785 591
rect 802 591 803 592
rect 807 591 808 595
rect 802 590 808 591
rect 810 595 816 596
rect 810 591 811 595
rect 815 594 816 595
rect 851 595 857 596
rect 851 594 852 595
rect 815 592 852 594
rect 815 591 816 592
rect 810 590 816 591
rect 851 591 852 592
rect 856 591 857 595
rect 851 590 857 591
rect 882 595 888 596
rect 882 591 883 595
rect 887 594 888 595
rect 915 595 921 596
rect 915 594 916 595
rect 887 592 916 594
rect 887 591 888 592
rect 882 590 888 591
rect 915 591 916 592
rect 920 591 921 595
rect 915 590 921 591
rect 946 595 952 596
rect 946 591 947 595
rect 951 594 952 595
rect 971 595 977 596
rect 971 594 972 595
rect 951 592 972 594
rect 951 591 952 592
rect 946 590 952 591
rect 971 591 972 592
rect 976 591 977 595
rect 971 590 977 591
rect 1002 595 1008 596
rect 1002 591 1003 595
rect 1007 594 1008 595
rect 1019 595 1025 596
rect 1019 594 1020 595
rect 1007 592 1020 594
rect 1007 591 1008 592
rect 1002 590 1008 591
rect 1019 591 1020 592
rect 1024 591 1025 595
rect 1019 590 1025 591
rect 1050 595 1056 596
rect 1050 591 1051 595
rect 1055 594 1056 595
rect 1075 595 1081 596
rect 1075 594 1076 595
rect 1055 592 1076 594
rect 1055 591 1056 592
rect 1050 590 1056 591
rect 1075 591 1076 592
rect 1080 591 1081 595
rect 1075 590 1081 591
rect 1106 595 1112 596
rect 1106 591 1107 595
rect 1111 594 1112 595
rect 1131 595 1137 596
rect 1131 594 1132 595
rect 1111 592 1132 594
rect 1111 591 1112 592
rect 1106 590 1112 591
rect 1131 591 1132 592
rect 1136 591 1137 595
rect 1131 590 1137 591
rect 1162 595 1168 596
rect 1162 591 1163 595
rect 1167 594 1168 595
rect 1187 595 1193 596
rect 1187 594 1188 595
rect 1167 592 1188 594
rect 1167 591 1168 592
rect 1162 590 1168 591
rect 1187 591 1188 592
rect 1192 591 1193 595
rect 1187 590 1193 591
rect 1411 595 1417 596
rect 1411 591 1412 595
rect 1416 594 1417 595
rect 1434 595 1440 596
rect 1434 594 1435 595
rect 1416 592 1435 594
rect 1416 591 1417 592
rect 1411 590 1417 591
rect 1434 591 1435 592
rect 1439 591 1440 595
rect 1434 590 1440 591
rect 1442 595 1448 596
rect 1442 591 1443 595
rect 1447 594 1448 595
rect 1451 595 1457 596
rect 1451 594 1452 595
rect 1447 592 1452 594
rect 1447 591 1448 592
rect 1442 590 1448 591
rect 1451 591 1452 592
rect 1456 591 1457 595
rect 1451 590 1457 591
rect 1482 595 1488 596
rect 1482 591 1483 595
rect 1487 594 1488 595
rect 1491 595 1497 596
rect 1491 594 1492 595
rect 1487 592 1492 594
rect 1487 591 1488 592
rect 1482 590 1488 591
rect 1491 591 1492 592
rect 1496 591 1497 595
rect 1491 590 1497 591
rect 1539 595 1545 596
rect 1539 591 1540 595
rect 1544 594 1545 595
rect 1582 595 1588 596
rect 1582 594 1583 595
rect 1544 592 1583 594
rect 1544 591 1545 592
rect 1539 590 1545 591
rect 1582 591 1583 592
rect 1587 591 1588 595
rect 1582 590 1588 591
rect 1590 595 1601 596
rect 1590 591 1591 595
rect 1595 591 1596 595
rect 1600 591 1601 595
rect 1590 590 1601 591
rect 1634 595 1640 596
rect 1634 591 1635 595
rect 1639 594 1640 595
rect 1659 595 1665 596
rect 1659 594 1660 595
rect 1639 592 1660 594
rect 1639 591 1640 592
rect 1634 590 1640 591
rect 1659 591 1660 592
rect 1664 591 1665 595
rect 1659 590 1665 591
rect 1690 595 1696 596
rect 1690 591 1691 595
rect 1695 594 1696 595
rect 1723 595 1729 596
rect 1723 594 1724 595
rect 1695 592 1724 594
rect 1695 591 1696 592
rect 1690 590 1696 591
rect 1723 591 1724 592
rect 1728 591 1729 595
rect 1723 590 1729 591
rect 1787 595 1793 596
rect 1787 591 1788 595
rect 1792 594 1793 595
rect 1823 595 1829 596
rect 1823 594 1824 595
rect 1792 592 1824 594
rect 1792 591 1793 592
rect 1787 590 1793 591
rect 1823 591 1824 592
rect 1828 591 1829 595
rect 1823 590 1829 591
rect 1831 595 1837 596
rect 1831 591 1832 595
rect 1836 594 1837 595
rect 1843 595 1849 596
rect 1843 594 1844 595
rect 1836 592 1844 594
rect 1836 591 1837 592
rect 1831 590 1837 591
rect 1843 591 1844 592
rect 1848 591 1849 595
rect 1843 590 1849 591
rect 1907 595 1913 596
rect 1907 591 1908 595
rect 1912 594 1913 595
rect 1951 595 1957 596
rect 1951 594 1952 595
rect 1912 592 1952 594
rect 1912 591 1913 592
rect 1907 590 1913 591
rect 1951 591 1952 592
rect 1956 591 1957 595
rect 1951 590 1957 591
rect 1971 595 1977 596
rect 1971 591 1972 595
rect 1976 594 1977 595
rect 2014 595 2020 596
rect 2014 594 2015 595
rect 1976 592 2015 594
rect 1976 591 1977 592
rect 1971 590 1977 591
rect 2014 591 2015 592
rect 2019 591 2020 595
rect 2014 590 2020 591
rect 2022 595 2028 596
rect 2022 591 2023 595
rect 2027 594 2028 595
rect 2043 595 2049 596
rect 2043 594 2044 595
rect 2027 592 2044 594
rect 2027 591 2028 592
rect 2022 590 2028 591
rect 2043 591 2044 592
rect 2048 591 2049 595
rect 2043 590 2049 591
rect 2074 595 2080 596
rect 2074 591 2075 595
rect 2079 594 2080 595
rect 2115 595 2121 596
rect 2115 594 2116 595
rect 2079 592 2116 594
rect 2079 591 2080 592
rect 2074 590 2080 591
rect 2115 591 2116 592
rect 2120 591 2121 595
rect 2115 590 2121 591
rect 2146 595 2152 596
rect 2146 591 2147 595
rect 2151 594 2152 595
rect 2195 595 2201 596
rect 2195 594 2196 595
rect 2151 592 2196 594
rect 2151 591 2152 592
rect 2146 590 2152 591
rect 2195 591 2196 592
rect 2200 591 2201 595
rect 2195 590 2201 591
rect 2283 595 2289 596
rect 2283 591 2284 595
rect 2288 594 2289 595
rect 2294 595 2300 596
rect 2294 594 2295 595
rect 2288 592 2295 594
rect 2288 591 2289 592
rect 2283 590 2289 591
rect 2294 591 2295 592
rect 2299 591 2300 595
rect 2294 590 2300 591
rect 2355 595 2361 596
rect 2355 591 2356 595
rect 2360 594 2361 595
rect 2370 595 2376 596
rect 2370 594 2371 595
rect 2360 592 2371 594
rect 2360 591 2361 592
rect 2355 590 2361 591
rect 2370 591 2371 592
rect 2375 591 2376 595
rect 2370 590 2376 591
rect 134 587 140 588
rect 134 583 135 587
rect 139 583 140 587
rect 134 582 140 583
rect 190 587 196 588
rect 190 583 191 587
rect 195 583 196 587
rect 190 582 196 583
rect 270 587 276 588
rect 270 583 271 587
rect 275 583 276 587
rect 270 582 276 583
rect 358 587 364 588
rect 358 583 359 587
rect 363 583 364 587
rect 358 582 364 583
rect 446 587 452 588
rect 446 583 447 587
rect 451 583 452 587
rect 446 582 452 583
rect 534 587 540 588
rect 534 583 535 587
rect 539 583 540 587
rect 534 582 540 583
rect 622 587 628 588
rect 622 583 623 587
rect 627 583 628 587
rect 622 582 628 583
rect 702 587 708 588
rect 702 583 703 587
rect 707 583 708 587
rect 702 582 708 583
rect 782 587 788 588
rect 782 583 783 587
rect 787 583 788 587
rect 782 582 788 583
rect 854 587 860 588
rect 854 583 855 587
rect 859 583 860 587
rect 854 582 860 583
rect 918 587 924 588
rect 918 583 919 587
rect 923 583 924 587
rect 918 582 924 583
rect 974 587 980 588
rect 974 583 975 587
rect 979 583 980 587
rect 974 582 980 583
rect 1022 587 1028 588
rect 1022 583 1023 587
rect 1027 583 1028 587
rect 1022 582 1028 583
rect 1078 587 1084 588
rect 1078 583 1079 587
rect 1083 583 1084 587
rect 1078 582 1084 583
rect 1134 587 1140 588
rect 1134 583 1135 587
rect 1139 583 1140 587
rect 1134 582 1140 583
rect 1190 587 1196 588
rect 1190 583 1191 587
rect 1195 583 1196 587
rect 1190 582 1196 583
rect 1414 587 1420 588
rect 1414 583 1415 587
rect 1419 583 1420 587
rect 1414 582 1420 583
rect 1454 587 1460 588
rect 1454 583 1455 587
rect 1459 583 1460 587
rect 1454 582 1460 583
rect 1494 587 1500 588
rect 1494 583 1495 587
rect 1499 583 1500 587
rect 1494 582 1500 583
rect 1542 587 1548 588
rect 1542 583 1543 587
rect 1547 583 1548 587
rect 1542 582 1548 583
rect 1598 587 1604 588
rect 1598 583 1599 587
rect 1603 583 1604 587
rect 1598 582 1604 583
rect 1662 587 1668 588
rect 1662 583 1663 587
rect 1667 583 1668 587
rect 1662 582 1668 583
rect 1726 587 1732 588
rect 1726 583 1727 587
rect 1731 583 1732 587
rect 1726 582 1732 583
rect 1790 587 1796 588
rect 1790 583 1791 587
rect 1795 583 1796 587
rect 1790 582 1796 583
rect 1846 587 1852 588
rect 1846 583 1847 587
rect 1851 583 1852 587
rect 1846 582 1852 583
rect 1910 587 1916 588
rect 1910 583 1911 587
rect 1915 583 1916 587
rect 1910 582 1916 583
rect 1974 587 1980 588
rect 1974 583 1975 587
rect 1979 583 1980 587
rect 1974 582 1980 583
rect 2046 587 2052 588
rect 2046 583 2047 587
rect 2051 583 2052 587
rect 2046 582 2052 583
rect 2118 587 2124 588
rect 2118 583 2119 587
rect 2123 583 2124 587
rect 2118 582 2124 583
rect 2198 587 2204 588
rect 2198 583 2199 587
rect 2203 583 2204 587
rect 2198 582 2204 583
rect 2286 587 2292 588
rect 2286 583 2287 587
rect 2291 583 2292 587
rect 2286 582 2292 583
rect 2358 587 2364 588
rect 2358 583 2359 587
rect 2363 583 2364 587
rect 2358 582 2364 583
rect 1582 571 1588 572
rect 378 567 384 568
rect 110 564 116 565
rect 110 560 111 564
rect 115 560 116 564
rect 378 563 379 567
rect 383 566 384 567
rect 1434 567 1440 568
rect 383 564 662 566
rect 383 563 384 564
rect 378 562 384 563
rect 110 559 116 560
rect 158 559 165 560
rect 158 555 159 559
rect 164 555 165 559
rect 158 554 165 555
rect 178 559 184 560
rect 178 555 179 559
rect 183 558 184 559
rect 215 559 221 560
rect 215 558 216 559
rect 183 556 216 558
rect 183 555 184 556
rect 178 554 184 555
rect 215 555 216 556
rect 220 555 221 559
rect 215 554 221 555
rect 258 559 264 560
rect 258 555 259 559
rect 263 558 264 559
rect 295 559 301 560
rect 295 558 296 559
rect 263 556 296 558
rect 263 555 264 556
rect 258 554 264 555
rect 295 555 296 556
rect 300 555 301 559
rect 295 554 301 555
rect 383 559 392 560
rect 383 555 384 559
rect 391 555 392 559
rect 383 554 392 555
rect 471 559 480 560
rect 471 555 472 559
rect 479 555 480 559
rect 471 554 480 555
rect 559 559 568 560
rect 559 555 560 559
rect 567 555 568 559
rect 559 554 568 555
rect 647 559 656 560
rect 647 555 648 559
rect 655 555 656 559
rect 660 558 662 564
rect 1238 564 1244 565
rect 1238 560 1239 564
rect 1243 560 1244 564
rect 727 559 733 560
rect 727 558 728 559
rect 660 556 728 558
rect 647 554 656 555
rect 727 555 728 556
rect 732 555 733 559
rect 727 554 733 555
rect 807 559 816 560
rect 807 555 808 559
rect 815 555 816 559
rect 807 554 816 555
rect 879 559 888 560
rect 879 555 880 559
rect 887 555 888 559
rect 879 554 888 555
rect 943 559 952 560
rect 943 555 944 559
rect 951 555 952 559
rect 943 554 952 555
rect 999 559 1008 560
rect 999 555 1000 559
rect 1007 555 1008 559
rect 999 554 1008 555
rect 1047 559 1056 560
rect 1047 555 1048 559
rect 1055 555 1056 559
rect 1047 554 1056 555
rect 1103 559 1112 560
rect 1103 555 1104 559
rect 1111 555 1112 559
rect 1103 554 1112 555
rect 1159 559 1168 560
rect 1159 555 1160 559
rect 1167 555 1168 559
rect 1159 554 1168 555
rect 1214 559 1221 560
rect 1238 559 1244 560
rect 1278 564 1284 565
rect 1278 560 1279 564
rect 1283 560 1284 564
rect 1434 563 1435 567
rect 1439 566 1440 567
rect 1582 567 1583 571
rect 1587 570 1588 571
rect 1823 571 1829 572
rect 1587 568 1702 570
rect 1587 567 1588 568
rect 1582 566 1588 567
rect 1439 564 1570 566
rect 1439 563 1440 564
rect 1434 562 1440 563
rect 1568 560 1570 564
rect 1634 563 1640 564
rect 1634 562 1635 563
rect 1623 561 1635 562
rect 1278 559 1284 560
rect 1439 559 1448 560
rect 1214 555 1215 559
rect 1220 555 1221 559
rect 1214 554 1221 555
rect 1439 555 1440 559
rect 1447 555 1448 559
rect 1439 554 1448 555
rect 1479 559 1488 560
rect 1479 555 1480 559
rect 1487 555 1488 559
rect 1479 554 1488 555
rect 1519 559 1525 560
rect 1519 555 1520 559
rect 1524 558 1525 559
rect 1558 559 1564 560
rect 1558 558 1559 559
rect 1524 556 1559 558
rect 1524 555 1525 556
rect 1519 554 1525 555
rect 1558 555 1559 556
rect 1563 555 1564 559
rect 1558 554 1564 555
rect 1567 559 1573 560
rect 1567 555 1568 559
rect 1572 555 1573 559
rect 1623 557 1624 561
rect 1628 560 1635 561
rect 1628 557 1629 560
rect 1634 559 1635 560
rect 1639 559 1640 563
rect 1634 558 1640 559
rect 1687 559 1696 560
rect 1623 556 1629 557
rect 1567 554 1573 555
rect 1687 555 1688 559
rect 1695 555 1696 559
rect 1700 558 1702 568
rect 1823 567 1824 571
rect 1828 570 1829 571
rect 1828 568 1906 570
rect 1828 567 1829 568
rect 1823 566 1829 567
rect 1831 563 1837 564
rect 1831 562 1832 563
rect 1815 561 1832 562
rect 1751 559 1757 560
rect 1751 558 1752 559
rect 1700 556 1752 558
rect 1687 554 1696 555
rect 1751 555 1752 556
rect 1756 555 1757 559
rect 1815 557 1816 561
rect 1820 560 1832 561
rect 1820 557 1821 560
rect 1831 559 1832 560
rect 1836 559 1837 563
rect 1831 558 1837 559
rect 1871 559 1877 560
rect 1815 556 1821 557
rect 1751 554 1757 555
rect 1871 555 1872 559
rect 1876 558 1877 559
rect 1894 559 1900 560
rect 1894 558 1895 559
rect 1876 556 1895 558
rect 1876 555 1877 556
rect 1871 554 1877 555
rect 1894 555 1895 556
rect 1899 555 1900 559
rect 1904 558 1906 568
rect 2014 567 2020 568
rect 2014 563 2015 567
rect 2019 566 2020 567
rect 2019 564 2158 566
rect 2019 563 2020 564
rect 2014 562 2020 563
rect 1935 559 1941 560
rect 1935 558 1936 559
rect 1904 556 1936 558
rect 1894 554 1900 555
rect 1935 555 1936 556
rect 1940 555 1941 559
rect 1935 554 1941 555
rect 1951 559 1957 560
rect 1951 555 1952 559
rect 1956 558 1957 559
rect 1999 559 2005 560
rect 1999 558 2000 559
rect 1956 556 2000 558
rect 1956 555 1957 556
rect 1951 554 1957 555
rect 1999 555 2000 556
rect 2004 555 2005 559
rect 1999 554 2005 555
rect 2071 559 2080 560
rect 2071 555 2072 559
rect 2079 555 2080 559
rect 2071 554 2080 555
rect 2143 559 2152 560
rect 2143 555 2144 559
rect 2151 555 2152 559
rect 2156 558 2158 564
rect 2406 564 2412 565
rect 2406 560 2407 564
rect 2411 560 2412 564
rect 2223 559 2229 560
rect 2223 558 2224 559
rect 2156 556 2224 558
rect 2143 554 2152 555
rect 2223 555 2224 556
rect 2228 555 2229 559
rect 2223 554 2229 555
rect 2302 559 2308 560
rect 2302 555 2303 559
rect 2307 558 2308 559
rect 2311 559 2317 560
rect 2311 558 2312 559
rect 2307 556 2312 558
rect 2307 555 2308 556
rect 2302 554 2308 555
rect 2311 555 2312 556
rect 2316 555 2317 559
rect 2311 554 2317 555
rect 2374 559 2380 560
rect 2374 555 2375 559
rect 2379 558 2380 559
rect 2383 559 2389 560
rect 2406 559 2412 560
rect 2383 558 2384 559
rect 2379 556 2384 558
rect 2379 555 2380 556
rect 2374 554 2380 555
rect 2383 555 2384 556
rect 2388 555 2389 559
rect 2383 554 2389 555
rect 110 547 116 548
rect 110 543 111 547
rect 115 543 116 547
rect 110 542 116 543
rect 1238 547 1244 548
rect 1238 543 1239 547
rect 1243 543 1244 547
rect 1238 542 1244 543
rect 1278 547 1284 548
rect 1278 543 1279 547
rect 1283 543 1284 547
rect 1278 542 1284 543
rect 2406 547 2412 548
rect 2406 543 2407 547
rect 2411 543 2412 547
rect 2406 542 2412 543
rect 134 540 140 541
rect 134 536 135 540
rect 139 536 140 540
rect 134 535 140 536
rect 190 540 196 541
rect 190 536 191 540
rect 195 536 196 540
rect 190 535 196 536
rect 270 540 276 541
rect 270 536 271 540
rect 275 536 276 540
rect 270 535 276 536
rect 358 540 364 541
rect 358 536 359 540
rect 363 536 364 540
rect 358 535 364 536
rect 446 540 452 541
rect 446 536 447 540
rect 451 536 452 540
rect 446 535 452 536
rect 534 540 540 541
rect 534 536 535 540
rect 539 536 540 540
rect 534 535 540 536
rect 622 540 628 541
rect 622 536 623 540
rect 627 536 628 540
rect 622 535 628 536
rect 702 540 708 541
rect 702 536 703 540
rect 707 536 708 540
rect 702 535 708 536
rect 782 540 788 541
rect 782 536 783 540
rect 787 536 788 540
rect 782 535 788 536
rect 854 540 860 541
rect 854 536 855 540
rect 859 536 860 540
rect 854 535 860 536
rect 918 540 924 541
rect 918 536 919 540
rect 923 536 924 540
rect 918 535 924 536
rect 974 540 980 541
rect 974 536 975 540
rect 979 536 980 540
rect 974 535 980 536
rect 1022 540 1028 541
rect 1022 536 1023 540
rect 1027 536 1028 540
rect 1022 535 1028 536
rect 1078 540 1084 541
rect 1078 536 1079 540
rect 1083 536 1084 540
rect 1078 535 1084 536
rect 1134 540 1140 541
rect 1134 536 1135 540
rect 1139 536 1140 540
rect 1134 535 1140 536
rect 1190 540 1196 541
rect 1190 536 1191 540
rect 1195 536 1196 540
rect 1190 535 1196 536
rect 1414 540 1420 541
rect 1414 536 1415 540
rect 1419 536 1420 540
rect 1414 535 1420 536
rect 1454 540 1460 541
rect 1454 536 1455 540
rect 1459 536 1460 540
rect 1454 535 1460 536
rect 1494 540 1500 541
rect 1494 536 1495 540
rect 1499 536 1500 540
rect 1494 535 1500 536
rect 1542 540 1548 541
rect 1542 536 1543 540
rect 1547 536 1548 540
rect 1542 535 1548 536
rect 1598 540 1604 541
rect 1598 536 1599 540
rect 1603 536 1604 540
rect 1598 535 1604 536
rect 1662 540 1668 541
rect 1662 536 1663 540
rect 1667 536 1668 540
rect 1662 535 1668 536
rect 1726 540 1732 541
rect 1726 536 1727 540
rect 1731 536 1732 540
rect 1726 535 1732 536
rect 1790 540 1796 541
rect 1790 536 1791 540
rect 1795 536 1796 540
rect 1790 535 1796 536
rect 1846 540 1852 541
rect 1846 536 1847 540
rect 1851 536 1852 540
rect 1846 535 1852 536
rect 1910 540 1916 541
rect 1910 536 1911 540
rect 1915 536 1916 540
rect 1910 535 1916 536
rect 1974 540 1980 541
rect 1974 536 1975 540
rect 1979 536 1980 540
rect 1974 535 1980 536
rect 2046 540 2052 541
rect 2046 536 2047 540
rect 2051 536 2052 540
rect 2046 535 2052 536
rect 2118 540 2124 541
rect 2118 536 2119 540
rect 2123 536 2124 540
rect 2118 535 2124 536
rect 2198 540 2204 541
rect 2198 536 2199 540
rect 2203 536 2204 540
rect 2198 535 2204 536
rect 2286 540 2292 541
rect 2286 536 2287 540
rect 2291 536 2292 540
rect 2286 535 2292 536
rect 2358 540 2364 541
rect 2358 536 2359 540
rect 2363 536 2364 540
rect 2358 535 2364 536
rect 1302 528 1308 529
rect 1302 524 1303 528
rect 1307 524 1308 528
rect 1302 523 1308 524
rect 1374 528 1380 529
rect 1374 524 1375 528
rect 1379 524 1380 528
rect 1374 523 1380 524
rect 1478 528 1484 529
rect 1478 524 1479 528
rect 1483 524 1484 528
rect 1478 523 1484 524
rect 1582 528 1588 529
rect 1582 524 1583 528
rect 1587 524 1588 528
rect 1582 523 1588 524
rect 1694 528 1700 529
rect 1694 524 1695 528
rect 1699 524 1700 528
rect 1694 523 1700 524
rect 1798 528 1804 529
rect 1798 524 1799 528
rect 1803 524 1804 528
rect 1798 523 1804 524
rect 1902 528 1908 529
rect 1902 524 1903 528
rect 1907 524 1908 528
rect 1902 523 1908 524
rect 2006 528 2012 529
rect 2006 524 2007 528
rect 2011 524 2012 528
rect 2006 523 2012 524
rect 2102 528 2108 529
rect 2102 524 2103 528
rect 2107 524 2108 528
rect 2102 523 2108 524
rect 2190 528 2196 529
rect 2190 524 2191 528
rect 2195 524 2196 528
rect 2190 523 2196 524
rect 2286 528 2292 529
rect 2286 524 2287 528
rect 2291 524 2292 528
rect 2286 523 2292 524
rect 2358 528 2364 529
rect 2358 524 2359 528
rect 2363 524 2364 528
rect 2358 523 2364 524
rect 1278 521 1284 522
rect 134 520 140 521
rect 134 516 135 520
rect 139 516 140 520
rect 134 515 140 516
rect 190 520 196 521
rect 190 516 191 520
rect 195 516 196 520
rect 190 515 196 516
rect 262 520 268 521
rect 262 516 263 520
rect 267 516 268 520
rect 262 515 268 516
rect 334 520 340 521
rect 334 516 335 520
rect 339 516 340 520
rect 334 515 340 516
rect 414 520 420 521
rect 414 516 415 520
rect 419 516 420 520
rect 414 515 420 516
rect 494 520 500 521
rect 494 516 495 520
rect 499 516 500 520
rect 494 515 500 516
rect 574 520 580 521
rect 574 516 575 520
rect 579 516 580 520
rect 574 515 580 516
rect 646 520 652 521
rect 646 516 647 520
rect 651 516 652 520
rect 646 515 652 516
rect 718 520 724 521
rect 718 516 719 520
rect 723 516 724 520
rect 718 515 724 516
rect 782 520 788 521
rect 782 516 783 520
rect 787 516 788 520
rect 782 515 788 516
rect 846 520 852 521
rect 846 516 847 520
rect 851 516 852 520
rect 846 515 852 516
rect 902 520 908 521
rect 902 516 903 520
rect 907 516 908 520
rect 902 515 908 516
rect 958 520 964 521
rect 958 516 959 520
rect 963 516 964 520
rect 958 515 964 516
rect 1022 520 1028 521
rect 1022 516 1023 520
rect 1027 516 1028 520
rect 1022 515 1028 516
rect 1086 520 1092 521
rect 1086 516 1087 520
rect 1091 516 1092 520
rect 1086 515 1092 516
rect 1150 520 1156 521
rect 1150 516 1151 520
rect 1155 516 1156 520
rect 1150 515 1156 516
rect 1190 520 1196 521
rect 1190 516 1191 520
rect 1195 516 1196 520
rect 1278 517 1279 521
rect 1283 517 1284 521
rect 1278 516 1284 517
rect 2406 521 2412 522
rect 2406 517 2407 521
rect 2411 517 2412 521
rect 2406 516 2412 517
rect 1190 515 1196 516
rect 110 513 116 514
rect 110 509 111 513
rect 115 509 116 513
rect 110 508 116 509
rect 1238 513 1244 514
rect 1238 509 1239 513
rect 1243 509 1244 513
rect 1238 508 1244 509
rect 802 507 808 508
rect 802 503 803 507
rect 807 506 808 507
rect 1310 507 1316 508
rect 807 504 1026 506
rect 807 503 808 504
rect 802 502 808 503
rect 159 499 165 500
rect 110 496 116 497
rect 110 492 111 496
rect 115 492 116 496
rect 159 495 160 499
rect 164 498 165 499
rect 175 499 181 500
rect 175 498 176 499
rect 164 496 176 498
rect 164 495 165 496
rect 159 494 165 495
rect 175 495 176 496
rect 180 495 181 499
rect 175 494 181 495
rect 215 499 221 500
rect 215 495 216 499
rect 220 498 221 499
rect 254 499 260 500
rect 254 498 255 499
rect 220 496 255 498
rect 220 495 221 496
rect 215 494 221 495
rect 254 495 255 496
rect 259 495 260 499
rect 254 494 260 495
rect 286 499 293 500
rect 286 495 287 499
rect 292 495 293 499
rect 286 494 293 495
rect 342 499 348 500
rect 342 495 343 499
rect 347 498 348 499
rect 359 499 365 500
rect 359 498 360 499
rect 347 496 360 498
rect 347 495 348 496
rect 342 494 348 495
rect 359 495 360 496
rect 364 495 365 499
rect 359 494 365 495
rect 367 499 373 500
rect 367 495 368 499
rect 372 498 373 499
rect 439 499 445 500
rect 439 498 440 499
rect 372 496 440 498
rect 372 495 373 496
rect 367 494 373 495
rect 439 495 440 496
rect 444 495 445 499
rect 439 494 445 495
rect 447 499 453 500
rect 447 495 448 499
rect 452 498 453 499
rect 519 499 525 500
rect 519 498 520 499
rect 452 496 520 498
rect 452 495 453 496
rect 447 494 453 495
rect 519 495 520 496
rect 524 495 525 499
rect 519 494 525 495
rect 527 499 533 500
rect 527 495 528 499
rect 532 498 533 499
rect 599 499 605 500
rect 599 498 600 499
rect 532 496 600 498
rect 532 495 533 496
rect 527 494 533 495
rect 599 495 600 496
rect 604 495 605 499
rect 599 494 605 495
rect 671 499 677 500
rect 671 495 672 499
rect 676 498 677 499
rect 710 499 716 500
rect 710 498 711 499
rect 676 496 711 498
rect 676 495 677 496
rect 671 494 677 495
rect 710 495 711 496
rect 715 495 716 499
rect 710 494 716 495
rect 743 499 749 500
rect 743 495 744 499
rect 748 498 749 499
rect 767 499 773 500
rect 767 498 768 499
rect 748 496 768 498
rect 748 495 749 496
rect 743 494 749 495
rect 767 495 768 496
rect 772 495 773 499
rect 767 494 773 495
rect 807 499 813 500
rect 807 495 808 499
rect 812 498 813 499
rect 838 499 844 500
rect 838 498 839 499
rect 812 496 839 498
rect 812 495 813 496
rect 807 494 813 495
rect 838 495 839 496
rect 843 495 844 499
rect 838 494 844 495
rect 871 499 877 500
rect 871 495 872 499
rect 876 498 877 499
rect 894 499 900 500
rect 894 498 895 499
rect 876 496 895 498
rect 876 495 877 496
rect 871 494 877 495
rect 894 495 895 496
rect 899 495 900 499
rect 894 494 900 495
rect 927 499 933 500
rect 927 495 928 499
rect 932 498 933 499
rect 950 499 956 500
rect 950 498 951 499
rect 932 496 951 498
rect 932 495 933 496
rect 927 494 933 495
rect 950 495 951 496
rect 955 495 956 499
rect 950 494 956 495
rect 983 499 989 500
rect 983 495 984 499
rect 988 498 989 499
rect 1014 499 1020 500
rect 1014 498 1015 499
rect 988 496 1015 498
rect 988 495 989 496
rect 983 494 989 495
rect 1014 495 1015 496
rect 1019 495 1020 499
rect 1024 498 1026 504
rect 1278 504 1284 505
rect 1278 500 1279 504
rect 1283 500 1284 504
rect 1310 503 1311 507
rect 1315 506 1316 507
rect 1327 507 1333 508
rect 1327 506 1328 507
rect 1315 504 1328 506
rect 1315 503 1316 504
rect 1310 502 1316 503
rect 1327 503 1328 504
rect 1332 503 1333 507
rect 1399 507 1405 508
rect 1399 506 1400 507
rect 1327 502 1333 503
rect 1336 504 1400 506
rect 1047 499 1053 500
rect 1047 498 1048 499
rect 1024 496 1048 498
rect 1014 494 1020 495
rect 1047 495 1048 496
rect 1052 495 1053 499
rect 1047 494 1053 495
rect 1111 499 1117 500
rect 1111 495 1112 499
rect 1116 498 1117 499
rect 1142 499 1148 500
rect 1142 498 1143 499
rect 1116 496 1143 498
rect 1116 495 1117 496
rect 1111 494 1117 495
rect 1142 495 1143 496
rect 1147 495 1148 499
rect 1142 494 1148 495
rect 1175 499 1184 500
rect 1175 495 1176 499
rect 1183 495 1184 499
rect 1175 494 1184 495
rect 1215 499 1221 500
rect 1215 495 1216 499
rect 1220 498 1221 499
rect 1230 499 1236 500
rect 1278 499 1284 500
rect 1230 498 1231 499
rect 1220 496 1231 498
rect 1220 495 1221 496
rect 1215 494 1221 495
rect 1230 495 1231 496
rect 1235 495 1236 499
rect 1230 494 1236 495
rect 1238 496 1244 497
rect 110 491 116 492
rect 1238 492 1239 496
rect 1243 492 1244 496
rect 1238 491 1244 492
rect 1336 490 1338 504
rect 1399 503 1400 504
rect 1404 503 1405 507
rect 1399 502 1405 503
rect 1407 507 1413 508
rect 1407 503 1408 507
rect 1412 506 1413 507
rect 1503 507 1509 508
rect 1503 506 1504 507
rect 1412 504 1504 506
rect 1412 503 1413 504
rect 1407 502 1413 503
rect 1503 503 1504 504
rect 1508 503 1509 507
rect 1503 502 1509 503
rect 1511 507 1517 508
rect 1511 503 1512 507
rect 1516 506 1517 507
rect 1607 507 1613 508
rect 1607 506 1608 507
rect 1516 504 1608 506
rect 1516 503 1517 504
rect 1511 502 1517 503
rect 1607 503 1608 504
rect 1612 503 1613 507
rect 1607 502 1613 503
rect 1719 507 1728 508
rect 1719 503 1720 507
rect 1727 503 1728 507
rect 1719 502 1728 503
rect 1730 507 1736 508
rect 1730 503 1731 507
rect 1735 506 1736 507
rect 1823 507 1829 508
rect 1823 506 1824 507
rect 1735 504 1824 506
rect 1735 503 1736 504
rect 1730 502 1736 503
rect 1823 503 1824 504
rect 1828 503 1829 507
rect 1823 502 1829 503
rect 1927 507 1933 508
rect 1927 503 1928 507
rect 1932 506 1933 507
rect 1998 507 2004 508
rect 1998 506 1999 507
rect 1932 504 1999 506
rect 1932 503 1933 504
rect 1927 502 1933 503
rect 1998 503 1999 504
rect 2003 503 2004 507
rect 2031 507 2037 508
rect 2031 506 2032 507
rect 1998 502 2004 503
rect 2016 504 2032 506
rect 1806 499 1812 500
rect 1806 495 1807 499
rect 1811 498 1812 499
rect 2016 498 2018 504
rect 2031 503 2032 504
rect 2036 503 2037 507
rect 2031 502 2037 503
rect 2127 507 2133 508
rect 2127 503 2128 507
rect 2132 506 2133 507
rect 2182 507 2188 508
rect 2182 506 2183 507
rect 2132 504 2183 506
rect 2132 503 2133 504
rect 2127 502 2133 503
rect 2182 503 2183 504
rect 2187 503 2188 507
rect 2182 502 2188 503
rect 2215 507 2221 508
rect 2215 503 2216 507
rect 2220 506 2221 507
rect 2278 507 2284 508
rect 2278 506 2279 507
rect 2220 504 2279 506
rect 2220 503 2221 504
rect 2215 502 2221 503
rect 2278 503 2279 504
rect 2283 503 2284 507
rect 2278 502 2284 503
rect 2294 507 2300 508
rect 2294 503 2295 507
rect 2299 506 2300 507
rect 2311 507 2317 508
rect 2311 506 2312 507
rect 2299 504 2312 506
rect 2299 503 2300 504
rect 2294 502 2300 503
rect 2311 503 2312 504
rect 2316 503 2317 507
rect 2311 502 2317 503
rect 2366 507 2372 508
rect 2366 503 2367 507
rect 2371 506 2372 507
rect 2383 507 2389 508
rect 2383 506 2384 507
rect 2371 504 2384 506
rect 2371 503 2372 504
rect 2366 502 2372 503
rect 2383 503 2384 504
rect 2388 503 2389 507
rect 2383 502 2389 503
rect 2406 504 2412 505
rect 2406 500 2407 504
rect 2411 500 2412 504
rect 2406 499 2412 500
rect 1811 496 2018 498
rect 1811 495 1812 496
rect 1806 494 1812 495
rect 1280 488 1338 490
rect 1094 487 1100 488
rect 1094 483 1095 487
rect 1099 486 1100 487
rect 1280 486 1282 488
rect 1099 484 1282 486
rect 1099 483 1100 484
rect 1094 482 1100 483
rect 1302 481 1308 482
rect 1302 477 1303 481
rect 1307 477 1308 481
rect 1302 476 1308 477
rect 1374 481 1380 482
rect 1374 477 1375 481
rect 1379 477 1380 481
rect 1374 476 1380 477
rect 1478 481 1484 482
rect 1478 477 1479 481
rect 1483 477 1484 481
rect 1478 476 1484 477
rect 1582 481 1588 482
rect 1582 477 1583 481
rect 1587 477 1588 481
rect 1582 476 1588 477
rect 1694 481 1700 482
rect 1694 477 1695 481
rect 1699 477 1700 481
rect 1694 476 1700 477
rect 1798 481 1804 482
rect 1798 477 1799 481
rect 1803 477 1804 481
rect 1798 476 1804 477
rect 1902 481 1908 482
rect 1902 477 1903 481
rect 1907 477 1908 481
rect 1902 476 1908 477
rect 2006 481 2012 482
rect 2006 477 2007 481
rect 2011 477 2012 481
rect 2006 476 2012 477
rect 2102 481 2108 482
rect 2102 477 2103 481
rect 2107 477 2108 481
rect 2102 476 2108 477
rect 2190 481 2196 482
rect 2190 477 2191 481
rect 2195 477 2196 481
rect 2190 476 2196 477
rect 2286 481 2292 482
rect 2286 477 2287 481
rect 2291 477 2292 481
rect 2286 476 2292 477
rect 2358 481 2364 482
rect 2358 477 2359 481
rect 2363 477 2364 481
rect 2358 476 2364 477
rect 134 473 140 474
rect 134 469 135 473
rect 139 469 140 473
rect 134 468 140 469
rect 190 473 196 474
rect 190 469 191 473
rect 195 469 196 473
rect 190 468 196 469
rect 262 473 268 474
rect 262 469 263 473
rect 267 469 268 473
rect 262 468 268 469
rect 334 473 340 474
rect 334 469 335 473
rect 339 469 340 473
rect 334 468 340 469
rect 414 473 420 474
rect 414 469 415 473
rect 419 469 420 473
rect 414 468 420 469
rect 494 473 500 474
rect 494 469 495 473
rect 499 469 500 473
rect 494 468 500 469
rect 574 473 580 474
rect 574 469 575 473
rect 579 469 580 473
rect 574 468 580 469
rect 646 473 652 474
rect 646 469 647 473
rect 651 469 652 473
rect 646 468 652 469
rect 718 473 724 474
rect 718 469 719 473
rect 723 469 724 473
rect 718 468 724 469
rect 782 473 788 474
rect 782 469 783 473
rect 787 469 788 473
rect 782 468 788 469
rect 846 473 852 474
rect 846 469 847 473
rect 851 469 852 473
rect 846 468 852 469
rect 902 473 908 474
rect 902 469 903 473
rect 907 469 908 473
rect 902 468 908 469
rect 958 473 964 474
rect 958 469 959 473
rect 963 469 964 473
rect 958 468 964 469
rect 1022 473 1028 474
rect 1022 469 1023 473
rect 1027 469 1028 473
rect 1022 468 1028 469
rect 1086 473 1092 474
rect 1086 469 1087 473
rect 1091 469 1092 473
rect 1086 468 1092 469
rect 1150 473 1156 474
rect 1150 469 1151 473
rect 1155 469 1156 473
rect 1150 468 1156 469
rect 1190 473 1196 474
rect 1190 469 1191 473
rect 1195 469 1196 473
rect 1190 468 1196 469
rect 1230 471 1236 472
rect 562 467 568 468
rect 131 463 137 464
rect 131 459 132 463
rect 136 462 137 463
rect 167 463 173 464
rect 167 462 168 463
rect 136 460 168 462
rect 136 459 137 460
rect 131 458 137 459
rect 167 459 168 460
rect 172 459 173 463
rect 167 458 173 459
rect 175 463 181 464
rect 175 459 176 463
rect 180 462 181 463
rect 187 463 193 464
rect 187 462 188 463
rect 180 460 188 462
rect 180 459 181 460
rect 175 458 181 459
rect 187 459 188 460
rect 192 459 193 463
rect 187 458 193 459
rect 254 463 265 464
rect 254 459 255 463
rect 259 459 260 463
rect 264 459 265 463
rect 254 458 265 459
rect 331 463 337 464
rect 331 459 332 463
rect 336 462 337 463
rect 367 463 373 464
rect 367 462 368 463
rect 336 460 368 462
rect 336 459 337 460
rect 331 458 337 459
rect 367 459 368 460
rect 372 459 373 463
rect 367 458 373 459
rect 411 463 417 464
rect 411 459 412 463
rect 416 462 417 463
rect 447 463 453 464
rect 447 462 448 463
rect 416 460 448 462
rect 416 459 417 460
rect 411 458 417 459
rect 447 459 448 460
rect 452 459 453 463
rect 447 458 453 459
rect 491 463 497 464
rect 491 459 492 463
rect 496 462 497 463
rect 527 463 533 464
rect 527 462 528 463
rect 496 460 528 462
rect 496 459 497 460
rect 491 458 497 459
rect 527 459 528 460
rect 532 459 533 463
rect 562 463 563 467
rect 567 466 568 467
rect 1230 467 1231 471
rect 1235 470 1236 471
rect 1299 471 1305 472
rect 1299 470 1300 471
rect 1235 468 1300 470
rect 1235 467 1236 468
rect 1230 466 1236 467
rect 1299 467 1300 468
rect 1304 467 1305 471
rect 1299 466 1305 467
rect 1371 471 1377 472
rect 1371 467 1372 471
rect 1376 470 1377 471
rect 1407 471 1413 472
rect 1407 470 1408 471
rect 1376 468 1408 470
rect 1376 467 1377 468
rect 1371 466 1377 467
rect 1407 467 1408 468
rect 1412 467 1413 471
rect 1407 466 1413 467
rect 1475 471 1481 472
rect 1475 467 1476 471
rect 1480 470 1481 471
rect 1511 471 1517 472
rect 1511 470 1512 471
rect 1480 468 1512 470
rect 1480 467 1481 468
rect 1475 466 1481 467
rect 1511 467 1512 468
rect 1516 467 1517 471
rect 1511 466 1517 467
rect 1558 471 1564 472
rect 1558 467 1559 471
rect 1563 470 1564 471
rect 1579 471 1585 472
rect 1579 470 1580 471
rect 1563 468 1580 470
rect 1563 467 1564 468
rect 1558 466 1564 467
rect 1579 467 1580 468
rect 1584 467 1585 471
rect 1579 466 1585 467
rect 1691 471 1697 472
rect 1691 467 1692 471
rect 1696 470 1697 471
rect 1730 471 1736 472
rect 1730 470 1731 471
rect 1696 468 1731 470
rect 1696 467 1697 468
rect 1691 466 1697 467
rect 1730 467 1731 468
rect 1735 467 1736 471
rect 1730 466 1736 467
rect 1795 471 1801 472
rect 1795 467 1796 471
rect 1800 470 1801 471
rect 1806 471 1812 472
rect 1806 470 1807 471
rect 1800 468 1807 470
rect 1800 467 1801 468
rect 1795 466 1801 467
rect 1806 467 1807 468
rect 1811 467 1812 471
rect 1806 466 1812 467
rect 1894 471 1905 472
rect 1894 467 1895 471
rect 1899 467 1900 471
rect 1904 467 1905 471
rect 1894 466 1905 467
rect 1998 471 2009 472
rect 1998 467 1999 471
rect 2003 467 2004 471
rect 2008 467 2009 471
rect 1998 466 2009 467
rect 2099 471 2105 472
rect 2099 467 2100 471
rect 2104 470 2105 471
rect 2174 471 2180 472
rect 2174 470 2175 471
rect 2104 468 2175 470
rect 2104 467 2105 468
rect 2099 466 2105 467
rect 2174 467 2175 468
rect 2179 467 2180 471
rect 2174 466 2180 467
rect 2182 471 2193 472
rect 2182 467 2183 471
rect 2187 467 2188 471
rect 2192 467 2193 471
rect 2182 466 2193 467
rect 2278 471 2289 472
rect 2278 467 2279 471
rect 2283 467 2284 471
rect 2288 467 2289 471
rect 2278 466 2289 467
rect 2355 471 2361 472
rect 2355 467 2356 471
rect 2360 470 2361 471
rect 2374 471 2380 472
rect 2374 470 2375 471
rect 2360 468 2375 470
rect 2360 467 2361 468
rect 2355 466 2361 467
rect 2374 467 2375 468
rect 2379 467 2380 471
rect 2374 466 2380 467
rect 567 465 577 466
rect 567 464 572 465
rect 567 463 568 464
rect 562 462 568 463
rect 571 461 572 464
rect 576 461 577 465
rect 571 460 577 461
rect 643 463 649 464
rect 527 458 533 459
rect 643 459 644 463
rect 648 462 649 463
rect 690 463 696 464
rect 690 462 691 463
rect 648 460 691 462
rect 648 459 649 460
rect 643 458 649 459
rect 690 459 691 460
rect 695 459 696 463
rect 690 458 696 459
rect 710 463 721 464
rect 710 459 711 463
rect 715 459 716 463
rect 720 459 721 463
rect 710 458 721 459
rect 767 463 773 464
rect 767 459 768 463
rect 772 462 773 463
rect 779 463 785 464
rect 779 462 780 463
rect 772 460 780 462
rect 772 459 773 460
rect 767 458 773 459
rect 779 459 780 460
rect 784 459 785 463
rect 779 458 785 459
rect 838 463 849 464
rect 838 459 839 463
rect 843 459 844 463
rect 848 459 849 463
rect 838 458 849 459
rect 894 463 905 464
rect 894 459 895 463
rect 899 459 900 463
rect 904 459 905 463
rect 894 458 905 459
rect 950 463 961 464
rect 950 459 951 463
rect 955 459 956 463
rect 960 459 961 463
rect 950 458 961 459
rect 1014 463 1025 464
rect 1014 459 1015 463
rect 1019 459 1020 463
rect 1024 459 1025 463
rect 1014 458 1025 459
rect 1083 463 1089 464
rect 1083 459 1084 463
rect 1088 462 1089 463
rect 1094 463 1100 464
rect 1094 462 1095 463
rect 1088 460 1095 462
rect 1088 459 1089 460
rect 1083 458 1089 459
rect 1094 459 1095 460
rect 1099 459 1100 463
rect 1094 458 1100 459
rect 1142 463 1153 464
rect 1142 459 1143 463
rect 1147 459 1148 463
rect 1152 459 1153 463
rect 1142 458 1153 459
rect 1178 463 1184 464
rect 1178 459 1179 463
rect 1183 462 1184 463
rect 1187 463 1193 464
rect 1187 462 1188 463
rect 1183 460 1188 462
rect 1183 459 1184 460
rect 1178 458 1184 459
rect 1187 459 1188 460
rect 1192 459 1193 463
rect 1187 458 1193 459
rect 1299 455 1305 456
rect 179 451 185 452
rect 179 447 180 451
rect 184 450 185 451
rect 210 451 216 452
rect 210 450 211 451
rect 184 448 211 450
rect 184 447 185 448
rect 179 446 185 447
rect 210 447 211 448
rect 215 447 216 451
rect 210 446 216 447
rect 219 451 225 452
rect 219 447 220 451
rect 224 450 225 451
rect 250 451 256 452
rect 250 450 251 451
rect 224 448 251 450
rect 224 447 225 448
rect 219 446 225 447
rect 250 447 251 448
rect 255 447 256 451
rect 250 446 256 447
rect 259 451 265 452
rect 259 447 260 451
rect 264 450 265 451
rect 298 451 304 452
rect 298 450 299 451
rect 264 448 299 450
rect 264 447 265 448
rect 259 446 265 447
rect 298 447 299 448
rect 303 447 304 451
rect 298 446 304 447
rect 307 451 313 452
rect 307 447 308 451
rect 312 450 313 451
rect 342 451 348 452
rect 342 450 343 451
rect 312 448 343 450
rect 312 447 313 448
rect 307 446 313 447
rect 342 447 343 448
rect 347 447 348 451
rect 342 446 348 447
rect 350 451 356 452
rect 350 447 351 451
rect 355 450 356 451
rect 363 451 369 452
rect 363 450 364 451
rect 355 448 364 450
rect 355 447 356 448
rect 350 446 356 447
rect 363 447 364 448
rect 368 447 369 451
rect 363 446 369 447
rect 394 451 400 452
rect 394 447 395 451
rect 399 450 400 451
rect 427 451 433 452
rect 427 450 428 451
rect 399 448 428 450
rect 399 447 400 448
rect 394 446 400 447
rect 427 447 428 448
rect 432 447 433 451
rect 427 446 433 447
rect 458 451 464 452
rect 458 447 459 451
rect 463 450 464 451
rect 491 451 497 452
rect 491 450 492 451
rect 463 448 492 450
rect 463 447 464 448
rect 458 446 464 447
rect 491 447 492 448
rect 496 447 497 451
rect 491 446 497 447
rect 555 451 561 452
rect 555 447 556 451
rect 560 450 561 451
rect 566 451 572 452
rect 566 450 567 451
rect 560 448 567 450
rect 560 447 561 448
rect 555 446 561 447
rect 566 447 567 448
rect 571 447 572 451
rect 566 446 572 447
rect 586 451 592 452
rect 586 447 587 451
rect 591 450 592 451
rect 611 451 617 452
rect 611 450 612 451
rect 591 448 612 450
rect 591 447 592 448
rect 586 446 592 447
rect 611 447 612 448
rect 616 447 617 451
rect 611 446 617 447
rect 647 451 653 452
rect 647 447 648 451
rect 652 450 653 451
rect 667 451 673 452
rect 667 450 668 451
rect 652 448 668 450
rect 652 447 653 448
rect 647 446 653 447
rect 667 447 668 448
rect 672 447 673 451
rect 667 446 673 447
rect 698 451 704 452
rect 698 447 699 451
rect 703 450 704 451
rect 715 451 721 452
rect 715 450 716 451
rect 703 448 716 450
rect 703 447 704 448
rect 698 446 704 447
rect 715 447 716 448
rect 720 447 721 451
rect 715 446 721 447
rect 759 451 765 452
rect 759 447 760 451
rect 764 450 765 451
rect 771 451 777 452
rect 771 450 772 451
rect 764 448 772 450
rect 764 447 765 448
rect 759 446 765 447
rect 771 447 772 448
rect 776 447 777 451
rect 771 446 777 447
rect 802 451 808 452
rect 802 447 803 451
rect 807 450 808 451
rect 827 451 833 452
rect 827 450 828 451
rect 807 448 828 450
rect 807 447 808 448
rect 802 446 808 447
rect 827 447 828 448
rect 832 447 833 451
rect 827 446 833 447
rect 858 451 864 452
rect 858 447 859 451
rect 863 450 864 451
rect 883 451 889 452
rect 883 450 884 451
rect 863 448 884 450
rect 863 447 864 448
rect 858 446 864 447
rect 883 447 884 448
rect 888 447 889 451
rect 1299 451 1300 455
rect 1304 454 1305 455
rect 1310 455 1316 456
rect 1310 454 1311 455
rect 1304 452 1311 454
rect 1304 451 1305 452
rect 1299 450 1305 451
rect 1310 451 1311 452
rect 1315 451 1316 455
rect 1310 450 1316 451
rect 1330 455 1336 456
rect 1330 451 1331 455
rect 1335 454 1336 455
rect 1339 455 1345 456
rect 1339 454 1340 455
rect 1335 452 1340 454
rect 1335 451 1336 452
rect 1330 450 1336 451
rect 1339 451 1340 452
rect 1344 451 1345 455
rect 1339 450 1345 451
rect 1375 455 1381 456
rect 1375 451 1376 455
rect 1380 454 1381 455
rect 1395 455 1401 456
rect 1395 454 1396 455
rect 1380 452 1396 454
rect 1380 451 1381 452
rect 1375 450 1381 451
rect 1395 451 1396 452
rect 1400 451 1401 455
rect 1395 450 1401 451
rect 1426 455 1432 456
rect 1426 451 1427 455
rect 1431 454 1432 455
rect 1459 455 1465 456
rect 1459 454 1460 455
rect 1431 452 1460 454
rect 1431 451 1432 452
rect 1426 450 1432 451
rect 1459 451 1460 452
rect 1464 451 1465 455
rect 1459 450 1465 451
rect 1490 455 1496 456
rect 1490 451 1491 455
rect 1495 454 1496 455
rect 1523 455 1529 456
rect 1523 454 1524 455
rect 1495 452 1524 454
rect 1495 451 1496 452
rect 1490 450 1496 451
rect 1523 451 1524 452
rect 1528 451 1529 455
rect 1523 450 1529 451
rect 1587 455 1593 456
rect 1587 451 1588 455
rect 1592 454 1593 455
rect 1634 455 1640 456
rect 1634 454 1635 455
rect 1592 452 1635 454
rect 1592 451 1593 452
rect 1587 450 1593 451
rect 1634 451 1635 452
rect 1639 451 1640 455
rect 1634 450 1640 451
rect 1659 455 1665 456
rect 1659 451 1660 455
rect 1664 454 1665 455
rect 1714 455 1720 456
rect 1714 454 1715 455
rect 1664 452 1715 454
rect 1664 451 1665 452
rect 1659 450 1665 451
rect 1714 451 1715 452
rect 1719 451 1720 455
rect 1714 450 1720 451
rect 1722 455 1728 456
rect 1722 451 1723 455
rect 1727 454 1728 455
rect 1731 455 1737 456
rect 1731 454 1732 455
rect 1727 452 1732 454
rect 1727 451 1728 452
rect 1722 450 1728 451
rect 1731 451 1732 452
rect 1736 451 1737 455
rect 1731 450 1737 451
rect 1762 455 1768 456
rect 1762 451 1763 455
rect 1767 454 1768 455
rect 1811 455 1817 456
rect 1811 454 1812 455
rect 1767 452 1812 454
rect 1767 451 1768 452
rect 1762 450 1768 451
rect 1811 451 1812 452
rect 1816 451 1817 455
rect 1811 450 1817 451
rect 1842 455 1848 456
rect 1842 451 1843 455
rect 1847 454 1848 455
rect 1891 455 1897 456
rect 1891 454 1892 455
rect 1847 452 1892 454
rect 1847 451 1848 452
rect 1842 450 1848 451
rect 1891 451 1892 452
rect 1896 451 1897 455
rect 1891 450 1897 451
rect 1922 455 1928 456
rect 1922 451 1923 455
rect 1927 454 1928 455
rect 1971 455 1977 456
rect 1971 454 1972 455
rect 1927 452 1972 454
rect 1927 451 1928 452
rect 1922 450 1928 451
rect 1971 451 1972 452
rect 1976 451 1977 455
rect 1971 450 1977 451
rect 2051 455 2057 456
rect 2051 451 2052 455
rect 2056 454 2057 455
rect 2062 455 2068 456
rect 2062 454 2063 455
rect 2056 452 2063 454
rect 2056 451 2057 452
rect 2051 450 2057 451
rect 2062 451 2063 452
rect 2067 451 2068 455
rect 2062 450 2068 451
rect 2082 455 2088 456
rect 2082 451 2083 455
rect 2087 454 2088 455
rect 2131 455 2137 456
rect 2131 454 2132 455
rect 2087 452 2132 454
rect 2087 451 2088 452
rect 2082 450 2088 451
rect 2131 451 2132 452
rect 2136 451 2137 455
rect 2131 450 2137 451
rect 2162 455 2168 456
rect 2162 451 2163 455
rect 2167 454 2168 455
rect 2211 455 2217 456
rect 2211 454 2212 455
rect 2167 452 2212 454
rect 2167 451 2168 452
rect 2162 450 2168 451
rect 2211 451 2212 452
rect 2216 451 2217 455
rect 2211 450 2217 451
rect 2291 455 2297 456
rect 2291 451 2292 455
rect 2296 454 2297 455
rect 2335 455 2341 456
rect 2335 454 2336 455
rect 2296 452 2336 454
rect 2296 451 2297 452
rect 2291 450 2297 451
rect 2335 451 2336 452
rect 2340 451 2341 455
rect 2335 450 2341 451
rect 2355 455 2361 456
rect 2355 451 2356 455
rect 2360 454 2361 455
rect 2366 455 2372 456
rect 2366 454 2367 455
rect 2360 452 2367 454
rect 2360 451 2361 452
rect 2355 450 2361 451
rect 2366 451 2367 452
rect 2371 451 2372 455
rect 2366 450 2372 451
rect 883 446 889 447
rect 1302 447 1308 448
rect 182 443 188 444
rect 182 439 183 443
rect 187 439 188 443
rect 182 438 188 439
rect 222 443 228 444
rect 222 439 223 443
rect 227 439 228 443
rect 222 438 228 439
rect 262 443 268 444
rect 262 439 263 443
rect 267 439 268 443
rect 262 438 268 439
rect 310 443 316 444
rect 310 439 311 443
rect 315 439 316 443
rect 310 438 316 439
rect 366 443 372 444
rect 366 439 367 443
rect 371 439 372 443
rect 366 438 372 439
rect 430 443 436 444
rect 430 439 431 443
rect 435 439 436 443
rect 430 438 436 439
rect 494 443 500 444
rect 494 439 495 443
rect 499 439 500 443
rect 494 438 500 439
rect 558 443 564 444
rect 558 439 559 443
rect 563 439 564 443
rect 558 438 564 439
rect 614 443 620 444
rect 614 439 615 443
rect 619 439 620 443
rect 614 438 620 439
rect 670 443 676 444
rect 670 439 671 443
rect 675 439 676 443
rect 670 438 676 439
rect 718 443 724 444
rect 718 439 719 443
rect 723 439 724 443
rect 718 438 724 439
rect 774 443 780 444
rect 774 439 775 443
rect 779 439 780 443
rect 774 438 780 439
rect 830 443 836 444
rect 830 439 831 443
rect 835 439 836 443
rect 830 438 836 439
rect 886 443 892 444
rect 886 439 887 443
rect 891 439 892 443
rect 1302 443 1303 447
rect 1307 443 1308 447
rect 1302 442 1308 443
rect 1342 447 1348 448
rect 1342 443 1343 447
rect 1347 443 1348 447
rect 1342 442 1348 443
rect 1398 447 1404 448
rect 1398 443 1399 447
rect 1403 443 1404 447
rect 1398 442 1404 443
rect 1462 447 1468 448
rect 1462 443 1463 447
rect 1467 443 1468 447
rect 1462 442 1468 443
rect 1526 447 1532 448
rect 1526 443 1527 447
rect 1531 443 1532 447
rect 1526 442 1532 443
rect 1590 447 1596 448
rect 1590 443 1591 447
rect 1595 443 1596 447
rect 1590 442 1596 443
rect 1662 447 1668 448
rect 1662 443 1663 447
rect 1667 443 1668 447
rect 1662 442 1668 443
rect 1734 447 1740 448
rect 1734 443 1735 447
rect 1739 443 1740 447
rect 1734 442 1740 443
rect 1814 447 1820 448
rect 1814 443 1815 447
rect 1819 443 1820 447
rect 1814 442 1820 443
rect 1894 447 1900 448
rect 1894 443 1895 447
rect 1899 443 1900 447
rect 1894 442 1900 443
rect 1974 447 1980 448
rect 1974 443 1975 447
rect 1979 443 1980 447
rect 1974 442 1980 443
rect 2054 447 2060 448
rect 2054 443 2055 447
rect 2059 443 2060 447
rect 2054 442 2060 443
rect 2134 447 2140 448
rect 2134 443 2135 447
rect 2139 443 2140 447
rect 2134 442 2140 443
rect 2214 447 2220 448
rect 2214 443 2215 447
rect 2219 443 2220 447
rect 2214 442 2220 443
rect 2294 447 2300 448
rect 2294 443 2295 447
rect 2299 443 2300 447
rect 2294 442 2300 443
rect 2358 447 2364 448
rect 2358 443 2359 447
rect 2363 443 2364 447
rect 2358 442 2364 443
rect 886 438 892 439
rect 1634 427 1640 428
rect 1278 424 1284 425
rect 690 423 696 424
rect 110 420 116 421
rect 110 416 111 420
rect 115 416 116 420
rect 690 419 691 423
rect 695 422 696 423
rect 695 420 870 422
rect 695 419 696 420
rect 690 418 696 419
rect 110 415 116 416
rect 167 415 173 416
rect 167 411 168 415
rect 172 414 173 415
rect 207 415 213 416
rect 207 414 208 415
rect 172 412 208 414
rect 172 411 173 412
rect 167 410 173 411
rect 207 411 208 412
rect 212 411 213 415
rect 207 410 213 411
rect 218 415 224 416
rect 218 411 219 415
rect 223 414 224 415
rect 247 415 253 416
rect 247 414 248 415
rect 223 412 248 414
rect 223 411 224 412
rect 218 410 224 411
rect 247 411 248 412
rect 252 411 253 415
rect 247 410 253 411
rect 258 415 264 416
rect 258 411 259 415
rect 263 414 264 415
rect 287 415 293 416
rect 287 414 288 415
rect 263 412 288 414
rect 263 411 264 412
rect 258 410 264 411
rect 287 411 288 412
rect 292 411 293 415
rect 287 410 293 411
rect 335 415 341 416
rect 335 411 336 415
rect 340 414 341 415
rect 350 415 356 416
rect 350 414 351 415
rect 340 412 351 414
rect 340 411 341 412
rect 335 410 341 411
rect 350 411 351 412
rect 355 411 356 415
rect 350 410 356 411
rect 391 415 400 416
rect 391 411 392 415
rect 399 411 400 415
rect 391 410 400 411
rect 455 415 464 416
rect 455 411 456 415
rect 463 411 464 415
rect 455 410 464 411
rect 466 415 472 416
rect 466 411 467 415
rect 471 414 472 415
rect 519 415 525 416
rect 519 414 520 415
rect 471 412 520 414
rect 471 411 472 412
rect 466 410 472 411
rect 519 411 520 412
rect 524 411 525 415
rect 519 410 525 411
rect 583 415 592 416
rect 583 411 584 415
rect 591 411 592 415
rect 583 410 592 411
rect 639 415 645 416
rect 639 411 640 415
rect 644 414 645 415
rect 647 415 653 416
rect 647 414 648 415
rect 644 412 648 414
rect 644 411 645 412
rect 639 410 645 411
rect 647 411 648 412
rect 652 411 653 415
rect 647 410 653 411
rect 695 415 704 416
rect 695 411 696 415
rect 703 411 704 415
rect 695 410 704 411
rect 743 415 749 416
rect 743 411 744 415
rect 748 414 749 415
rect 759 415 765 416
rect 759 414 760 415
rect 748 412 760 414
rect 748 411 749 412
rect 743 410 749 411
rect 759 411 760 412
rect 764 411 765 415
rect 759 410 765 411
rect 799 415 808 416
rect 799 411 800 415
rect 807 411 808 415
rect 799 410 808 411
rect 855 415 864 416
rect 855 411 856 415
rect 863 411 864 415
rect 868 414 870 420
rect 1238 420 1244 421
rect 1238 416 1239 420
rect 1243 416 1244 420
rect 1278 420 1279 424
rect 1283 420 1284 424
rect 1634 423 1635 427
rect 1639 426 1640 427
rect 2335 427 2341 428
rect 1639 424 1666 426
rect 1639 423 1640 424
rect 1634 422 1640 423
rect 1278 419 1284 420
rect 1327 419 1336 420
rect 911 415 917 416
rect 1238 415 1244 416
rect 1327 415 1328 419
rect 1335 415 1336 419
rect 911 414 912 415
rect 868 412 912 414
rect 855 410 864 411
rect 911 411 912 412
rect 916 411 917 415
rect 1327 414 1336 415
rect 1367 419 1373 420
rect 1367 415 1368 419
rect 1372 418 1373 419
rect 1375 419 1381 420
rect 1375 418 1376 419
rect 1372 416 1376 418
rect 1372 415 1373 416
rect 1367 414 1373 415
rect 1375 415 1376 416
rect 1380 415 1381 419
rect 1375 414 1381 415
rect 1423 419 1432 420
rect 1423 415 1424 419
rect 1431 415 1432 419
rect 1423 414 1432 415
rect 1487 419 1496 420
rect 1487 415 1488 419
rect 1495 415 1496 419
rect 1551 419 1557 420
rect 1551 418 1552 419
rect 1487 414 1496 415
rect 1500 416 1552 418
rect 911 410 917 411
rect 1454 411 1460 412
rect 1278 407 1284 408
rect 110 403 116 404
rect 110 399 111 403
rect 115 399 116 403
rect 110 398 116 399
rect 1238 403 1244 404
rect 1238 399 1239 403
rect 1243 399 1244 403
rect 1278 403 1279 407
rect 1283 403 1284 407
rect 1454 407 1455 411
rect 1459 410 1460 411
rect 1500 410 1502 416
rect 1551 415 1552 416
rect 1556 415 1557 419
rect 1551 414 1557 415
rect 1615 419 1621 420
rect 1615 415 1616 419
rect 1620 418 1621 419
rect 1654 419 1660 420
rect 1654 418 1655 419
rect 1620 416 1655 418
rect 1620 415 1621 416
rect 1615 414 1621 415
rect 1654 415 1655 416
rect 1659 415 1660 419
rect 1664 418 1666 424
rect 2335 423 2336 427
rect 2340 426 2341 427
rect 2340 424 2362 426
rect 2340 423 2341 424
rect 2335 422 2341 423
rect 1687 419 1693 420
rect 1687 418 1688 419
rect 1664 416 1688 418
rect 1654 414 1660 415
rect 1687 415 1688 416
rect 1692 415 1693 419
rect 1687 414 1693 415
rect 1759 419 1768 420
rect 1759 415 1760 419
rect 1767 415 1768 419
rect 1759 414 1768 415
rect 1839 419 1848 420
rect 1839 415 1840 419
rect 1847 415 1848 419
rect 1839 414 1848 415
rect 1919 419 1928 420
rect 1919 415 1920 419
rect 1927 415 1928 419
rect 1919 414 1928 415
rect 1930 419 1936 420
rect 1930 415 1931 419
rect 1935 418 1936 419
rect 1999 419 2005 420
rect 1999 418 2000 419
rect 1935 416 2000 418
rect 1935 415 1936 416
rect 1930 414 1936 415
rect 1999 415 2000 416
rect 2004 415 2005 419
rect 1999 414 2005 415
rect 2079 419 2088 420
rect 2079 415 2080 419
rect 2087 415 2088 419
rect 2079 414 2088 415
rect 2159 419 2168 420
rect 2159 415 2160 419
rect 2167 415 2168 419
rect 2159 414 2168 415
rect 2174 419 2180 420
rect 2174 415 2175 419
rect 2179 418 2180 419
rect 2239 419 2245 420
rect 2239 418 2240 419
rect 2179 416 2240 418
rect 2179 415 2180 416
rect 2174 414 2180 415
rect 2239 415 2240 416
rect 2244 415 2245 419
rect 2239 414 2245 415
rect 2319 419 2325 420
rect 2319 415 2320 419
rect 2324 418 2325 419
rect 2350 419 2356 420
rect 2350 418 2351 419
rect 2324 416 2351 418
rect 2324 415 2325 416
rect 2319 414 2325 415
rect 2350 415 2351 416
rect 2355 415 2356 419
rect 2360 418 2362 424
rect 2406 424 2412 425
rect 2406 420 2407 424
rect 2411 420 2412 424
rect 2383 419 2389 420
rect 2406 419 2412 420
rect 2383 418 2384 419
rect 2360 416 2384 418
rect 2350 414 2356 415
rect 2383 415 2384 416
rect 2388 415 2389 419
rect 2383 414 2389 415
rect 1459 408 1502 410
rect 1459 407 1460 408
rect 1454 406 1460 407
rect 2406 407 2412 408
rect 1278 402 1284 403
rect 2406 403 2407 407
rect 2411 403 2412 407
rect 2406 402 2412 403
rect 1238 398 1244 399
rect 1302 400 1308 401
rect 182 396 188 397
rect 182 392 183 396
rect 187 392 188 396
rect 182 391 188 392
rect 222 396 228 397
rect 222 392 223 396
rect 227 392 228 396
rect 222 391 228 392
rect 262 396 268 397
rect 262 392 263 396
rect 267 392 268 396
rect 262 391 268 392
rect 310 396 316 397
rect 310 392 311 396
rect 315 392 316 396
rect 310 391 316 392
rect 366 396 372 397
rect 366 392 367 396
rect 371 392 372 396
rect 366 391 372 392
rect 430 396 436 397
rect 430 392 431 396
rect 435 392 436 396
rect 430 391 436 392
rect 494 396 500 397
rect 494 392 495 396
rect 499 392 500 396
rect 494 391 500 392
rect 558 396 564 397
rect 558 392 559 396
rect 563 392 564 396
rect 558 391 564 392
rect 614 396 620 397
rect 614 392 615 396
rect 619 392 620 396
rect 614 391 620 392
rect 670 396 676 397
rect 670 392 671 396
rect 675 392 676 396
rect 670 391 676 392
rect 718 396 724 397
rect 718 392 719 396
rect 723 392 724 396
rect 718 391 724 392
rect 774 396 780 397
rect 774 392 775 396
rect 779 392 780 396
rect 774 391 780 392
rect 830 396 836 397
rect 830 392 831 396
rect 835 392 836 396
rect 830 391 836 392
rect 886 396 892 397
rect 886 392 887 396
rect 891 392 892 396
rect 1302 396 1303 400
rect 1307 396 1308 400
rect 1302 395 1308 396
rect 1342 400 1348 401
rect 1342 396 1343 400
rect 1347 396 1348 400
rect 1342 395 1348 396
rect 1398 400 1404 401
rect 1398 396 1399 400
rect 1403 396 1404 400
rect 1398 395 1404 396
rect 1462 400 1468 401
rect 1462 396 1463 400
rect 1467 396 1468 400
rect 1462 395 1468 396
rect 1526 400 1532 401
rect 1526 396 1527 400
rect 1531 396 1532 400
rect 1526 395 1532 396
rect 1590 400 1596 401
rect 1590 396 1591 400
rect 1595 396 1596 400
rect 1590 395 1596 396
rect 1662 400 1668 401
rect 1662 396 1663 400
rect 1667 396 1668 400
rect 1662 395 1668 396
rect 1734 400 1740 401
rect 1734 396 1735 400
rect 1739 396 1740 400
rect 1734 395 1740 396
rect 1814 400 1820 401
rect 1814 396 1815 400
rect 1819 396 1820 400
rect 1814 395 1820 396
rect 1894 400 1900 401
rect 1894 396 1895 400
rect 1899 396 1900 400
rect 1894 395 1900 396
rect 1974 400 1980 401
rect 1974 396 1975 400
rect 1979 396 1980 400
rect 1974 395 1980 396
rect 2054 400 2060 401
rect 2054 396 2055 400
rect 2059 396 2060 400
rect 2054 395 2060 396
rect 2134 400 2140 401
rect 2134 396 2135 400
rect 2139 396 2140 400
rect 2134 395 2140 396
rect 2214 400 2220 401
rect 2214 396 2215 400
rect 2219 396 2220 400
rect 2214 395 2220 396
rect 2294 400 2300 401
rect 2294 396 2295 400
rect 2299 396 2300 400
rect 2294 395 2300 396
rect 2358 400 2364 401
rect 2358 396 2359 400
rect 2363 396 2364 400
rect 2358 395 2364 396
rect 886 391 892 392
rect 134 384 140 385
rect 134 380 135 384
rect 139 380 140 384
rect 134 379 140 380
rect 174 384 180 385
rect 174 380 175 384
rect 179 380 180 384
rect 174 379 180 380
rect 230 384 236 385
rect 230 380 231 384
rect 235 380 236 384
rect 230 379 236 380
rect 286 384 292 385
rect 286 380 287 384
rect 291 380 292 384
rect 286 379 292 380
rect 342 384 348 385
rect 342 380 343 384
rect 347 380 348 384
rect 342 379 348 380
rect 390 384 396 385
rect 390 380 391 384
rect 395 380 396 384
rect 390 379 396 380
rect 438 384 444 385
rect 438 380 439 384
rect 443 380 444 384
rect 438 379 444 380
rect 486 384 492 385
rect 486 380 487 384
rect 491 380 492 384
rect 486 379 492 380
rect 534 384 540 385
rect 534 380 535 384
rect 539 380 540 384
rect 534 379 540 380
rect 582 384 588 385
rect 582 380 583 384
rect 587 380 588 384
rect 582 379 588 380
rect 630 384 636 385
rect 630 380 631 384
rect 635 380 636 384
rect 630 379 636 380
rect 678 384 684 385
rect 678 380 679 384
rect 683 380 684 384
rect 678 379 684 380
rect 726 384 732 385
rect 726 380 727 384
rect 731 380 732 384
rect 726 379 732 380
rect 774 384 780 385
rect 774 380 775 384
rect 779 380 780 384
rect 774 379 780 380
rect 1446 384 1452 385
rect 1446 380 1447 384
rect 1451 380 1452 384
rect 1446 379 1452 380
rect 1486 384 1492 385
rect 1486 380 1487 384
rect 1491 380 1492 384
rect 1486 379 1492 380
rect 1534 384 1540 385
rect 1534 380 1535 384
rect 1539 380 1540 384
rect 1534 379 1540 380
rect 1590 384 1596 385
rect 1590 380 1591 384
rect 1595 380 1596 384
rect 1590 379 1596 380
rect 1662 384 1668 385
rect 1662 380 1663 384
rect 1667 380 1668 384
rect 1662 379 1668 380
rect 1734 384 1740 385
rect 1734 380 1735 384
rect 1739 380 1740 384
rect 1734 379 1740 380
rect 1814 384 1820 385
rect 1814 380 1815 384
rect 1819 380 1820 384
rect 1814 379 1820 380
rect 1894 384 1900 385
rect 1894 380 1895 384
rect 1899 380 1900 384
rect 1894 379 1900 380
rect 1966 384 1972 385
rect 1966 380 1967 384
rect 1971 380 1972 384
rect 1966 379 1972 380
rect 2038 384 2044 385
rect 2038 380 2039 384
rect 2043 380 2044 384
rect 2038 379 2044 380
rect 2110 384 2116 385
rect 2110 380 2111 384
rect 2115 380 2116 384
rect 2110 379 2116 380
rect 2174 384 2180 385
rect 2174 380 2175 384
rect 2179 380 2180 384
rect 2174 379 2180 380
rect 2238 384 2244 385
rect 2238 380 2239 384
rect 2243 380 2244 384
rect 2238 379 2244 380
rect 2302 384 2308 385
rect 2302 380 2303 384
rect 2307 380 2308 384
rect 2302 379 2308 380
rect 2358 384 2364 385
rect 2358 380 2359 384
rect 2363 380 2364 384
rect 2358 379 2364 380
rect 110 377 116 378
rect 110 373 111 377
rect 115 373 116 377
rect 1238 377 1244 378
rect 110 372 116 373
rect 566 375 572 376
rect 566 371 567 375
rect 571 374 572 375
rect 571 372 778 374
rect 1238 373 1239 377
rect 1243 373 1244 377
rect 1238 372 1244 373
rect 1278 377 1284 378
rect 1278 373 1279 377
rect 1283 373 1284 377
rect 1278 372 1284 373
rect 2406 377 2412 378
rect 2406 373 2407 377
rect 2411 373 2412 377
rect 2406 372 2412 373
rect 571 371 572 372
rect 566 370 572 371
rect 159 363 168 364
rect 110 360 116 361
rect 110 356 111 360
rect 115 356 116 360
rect 159 359 160 363
rect 167 359 168 363
rect 159 358 168 359
rect 199 363 205 364
rect 199 359 200 363
rect 204 362 205 363
rect 222 363 228 364
rect 222 362 223 363
rect 204 360 223 362
rect 204 359 205 360
rect 199 358 205 359
rect 222 359 223 360
rect 227 359 228 363
rect 222 358 228 359
rect 255 363 261 364
rect 255 359 256 363
rect 260 362 261 363
rect 278 363 284 364
rect 278 362 279 363
rect 260 360 279 362
rect 260 359 261 360
rect 255 358 261 359
rect 278 359 279 360
rect 283 359 284 363
rect 278 358 284 359
rect 298 363 304 364
rect 298 359 299 363
rect 303 362 304 363
rect 311 363 317 364
rect 311 362 312 363
rect 303 360 312 362
rect 303 359 304 360
rect 298 358 304 359
rect 311 359 312 360
rect 316 359 317 363
rect 311 358 317 359
rect 334 363 340 364
rect 334 359 335 363
rect 339 362 340 363
rect 367 363 373 364
rect 367 362 368 363
rect 339 360 368 362
rect 339 359 340 360
rect 334 358 340 359
rect 367 359 368 360
rect 372 359 373 363
rect 367 358 373 359
rect 375 363 381 364
rect 375 359 376 363
rect 380 362 381 363
rect 415 363 421 364
rect 415 362 416 363
rect 380 360 416 362
rect 380 359 381 360
rect 375 358 381 359
rect 415 359 416 360
rect 420 359 421 363
rect 415 358 421 359
rect 423 363 429 364
rect 423 359 424 363
rect 428 362 429 363
rect 463 363 469 364
rect 463 362 464 363
rect 428 360 464 362
rect 428 359 429 360
rect 423 358 429 359
rect 463 359 464 360
rect 468 359 469 363
rect 463 358 469 359
rect 511 363 517 364
rect 511 359 512 363
rect 516 362 517 363
rect 526 363 532 364
rect 526 362 527 363
rect 516 360 527 362
rect 516 359 517 360
rect 511 358 517 359
rect 526 359 527 360
rect 531 359 532 363
rect 526 358 532 359
rect 559 363 565 364
rect 559 359 560 363
rect 564 362 565 363
rect 574 363 580 364
rect 574 362 575 363
rect 564 360 575 362
rect 564 359 565 360
rect 559 358 565 359
rect 574 359 575 360
rect 579 359 580 363
rect 574 358 580 359
rect 607 363 613 364
rect 607 359 608 363
rect 612 362 613 363
rect 622 363 628 364
rect 622 362 623 363
rect 612 360 623 362
rect 612 359 613 360
rect 607 358 613 359
rect 622 359 623 360
rect 627 359 628 363
rect 622 358 628 359
rect 655 363 661 364
rect 655 359 656 363
rect 660 362 661 363
rect 670 363 676 364
rect 670 362 671 363
rect 660 360 671 362
rect 660 359 661 360
rect 655 358 661 359
rect 670 359 671 360
rect 675 359 676 363
rect 670 358 676 359
rect 703 363 709 364
rect 703 359 704 363
rect 708 362 709 363
rect 718 363 724 364
rect 718 362 719 363
rect 708 360 719 362
rect 708 359 709 360
rect 703 358 709 359
rect 718 359 719 360
rect 723 359 724 363
rect 718 358 724 359
rect 751 363 757 364
rect 751 359 752 363
rect 756 362 757 363
rect 766 363 772 364
rect 766 362 767 363
rect 756 360 767 362
rect 756 359 757 360
rect 751 358 757 359
rect 766 359 767 360
rect 771 359 772 363
rect 776 362 778 372
rect 1714 371 1720 372
rect 1714 367 1715 371
rect 1719 370 1720 371
rect 1719 368 1850 370
rect 1719 367 1720 368
rect 1714 366 1720 367
rect 799 363 805 364
rect 799 362 800 363
rect 776 360 800 362
rect 766 358 772 359
rect 799 359 800 360
rect 804 359 805 363
rect 1471 363 1480 364
rect 799 358 805 359
rect 1238 360 1244 361
rect 110 355 116 356
rect 1238 356 1239 360
rect 1243 356 1244 360
rect 1238 355 1244 356
rect 1278 360 1284 361
rect 1278 356 1279 360
rect 1283 356 1284 360
rect 1471 359 1472 363
rect 1479 359 1480 363
rect 1471 358 1480 359
rect 1511 363 1517 364
rect 1511 359 1512 363
rect 1516 362 1517 363
rect 1526 363 1532 364
rect 1526 362 1527 363
rect 1516 360 1527 362
rect 1516 359 1517 360
rect 1511 358 1517 359
rect 1526 359 1527 360
rect 1531 359 1532 363
rect 1526 358 1532 359
rect 1559 363 1565 364
rect 1559 359 1560 363
rect 1564 362 1565 363
rect 1582 363 1588 364
rect 1582 362 1583 363
rect 1564 360 1583 362
rect 1564 359 1565 360
rect 1559 358 1565 359
rect 1582 359 1583 360
rect 1587 359 1588 363
rect 1582 358 1588 359
rect 1598 363 1604 364
rect 1598 359 1599 363
rect 1603 362 1604 363
rect 1615 363 1621 364
rect 1615 362 1616 363
rect 1603 360 1616 362
rect 1603 359 1604 360
rect 1598 358 1604 359
rect 1615 359 1616 360
rect 1620 359 1621 363
rect 1615 358 1621 359
rect 1687 363 1693 364
rect 1687 359 1688 363
rect 1692 362 1693 363
rect 1726 363 1732 364
rect 1726 362 1727 363
rect 1692 360 1727 362
rect 1692 359 1693 360
rect 1687 358 1693 359
rect 1726 359 1727 360
rect 1731 359 1732 363
rect 1726 358 1732 359
rect 1759 363 1765 364
rect 1759 359 1760 363
rect 1764 362 1765 363
rect 1806 363 1812 364
rect 1806 362 1807 363
rect 1764 360 1807 362
rect 1764 359 1765 360
rect 1759 358 1765 359
rect 1806 359 1807 360
rect 1811 359 1812 363
rect 1806 358 1812 359
rect 1822 363 1828 364
rect 1822 359 1823 363
rect 1827 362 1828 363
rect 1839 363 1845 364
rect 1839 362 1840 363
rect 1827 360 1840 362
rect 1827 359 1828 360
rect 1822 358 1828 359
rect 1839 359 1840 360
rect 1844 359 1845 363
rect 1848 362 1850 368
rect 1919 363 1925 364
rect 1919 362 1920 363
rect 1848 360 1920 362
rect 1839 358 1845 359
rect 1919 359 1920 360
rect 1924 359 1925 363
rect 1919 358 1925 359
rect 1991 363 1997 364
rect 1991 359 1992 363
rect 1996 362 1997 363
rect 2030 363 2036 364
rect 2030 362 2031 363
rect 1996 360 2031 362
rect 1996 359 1997 360
rect 1991 358 1997 359
rect 2030 359 2031 360
rect 2035 359 2036 363
rect 2030 358 2036 359
rect 2062 363 2069 364
rect 2062 359 2063 363
rect 2068 359 2069 363
rect 2135 363 2141 364
rect 2135 362 2136 363
rect 2062 358 2069 359
rect 2072 360 2136 362
rect 1278 355 1284 356
rect 1974 355 1980 356
rect 1974 351 1975 355
rect 1979 354 1980 355
rect 2072 354 2074 360
rect 2135 359 2136 360
rect 2140 359 2141 363
rect 2135 358 2141 359
rect 2143 363 2149 364
rect 2143 359 2144 363
rect 2148 362 2149 363
rect 2199 363 2205 364
rect 2199 362 2200 363
rect 2148 360 2200 362
rect 2148 359 2149 360
rect 2143 358 2149 359
rect 2199 359 2200 360
rect 2204 359 2205 363
rect 2199 358 2205 359
rect 2207 363 2213 364
rect 2207 359 2208 363
rect 2212 362 2213 363
rect 2263 363 2269 364
rect 2263 362 2264 363
rect 2212 360 2264 362
rect 2212 359 2213 360
rect 2207 358 2213 359
rect 2263 359 2264 360
rect 2268 359 2269 363
rect 2263 358 2269 359
rect 2271 363 2277 364
rect 2271 359 2272 363
rect 2276 362 2277 363
rect 2327 363 2333 364
rect 2327 362 2328 363
rect 2276 360 2328 362
rect 2276 359 2277 360
rect 2271 358 2277 359
rect 2327 359 2328 360
rect 2332 359 2333 363
rect 2327 358 2333 359
rect 2338 363 2344 364
rect 2338 359 2339 363
rect 2343 362 2344 363
rect 2383 363 2389 364
rect 2383 362 2384 363
rect 2343 360 2384 362
rect 2343 359 2344 360
rect 2338 358 2344 359
rect 2383 359 2384 360
rect 2388 359 2389 363
rect 2383 358 2389 359
rect 2406 360 2412 361
rect 2406 356 2407 360
rect 2411 356 2412 360
rect 2406 355 2412 356
rect 1979 352 2074 354
rect 1979 351 1980 352
rect 1974 350 1980 351
rect 134 337 140 338
rect 134 333 135 337
rect 139 333 140 337
rect 134 332 140 333
rect 174 337 180 338
rect 174 333 175 337
rect 179 333 180 337
rect 174 332 180 333
rect 230 337 236 338
rect 230 333 231 337
rect 235 333 236 337
rect 230 332 236 333
rect 286 337 292 338
rect 286 333 287 337
rect 291 333 292 337
rect 286 332 292 333
rect 342 337 348 338
rect 342 333 343 337
rect 347 333 348 337
rect 342 332 348 333
rect 390 337 396 338
rect 390 333 391 337
rect 395 333 396 337
rect 390 332 396 333
rect 438 337 444 338
rect 438 333 439 337
rect 443 333 444 337
rect 438 332 444 333
rect 486 337 492 338
rect 486 333 487 337
rect 491 333 492 337
rect 486 332 492 333
rect 534 337 540 338
rect 534 333 535 337
rect 539 333 540 337
rect 534 332 540 333
rect 582 337 588 338
rect 582 333 583 337
rect 587 333 588 337
rect 582 332 588 333
rect 630 337 636 338
rect 630 333 631 337
rect 635 333 636 337
rect 630 332 636 333
rect 678 337 684 338
rect 678 333 679 337
rect 683 333 684 337
rect 678 332 684 333
rect 726 337 732 338
rect 726 333 727 337
rect 731 333 732 337
rect 726 332 732 333
rect 774 337 780 338
rect 774 333 775 337
rect 779 333 780 337
rect 774 332 780 333
rect 1446 337 1452 338
rect 1446 333 1447 337
rect 1451 333 1452 337
rect 1446 332 1452 333
rect 1486 337 1492 338
rect 1486 333 1487 337
rect 1491 333 1492 337
rect 1486 332 1492 333
rect 1534 337 1540 338
rect 1534 333 1535 337
rect 1539 333 1540 337
rect 1534 332 1540 333
rect 1590 337 1596 338
rect 1590 333 1591 337
rect 1595 333 1596 337
rect 1590 332 1596 333
rect 1662 337 1668 338
rect 1662 333 1663 337
rect 1667 333 1668 337
rect 1662 332 1668 333
rect 1734 337 1740 338
rect 1734 333 1735 337
rect 1739 333 1740 337
rect 1734 332 1740 333
rect 1814 337 1820 338
rect 1814 333 1815 337
rect 1819 333 1820 337
rect 1814 332 1820 333
rect 1894 337 1900 338
rect 1894 333 1895 337
rect 1899 333 1900 337
rect 1894 332 1900 333
rect 1966 337 1972 338
rect 1966 333 1967 337
rect 1971 333 1972 337
rect 1966 332 1972 333
rect 2038 337 2044 338
rect 2038 333 2039 337
rect 2043 333 2044 337
rect 2038 332 2044 333
rect 2110 337 2116 338
rect 2110 333 2111 337
rect 2115 333 2116 337
rect 2110 332 2116 333
rect 2174 337 2180 338
rect 2174 333 2175 337
rect 2179 333 2180 337
rect 2174 332 2180 333
rect 2238 337 2244 338
rect 2238 333 2239 337
rect 2243 333 2244 337
rect 2238 332 2244 333
rect 2302 337 2308 338
rect 2302 333 2303 337
rect 2307 333 2308 337
rect 2302 332 2308 333
rect 2358 337 2364 338
rect 2358 333 2359 337
rect 2363 333 2364 337
rect 2358 332 2364 333
rect 131 327 137 328
rect 131 323 132 327
rect 136 323 137 327
rect 131 322 137 323
rect 162 327 168 328
rect 162 323 163 327
rect 167 326 168 327
rect 171 327 177 328
rect 171 326 172 327
rect 167 324 172 326
rect 167 323 168 324
rect 162 322 168 323
rect 171 323 172 324
rect 176 323 177 327
rect 171 322 177 323
rect 222 327 233 328
rect 222 323 223 327
rect 227 323 228 327
rect 232 323 233 327
rect 222 322 233 323
rect 278 327 289 328
rect 278 323 279 327
rect 283 323 284 327
rect 288 323 289 327
rect 278 322 289 323
rect 339 327 345 328
rect 339 323 340 327
rect 344 326 345 327
rect 375 327 381 328
rect 375 326 376 327
rect 344 324 376 326
rect 344 323 345 324
rect 339 322 345 323
rect 375 323 376 324
rect 380 323 381 327
rect 375 322 381 323
rect 387 327 393 328
rect 387 323 388 327
rect 392 326 393 327
rect 423 327 429 328
rect 423 326 424 327
rect 392 324 424 326
rect 392 323 393 324
rect 387 322 393 323
rect 423 323 424 324
rect 428 323 429 327
rect 423 322 429 323
rect 435 327 441 328
rect 435 323 436 327
rect 440 326 441 327
rect 466 327 472 328
rect 466 326 467 327
rect 440 324 467 326
rect 440 323 441 324
rect 435 322 441 323
rect 466 323 467 324
rect 471 323 472 327
rect 466 322 472 323
rect 483 327 489 328
rect 483 323 484 327
rect 488 326 489 327
rect 526 327 537 328
rect 488 324 522 326
rect 488 323 489 324
rect 483 322 489 323
rect 133 318 135 322
rect 278 319 284 320
rect 278 318 279 319
rect 133 316 279 318
rect 278 315 279 316
rect 283 315 284 319
rect 520 318 522 324
rect 526 323 527 327
rect 531 323 532 327
rect 536 323 537 327
rect 526 322 537 323
rect 574 327 585 328
rect 574 323 575 327
rect 579 323 580 327
rect 584 323 585 327
rect 574 322 585 323
rect 622 327 633 328
rect 622 323 623 327
rect 627 323 628 327
rect 632 323 633 327
rect 622 322 633 323
rect 670 327 681 328
rect 670 323 671 327
rect 675 323 676 327
rect 680 323 681 327
rect 670 322 681 323
rect 718 327 729 328
rect 718 323 719 327
rect 723 323 724 327
rect 728 323 729 327
rect 718 322 729 323
rect 766 327 777 328
rect 766 323 767 327
rect 771 323 772 327
rect 776 323 777 327
rect 766 322 777 323
rect 1443 327 1449 328
rect 1443 323 1444 327
rect 1448 326 1449 327
rect 1454 327 1460 328
rect 1454 326 1455 327
rect 1448 324 1455 326
rect 1448 323 1449 324
rect 1443 322 1449 323
rect 1454 323 1455 324
rect 1459 323 1460 327
rect 1454 322 1460 323
rect 1474 327 1480 328
rect 1474 323 1475 327
rect 1479 326 1480 327
rect 1483 327 1489 328
rect 1483 326 1484 327
rect 1479 324 1484 326
rect 1479 323 1480 324
rect 1474 322 1480 323
rect 1483 323 1484 324
rect 1488 323 1489 327
rect 1483 322 1489 323
rect 1526 327 1537 328
rect 1526 323 1527 327
rect 1531 323 1532 327
rect 1536 323 1537 327
rect 1526 322 1537 323
rect 1582 327 1593 328
rect 1582 323 1583 327
rect 1587 323 1588 327
rect 1592 323 1593 327
rect 1582 322 1593 323
rect 1654 327 1665 328
rect 1654 323 1655 327
rect 1659 323 1660 327
rect 1664 323 1665 327
rect 1654 322 1665 323
rect 1726 327 1737 328
rect 1726 323 1727 327
rect 1731 323 1732 327
rect 1736 323 1737 327
rect 1726 322 1737 323
rect 1806 327 1817 328
rect 1806 323 1807 327
rect 1811 323 1812 327
rect 1816 323 1817 327
rect 1806 322 1817 323
rect 1891 327 1897 328
rect 1891 323 1892 327
rect 1896 326 1897 327
rect 1930 327 1936 328
rect 1930 326 1931 327
rect 1896 324 1931 326
rect 1896 323 1897 324
rect 1891 322 1897 323
rect 1930 323 1931 324
rect 1935 323 1936 327
rect 1930 322 1936 323
rect 1963 327 1969 328
rect 1963 323 1964 327
rect 1968 326 1969 327
rect 1974 327 1980 328
rect 1974 326 1975 327
rect 1968 324 1975 326
rect 1968 323 1969 324
rect 1963 322 1969 323
rect 1974 323 1975 324
rect 1979 323 1980 327
rect 1974 322 1980 323
rect 2030 327 2041 328
rect 2030 323 2031 327
rect 2035 323 2036 327
rect 2040 323 2041 327
rect 2030 322 2041 323
rect 2107 327 2113 328
rect 2107 323 2108 327
rect 2112 326 2113 327
rect 2143 327 2149 328
rect 2143 326 2144 327
rect 2112 324 2144 326
rect 2112 323 2113 324
rect 2107 322 2113 323
rect 2143 323 2144 324
rect 2148 323 2149 327
rect 2143 322 2149 323
rect 2171 327 2177 328
rect 2171 323 2172 327
rect 2176 326 2177 327
rect 2207 327 2213 328
rect 2207 326 2208 327
rect 2176 324 2208 326
rect 2176 323 2177 324
rect 2171 322 2177 323
rect 2207 323 2208 324
rect 2212 323 2213 327
rect 2207 322 2213 323
rect 2235 327 2241 328
rect 2235 323 2236 327
rect 2240 326 2241 327
rect 2271 327 2277 328
rect 2271 326 2272 327
rect 2240 324 2272 326
rect 2240 323 2241 324
rect 2235 322 2241 323
rect 2271 323 2272 324
rect 2276 323 2277 327
rect 2271 322 2277 323
rect 2282 327 2288 328
rect 2282 323 2283 327
rect 2287 326 2288 327
rect 2299 327 2305 328
rect 2299 326 2300 327
rect 2287 324 2300 326
rect 2287 323 2288 324
rect 2282 322 2288 323
rect 2299 323 2300 324
rect 2304 323 2305 327
rect 2299 322 2305 323
rect 2350 327 2361 328
rect 2350 323 2351 327
rect 2355 323 2356 327
rect 2360 323 2361 327
rect 2350 322 2361 323
rect 610 319 616 320
rect 610 318 611 319
rect 520 316 611 318
rect 278 314 284 315
rect 610 315 611 316
rect 615 315 616 319
rect 1598 319 1604 320
rect 1598 318 1599 319
rect 610 314 616 315
rect 1492 316 1599 318
rect 1492 314 1494 316
rect 1598 315 1599 316
rect 1603 315 1604 319
rect 1822 319 1828 320
rect 1822 318 1823 319
rect 1598 314 1604 315
rect 1796 316 1823 318
rect 1796 314 1798 316
rect 1822 315 1823 316
rect 1827 315 1828 319
rect 1822 314 1828 315
rect 1491 313 1497 314
rect 131 311 137 312
rect 131 307 132 311
rect 136 310 137 311
rect 154 311 160 312
rect 154 310 155 311
rect 136 308 155 310
rect 136 307 137 308
rect 131 306 137 307
rect 154 307 155 308
rect 159 307 160 311
rect 154 306 160 307
rect 162 311 168 312
rect 162 307 163 311
rect 167 310 168 311
rect 179 311 185 312
rect 179 310 180 311
rect 167 308 180 310
rect 167 307 168 308
rect 162 306 168 307
rect 179 307 180 308
rect 184 307 185 311
rect 179 306 185 307
rect 210 311 216 312
rect 210 307 211 311
rect 215 310 216 311
rect 251 311 257 312
rect 251 310 252 311
rect 215 308 252 310
rect 215 307 216 308
rect 210 306 216 307
rect 251 307 252 308
rect 256 307 257 311
rect 251 306 257 307
rect 323 311 329 312
rect 323 307 324 311
rect 328 310 329 311
rect 334 311 340 312
rect 334 310 335 311
rect 328 308 335 310
rect 328 307 329 308
rect 323 306 329 307
rect 334 307 335 308
rect 339 307 340 311
rect 334 306 340 307
rect 354 311 360 312
rect 354 307 355 311
rect 359 310 360 311
rect 387 311 393 312
rect 387 310 388 311
rect 359 308 388 310
rect 359 307 360 308
rect 354 306 360 307
rect 387 307 388 308
rect 392 307 393 311
rect 387 306 393 307
rect 418 311 424 312
rect 418 307 419 311
rect 423 310 424 311
rect 443 311 449 312
rect 443 310 444 311
rect 423 308 444 310
rect 423 307 424 308
rect 418 306 424 307
rect 443 307 444 308
rect 448 307 449 311
rect 443 306 449 307
rect 474 311 480 312
rect 474 307 475 311
rect 479 310 480 311
rect 499 311 505 312
rect 499 310 500 311
rect 479 308 500 310
rect 479 307 480 308
rect 474 306 480 307
rect 499 307 500 308
rect 504 307 505 311
rect 499 306 505 307
rect 535 311 541 312
rect 535 307 536 311
rect 540 310 541 311
rect 547 311 553 312
rect 547 310 548 311
rect 540 308 548 310
rect 540 307 541 308
rect 535 306 541 307
rect 547 307 548 308
rect 552 307 553 311
rect 547 306 553 307
rect 587 311 593 312
rect 587 307 588 311
rect 592 310 593 311
rect 618 311 624 312
rect 618 310 619 311
rect 592 308 619 310
rect 592 307 593 308
rect 587 306 593 307
rect 618 307 619 308
rect 623 307 624 311
rect 618 306 624 307
rect 627 311 633 312
rect 627 307 628 311
rect 632 310 633 311
rect 666 311 672 312
rect 666 310 667 311
rect 632 308 667 310
rect 632 307 633 308
rect 627 306 633 307
rect 666 307 667 308
rect 671 307 672 311
rect 666 306 672 307
rect 675 311 681 312
rect 675 307 676 311
rect 680 310 681 311
rect 714 311 720 312
rect 714 310 715 311
rect 680 308 715 310
rect 680 307 681 308
rect 675 306 681 307
rect 714 307 715 308
rect 719 307 720 311
rect 714 306 720 307
rect 723 311 729 312
rect 723 307 724 311
rect 728 310 729 311
rect 762 311 768 312
rect 762 310 763 311
rect 728 308 763 310
rect 728 307 729 308
rect 723 306 729 307
rect 762 307 763 308
rect 767 307 768 311
rect 762 306 768 307
rect 771 311 777 312
rect 771 307 772 311
rect 776 310 777 311
rect 806 311 812 312
rect 806 310 807 311
rect 776 308 807 310
rect 776 307 777 308
rect 771 306 777 307
rect 806 307 807 308
rect 811 307 812 311
rect 806 306 812 307
rect 814 311 825 312
rect 814 307 815 311
rect 819 307 820 311
rect 824 307 825 311
rect 814 306 825 307
rect 858 311 864 312
rect 858 307 859 311
rect 863 310 864 311
rect 867 311 873 312
rect 867 310 868 311
rect 863 308 868 310
rect 863 307 864 308
rect 858 306 864 307
rect 867 307 868 308
rect 872 307 873 311
rect 867 306 873 307
rect 906 311 912 312
rect 906 307 907 311
rect 911 310 912 311
rect 915 311 921 312
rect 915 310 916 311
rect 911 308 916 310
rect 911 307 912 308
rect 906 306 912 307
rect 915 307 916 308
rect 920 307 921 311
rect 1491 309 1492 313
rect 1496 309 1497 313
rect 1795 313 1801 314
rect 1491 308 1497 309
rect 1522 311 1528 312
rect 915 306 921 307
rect 1522 307 1523 311
rect 1527 310 1528 311
rect 1531 311 1537 312
rect 1531 310 1532 311
rect 1527 308 1532 310
rect 1527 307 1528 308
rect 1522 306 1528 307
rect 1531 307 1532 308
rect 1536 307 1537 311
rect 1531 306 1537 307
rect 1562 311 1568 312
rect 1562 307 1563 311
rect 1567 310 1568 311
rect 1571 311 1577 312
rect 1571 310 1572 311
rect 1567 308 1572 310
rect 1567 307 1568 308
rect 1562 306 1568 307
rect 1571 307 1572 308
rect 1576 307 1577 311
rect 1571 306 1577 307
rect 1602 311 1608 312
rect 1602 307 1603 311
rect 1607 310 1608 311
rect 1611 311 1617 312
rect 1611 310 1612 311
rect 1607 308 1612 310
rect 1607 307 1608 308
rect 1602 306 1608 307
rect 1611 307 1612 308
rect 1616 307 1617 311
rect 1611 306 1617 307
rect 1642 311 1648 312
rect 1642 307 1643 311
rect 1647 310 1648 311
rect 1651 311 1657 312
rect 1651 310 1652 311
rect 1647 308 1652 310
rect 1647 307 1648 308
rect 1642 306 1648 307
rect 1651 307 1652 308
rect 1656 307 1657 311
rect 1651 306 1657 307
rect 1682 311 1688 312
rect 1682 307 1683 311
rect 1687 310 1688 311
rect 1691 311 1697 312
rect 1691 310 1692 311
rect 1687 308 1692 310
rect 1687 307 1688 308
rect 1682 306 1688 307
rect 1691 307 1692 308
rect 1696 307 1697 311
rect 1691 306 1697 307
rect 1722 311 1728 312
rect 1722 307 1723 311
rect 1727 310 1728 311
rect 1739 311 1745 312
rect 1739 310 1740 311
rect 1727 308 1740 310
rect 1727 307 1728 308
rect 1722 306 1728 307
rect 1739 307 1740 308
rect 1744 307 1745 311
rect 1795 309 1796 313
rect 1800 309 1801 313
rect 1795 308 1801 309
rect 1826 311 1832 312
rect 1739 306 1745 307
rect 1826 307 1827 311
rect 1831 310 1832 311
rect 1859 311 1865 312
rect 1859 310 1860 311
rect 1831 308 1860 310
rect 1831 307 1832 308
rect 1826 306 1832 307
rect 1859 307 1860 308
rect 1864 307 1865 311
rect 1859 306 1865 307
rect 1895 311 1901 312
rect 1895 307 1896 311
rect 1900 310 1901 311
rect 1931 311 1937 312
rect 1931 310 1932 311
rect 1900 308 1932 310
rect 1900 307 1901 308
rect 1895 306 1901 307
rect 1931 307 1932 308
rect 1936 307 1937 311
rect 1931 306 1937 307
rect 1974 311 1980 312
rect 1974 307 1975 311
rect 1979 310 1980 311
rect 2003 311 2009 312
rect 2003 310 2004 311
rect 1979 308 2004 310
rect 1979 307 1980 308
rect 1974 306 1980 307
rect 2003 307 2004 308
rect 2008 307 2009 311
rect 2003 306 2009 307
rect 2067 311 2073 312
rect 2067 307 2068 311
rect 2072 310 2073 311
rect 2090 311 2096 312
rect 2090 310 2091 311
rect 2072 308 2091 310
rect 2072 307 2073 308
rect 2067 306 2073 307
rect 2090 307 2091 308
rect 2095 307 2096 311
rect 2090 306 2096 307
rect 2098 311 2104 312
rect 2098 307 2099 311
rect 2103 310 2104 311
rect 2131 311 2137 312
rect 2131 310 2132 311
rect 2103 308 2132 310
rect 2103 307 2104 308
rect 2098 306 2104 307
rect 2131 307 2132 308
rect 2136 307 2137 311
rect 2131 306 2137 307
rect 2162 311 2168 312
rect 2162 307 2163 311
rect 2167 310 2168 311
rect 2187 311 2193 312
rect 2187 310 2188 311
rect 2167 308 2188 310
rect 2167 307 2168 308
rect 2162 306 2168 307
rect 2187 307 2188 308
rect 2192 307 2193 311
rect 2187 306 2193 307
rect 2218 311 2224 312
rect 2218 307 2219 311
rect 2223 310 2224 311
rect 2251 311 2257 312
rect 2251 310 2252 311
rect 2223 308 2252 310
rect 2223 307 2224 308
rect 2218 306 2224 307
rect 2251 307 2252 308
rect 2256 307 2257 311
rect 2251 306 2257 307
rect 2315 311 2321 312
rect 2315 307 2316 311
rect 2320 310 2321 311
rect 2338 311 2344 312
rect 2338 310 2339 311
rect 2320 308 2339 310
rect 2320 307 2321 308
rect 2315 306 2321 307
rect 2338 307 2339 308
rect 2343 307 2344 311
rect 2338 306 2344 307
rect 2346 311 2352 312
rect 2346 307 2347 311
rect 2351 310 2352 311
rect 2355 311 2361 312
rect 2355 310 2356 311
rect 2351 308 2356 310
rect 2351 307 2352 308
rect 2346 306 2352 307
rect 2355 307 2356 308
rect 2360 307 2361 311
rect 2355 306 2361 307
rect 134 303 140 304
rect 134 299 135 303
rect 139 299 140 303
rect 134 298 140 299
rect 182 303 188 304
rect 182 299 183 303
rect 187 299 188 303
rect 182 298 188 299
rect 254 303 260 304
rect 254 299 255 303
rect 259 299 260 303
rect 254 298 260 299
rect 326 303 332 304
rect 326 299 327 303
rect 331 299 332 303
rect 326 298 332 299
rect 390 303 396 304
rect 390 299 391 303
rect 395 299 396 303
rect 390 298 396 299
rect 446 303 452 304
rect 446 299 447 303
rect 451 299 452 303
rect 446 298 452 299
rect 502 303 508 304
rect 502 299 503 303
rect 507 299 508 303
rect 502 298 508 299
rect 550 303 556 304
rect 550 299 551 303
rect 555 299 556 303
rect 550 298 556 299
rect 590 303 596 304
rect 590 299 591 303
rect 595 299 596 303
rect 590 298 596 299
rect 630 303 636 304
rect 630 299 631 303
rect 635 299 636 303
rect 630 298 636 299
rect 678 303 684 304
rect 678 299 679 303
rect 683 299 684 303
rect 678 298 684 299
rect 726 303 732 304
rect 726 299 727 303
rect 731 299 732 303
rect 726 298 732 299
rect 774 303 780 304
rect 774 299 775 303
rect 779 299 780 303
rect 774 298 780 299
rect 822 303 828 304
rect 822 299 823 303
rect 827 299 828 303
rect 822 298 828 299
rect 870 303 876 304
rect 870 299 871 303
rect 875 299 876 303
rect 870 298 876 299
rect 918 303 924 304
rect 918 299 919 303
rect 923 299 924 303
rect 918 298 924 299
rect 1494 303 1500 304
rect 1494 299 1495 303
rect 1499 299 1500 303
rect 1494 298 1500 299
rect 1534 303 1540 304
rect 1534 299 1535 303
rect 1539 299 1540 303
rect 1534 298 1540 299
rect 1574 303 1580 304
rect 1574 299 1575 303
rect 1579 299 1580 303
rect 1574 298 1580 299
rect 1614 303 1620 304
rect 1614 299 1615 303
rect 1619 299 1620 303
rect 1614 298 1620 299
rect 1654 303 1660 304
rect 1654 299 1655 303
rect 1659 299 1660 303
rect 1654 298 1660 299
rect 1694 303 1700 304
rect 1694 299 1695 303
rect 1699 299 1700 303
rect 1694 298 1700 299
rect 1742 303 1748 304
rect 1742 299 1743 303
rect 1747 299 1748 303
rect 1742 298 1748 299
rect 1798 303 1804 304
rect 1798 299 1799 303
rect 1803 299 1804 303
rect 1798 298 1804 299
rect 1862 303 1868 304
rect 1862 299 1863 303
rect 1867 299 1868 303
rect 1862 298 1868 299
rect 1934 303 1940 304
rect 1934 299 1935 303
rect 1939 299 1940 303
rect 1934 298 1940 299
rect 2006 303 2012 304
rect 2006 299 2007 303
rect 2011 299 2012 303
rect 2006 298 2012 299
rect 2070 303 2076 304
rect 2070 299 2071 303
rect 2075 299 2076 303
rect 2070 298 2076 299
rect 2134 303 2140 304
rect 2134 299 2135 303
rect 2139 299 2140 303
rect 2134 298 2140 299
rect 2190 303 2196 304
rect 2190 299 2191 303
rect 2195 299 2196 303
rect 2190 298 2196 299
rect 2254 303 2260 304
rect 2254 299 2255 303
rect 2259 299 2260 303
rect 2254 298 2260 299
rect 2318 303 2324 304
rect 2318 299 2319 303
rect 2323 299 2324 303
rect 2318 298 2324 299
rect 2358 303 2364 304
rect 2358 299 2359 303
rect 2363 299 2364 303
rect 2358 298 2364 299
rect 806 283 812 284
rect 110 280 116 281
rect 110 276 111 280
rect 115 276 116 280
rect 806 279 807 283
rect 811 282 812 283
rect 811 280 918 282
rect 811 279 812 280
rect 806 278 812 279
rect 110 275 116 276
rect 159 275 168 276
rect 159 271 160 275
rect 167 271 168 275
rect 159 270 168 271
rect 207 275 216 276
rect 207 271 208 275
rect 215 271 216 275
rect 207 270 216 271
rect 278 275 285 276
rect 278 271 279 275
rect 284 271 285 275
rect 278 270 285 271
rect 351 275 360 276
rect 351 271 352 275
rect 359 271 360 275
rect 351 270 360 271
rect 415 275 424 276
rect 415 271 416 275
rect 423 271 424 275
rect 415 270 424 271
rect 471 275 480 276
rect 471 271 472 275
rect 479 271 480 275
rect 471 270 480 271
rect 527 275 533 276
rect 527 271 528 275
rect 532 274 533 275
rect 535 275 541 276
rect 535 274 536 275
rect 532 272 536 274
rect 532 271 533 272
rect 527 270 533 271
rect 535 271 536 272
rect 540 271 541 275
rect 535 270 541 271
rect 566 275 572 276
rect 566 271 567 275
rect 571 274 572 275
rect 575 275 581 276
rect 575 274 576 275
rect 571 272 576 274
rect 571 271 572 272
rect 566 270 572 271
rect 575 271 576 272
rect 580 271 581 275
rect 575 270 581 271
rect 610 275 621 276
rect 610 271 611 275
rect 615 271 616 275
rect 620 271 621 275
rect 610 270 621 271
rect 626 275 632 276
rect 626 271 627 275
rect 631 274 632 275
rect 655 275 661 276
rect 655 274 656 275
rect 631 272 656 274
rect 631 271 632 272
rect 626 270 632 271
rect 655 271 656 272
rect 660 271 661 275
rect 655 270 661 271
rect 666 275 672 276
rect 666 271 667 275
rect 671 274 672 275
rect 703 275 709 276
rect 703 274 704 275
rect 671 272 704 274
rect 671 271 672 272
rect 666 270 672 271
rect 703 271 704 272
rect 708 271 709 275
rect 703 270 709 271
rect 714 275 720 276
rect 714 271 715 275
rect 719 274 720 275
rect 751 275 757 276
rect 751 274 752 275
rect 719 272 752 274
rect 719 271 720 272
rect 714 270 720 271
rect 751 271 752 272
rect 756 271 757 275
rect 751 270 757 271
rect 762 275 768 276
rect 762 271 763 275
rect 767 274 768 275
rect 799 275 805 276
rect 799 274 800 275
rect 767 272 800 274
rect 767 271 768 272
rect 762 270 768 271
rect 799 271 800 272
rect 804 271 805 275
rect 799 270 805 271
rect 847 275 853 276
rect 847 271 848 275
rect 852 274 853 275
rect 858 275 864 276
rect 858 274 859 275
rect 852 272 859 274
rect 852 271 853 272
rect 847 270 853 271
rect 858 271 859 272
rect 863 271 864 275
rect 858 270 864 271
rect 895 275 901 276
rect 895 271 896 275
rect 900 274 901 275
rect 906 275 912 276
rect 906 274 907 275
rect 900 272 907 274
rect 900 271 901 272
rect 895 270 901 271
rect 906 271 907 272
rect 911 271 912 275
rect 916 274 918 280
rect 1238 280 1244 281
rect 1238 276 1239 280
rect 1243 276 1244 280
rect 943 275 949 276
rect 1238 275 1244 276
rect 1278 280 1284 281
rect 1278 276 1279 280
rect 1283 276 1284 280
rect 2406 280 2412 281
rect 2406 276 2407 280
rect 2411 276 2412 280
rect 1278 275 1284 276
rect 1519 275 1528 276
rect 943 274 944 275
rect 916 272 944 274
rect 906 270 912 271
rect 943 271 944 272
rect 948 271 949 275
rect 943 270 949 271
rect 1519 271 1520 275
rect 1527 271 1528 275
rect 1519 270 1528 271
rect 1559 275 1568 276
rect 1559 271 1560 275
rect 1567 271 1568 275
rect 1559 270 1568 271
rect 1599 275 1608 276
rect 1599 271 1600 275
rect 1607 271 1608 275
rect 1599 270 1608 271
rect 1639 275 1648 276
rect 1639 271 1640 275
rect 1647 271 1648 275
rect 1639 270 1648 271
rect 1679 275 1688 276
rect 1679 271 1680 275
rect 1687 271 1688 275
rect 1679 270 1688 271
rect 1719 275 1728 276
rect 1719 271 1720 275
rect 1727 271 1728 275
rect 1767 275 1773 276
rect 1767 274 1768 275
rect 1719 270 1728 271
rect 1732 272 1768 274
rect 1710 267 1716 268
rect 110 263 116 264
rect 110 259 111 263
rect 115 259 116 263
rect 110 258 116 259
rect 1238 263 1244 264
rect 1238 259 1239 263
rect 1243 259 1244 263
rect 1238 258 1244 259
rect 1278 263 1284 264
rect 1278 259 1279 263
rect 1283 259 1284 263
rect 1710 263 1711 267
rect 1715 266 1716 267
rect 1732 266 1734 272
rect 1767 271 1768 272
rect 1772 271 1773 275
rect 1767 270 1773 271
rect 1823 275 1832 276
rect 1823 271 1824 275
rect 1831 271 1832 275
rect 1823 270 1832 271
rect 1887 275 1893 276
rect 1887 271 1888 275
rect 1892 274 1893 275
rect 1895 275 1901 276
rect 1895 274 1896 275
rect 1892 272 1896 274
rect 1892 271 1893 272
rect 1887 270 1893 271
rect 1895 271 1896 272
rect 1900 271 1901 275
rect 1895 270 1901 271
rect 1959 275 1965 276
rect 1959 271 1960 275
rect 1964 274 1965 275
rect 1974 275 1980 276
rect 1974 274 1975 275
rect 1964 272 1975 274
rect 1964 271 1965 272
rect 1959 270 1965 271
rect 1974 271 1975 272
rect 1979 271 1980 275
rect 1974 270 1980 271
rect 1982 275 1988 276
rect 1982 271 1983 275
rect 1987 274 1988 275
rect 2031 275 2037 276
rect 2031 274 2032 275
rect 1987 272 2032 274
rect 1987 271 1988 272
rect 1982 270 1988 271
rect 2031 271 2032 272
rect 2036 271 2037 275
rect 2031 270 2037 271
rect 2095 275 2104 276
rect 2095 271 2096 275
rect 2103 271 2104 275
rect 2095 270 2104 271
rect 2159 275 2168 276
rect 2159 271 2160 275
rect 2167 271 2168 275
rect 2159 270 2168 271
rect 2215 275 2224 276
rect 2215 271 2216 275
rect 2223 271 2224 275
rect 2215 270 2224 271
rect 2279 275 2288 276
rect 2279 271 2280 275
rect 2287 271 2288 275
rect 2279 270 2288 271
rect 2343 275 2352 276
rect 2343 271 2344 275
rect 2351 271 2352 275
rect 2343 270 2352 271
rect 2374 275 2380 276
rect 2374 271 2375 275
rect 2379 274 2380 275
rect 2383 275 2389 276
rect 2406 275 2412 276
rect 2383 274 2384 275
rect 2379 272 2384 274
rect 2379 271 2380 272
rect 2374 270 2380 271
rect 2383 271 2384 272
rect 2388 271 2389 275
rect 2383 270 2389 271
rect 1715 264 1734 266
rect 1715 263 1716 264
rect 1710 262 1716 263
rect 2406 263 2412 264
rect 1278 258 1284 259
rect 2406 259 2407 263
rect 2411 259 2412 263
rect 2406 258 2412 259
rect 134 256 140 257
rect 134 252 135 256
rect 139 252 140 256
rect 134 251 140 252
rect 182 256 188 257
rect 182 252 183 256
rect 187 252 188 256
rect 182 251 188 252
rect 254 256 260 257
rect 254 252 255 256
rect 259 252 260 256
rect 254 251 260 252
rect 326 256 332 257
rect 326 252 327 256
rect 331 252 332 256
rect 326 251 332 252
rect 390 256 396 257
rect 390 252 391 256
rect 395 252 396 256
rect 390 251 396 252
rect 446 256 452 257
rect 446 252 447 256
rect 451 252 452 256
rect 446 251 452 252
rect 502 256 508 257
rect 502 252 503 256
rect 507 252 508 256
rect 502 251 508 252
rect 550 256 556 257
rect 550 252 551 256
rect 555 252 556 256
rect 550 251 556 252
rect 590 256 596 257
rect 590 252 591 256
rect 595 252 596 256
rect 590 251 596 252
rect 630 256 636 257
rect 630 252 631 256
rect 635 252 636 256
rect 630 251 636 252
rect 678 256 684 257
rect 678 252 679 256
rect 683 252 684 256
rect 678 251 684 252
rect 726 256 732 257
rect 726 252 727 256
rect 731 252 732 256
rect 726 251 732 252
rect 774 256 780 257
rect 774 252 775 256
rect 779 252 780 256
rect 774 251 780 252
rect 822 256 828 257
rect 822 252 823 256
rect 827 252 828 256
rect 822 251 828 252
rect 870 256 876 257
rect 870 252 871 256
rect 875 252 876 256
rect 870 251 876 252
rect 918 256 924 257
rect 918 252 919 256
rect 923 252 924 256
rect 918 251 924 252
rect 1494 256 1500 257
rect 1494 252 1495 256
rect 1499 252 1500 256
rect 1494 251 1500 252
rect 1534 256 1540 257
rect 1534 252 1535 256
rect 1539 252 1540 256
rect 1534 251 1540 252
rect 1574 256 1580 257
rect 1574 252 1575 256
rect 1579 252 1580 256
rect 1574 251 1580 252
rect 1614 256 1620 257
rect 1614 252 1615 256
rect 1619 252 1620 256
rect 1614 251 1620 252
rect 1654 256 1660 257
rect 1654 252 1655 256
rect 1659 252 1660 256
rect 1654 251 1660 252
rect 1694 256 1700 257
rect 1694 252 1695 256
rect 1699 252 1700 256
rect 1694 251 1700 252
rect 1742 256 1748 257
rect 1742 252 1743 256
rect 1747 252 1748 256
rect 1742 251 1748 252
rect 1798 256 1804 257
rect 1798 252 1799 256
rect 1803 252 1804 256
rect 1798 251 1804 252
rect 1862 256 1868 257
rect 1862 252 1863 256
rect 1867 252 1868 256
rect 1862 251 1868 252
rect 1934 256 1940 257
rect 1934 252 1935 256
rect 1939 252 1940 256
rect 1934 251 1940 252
rect 2006 256 2012 257
rect 2006 252 2007 256
rect 2011 252 2012 256
rect 2006 251 2012 252
rect 2070 256 2076 257
rect 2070 252 2071 256
rect 2075 252 2076 256
rect 2070 251 2076 252
rect 2134 256 2140 257
rect 2134 252 2135 256
rect 2139 252 2140 256
rect 2134 251 2140 252
rect 2190 256 2196 257
rect 2190 252 2191 256
rect 2195 252 2196 256
rect 2190 251 2196 252
rect 2254 256 2260 257
rect 2254 252 2255 256
rect 2259 252 2260 256
rect 2254 251 2260 252
rect 2318 256 2324 257
rect 2318 252 2319 256
rect 2323 252 2324 256
rect 2318 251 2324 252
rect 2358 256 2364 257
rect 2358 252 2359 256
rect 2363 252 2364 256
rect 2358 251 2364 252
rect 1366 240 1372 241
rect 134 236 140 237
rect 134 232 135 236
rect 139 232 140 236
rect 134 231 140 232
rect 174 236 180 237
rect 174 232 175 236
rect 179 232 180 236
rect 174 231 180 232
rect 246 236 252 237
rect 246 232 247 236
rect 251 232 252 236
rect 246 231 252 232
rect 326 236 332 237
rect 326 232 327 236
rect 331 232 332 236
rect 326 231 332 232
rect 414 236 420 237
rect 414 232 415 236
rect 419 232 420 236
rect 414 231 420 232
rect 494 236 500 237
rect 494 232 495 236
rect 499 232 500 236
rect 494 231 500 232
rect 574 236 580 237
rect 574 232 575 236
rect 579 232 580 236
rect 574 231 580 232
rect 654 236 660 237
rect 654 232 655 236
rect 659 232 660 236
rect 654 231 660 232
rect 726 236 732 237
rect 726 232 727 236
rect 731 232 732 236
rect 726 231 732 232
rect 790 236 796 237
rect 790 232 791 236
rect 795 232 796 236
rect 790 231 796 232
rect 846 236 852 237
rect 846 232 847 236
rect 851 232 852 236
rect 846 231 852 232
rect 902 236 908 237
rect 902 232 903 236
rect 907 232 908 236
rect 902 231 908 232
rect 958 236 964 237
rect 958 232 959 236
rect 963 232 964 236
rect 958 231 964 232
rect 1022 236 1028 237
rect 1022 232 1023 236
rect 1027 232 1028 236
rect 1366 236 1367 240
rect 1371 236 1372 240
rect 1366 235 1372 236
rect 1406 240 1412 241
rect 1406 236 1407 240
rect 1411 236 1412 240
rect 1406 235 1412 236
rect 1446 240 1452 241
rect 1446 236 1447 240
rect 1451 236 1452 240
rect 1446 235 1452 236
rect 1494 240 1500 241
rect 1494 236 1495 240
rect 1499 236 1500 240
rect 1494 235 1500 236
rect 1550 240 1556 241
rect 1550 236 1551 240
rect 1555 236 1556 240
rect 1550 235 1556 236
rect 1606 240 1612 241
rect 1606 236 1607 240
rect 1611 236 1612 240
rect 1606 235 1612 236
rect 1670 240 1676 241
rect 1670 236 1671 240
rect 1675 236 1676 240
rect 1670 235 1676 236
rect 1734 240 1740 241
rect 1734 236 1735 240
rect 1739 236 1740 240
rect 1734 235 1740 236
rect 1806 240 1812 241
rect 1806 236 1807 240
rect 1811 236 1812 240
rect 1806 235 1812 236
rect 1886 240 1892 241
rect 1886 236 1887 240
rect 1891 236 1892 240
rect 1886 235 1892 236
rect 1974 240 1980 241
rect 1974 236 1975 240
rect 1979 236 1980 240
rect 1974 235 1980 236
rect 2070 240 2076 241
rect 2070 236 2071 240
rect 2075 236 2076 240
rect 2070 235 2076 236
rect 2166 240 2172 241
rect 2166 236 2167 240
rect 2171 236 2172 240
rect 2166 235 2172 236
rect 2270 240 2276 241
rect 2270 236 2271 240
rect 2275 236 2276 240
rect 2270 235 2276 236
rect 2358 240 2364 241
rect 2358 236 2359 240
rect 2363 236 2364 240
rect 2358 235 2364 236
rect 1022 231 1028 232
rect 1278 233 1284 234
rect 110 229 116 230
rect 110 225 111 229
rect 115 225 116 229
rect 110 224 116 225
rect 1238 229 1244 230
rect 1238 225 1239 229
rect 1243 225 1244 229
rect 1278 229 1279 233
rect 1283 229 1284 233
rect 1278 228 1284 229
rect 2406 233 2412 234
rect 2406 229 2407 233
rect 2411 229 2412 233
rect 2406 228 2412 229
rect 1238 224 1244 225
rect 1391 219 1400 220
rect 1278 216 1284 217
rect 154 215 165 216
rect 110 212 116 213
rect 110 208 111 212
rect 115 208 116 212
rect 154 211 155 215
rect 159 211 160 215
rect 164 211 165 215
rect 154 210 165 211
rect 170 215 176 216
rect 170 211 171 215
rect 175 214 176 215
rect 199 215 205 216
rect 199 214 200 215
rect 175 212 200 214
rect 175 211 176 212
rect 170 210 176 211
rect 199 211 200 212
rect 204 211 205 215
rect 199 210 205 211
rect 271 215 277 216
rect 271 211 272 215
rect 276 214 277 215
rect 318 215 324 216
rect 318 214 319 215
rect 276 212 319 214
rect 276 211 277 212
rect 271 210 277 211
rect 318 211 319 212
rect 323 211 324 215
rect 318 210 324 211
rect 351 215 357 216
rect 351 211 352 215
rect 356 211 357 215
rect 351 210 357 211
rect 439 215 445 216
rect 439 211 440 215
rect 444 214 445 215
rect 486 215 492 216
rect 486 214 487 215
rect 444 212 487 214
rect 444 211 445 212
rect 439 210 445 211
rect 486 211 487 212
rect 491 211 492 215
rect 486 210 492 211
rect 518 215 525 216
rect 518 211 519 215
rect 524 211 525 215
rect 599 215 605 216
rect 599 214 600 215
rect 518 210 525 211
rect 528 212 600 214
rect 110 207 116 208
rect 182 207 188 208
rect 182 203 183 207
rect 187 206 188 207
rect 353 206 355 210
rect 187 204 355 206
rect 422 207 428 208
rect 187 203 188 204
rect 182 202 188 203
rect 422 203 423 207
rect 427 206 428 207
rect 528 206 530 212
rect 599 211 600 212
rect 604 211 605 215
rect 599 210 605 211
rect 679 215 685 216
rect 679 211 680 215
rect 684 214 685 215
rect 718 215 724 216
rect 718 214 719 215
rect 684 212 719 214
rect 684 211 685 212
rect 679 210 685 211
rect 718 211 719 212
rect 723 211 724 215
rect 718 210 724 211
rect 751 215 757 216
rect 751 211 752 215
rect 756 214 757 215
rect 782 215 788 216
rect 782 214 783 215
rect 756 212 783 214
rect 756 211 757 212
rect 751 210 757 211
rect 782 211 783 212
rect 787 211 788 215
rect 782 210 788 211
rect 814 215 821 216
rect 814 211 815 215
rect 820 211 821 215
rect 871 215 877 216
rect 871 214 872 215
rect 814 210 821 211
rect 824 212 872 214
rect 427 204 530 206
rect 662 207 668 208
rect 427 203 428 204
rect 422 202 428 203
rect 662 203 663 207
rect 667 206 668 207
rect 824 206 826 212
rect 871 211 872 212
rect 876 211 877 215
rect 871 210 877 211
rect 927 215 933 216
rect 927 211 928 215
rect 932 214 933 215
rect 942 215 948 216
rect 942 214 943 215
rect 932 212 943 214
rect 932 211 933 212
rect 927 210 933 211
rect 942 211 943 212
rect 947 211 948 215
rect 942 210 948 211
rect 983 215 989 216
rect 983 211 984 215
rect 988 214 989 215
rect 1014 215 1020 216
rect 1014 214 1015 215
rect 988 212 1015 214
rect 988 211 989 212
rect 983 210 989 211
rect 1014 211 1015 212
rect 1019 211 1020 215
rect 1047 215 1053 216
rect 1047 214 1048 215
rect 1014 210 1020 211
rect 1024 212 1048 214
rect 667 204 826 206
rect 854 207 860 208
rect 667 203 668 204
rect 662 202 668 203
rect 854 203 855 207
rect 859 206 860 207
rect 1024 206 1026 212
rect 1047 211 1048 212
rect 1052 211 1053 215
rect 1047 210 1053 211
rect 1238 212 1244 213
rect 1238 208 1239 212
rect 1243 208 1244 212
rect 1278 212 1279 216
rect 1283 212 1284 216
rect 1391 215 1392 219
rect 1399 215 1400 219
rect 1391 214 1400 215
rect 1431 219 1440 220
rect 1431 215 1432 219
rect 1439 215 1440 219
rect 1431 214 1440 215
rect 1471 219 1477 220
rect 1471 215 1472 219
rect 1476 218 1477 219
rect 1510 219 1516 220
rect 1510 218 1511 219
rect 1476 216 1511 218
rect 1476 215 1477 216
rect 1471 214 1477 215
rect 1510 215 1511 216
rect 1515 215 1516 219
rect 1510 214 1516 215
rect 1519 219 1525 220
rect 1519 215 1520 219
rect 1524 215 1525 219
rect 1519 214 1525 215
rect 1527 219 1533 220
rect 1527 215 1528 219
rect 1532 218 1533 219
rect 1575 219 1581 220
rect 1575 218 1576 219
rect 1532 216 1576 218
rect 1532 215 1533 216
rect 1527 214 1533 215
rect 1575 215 1576 216
rect 1580 215 1581 219
rect 1575 214 1581 215
rect 1583 219 1589 220
rect 1583 215 1584 219
rect 1588 218 1589 219
rect 1631 219 1637 220
rect 1631 218 1632 219
rect 1588 216 1632 218
rect 1588 215 1589 216
rect 1583 214 1589 215
rect 1631 215 1632 216
rect 1636 215 1637 219
rect 1631 214 1637 215
rect 1642 219 1648 220
rect 1642 215 1643 219
rect 1647 218 1648 219
rect 1695 219 1701 220
rect 1695 218 1696 219
rect 1647 216 1696 218
rect 1647 215 1648 216
rect 1642 214 1648 215
rect 1695 215 1696 216
rect 1700 215 1701 219
rect 1695 214 1701 215
rect 1759 219 1765 220
rect 1759 215 1760 219
rect 1764 218 1765 219
rect 1798 219 1804 220
rect 1798 218 1799 219
rect 1764 216 1799 218
rect 1764 215 1765 216
rect 1759 214 1765 215
rect 1798 215 1799 216
rect 1803 215 1804 219
rect 1798 214 1804 215
rect 1831 219 1837 220
rect 1831 215 1832 219
rect 1836 218 1837 219
rect 1878 219 1884 220
rect 1878 218 1879 219
rect 1836 216 1879 218
rect 1836 215 1837 216
rect 1831 214 1837 215
rect 1878 215 1879 216
rect 1883 215 1884 219
rect 1878 214 1884 215
rect 1911 219 1917 220
rect 1911 215 1912 219
rect 1916 218 1917 219
rect 1966 219 1972 220
rect 1966 218 1967 219
rect 1916 216 1967 218
rect 1916 215 1917 216
rect 1911 214 1917 215
rect 1966 215 1967 216
rect 1971 215 1972 219
rect 1966 214 1972 215
rect 1990 219 1996 220
rect 1990 215 1991 219
rect 1995 218 1996 219
rect 1999 219 2005 220
rect 1999 218 2000 219
rect 1995 216 2000 218
rect 1995 215 1996 216
rect 1990 214 1996 215
rect 1999 215 2000 216
rect 2004 215 2005 219
rect 1999 214 2005 215
rect 2090 219 2101 220
rect 2090 215 2091 219
rect 2095 215 2096 219
rect 2100 215 2101 219
rect 2090 214 2101 215
rect 2103 219 2109 220
rect 2103 215 2104 219
rect 2108 218 2109 219
rect 2191 219 2197 220
rect 2191 218 2192 219
rect 2108 216 2192 218
rect 2108 215 2109 216
rect 2103 214 2109 215
rect 2191 215 2192 216
rect 2196 215 2197 219
rect 2191 214 2197 215
rect 2199 219 2205 220
rect 2199 215 2200 219
rect 2204 218 2205 219
rect 2295 219 2301 220
rect 2295 218 2296 219
rect 2204 216 2296 218
rect 2204 215 2205 216
rect 2199 214 2205 215
rect 2295 215 2296 216
rect 2300 215 2301 219
rect 2295 214 2301 215
rect 2366 219 2372 220
rect 2366 215 2367 219
rect 2371 218 2372 219
rect 2383 219 2389 220
rect 2383 218 2384 219
rect 2371 216 2384 218
rect 2371 215 2372 216
rect 2366 214 2372 215
rect 2383 215 2384 216
rect 2388 215 2389 219
rect 2383 214 2389 215
rect 2406 216 2412 217
rect 1278 211 1284 212
rect 1374 211 1380 212
rect 1238 207 1244 208
rect 1374 207 1375 211
rect 1379 210 1380 211
rect 1521 210 1523 214
rect 2406 212 2407 216
rect 2411 212 2412 216
rect 2406 211 2412 212
rect 1379 208 1523 210
rect 1379 207 1380 208
rect 1374 206 1380 207
rect 859 204 1026 206
rect 859 203 860 204
rect 854 202 860 203
rect 1366 193 1372 194
rect 134 189 140 190
rect 134 185 135 189
rect 139 185 140 189
rect 134 184 140 185
rect 174 189 180 190
rect 174 185 175 189
rect 179 185 180 189
rect 174 184 180 185
rect 246 189 252 190
rect 246 185 247 189
rect 251 185 252 189
rect 246 184 252 185
rect 326 189 332 190
rect 326 185 327 189
rect 331 185 332 189
rect 326 184 332 185
rect 414 189 420 190
rect 414 185 415 189
rect 419 185 420 189
rect 414 184 420 185
rect 494 189 500 190
rect 494 185 495 189
rect 499 185 500 189
rect 494 184 500 185
rect 574 189 580 190
rect 574 185 575 189
rect 579 185 580 189
rect 574 184 580 185
rect 654 189 660 190
rect 654 185 655 189
rect 659 185 660 189
rect 654 184 660 185
rect 726 189 732 190
rect 726 185 727 189
rect 731 185 732 189
rect 726 184 732 185
rect 790 189 796 190
rect 790 185 791 189
rect 795 185 796 189
rect 790 184 796 185
rect 846 189 852 190
rect 846 185 847 189
rect 851 185 852 189
rect 846 184 852 185
rect 902 189 908 190
rect 902 185 903 189
rect 907 185 908 189
rect 902 184 908 185
rect 958 189 964 190
rect 958 185 959 189
rect 963 185 964 189
rect 958 184 964 185
rect 1022 189 1028 190
rect 1022 185 1023 189
rect 1027 185 1028 189
rect 1366 189 1367 193
rect 1371 189 1372 193
rect 1366 188 1372 189
rect 1406 193 1412 194
rect 1406 189 1407 193
rect 1411 189 1412 193
rect 1406 188 1412 189
rect 1446 193 1452 194
rect 1446 189 1447 193
rect 1451 189 1452 193
rect 1446 188 1452 189
rect 1494 193 1500 194
rect 1494 189 1495 193
rect 1499 189 1500 193
rect 1494 188 1500 189
rect 1550 193 1556 194
rect 1550 189 1551 193
rect 1555 189 1556 193
rect 1550 188 1556 189
rect 1606 193 1612 194
rect 1606 189 1607 193
rect 1611 189 1612 193
rect 1606 188 1612 189
rect 1670 193 1676 194
rect 1670 189 1671 193
rect 1675 189 1676 193
rect 1670 188 1676 189
rect 1734 193 1740 194
rect 1734 189 1735 193
rect 1739 189 1740 193
rect 1734 188 1740 189
rect 1806 193 1812 194
rect 1806 189 1807 193
rect 1811 189 1812 193
rect 1806 188 1812 189
rect 1886 193 1892 194
rect 1886 189 1887 193
rect 1891 189 1892 193
rect 1886 188 1892 189
rect 1974 193 1980 194
rect 1974 189 1975 193
rect 1979 189 1980 193
rect 1974 188 1980 189
rect 2070 193 2076 194
rect 2070 189 2071 193
rect 2075 189 2076 193
rect 2070 188 2076 189
rect 2166 193 2172 194
rect 2166 189 2167 193
rect 2171 189 2172 193
rect 2166 188 2172 189
rect 2270 193 2276 194
rect 2270 189 2271 193
rect 2275 189 2276 193
rect 2270 188 2276 189
rect 2358 193 2364 194
rect 2358 189 2359 193
rect 2363 189 2364 193
rect 2358 188 2364 189
rect 1022 184 1028 185
rect 1363 183 1369 184
rect 131 179 137 180
rect 131 175 132 179
rect 136 178 137 179
rect 162 179 168 180
rect 162 178 163 179
rect 136 176 163 178
rect 136 175 137 176
rect 131 174 137 175
rect 162 175 163 176
rect 167 175 168 179
rect 162 174 168 175
rect 171 179 177 180
rect 171 175 172 179
rect 176 178 177 179
rect 182 179 188 180
rect 182 178 183 179
rect 176 176 183 178
rect 176 175 177 176
rect 171 174 177 175
rect 182 175 183 176
rect 187 175 188 179
rect 182 174 188 175
rect 238 179 249 180
rect 238 175 239 179
rect 243 175 244 179
rect 248 175 249 179
rect 238 174 249 175
rect 318 179 329 180
rect 318 175 319 179
rect 323 175 324 179
rect 328 175 329 179
rect 318 174 329 175
rect 411 179 417 180
rect 411 175 412 179
rect 416 178 417 179
rect 422 179 428 180
rect 422 178 423 179
rect 416 176 423 178
rect 416 175 417 176
rect 411 174 417 175
rect 422 175 423 176
rect 427 175 428 179
rect 422 174 428 175
rect 486 179 497 180
rect 486 175 487 179
rect 491 175 492 179
rect 496 175 497 179
rect 486 174 497 175
rect 566 179 577 180
rect 566 175 567 179
rect 571 175 572 179
rect 576 175 577 179
rect 566 174 577 175
rect 651 179 657 180
rect 651 175 652 179
rect 656 178 657 179
rect 662 179 668 180
rect 662 178 663 179
rect 656 176 663 178
rect 656 175 657 176
rect 651 174 657 175
rect 662 175 663 176
rect 667 175 668 179
rect 662 174 668 175
rect 718 179 729 180
rect 718 175 719 179
rect 723 175 724 179
rect 728 175 729 179
rect 718 174 729 175
rect 782 179 793 180
rect 782 175 783 179
rect 787 175 788 179
rect 792 175 793 179
rect 782 174 793 175
rect 843 179 849 180
rect 843 175 844 179
rect 848 178 849 179
rect 854 179 860 180
rect 854 178 855 179
rect 848 176 855 178
rect 848 175 849 176
rect 843 174 849 175
rect 854 175 855 176
rect 859 175 860 179
rect 899 179 905 180
rect 899 178 900 179
rect 854 174 860 175
rect 864 176 900 178
rect 750 171 756 172
rect 750 167 751 171
rect 755 170 756 171
rect 864 170 866 176
rect 899 175 900 176
rect 904 175 905 179
rect 899 174 905 175
rect 942 179 948 180
rect 942 175 943 179
rect 947 178 948 179
rect 955 179 961 180
rect 955 178 956 179
rect 947 176 956 178
rect 947 175 948 176
rect 942 174 948 175
rect 955 175 956 176
rect 960 175 961 179
rect 955 174 961 175
rect 1014 179 1025 180
rect 1014 175 1015 179
rect 1019 175 1020 179
rect 1024 175 1025 179
rect 1363 179 1364 183
rect 1368 182 1369 183
rect 1374 183 1380 184
rect 1374 182 1375 183
rect 1368 180 1375 182
rect 1368 179 1369 180
rect 1363 178 1369 179
rect 1374 179 1375 180
rect 1379 179 1380 183
rect 1374 178 1380 179
rect 1394 183 1400 184
rect 1394 179 1395 183
rect 1399 182 1400 183
rect 1403 183 1409 184
rect 1403 182 1404 183
rect 1399 180 1404 182
rect 1399 179 1400 180
rect 1394 178 1400 179
rect 1403 179 1404 180
rect 1408 179 1409 183
rect 1403 178 1409 179
rect 1434 183 1440 184
rect 1434 179 1435 183
rect 1439 182 1440 183
rect 1443 183 1449 184
rect 1443 182 1444 183
rect 1439 180 1444 182
rect 1439 179 1440 180
rect 1434 178 1440 179
rect 1443 179 1444 180
rect 1448 179 1449 183
rect 1443 178 1449 179
rect 1491 183 1497 184
rect 1491 179 1492 183
rect 1496 182 1497 183
rect 1527 183 1533 184
rect 1527 182 1528 183
rect 1496 180 1528 182
rect 1496 179 1497 180
rect 1491 178 1497 179
rect 1527 179 1528 180
rect 1532 179 1533 183
rect 1527 178 1533 179
rect 1547 183 1553 184
rect 1547 179 1548 183
rect 1552 182 1553 183
rect 1583 183 1589 184
rect 1583 182 1584 183
rect 1552 180 1584 182
rect 1552 179 1553 180
rect 1547 178 1553 179
rect 1583 179 1584 180
rect 1588 179 1589 183
rect 1583 178 1589 179
rect 1603 183 1609 184
rect 1603 179 1604 183
rect 1608 182 1609 183
rect 1642 183 1648 184
rect 1642 182 1643 183
rect 1608 180 1643 182
rect 1608 179 1609 180
rect 1603 178 1609 179
rect 1642 179 1643 180
rect 1647 179 1648 183
rect 1642 178 1648 179
rect 1667 183 1673 184
rect 1667 179 1668 183
rect 1672 182 1673 183
rect 1710 183 1716 184
rect 1710 182 1711 183
rect 1672 180 1711 182
rect 1672 179 1673 180
rect 1667 178 1673 179
rect 1710 179 1711 180
rect 1715 179 1716 183
rect 1710 178 1716 179
rect 1731 183 1737 184
rect 1731 179 1732 183
rect 1736 182 1737 183
rect 1742 183 1748 184
rect 1742 182 1743 183
rect 1736 180 1743 182
rect 1736 179 1737 180
rect 1731 178 1737 179
rect 1742 179 1743 180
rect 1747 179 1748 183
rect 1742 178 1748 179
rect 1798 183 1809 184
rect 1798 179 1799 183
rect 1803 179 1804 183
rect 1808 179 1809 183
rect 1798 178 1809 179
rect 1878 183 1889 184
rect 1878 179 1879 183
rect 1883 179 1884 183
rect 1888 179 1889 183
rect 1878 178 1889 179
rect 1966 183 1977 184
rect 1966 179 1967 183
rect 1971 179 1972 183
rect 1976 179 1977 183
rect 1966 178 1977 179
rect 2067 183 2073 184
rect 2067 179 2068 183
rect 2072 182 2073 183
rect 2103 183 2109 184
rect 2103 182 2104 183
rect 2072 180 2104 182
rect 2072 179 2073 180
rect 2067 178 2073 179
rect 2103 179 2104 180
rect 2108 179 2109 183
rect 2103 178 2109 179
rect 2163 183 2169 184
rect 2163 179 2164 183
rect 2168 182 2169 183
rect 2199 183 2205 184
rect 2199 182 2200 183
rect 2168 180 2200 182
rect 2168 179 2169 180
rect 2163 178 2169 179
rect 2199 179 2200 180
rect 2204 179 2205 183
rect 2199 178 2205 179
rect 2242 183 2248 184
rect 2242 179 2243 183
rect 2247 182 2248 183
rect 2267 183 2273 184
rect 2267 182 2268 183
rect 2247 180 2268 182
rect 2247 179 2248 180
rect 2242 178 2248 179
rect 2267 179 2268 180
rect 2272 179 2273 183
rect 2267 178 2273 179
rect 2355 183 2361 184
rect 2355 179 2356 183
rect 2360 182 2361 183
rect 2374 183 2380 184
rect 2374 182 2375 183
rect 2360 180 2375 182
rect 2360 179 2361 180
rect 2355 178 2361 179
rect 2374 179 2375 180
rect 2379 179 2380 183
rect 2374 178 2380 179
rect 1014 174 1025 175
rect 755 168 866 170
rect 755 167 756 168
rect 750 166 756 167
rect 1990 163 1996 164
rect 1990 162 1991 163
rect 1708 160 1991 162
rect 1708 158 1710 160
rect 1990 159 1991 160
rect 1995 159 1996 163
rect 1990 158 1996 159
rect 1707 157 1713 158
rect 1299 155 1305 156
rect 1299 151 1300 155
rect 1304 154 1305 155
rect 1330 155 1336 156
rect 1330 154 1331 155
rect 1304 152 1331 154
rect 1304 151 1305 152
rect 1299 150 1305 151
rect 1330 151 1331 152
rect 1335 151 1336 155
rect 1330 150 1336 151
rect 1339 155 1345 156
rect 1339 151 1340 155
rect 1344 154 1345 155
rect 1358 155 1364 156
rect 1358 154 1359 155
rect 1344 152 1359 154
rect 1344 151 1345 152
rect 1339 150 1345 151
rect 1358 151 1359 152
rect 1363 151 1364 155
rect 1358 150 1364 151
rect 1379 155 1385 156
rect 1379 151 1380 155
rect 1384 154 1385 155
rect 1398 155 1404 156
rect 1398 154 1399 155
rect 1384 152 1399 154
rect 1384 151 1385 152
rect 1379 150 1385 151
rect 1398 151 1399 152
rect 1403 151 1404 155
rect 1398 150 1404 151
rect 1419 155 1425 156
rect 1419 151 1420 155
rect 1424 154 1425 155
rect 1438 155 1444 156
rect 1438 154 1439 155
rect 1424 152 1439 154
rect 1424 151 1425 152
rect 1419 150 1425 151
rect 1438 151 1439 152
rect 1443 151 1444 155
rect 1438 150 1444 151
rect 1459 155 1465 156
rect 1459 151 1460 155
rect 1464 154 1465 155
rect 1502 155 1508 156
rect 1502 154 1503 155
rect 1464 152 1503 154
rect 1464 151 1465 152
rect 1459 150 1465 151
rect 1502 151 1503 152
rect 1507 151 1508 155
rect 1502 150 1508 151
rect 1510 155 1521 156
rect 1510 151 1511 155
rect 1515 151 1516 155
rect 1520 151 1521 155
rect 1510 150 1521 151
rect 1551 155 1557 156
rect 1551 151 1552 155
rect 1556 154 1557 155
rect 1579 155 1585 156
rect 1579 154 1580 155
rect 1556 152 1580 154
rect 1556 151 1557 152
rect 1551 150 1557 151
rect 1579 151 1580 152
rect 1584 151 1585 155
rect 1579 150 1585 151
rect 1615 155 1621 156
rect 1615 151 1616 155
rect 1620 154 1621 155
rect 1643 155 1649 156
rect 1643 154 1644 155
rect 1620 152 1644 154
rect 1620 151 1621 152
rect 1615 150 1621 151
rect 1643 151 1644 152
rect 1648 151 1649 155
rect 1707 153 1708 157
rect 1712 153 1713 157
rect 1707 152 1713 153
rect 1751 155 1757 156
rect 1643 150 1649 151
rect 1751 151 1752 155
rect 1756 154 1757 155
rect 1763 155 1769 156
rect 1763 154 1764 155
rect 1756 152 1764 154
rect 1756 151 1757 152
rect 1751 150 1757 151
rect 1763 151 1764 152
rect 1768 151 1769 155
rect 1763 150 1769 151
rect 1799 155 1805 156
rect 1799 151 1800 155
rect 1804 154 1805 155
rect 1819 155 1825 156
rect 1819 154 1820 155
rect 1804 152 1820 154
rect 1804 151 1805 152
rect 1799 150 1805 151
rect 1819 151 1820 152
rect 1824 151 1825 155
rect 1819 150 1825 151
rect 1850 155 1856 156
rect 1850 151 1851 155
rect 1855 154 1856 155
rect 1867 155 1873 156
rect 1867 154 1868 155
rect 1855 152 1868 154
rect 1855 151 1856 152
rect 1850 150 1856 151
rect 1867 151 1868 152
rect 1872 151 1873 155
rect 1867 150 1873 151
rect 1898 155 1904 156
rect 1898 151 1899 155
rect 1903 154 1904 155
rect 1915 155 1921 156
rect 1915 154 1916 155
rect 1903 152 1916 154
rect 1903 151 1904 152
rect 1898 150 1904 151
rect 1915 151 1916 152
rect 1920 151 1921 155
rect 1915 150 1921 151
rect 1946 155 1952 156
rect 1946 151 1947 155
rect 1951 154 1952 155
rect 1963 155 1969 156
rect 1963 154 1964 155
rect 1951 152 1964 154
rect 1951 151 1952 152
rect 1946 150 1952 151
rect 1963 151 1964 152
rect 1968 151 1969 155
rect 1963 150 1969 151
rect 1994 155 2000 156
rect 1994 151 1995 155
rect 1999 154 2000 155
rect 2011 155 2017 156
rect 2011 154 2012 155
rect 1999 152 2012 154
rect 1999 151 2000 152
rect 1994 150 2000 151
rect 2011 151 2012 152
rect 2016 151 2017 155
rect 2011 150 2017 151
rect 2042 155 2048 156
rect 2042 151 2043 155
rect 2047 154 2048 155
rect 2059 155 2065 156
rect 2059 154 2060 155
rect 2047 152 2060 154
rect 2047 151 2048 152
rect 2042 150 2048 151
rect 2059 151 2060 152
rect 2064 151 2065 155
rect 2059 150 2065 151
rect 2090 155 2096 156
rect 2090 151 2091 155
rect 2095 154 2096 155
rect 2107 155 2113 156
rect 2107 154 2108 155
rect 2095 152 2108 154
rect 2095 151 2096 152
rect 2090 150 2096 151
rect 2107 151 2108 152
rect 2112 151 2113 155
rect 2107 150 2113 151
rect 2138 155 2144 156
rect 2138 151 2139 155
rect 2143 154 2144 155
rect 2155 155 2161 156
rect 2155 154 2156 155
rect 2143 152 2156 154
rect 2143 151 2144 152
rect 2138 150 2144 151
rect 2155 151 2156 152
rect 2160 151 2161 155
rect 2155 150 2161 151
rect 2186 155 2192 156
rect 2186 151 2187 155
rect 2191 154 2192 155
rect 2211 155 2217 156
rect 2211 154 2212 155
rect 2191 152 2212 154
rect 2191 151 2192 152
rect 2186 150 2192 151
rect 2211 151 2212 152
rect 2216 151 2217 155
rect 2211 150 2217 151
rect 2267 155 2273 156
rect 2267 151 2268 155
rect 2272 154 2273 155
rect 2306 155 2312 156
rect 2306 154 2307 155
rect 2272 152 2307 154
rect 2272 151 2273 152
rect 2267 150 2273 151
rect 2306 151 2307 152
rect 2311 151 2312 155
rect 2306 150 2312 151
rect 2315 155 2321 156
rect 2315 151 2316 155
rect 2320 154 2321 155
rect 2346 155 2352 156
rect 2346 154 2347 155
rect 2320 152 2347 154
rect 2320 151 2321 152
rect 2315 150 2321 151
rect 2346 151 2347 152
rect 2351 151 2352 155
rect 2346 150 2352 151
rect 2355 155 2361 156
rect 2355 151 2356 155
rect 2360 154 2361 155
rect 2366 155 2372 156
rect 2366 154 2367 155
rect 2360 152 2367 154
rect 2360 151 2361 152
rect 2355 150 2361 151
rect 2366 151 2367 152
rect 2371 151 2372 155
rect 2366 150 2372 151
rect 131 147 137 148
rect 131 143 132 147
rect 136 146 137 147
rect 150 147 156 148
rect 150 146 151 147
rect 136 144 151 146
rect 136 143 137 144
rect 131 142 137 143
rect 150 143 151 144
rect 155 143 156 147
rect 150 142 156 143
rect 158 147 164 148
rect 158 143 159 147
rect 163 146 164 147
rect 171 147 177 148
rect 171 146 172 147
rect 163 144 172 146
rect 163 143 164 144
rect 158 142 164 143
rect 171 143 172 144
rect 176 143 177 147
rect 171 142 177 143
rect 202 147 208 148
rect 202 143 203 147
rect 207 146 208 147
rect 211 147 217 148
rect 211 146 212 147
rect 207 144 212 146
rect 207 143 208 144
rect 202 142 208 143
rect 211 143 212 144
rect 216 143 217 147
rect 211 142 217 143
rect 251 147 257 148
rect 251 143 252 147
rect 256 146 257 147
rect 282 147 288 148
rect 282 146 283 147
rect 256 144 283 146
rect 256 143 257 144
rect 251 142 257 143
rect 282 143 283 144
rect 287 143 288 147
rect 282 142 288 143
rect 291 147 297 148
rect 291 143 292 147
rect 296 146 297 147
rect 318 147 324 148
rect 318 146 319 147
rect 296 144 319 146
rect 296 143 297 144
rect 291 142 297 143
rect 318 143 319 144
rect 323 143 324 147
rect 318 142 324 143
rect 331 147 337 148
rect 331 143 332 147
rect 336 146 337 147
rect 362 147 368 148
rect 362 146 363 147
rect 336 144 363 146
rect 336 143 337 144
rect 331 142 337 143
rect 362 143 363 144
rect 367 143 368 147
rect 362 142 368 143
rect 371 147 377 148
rect 371 143 372 147
rect 376 146 377 147
rect 407 147 413 148
rect 407 146 408 147
rect 376 144 408 146
rect 376 143 377 144
rect 371 142 377 143
rect 407 143 408 144
rect 412 143 413 147
rect 407 142 413 143
rect 419 147 425 148
rect 419 143 420 147
rect 424 146 425 147
rect 458 147 464 148
rect 458 146 459 147
rect 424 144 459 146
rect 424 143 425 144
rect 419 142 425 143
rect 458 143 459 144
rect 463 143 464 147
rect 458 142 464 143
rect 467 147 473 148
rect 467 143 468 147
rect 472 146 473 147
rect 510 147 516 148
rect 510 146 511 147
rect 472 144 511 146
rect 472 143 473 144
rect 467 142 473 143
rect 510 143 511 144
rect 515 143 516 147
rect 510 142 516 143
rect 518 147 529 148
rect 518 143 519 147
rect 523 143 524 147
rect 528 143 529 147
rect 518 142 529 143
rect 554 147 560 148
rect 554 143 555 147
rect 559 146 560 147
rect 579 147 585 148
rect 579 146 580 147
rect 559 144 580 146
rect 559 143 560 144
rect 554 142 560 143
rect 579 143 580 144
rect 584 143 585 147
rect 579 142 585 143
rect 627 147 633 148
rect 627 143 628 147
rect 632 146 633 147
rect 646 147 652 148
rect 646 146 647 147
rect 632 144 647 146
rect 632 143 633 144
rect 627 142 633 143
rect 646 143 647 144
rect 651 143 652 147
rect 646 142 652 143
rect 663 147 669 148
rect 663 143 664 147
rect 668 146 669 147
rect 675 147 681 148
rect 675 146 676 147
rect 668 144 676 146
rect 668 143 669 144
rect 663 142 669 143
rect 675 143 676 144
rect 680 143 681 147
rect 675 142 681 143
rect 706 147 712 148
rect 706 143 707 147
rect 711 146 712 147
rect 723 147 729 148
rect 723 146 724 147
rect 711 144 724 146
rect 711 143 712 144
rect 706 142 712 143
rect 723 143 724 144
rect 728 143 729 147
rect 723 142 729 143
rect 763 147 769 148
rect 763 143 764 147
rect 768 146 769 147
rect 782 147 788 148
rect 782 146 783 147
rect 768 144 783 146
rect 768 143 769 144
rect 763 142 769 143
rect 782 143 783 144
rect 787 143 788 147
rect 782 142 788 143
rect 803 147 809 148
rect 803 143 804 147
rect 808 146 809 147
rect 834 147 840 148
rect 834 146 835 147
rect 808 144 835 146
rect 808 143 809 144
rect 803 142 809 143
rect 834 143 835 144
rect 839 143 840 147
rect 834 142 840 143
rect 843 147 849 148
rect 843 143 844 147
rect 848 146 849 147
rect 874 147 880 148
rect 874 146 875 147
rect 848 144 875 146
rect 848 143 849 144
rect 843 142 849 143
rect 874 143 875 144
rect 879 143 880 147
rect 874 142 880 143
rect 883 147 889 148
rect 883 143 884 147
rect 888 146 889 147
rect 914 147 920 148
rect 914 146 915 147
rect 888 144 915 146
rect 888 143 889 144
rect 883 142 889 143
rect 914 143 915 144
rect 919 143 920 147
rect 914 142 920 143
rect 923 147 929 148
rect 923 143 924 147
rect 928 146 929 147
rect 959 147 965 148
rect 959 146 960 147
rect 928 144 960 146
rect 928 143 929 144
rect 923 142 929 143
rect 959 143 960 144
rect 964 143 965 147
rect 959 142 965 143
rect 971 147 977 148
rect 971 143 972 147
rect 976 146 977 147
rect 1010 147 1016 148
rect 1010 146 1011 147
rect 976 144 1011 146
rect 976 143 977 144
rect 971 142 977 143
rect 1010 143 1011 144
rect 1015 143 1016 147
rect 1010 142 1016 143
rect 1019 147 1025 148
rect 1019 143 1020 147
rect 1024 146 1025 147
rect 1058 147 1064 148
rect 1058 146 1059 147
rect 1024 144 1059 146
rect 1024 143 1025 144
rect 1019 142 1025 143
rect 1058 143 1059 144
rect 1063 143 1064 147
rect 1058 142 1064 143
rect 1067 147 1073 148
rect 1067 143 1068 147
rect 1072 146 1073 147
rect 1098 147 1104 148
rect 1098 146 1099 147
rect 1072 144 1099 146
rect 1072 143 1073 144
rect 1067 142 1073 143
rect 1098 143 1099 144
rect 1103 143 1104 147
rect 1098 142 1104 143
rect 1107 147 1113 148
rect 1107 143 1108 147
rect 1112 146 1113 147
rect 1134 147 1140 148
rect 1134 146 1135 147
rect 1112 144 1135 146
rect 1112 143 1113 144
rect 1107 142 1113 143
rect 1134 143 1135 144
rect 1139 143 1140 147
rect 1134 142 1140 143
rect 1147 147 1153 148
rect 1147 143 1148 147
rect 1152 146 1153 147
rect 1178 147 1184 148
rect 1178 146 1179 147
rect 1152 144 1179 146
rect 1152 143 1153 144
rect 1147 142 1153 143
rect 1178 143 1179 144
rect 1183 143 1184 147
rect 1178 142 1184 143
rect 1187 147 1193 148
rect 1187 143 1188 147
rect 1192 146 1193 147
rect 1294 147 1300 148
rect 1294 146 1295 147
rect 1192 144 1295 146
rect 1192 143 1193 144
rect 1187 142 1193 143
rect 1294 143 1295 144
rect 1299 143 1300 147
rect 1294 142 1300 143
rect 1302 147 1308 148
rect 1302 143 1303 147
rect 1307 143 1308 147
rect 1302 142 1308 143
rect 1342 147 1348 148
rect 1342 143 1343 147
rect 1347 143 1348 147
rect 1342 142 1348 143
rect 1382 147 1388 148
rect 1382 143 1383 147
rect 1387 143 1388 147
rect 1382 142 1388 143
rect 1422 147 1428 148
rect 1422 143 1423 147
rect 1427 143 1428 147
rect 1422 142 1428 143
rect 1462 147 1468 148
rect 1462 143 1463 147
rect 1467 143 1468 147
rect 1462 142 1468 143
rect 1518 147 1524 148
rect 1518 143 1519 147
rect 1523 143 1524 147
rect 1518 142 1524 143
rect 1582 147 1588 148
rect 1582 143 1583 147
rect 1587 143 1588 147
rect 1582 142 1588 143
rect 1646 147 1652 148
rect 1646 143 1647 147
rect 1651 143 1652 147
rect 1646 142 1652 143
rect 1710 147 1716 148
rect 1710 143 1711 147
rect 1715 143 1716 147
rect 1710 142 1716 143
rect 1766 147 1772 148
rect 1766 143 1767 147
rect 1771 143 1772 147
rect 1766 142 1772 143
rect 1822 147 1828 148
rect 1822 143 1823 147
rect 1827 143 1828 147
rect 1822 142 1828 143
rect 1870 147 1876 148
rect 1870 143 1871 147
rect 1875 143 1876 147
rect 1870 142 1876 143
rect 1918 147 1924 148
rect 1918 143 1919 147
rect 1923 143 1924 147
rect 1918 142 1924 143
rect 1966 147 1972 148
rect 1966 143 1967 147
rect 1971 143 1972 147
rect 1966 142 1972 143
rect 2014 147 2020 148
rect 2014 143 2015 147
rect 2019 143 2020 147
rect 2014 142 2020 143
rect 2062 147 2068 148
rect 2062 143 2063 147
rect 2067 143 2068 147
rect 2062 142 2068 143
rect 2110 147 2116 148
rect 2110 143 2111 147
rect 2115 143 2116 147
rect 2110 142 2116 143
rect 2158 147 2164 148
rect 2158 143 2159 147
rect 2163 143 2164 147
rect 2158 142 2164 143
rect 2214 147 2220 148
rect 2214 143 2215 147
rect 2219 143 2220 147
rect 2214 142 2220 143
rect 2270 147 2276 148
rect 2270 143 2271 147
rect 2275 143 2276 147
rect 2270 142 2276 143
rect 2318 147 2324 148
rect 2318 143 2319 147
rect 2323 143 2324 147
rect 2318 142 2324 143
rect 2358 147 2364 148
rect 2358 143 2359 147
rect 2363 143 2364 147
rect 2358 142 2364 143
rect 134 139 140 140
rect 134 135 135 139
rect 139 135 140 139
rect 134 134 140 135
rect 174 139 180 140
rect 174 135 175 139
rect 179 135 180 139
rect 174 134 180 135
rect 214 139 220 140
rect 214 135 215 139
rect 219 135 220 139
rect 214 134 220 135
rect 254 139 260 140
rect 254 135 255 139
rect 259 135 260 139
rect 254 134 260 135
rect 294 139 300 140
rect 294 135 295 139
rect 299 135 300 139
rect 294 134 300 135
rect 334 139 340 140
rect 334 135 335 139
rect 339 135 340 139
rect 334 134 340 135
rect 374 139 380 140
rect 374 135 375 139
rect 379 135 380 139
rect 374 134 380 135
rect 422 139 428 140
rect 422 135 423 139
rect 427 135 428 139
rect 422 134 428 135
rect 470 139 476 140
rect 470 135 471 139
rect 475 135 476 139
rect 470 134 476 135
rect 526 139 532 140
rect 526 135 527 139
rect 531 135 532 139
rect 526 134 532 135
rect 582 139 588 140
rect 582 135 583 139
rect 587 135 588 139
rect 582 134 588 135
rect 630 139 636 140
rect 630 135 631 139
rect 635 135 636 139
rect 630 134 636 135
rect 678 139 684 140
rect 678 135 679 139
rect 683 135 684 139
rect 678 134 684 135
rect 726 139 732 140
rect 726 135 727 139
rect 731 135 732 139
rect 726 134 732 135
rect 766 139 772 140
rect 766 135 767 139
rect 771 135 772 139
rect 766 134 772 135
rect 806 139 812 140
rect 806 135 807 139
rect 811 135 812 139
rect 806 134 812 135
rect 846 139 852 140
rect 846 135 847 139
rect 851 135 852 139
rect 846 134 852 135
rect 886 139 892 140
rect 886 135 887 139
rect 891 135 892 139
rect 886 134 892 135
rect 926 139 932 140
rect 926 135 927 139
rect 931 135 932 139
rect 926 134 932 135
rect 974 139 980 140
rect 974 135 975 139
rect 979 135 980 139
rect 974 134 980 135
rect 1022 139 1028 140
rect 1022 135 1023 139
rect 1027 135 1028 139
rect 1022 134 1028 135
rect 1070 139 1076 140
rect 1070 135 1071 139
rect 1075 135 1076 139
rect 1070 134 1076 135
rect 1110 139 1116 140
rect 1110 135 1111 139
rect 1115 135 1116 139
rect 1110 134 1116 135
rect 1150 139 1156 140
rect 1150 135 1151 139
rect 1155 135 1156 139
rect 1150 134 1156 135
rect 1190 139 1196 140
rect 1190 135 1191 139
rect 1195 135 1196 139
rect 1190 134 1196 135
rect 1502 131 1508 132
rect 1358 127 1364 128
rect 1278 124 1284 125
rect 646 123 652 124
rect 150 119 156 120
rect 110 116 116 117
rect 110 112 111 116
rect 115 112 116 116
rect 150 115 151 119
rect 155 118 156 119
rect 282 119 288 120
rect 155 116 250 118
rect 155 115 156 116
rect 150 114 156 115
rect 110 111 116 112
rect 158 111 165 112
rect 158 107 159 111
rect 164 107 165 111
rect 158 106 165 107
rect 199 111 208 112
rect 199 107 200 111
rect 207 107 208 111
rect 199 106 208 107
rect 238 111 245 112
rect 238 107 239 111
rect 244 107 245 111
rect 248 110 250 116
rect 282 115 283 119
rect 287 118 288 119
rect 318 119 324 120
rect 287 115 290 118
rect 282 114 290 115
rect 318 115 319 119
rect 323 118 324 119
rect 362 119 368 120
rect 323 116 342 118
rect 323 115 324 116
rect 318 114 324 115
rect 279 111 285 112
rect 279 110 280 111
rect 248 108 280 110
rect 238 106 245 107
rect 279 107 280 108
rect 284 107 285 111
rect 288 110 290 114
rect 319 111 325 112
rect 319 110 320 111
rect 288 108 320 110
rect 279 106 285 107
rect 319 107 320 108
rect 324 107 325 111
rect 340 110 342 116
rect 362 115 363 119
rect 367 118 368 119
rect 510 119 516 120
rect 367 115 370 118
rect 362 114 370 115
rect 510 115 511 119
rect 515 118 516 119
rect 646 119 647 123
rect 651 122 652 123
rect 651 120 762 122
rect 1278 120 1279 124
rect 1283 120 1284 124
rect 1358 123 1359 127
rect 1363 126 1364 127
rect 1398 127 1404 128
rect 1363 124 1378 126
rect 1363 123 1364 124
rect 1358 122 1364 123
rect 651 119 652 120
rect 646 118 652 119
rect 515 116 566 118
rect 515 115 516 116
rect 510 114 516 115
rect 359 111 365 112
rect 359 110 360 111
rect 340 108 360 110
rect 319 106 325 107
rect 359 107 360 108
rect 364 107 365 111
rect 368 110 370 114
rect 399 111 405 112
rect 399 110 400 111
rect 368 108 400 110
rect 359 106 365 107
rect 399 107 400 108
rect 404 107 405 111
rect 399 106 405 107
rect 407 111 413 112
rect 407 107 408 111
rect 412 110 413 111
rect 447 111 453 112
rect 447 110 448 111
rect 412 108 448 110
rect 412 107 413 108
rect 407 106 413 107
rect 447 107 448 108
rect 452 107 453 111
rect 447 106 453 107
rect 458 111 464 112
rect 458 107 459 111
rect 463 110 464 111
rect 495 111 501 112
rect 495 110 496 111
rect 463 108 496 110
rect 463 107 464 108
rect 458 106 464 107
rect 495 107 496 108
rect 500 107 501 111
rect 495 106 501 107
rect 551 111 560 112
rect 551 107 552 111
rect 559 107 560 111
rect 564 110 566 116
rect 663 115 669 116
rect 663 114 664 115
rect 655 113 664 114
rect 607 111 613 112
rect 607 110 608 111
rect 564 108 608 110
rect 551 106 560 107
rect 607 107 608 108
rect 612 107 613 111
rect 655 109 656 113
rect 660 112 664 113
rect 660 109 661 112
rect 663 111 664 112
rect 668 111 669 115
rect 663 110 669 111
rect 703 111 712 112
rect 655 108 661 109
rect 607 106 613 107
rect 703 107 704 111
rect 711 107 712 111
rect 703 106 712 107
rect 750 111 757 112
rect 750 107 751 111
rect 756 107 757 111
rect 760 110 762 120
rect 782 119 788 120
rect 782 115 783 119
rect 787 118 788 119
rect 834 119 840 120
rect 787 116 802 118
rect 787 115 788 116
rect 782 114 788 115
rect 791 111 797 112
rect 791 110 792 111
rect 760 108 792 110
rect 750 106 757 107
rect 791 107 792 108
rect 796 107 797 111
rect 800 110 802 116
rect 834 115 835 119
rect 839 118 840 119
rect 874 119 880 120
rect 839 115 842 118
rect 834 114 842 115
rect 874 115 875 119
rect 879 118 880 119
rect 914 119 920 120
rect 879 115 882 118
rect 874 114 882 115
rect 914 115 915 119
rect 919 118 920 119
rect 1098 119 1104 120
rect 919 115 922 118
rect 914 114 922 115
rect 1098 115 1099 119
rect 1103 118 1104 119
rect 1134 119 1140 120
rect 1103 115 1106 118
rect 1098 114 1106 115
rect 1134 115 1135 119
rect 1139 118 1140 119
rect 1178 119 1184 120
rect 1278 119 1284 120
rect 1294 119 1300 120
rect 1139 116 1161 118
rect 1139 115 1140 116
rect 1134 114 1140 115
rect 831 111 837 112
rect 831 110 832 111
rect 800 108 832 110
rect 791 106 797 107
rect 831 107 832 108
rect 836 107 837 111
rect 840 110 842 114
rect 871 111 877 112
rect 871 110 872 111
rect 840 108 872 110
rect 831 106 837 107
rect 871 107 872 108
rect 876 107 877 111
rect 880 110 882 114
rect 911 111 917 112
rect 911 110 912 111
rect 880 108 912 110
rect 871 106 877 107
rect 911 107 912 108
rect 916 107 917 111
rect 920 110 922 114
rect 951 111 957 112
rect 951 110 952 111
rect 920 108 952 110
rect 911 106 917 107
rect 951 107 952 108
rect 956 107 957 111
rect 951 106 957 107
rect 959 111 965 112
rect 959 107 960 111
rect 964 110 965 111
rect 999 111 1005 112
rect 999 110 1000 111
rect 964 108 1000 110
rect 964 107 965 108
rect 959 106 965 107
rect 999 107 1000 108
rect 1004 107 1005 111
rect 999 106 1005 107
rect 1010 111 1016 112
rect 1010 107 1011 111
rect 1015 110 1016 111
rect 1047 111 1053 112
rect 1047 110 1048 111
rect 1015 108 1048 110
rect 1015 107 1016 108
rect 1010 106 1016 107
rect 1047 107 1048 108
rect 1052 107 1053 111
rect 1047 106 1053 107
rect 1058 111 1064 112
rect 1058 107 1059 111
rect 1063 110 1064 111
rect 1095 111 1101 112
rect 1095 110 1096 111
rect 1063 108 1096 110
rect 1063 107 1064 108
rect 1058 106 1064 107
rect 1095 107 1096 108
rect 1100 107 1101 111
rect 1104 110 1106 114
rect 1135 111 1141 112
rect 1135 110 1136 111
rect 1104 108 1136 110
rect 1095 106 1101 107
rect 1135 107 1136 108
rect 1140 107 1141 111
rect 1159 110 1161 116
rect 1178 115 1179 119
rect 1183 118 1184 119
rect 1183 116 1190 118
rect 1183 115 1184 116
rect 1178 114 1184 115
rect 1175 111 1181 112
rect 1175 110 1176 111
rect 1159 108 1176 110
rect 1135 106 1141 107
rect 1175 107 1176 108
rect 1180 107 1181 111
rect 1188 110 1190 116
rect 1238 116 1244 117
rect 1238 112 1239 116
rect 1243 112 1244 116
rect 1294 115 1295 119
rect 1299 118 1300 119
rect 1327 119 1333 120
rect 1327 118 1328 119
rect 1299 116 1328 118
rect 1299 115 1300 116
rect 1294 114 1300 115
rect 1327 115 1328 116
rect 1332 115 1333 119
rect 1327 114 1333 115
rect 1338 119 1344 120
rect 1338 115 1339 119
rect 1343 118 1344 119
rect 1367 119 1373 120
rect 1367 118 1368 119
rect 1343 116 1368 118
rect 1343 115 1344 116
rect 1338 114 1344 115
rect 1367 115 1368 116
rect 1372 115 1373 119
rect 1376 118 1378 124
rect 1398 123 1399 127
rect 1403 126 1404 127
rect 1438 127 1444 128
rect 1403 124 1418 126
rect 1403 123 1404 124
rect 1398 122 1404 123
rect 1407 119 1413 120
rect 1407 118 1408 119
rect 1376 116 1408 118
rect 1367 114 1373 115
rect 1407 115 1408 116
rect 1412 115 1413 119
rect 1416 118 1418 124
rect 1438 123 1439 127
rect 1443 126 1444 127
rect 1502 127 1503 131
rect 1507 130 1508 131
rect 1507 128 1626 130
rect 1507 127 1508 128
rect 1502 126 1508 127
rect 1443 124 1458 126
rect 1443 123 1444 124
rect 1438 122 1444 123
rect 1447 119 1453 120
rect 1447 118 1448 119
rect 1416 116 1448 118
rect 1407 114 1413 115
rect 1447 115 1448 116
rect 1452 115 1453 119
rect 1456 118 1458 124
rect 1615 123 1621 124
rect 1615 122 1616 123
rect 1607 121 1616 122
rect 1487 119 1493 120
rect 1487 118 1488 119
rect 1456 116 1488 118
rect 1447 114 1453 115
rect 1487 115 1488 116
rect 1492 115 1493 119
rect 1487 114 1493 115
rect 1543 119 1549 120
rect 1543 115 1544 119
rect 1548 118 1549 119
rect 1551 119 1557 120
rect 1551 118 1552 119
rect 1548 116 1552 118
rect 1548 115 1549 116
rect 1543 114 1549 115
rect 1551 115 1552 116
rect 1556 115 1557 119
rect 1607 117 1608 121
rect 1612 120 1616 121
rect 1612 117 1613 120
rect 1615 119 1616 120
rect 1620 119 1621 123
rect 1615 118 1621 119
rect 1624 118 1626 128
rect 2346 127 2352 128
rect 1751 123 1757 124
rect 1751 122 1752 123
rect 1735 121 1752 122
rect 1671 119 1677 120
rect 1671 118 1672 119
rect 1607 116 1613 117
rect 1624 116 1672 118
rect 1551 114 1557 115
rect 1671 115 1672 116
rect 1676 115 1677 119
rect 1735 117 1736 121
rect 1740 120 1752 121
rect 1740 117 1741 120
rect 1751 119 1752 120
rect 1756 119 1757 123
rect 2346 123 2347 127
rect 2351 126 2352 127
rect 2351 124 2387 126
rect 2351 123 2352 124
rect 2346 122 2352 123
rect 2385 120 2387 124
rect 2406 124 2412 125
rect 2406 120 2407 124
rect 2411 120 2412 124
rect 1751 118 1757 119
rect 1791 119 1797 120
rect 1735 116 1741 117
rect 1671 114 1677 115
rect 1791 115 1792 119
rect 1796 118 1797 119
rect 1799 119 1805 120
rect 1799 118 1800 119
rect 1796 116 1800 118
rect 1796 115 1797 116
rect 1791 114 1797 115
rect 1799 115 1800 116
rect 1804 115 1805 119
rect 1799 114 1805 115
rect 1847 119 1856 120
rect 1847 115 1848 119
rect 1855 115 1856 119
rect 1847 114 1856 115
rect 1895 119 1904 120
rect 1895 115 1896 119
rect 1903 115 1904 119
rect 1895 114 1904 115
rect 1943 119 1952 120
rect 1943 115 1944 119
rect 1951 115 1952 119
rect 1943 114 1952 115
rect 1991 119 2000 120
rect 1991 115 1992 119
rect 1999 115 2000 119
rect 1991 114 2000 115
rect 2039 119 2048 120
rect 2039 115 2040 119
rect 2047 115 2048 119
rect 2039 114 2048 115
rect 2087 119 2096 120
rect 2087 115 2088 119
rect 2095 115 2096 119
rect 2087 114 2096 115
rect 2135 119 2144 120
rect 2135 115 2136 119
rect 2143 115 2144 119
rect 2135 114 2144 115
rect 2183 119 2192 120
rect 2183 115 2184 119
rect 2191 115 2192 119
rect 2183 114 2192 115
rect 2239 119 2248 120
rect 2239 115 2240 119
rect 2247 115 2248 119
rect 2239 114 2248 115
rect 2306 119 2312 120
rect 2306 115 2307 119
rect 2311 118 2312 119
rect 2343 119 2349 120
rect 2343 118 2344 119
rect 2311 116 2344 118
rect 2311 115 2312 116
rect 2306 114 2312 115
rect 2343 115 2344 116
rect 2348 115 2349 119
rect 2343 114 2349 115
rect 2383 119 2389 120
rect 2406 119 2412 120
rect 2383 115 2384 119
rect 2388 115 2389 119
rect 2383 114 2389 115
rect 1215 111 1221 112
rect 1238 111 1244 112
rect 1215 110 1216 111
rect 1188 108 1216 110
rect 1175 106 1181 107
rect 1215 107 1216 108
rect 1220 107 1221 111
rect 1215 106 1221 107
rect 1278 107 1284 108
rect 1278 103 1279 107
rect 1283 103 1284 107
rect 1278 102 1284 103
rect 2406 107 2412 108
rect 2406 103 2407 107
rect 2411 103 2412 107
rect 2406 102 2412 103
rect 1302 100 1308 101
rect 110 99 116 100
rect 110 95 111 99
rect 115 95 116 99
rect 110 94 116 95
rect 1238 99 1244 100
rect 1238 95 1239 99
rect 1243 95 1244 99
rect 1302 96 1303 100
rect 1307 96 1308 100
rect 1302 95 1308 96
rect 1342 100 1348 101
rect 1342 96 1343 100
rect 1347 96 1348 100
rect 1342 95 1348 96
rect 1382 100 1388 101
rect 1382 96 1383 100
rect 1387 96 1388 100
rect 1382 95 1388 96
rect 1422 100 1428 101
rect 1422 96 1423 100
rect 1427 96 1428 100
rect 1422 95 1428 96
rect 1462 100 1468 101
rect 1462 96 1463 100
rect 1467 96 1468 100
rect 1462 95 1468 96
rect 1518 100 1524 101
rect 1518 96 1519 100
rect 1523 96 1524 100
rect 1518 95 1524 96
rect 1582 100 1588 101
rect 1582 96 1583 100
rect 1587 96 1588 100
rect 1582 95 1588 96
rect 1646 100 1652 101
rect 1646 96 1647 100
rect 1651 96 1652 100
rect 1646 95 1652 96
rect 1710 100 1716 101
rect 1710 96 1711 100
rect 1715 96 1716 100
rect 1710 95 1716 96
rect 1766 100 1772 101
rect 1766 96 1767 100
rect 1771 96 1772 100
rect 1766 95 1772 96
rect 1822 100 1828 101
rect 1822 96 1823 100
rect 1827 96 1828 100
rect 1822 95 1828 96
rect 1870 100 1876 101
rect 1870 96 1871 100
rect 1875 96 1876 100
rect 1870 95 1876 96
rect 1918 100 1924 101
rect 1918 96 1919 100
rect 1923 96 1924 100
rect 1918 95 1924 96
rect 1966 100 1972 101
rect 1966 96 1967 100
rect 1971 96 1972 100
rect 1966 95 1972 96
rect 2014 100 2020 101
rect 2014 96 2015 100
rect 2019 96 2020 100
rect 2014 95 2020 96
rect 2062 100 2068 101
rect 2062 96 2063 100
rect 2067 96 2068 100
rect 2062 95 2068 96
rect 2110 100 2116 101
rect 2110 96 2111 100
rect 2115 96 2116 100
rect 2110 95 2116 96
rect 2158 100 2164 101
rect 2158 96 2159 100
rect 2163 96 2164 100
rect 2158 95 2164 96
rect 2214 100 2220 101
rect 2214 96 2215 100
rect 2219 96 2220 100
rect 2214 95 2220 96
rect 2270 100 2276 101
rect 2270 96 2271 100
rect 2275 96 2276 100
rect 2270 95 2276 96
rect 2318 100 2324 101
rect 2318 96 2319 100
rect 2323 96 2324 100
rect 2318 95 2324 96
rect 2358 100 2364 101
rect 2358 96 2359 100
rect 2363 96 2364 100
rect 2358 95 2364 96
rect 1238 94 1244 95
rect 134 92 140 93
rect 134 88 135 92
rect 139 88 140 92
rect 134 87 140 88
rect 174 92 180 93
rect 174 88 175 92
rect 179 88 180 92
rect 174 87 180 88
rect 214 92 220 93
rect 214 88 215 92
rect 219 88 220 92
rect 214 87 220 88
rect 254 92 260 93
rect 254 88 255 92
rect 259 88 260 92
rect 254 87 260 88
rect 294 92 300 93
rect 294 88 295 92
rect 299 88 300 92
rect 294 87 300 88
rect 334 92 340 93
rect 334 88 335 92
rect 339 88 340 92
rect 334 87 340 88
rect 374 92 380 93
rect 374 88 375 92
rect 379 88 380 92
rect 374 87 380 88
rect 422 92 428 93
rect 422 88 423 92
rect 427 88 428 92
rect 422 87 428 88
rect 470 92 476 93
rect 470 88 471 92
rect 475 88 476 92
rect 470 87 476 88
rect 526 92 532 93
rect 526 88 527 92
rect 531 88 532 92
rect 526 87 532 88
rect 582 92 588 93
rect 582 88 583 92
rect 587 88 588 92
rect 582 87 588 88
rect 630 92 636 93
rect 630 88 631 92
rect 635 88 636 92
rect 630 87 636 88
rect 678 92 684 93
rect 678 88 679 92
rect 683 88 684 92
rect 678 87 684 88
rect 726 92 732 93
rect 726 88 727 92
rect 731 88 732 92
rect 726 87 732 88
rect 766 92 772 93
rect 766 88 767 92
rect 771 88 772 92
rect 766 87 772 88
rect 806 92 812 93
rect 806 88 807 92
rect 811 88 812 92
rect 806 87 812 88
rect 846 92 852 93
rect 846 88 847 92
rect 851 88 852 92
rect 846 87 852 88
rect 886 92 892 93
rect 886 88 887 92
rect 891 88 892 92
rect 886 87 892 88
rect 926 92 932 93
rect 926 88 927 92
rect 931 88 932 92
rect 926 87 932 88
rect 974 92 980 93
rect 974 88 975 92
rect 979 88 980 92
rect 974 87 980 88
rect 1022 92 1028 93
rect 1022 88 1023 92
rect 1027 88 1028 92
rect 1022 87 1028 88
rect 1070 92 1076 93
rect 1070 88 1071 92
rect 1075 88 1076 92
rect 1070 87 1076 88
rect 1110 92 1116 93
rect 1110 88 1111 92
rect 1115 88 1116 92
rect 1110 87 1116 88
rect 1150 92 1156 93
rect 1150 88 1151 92
rect 1155 88 1156 92
rect 1150 87 1156 88
rect 1190 92 1196 93
rect 1190 88 1191 92
rect 1195 88 1196 92
rect 1190 87 1196 88
<< m3c >>
rect 1535 2504 1539 2508
rect 1575 2504 1579 2508
rect 1615 2504 1619 2508
rect 1655 2504 1659 2508
rect 1695 2504 1699 2508
rect 1735 2504 1739 2508
rect 1775 2504 1779 2508
rect 1815 2504 1819 2508
rect 1855 2504 1859 2508
rect 1895 2504 1899 2508
rect 1935 2504 1939 2508
rect 1975 2504 1979 2508
rect 1279 2497 1283 2501
rect 2407 2497 2411 2501
rect 159 2491 163 2495
rect 203 2491 207 2495
rect 243 2491 247 2495
rect 283 2491 287 2495
rect 339 2491 343 2495
rect 419 2491 423 2495
rect 507 2491 511 2495
rect 671 2491 675 2495
rect 683 2491 687 2495
rect 799 2491 803 2495
rect 859 2491 863 2495
rect 135 2483 139 2487
rect 175 2483 179 2487
rect 215 2483 219 2487
rect 255 2483 259 2487
rect 311 2483 315 2487
rect 391 2483 395 2487
rect 479 2483 483 2487
rect 567 2483 571 2487
rect 655 2483 659 2487
rect 743 2483 747 2487
rect 831 2483 835 2487
rect 927 2483 931 2487
rect 1279 2480 1283 2484
rect 1563 2483 1564 2487
rect 1564 2483 1567 2487
rect 1603 2483 1604 2487
rect 1604 2483 1607 2487
rect 1643 2483 1644 2487
rect 1644 2483 1647 2487
rect 1683 2483 1684 2487
rect 1684 2483 1687 2487
rect 1723 2483 1724 2487
rect 1724 2483 1727 2487
rect 1763 2483 1764 2487
rect 1764 2483 1767 2487
rect 1803 2483 1804 2487
rect 1804 2483 1807 2487
rect 1843 2483 1844 2487
rect 1844 2483 1847 2487
rect 1883 2483 1884 2487
rect 1884 2483 1887 2487
rect 1923 2483 1924 2487
rect 1924 2483 1927 2487
rect 1963 2483 1964 2487
rect 1964 2483 1967 2487
rect 1831 2475 1835 2479
rect 2407 2480 2411 2484
rect 111 2460 115 2464
rect 1239 2460 1243 2464
rect 159 2455 160 2459
rect 160 2455 163 2459
rect 203 2455 204 2459
rect 204 2455 207 2459
rect 243 2455 244 2459
rect 244 2455 247 2459
rect 283 2455 284 2459
rect 284 2455 287 2459
rect 339 2455 340 2459
rect 340 2455 343 2459
rect 419 2455 420 2459
rect 420 2455 423 2459
rect 507 2455 508 2459
rect 508 2455 511 2459
rect 111 2443 115 2447
rect 143 2447 147 2451
rect 683 2455 684 2459
rect 684 2455 687 2459
rect 799 2455 803 2459
rect 859 2455 860 2459
rect 860 2455 863 2459
rect 867 2455 871 2459
rect 1535 2457 1539 2461
rect 1575 2457 1579 2461
rect 1615 2457 1619 2461
rect 1655 2457 1659 2461
rect 1695 2457 1699 2461
rect 1735 2457 1739 2461
rect 1775 2457 1779 2461
rect 1815 2457 1819 2461
rect 1855 2457 1859 2461
rect 1895 2457 1899 2461
rect 1935 2457 1939 2461
rect 1975 2457 1979 2461
rect 1239 2443 1243 2447
rect 1555 2447 1559 2451
rect 1563 2447 1567 2451
rect 1603 2451 1607 2455
rect 1643 2447 1647 2451
rect 1683 2451 1687 2455
rect 1723 2447 1727 2451
rect 1763 2451 1767 2455
rect 1803 2447 1807 2451
rect 1843 2451 1847 2455
rect 1883 2447 1887 2451
rect 1923 2451 1927 2455
rect 1963 2447 1967 2451
rect 135 2436 139 2440
rect 175 2436 179 2440
rect 215 2436 219 2440
rect 255 2436 259 2440
rect 311 2436 315 2440
rect 391 2436 395 2440
rect 479 2436 483 2440
rect 567 2436 571 2440
rect 655 2436 659 2440
rect 743 2436 747 2440
rect 831 2436 835 2440
rect 927 2436 931 2440
rect 1379 2435 1383 2439
rect 1387 2435 1391 2439
rect 1427 2435 1431 2439
rect 1483 2435 1487 2439
rect 1547 2435 1551 2439
rect 1627 2435 1631 2439
rect 1707 2435 1711 2439
rect 1831 2435 1835 2439
rect 1867 2435 1871 2439
rect 1947 2435 1951 2439
rect 2027 2435 2031 2439
rect 2107 2435 2111 2439
rect 2183 2435 2187 2439
rect 2291 2435 2295 2439
rect 135 2424 139 2428
rect 183 2424 187 2428
rect 247 2424 251 2428
rect 319 2424 323 2428
rect 391 2424 395 2428
rect 471 2424 475 2428
rect 543 2424 547 2428
rect 615 2424 619 2428
rect 679 2424 683 2428
rect 735 2424 739 2428
rect 791 2424 795 2428
rect 839 2424 843 2428
rect 887 2424 891 2428
rect 935 2424 939 2428
rect 991 2424 995 2428
rect 1047 2424 1051 2428
rect 1359 2427 1363 2431
rect 1399 2427 1403 2431
rect 1455 2427 1459 2431
rect 1519 2427 1523 2431
rect 1599 2427 1603 2431
rect 1679 2427 1683 2431
rect 1759 2427 1763 2431
rect 1839 2427 1843 2431
rect 1919 2427 1923 2431
rect 1999 2427 2003 2431
rect 2079 2427 2083 2431
rect 2159 2427 2163 2431
rect 2247 2427 2251 2431
rect 2335 2427 2339 2431
rect 111 2417 115 2421
rect 1239 2417 1243 2421
rect 671 2411 675 2415
rect 111 2400 115 2404
rect 175 2403 179 2407
rect 239 2403 243 2407
rect 311 2403 315 2407
rect 383 2403 387 2407
rect 463 2403 467 2407
rect 511 2403 515 2407
rect 607 2403 611 2407
rect 671 2403 675 2407
rect 727 2403 731 2407
rect 783 2403 787 2407
rect 879 2403 883 2407
rect 927 2403 931 2407
rect 975 2403 979 2407
rect 1039 2403 1043 2407
rect 1055 2403 1059 2407
rect 1239 2400 1243 2404
rect 1279 2404 1283 2408
rect 1555 2407 1559 2411
rect 1387 2399 1388 2403
rect 1388 2399 1391 2403
rect 1427 2399 1428 2403
rect 1428 2399 1431 2403
rect 1483 2399 1484 2403
rect 1484 2399 1487 2403
rect 1547 2399 1548 2403
rect 1548 2399 1551 2403
rect 1627 2399 1628 2403
rect 1628 2399 1631 2403
rect 1707 2399 1708 2403
rect 1708 2399 1711 2403
rect 2407 2404 2411 2408
rect 1867 2399 1868 2403
rect 1868 2399 1871 2403
rect 1947 2399 1948 2403
rect 1948 2399 1951 2403
rect 2027 2399 2028 2403
rect 2028 2399 2031 2403
rect 2107 2399 2108 2403
rect 2108 2399 2111 2403
rect 2183 2399 2184 2403
rect 2184 2399 2187 2403
rect 2351 2399 2355 2403
rect 1279 2387 1283 2391
rect 2407 2387 2411 2391
rect 135 2377 139 2381
rect 183 2377 187 2381
rect 247 2377 251 2381
rect 319 2377 323 2381
rect 391 2377 395 2381
rect 471 2377 475 2381
rect 543 2377 547 2381
rect 615 2377 619 2381
rect 679 2377 683 2381
rect 735 2377 739 2381
rect 791 2377 795 2381
rect 839 2377 843 2381
rect 887 2377 891 2381
rect 935 2377 939 2381
rect 991 2377 995 2381
rect 1047 2377 1051 2381
rect 1359 2380 1363 2384
rect 1399 2380 1403 2384
rect 1455 2380 1459 2384
rect 1519 2380 1523 2384
rect 1599 2380 1603 2384
rect 1679 2380 1683 2384
rect 1759 2380 1763 2384
rect 1839 2380 1843 2384
rect 1919 2380 1923 2384
rect 1999 2380 2003 2384
rect 2079 2380 2083 2384
rect 2159 2380 2163 2384
rect 2247 2380 2251 2384
rect 2335 2380 2339 2384
rect 143 2367 147 2371
rect 175 2367 179 2371
rect 239 2367 243 2371
rect 311 2367 315 2371
rect 383 2367 387 2371
rect 463 2367 467 2371
rect 591 2367 595 2371
rect 607 2367 611 2371
rect 671 2367 675 2371
rect 727 2367 731 2371
rect 783 2367 787 2371
rect 867 2367 871 2371
rect 879 2367 883 2371
rect 927 2367 931 2371
rect 975 2367 979 2371
rect 1039 2367 1043 2371
rect 1359 2368 1363 2372
rect 1407 2368 1411 2372
rect 1471 2368 1475 2372
rect 1543 2368 1547 2372
rect 1615 2368 1619 2372
rect 1695 2368 1699 2372
rect 1775 2368 1779 2372
rect 1855 2368 1859 2372
rect 1927 2368 1931 2372
rect 1999 2368 2003 2372
rect 2071 2368 2075 2372
rect 2143 2368 2147 2372
rect 2223 2368 2227 2372
rect 2303 2368 2307 2372
rect 2359 2368 2363 2372
rect 1279 2361 1283 2365
rect 2407 2361 2411 2365
rect 1055 2355 1059 2359
rect 155 2347 159 2351
rect 163 2347 167 2351
rect 203 2347 207 2351
rect 419 2347 423 2351
rect 503 2347 507 2351
rect 511 2347 515 2351
rect 667 2347 671 2351
rect 727 2347 731 2351
rect 783 2347 787 2351
rect 851 2347 855 2351
rect 915 2347 919 2351
rect 1279 2344 1283 2348
rect 1379 2347 1383 2351
rect 1687 2347 1691 2351
rect 135 2339 139 2343
rect 175 2339 179 2343
rect 215 2339 219 2343
rect 271 2339 275 2343
rect 351 2339 355 2343
rect 431 2339 435 2343
rect 519 2339 523 2343
rect 599 2339 603 2343
rect 679 2339 683 2343
rect 751 2339 755 2343
rect 823 2339 827 2343
rect 887 2339 891 2343
rect 959 2339 963 2343
rect 1031 2339 1035 2343
rect 1551 2339 1555 2343
rect 1767 2347 1771 2351
rect 2047 2347 2051 2351
rect 2291 2351 2295 2355
rect 2311 2347 2315 2351
rect 2407 2344 2411 2348
rect 111 2316 115 2320
rect 155 2319 159 2323
rect 1359 2321 1363 2325
rect 163 2311 164 2315
rect 164 2311 167 2315
rect 203 2311 204 2315
rect 204 2311 207 2315
rect 111 2299 115 2303
rect 143 2303 147 2307
rect 1407 2321 1411 2325
rect 1471 2321 1475 2325
rect 1543 2321 1547 2325
rect 1615 2321 1619 2325
rect 1695 2321 1699 2325
rect 1775 2321 1779 2325
rect 1855 2321 1859 2325
rect 1927 2321 1931 2325
rect 1999 2321 2003 2325
rect 2071 2321 2075 2325
rect 2143 2321 2147 2325
rect 2223 2321 2227 2325
rect 2303 2321 2307 2325
rect 2359 2321 2363 2325
rect 1239 2316 1243 2320
rect 419 2311 423 2315
rect 503 2311 507 2315
rect 591 2311 595 2315
rect 667 2311 671 2315
rect 727 2311 731 2315
rect 851 2311 852 2315
rect 852 2311 855 2315
rect 915 2311 916 2315
rect 916 2311 919 2315
rect 1003 2311 1007 2315
rect 1551 2311 1555 2315
rect 1607 2311 1611 2315
rect 1687 2311 1691 2315
rect 2047 2311 2051 2315
rect 2231 2311 2235 2315
rect 2351 2311 2355 2315
rect 1239 2299 1243 2303
rect 135 2292 139 2296
rect 175 2292 179 2296
rect 215 2292 219 2296
rect 271 2292 275 2296
rect 351 2292 355 2296
rect 431 2292 435 2296
rect 519 2292 523 2296
rect 599 2292 603 2296
rect 679 2292 683 2296
rect 751 2292 755 2296
rect 823 2292 827 2296
rect 887 2292 891 2296
rect 959 2292 963 2296
rect 1031 2292 1035 2296
rect 1523 2295 1527 2299
rect 1531 2295 1535 2299
rect 1567 2295 1571 2299
rect 1647 2295 1651 2299
rect 1655 2295 1659 2299
rect 1687 2295 1691 2299
rect 1767 2295 1771 2299
rect 1787 2295 1791 2299
rect 2019 2295 2023 2299
rect 2135 2295 2139 2299
rect 2155 2295 2159 2299
rect 2311 2295 2315 2299
rect 2323 2295 2327 2299
rect 1503 2287 1507 2291
rect 1543 2287 1547 2291
rect 1583 2287 1587 2291
rect 1623 2287 1627 2291
rect 1663 2287 1667 2291
rect 1703 2287 1707 2291
rect 1759 2287 1763 2291
rect 1823 2287 1827 2291
rect 1895 2287 1899 2291
rect 1967 2287 1971 2291
rect 2047 2287 2051 2291
rect 2127 2287 2131 2291
rect 2207 2287 2211 2291
rect 2295 2287 2299 2291
rect 2359 2287 2363 2291
rect 135 2276 139 2280
rect 175 2276 179 2280
rect 231 2276 235 2280
rect 303 2276 307 2280
rect 375 2276 379 2280
rect 455 2276 459 2280
rect 535 2276 539 2280
rect 615 2276 619 2280
rect 687 2276 691 2280
rect 759 2276 763 2280
rect 831 2276 835 2280
rect 911 2276 915 2280
rect 991 2276 995 2280
rect 111 2269 115 2273
rect 1239 2269 1243 2273
rect 1279 2264 1283 2268
rect 1523 2267 1527 2271
rect 111 2252 115 2256
rect 163 2255 164 2259
rect 164 2255 167 2259
rect 215 2255 219 2259
rect 295 2255 299 2259
rect 367 2255 371 2259
rect 447 2255 451 2259
rect 255 2247 259 2251
rect 679 2255 683 2259
rect 751 2255 755 2259
rect 783 2255 784 2259
rect 784 2255 787 2259
rect 855 2255 856 2259
rect 856 2255 859 2259
rect 1531 2259 1532 2263
rect 1532 2259 1535 2263
rect 1567 2259 1568 2263
rect 1568 2259 1571 2263
rect 1607 2259 1608 2263
rect 1608 2259 1611 2263
rect 1647 2267 1651 2271
rect 1687 2259 1688 2263
rect 1688 2259 1691 2263
rect 2407 2264 2411 2268
rect 1787 2259 1788 2263
rect 1788 2259 1791 2263
rect 2019 2259 2023 2263
rect 1239 2252 1243 2256
rect 1279 2247 1283 2251
rect 1791 2251 1795 2255
rect 2155 2259 2156 2263
rect 2156 2259 2159 2263
rect 2231 2259 2232 2263
rect 2232 2259 2235 2263
rect 2323 2259 2324 2263
rect 2324 2259 2327 2263
rect 2367 2259 2371 2263
rect 2407 2247 2411 2251
rect 1503 2240 1507 2244
rect 1543 2240 1547 2244
rect 1583 2240 1587 2244
rect 1623 2240 1627 2244
rect 1663 2240 1667 2244
rect 1703 2240 1707 2244
rect 1759 2240 1763 2244
rect 1823 2240 1827 2244
rect 1895 2240 1899 2244
rect 1967 2240 1971 2244
rect 2047 2240 2051 2244
rect 2127 2240 2131 2244
rect 2207 2240 2211 2244
rect 2295 2240 2299 2244
rect 2359 2240 2363 2244
rect 135 2229 139 2233
rect 175 2229 179 2233
rect 231 2229 235 2233
rect 303 2229 307 2233
rect 375 2229 379 2233
rect 455 2229 459 2233
rect 535 2229 539 2233
rect 615 2229 619 2233
rect 687 2229 691 2233
rect 759 2229 763 2233
rect 831 2229 835 2233
rect 911 2229 915 2233
rect 991 2229 995 2233
rect 143 2219 147 2223
rect 163 2219 167 2223
rect 215 2219 219 2223
rect 295 2219 299 2223
rect 367 2219 371 2223
rect 447 2219 451 2223
rect 679 2219 683 2223
rect 751 2219 755 2223
rect 1003 2219 1007 2223
rect 1303 2220 1307 2224
rect 1343 2220 1347 2224
rect 1383 2220 1387 2224
rect 1431 2220 1435 2224
rect 1495 2220 1499 2224
rect 1567 2220 1571 2224
rect 1639 2220 1643 2224
rect 1711 2220 1715 2224
rect 1783 2220 1787 2224
rect 1855 2220 1859 2224
rect 1935 2220 1939 2224
rect 2015 2220 2019 2224
rect 2095 2220 2099 2224
rect 2183 2220 2187 2224
rect 2279 2220 2283 2224
rect 2359 2220 2363 2224
rect 1279 2213 1283 2217
rect 2407 2213 2411 2217
rect 255 2207 259 2211
rect 275 2207 279 2211
rect 315 2207 319 2211
rect 351 2207 355 2211
rect 403 2207 407 2211
rect 463 2207 467 2211
rect 571 2207 575 2211
rect 579 2207 583 2211
rect 635 2207 639 2211
rect 739 2207 743 2211
rect 747 2207 751 2211
rect 855 2207 859 2211
rect 875 2207 879 2211
rect 247 2199 251 2203
rect 287 2199 291 2203
rect 327 2199 331 2203
rect 375 2199 379 2203
rect 431 2199 435 2203
rect 495 2199 499 2203
rect 551 2199 555 2203
rect 607 2199 611 2203
rect 663 2199 667 2203
rect 719 2199 723 2203
rect 783 2199 787 2203
rect 847 2199 851 2203
rect 911 2199 915 2203
rect 1279 2196 1283 2200
rect 1331 2199 1332 2203
rect 1332 2199 1335 2203
rect 1371 2199 1372 2203
rect 1372 2199 1375 2203
rect 1423 2199 1427 2203
rect 1487 2199 1491 2203
rect 1559 2199 1563 2203
rect 1623 2199 1627 2203
rect 1655 2199 1659 2203
rect 1847 2199 1851 2203
rect 1927 2199 1931 2203
rect 2007 2199 2011 2203
rect 2087 2199 2091 2203
rect 1823 2191 1827 2195
rect 2135 2199 2139 2203
rect 2319 2199 2323 2203
rect 2407 2196 2411 2200
rect 111 2176 115 2180
rect 275 2171 276 2175
rect 276 2171 279 2175
rect 315 2171 316 2175
rect 316 2171 319 2175
rect 351 2171 352 2175
rect 352 2171 355 2175
rect 403 2171 404 2175
rect 404 2171 407 2175
rect 459 2171 460 2175
rect 460 2171 463 2175
rect 111 2159 115 2163
rect 391 2163 395 2167
rect 579 2171 580 2175
rect 580 2171 583 2175
rect 635 2171 636 2175
rect 636 2171 639 2175
rect 739 2179 743 2183
rect 747 2171 748 2175
rect 748 2171 751 2175
rect 807 2171 808 2175
rect 808 2171 811 2175
rect 875 2171 876 2175
rect 876 2171 879 2175
rect 1239 2176 1243 2180
rect 1303 2173 1307 2177
rect 1343 2173 1347 2177
rect 1383 2173 1387 2177
rect 1431 2173 1435 2177
rect 1495 2173 1499 2177
rect 1567 2173 1571 2177
rect 1639 2173 1643 2177
rect 1711 2173 1715 2177
rect 1783 2173 1787 2177
rect 1855 2173 1859 2177
rect 1935 2173 1939 2177
rect 2015 2173 2019 2177
rect 2095 2173 2099 2177
rect 2183 2173 2187 2177
rect 2279 2173 2283 2177
rect 2359 2173 2363 2177
rect 1239 2159 1243 2163
rect 1315 2163 1319 2167
rect 1331 2163 1335 2167
rect 1371 2163 1375 2167
rect 1423 2163 1427 2167
rect 1487 2163 1491 2167
rect 1559 2163 1563 2167
rect 1751 2163 1755 2167
rect 1791 2163 1795 2167
rect 1847 2163 1851 2167
rect 1927 2163 1931 2167
rect 2007 2163 2011 2167
rect 2087 2163 2091 2167
rect 2267 2163 2271 2167
rect 2367 2163 2371 2167
rect 247 2152 251 2156
rect 287 2152 291 2156
rect 327 2152 331 2156
rect 375 2152 379 2156
rect 431 2152 435 2156
rect 495 2152 499 2156
rect 551 2152 555 2156
rect 607 2152 611 2156
rect 663 2152 667 2156
rect 719 2152 723 2156
rect 783 2152 787 2156
rect 847 2152 851 2156
rect 911 2152 915 2156
rect 1323 2151 1327 2155
rect 1331 2151 1335 2155
rect 1523 2151 1527 2155
rect 1615 2151 1619 2155
rect 1623 2151 1627 2155
rect 1775 2151 1779 2155
rect 1823 2151 1827 2155
rect 1843 2151 1847 2155
rect 1999 2151 2003 2155
rect 2055 2151 2059 2155
rect 2139 2151 2143 2155
rect 2203 2151 2207 2155
rect 2319 2151 2323 2155
rect 2339 2151 2343 2155
rect 1303 2143 1307 2147
rect 1351 2143 1355 2147
rect 1439 2143 1443 2147
rect 1535 2143 1539 2147
rect 1631 2143 1635 2147
rect 1727 2143 1731 2147
rect 1815 2143 1819 2147
rect 1895 2143 1899 2147
rect 1975 2143 1979 2147
rect 2047 2143 2051 2147
rect 2111 2143 2115 2147
rect 2175 2143 2179 2147
rect 2239 2143 2243 2147
rect 2311 2143 2315 2147
rect 2359 2143 2363 2147
rect 383 2132 387 2136
rect 423 2132 427 2136
rect 463 2132 467 2136
rect 503 2132 507 2136
rect 551 2132 555 2136
rect 607 2132 611 2136
rect 663 2132 667 2136
rect 727 2132 731 2136
rect 791 2132 795 2136
rect 855 2132 859 2136
rect 911 2132 915 2136
rect 967 2132 971 2136
rect 1023 2132 1027 2136
rect 1079 2132 1083 2136
rect 1143 2132 1147 2136
rect 111 2125 115 2129
rect 1239 2125 1243 2129
rect 1279 2120 1283 2124
rect 1315 2123 1319 2127
rect 111 2108 115 2112
rect 411 2111 412 2115
rect 412 2111 415 2115
rect 451 2111 452 2115
rect 452 2111 455 2115
rect 491 2111 492 2115
rect 492 2111 495 2115
rect 399 2103 403 2107
rect 571 2111 575 2115
rect 751 2111 752 2115
rect 752 2111 755 2115
rect 771 2111 775 2115
rect 895 2111 899 2115
rect 951 2111 955 2115
rect 1007 2111 1011 2115
rect 1063 2111 1067 2115
rect 1135 2111 1139 2115
rect 1151 2111 1155 2115
rect 1331 2115 1332 2119
rect 1332 2115 1335 2119
rect 2407 2120 2411 2124
rect 1407 2115 1411 2119
rect 1523 2115 1527 2119
rect 1615 2115 1619 2119
rect 1751 2115 1752 2119
rect 1752 2115 1755 2119
rect 1843 2115 1844 2119
rect 1844 2115 1847 2119
rect 1999 2115 2000 2119
rect 2000 2115 2003 2119
rect 1239 2108 1243 2112
rect 1279 2103 1283 2107
rect 1943 2107 1947 2111
rect 2139 2115 2140 2119
rect 2140 2115 2143 2119
rect 2203 2115 2204 2119
rect 2204 2115 2207 2119
rect 2267 2115 2268 2119
rect 2268 2115 2271 2119
rect 2339 2115 2340 2119
rect 2340 2115 2343 2119
rect 2367 2115 2371 2119
rect 2407 2103 2411 2107
rect 1303 2096 1307 2100
rect 1351 2096 1355 2100
rect 1439 2096 1443 2100
rect 1535 2096 1539 2100
rect 1631 2096 1635 2100
rect 1727 2096 1731 2100
rect 1815 2096 1819 2100
rect 1895 2096 1899 2100
rect 1975 2096 1979 2100
rect 2047 2096 2051 2100
rect 2111 2096 2115 2100
rect 2175 2096 2179 2100
rect 2239 2096 2243 2100
rect 2311 2096 2315 2100
rect 2359 2096 2363 2100
rect 383 2085 387 2089
rect 423 2085 427 2089
rect 463 2085 467 2089
rect 503 2085 507 2089
rect 551 2085 555 2089
rect 607 2085 611 2089
rect 663 2085 667 2089
rect 727 2085 731 2089
rect 791 2085 795 2089
rect 855 2085 859 2089
rect 911 2085 915 2089
rect 967 2085 971 2089
rect 1023 2085 1027 2089
rect 1079 2085 1083 2089
rect 1143 2085 1147 2089
rect 1303 2080 1307 2084
rect 391 2075 395 2079
rect 411 2075 415 2079
rect 451 2075 455 2079
rect 491 2075 495 2079
rect 655 2075 659 2079
rect 771 2075 775 2079
rect 807 2075 811 2079
rect 887 2075 891 2079
rect 895 2075 899 2079
rect 951 2075 955 2079
rect 1007 2075 1011 2079
rect 1063 2075 1067 2079
rect 1343 2080 1347 2084
rect 1399 2080 1403 2084
rect 1479 2080 1483 2084
rect 1567 2080 1571 2084
rect 1663 2080 1667 2084
rect 1759 2080 1763 2084
rect 1847 2080 1851 2084
rect 1935 2080 1939 2084
rect 2015 2080 2019 2084
rect 2095 2080 2099 2084
rect 2167 2080 2171 2084
rect 2239 2080 2243 2084
rect 2311 2080 2315 2084
rect 2359 2080 2363 2084
rect 1135 2075 1139 2079
rect 1279 2073 1283 2077
rect 2407 2073 2411 2077
rect 399 2063 403 2067
rect 411 2063 415 2067
rect 447 2063 451 2067
rect 491 2063 495 2067
rect 527 2063 531 2067
rect 571 2063 575 2067
rect 615 2063 619 2067
rect 751 2063 755 2067
rect 783 2063 787 2067
rect 827 2063 831 2067
rect 875 2063 879 2067
rect 1003 2063 1007 2067
rect 1059 2063 1063 2067
rect 1151 2063 1155 2067
rect 383 2055 387 2059
rect 423 2055 427 2059
rect 463 2055 467 2059
rect 503 2055 507 2059
rect 543 2055 547 2059
rect 583 2055 587 2059
rect 631 2055 635 2059
rect 687 2055 691 2059
rect 743 2055 747 2059
rect 799 2055 803 2059
rect 847 2055 851 2059
rect 903 2055 907 2059
rect 959 2055 963 2059
rect 1015 2055 1019 2059
rect 1071 2055 1075 2059
rect 1279 2056 1283 2060
rect 1323 2059 1327 2063
rect 1339 2059 1343 2063
rect 1471 2059 1475 2063
rect 1547 2059 1551 2063
rect 1655 2059 1659 2063
rect 1671 2059 1675 2063
rect 1775 2059 1779 2063
rect 2007 2059 2011 2063
rect 2055 2059 2059 2063
rect 2159 2059 2163 2063
rect 2183 2059 2187 2063
rect 2103 2051 2107 2055
rect 2275 2059 2279 2063
rect 2407 2056 2411 2060
rect 111 2032 115 2036
rect 1239 2032 1243 2036
rect 1303 2033 1307 2037
rect 1343 2033 1347 2037
rect 1399 2033 1403 2037
rect 1479 2033 1483 2037
rect 1567 2033 1571 2037
rect 1663 2033 1667 2037
rect 1759 2033 1763 2037
rect 1847 2033 1851 2037
rect 1935 2033 1939 2037
rect 2015 2033 2019 2037
rect 2095 2033 2099 2037
rect 2167 2033 2171 2037
rect 2239 2033 2243 2037
rect 2311 2033 2315 2037
rect 2359 2033 2363 2037
rect 411 2027 412 2031
rect 412 2027 415 2031
rect 447 2027 448 2031
rect 448 2027 451 2031
rect 491 2027 492 2031
rect 492 2027 495 2031
rect 527 2027 528 2031
rect 528 2027 531 2031
rect 571 2027 572 2031
rect 572 2027 575 2031
rect 611 2027 612 2031
rect 612 2027 615 2031
rect 655 2027 656 2031
rect 656 2027 659 2031
rect 827 2027 828 2031
rect 828 2027 831 2031
rect 875 2027 876 2031
rect 876 2027 879 2031
rect 887 2027 891 2031
rect 111 2015 115 2019
rect 879 2019 883 2023
rect 1003 2027 1007 2031
rect 1059 2027 1063 2031
rect 1331 2023 1335 2027
rect 1375 2023 1379 2027
rect 1407 2023 1411 2027
rect 1471 2023 1475 2027
rect 1547 2023 1551 2027
rect 1655 2023 1659 2027
rect 1863 2023 1867 2027
rect 1943 2023 1947 2027
rect 2007 2023 2011 2027
rect 2103 2023 2107 2027
rect 2159 2023 2163 2027
rect 2275 2023 2279 2027
rect 2343 2023 2347 2027
rect 2367 2023 2371 2027
rect 1239 2015 1243 2019
rect 383 2008 387 2012
rect 423 2008 427 2012
rect 463 2008 467 2012
rect 503 2008 507 2012
rect 543 2008 547 2012
rect 583 2008 587 2012
rect 631 2008 635 2012
rect 687 2008 691 2012
rect 743 2008 747 2012
rect 799 2008 803 2012
rect 847 2008 851 2012
rect 903 2008 907 2012
rect 959 2008 963 2012
rect 1015 2008 1019 2012
rect 1071 2008 1075 2012
rect 1671 2011 1675 2015
rect 1323 2003 1327 2007
rect 1331 2003 1335 2007
rect 1443 2003 1447 2007
rect 1451 2003 1455 2007
rect 1303 1995 1307 1999
rect 1351 1995 1355 1999
rect 1423 1995 1427 1999
rect 1495 1995 1499 1999
rect 1575 1995 1579 1999
rect 1663 1995 1667 1999
rect 1691 2003 1695 2007
rect 1779 2003 1783 2007
rect 1927 2003 1931 2007
rect 1947 2003 1951 2007
rect 2123 2003 2127 2007
rect 2175 2003 2179 2007
rect 2183 2003 2187 2007
rect 2335 2003 2339 2007
rect 2383 2003 2387 2007
rect 1735 1995 1739 1999
rect 1751 1995 1755 1999
rect 1839 1995 1843 1999
rect 1919 1995 1923 1999
rect 1999 1995 2003 1999
rect 2071 1995 2075 1999
rect 2135 1995 2139 1999
rect 2191 1995 2195 1999
rect 2255 1995 2259 1999
rect 2319 1995 2323 1999
rect 2359 1995 2363 1999
rect 367 1988 371 1992
rect 407 1988 411 1992
rect 455 1988 459 1992
rect 511 1988 515 1992
rect 567 1988 571 1992
rect 631 1988 635 1992
rect 695 1988 699 1992
rect 759 1988 763 1992
rect 815 1988 819 1992
rect 871 1988 875 1992
rect 935 1988 939 1992
rect 999 1988 1003 1992
rect 1063 1988 1067 1992
rect 111 1981 115 1985
rect 1239 1981 1243 1985
rect 1279 1972 1283 1976
rect 1443 1975 1447 1979
rect 111 1964 115 1968
rect 395 1967 396 1971
rect 396 1967 399 1971
rect 447 1967 451 1971
rect 479 1967 480 1971
rect 480 1967 483 1971
rect 375 1959 379 1963
rect 603 1967 607 1971
rect 751 1967 755 1971
rect 783 1967 784 1971
rect 784 1967 787 1971
rect 703 1959 707 1963
rect 927 1967 931 1971
rect 991 1967 995 1971
rect 1055 1967 1059 1971
rect 1071 1967 1075 1971
rect 1239 1964 1243 1968
rect 1331 1967 1332 1971
rect 1332 1967 1335 1971
rect 1375 1967 1376 1971
rect 1376 1967 1379 1971
rect 1451 1967 1452 1971
rect 1452 1967 1455 1971
rect 1523 1967 1524 1971
rect 1524 1967 1527 1971
rect 1927 1975 1931 1979
rect 1691 1967 1692 1971
rect 1692 1967 1695 1971
rect 1779 1967 1780 1971
rect 1780 1967 1783 1971
rect 1863 1967 1864 1971
rect 1864 1967 1867 1971
rect 1947 1967 1948 1971
rect 1948 1967 1951 1971
rect 2335 1975 2339 1979
rect 2407 1972 2411 1976
rect 2123 1967 2127 1971
rect 2175 1967 2179 1971
rect 2231 1967 2235 1971
rect 2343 1967 2344 1971
rect 2344 1967 2347 1971
rect 1279 1955 1283 1959
rect 2407 1955 2411 1959
rect 1303 1948 1307 1952
rect 1351 1948 1355 1952
rect 1423 1948 1427 1952
rect 1495 1948 1499 1952
rect 1575 1948 1579 1952
rect 1663 1948 1667 1952
rect 1751 1948 1755 1952
rect 1839 1948 1843 1952
rect 1919 1948 1923 1952
rect 1999 1948 2003 1952
rect 2071 1948 2075 1952
rect 2135 1948 2139 1952
rect 2191 1948 2195 1952
rect 2255 1948 2259 1952
rect 2319 1948 2323 1952
rect 2359 1948 2363 1952
rect 367 1941 371 1945
rect 407 1941 411 1945
rect 455 1941 459 1945
rect 511 1941 515 1945
rect 567 1941 571 1945
rect 631 1941 635 1945
rect 695 1941 699 1945
rect 759 1941 763 1945
rect 815 1941 819 1945
rect 871 1941 875 1945
rect 935 1941 939 1945
rect 999 1941 1003 1945
rect 1063 1941 1067 1945
rect 1303 1936 1307 1940
rect 375 1931 379 1935
rect 395 1931 399 1935
rect 447 1931 451 1935
rect 603 1931 607 1935
rect 703 1931 707 1935
rect 751 1931 755 1935
rect 823 1931 827 1935
rect 879 1931 883 1935
rect 927 1931 931 1935
rect 991 1931 995 1935
rect 1359 1936 1363 1940
rect 1447 1936 1451 1940
rect 1535 1936 1539 1940
rect 1623 1936 1627 1940
rect 1711 1936 1715 1940
rect 1791 1936 1795 1940
rect 1863 1936 1867 1940
rect 1935 1936 1939 1940
rect 2007 1936 2011 1940
rect 2079 1936 2083 1940
rect 2151 1936 2155 1940
rect 2223 1936 2227 1940
rect 2303 1936 2307 1940
rect 2359 1936 2363 1940
rect 1055 1931 1059 1935
rect 1279 1929 1283 1933
rect 2407 1929 2411 1933
rect 1071 1923 1075 1927
rect 191 1915 195 1919
rect 199 1915 203 1919
rect 379 1915 383 1919
rect 479 1915 483 1919
rect 499 1915 503 1919
rect 655 1915 659 1919
rect 747 1915 751 1919
rect 903 1915 907 1919
rect 987 1915 991 1919
rect 1071 1915 1075 1919
rect 1279 1912 1283 1916
rect 1323 1915 1327 1919
rect 1703 1915 1707 1919
rect 1735 1915 1736 1919
rect 1736 1915 1739 1919
rect 1855 1915 1859 1919
rect 1927 1915 1931 1919
rect 1963 1915 1964 1919
rect 1964 1915 1967 1919
rect 175 1907 179 1911
rect 215 1907 219 1911
rect 263 1907 267 1911
rect 319 1907 323 1911
rect 391 1907 395 1911
rect 471 1907 475 1911
rect 551 1907 555 1911
rect 639 1907 643 1911
rect 719 1907 723 1911
rect 799 1907 803 1911
rect 879 1907 883 1911
rect 959 1907 963 1911
rect 1039 1907 1043 1911
rect 1119 1907 1123 1911
rect 1799 1907 1803 1911
rect 2143 1915 2147 1919
rect 2015 1907 2019 1911
rect 2295 1915 2299 1919
rect 2351 1915 2355 1919
rect 2383 1915 2384 1919
rect 2384 1915 2387 1919
rect 2407 1912 2411 1916
rect 111 1884 115 1888
rect 191 1887 195 1891
rect 1303 1889 1307 1893
rect 199 1879 200 1883
rect 200 1879 203 1883
rect 335 1879 339 1883
rect 379 1879 383 1883
rect 499 1879 500 1883
rect 500 1879 503 1883
rect 1359 1889 1363 1893
rect 1447 1889 1451 1893
rect 1535 1889 1539 1893
rect 1623 1889 1627 1893
rect 1711 1889 1715 1893
rect 1791 1889 1795 1893
rect 1863 1889 1867 1893
rect 1935 1889 1939 1893
rect 2007 1889 2011 1893
rect 2079 1889 2083 1893
rect 2151 1889 2155 1893
rect 2223 1889 2227 1893
rect 2303 1889 2307 1893
rect 2359 1889 2363 1893
rect 1239 1884 1243 1888
rect 747 1879 748 1883
rect 748 1879 751 1883
rect 823 1879 824 1883
rect 824 1879 827 1883
rect 903 1879 904 1883
rect 904 1879 907 1883
rect 987 1879 988 1883
rect 988 1879 991 1883
rect 1067 1879 1068 1883
rect 1068 1879 1071 1883
rect 111 1867 115 1871
rect 919 1871 923 1875
rect 1439 1879 1443 1883
rect 1523 1879 1527 1883
rect 1703 1879 1707 1883
rect 1799 1879 1803 1883
rect 1855 1879 1859 1883
rect 1927 1879 1931 1883
rect 2015 1879 2019 1883
rect 2143 1879 2147 1883
rect 2231 1879 2235 1883
rect 2295 1879 2299 1883
rect 2383 1879 2387 1883
rect 1239 1867 1243 1871
rect 1331 1867 1335 1871
rect 1339 1867 1343 1871
rect 1387 1867 1391 1871
rect 1599 1867 1603 1871
rect 1607 1867 1611 1871
rect 1755 1867 1759 1871
rect 1851 1867 1855 1871
rect 1963 1867 1967 1871
rect 2123 1867 2127 1871
rect 2351 1867 2355 1871
rect 175 1860 179 1864
rect 215 1860 219 1864
rect 263 1860 267 1864
rect 319 1860 323 1864
rect 391 1860 395 1864
rect 471 1860 475 1864
rect 551 1860 555 1864
rect 639 1860 643 1864
rect 719 1860 723 1864
rect 799 1860 803 1864
rect 879 1860 883 1864
rect 959 1860 963 1864
rect 1039 1860 1043 1864
rect 1119 1860 1123 1864
rect 1311 1859 1315 1863
rect 1359 1859 1363 1863
rect 1415 1859 1419 1863
rect 1479 1859 1483 1863
rect 1543 1859 1547 1863
rect 1615 1859 1619 1863
rect 1687 1859 1691 1863
rect 1767 1859 1771 1863
rect 1863 1859 1867 1863
rect 1975 1859 1979 1863
rect 2095 1859 2099 1863
rect 2223 1859 2227 1863
rect 2359 1859 2363 1863
rect 135 1840 139 1844
rect 175 1840 179 1844
rect 215 1840 219 1844
rect 271 1840 275 1844
rect 351 1840 355 1844
rect 439 1840 443 1844
rect 535 1840 539 1844
rect 631 1840 635 1844
rect 727 1840 731 1844
rect 823 1840 827 1844
rect 911 1840 915 1844
rect 991 1840 995 1844
rect 1063 1840 1067 1844
rect 1135 1840 1139 1844
rect 1191 1840 1195 1844
rect 111 1833 115 1837
rect 1239 1833 1243 1837
rect 1279 1836 1283 1840
rect 1331 1839 1335 1843
rect 1339 1831 1340 1835
rect 1340 1831 1343 1835
rect 1387 1831 1388 1835
rect 1388 1831 1391 1835
rect 1439 1831 1440 1835
rect 1440 1831 1443 1835
rect 1599 1831 1603 1835
rect 1671 1831 1675 1835
rect 1755 1831 1759 1835
rect 1851 1831 1855 1835
rect 2123 1831 2124 1835
rect 2124 1831 2127 1835
rect 2407 1836 2411 1840
rect 2383 1831 2384 1835
rect 2384 1831 2387 1835
rect 111 1816 115 1820
rect 143 1819 147 1823
rect 151 1811 155 1815
rect 183 1811 187 1815
rect 431 1819 435 1823
rect 527 1819 531 1823
rect 295 1811 299 1815
rect 655 1819 656 1823
rect 656 1819 659 1823
rect 983 1819 987 1823
rect 1055 1819 1059 1823
rect 1127 1819 1131 1823
rect 1183 1819 1187 1823
rect 1039 1811 1043 1815
rect 1239 1816 1243 1820
rect 1279 1819 1283 1823
rect 2407 1819 2411 1823
rect 1311 1812 1315 1816
rect 1359 1812 1363 1816
rect 1415 1812 1419 1816
rect 1479 1812 1483 1816
rect 1543 1812 1547 1816
rect 1615 1812 1619 1816
rect 1687 1812 1691 1816
rect 1767 1812 1771 1816
rect 1863 1812 1867 1816
rect 1975 1812 1979 1816
rect 2095 1812 2099 1816
rect 2223 1812 2227 1816
rect 2359 1812 2363 1816
rect 135 1793 139 1797
rect 175 1793 179 1797
rect 215 1793 219 1797
rect 271 1793 275 1797
rect 351 1793 355 1797
rect 439 1793 443 1797
rect 535 1793 539 1797
rect 631 1793 635 1797
rect 727 1793 731 1797
rect 823 1793 827 1797
rect 911 1793 915 1797
rect 991 1793 995 1797
rect 1063 1793 1067 1797
rect 1135 1793 1139 1797
rect 1191 1793 1195 1797
rect 1407 1796 1411 1800
rect 1471 1796 1475 1800
rect 1535 1796 1539 1800
rect 1599 1796 1603 1800
rect 1663 1796 1667 1800
rect 1727 1796 1731 1800
rect 1783 1796 1787 1800
rect 1839 1796 1843 1800
rect 1895 1796 1899 1800
rect 1959 1796 1963 1800
rect 1279 1789 1283 1793
rect 2407 1789 2411 1793
rect 151 1783 155 1787
rect 183 1783 187 1787
rect 295 1783 299 1787
rect 335 1783 339 1787
rect 431 1783 435 1787
rect 527 1783 531 1787
rect 779 1783 783 1787
rect 919 1783 923 1787
rect 983 1783 987 1787
rect 1055 1783 1059 1787
rect 1127 1783 1131 1787
rect 1183 1783 1187 1787
rect 143 1771 147 1775
rect 159 1771 163 1775
rect 199 1771 203 1775
rect 243 1771 247 1775
rect 315 1771 319 1775
rect 403 1771 407 1775
rect 499 1771 503 1775
rect 683 1771 687 1775
rect 691 1771 695 1775
rect 891 1771 895 1775
rect 955 1771 959 1775
rect 1007 1771 1011 1775
rect 1039 1771 1043 1775
rect 1115 1771 1119 1775
rect 1175 1771 1179 1775
rect 1279 1772 1283 1776
rect 1463 1775 1467 1779
rect 1527 1775 1531 1779
rect 1591 1775 1595 1779
rect 1607 1775 1611 1779
rect 1719 1775 1723 1779
rect 1775 1775 1779 1779
rect 1831 1775 1835 1779
rect 1887 1775 1891 1779
rect 1951 1775 1955 1779
rect 135 1763 139 1767
rect 175 1763 179 1767
rect 215 1763 219 1767
rect 287 1763 291 1767
rect 375 1763 379 1767
rect 471 1763 475 1767
rect 567 1763 571 1767
rect 663 1763 667 1767
rect 751 1763 755 1767
rect 831 1763 835 1767
rect 903 1763 907 1767
rect 967 1763 971 1767
rect 1031 1763 1035 1767
rect 1087 1763 1091 1767
rect 1151 1763 1155 1767
rect 1191 1763 1195 1767
rect 1743 1767 1747 1771
rect 2407 1772 2411 1776
rect 1407 1749 1411 1753
rect 1471 1749 1475 1753
rect 1535 1749 1539 1753
rect 1599 1749 1603 1753
rect 1663 1749 1667 1753
rect 1727 1749 1731 1753
rect 1783 1749 1787 1753
rect 1839 1749 1843 1753
rect 1895 1749 1899 1753
rect 1959 1749 1963 1753
rect 111 1740 115 1744
rect 683 1743 687 1747
rect 159 1735 160 1739
rect 160 1735 163 1739
rect 199 1735 200 1739
rect 200 1735 203 1739
rect 243 1735 244 1739
rect 244 1735 247 1739
rect 315 1735 316 1739
rect 316 1735 319 1739
rect 403 1735 404 1739
rect 404 1735 407 1739
rect 499 1735 500 1739
rect 500 1735 503 1739
rect 111 1723 115 1727
rect 143 1727 147 1731
rect 691 1735 692 1739
rect 692 1735 695 1739
rect 779 1735 780 1739
rect 780 1735 783 1739
rect 1239 1740 1243 1744
rect 891 1735 895 1739
rect 955 1735 959 1739
rect 1115 1735 1116 1739
rect 1116 1735 1119 1739
rect 1175 1735 1176 1739
rect 1176 1735 1179 1739
rect 1447 1739 1451 1743
rect 1463 1739 1467 1743
rect 1527 1739 1531 1743
rect 1591 1739 1595 1743
rect 1671 1739 1675 1743
rect 1719 1739 1723 1743
rect 1775 1739 1779 1743
rect 1831 1739 1835 1743
rect 1887 1739 1891 1743
rect 1951 1739 1955 1743
rect 1239 1723 1243 1727
rect 1331 1727 1335 1731
rect 1487 1727 1491 1731
rect 1571 1727 1575 1731
rect 1651 1727 1655 1731
rect 1743 1727 1747 1731
rect 1763 1727 1767 1731
rect 1919 1727 1923 1731
rect 1967 1727 1971 1731
rect 2027 1727 2031 1731
rect 135 1716 139 1720
rect 175 1716 179 1720
rect 215 1716 219 1720
rect 287 1716 291 1720
rect 375 1716 379 1720
rect 471 1716 475 1720
rect 567 1716 571 1720
rect 663 1716 667 1720
rect 751 1716 755 1720
rect 831 1716 835 1720
rect 903 1716 907 1720
rect 967 1716 971 1720
rect 1031 1716 1035 1720
rect 1087 1716 1091 1720
rect 1151 1716 1155 1720
rect 1191 1716 1195 1720
rect 1303 1719 1307 1723
rect 1351 1719 1355 1723
rect 1423 1719 1427 1723
rect 1503 1719 1507 1723
rect 1583 1719 1587 1723
rect 1663 1719 1667 1723
rect 1735 1719 1739 1723
rect 1807 1719 1811 1723
rect 1871 1719 1875 1723
rect 1935 1719 1939 1723
rect 1999 1719 2003 1723
rect 2063 1719 2067 1723
rect 135 1700 139 1704
rect 175 1700 179 1704
rect 239 1700 243 1704
rect 319 1700 323 1704
rect 415 1700 419 1704
rect 511 1700 515 1704
rect 615 1700 619 1704
rect 711 1700 715 1704
rect 799 1700 803 1704
rect 879 1700 883 1704
rect 951 1700 955 1704
rect 1015 1700 1019 1704
rect 1087 1700 1091 1704
rect 1159 1700 1163 1704
rect 111 1693 115 1697
rect 1239 1693 1243 1697
rect 1279 1696 1283 1700
rect 1007 1687 1011 1691
rect 1331 1691 1332 1695
rect 1332 1691 1335 1695
rect 1339 1691 1343 1695
rect 1447 1691 1448 1695
rect 1448 1691 1451 1695
rect 1487 1691 1491 1695
rect 1571 1691 1575 1695
rect 1651 1691 1655 1695
rect 1763 1691 1764 1695
rect 1764 1691 1767 1695
rect 1919 1695 1923 1699
rect 2407 1696 2411 1700
rect 1963 1691 1964 1695
rect 1964 1691 1967 1695
rect 2027 1691 2028 1695
rect 2028 1691 2031 1695
rect 111 1676 115 1680
rect 163 1679 164 1683
rect 164 1679 167 1683
rect 231 1679 235 1683
rect 311 1679 315 1683
rect 407 1679 411 1683
rect 503 1679 507 1683
rect 607 1679 611 1683
rect 623 1679 627 1683
rect 791 1679 795 1683
rect 871 1679 875 1683
rect 943 1679 947 1683
rect 1007 1679 1011 1683
rect 1079 1679 1083 1683
rect 1151 1679 1155 1683
rect 1239 1676 1243 1680
rect 1279 1679 1283 1683
rect 1823 1683 1827 1687
rect 2407 1679 2411 1683
rect 1303 1672 1307 1676
rect 1351 1672 1355 1676
rect 1423 1672 1427 1676
rect 1503 1672 1507 1676
rect 1583 1672 1587 1676
rect 1663 1672 1667 1676
rect 1735 1672 1739 1676
rect 1807 1672 1811 1676
rect 1871 1672 1875 1676
rect 1935 1672 1939 1676
rect 1999 1672 2003 1676
rect 2063 1672 2067 1676
rect 1303 1660 1307 1664
rect 1359 1660 1363 1664
rect 1447 1660 1451 1664
rect 1543 1660 1547 1664
rect 1639 1660 1643 1664
rect 1727 1660 1731 1664
rect 1815 1660 1819 1664
rect 1895 1660 1899 1664
rect 1967 1660 1971 1664
rect 2031 1660 2035 1664
rect 2095 1660 2099 1664
rect 2159 1660 2163 1664
rect 2223 1660 2227 1664
rect 135 1653 139 1657
rect 175 1653 179 1657
rect 239 1653 243 1657
rect 319 1653 323 1657
rect 415 1653 419 1657
rect 511 1653 515 1657
rect 615 1653 619 1657
rect 711 1653 715 1657
rect 799 1653 803 1657
rect 879 1653 883 1657
rect 951 1653 955 1657
rect 1015 1653 1019 1657
rect 1087 1653 1091 1657
rect 1159 1653 1163 1657
rect 1279 1653 1283 1657
rect 2407 1653 2411 1657
rect 143 1643 147 1647
rect 163 1643 167 1647
rect 231 1643 235 1647
rect 311 1643 315 1647
rect 407 1643 411 1647
rect 503 1643 507 1647
rect 607 1643 611 1647
rect 767 1635 771 1639
rect 791 1643 795 1647
rect 871 1643 875 1647
rect 943 1643 947 1647
rect 1007 1643 1011 1647
rect 1079 1643 1083 1647
rect 1151 1643 1155 1647
rect 1023 1635 1027 1639
rect 1279 1636 1283 1640
rect 1351 1639 1355 1643
rect 1439 1639 1443 1643
rect 1455 1639 1459 1643
rect 1631 1639 1635 1643
rect 1719 1639 1723 1643
rect 1887 1639 1891 1643
rect 1959 1639 1963 1643
rect 2023 1639 2027 1643
rect 2087 1639 2091 1643
rect 2151 1639 2155 1643
rect 2207 1639 2211 1643
rect 279 1627 283 1631
rect 299 1627 303 1631
rect 339 1627 343 1631
rect 395 1627 399 1631
rect 443 1627 447 1631
rect 499 1627 503 1631
rect 563 1627 567 1631
rect 691 1627 695 1631
rect 747 1627 751 1631
rect 811 1627 815 1631
rect 859 1627 863 1631
rect 915 1627 919 1631
rect 971 1627 975 1631
rect 1919 1631 1923 1635
rect 2407 1636 2411 1640
rect 271 1619 275 1623
rect 311 1619 315 1623
rect 359 1619 363 1623
rect 415 1619 419 1623
rect 471 1619 475 1623
rect 535 1619 539 1623
rect 599 1619 603 1623
rect 663 1619 667 1623
rect 719 1619 723 1623
rect 775 1619 779 1623
rect 831 1619 835 1623
rect 887 1619 891 1623
rect 943 1619 947 1623
rect 999 1619 1003 1623
rect 1303 1613 1307 1617
rect 1359 1613 1363 1617
rect 1447 1613 1451 1617
rect 1543 1613 1547 1617
rect 1639 1613 1643 1617
rect 1727 1613 1731 1617
rect 1815 1613 1819 1617
rect 1895 1613 1899 1617
rect 1967 1613 1971 1617
rect 2031 1613 2035 1617
rect 2095 1613 2099 1617
rect 2159 1613 2163 1617
rect 2223 1613 2227 1617
rect 1339 1603 1343 1607
rect 1351 1603 1355 1607
rect 1439 1603 1443 1607
rect 1507 1603 1511 1607
rect 1631 1603 1635 1607
rect 1719 1603 1723 1607
rect 1823 1603 1827 1607
rect 1887 1603 1891 1607
rect 1959 1603 1963 1607
rect 2023 1603 2027 1607
rect 2087 1603 2091 1607
rect 2151 1603 2155 1607
rect 2207 1603 2211 1607
rect 111 1596 115 1600
rect 1239 1596 1243 1600
rect 299 1591 300 1595
rect 300 1591 303 1595
rect 339 1591 340 1595
rect 340 1591 343 1595
rect 395 1591 399 1595
rect 443 1591 444 1595
rect 444 1591 447 1595
rect 499 1591 500 1595
rect 500 1591 503 1595
rect 563 1591 564 1595
rect 564 1591 567 1595
rect 691 1591 692 1595
rect 692 1591 695 1595
rect 747 1591 748 1595
rect 748 1591 751 1595
rect 811 1591 815 1595
rect 859 1591 860 1595
rect 860 1591 863 1595
rect 915 1591 916 1595
rect 916 1591 919 1595
rect 971 1591 972 1595
rect 972 1591 975 1595
rect 1023 1591 1024 1595
rect 1024 1591 1027 1595
rect 1383 1591 1387 1595
rect 1455 1591 1459 1595
rect 1555 1591 1559 1595
rect 1719 1591 1723 1595
rect 1919 1591 1923 1595
rect 1939 1591 1943 1595
rect 2011 1591 2015 1595
rect 2075 1591 2079 1595
rect 2151 1591 2155 1595
rect 2195 1591 2199 1595
rect 2243 1591 2247 1595
rect 2299 1591 2303 1595
rect 2347 1591 2351 1595
rect 111 1579 115 1583
rect 347 1583 351 1587
rect 767 1583 771 1587
rect 951 1583 955 1587
rect 1239 1579 1243 1583
rect 1327 1583 1331 1587
rect 1399 1583 1403 1587
rect 1479 1583 1483 1587
rect 1567 1583 1571 1587
rect 1655 1583 1659 1587
rect 1743 1583 1747 1587
rect 1831 1583 1835 1587
rect 1911 1583 1915 1587
rect 1983 1583 1987 1587
rect 2047 1583 2051 1587
rect 2111 1583 2115 1587
rect 2167 1583 2171 1587
rect 2215 1583 2219 1587
rect 2271 1583 2275 1587
rect 2319 1583 2323 1587
rect 2359 1583 2363 1587
rect 271 1572 275 1576
rect 311 1572 315 1576
rect 359 1572 363 1576
rect 415 1572 419 1576
rect 471 1572 475 1576
rect 535 1572 539 1576
rect 599 1572 603 1576
rect 663 1572 667 1576
rect 719 1572 723 1576
rect 775 1572 779 1576
rect 831 1572 835 1576
rect 887 1572 891 1576
rect 943 1572 947 1576
rect 999 1572 1003 1576
rect 1279 1560 1283 1564
rect 2407 1560 2411 1564
rect 327 1552 331 1556
rect 367 1552 371 1556
rect 407 1552 411 1556
rect 447 1552 451 1556
rect 487 1552 491 1556
rect 527 1552 531 1556
rect 567 1552 571 1556
rect 607 1552 611 1556
rect 647 1552 651 1556
rect 687 1552 691 1556
rect 727 1552 731 1556
rect 767 1552 771 1556
rect 807 1552 811 1556
rect 847 1552 851 1556
rect 887 1552 891 1556
rect 927 1552 931 1556
rect 1343 1555 1347 1559
rect 1383 1555 1387 1559
rect 1507 1555 1508 1559
rect 1508 1555 1511 1559
rect 1555 1555 1559 1559
rect 1719 1555 1723 1559
rect 1939 1555 1940 1559
rect 1940 1555 1943 1559
rect 2011 1555 2012 1559
rect 2012 1555 2015 1559
rect 2075 1555 2076 1559
rect 2076 1555 2079 1559
rect 2151 1555 2155 1559
rect 2195 1555 2196 1559
rect 2196 1555 2199 1559
rect 2243 1555 2244 1559
rect 2244 1555 2247 1559
rect 2299 1555 2300 1559
rect 2300 1555 2303 1559
rect 2347 1555 2348 1559
rect 2348 1555 2351 1559
rect 111 1545 115 1549
rect 1239 1545 1243 1549
rect 1279 1543 1283 1547
rect 2223 1547 2227 1551
rect 2407 1543 2411 1547
rect 1327 1536 1331 1540
rect 111 1528 115 1532
rect 355 1531 356 1535
rect 356 1531 359 1535
rect 395 1531 396 1535
rect 396 1531 399 1535
rect 435 1531 436 1535
rect 436 1531 439 1535
rect 475 1531 476 1535
rect 476 1531 479 1535
rect 515 1531 516 1535
rect 516 1531 519 1535
rect 555 1531 556 1535
rect 556 1531 559 1535
rect 595 1531 596 1535
rect 596 1531 599 1535
rect 635 1531 636 1535
rect 636 1531 639 1535
rect 675 1531 676 1535
rect 676 1531 679 1535
rect 715 1531 716 1535
rect 716 1531 719 1535
rect 755 1531 756 1535
rect 756 1531 759 1535
rect 795 1531 796 1535
rect 796 1531 799 1535
rect 835 1531 836 1535
rect 836 1531 839 1535
rect 875 1531 876 1535
rect 876 1531 879 1535
rect 915 1531 916 1535
rect 916 1531 919 1535
rect 1399 1536 1403 1540
rect 1479 1536 1483 1540
rect 1567 1536 1571 1540
rect 1655 1536 1659 1540
rect 1743 1536 1747 1540
rect 1831 1536 1835 1540
rect 1911 1536 1915 1540
rect 1983 1536 1987 1540
rect 2047 1536 2051 1540
rect 2111 1536 2115 1540
rect 2167 1536 2171 1540
rect 2215 1536 2219 1540
rect 2271 1536 2275 1540
rect 2319 1536 2323 1540
rect 2359 1536 2363 1540
rect 951 1531 952 1535
rect 952 1531 955 1535
rect 1239 1528 1243 1532
rect 1335 1520 1339 1524
rect 1415 1520 1419 1524
rect 1503 1520 1507 1524
rect 1615 1520 1619 1524
rect 1743 1520 1747 1524
rect 1887 1520 1891 1524
rect 2047 1520 2051 1524
rect 2215 1520 2219 1524
rect 2359 1520 2363 1524
rect 1279 1513 1283 1517
rect 2407 1513 2411 1517
rect 327 1505 331 1509
rect 367 1505 371 1509
rect 407 1505 411 1509
rect 447 1505 451 1509
rect 487 1505 491 1509
rect 527 1505 531 1509
rect 567 1505 571 1509
rect 607 1505 611 1509
rect 647 1505 651 1509
rect 687 1505 691 1509
rect 727 1505 731 1509
rect 767 1505 771 1509
rect 807 1505 811 1509
rect 847 1505 851 1509
rect 887 1505 891 1509
rect 927 1505 931 1509
rect 347 1495 351 1499
rect 355 1495 359 1499
rect 395 1495 399 1499
rect 435 1495 439 1499
rect 475 1495 479 1499
rect 515 1495 519 1499
rect 555 1495 559 1499
rect 595 1495 599 1499
rect 635 1495 639 1499
rect 675 1495 679 1499
rect 715 1495 719 1499
rect 755 1495 759 1499
rect 795 1495 799 1499
rect 835 1495 839 1499
rect 875 1495 879 1499
rect 915 1495 919 1499
rect 1279 1496 1283 1500
rect 1407 1499 1411 1503
rect 1487 1499 1491 1503
rect 1495 1499 1499 1503
rect 1735 1499 1739 1503
rect 2039 1499 2043 1503
rect 2351 1499 2355 1503
rect 2367 1499 2371 1503
rect 2407 1496 2411 1500
rect 1335 1473 1339 1477
rect 1415 1473 1419 1477
rect 1503 1473 1507 1477
rect 1615 1473 1619 1477
rect 1743 1473 1747 1477
rect 1887 1473 1891 1477
rect 2047 1473 2051 1477
rect 2215 1473 2219 1477
rect 2359 1473 2363 1477
rect 1343 1463 1347 1467
rect 1407 1463 1411 1467
rect 1487 1463 1491 1467
rect 1719 1463 1723 1467
rect 1735 1463 1739 1467
rect 2039 1463 2043 1467
rect 2223 1463 2227 1467
rect 2351 1463 2355 1467
rect 1451 1451 1455 1455
rect 1495 1451 1499 1455
rect 1559 1451 1563 1455
rect 1579 1451 1583 1455
rect 1667 1451 1671 1455
rect 1827 1451 1831 1455
rect 1835 1451 1839 1455
rect 1907 1451 1911 1455
rect 2035 1451 2039 1455
rect 2083 1451 2087 1455
rect 2131 1451 2135 1455
rect 2179 1451 2183 1455
rect 2227 1451 2231 1455
rect 2267 1451 2271 1455
rect 2303 1451 2307 1455
rect 2311 1451 2315 1455
rect 2367 1451 2371 1455
rect 159 1443 163 1447
rect 167 1443 171 1447
rect 207 1443 211 1447
rect 251 1443 255 1447
rect 347 1443 351 1447
rect 419 1443 423 1447
rect 499 1443 503 1447
rect 587 1443 591 1447
rect 743 1443 747 1447
rect 755 1443 759 1447
rect 835 1443 839 1447
rect 907 1443 911 1447
rect 971 1443 975 1447
rect 1027 1443 1031 1447
rect 1075 1443 1079 1447
rect 1139 1443 1143 1447
rect 1175 1443 1179 1447
rect 1375 1443 1379 1447
rect 1463 1443 1467 1447
rect 1551 1443 1555 1447
rect 1639 1443 1643 1447
rect 1727 1443 1731 1447
rect 1807 1443 1811 1447
rect 1879 1443 1883 1447
rect 1943 1443 1947 1447
rect 1999 1443 2003 1447
rect 2047 1443 2051 1447
rect 2095 1443 2099 1447
rect 2143 1443 2147 1447
rect 2191 1443 2195 1447
rect 2239 1443 2243 1447
rect 2279 1443 2283 1447
rect 2319 1443 2323 1447
rect 2359 1443 2363 1447
rect 143 1435 147 1439
rect 183 1435 187 1439
rect 223 1435 227 1439
rect 263 1435 267 1439
rect 319 1435 323 1439
rect 391 1435 395 1439
rect 471 1435 475 1439
rect 559 1435 563 1439
rect 647 1435 651 1439
rect 727 1435 731 1439
rect 807 1435 811 1439
rect 879 1435 883 1439
rect 943 1435 947 1439
rect 999 1435 1003 1439
rect 1047 1435 1051 1439
rect 1103 1435 1107 1439
rect 1151 1435 1155 1439
rect 1191 1435 1195 1439
rect 1279 1420 1283 1424
rect 1827 1423 1831 1427
rect 2267 1423 2271 1427
rect 2303 1423 2307 1427
rect 111 1412 115 1416
rect 1239 1412 1243 1416
rect 1351 1415 1355 1419
rect 1451 1415 1455 1419
rect 1579 1415 1580 1419
rect 1580 1415 1583 1419
rect 1667 1415 1668 1419
rect 1668 1415 1671 1419
rect 1719 1415 1723 1419
rect 1835 1415 1836 1419
rect 1836 1415 1839 1419
rect 1907 1415 1908 1419
rect 1908 1415 1911 1419
rect 167 1407 168 1411
rect 168 1407 171 1411
rect 207 1407 208 1411
rect 208 1407 211 1411
rect 251 1407 252 1411
rect 252 1407 255 1411
rect 347 1407 348 1411
rect 348 1407 351 1411
rect 419 1407 420 1411
rect 420 1407 423 1411
rect 499 1407 500 1411
rect 500 1407 503 1411
rect 587 1407 588 1411
rect 588 1407 591 1411
rect 111 1395 115 1399
rect 375 1399 379 1403
rect 755 1407 756 1411
rect 756 1407 759 1411
rect 835 1407 836 1411
rect 836 1407 839 1411
rect 907 1407 908 1411
rect 908 1407 911 1411
rect 971 1407 972 1411
rect 972 1407 975 1411
rect 1027 1407 1028 1411
rect 1028 1407 1031 1411
rect 1075 1407 1076 1411
rect 1076 1407 1079 1411
rect 1139 1407 1143 1411
rect 1175 1407 1176 1411
rect 1176 1407 1179 1411
rect 1087 1399 1091 1403
rect 2035 1415 2039 1419
rect 2083 1415 2087 1419
rect 2131 1415 2135 1419
rect 2179 1415 2183 1419
rect 2227 1415 2231 1419
rect 2407 1420 2411 1424
rect 2375 1415 2379 1419
rect 1279 1403 1283 1407
rect 2015 1407 2019 1411
rect 2407 1403 2411 1407
rect 1239 1395 1243 1399
rect 1375 1396 1379 1400
rect 1463 1396 1467 1400
rect 1551 1396 1555 1400
rect 1639 1396 1643 1400
rect 1727 1396 1731 1400
rect 1807 1396 1811 1400
rect 1879 1396 1883 1400
rect 1943 1396 1947 1400
rect 1999 1396 2003 1400
rect 2047 1396 2051 1400
rect 2095 1396 2099 1400
rect 2143 1396 2147 1400
rect 2191 1396 2195 1400
rect 2239 1396 2243 1400
rect 2279 1396 2283 1400
rect 2319 1396 2323 1400
rect 2359 1396 2363 1400
rect 143 1388 147 1392
rect 183 1388 187 1392
rect 223 1388 227 1392
rect 263 1388 267 1392
rect 319 1388 323 1392
rect 391 1388 395 1392
rect 471 1388 475 1392
rect 559 1388 563 1392
rect 647 1388 651 1392
rect 727 1388 731 1392
rect 807 1388 811 1392
rect 879 1388 883 1392
rect 943 1388 947 1392
rect 999 1388 1003 1392
rect 1047 1388 1051 1392
rect 1103 1388 1107 1392
rect 1151 1388 1155 1392
rect 1191 1388 1195 1392
rect 167 1376 171 1380
rect 207 1376 211 1380
rect 247 1376 251 1380
rect 303 1376 307 1380
rect 367 1376 371 1380
rect 439 1376 443 1380
rect 519 1376 523 1380
rect 599 1376 603 1380
rect 679 1376 683 1380
rect 751 1376 755 1380
rect 823 1376 827 1380
rect 887 1376 891 1380
rect 951 1376 955 1380
rect 1015 1376 1019 1380
rect 1079 1376 1083 1380
rect 1143 1376 1147 1380
rect 1191 1376 1195 1380
rect 1303 1376 1307 1380
rect 1343 1376 1347 1380
rect 1399 1376 1403 1380
rect 1463 1376 1467 1380
rect 1535 1376 1539 1380
rect 1607 1376 1611 1380
rect 1687 1376 1691 1380
rect 1767 1376 1771 1380
rect 1847 1376 1851 1380
rect 1935 1376 1939 1380
rect 2023 1376 2027 1380
rect 2111 1376 2115 1380
rect 2199 1376 2203 1380
rect 2287 1376 2291 1380
rect 2359 1376 2363 1380
rect 111 1369 115 1373
rect 1239 1369 1243 1373
rect 1279 1369 1283 1373
rect 2407 1369 2411 1373
rect 159 1363 163 1367
rect 111 1352 115 1356
rect 195 1355 196 1359
rect 196 1355 199 1359
rect 235 1355 236 1359
rect 236 1355 239 1359
rect 295 1355 299 1359
rect 743 1363 747 1367
rect 431 1355 435 1359
rect 511 1355 515 1359
rect 591 1355 595 1359
rect 607 1355 611 1359
rect 743 1355 747 1359
rect 815 1355 819 1359
rect 879 1355 883 1359
rect 943 1355 947 1359
rect 1007 1355 1011 1359
rect 1135 1355 1139 1359
rect 1183 1355 1187 1359
rect 1231 1355 1235 1359
rect 1239 1352 1243 1356
rect 1279 1352 1283 1356
rect 1311 1355 1315 1359
rect 1391 1355 1395 1359
rect 1455 1355 1459 1359
rect 1491 1355 1492 1359
rect 1492 1355 1495 1359
rect 1559 1355 1560 1359
rect 1560 1355 1563 1359
rect 1783 1355 1787 1359
rect 2103 1355 2107 1359
rect 1943 1347 1947 1351
rect 2271 1355 2275 1359
rect 2311 1355 2312 1359
rect 2312 1355 2315 1359
rect 2367 1355 2371 1359
rect 2407 1352 2411 1356
rect 167 1329 171 1333
rect 207 1329 211 1333
rect 247 1329 251 1333
rect 303 1329 307 1333
rect 367 1329 371 1333
rect 439 1329 443 1333
rect 519 1329 523 1333
rect 599 1329 603 1333
rect 679 1329 683 1333
rect 751 1329 755 1333
rect 823 1329 827 1333
rect 887 1329 891 1333
rect 951 1329 955 1333
rect 1015 1329 1019 1333
rect 1079 1329 1083 1333
rect 1143 1329 1147 1333
rect 1191 1329 1195 1333
rect 1303 1329 1307 1333
rect 1343 1329 1347 1333
rect 1399 1329 1403 1333
rect 1463 1329 1467 1333
rect 1535 1329 1539 1333
rect 1607 1329 1611 1333
rect 1687 1329 1691 1333
rect 1767 1329 1771 1333
rect 1847 1329 1851 1333
rect 1935 1329 1939 1333
rect 2023 1329 2027 1333
rect 2111 1329 2115 1333
rect 2199 1329 2203 1333
rect 2287 1329 2291 1333
rect 2359 1329 2363 1333
rect 175 1319 179 1323
rect 195 1319 199 1323
rect 235 1319 239 1323
rect 295 1319 299 1323
rect 375 1319 379 1323
rect 431 1319 435 1323
rect 511 1319 515 1323
rect 591 1319 595 1323
rect 743 1319 747 1323
rect 815 1319 819 1323
rect 879 1319 883 1323
rect 943 1319 947 1323
rect 1007 1319 1011 1323
rect 1087 1319 1091 1323
rect 1135 1319 1139 1323
rect 1183 1319 1187 1323
rect 1231 1319 1235 1323
rect 1351 1319 1355 1323
rect 1391 1319 1395 1323
rect 1455 1319 1459 1323
rect 1755 1319 1759 1323
rect 1943 1319 1947 1323
rect 2015 1319 2019 1323
rect 2103 1319 2107 1323
rect 2263 1319 2267 1323
rect 2271 1319 2275 1323
rect 2375 1319 2379 1323
rect 1023 1311 1027 1315
rect 219 1303 223 1307
rect 255 1303 259 1307
rect 279 1303 283 1307
rect 315 1303 319 1307
rect 379 1303 383 1307
rect 451 1303 455 1307
rect 655 1303 659 1307
rect 667 1303 671 1307
rect 731 1303 735 1307
rect 795 1303 799 1307
rect 851 1303 855 1307
rect 907 1303 911 1307
rect 963 1303 967 1307
rect 1311 1307 1315 1311
rect 1331 1307 1335 1311
rect 1371 1307 1375 1311
rect 1411 1307 1415 1311
rect 1447 1307 1451 1311
rect 1491 1307 1495 1311
rect 1527 1307 1531 1311
rect 1551 1307 1555 1311
rect 1615 1307 1619 1311
rect 1651 1307 1655 1311
rect 1783 1307 1787 1311
rect 1819 1307 1823 1311
rect 1875 1307 1879 1311
rect 1995 1307 1999 1311
rect 2067 1307 2071 1311
rect 2147 1307 2151 1311
rect 2251 1307 2255 1311
rect 2367 1307 2371 1311
rect 183 1295 187 1299
rect 231 1295 235 1299
rect 287 1295 291 1299
rect 351 1295 355 1299
rect 423 1295 427 1299
rect 495 1295 499 1299
rect 567 1295 571 1299
rect 639 1295 643 1299
rect 703 1295 707 1299
rect 767 1295 771 1299
rect 823 1295 827 1299
rect 879 1295 883 1299
rect 935 1295 939 1299
rect 999 1295 1003 1299
rect 1303 1299 1307 1303
rect 1343 1299 1347 1303
rect 1383 1299 1387 1303
rect 1423 1299 1427 1303
rect 1463 1299 1467 1303
rect 1503 1299 1507 1303
rect 1543 1299 1547 1303
rect 1583 1299 1587 1303
rect 1623 1299 1627 1303
rect 1679 1299 1683 1303
rect 1735 1299 1739 1303
rect 1791 1299 1795 1303
rect 1847 1299 1851 1303
rect 1903 1299 1907 1303
rect 1967 1299 1971 1303
rect 2039 1299 2043 1303
rect 2119 1299 2123 1303
rect 2199 1299 2203 1303
rect 2287 1299 2291 1303
rect 2359 1299 2363 1303
rect 111 1272 115 1276
rect 175 1267 179 1271
rect 219 1267 223 1271
rect 315 1267 316 1271
rect 316 1267 319 1271
rect 379 1267 380 1271
rect 380 1267 383 1271
rect 451 1267 452 1271
rect 452 1267 455 1271
rect 1239 1272 1243 1276
rect 1279 1276 1283 1280
rect 583 1267 587 1271
rect 667 1267 668 1271
rect 668 1267 671 1271
rect 731 1267 732 1271
rect 732 1267 735 1271
rect 795 1267 796 1271
rect 796 1267 799 1271
rect 851 1267 852 1271
rect 852 1267 855 1271
rect 907 1267 908 1271
rect 908 1267 911 1271
rect 963 1267 964 1271
rect 964 1267 967 1271
rect 1331 1271 1332 1275
rect 1332 1271 1335 1275
rect 1023 1267 1024 1271
rect 1024 1267 1027 1271
rect 1371 1271 1372 1275
rect 1372 1271 1375 1275
rect 1411 1271 1412 1275
rect 1412 1271 1415 1275
rect 1447 1271 1448 1275
rect 1448 1271 1451 1275
rect 1551 1279 1555 1283
rect 2407 1276 2411 1280
rect 1527 1271 1528 1275
rect 1528 1271 1531 1275
rect 1571 1271 1572 1275
rect 1572 1271 1575 1275
rect 1611 1271 1612 1275
rect 1612 1271 1615 1275
rect 1651 1271 1652 1275
rect 1652 1271 1655 1275
rect 1755 1271 1759 1275
rect 1819 1271 1820 1275
rect 1820 1271 1823 1275
rect 1875 1271 1876 1275
rect 1876 1271 1879 1275
rect 1995 1271 1996 1275
rect 1996 1271 1999 1275
rect 2067 1271 2068 1275
rect 2068 1271 2071 1275
rect 2147 1271 2148 1275
rect 2148 1271 2151 1275
rect 111 1255 115 1259
rect 1239 1255 1243 1259
rect 1279 1259 1283 1263
rect 1807 1263 1811 1267
rect 2263 1271 2267 1275
rect 2367 1271 2371 1275
rect 2407 1259 2411 1263
rect 183 1248 187 1252
rect 231 1248 235 1252
rect 287 1248 291 1252
rect 351 1248 355 1252
rect 423 1248 427 1252
rect 495 1248 499 1252
rect 567 1248 571 1252
rect 639 1248 643 1252
rect 703 1248 707 1252
rect 767 1248 771 1252
rect 823 1248 827 1252
rect 879 1248 883 1252
rect 935 1248 939 1252
rect 999 1248 1003 1252
rect 1303 1252 1307 1256
rect 1343 1252 1347 1256
rect 1383 1252 1387 1256
rect 1423 1252 1427 1256
rect 1463 1252 1467 1256
rect 1503 1252 1507 1256
rect 1543 1252 1547 1256
rect 1583 1252 1587 1256
rect 1623 1252 1627 1256
rect 1679 1252 1683 1256
rect 1735 1252 1739 1256
rect 1791 1252 1795 1256
rect 1847 1252 1851 1256
rect 1903 1252 1907 1256
rect 1967 1252 1971 1256
rect 2039 1252 2043 1256
rect 2119 1252 2123 1256
rect 2199 1252 2203 1256
rect 2287 1252 2291 1256
rect 2359 1252 2363 1256
rect 135 1232 139 1236
rect 175 1232 179 1236
rect 231 1232 235 1236
rect 311 1232 315 1236
rect 399 1232 403 1236
rect 487 1232 491 1236
rect 575 1232 579 1236
rect 663 1232 667 1236
rect 743 1232 747 1236
rect 815 1232 819 1236
rect 879 1232 883 1236
rect 943 1232 947 1236
rect 1007 1232 1011 1236
rect 1071 1232 1075 1236
rect 1303 1232 1307 1236
rect 1375 1232 1379 1236
rect 1479 1232 1483 1236
rect 1583 1232 1587 1236
rect 1687 1232 1691 1236
rect 1791 1232 1795 1236
rect 1887 1232 1891 1236
rect 1983 1232 1987 1236
rect 2071 1232 2075 1236
rect 2151 1232 2155 1236
rect 2223 1232 2227 1236
rect 2303 1232 2307 1236
rect 2359 1232 2363 1236
rect 111 1225 115 1229
rect 1239 1225 1243 1229
rect 1279 1225 1283 1229
rect 2407 1225 2411 1229
rect 111 1208 115 1212
rect 163 1211 164 1215
rect 164 1211 167 1215
rect 223 1211 227 1215
rect 255 1211 256 1215
rect 256 1211 259 1215
rect 655 1211 659 1215
rect 711 1211 715 1215
rect 1239 1208 1243 1212
rect 1279 1208 1283 1212
rect 1311 1211 1315 1215
rect 1679 1211 1683 1215
rect 1495 1203 1499 1207
rect 1879 1211 1883 1215
rect 1975 1211 1979 1215
rect 2063 1211 2067 1215
rect 2143 1211 2147 1215
rect 1911 1203 1915 1207
rect 2251 1211 2252 1215
rect 2252 1211 2255 1215
rect 2351 1211 2355 1215
rect 2311 1203 2315 1207
rect 2407 1208 2411 1212
rect 135 1185 139 1189
rect 175 1185 179 1189
rect 231 1185 235 1189
rect 311 1185 315 1189
rect 399 1185 403 1189
rect 487 1185 491 1189
rect 575 1185 579 1189
rect 663 1185 667 1189
rect 743 1185 747 1189
rect 815 1185 819 1189
rect 879 1185 883 1189
rect 943 1185 947 1189
rect 1007 1185 1011 1189
rect 1071 1185 1075 1189
rect 1303 1185 1307 1189
rect 1375 1185 1379 1189
rect 1479 1185 1483 1189
rect 1583 1185 1587 1189
rect 1687 1185 1691 1189
rect 1791 1185 1795 1189
rect 1887 1185 1891 1189
rect 1983 1185 1987 1189
rect 2071 1185 2075 1189
rect 2151 1185 2155 1189
rect 2223 1185 2227 1189
rect 2303 1185 2307 1189
rect 2359 1185 2363 1189
rect 155 1175 159 1179
rect 163 1175 167 1179
rect 223 1175 227 1179
rect 583 1175 587 1179
rect 711 1175 715 1179
rect 1215 1175 1219 1179
rect 1495 1175 1499 1179
rect 1571 1175 1575 1179
rect 1679 1175 1683 1179
rect 1807 1175 1811 1179
rect 1879 1175 1883 1179
rect 1975 1175 1979 1179
rect 2063 1175 2067 1179
rect 2143 1175 2147 1179
rect 2187 1175 2191 1179
rect 2311 1175 2315 1179
rect 2367 1175 2371 1179
rect 147 1163 151 1167
rect 163 1163 167 1167
rect 355 1163 359 1167
rect 459 1163 463 1167
rect 563 1163 567 1167
rect 763 1163 767 1167
rect 771 1163 775 1167
rect 867 1163 871 1167
rect 971 1163 975 1167
rect 1027 1163 1031 1167
rect 1099 1163 1103 1167
rect 1171 1163 1175 1167
rect 1311 1163 1315 1167
rect 1331 1163 1335 1167
rect 1435 1163 1439 1167
rect 1515 1163 1519 1167
rect 1611 1163 1615 1167
rect 1715 1163 1719 1167
rect 1911 1163 1915 1167
rect 1931 1163 1935 1167
rect 2027 1163 2031 1167
rect 2291 1163 2295 1167
rect 2343 1163 2347 1167
rect 2351 1163 2355 1167
rect 135 1155 139 1159
rect 175 1155 179 1159
rect 239 1155 243 1159
rect 327 1155 331 1159
rect 431 1155 435 1159
rect 535 1155 539 1159
rect 639 1155 643 1159
rect 743 1155 747 1159
rect 839 1155 843 1159
rect 919 1155 923 1159
rect 999 1155 1003 1159
rect 1071 1155 1075 1159
rect 1143 1155 1147 1159
rect 1191 1155 1195 1159
rect 1303 1155 1307 1159
rect 1343 1155 1347 1159
rect 1407 1155 1411 1159
rect 1487 1155 1491 1159
rect 1583 1155 1587 1159
rect 1687 1155 1691 1159
rect 1799 1155 1803 1159
rect 1903 1155 1907 1159
rect 1999 1155 2003 1159
rect 2079 1155 2083 1159
rect 2159 1155 2163 1159
rect 2231 1155 2235 1159
rect 2303 1155 2307 1159
rect 2359 1155 2363 1159
rect 111 1132 115 1136
rect 147 1135 151 1139
rect 1239 1132 1243 1136
rect 155 1127 159 1131
rect 355 1127 356 1131
rect 356 1127 359 1131
rect 459 1127 460 1131
rect 460 1127 463 1131
rect 563 1127 564 1131
rect 564 1127 567 1131
rect 771 1127 772 1131
rect 772 1127 775 1131
rect 867 1127 868 1131
rect 868 1127 871 1131
rect 971 1127 975 1131
rect 1027 1127 1028 1131
rect 1028 1127 1031 1131
rect 1099 1127 1100 1131
rect 1100 1127 1103 1131
rect 1171 1127 1172 1131
rect 1172 1127 1175 1131
rect 1279 1132 1283 1136
rect 2407 1132 2411 1136
rect 1215 1127 1216 1131
rect 1216 1127 1219 1131
rect 1331 1127 1332 1131
rect 1332 1127 1335 1131
rect 1435 1127 1436 1131
rect 1436 1127 1439 1131
rect 1515 1127 1516 1131
rect 1516 1127 1519 1131
rect 1611 1127 1612 1131
rect 1612 1127 1615 1131
rect 1715 1127 1716 1131
rect 1716 1127 1719 1131
rect 1735 1127 1739 1131
rect 1931 1127 1932 1131
rect 1932 1127 1935 1131
rect 2027 1127 2028 1131
rect 2028 1127 2031 1131
rect 2167 1127 2171 1131
rect 2187 1127 2188 1131
rect 2188 1127 2191 1131
rect 2291 1127 2295 1131
rect 2343 1127 2347 1131
rect 111 1115 115 1119
rect 347 1119 351 1123
rect 1239 1115 1243 1119
rect 1279 1115 1283 1119
rect 2407 1115 2411 1119
rect 135 1108 139 1112
rect 175 1108 179 1112
rect 239 1108 243 1112
rect 327 1108 331 1112
rect 431 1108 435 1112
rect 535 1108 539 1112
rect 639 1108 643 1112
rect 743 1108 747 1112
rect 839 1108 843 1112
rect 919 1108 923 1112
rect 999 1108 1003 1112
rect 1071 1108 1075 1112
rect 1143 1108 1147 1112
rect 1191 1108 1195 1112
rect 1303 1108 1307 1112
rect 1343 1108 1347 1112
rect 1407 1108 1411 1112
rect 1487 1108 1491 1112
rect 1583 1108 1587 1112
rect 1687 1108 1691 1112
rect 1799 1108 1803 1112
rect 1903 1108 1907 1112
rect 1999 1108 2003 1112
rect 2079 1108 2083 1112
rect 2159 1108 2163 1112
rect 2231 1108 2235 1112
rect 2303 1108 2307 1112
rect 2359 1108 2363 1112
rect 135 1092 139 1096
rect 175 1092 179 1096
rect 247 1092 251 1096
rect 327 1092 331 1096
rect 415 1092 419 1096
rect 503 1092 507 1096
rect 583 1092 587 1096
rect 663 1092 667 1096
rect 735 1092 739 1096
rect 799 1092 803 1096
rect 863 1092 867 1096
rect 919 1092 923 1096
rect 983 1092 987 1096
rect 1047 1092 1051 1096
rect 1431 1096 1435 1100
rect 1471 1096 1475 1100
rect 1511 1096 1515 1100
rect 1559 1096 1563 1100
rect 1615 1096 1619 1100
rect 1671 1096 1675 1100
rect 1727 1096 1731 1100
rect 1775 1096 1779 1100
rect 1823 1096 1827 1100
rect 1871 1096 1875 1100
rect 1919 1096 1923 1100
rect 1967 1096 1971 1100
rect 2015 1096 2019 1100
rect 2063 1096 2067 1100
rect 2119 1096 2123 1100
rect 2175 1096 2179 1100
rect 2231 1096 2235 1100
rect 111 1085 115 1089
rect 1239 1085 1243 1089
rect 1279 1089 1283 1093
rect 2407 1089 2411 1093
rect 111 1068 115 1072
rect 163 1071 164 1075
rect 164 1071 167 1075
rect 239 1071 243 1075
rect 143 1063 147 1067
rect 407 1071 411 1075
rect 495 1071 499 1075
rect 335 1063 339 1067
rect 727 1071 731 1075
rect 791 1071 795 1075
rect 855 1071 859 1075
rect 911 1071 915 1075
rect 975 1071 979 1075
rect 1039 1071 1043 1075
rect 1071 1071 1072 1075
rect 1072 1071 1075 1075
rect 1239 1068 1243 1072
rect 1279 1072 1283 1076
rect 1459 1075 1460 1079
rect 1460 1075 1463 1079
rect 1499 1075 1500 1079
rect 1500 1075 1503 1079
rect 1551 1075 1555 1079
rect 1607 1075 1611 1079
rect 1663 1075 1667 1079
rect 1715 1075 1719 1079
rect 1583 1067 1587 1071
rect 1815 1075 1819 1079
rect 1783 1067 1787 1071
rect 2003 1075 2007 1079
rect 2223 1075 2227 1079
rect 2247 1075 2251 1079
rect 2407 1072 2411 1076
rect 135 1045 139 1049
rect 175 1045 179 1049
rect 247 1045 251 1049
rect 327 1045 331 1049
rect 415 1045 419 1049
rect 503 1045 507 1049
rect 583 1045 587 1049
rect 663 1045 667 1049
rect 735 1045 739 1049
rect 799 1045 803 1049
rect 863 1045 867 1049
rect 919 1045 923 1049
rect 983 1045 987 1049
rect 1047 1045 1051 1049
rect 1431 1049 1435 1053
rect 1471 1049 1475 1053
rect 1511 1049 1515 1053
rect 1559 1049 1563 1053
rect 1615 1049 1619 1053
rect 1671 1049 1675 1053
rect 1727 1049 1731 1053
rect 1775 1049 1779 1053
rect 1823 1049 1827 1053
rect 1871 1049 1875 1053
rect 1919 1049 1923 1053
rect 1967 1049 1971 1053
rect 2015 1049 2019 1053
rect 2063 1049 2067 1053
rect 2119 1049 2123 1053
rect 2175 1049 2179 1053
rect 2231 1049 2235 1053
rect 143 1035 147 1039
rect 199 1035 203 1039
rect 239 1035 243 1039
rect 347 1035 351 1039
rect 407 1035 411 1039
rect 495 1035 499 1039
rect 719 1035 723 1039
rect 727 1035 731 1039
rect 791 1035 795 1039
rect 855 1035 859 1039
rect 911 1035 915 1039
rect 975 1035 979 1039
rect 1039 1035 1043 1039
rect 1439 1039 1443 1043
rect 1459 1039 1463 1043
rect 1499 1039 1503 1043
rect 1551 1039 1555 1043
rect 1607 1039 1611 1043
rect 1663 1039 1667 1043
rect 1715 1039 1719 1043
rect 1783 1039 1787 1043
rect 2003 1039 2007 1043
rect 2111 1039 2115 1043
rect 2167 1039 2171 1043
rect 2223 1039 2227 1043
rect 239 1023 243 1027
rect 279 1023 283 1027
rect 335 1023 339 1027
rect 355 1023 359 1027
rect 427 1023 431 1027
rect 491 1023 495 1027
rect 547 1023 551 1027
rect 631 1023 635 1027
rect 651 1023 655 1027
rect 699 1023 703 1027
rect 763 1023 767 1027
rect 835 1023 839 1027
rect 927 1023 931 1027
rect 1027 1023 1031 1027
rect 1215 1023 1219 1027
rect 1583 1027 1587 1031
rect 1603 1027 1607 1031
rect 1643 1027 1647 1031
rect 1683 1027 1687 1031
rect 1719 1027 1723 1031
rect 1763 1027 1767 1031
rect 1815 1027 1819 1031
rect 1851 1027 1855 1031
rect 1907 1027 1911 1031
rect 2127 1027 2131 1031
rect 2239 1027 2243 1031
rect 2247 1027 2251 1031
rect 175 1015 179 1019
rect 255 1015 259 1019
rect 327 1015 331 1019
rect 399 1015 403 1019
rect 463 1015 467 1019
rect 519 1015 523 1019
rect 575 1015 579 1019
rect 623 1015 627 1019
rect 671 1015 675 1019
rect 735 1015 739 1019
rect 807 1015 811 1019
rect 895 1015 899 1019
rect 999 1015 1003 1019
rect 1103 1015 1107 1019
rect 1191 1015 1195 1019
rect 1575 1019 1579 1023
rect 1615 1019 1619 1023
rect 1655 1019 1659 1023
rect 1695 1019 1699 1023
rect 1735 1019 1739 1023
rect 1775 1019 1779 1023
rect 1823 1019 1827 1023
rect 1879 1019 1883 1023
rect 1943 1019 1947 1023
rect 2015 1019 2019 1023
rect 2095 1019 2099 1023
rect 2175 1019 2179 1023
rect 2255 1019 2259 1023
rect 111 992 115 996
rect 1239 992 1243 996
rect 1279 996 1283 1000
rect 199 987 200 991
rect 200 987 203 991
rect 239 987 243 991
rect 355 987 356 991
rect 356 987 359 991
rect 427 987 428 991
rect 428 987 431 991
rect 491 987 492 991
rect 492 987 495 991
rect 547 987 548 991
rect 548 987 551 991
rect 111 975 115 979
rect 471 979 475 983
rect 651 987 652 991
rect 652 987 655 991
rect 699 987 700 991
rect 700 987 703 991
rect 763 987 764 991
rect 764 987 767 991
rect 835 987 836 991
rect 836 987 839 991
rect 923 987 924 991
rect 924 987 927 991
rect 1027 987 1028 991
rect 1028 987 1031 991
rect 1127 987 1128 991
rect 1128 987 1131 991
rect 1151 987 1155 991
rect 1603 991 1604 995
rect 1604 991 1607 995
rect 1643 991 1644 995
rect 1644 991 1647 995
rect 1683 991 1684 995
rect 1684 991 1687 995
rect 1719 991 1720 995
rect 1720 991 1723 995
rect 1763 991 1764 995
rect 1764 991 1767 995
rect 1239 975 1243 979
rect 1279 979 1283 983
rect 1687 983 1691 987
rect 1851 991 1852 995
rect 1852 991 1855 995
rect 1907 991 1908 995
rect 1908 991 1911 995
rect 2407 996 2411 1000
rect 2111 991 2115 995
rect 2191 991 2195 995
rect 2239 991 2243 995
rect 2407 979 2411 983
rect 175 968 179 972
rect 255 968 259 972
rect 327 968 331 972
rect 399 968 403 972
rect 463 968 467 972
rect 519 968 523 972
rect 575 968 579 972
rect 623 968 627 972
rect 671 968 675 972
rect 735 968 739 972
rect 807 968 811 972
rect 895 968 899 972
rect 999 968 1003 972
rect 1103 968 1107 972
rect 1191 968 1195 972
rect 1575 972 1579 976
rect 1615 972 1619 976
rect 1655 972 1659 976
rect 1695 972 1699 976
rect 1735 972 1739 976
rect 1775 972 1779 976
rect 1823 972 1827 976
rect 1879 972 1883 976
rect 1943 972 1947 976
rect 2015 972 2019 976
rect 2095 972 2099 976
rect 2175 972 2179 976
rect 2255 972 2259 976
rect 215 956 219 960
rect 255 956 259 960
rect 303 956 307 960
rect 359 956 363 960
rect 415 956 419 960
rect 463 956 467 960
rect 519 956 523 960
rect 575 956 579 960
rect 639 956 643 960
rect 711 956 715 960
rect 783 956 787 960
rect 855 956 859 960
rect 927 956 931 960
rect 999 956 1003 960
rect 1071 956 1075 960
rect 1143 956 1147 960
rect 1191 956 1195 960
rect 111 949 115 953
rect 1239 949 1243 953
rect 1303 952 1307 956
rect 1351 952 1355 956
rect 1431 952 1435 956
rect 1511 952 1515 956
rect 1591 952 1595 956
rect 1679 952 1683 956
rect 1767 952 1771 956
rect 1855 952 1859 956
rect 1943 952 1947 956
rect 2023 952 2027 956
rect 2103 952 2107 956
rect 2183 952 2187 956
rect 2271 952 2275 956
rect 631 943 635 947
rect 1279 945 1283 949
rect 2407 945 2411 949
rect 111 932 115 936
rect 243 935 244 939
rect 244 935 247 939
rect 279 935 280 939
rect 280 935 283 939
rect 223 927 227 931
rect 347 935 351 939
rect 503 935 507 939
rect 559 935 563 939
rect 631 935 635 939
rect 703 935 707 939
rect 775 935 779 939
rect 847 935 851 939
rect 991 935 995 939
rect 1015 935 1019 939
rect 939 927 943 931
rect 1215 935 1216 939
rect 1216 935 1219 939
rect 1239 932 1243 936
rect 1279 928 1283 932
rect 1287 931 1291 935
rect 1647 931 1651 935
rect 1783 931 1787 935
rect 2095 931 2099 935
rect 2127 931 2128 935
rect 2128 931 2131 935
rect 2263 931 2267 935
rect 2287 931 2291 935
rect 2407 928 2411 932
rect 215 909 219 913
rect 255 909 259 913
rect 303 909 307 913
rect 359 909 363 913
rect 415 909 419 913
rect 463 909 467 913
rect 519 909 523 913
rect 575 909 579 913
rect 639 909 643 913
rect 711 909 715 913
rect 783 909 787 913
rect 855 909 859 913
rect 927 909 931 913
rect 999 909 1003 913
rect 1071 909 1075 913
rect 1143 909 1147 913
rect 1191 909 1195 913
rect 1303 905 1307 909
rect 1351 905 1355 909
rect 1431 905 1435 909
rect 1511 905 1515 909
rect 1591 905 1595 909
rect 1679 905 1683 909
rect 1767 905 1771 909
rect 1855 905 1859 909
rect 1943 905 1947 909
rect 2023 905 2027 909
rect 2103 905 2107 909
rect 2183 905 2187 909
rect 2271 905 2275 909
rect 223 899 227 903
rect 243 899 247 903
rect 347 899 351 903
rect 471 899 475 903
rect 503 899 507 903
rect 559 899 563 903
rect 631 899 635 903
rect 703 899 707 903
rect 775 899 779 903
rect 847 899 851 903
rect 939 899 943 903
rect 991 899 995 903
rect 1151 899 1155 903
rect 1287 899 1291 903
rect 275 887 279 891
rect 663 891 667 895
rect 1571 895 1575 899
rect 1687 895 1691 899
rect 2087 895 2091 899
rect 2095 895 2099 899
rect 2191 895 2195 899
rect 2263 895 2267 899
rect 191 871 195 875
rect 215 875 219 879
rect 231 871 235 875
rect 255 875 259 879
rect 387 879 391 883
rect 499 879 503 883
rect 603 879 607 883
rect 747 879 751 883
rect 755 879 759 883
rect 947 879 951 883
rect 1007 879 1011 883
rect 1015 879 1019 883
rect 1051 879 1055 883
rect 1115 879 1119 883
rect 1455 883 1459 887
rect 1463 883 1467 887
rect 1503 883 1507 887
rect 1547 883 1551 887
rect 1647 883 1651 887
rect 1783 883 1787 887
rect 1803 883 1807 887
rect 1875 883 1879 887
rect 2111 883 2115 887
rect 2203 883 2207 887
rect 2279 883 2283 887
rect 2287 883 2291 887
rect 287 871 291 875
rect 359 871 363 875
rect 447 871 451 875
rect 543 871 547 875
rect 639 871 643 875
rect 727 871 731 875
rect 807 871 811 875
rect 887 871 891 875
rect 959 871 963 875
rect 1023 871 1027 875
rect 1087 871 1091 875
rect 1159 871 1163 875
rect 1439 875 1443 879
rect 1479 875 1483 879
rect 1519 875 1523 879
rect 1559 875 1563 879
rect 1607 875 1611 879
rect 1655 875 1659 879
rect 1711 875 1715 879
rect 1775 875 1779 879
rect 1847 875 1851 879
rect 1919 875 1923 879
rect 1991 875 1995 879
rect 2063 875 2067 879
rect 2135 875 2139 879
rect 2215 875 2219 879
rect 2295 875 2299 879
rect 111 848 115 852
rect 747 851 751 855
rect 215 843 216 847
rect 216 843 219 847
rect 255 843 256 847
rect 256 843 259 847
rect 387 843 388 847
rect 388 843 391 847
rect 499 843 503 847
rect 603 843 607 847
rect 663 843 664 847
rect 664 843 667 847
rect 755 843 756 847
rect 756 843 759 847
rect 871 843 875 847
rect 1007 851 1011 855
rect 947 843 951 847
rect 1051 843 1052 847
rect 1052 843 1055 847
rect 1115 843 1116 847
rect 1116 843 1119 847
rect 1239 848 1243 852
rect 1279 852 1283 856
rect 1571 855 1575 859
rect 1463 847 1464 851
rect 1464 847 1467 851
rect 1503 847 1504 851
rect 1504 847 1507 851
rect 1547 847 1548 851
rect 1548 847 1551 851
rect 1719 847 1723 851
rect 1803 847 1804 851
rect 1804 847 1807 851
rect 1875 847 1876 851
rect 1876 847 1879 851
rect 2407 852 2411 856
rect 111 831 115 835
rect 1239 831 1243 835
rect 1279 835 1283 839
rect 1767 839 1771 843
rect 2087 847 2088 851
rect 2088 847 2091 851
rect 2111 847 2115 851
rect 2203 847 2207 851
rect 2279 847 2283 851
rect 2407 835 2411 839
rect 191 824 195 828
rect 231 824 235 828
rect 287 824 291 828
rect 359 824 363 828
rect 447 824 451 828
rect 543 824 547 828
rect 639 824 643 828
rect 727 824 731 828
rect 807 824 811 828
rect 887 824 891 828
rect 959 824 963 828
rect 1023 824 1027 828
rect 1087 824 1091 828
rect 1159 824 1163 828
rect 1439 828 1443 832
rect 1479 828 1483 832
rect 1519 828 1523 832
rect 1559 828 1563 832
rect 1607 828 1611 832
rect 1655 828 1659 832
rect 1711 828 1715 832
rect 1775 828 1779 832
rect 1847 828 1851 832
rect 1919 828 1923 832
rect 1991 828 1995 832
rect 2063 828 2067 832
rect 2135 828 2139 832
rect 2215 828 2219 832
rect 2295 828 2299 832
rect 135 812 139 816
rect 175 812 179 816
rect 239 812 243 816
rect 327 812 331 816
rect 415 812 419 816
rect 503 812 507 816
rect 591 812 595 816
rect 671 812 675 816
rect 743 812 747 816
rect 815 812 819 816
rect 879 812 883 816
rect 943 812 947 816
rect 1015 812 1019 816
rect 111 805 115 809
rect 1239 805 1243 809
rect 1359 804 1363 808
rect 1415 804 1419 808
rect 1471 804 1475 808
rect 1535 804 1539 808
rect 1591 804 1595 808
rect 1647 804 1651 808
rect 1703 804 1707 808
rect 1759 804 1763 808
rect 1815 804 1819 808
rect 1871 804 1875 808
rect 1935 804 1939 808
rect 1999 804 2003 808
rect 2071 804 2075 808
rect 2143 804 2147 808
rect 2223 804 2227 808
rect 2303 804 2307 808
rect 2359 804 2363 808
rect 275 799 279 803
rect 111 788 115 792
rect 163 791 164 795
rect 164 791 167 795
rect 231 791 235 795
rect 319 791 323 795
rect 407 791 411 795
rect 495 791 499 795
rect 1279 797 1283 801
rect 2407 797 2411 801
rect 663 791 667 795
rect 735 791 739 795
rect 807 791 811 795
rect 607 783 611 787
rect 935 791 939 795
rect 1007 791 1011 795
rect 823 783 827 787
rect 1239 788 1243 792
rect 1455 791 1459 795
rect 1279 780 1283 784
rect 1399 783 1403 787
rect 1463 783 1467 787
rect 1527 783 1531 787
rect 1639 783 1643 787
rect 1671 783 1672 787
rect 1672 783 1675 787
rect 1599 775 1603 779
rect 1799 783 1803 787
rect 1863 783 1867 787
rect 1927 783 1931 787
rect 1983 783 1987 787
rect 2063 783 2067 787
rect 2135 783 2139 787
rect 2151 783 2155 787
rect 2295 783 2299 787
rect 2351 783 2355 787
rect 2371 783 2375 787
rect 2407 780 2411 784
rect 135 765 139 769
rect 175 765 179 769
rect 239 765 243 769
rect 327 765 331 769
rect 415 765 419 769
rect 503 765 507 769
rect 591 765 595 769
rect 671 765 675 769
rect 743 765 747 769
rect 815 765 819 769
rect 879 765 883 769
rect 943 765 947 769
rect 1015 765 1019 769
rect 155 755 159 759
rect 163 755 167 759
rect 231 755 235 759
rect 319 755 323 759
rect 407 755 411 759
rect 495 755 499 759
rect 607 755 611 759
rect 663 755 667 759
rect 735 755 739 759
rect 823 755 827 759
rect 871 755 875 759
rect 935 755 939 759
rect 1007 755 1011 759
rect 1359 757 1363 761
rect 1415 757 1419 761
rect 1471 757 1475 761
rect 1535 757 1539 761
rect 1591 757 1595 761
rect 1647 757 1651 761
rect 1703 757 1707 761
rect 1759 757 1763 761
rect 1815 757 1819 761
rect 1871 757 1875 761
rect 1935 757 1939 761
rect 1999 757 2003 761
rect 2071 757 2075 761
rect 2143 757 2147 761
rect 2223 757 2227 761
rect 2303 757 2307 761
rect 2359 757 2363 761
rect 1391 747 1395 751
rect 1399 747 1403 751
rect 1463 747 1467 751
rect 1527 747 1531 751
rect 1599 747 1603 751
rect 1639 747 1643 751
rect 1719 747 1723 751
rect 1767 747 1771 751
rect 1799 747 1803 751
rect 1863 747 1867 751
rect 1927 747 1931 751
rect 1983 747 1987 751
rect 2063 747 2067 751
rect 2135 747 2139 751
rect 2287 747 2291 751
rect 2295 747 2299 751
rect 2351 747 2355 751
rect 223 739 227 743
rect 387 739 391 743
rect 443 739 447 743
rect 491 739 495 743
rect 531 739 535 743
rect 571 739 575 743
rect 611 739 615 743
rect 659 739 663 743
rect 699 739 703 743
rect 707 739 711 743
rect 755 739 759 743
rect 807 739 811 743
rect 851 739 855 743
rect 899 739 903 743
rect 135 731 139 735
rect 191 731 195 735
rect 263 731 267 735
rect 335 731 339 735
rect 399 731 403 735
rect 455 731 459 735
rect 503 731 507 735
rect 543 731 547 735
rect 583 731 587 735
rect 623 731 627 735
rect 671 731 675 735
rect 719 731 723 735
rect 767 731 771 735
rect 815 731 819 735
rect 863 731 867 735
rect 911 731 915 735
rect 1323 735 1327 739
rect 1331 735 1335 739
rect 1371 735 1375 739
rect 1435 735 1439 739
rect 1515 735 1519 739
rect 1671 735 1675 739
rect 1691 735 1695 739
rect 1839 735 1843 739
rect 1859 735 1863 739
rect 1303 727 1307 731
rect 1343 727 1347 731
rect 1407 727 1411 731
rect 1487 727 1491 731
rect 1575 727 1579 731
rect 1663 727 1667 731
rect 1751 727 1755 731
rect 1831 727 1835 731
rect 1911 727 1915 731
rect 1935 731 1939 735
rect 2019 735 2023 739
rect 2107 735 2111 739
rect 2203 735 2207 739
rect 2371 735 2375 739
rect 1991 727 1995 731
rect 2079 727 2083 731
rect 2175 727 2179 731
rect 2279 727 2283 731
rect 2359 727 2363 731
rect 699 715 703 719
rect 111 708 115 712
rect 155 703 159 707
rect 287 703 288 707
rect 288 703 291 707
rect 387 703 391 707
rect 443 703 447 707
rect 491 703 495 707
rect 539 703 543 707
rect 579 703 583 707
rect 619 703 623 707
rect 707 703 711 707
rect 755 707 759 711
rect 791 703 792 707
rect 792 703 795 707
rect 851 703 855 707
rect 899 703 903 707
rect 1239 708 1243 712
rect 1279 704 1283 708
rect 1391 707 1395 711
rect 1331 699 1332 703
rect 1332 699 1335 703
rect 1371 699 1372 703
rect 1372 699 1375 703
rect 1435 699 1436 703
rect 1436 699 1439 703
rect 1515 699 1516 703
rect 1516 699 1519 703
rect 2407 704 2411 708
rect 1691 699 1692 703
rect 1692 699 1695 703
rect 1735 699 1739 703
rect 1859 699 1860 703
rect 1860 699 1863 703
rect 1935 699 1936 703
rect 1936 699 1939 703
rect 2019 699 2020 703
rect 2020 699 2023 703
rect 2107 699 2108 703
rect 2108 699 2111 703
rect 2203 699 2204 703
rect 2204 699 2207 703
rect 2247 699 2251 703
rect 2379 699 2383 703
rect 111 691 115 695
rect 1239 691 1243 695
rect 135 684 139 688
rect 191 684 195 688
rect 263 684 267 688
rect 335 684 339 688
rect 399 684 403 688
rect 455 684 459 688
rect 503 684 507 688
rect 543 684 547 688
rect 583 684 587 688
rect 623 684 627 688
rect 671 684 675 688
rect 719 684 723 688
rect 767 684 771 688
rect 815 684 819 688
rect 863 684 867 688
rect 911 684 915 688
rect 1279 687 1283 691
rect 2407 687 2411 691
rect 1303 680 1307 684
rect 1343 680 1347 684
rect 1407 680 1411 684
rect 1487 680 1491 684
rect 1575 680 1579 684
rect 1663 680 1667 684
rect 1751 680 1755 684
rect 1831 680 1835 684
rect 1911 680 1915 684
rect 1991 680 1995 684
rect 2079 680 2083 684
rect 2175 680 2179 684
rect 2279 680 2283 684
rect 2359 680 2363 684
rect 135 668 139 672
rect 199 668 203 672
rect 279 668 283 672
rect 351 668 355 672
rect 415 668 419 672
rect 487 668 491 672
rect 559 668 563 672
rect 639 668 643 672
rect 711 668 715 672
rect 783 668 787 672
rect 855 668 859 672
rect 919 668 923 672
rect 983 668 987 672
rect 1039 668 1043 672
rect 1095 668 1099 672
rect 1151 668 1155 672
rect 1191 668 1195 672
rect 111 661 115 665
rect 1239 661 1243 665
rect 1303 664 1307 668
rect 1399 664 1403 668
rect 1511 664 1515 668
rect 1623 664 1627 668
rect 1727 664 1731 668
rect 1815 664 1819 668
rect 1895 664 1899 668
rect 1975 664 1979 668
rect 2047 664 2051 668
rect 2111 664 2115 668
rect 2175 664 2179 668
rect 2239 664 2243 668
rect 2311 664 2315 668
rect 2359 664 2363 668
rect 1279 657 1283 661
rect 2407 657 2411 661
rect 111 644 115 648
rect 191 647 195 651
rect 223 647 224 651
rect 224 647 227 651
rect 343 647 347 651
rect 407 647 411 651
rect 479 647 483 651
rect 551 647 555 651
rect 615 647 619 651
rect 659 647 663 651
rect 911 647 915 651
rect 975 647 979 651
rect 1023 647 1027 651
rect 1087 647 1091 651
rect 1143 647 1147 651
rect 1179 647 1180 651
rect 1180 647 1183 651
rect 1231 647 1235 651
rect 1239 644 1243 648
rect 1279 640 1283 644
rect 1323 643 1327 647
rect 1503 643 1507 647
rect 1591 643 1595 647
rect 1407 635 1411 639
rect 1887 643 1891 647
rect 1967 643 1971 647
rect 2023 643 2027 647
rect 1823 635 1827 639
rect 2287 643 2291 647
rect 2371 643 2375 647
rect 2407 640 2411 644
rect 135 621 139 625
rect 199 621 203 625
rect 279 621 283 625
rect 351 621 355 625
rect 415 621 419 625
rect 487 621 491 625
rect 559 621 563 625
rect 639 621 643 625
rect 711 621 715 625
rect 783 621 787 625
rect 855 621 859 625
rect 919 621 923 625
rect 983 621 987 625
rect 1039 621 1043 625
rect 1095 621 1099 625
rect 1151 621 1155 625
rect 1191 621 1195 625
rect 1303 617 1307 621
rect 1399 617 1403 621
rect 1511 617 1515 621
rect 1623 617 1627 621
rect 1727 617 1731 621
rect 1815 617 1819 621
rect 1895 617 1899 621
rect 1975 617 1979 621
rect 2047 617 2051 621
rect 2111 617 2115 621
rect 2175 617 2179 621
rect 2239 617 2243 621
rect 2311 617 2315 621
rect 2359 617 2363 621
rect 159 611 163 615
rect 191 611 195 615
rect 287 611 291 615
rect 343 611 347 615
rect 407 611 411 615
rect 479 611 483 615
rect 551 611 555 615
rect 791 611 795 615
rect 903 611 907 615
rect 911 611 915 615
rect 975 611 979 615
rect 1023 611 1027 615
rect 1087 611 1091 615
rect 1143 611 1147 615
rect 1179 611 1183 615
rect 1231 607 1235 611
rect 1407 607 1411 611
rect 1503 607 1507 611
rect 1735 607 1739 611
rect 1823 607 1827 611
rect 1887 607 1891 611
rect 1967 607 1971 611
rect 2247 607 2251 611
rect 2303 607 2307 611
rect 2379 607 2383 611
rect 179 591 183 595
rect 259 591 263 595
rect 287 591 291 595
rect 379 591 383 595
rect 387 591 391 595
rect 475 591 479 595
rect 615 591 619 595
rect 651 591 655 595
rect 803 591 807 595
rect 811 591 815 595
rect 883 591 887 595
rect 947 591 951 595
rect 1003 591 1007 595
rect 1051 591 1055 595
rect 1107 591 1111 595
rect 1163 591 1167 595
rect 1435 591 1439 595
rect 1443 591 1447 595
rect 1483 591 1487 595
rect 1583 591 1587 595
rect 1591 591 1595 595
rect 1635 591 1639 595
rect 1691 591 1695 595
rect 2015 591 2019 595
rect 2023 591 2027 595
rect 2075 591 2079 595
rect 2147 591 2151 595
rect 2295 591 2299 595
rect 2371 591 2375 595
rect 135 583 139 587
rect 191 583 195 587
rect 271 583 275 587
rect 359 583 363 587
rect 447 583 451 587
rect 535 583 539 587
rect 623 583 627 587
rect 703 583 707 587
rect 783 583 787 587
rect 855 583 859 587
rect 919 583 923 587
rect 975 583 979 587
rect 1023 583 1027 587
rect 1079 583 1083 587
rect 1135 583 1139 587
rect 1191 583 1195 587
rect 1415 583 1419 587
rect 1455 583 1459 587
rect 1495 583 1499 587
rect 1543 583 1547 587
rect 1599 583 1603 587
rect 1663 583 1667 587
rect 1727 583 1731 587
rect 1791 583 1795 587
rect 1847 583 1851 587
rect 1911 583 1915 587
rect 1975 583 1979 587
rect 2047 583 2051 587
rect 2119 583 2123 587
rect 2199 583 2203 587
rect 2287 583 2291 587
rect 2359 583 2363 587
rect 111 560 115 564
rect 379 563 383 567
rect 159 555 160 559
rect 160 555 163 559
rect 179 555 183 559
rect 259 555 263 559
rect 387 555 388 559
rect 388 555 391 559
rect 475 555 476 559
rect 476 555 479 559
rect 563 555 564 559
rect 564 555 567 559
rect 651 555 652 559
rect 652 555 655 559
rect 1239 560 1243 564
rect 811 555 812 559
rect 812 555 815 559
rect 883 555 884 559
rect 884 555 887 559
rect 947 555 948 559
rect 948 555 951 559
rect 1003 555 1004 559
rect 1004 555 1007 559
rect 1051 555 1052 559
rect 1052 555 1055 559
rect 1107 555 1108 559
rect 1108 555 1111 559
rect 1163 555 1164 559
rect 1164 555 1167 559
rect 1279 560 1283 564
rect 1435 563 1439 567
rect 1583 567 1587 571
rect 1215 555 1216 559
rect 1216 555 1219 559
rect 1443 555 1444 559
rect 1444 555 1447 559
rect 1483 555 1484 559
rect 1484 555 1487 559
rect 1559 555 1563 559
rect 1635 559 1639 563
rect 1691 555 1692 559
rect 1692 555 1695 559
rect 1895 555 1899 559
rect 2015 563 2019 567
rect 2075 555 2076 559
rect 2076 555 2079 559
rect 2147 555 2148 559
rect 2148 555 2151 559
rect 2407 560 2411 564
rect 2303 555 2307 559
rect 2375 555 2379 559
rect 111 543 115 547
rect 1239 543 1243 547
rect 1279 543 1283 547
rect 2407 543 2411 547
rect 135 536 139 540
rect 191 536 195 540
rect 271 536 275 540
rect 359 536 363 540
rect 447 536 451 540
rect 535 536 539 540
rect 623 536 627 540
rect 703 536 707 540
rect 783 536 787 540
rect 855 536 859 540
rect 919 536 923 540
rect 975 536 979 540
rect 1023 536 1027 540
rect 1079 536 1083 540
rect 1135 536 1139 540
rect 1191 536 1195 540
rect 1415 536 1419 540
rect 1455 536 1459 540
rect 1495 536 1499 540
rect 1543 536 1547 540
rect 1599 536 1603 540
rect 1663 536 1667 540
rect 1727 536 1731 540
rect 1791 536 1795 540
rect 1847 536 1851 540
rect 1911 536 1915 540
rect 1975 536 1979 540
rect 2047 536 2051 540
rect 2119 536 2123 540
rect 2199 536 2203 540
rect 2287 536 2291 540
rect 2359 536 2363 540
rect 1303 524 1307 528
rect 1375 524 1379 528
rect 1479 524 1483 528
rect 1583 524 1587 528
rect 1695 524 1699 528
rect 1799 524 1803 528
rect 1903 524 1907 528
rect 2007 524 2011 528
rect 2103 524 2107 528
rect 2191 524 2195 528
rect 2287 524 2291 528
rect 2359 524 2363 528
rect 135 516 139 520
rect 191 516 195 520
rect 263 516 267 520
rect 335 516 339 520
rect 415 516 419 520
rect 495 516 499 520
rect 575 516 579 520
rect 647 516 651 520
rect 719 516 723 520
rect 783 516 787 520
rect 847 516 851 520
rect 903 516 907 520
rect 959 516 963 520
rect 1023 516 1027 520
rect 1087 516 1091 520
rect 1151 516 1155 520
rect 1191 516 1195 520
rect 1279 517 1283 521
rect 2407 517 2411 521
rect 111 509 115 513
rect 1239 509 1243 513
rect 803 503 807 507
rect 111 492 115 496
rect 255 495 259 499
rect 287 495 288 499
rect 288 495 291 499
rect 343 495 347 499
rect 711 495 715 499
rect 839 495 843 499
rect 895 495 899 499
rect 951 495 955 499
rect 1015 495 1019 499
rect 1279 500 1283 504
rect 1311 503 1315 507
rect 1143 495 1147 499
rect 1179 495 1180 499
rect 1180 495 1183 499
rect 1231 495 1235 499
rect 1239 492 1243 496
rect 1723 503 1724 507
rect 1724 503 1727 507
rect 1731 503 1735 507
rect 1999 503 2003 507
rect 1807 495 1811 499
rect 2183 503 2187 507
rect 2279 503 2283 507
rect 2295 503 2299 507
rect 2367 503 2371 507
rect 2407 500 2411 504
rect 1095 483 1099 487
rect 1303 477 1307 481
rect 1375 477 1379 481
rect 1479 477 1483 481
rect 1583 477 1587 481
rect 1695 477 1699 481
rect 1799 477 1803 481
rect 1903 477 1907 481
rect 2007 477 2011 481
rect 2103 477 2107 481
rect 2191 477 2195 481
rect 2287 477 2291 481
rect 2359 477 2363 481
rect 135 469 139 473
rect 191 469 195 473
rect 263 469 267 473
rect 335 469 339 473
rect 415 469 419 473
rect 495 469 499 473
rect 575 469 579 473
rect 647 469 651 473
rect 719 469 723 473
rect 783 469 787 473
rect 847 469 851 473
rect 903 469 907 473
rect 959 469 963 473
rect 1023 469 1027 473
rect 1087 469 1091 473
rect 1151 469 1155 473
rect 1191 469 1195 473
rect 255 459 259 463
rect 563 463 567 467
rect 1231 467 1235 471
rect 1559 467 1563 471
rect 1731 467 1735 471
rect 1807 467 1811 471
rect 1895 467 1899 471
rect 1999 467 2003 471
rect 2175 467 2179 471
rect 2183 467 2187 471
rect 2279 467 2283 471
rect 2375 467 2379 471
rect 691 459 695 463
rect 711 459 715 463
rect 839 459 843 463
rect 895 459 899 463
rect 951 459 955 463
rect 1015 459 1019 463
rect 1095 459 1099 463
rect 1143 459 1147 463
rect 1179 459 1183 463
rect 211 447 215 451
rect 251 447 255 451
rect 299 447 303 451
rect 343 447 347 451
rect 351 447 355 451
rect 395 447 399 451
rect 459 447 463 451
rect 567 447 571 451
rect 587 447 591 451
rect 699 447 703 451
rect 803 447 807 451
rect 859 447 863 451
rect 1311 451 1315 455
rect 1331 451 1335 455
rect 1427 451 1431 455
rect 1491 451 1495 455
rect 1635 451 1639 455
rect 1715 451 1719 455
rect 1723 451 1727 455
rect 1763 451 1767 455
rect 1843 451 1847 455
rect 1923 451 1927 455
rect 2063 451 2067 455
rect 2083 451 2087 455
rect 2163 451 2167 455
rect 2367 451 2371 455
rect 183 439 187 443
rect 223 439 227 443
rect 263 439 267 443
rect 311 439 315 443
rect 367 439 371 443
rect 431 439 435 443
rect 495 439 499 443
rect 559 439 563 443
rect 615 439 619 443
rect 671 439 675 443
rect 719 439 723 443
rect 775 439 779 443
rect 831 439 835 443
rect 887 439 891 443
rect 1303 443 1307 447
rect 1343 443 1347 447
rect 1399 443 1403 447
rect 1463 443 1467 447
rect 1527 443 1531 447
rect 1591 443 1595 447
rect 1663 443 1667 447
rect 1735 443 1739 447
rect 1815 443 1819 447
rect 1895 443 1899 447
rect 1975 443 1979 447
rect 2055 443 2059 447
rect 2135 443 2139 447
rect 2215 443 2219 447
rect 2295 443 2299 447
rect 2359 443 2363 447
rect 111 416 115 420
rect 691 419 695 423
rect 219 411 223 415
rect 259 411 263 415
rect 351 411 355 415
rect 395 411 396 415
rect 396 411 399 415
rect 459 411 460 415
rect 460 411 463 415
rect 467 411 471 415
rect 587 411 588 415
rect 588 411 591 415
rect 699 411 700 415
rect 700 411 703 415
rect 803 411 804 415
rect 804 411 807 415
rect 859 411 860 415
rect 860 411 863 415
rect 1239 416 1243 420
rect 1279 420 1283 424
rect 1635 423 1639 427
rect 1331 415 1332 419
rect 1332 415 1335 419
rect 1427 415 1428 419
rect 1428 415 1431 419
rect 1491 415 1492 419
rect 1492 415 1495 419
rect 111 399 115 403
rect 1239 399 1243 403
rect 1279 403 1283 407
rect 1455 407 1459 411
rect 1655 415 1659 419
rect 1763 415 1764 419
rect 1764 415 1767 419
rect 1843 415 1844 419
rect 1844 415 1847 419
rect 1923 415 1924 419
rect 1924 415 1927 419
rect 1931 415 1935 419
rect 2083 415 2084 419
rect 2084 415 2087 419
rect 2163 415 2164 419
rect 2164 415 2167 419
rect 2175 415 2179 419
rect 2351 415 2355 419
rect 2407 420 2411 424
rect 2407 403 2411 407
rect 183 392 187 396
rect 223 392 227 396
rect 263 392 267 396
rect 311 392 315 396
rect 367 392 371 396
rect 431 392 435 396
rect 495 392 499 396
rect 559 392 563 396
rect 615 392 619 396
rect 671 392 675 396
rect 719 392 723 396
rect 775 392 779 396
rect 831 392 835 396
rect 887 392 891 396
rect 1303 396 1307 400
rect 1343 396 1347 400
rect 1399 396 1403 400
rect 1463 396 1467 400
rect 1527 396 1531 400
rect 1591 396 1595 400
rect 1663 396 1667 400
rect 1735 396 1739 400
rect 1815 396 1819 400
rect 1895 396 1899 400
rect 1975 396 1979 400
rect 2055 396 2059 400
rect 2135 396 2139 400
rect 2215 396 2219 400
rect 2295 396 2299 400
rect 2359 396 2363 400
rect 135 380 139 384
rect 175 380 179 384
rect 231 380 235 384
rect 287 380 291 384
rect 343 380 347 384
rect 391 380 395 384
rect 439 380 443 384
rect 487 380 491 384
rect 535 380 539 384
rect 583 380 587 384
rect 631 380 635 384
rect 679 380 683 384
rect 727 380 731 384
rect 775 380 779 384
rect 1447 380 1451 384
rect 1487 380 1491 384
rect 1535 380 1539 384
rect 1591 380 1595 384
rect 1663 380 1667 384
rect 1735 380 1739 384
rect 1815 380 1819 384
rect 1895 380 1899 384
rect 1967 380 1971 384
rect 2039 380 2043 384
rect 2111 380 2115 384
rect 2175 380 2179 384
rect 2239 380 2243 384
rect 2303 380 2307 384
rect 2359 380 2363 384
rect 111 373 115 377
rect 567 371 571 375
rect 1239 373 1243 377
rect 1279 373 1283 377
rect 2407 373 2411 377
rect 111 356 115 360
rect 163 359 164 363
rect 164 359 167 363
rect 223 359 227 363
rect 279 359 283 363
rect 299 359 303 363
rect 335 359 339 363
rect 527 359 531 363
rect 575 359 579 363
rect 623 359 627 363
rect 671 359 675 363
rect 719 359 723 363
rect 767 359 771 363
rect 1715 367 1719 371
rect 1239 356 1243 360
rect 1279 356 1283 360
rect 1475 359 1476 363
rect 1476 359 1479 363
rect 1527 359 1531 363
rect 1583 359 1587 363
rect 1599 359 1603 363
rect 1727 359 1731 363
rect 1807 359 1811 363
rect 1823 359 1827 363
rect 2031 359 2035 363
rect 2063 359 2064 363
rect 2064 359 2067 363
rect 1975 351 1979 355
rect 2339 359 2343 363
rect 2407 356 2411 360
rect 135 333 139 337
rect 175 333 179 337
rect 231 333 235 337
rect 287 333 291 337
rect 343 333 347 337
rect 391 333 395 337
rect 439 333 443 337
rect 487 333 491 337
rect 535 333 539 337
rect 583 333 587 337
rect 631 333 635 337
rect 679 333 683 337
rect 727 333 731 337
rect 775 333 779 337
rect 1447 333 1451 337
rect 1487 333 1491 337
rect 1535 333 1539 337
rect 1591 333 1595 337
rect 1663 333 1667 337
rect 1735 333 1739 337
rect 1815 333 1819 337
rect 1895 333 1899 337
rect 1967 333 1971 337
rect 2039 333 2043 337
rect 2111 333 2115 337
rect 2175 333 2179 337
rect 2239 333 2243 337
rect 2303 333 2307 337
rect 2359 333 2363 337
rect 163 323 167 327
rect 223 323 227 327
rect 279 323 283 327
rect 467 323 471 327
rect 279 315 283 319
rect 527 323 531 327
rect 575 323 579 327
rect 623 323 627 327
rect 671 323 675 327
rect 719 323 723 327
rect 767 323 771 327
rect 1455 323 1459 327
rect 1475 323 1479 327
rect 1527 323 1531 327
rect 1583 323 1587 327
rect 1655 323 1659 327
rect 1727 323 1731 327
rect 1807 323 1811 327
rect 1931 323 1935 327
rect 1975 323 1979 327
rect 2031 323 2035 327
rect 2283 323 2287 327
rect 2351 323 2355 327
rect 611 315 615 319
rect 1599 315 1603 319
rect 1823 315 1827 319
rect 155 307 159 311
rect 163 307 167 311
rect 211 307 215 311
rect 335 307 339 311
rect 355 307 359 311
rect 419 307 423 311
rect 475 307 479 311
rect 619 307 623 311
rect 667 307 671 311
rect 715 307 719 311
rect 763 307 767 311
rect 807 307 811 311
rect 815 307 819 311
rect 859 307 863 311
rect 907 307 911 311
rect 1523 307 1527 311
rect 1563 307 1567 311
rect 1603 307 1607 311
rect 1643 307 1647 311
rect 1683 307 1687 311
rect 1723 307 1727 311
rect 1827 307 1831 311
rect 1975 307 1979 311
rect 2091 307 2095 311
rect 2099 307 2103 311
rect 2163 307 2167 311
rect 2219 307 2223 311
rect 2339 307 2343 311
rect 2347 307 2351 311
rect 135 299 139 303
rect 183 299 187 303
rect 255 299 259 303
rect 327 299 331 303
rect 391 299 395 303
rect 447 299 451 303
rect 503 299 507 303
rect 551 299 555 303
rect 591 299 595 303
rect 631 299 635 303
rect 679 299 683 303
rect 727 299 731 303
rect 775 299 779 303
rect 823 299 827 303
rect 871 299 875 303
rect 919 299 923 303
rect 1495 299 1499 303
rect 1535 299 1539 303
rect 1575 299 1579 303
rect 1615 299 1619 303
rect 1655 299 1659 303
rect 1695 299 1699 303
rect 1743 299 1747 303
rect 1799 299 1803 303
rect 1863 299 1867 303
rect 1935 299 1939 303
rect 2007 299 2011 303
rect 2071 299 2075 303
rect 2135 299 2139 303
rect 2191 299 2195 303
rect 2255 299 2259 303
rect 2319 299 2323 303
rect 2359 299 2363 303
rect 111 276 115 280
rect 807 279 811 283
rect 163 271 164 275
rect 164 271 167 275
rect 211 271 212 275
rect 212 271 215 275
rect 279 271 280 275
rect 280 271 283 275
rect 355 271 356 275
rect 356 271 359 275
rect 419 271 420 275
rect 420 271 423 275
rect 475 271 476 275
rect 476 271 479 275
rect 567 271 571 275
rect 611 271 615 275
rect 627 271 631 275
rect 667 271 671 275
rect 715 271 719 275
rect 763 271 767 275
rect 859 271 863 275
rect 907 271 911 275
rect 1239 276 1243 280
rect 1279 276 1283 280
rect 2407 276 2411 280
rect 1523 271 1524 275
rect 1524 271 1527 275
rect 1563 271 1564 275
rect 1564 271 1567 275
rect 1603 271 1604 275
rect 1604 271 1607 275
rect 1643 271 1644 275
rect 1644 271 1647 275
rect 1683 271 1684 275
rect 1684 271 1687 275
rect 1723 271 1724 275
rect 1724 271 1727 275
rect 111 259 115 263
rect 1239 259 1243 263
rect 1279 259 1283 263
rect 1711 263 1715 267
rect 1827 271 1828 275
rect 1828 271 1831 275
rect 1975 271 1979 275
rect 1983 271 1987 275
rect 2099 271 2100 275
rect 2100 271 2103 275
rect 2163 271 2164 275
rect 2164 271 2167 275
rect 2219 271 2220 275
rect 2220 271 2223 275
rect 2283 271 2284 275
rect 2284 271 2287 275
rect 2347 271 2348 275
rect 2348 271 2351 275
rect 2375 271 2379 275
rect 2407 259 2411 263
rect 135 252 139 256
rect 183 252 187 256
rect 255 252 259 256
rect 327 252 331 256
rect 391 252 395 256
rect 447 252 451 256
rect 503 252 507 256
rect 551 252 555 256
rect 591 252 595 256
rect 631 252 635 256
rect 679 252 683 256
rect 727 252 731 256
rect 775 252 779 256
rect 823 252 827 256
rect 871 252 875 256
rect 919 252 923 256
rect 1495 252 1499 256
rect 1535 252 1539 256
rect 1575 252 1579 256
rect 1615 252 1619 256
rect 1655 252 1659 256
rect 1695 252 1699 256
rect 1743 252 1747 256
rect 1799 252 1803 256
rect 1863 252 1867 256
rect 1935 252 1939 256
rect 2007 252 2011 256
rect 2071 252 2075 256
rect 2135 252 2139 256
rect 2191 252 2195 256
rect 2255 252 2259 256
rect 2319 252 2323 256
rect 2359 252 2363 256
rect 135 232 139 236
rect 175 232 179 236
rect 247 232 251 236
rect 327 232 331 236
rect 415 232 419 236
rect 495 232 499 236
rect 575 232 579 236
rect 655 232 659 236
rect 727 232 731 236
rect 791 232 795 236
rect 847 232 851 236
rect 903 232 907 236
rect 959 232 963 236
rect 1023 232 1027 236
rect 1367 236 1371 240
rect 1407 236 1411 240
rect 1447 236 1451 240
rect 1495 236 1499 240
rect 1551 236 1555 240
rect 1607 236 1611 240
rect 1671 236 1675 240
rect 1735 236 1739 240
rect 1807 236 1811 240
rect 1887 236 1891 240
rect 1975 236 1979 240
rect 2071 236 2075 240
rect 2167 236 2171 240
rect 2271 236 2275 240
rect 2359 236 2363 240
rect 111 225 115 229
rect 1239 225 1243 229
rect 1279 229 1283 233
rect 2407 229 2411 233
rect 111 208 115 212
rect 155 211 159 215
rect 171 211 175 215
rect 319 211 323 215
rect 487 211 491 215
rect 519 211 520 215
rect 520 211 523 215
rect 183 203 187 207
rect 423 203 427 207
rect 719 211 723 215
rect 783 211 787 215
rect 815 211 816 215
rect 816 211 819 215
rect 663 203 667 207
rect 943 211 947 215
rect 1015 211 1019 215
rect 855 203 859 207
rect 1239 208 1243 212
rect 1279 212 1283 216
rect 1395 215 1396 219
rect 1396 215 1399 219
rect 1435 215 1436 219
rect 1436 215 1439 219
rect 1511 215 1515 219
rect 1643 215 1647 219
rect 1799 215 1803 219
rect 1879 215 1883 219
rect 1967 215 1971 219
rect 1991 215 1995 219
rect 2091 215 2095 219
rect 2367 215 2371 219
rect 1375 207 1379 211
rect 2407 212 2411 216
rect 135 185 139 189
rect 175 185 179 189
rect 247 185 251 189
rect 327 185 331 189
rect 415 185 419 189
rect 495 185 499 189
rect 575 185 579 189
rect 655 185 659 189
rect 727 185 731 189
rect 791 185 795 189
rect 847 185 851 189
rect 903 185 907 189
rect 959 185 963 189
rect 1023 185 1027 189
rect 1367 189 1371 193
rect 1407 189 1411 193
rect 1447 189 1451 193
rect 1495 189 1499 193
rect 1551 189 1555 193
rect 1607 189 1611 193
rect 1671 189 1675 193
rect 1735 189 1739 193
rect 1807 189 1811 193
rect 1887 189 1891 193
rect 1975 189 1979 193
rect 2071 189 2075 193
rect 2167 189 2171 193
rect 2271 189 2275 193
rect 2359 189 2363 193
rect 163 175 167 179
rect 183 175 187 179
rect 239 175 243 179
rect 319 175 323 179
rect 423 175 427 179
rect 487 175 491 179
rect 567 175 571 179
rect 663 175 667 179
rect 719 175 723 179
rect 783 175 787 179
rect 855 175 859 179
rect 751 167 755 171
rect 943 175 947 179
rect 1015 175 1019 179
rect 1375 179 1379 183
rect 1395 179 1399 183
rect 1435 179 1439 183
rect 1643 179 1647 183
rect 1711 179 1715 183
rect 1743 179 1747 183
rect 1799 179 1803 183
rect 1879 179 1883 183
rect 1967 179 1971 183
rect 2243 179 2247 183
rect 2375 179 2379 183
rect 1991 159 1995 163
rect 1331 151 1335 155
rect 1359 151 1363 155
rect 1399 151 1403 155
rect 1439 151 1443 155
rect 1503 151 1507 155
rect 1511 151 1515 155
rect 1851 151 1855 155
rect 1899 151 1903 155
rect 1947 151 1951 155
rect 1995 151 1999 155
rect 2043 151 2047 155
rect 2091 151 2095 155
rect 2139 151 2143 155
rect 2187 151 2191 155
rect 2307 151 2311 155
rect 2347 151 2351 155
rect 2367 151 2371 155
rect 151 143 155 147
rect 159 143 163 147
rect 203 143 207 147
rect 283 143 287 147
rect 319 143 323 147
rect 363 143 367 147
rect 459 143 463 147
rect 511 143 515 147
rect 519 143 523 147
rect 555 143 559 147
rect 647 143 651 147
rect 707 143 711 147
rect 783 143 787 147
rect 835 143 839 147
rect 875 143 879 147
rect 915 143 919 147
rect 1011 143 1015 147
rect 1059 143 1063 147
rect 1099 143 1103 147
rect 1135 143 1139 147
rect 1179 143 1183 147
rect 1295 143 1299 147
rect 1303 143 1307 147
rect 1343 143 1347 147
rect 1383 143 1387 147
rect 1423 143 1427 147
rect 1463 143 1467 147
rect 1519 143 1523 147
rect 1583 143 1587 147
rect 1647 143 1651 147
rect 1711 143 1715 147
rect 1767 143 1771 147
rect 1823 143 1827 147
rect 1871 143 1875 147
rect 1919 143 1923 147
rect 1967 143 1971 147
rect 2015 143 2019 147
rect 2063 143 2067 147
rect 2111 143 2115 147
rect 2159 143 2163 147
rect 2215 143 2219 147
rect 2271 143 2275 147
rect 2319 143 2323 147
rect 2359 143 2363 147
rect 135 135 139 139
rect 175 135 179 139
rect 215 135 219 139
rect 255 135 259 139
rect 295 135 299 139
rect 335 135 339 139
rect 375 135 379 139
rect 423 135 427 139
rect 471 135 475 139
rect 527 135 531 139
rect 583 135 587 139
rect 631 135 635 139
rect 679 135 683 139
rect 727 135 731 139
rect 767 135 771 139
rect 807 135 811 139
rect 847 135 851 139
rect 887 135 891 139
rect 927 135 931 139
rect 975 135 979 139
rect 1023 135 1027 139
rect 1071 135 1075 139
rect 1111 135 1115 139
rect 1151 135 1155 139
rect 1191 135 1195 139
rect 111 112 115 116
rect 151 115 155 119
rect 159 107 160 111
rect 160 107 163 111
rect 203 107 204 111
rect 204 107 207 111
rect 239 107 240 111
rect 240 107 243 111
rect 283 115 287 119
rect 319 115 323 119
rect 363 115 367 119
rect 511 115 515 119
rect 647 119 651 123
rect 1279 120 1283 124
rect 1359 123 1363 127
rect 459 107 463 111
rect 555 107 556 111
rect 556 107 559 111
rect 707 107 708 111
rect 708 107 711 111
rect 751 107 752 111
rect 752 107 755 111
rect 783 115 787 119
rect 835 115 839 119
rect 875 115 879 119
rect 915 115 919 119
rect 1099 115 1103 119
rect 1135 115 1139 119
rect 1011 107 1015 111
rect 1059 107 1063 111
rect 1179 115 1183 119
rect 1239 112 1243 116
rect 1295 115 1299 119
rect 1339 115 1343 119
rect 1399 123 1403 127
rect 1439 123 1443 127
rect 1503 127 1507 131
rect 2347 123 2351 127
rect 2407 120 2411 124
rect 1851 115 1852 119
rect 1852 115 1855 119
rect 1899 115 1900 119
rect 1900 115 1903 119
rect 1947 115 1948 119
rect 1948 115 1951 119
rect 1995 115 1996 119
rect 1996 115 1999 119
rect 2043 115 2044 119
rect 2044 115 2047 119
rect 2091 115 2092 119
rect 2092 115 2095 119
rect 2139 115 2140 119
rect 2140 115 2143 119
rect 2187 115 2188 119
rect 2188 115 2191 119
rect 2243 115 2244 119
rect 2244 115 2247 119
rect 2307 115 2311 119
rect 1279 103 1283 107
rect 2407 103 2411 107
rect 111 95 115 99
rect 1239 95 1243 99
rect 1303 96 1307 100
rect 1343 96 1347 100
rect 1383 96 1387 100
rect 1423 96 1427 100
rect 1463 96 1467 100
rect 1519 96 1523 100
rect 1583 96 1587 100
rect 1647 96 1651 100
rect 1711 96 1715 100
rect 1767 96 1771 100
rect 1823 96 1827 100
rect 1871 96 1875 100
rect 1919 96 1923 100
rect 1967 96 1971 100
rect 2015 96 2019 100
rect 2063 96 2067 100
rect 2111 96 2115 100
rect 2159 96 2163 100
rect 2215 96 2219 100
rect 2271 96 2275 100
rect 2319 96 2323 100
rect 2359 96 2363 100
rect 135 88 139 92
rect 175 88 179 92
rect 215 88 219 92
rect 255 88 259 92
rect 295 88 299 92
rect 335 88 339 92
rect 375 88 379 92
rect 423 88 427 92
rect 471 88 475 92
rect 527 88 531 92
rect 583 88 587 92
rect 631 88 635 92
rect 679 88 683 92
rect 727 88 731 92
rect 767 88 771 92
rect 807 88 811 92
rect 847 88 851 92
rect 887 88 891 92
rect 927 88 931 92
rect 975 88 979 92
rect 1023 88 1027 92
rect 1071 88 1075 92
rect 1111 88 1115 92
rect 1151 88 1155 92
rect 1191 88 1195 92
<< m3 >>
rect 1279 2514 1283 2515
rect 1279 2509 1283 2510
rect 1535 2514 1539 2515
rect 1535 2509 1539 2510
rect 1575 2514 1579 2515
rect 1575 2509 1579 2510
rect 1615 2514 1619 2515
rect 1615 2509 1619 2510
rect 1655 2514 1659 2515
rect 1655 2509 1659 2510
rect 1695 2514 1699 2515
rect 1695 2509 1699 2510
rect 1735 2514 1739 2515
rect 1735 2509 1739 2510
rect 1775 2514 1779 2515
rect 1775 2509 1779 2510
rect 1815 2514 1819 2515
rect 1815 2509 1819 2510
rect 1855 2514 1859 2515
rect 1855 2509 1859 2510
rect 1895 2514 1899 2515
rect 1895 2509 1899 2510
rect 1935 2514 1939 2515
rect 1935 2509 1939 2510
rect 1975 2514 1979 2515
rect 1975 2509 1979 2510
rect 2407 2514 2411 2515
rect 2407 2509 2411 2510
rect 111 2502 115 2503
rect 111 2497 115 2498
rect 135 2502 139 2503
rect 135 2497 139 2498
rect 175 2502 179 2503
rect 175 2497 179 2498
rect 215 2502 219 2503
rect 215 2497 219 2498
rect 255 2502 259 2503
rect 255 2497 259 2498
rect 311 2502 315 2503
rect 311 2497 315 2498
rect 391 2502 395 2503
rect 391 2497 395 2498
rect 479 2502 483 2503
rect 479 2497 483 2498
rect 567 2502 571 2503
rect 567 2497 571 2498
rect 655 2502 659 2503
rect 655 2497 659 2498
rect 743 2502 747 2503
rect 743 2497 747 2498
rect 831 2502 835 2503
rect 831 2497 835 2498
rect 927 2502 931 2503
rect 927 2497 931 2498
rect 1239 2502 1243 2503
rect 1280 2502 1282 2509
rect 1534 2508 1540 2509
rect 1534 2504 1535 2508
rect 1539 2504 1540 2508
rect 1534 2503 1540 2504
rect 1574 2508 1580 2509
rect 1574 2504 1575 2508
rect 1579 2504 1580 2508
rect 1574 2503 1580 2504
rect 1614 2508 1620 2509
rect 1614 2504 1615 2508
rect 1619 2504 1620 2508
rect 1614 2503 1620 2504
rect 1654 2508 1660 2509
rect 1654 2504 1655 2508
rect 1659 2504 1660 2508
rect 1654 2503 1660 2504
rect 1694 2508 1700 2509
rect 1694 2504 1695 2508
rect 1699 2504 1700 2508
rect 1694 2503 1700 2504
rect 1734 2508 1740 2509
rect 1734 2504 1735 2508
rect 1739 2504 1740 2508
rect 1734 2503 1740 2504
rect 1774 2508 1780 2509
rect 1774 2504 1775 2508
rect 1779 2504 1780 2508
rect 1774 2503 1780 2504
rect 1814 2508 1820 2509
rect 1814 2504 1815 2508
rect 1819 2504 1820 2508
rect 1814 2503 1820 2504
rect 1854 2508 1860 2509
rect 1854 2504 1855 2508
rect 1859 2504 1860 2508
rect 1854 2503 1860 2504
rect 1894 2508 1900 2509
rect 1894 2504 1895 2508
rect 1899 2504 1900 2508
rect 1894 2503 1900 2504
rect 1934 2508 1940 2509
rect 1934 2504 1935 2508
rect 1939 2504 1940 2508
rect 1934 2503 1940 2504
rect 1974 2508 1980 2509
rect 1974 2504 1975 2508
rect 1979 2504 1980 2508
rect 1974 2503 1980 2504
rect 2408 2502 2410 2509
rect 1239 2497 1243 2498
rect 1278 2501 1284 2502
rect 1278 2497 1279 2501
rect 1283 2497 1284 2501
rect 112 2465 114 2497
rect 136 2488 138 2497
rect 158 2495 164 2496
rect 158 2491 159 2495
rect 163 2491 164 2495
rect 158 2490 164 2491
rect 134 2487 140 2488
rect 134 2483 135 2487
rect 139 2483 140 2487
rect 134 2482 140 2483
rect 110 2464 116 2465
rect 110 2460 111 2464
rect 115 2460 116 2464
rect 160 2460 162 2490
rect 176 2488 178 2497
rect 202 2495 208 2496
rect 202 2491 203 2495
rect 207 2491 208 2495
rect 202 2490 208 2491
rect 174 2487 180 2488
rect 174 2483 175 2487
rect 179 2483 180 2487
rect 174 2482 180 2483
rect 204 2460 206 2490
rect 216 2488 218 2497
rect 242 2495 248 2496
rect 242 2491 243 2495
rect 247 2491 248 2495
rect 242 2490 248 2491
rect 214 2487 220 2488
rect 214 2483 215 2487
rect 219 2483 220 2487
rect 214 2482 220 2483
rect 244 2460 246 2490
rect 256 2488 258 2497
rect 282 2495 288 2496
rect 282 2491 283 2495
rect 287 2491 288 2495
rect 282 2490 288 2491
rect 254 2487 260 2488
rect 254 2483 255 2487
rect 259 2483 260 2487
rect 254 2482 260 2483
rect 284 2460 286 2490
rect 312 2488 314 2497
rect 338 2495 344 2496
rect 338 2491 339 2495
rect 343 2491 344 2495
rect 338 2490 344 2491
rect 310 2487 316 2488
rect 310 2483 311 2487
rect 315 2483 316 2487
rect 310 2482 316 2483
rect 340 2460 342 2490
rect 392 2488 394 2497
rect 418 2495 424 2496
rect 418 2491 419 2495
rect 423 2491 424 2495
rect 418 2490 424 2491
rect 390 2487 396 2488
rect 390 2483 391 2487
rect 395 2483 396 2487
rect 390 2482 396 2483
rect 420 2460 422 2490
rect 480 2488 482 2497
rect 506 2495 512 2496
rect 506 2491 507 2495
rect 511 2491 512 2495
rect 506 2490 512 2491
rect 478 2487 484 2488
rect 478 2483 479 2487
rect 483 2483 484 2487
rect 478 2482 484 2483
rect 508 2460 510 2490
rect 568 2488 570 2497
rect 656 2488 658 2497
rect 670 2495 676 2496
rect 670 2491 671 2495
rect 675 2491 676 2495
rect 670 2490 676 2491
rect 682 2495 688 2496
rect 682 2491 683 2495
rect 687 2491 688 2495
rect 682 2490 688 2491
rect 566 2487 572 2488
rect 566 2483 567 2487
rect 571 2483 572 2487
rect 566 2482 572 2483
rect 654 2487 660 2488
rect 654 2483 655 2487
rect 659 2483 660 2487
rect 654 2482 660 2483
rect 110 2459 116 2460
rect 158 2459 164 2460
rect 158 2455 159 2459
rect 163 2455 164 2459
rect 158 2454 164 2455
rect 202 2459 208 2460
rect 202 2455 203 2459
rect 207 2455 208 2459
rect 202 2454 208 2455
rect 242 2459 248 2460
rect 242 2455 243 2459
rect 247 2455 248 2459
rect 242 2454 248 2455
rect 282 2459 288 2460
rect 282 2455 283 2459
rect 287 2455 288 2459
rect 282 2454 288 2455
rect 338 2459 344 2460
rect 338 2455 339 2459
rect 343 2455 344 2459
rect 338 2454 344 2455
rect 418 2459 424 2460
rect 418 2455 419 2459
rect 423 2455 424 2459
rect 418 2454 424 2455
rect 506 2459 512 2460
rect 506 2455 507 2459
rect 511 2455 512 2459
rect 506 2454 512 2455
rect 142 2451 148 2452
rect 110 2447 116 2448
rect 110 2443 111 2447
rect 115 2443 116 2447
rect 142 2447 143 2451
rect 147 2447 148 2451
rect 142 2446 148 2447
rect 110 2442 116 2443
rect 112 2435 114 2442
rect 134 2440 140 2441
rect 134 2436 135 2440
rect 139 2436 140 2440
rect 134 2435 140 2436
rect 111 2434 115 2435
rect 111 2429 115 2430
rect 135 2434 139 2435
rect 135 2429 139 2430
rect 112 2422 114 2429
rect 134 2428 140 2429
rect 134 2424 135 2428
rect 139 2424 140 2428
rect 134 2423 140 2424
rect 110 2421 116 2422
rect 110 2417 111 2421
rect 115 2417 116 2421
rect 110 2416 116 2417
rect 110 2404 116 2405
rect 110 2400 111 2404
rect 115 2400 116 2404
rect 110 2399 116 2400
rect 112 2359 114 2399
rect 134 2381 140 2382
rect 134 2377 135 2381
rect 139 2377 140 2381
rect 134 2376 140 2377
rect 136 2359 138 2376
rect 144 2372 146 2446
rect 174 2440 180 2441
rect 174 2436 175 2440
rect 179 2436 180 2440
rect 174 2435 180 2436
rect 214 2440 220 2441
rect 214 2436 215 2440
rect 219 2436 220 2440
rect 214 2435 220 2436
rect 254 2440 260 2441
rect 254 2436 255 2440
rect 259 2436 260 2440
rect 254 2435 260 2436
rect 310 2440 316 2441
rect 310 2436 311 2440
rect 315 2436 316 2440
rect 310 2435 316 2436
rect 390 2440 396 2441
rect 390 2436 391 2440
rect 395 2436 396 2440
rect 390 2435 396 2436
rect 478 2440 484 2441
rect 478 2436 479 2440
rect 483 2436 484 2440
rect 478 2435 484 2436
rect 566 2440 572 2441
rect 566 2436 567 2440
rect 571 2436 572 2440
rect 566 2435 572 2436
rect 654 2440 660 2441
rect 654 2436 655 2440
rect 659 2436 660 2440
rect 654 2435 660 2436
rect 175 2434 179 2435
rect 175 2429 179 2430
rect 183 2434 187 2435
rect 183 2429 187 2430
rect 215 2434 219 2435
rect 215 2429 219 2430
rect 247 2434 251 2435
rect 247 2429 251 2430
rect 255 2434 259 2435
rect 255 2429 259 2430
rect 311 2434 315 2435
rect 311 2429 315 2430
rect 319 2434 323 2435
rect 319 2429 323 2430
rect 391 2434 395 2435
rect 391 2429 395 2430
rect 471 2434 475 2435
rect 471 2429 475 2430
rect 479 2434 483 2435
rect 479 2429 483 2430
rect 543 2434 547 2435
rect 543 2429 547 2430
rect 567 2434 571 2435
rect 567 2429 571 2430
rect 615 2434 619 2435
rect 615 2429 619 2430
rect 655 2434 659 2435
rect 655 2429 659 2430
rect 182 2428 188 2429
rect 182 2424 183 2428
rect 187 2424 188 2428
rect 182 2423 188 2424
rect 246 2428 252 2429
rect 246 2424 247 2428
rect 251 2424 252 2428
rect 246 2423 252 2424
rect 318 2428 324 2429
rect 318 2424 319 2428
rect 323 2424 324 2428
rect 318 2423 324 2424
rect 390 2428 396 2429
rect 390 2424 391 2428
rect 395 2424 396 2428
rect 390 2423 396 2424
rect 470 2428 476 2429
rect 470 2424 471 2428
rect 475 2424 476 2428
rect 470 2423 476 2424
rect 542 2428 548 2429
rect 542 2424 543 2428
rect 547 2424 548 2428
rect 542 2423 548 2424
rect 614 2428 620 2429
rect 614 2424 615 2428
rect 619 2424 620 2428
rect 614 2423 620 2424
rect 672 2416 674 2490
rect 684 2460 686 2490
rect 744 2488 746 2497
rect 798 2495 804 2496
rect 798 2491 799 2495
rect 803 2491 804 2495
rect 798 2490 804 2491
rect 742 2487 748 2488
rect 742 2483 743 2487
rect 747 2483 748 2487
rect 742 2482 748 2483
rect 800 2460 802 2490
rect 832 2488 834 2497
rect 858 2495 864 2496
rect 858 2491 859 2495
rect 863 2491 864 2495
rect 858 2490 864 2491
rect 830 2487 836 2488
rect 830 2483 831 2487
rect 835 2483 836 2487
rect 830 2482 836 2483
rect 860 2460 862 2490
rect 928 2488 930 2497
rect 926 2487 932 2488
rect 926 2483 927 2487
rect 931 2483 932 2487
rect 926 2482 932 2483
rect 1240 2465 1242 2497
rect 1278 2496 1284 2497
rect 2406 2501 2412 2502
rect 2406 2497 2407 2501
rect 2411 2497 2412 2501
rect 2406 2496 2412 2497
rect 1562 2487 1568 2488
rect 1278 2484 1284 2485
rect 1278 2480 1279 2484
rect 1283 2480 1284 2484
rect 1562 2483 1563 2487
rect 1567 2483 1568 2487
rect 1562 2482 1568 2483
rect 1602 2487 1608 2488
rect 1602 2483 1603 2487
rect 1607 2483 1608 2487
rect 1602 2482 1608 2483
rect 1642 2487 1648 2488
rect 1642 2483 1643 2487
rect 1647 2483 1648 2487
rect 1642 2482 1648 2483
rect 1682 2487 1688 2488
rect 1682 2483 1683 2487
rect 1687 2483 1688 2487
rect 1682 2482 1688 2483
rect 1722 2487 1728 2488
rect 1722 2483 1723 2487
rect 1727 2483 1728 2487
rect 1722 2482 1728 2483
rect 1762 2487 1768 2488
rect 1762 2483 1763 2487
rect 1767 2483 1768 2487
rect 1762 2482 1768 2483
rect 1802 2487 1808 2488
rect 1802 2483 1803 2487
rect 1807 2483 1808 2487
rect 1802 2482 1808 2483
rect 1842 2487 1848 2488
rect 1842 2483 1843 2487
rect 1847 2483 1848 2487
rect 1842 2482 1848 2483
rect 1882 2487 1888 2488
rect 1882 2483 1883 2487
rect 1887 2483 1888 2487
rect 1882 2482 1888 2483
rect 1922 2487 1928 2488
rect 1922 2483 1923 2487
rect 1927 2483 1928 2487
rect 1922 2482 1928 2483
rect 1962 2487 1968 2488
rect 1962 2483 1963 2487
rect 1967 2483 1968 2487
rect 1962 2482 1968 2483
rect 2406 2484 2412 2485
rect 1278 2479 1284 2480
rect 1238 2464 1244 2465
rect 1238 2460 1239 2464
rect 1243 2460 1244 2464
rect 682 2459 688 2460
rect 682 2455 683 2459
rect 687 2455 688 2459
rect 682 2454 688 2455
rect 798 2459 804 2460
rect 798 2455 799 2459
rect 803 2455 804 2459
rect 798 2454 804 2455
rect 858 2459 864 2460
rect 858 2455 859 2459
rect 863 2455 864 2459
rect 858 2454 864 2455
rect 866 2459 872 2460
rect 1238 2459 1244 2460
rect 866 2455 867 2459
rect 871 2455 872 2459
rect 866 2454 872 2455
rect 742 2440 748 2441
rect 742 2436 743 2440
rect 747 2436 748 2440
rect 742 2435 748 2436
rect 830 2440 836 2441
rect 830 2436 831 2440
rect 835 2436 836 2440
rect 830 2435 836 2436
rect 679 2434 683 2435
rect 679 2429 683 2430
rect 735 2434 739 2435
rect 735 2429 739 2430
rect 743 2434 747 2435
rect 743 2429 747 2430
rect 791 2434 795 2435
rect 791 2429 795 2430
rect 831 2434 835 2435
rect 831 2429 835 2430
rect 839 2434 843 2435
rect 839 2429 843 2430
rect 678 2428 684 2429
rect 678 2424 679 2428
rect 683 2424 684 2428
rect 678 2423 684 2424
rect 734 2428 740 2429
rect 734 2424 735 2428
rect 739 2424 740 2428
rect 734 2423 740 2424
rect 790 2428 796 2429
rect 790 2424 791 2428
rect 795 2424 796 2428
rect 790 2423 796 2424
rect 838 2428 844 2429
rect 838 2424 839 2428
rect 843 2424 844 2428
rect 838 2423 844 2424
rect 670 2415 676 2416
rect 670 2411 671 2415
rect 675 2411 676 2415
rect 670 2410 676 2411
rect 174 2407 180 2408
rect 174 2403 175 2407
rect 179 2403 180 2407
rect 174 2402 180 2403
rect 238 2407 244 2408
rect 238 2403 239 2407
rect 243 2403 244 2407
rect 238 2402 244 2403
rect 310 2407 316 2408
rect 310 2403 311 2407
rect 315 2403 316 2407
rect 310 2402 316 2403
rect 382 2407 388 2408
rect 382 2403 383 2407
rect 387 2403 388 2407
rect 382 2402 388 2403
rect 462 2407 468 2408
rect 462 2403 463 2407
rect 467 2403 468 2407
rect 462 2402 468 2403
rect 510 2407 516 2408
rect 510 2403 511 2407
rect 515 2403 516 2407
rect 510 2402 516 2403
rect 606 2407 612 2408
rect 606 2403 607 2407
rect 611 2403 612 2407
rect 606 2402 612 2403
rect 670 2407 676 2408
rect 670 2403 671 2407
rect 675 2403 676 2407
rect 670 2402 676 2403
rect 726 2407 732 2408
rect 726 2403 727 2407
rect 731 2403 732 2407
rect 726 2402 732 2403
rect 782 2407 788 2408
rect 782 2403 783 2407
rect 787 2403 788 2407
rect 782 2402 788 2403
rect 176 2372 178 2402
rect 182 2381 188 2382
rect 182 2377 183 2381
rect 187 2377 188 2381
rect 182 2376 188 2377
rect 142 2371 148 2372
rect 142 2367 143 2371
rect 147 2367 148 2371
rect 142 2366 148 2367
rect 174 2371 180 2372
rect 174 2367 175 2371
rect 179 2367 180 2371
rect 174 2366 180 2367
rect 184 2359 186 2376
rect 240 2372 242 2402
rect 246 2381 252 2382
rect 246 2377 247 2381
rect 251 2377 252 2381
rect 246 2376 252 2377
rect 238 2371 244 2372
rect 238 2367 239 2371
rect 243 2367 244 2371
rect 238 2366 244 2367
rect 248 2359 250 2376
rect 312 2372 314 2402
rect 318 2381 324 2382
rect 318 2377 319 2381
rect 323 2377 324 2381
rect 318 2376 324 2377
rect 310 2371 316 2372
rect 310 2367 311 2371
rect 315 2367 316 2371
rect 310 2366 316 2367
rect 320 2359 322 2376
rect 384 2372 386 2402
rect 390 2381 396 2382
rect 390 2377 391 2381
rect 395 2377 396 2381
rect 390 2376 396 2377
rect 382 2371 388 2372
rect 382 2367 383 2371
rect 387 2367 388 2371
rect 382 2366 388 2367
rect 392 2359 394 2376
rect 464 2372 466 2402
rect 470 2381 476 2382
rect 470 2377 471 2381
rect 475 2377 476 2381
rect 470 2376 476 2377
rect 462 2371 468 2372
rect 462 2367 463 2371
rect 467 2367 468 2371
rect 462 2366 468 2367
rect 472 2359 474 2376
rect 111 2358 115 2359
rect 111 2353 115 2354
rect 135 2358 139 2359
rect 135 2353 139 2354
rect 175 2358 179 2359
rect 175 2353 179 2354
rect 183 2358 187 2359
rect 183 2353 187 2354
rect 215 2358 219 2359
rect 215 2353 219 2354
rect 247 2358 251 2359
rect 247 2353 251 2354
rect 271 2358 275 2359
rect 271 2353 275 2354
rect 319 2358 323 2359
rect 319 2353 323 2354
rect 351 2358 355 2359
rect 351 2353 355 2354
rect 391 2358 395 2359
rect 391 2353 395 2354
rect 431 2358 435 2359
rect 431 2353 435 2354
rect 471 2358 475 2359
rect 471 2353 475 2354
rect 112 2321 114 2353
rect 136 2344 138 2353
rect 154 2351 160 2352
rect 154 2347 155 2351
rect 159 2347 160 2351
rect 154 2346 160 2347
rect 162 2351 168 2352
rect 162 2347 163 2351
rect 167 2347 168 2351
rect 162 2346 168 2347
rect 134 2343 140 2344
rect 134 2339 135 2343
rect 139 2339 140 2343
rect 134 2338 140 2339
rect 156 2324 158 2346
rect 154 2323 160 2324
rect 110 2320 116 2321
rect 110 2316 111 2320
rect 115 2316 116 2320
rect 154 2319 155 2323
rect 159 2319 160 2323
rect 154 2318 160 2319
rect 164 2316 166 2346
rect 176 2344 178 2353
rect 202 2351 208 2352
rect 202 2347 203 2351
rect 207 2347 208 2351
rect 202 2346 208 2347
rect 174 2343 180 2344
rect 174 2339 175 2343
rect 179 2339 180 2343
rect 174 2338 180 2339
rect 204 2316 206 2346
rect 216 2344 218 2353
rect 272 2344 274 2353
rect 352 2344 354 2353
rect 418 2351 424 2352
rect 418 2347 419 2351
rect 423 2347 424 2351
rect 418 2346 424 2347
rect 214 2343 220 2344
rect 214 2339 215 2343
rect 219 2339 220 2343
rect 214 2338 220 2339
rect 270 2343 276 2344
rect 270 2339 271 2343
rect 275 2339 276 2343
rect 270 2338 276 2339
rect 350 2343 356 2344
rect 350 2339 351 2343
rect 355 2339 356 2343
rect 350 2338 356 2339
rect 420 2316 422 2346
rect 432 2344 434 2353
rect 512 2352 514 2402
rect 542 2381 548 2382
rect 542 2377 543 2381
rect 547 2377 548 2381
rect 542 2376 548 2377
rect 544 2359 546 2376
rect 608 2372 610 2402
rect 614 2381 620 2382
rect 614 2377 615 2381
rect 619 2377 620 2381
rect 614 2376 620 2377
rect 590 2371 596 2372
rect 590 2367 591 2371
rect 595 2367 596 2371
rect 590 2366 596 2367
rect 606 2371 612 2372
rect 606 2367 607 2371
rect 611 2367 612 2371
rect 606 2366 612 2367
rect 519 2358 523 2359
rect 519 2353 523 2354
rect 543 2358 547 2359
rect 543 2353 547 2354
rect 502 2351 508 2352
rect 502 2347 503 2351
rect 507 2347 508 2351
rect 502 2346 508 2347
rect 510 2351 516 2352
rect 510 2347 511 2351
rect 515 2347 516 2351
rect 510 2346 516 2347
rect 430 2343 436 2344
rect 430 2339 431 2343
rect 435 2339 436 2343
rect 430 2338 436 2339
rect 504 2316 506 2346
rect 520 2344 522 2353
rect 518 2343 524 2344
rect 518 2339 519 2343
rect 523 2339 524 2343
rect 518 2338 524 2339
rect 592 2316 594 2366
rect 616 2359 618 2376
rect 672 2372 674 2402
rect 678 2381 684 2382
rect 678 2377 679 2381
rect 683 2377 684 2381
rect 678 2376 684 2377
rect 670 2371 676 2372
rect 670 2367 671 2371
rect 675 2367 676 2371
rect 670 2366 676 2367
rect 680 2359 682 2376
rect 728 2372 730 2402
rect 734 2381 740 2382
rect 734 2377 735 2381
rect 739 2377 740 2381
rect 734 2376 740 2377
rect 726 2371 732 2372
rect 726 2367 727 2371
rect 731 2367 732 2371
rect 726 2366 732 2367
rect 736 2359 738 2376
rect 784 2372 786 2402
rect 790 2381 796 2382
rect 790 2377 791 2381
rect 795 2377 796 2381
rect 790 2376 796 2377
rect 838 2381 844 2382
rect 838 2377 839 2381
rect 843 2377 844 2381
rect 838 2376 844 2377
rect 782 2371 788 2372
rect 782 2367 783 2371
rect 787 2367 788 2371
rect 782 2366 788 2367
rect 792 2359 794 2376
rect 840 2359 842 2376
rect 868 2372 870 2454
rect 1238 2447 1244 2448
rect 1280 2447 1282 2479
rect 1534 2461 1540 2462
rect 1534 2457 1535 2461
rect 1539 2457 1540 2461
rect 1534 2456 1540 2457
rect 1536 2447 1538 2456
rect 1564 2452 1566 2482
rect 1574 2461 1580 2462
rect 1574 2457 1575 2461
rect 1579 2457 1580 2461
rect 1574 2456 1580 2457
rect 1604 2456 1606 2482
rect 1614 2461 1620 2462
rect 1614 2457 1615 2461
rect 1619 2457 1620 2461
rect 1614 2456 1620 2457
rect 1554 2451 1560 2452
rect 1554 2447 1555 2451
rect 1559 2447 1560 2451
rect 1238 2443 1239 2447
rect 1243 2443 1244 2447
rect 1238 2442 1244 2443
rect 1279 2446 1283 2447
rect 926 2440 932 2441
rect 926 2436 927 2440
rect 931 2436 932 2440
rect 926 2435 932 2436
rect 1240 2435 1242 2442
rect 1279 2441 1283 2442
rect 1359 2446 1363 2447
rect 1359 2441 1363 2442
rect 1399 2446 1403 2447
rect 1399 2441 1403 2442
rect 1455 2446 1459 2447
rect 1455 2441 1459 2442
rect 1519 2446 1523 2447
rect 1519 2441 1523 2442
rect 1535 2446 1539 2447
rect 1554 2446 1560 2447
rect 1562 2451 1568 2452
rect 1562 2447 1563 2451
rect 1567 2447 1568 2451
rect 1576 2447 1578 2456
rect 1602 2455 1608 2456
rect 1602 2451 1603 2455
rect 1607 2451 1608 2455
rect 1602 2450 1608 2451
rect 1616 2447 1618 2456
rect 1644 2452 1646 2482
rect 1654 2461 1660 2462
rect 1654 2457 1655 2461
rect 1659 2457 1660 2461
rect 1654 2456 1660 2457
rect 1684 2456 1686 2482
rect 1694 2461 1700 2462
rect 1694 2457 1695 2461
rect 1699 2457 1700 2461
rect 1694 2456 1700 2457
rect 1642 2451 1648 2452
rect 1642 2447 1643 2451
rect 1647 2447 1648 2451
rect 1656 2447 1658 2456
rect 1682 2455 1688 2456
rect 1682 2451 1683 2455
rect 1687 2451 1688 2455
rect 1682 2450 1688 2451
rect 1696 2447 1698 2456
rect 1724 2452 1726 2482
rect 1734 2461 1740 2462
rect 1734 2457 1735 2461
rect 1739 2457 1740 2461
rect 1734 2456 1740 2457
rect 1764 2456 1766 2482
rect 1774 2461 1780 2462
rect 1774 2457 1775 2461
rect 1779 2457 1780 2461
rect 1774 2456 1780 2457
rect 1722 2451 1728 2452
rect 1722 2447 1723 2451
rect 1727 2447 1728 2451
rect 1736 2447 1738 2456
rect 1762 2455 1768 2456
rect 1762 2451 1763 2455
rect 1767 2451 1768 2455
rect 1762 2450 1768 2451
rect 1776 2447 1778 2456
rect 1804 2452 1806 2482
rect 1830 2479 1836 2480
rect 1830 2475 1831 2479
rect 1835 2475 1836 2479
rect 1830 2474 1836 2475
rect 1814 2461 1820 2462
rect 1814 2457 1815 2461
rect 1819 2457 1820 2461
rect 1814 2456 1820 2457
rect 1802 2451 1808 2452
rect 1802 2447 1803 2451
rect 1807 2447 1808 2451
rect 1816 2447 1818 2456
rect 1562 2446 1568 2447
rect 1575 2446 1579 2447
rect 1535 2441 1539 2442
rect 887 2434 891 2435
rect 887 2429 891 2430
rect 927 2434 931 2435
rect 927 2429 931 2430
rect 935 2434 939 2435
rect 935 2429 939 2430
rect 991 2434 995 2435
rect 991 2429 995 2430
rect 1047 2434 1051 2435
rect 1047 2429 1051 2430
rect 1239 2434 1243 2435
rect 1239 2429 1243 2430
rect 886 2428 892 2429
rect 886 2424 887 2428
rect 891 2424 892 2428
rect 886 2423 892 2424
rect 934 2428 940 2429
rect 934 2424 935 2428
rect 939 2424 940 2428
rect 934 2423 940 2424
rect 990 2428 996 2429
rect 990 2424 991 2428
rect 995 2424 996 2428
rect 990 2423 996 2424
rect 1046 2428 1052 2429
rect 1046 2424 1047 2428
rect 1051 2424 1052 2428
rect 1046 2423 1052 2424
rect 1240 2422 1242 2429
rect 1238 2421 1244 2422
rect 1238 2417 1239 2421
rect 1243 2417 1244 2421
rect 1238 2416 1244 2417
rect 1280 2409 1282 2441
rect 1360 2432 1362 2441
rect 1378 2439 1384 2440
rect 1378 2435 1379 2439
rect 1383 2435 1384 2439
rect 1378 2434 1384 2435
rect 1386 2439 1392 2440
rect 1386 2435 1387 2439
rect 1391 2435 1392 2439
rect 1386 2434 1392 2435
rect 1358 2431 1364 2432
rect 1358 2427 1359 2431
rect 1363 2427 1364 2431
rect 1358 2426 1364 2427
rect 1278 2408 1284 2409
rect 878 2407 884 2408
rect 878 2403 879 2407
rect 883 2403 884 2407
rect 878 2402 884 2403
rect 926 2407 932 2408
rect 926 2403 927 2407
rect 931 2403 932 2407
rect 926 2402 932 2403
rect 974 2407 980 2408
rect 974 2403 975 2407
rect 979 2403 980 2407
rect 974 2402 980 2403
rect 1038 2407 1044 2408
rect 1038 2403 1039 2407
rect 1043 2403 1044 2407
rect 1038 2402 1044 2403
rect 1054 2407 1060 2408
rect 1054 2403 1055 2407
rect 1059 2403 1060 2407
rect 1054 2402 1060 2403
rect 1238 2404 1244 2405
rect 880 2372 882 2402
rect 886 2381 892 2382
rect 886 2377 887 2381
rect 891 2377 892 2381
rect 886 2376 892 2377
rect 866 2371 872 2372
rect 866 2367 867 2371
rect 871 2367 872 2371
rect 866 2366 872 2367
rect 878 2371 884 2372
rect 878 2367 879 2371
rect 883 2367 884 2371
rect 878 2366 884 2367
rect 888 2359 890 2376
rect 928 2372 930 2402
rect 934 2381 940 2382
rect 934 2377 935 2381
rect 939 2377 940 2381
rect 934 2376 940 2377
rect 926 2371 932 2372
rect 926 2367 927 2371
rect 931 2367 932 2371
rect 926 2366 932 2367
rect 936 2359 938 2376
rect 976 2372 978 2402
rect 990 2381 996 2382
rect 990 2377 991 2381
rect 995 2377 996 2381
rect 990 2376 996 2377
rect 974 2371 980 2372
rect 974 2367 975 2371
rect 979 2367 980 2371
rect 974 2366 980 2367
rect 992 2359 994 2376
rect 1040 2372 1042 2402
rect 1046 2381 1052 2382
rect 1046 2377 1047 2381
rect 1051 2377 1052 2381
rect 1046 2376 1052 2377
rect 1038 2371 1044 2372
rect 1038 2367 1039 2371
rect 1043 2367 1044 2371
rect 1038 2366 1044 2367
rect 1048 2359 1050 2376
rect 1056 2360 1058 2402
rect 1238 2400 1239 2404
rect 1243 2400 1244 2404
rect 1278 2404 1279 2408
rect 1283 2404 1284 2408
rect 1278 2403 1284 2404
rect 1238 2399 1244 2400
rect 1054 2359 1060 2360
rect 1240 2359 1242 2399
rect 1278 2391 1284 2392
rect 1278 2387 1279 2391
rect 1283 2387 1284 2391
rect 1278 2386 1284 2387
rect 1280 2379 1282 2386
rect 1358 2384 1364 2385
rect 1358 2380 1359 2384
rect 1363 2380 1364 2384
rect 1358 2379 1364 2380
rect 1279 2378 1283 2379
rect 1279 2373 1283 2374
rect 1359 2378 1363 2379
rect 1359 2373 1363 2374
rect 1280 2366 1282 2373
rect 1358 2372 1364 2373
rect 1358 2368 1359 2372
rect 1363 2368 1364 2372
rect 1358 2367 1364 2368
rect 1278 2365 1284 2366
rect 1278 2361 1279 2365
rect 1283 2361 1284 2365
rect 1278 2360 1284 2361
rect 599 2358 603 2359
rect 599 2353 603 2354
rect 615 2358 619 2359
rect 615 2353 619 2354
rect 679 2358 683 2359
rect 679 2353 683 2354
rect 735 2358 739 2359
rect 735 2353 739 2354
rect 751 2358 755 2359
rect 751 2353 755 2354
rect 791 2358 795 2359
rect 791 2353 795 2354
rect 823 2358 827 2359
rect 823 2353 827 2354
rect 839 2358 843 2359
rect 839 2353 843 2354
rect 887 2358 891 2359
rect 887 2353 891 2354
rect 935 2358 939 2359
rect 935 2353 939 2354
rect 959 2358 963 2359
rect 959 2353 963 2354
rect 991 2358 995 2359
rect 991 2353 995 2354
rect 1031 2358 1035 2359
rect 1031 2353 1035 2354
rect 1047 2358 1051 2359
rect 1054 2355 1055 2359
rect 1059 2355 1060 2359
rect 1054 2354 1060 2355
rect 1239 2358 1243 2359
rect 1047 2353 1051 2354
rect 1239 2353 1243 2354
rect 600 2344 602 2353
rect 666 2351 672 2352
rect 666 2347 667 2351
rect 671 2347 672 2351
rect 666 2346 672 2347
rect 598 2343 604 2344
rect 598 2339 599 2343
rect 603 2339 604 2343
rect 598 2338 604 2339
rect 668 2316 670 2346
rect 680 2344 682 2353
rect 726 2351 732 2352
rect 726 2347 727 2351
rect 731 2347 732 2351
rect 726 2346 732 2347
rect 678 2343 684 2344
rect 678 2339 679 2343
rect 683 2339 684 2343
rect 678 2338 684 2339
rect 728 2316 730 2346
rect 752 2344 754 2353
rect 782 2351 788 2352
rect 782 2347 783 2351
rect 787 2347 788 2351
rect 782 2346 788 2347
rect 750 2343 756 2344
rect 750 2339 751 2343
rect 755 2339 756 2343
rect 750 2338 756 2339
rect 110 2315 116 2316
rect 162 2315 168 2316
rect 162 2311 163 2315
rect 167 2311 168 2315
rect 162 2310 168 2311
rect 202 2315 208 2316
rect 202 2311 203 2315
rect 207 2311 208 2315
rect 202 2310 208 2311
rect 418 2315 424 2316
rect 418 2311 419 2315
rect 423 2311 424 2315
rect 418 2310 424 2311
rect 502 2315 508 2316
rect 502 2311 503 2315
rect 507 2311 508 2315
rect 502 2310 508 2311
rect 590 2315 596 2316
rect 590 2311 591 2315
rect 595 2311 596 2315
rect 590 2310 596 2311
rect 666 2315 672 2316
rect 666 2311 667 2315
rect 671 2311 672 2315
rect 666 2310 672 2311
rect 726 2315 732 2316
rect 726 2311 727 2315
rect 731 2311 732 2315
rect 726 2310 732 2311
rect 142 2307 148 2308
rect 110 2303 116 2304
rect 110 2299 111 2303
rect 115 2299 116 2303
rect 142 2303 143 2307
rect 147 2303 148 2307
rect 142 2302 148 2303
rect 110 2298 116 2299
rect 112 2287 114 2298
rect 134 2296 140 2297
rect 134 2292 135 2296
rect 139 2292 140 2296
rect 134 2291 140 2292
rect 136 2287 138 2291
rect 111 2286 115 2287
rect 111 2281 115 2282
rect 135 2286 139 2287
rect 135 2281 139 2282
rect 112 2274 114 2281
rect 134 2280 140 2281
rect 134 2276 135 2280
rect 139 2276 140 2280
rect 134 2275 140 2276
rect 110 2273 116 2274
rect 110 2269 111 2273
rect 115 2269 116 2273
rect 110 2268 116 2269
rect 110 2256 116 2257
rect 110 2252 111 2256
rect 115 2252 116 2256
rect 110 2251 116 2252
rect 112 2219 114 2251
rect 134 2233 140 2234
rect 134 2229 135 2233
rect 139 2229 140 2233
rect 134 2228 140 2229
rect 136 2219 138 2228
rect 144 2224 146 2302
rect 174 2296 180 2297
rect 174 2292 175 2296
rect 179 2292 180 2296
rect 174 2291 180 2292
rect 214 2296 220 2297
rect 214 2292 215 2296
rect 219 2292 220 2296
rect 214 2291 220 2292
rect 270 2296 276 2297
rect 270 2292 271 2296
rect 275 2292 276 2296
rect 270 2291 276 2292
rect 350 2296 356 2297
rect 350 2292 351 2296
rect 355 2292 356 2296
rect 350 2291 356 2292
rect 430 2296 436 2297
rect 430 2292 431 2296
rect 435 2292 436 2296
rect 430 2291 436 2292
rect 518 2296 524 2297
rect 518 2292 519 2296
rect 523 2292 524 2296
rect 518 2291 524 2292
rect 598 2296 604 2297
rect 598 2292 599 2296
rect 603 2292 604 2296
rect 598 2291 604 2292
rect 678 2296 684 2297
rect 678 2292 679 2296
rect 683 2292 684 2296
rect 678 2291 684 2292
rect 750 2296 756 2297
rect 750 2292 751 2296
rect 755 2292 756 2296
rect 750 2291 756 2292
rect 176 2287 178 2291
rect 216 2287 218 2291
rect 272 2287 274 2291
rect 352 2287 354 2291
rect 432 2287 434 2291
rect 520 2287 522 2291
rect 600 2287 602 2291
rect 680 2287 682 2291
rect 752 2287 754 2291
rect 175 2286 179 2287
rect 175 2281 179 2282
rect 215 2286 219 2287
rect 215 2281 219 2282
rect 231 2286 235 2287
rect 231 2281 235 2282
rect 271 2286 275 2287
rect 271 2281 275 2282
rect 303 2286 307 2287
rect 303 2281 307 2282
rect 351 2286 355 2287
rect 351 2281 355 2282
rect 375 2286 379 2287
rect 375 2281 379 2282
rect 431 2286 435 2287
rect 431 2281 435 2282
rect 455 2286 459 2287
rect 455 2281 459 2282
rect 519 2286 523 2287
rect 519 2281 523 2282
rect 535 2286 539 2287
rect 535 2281 539 2282
rect 599 2286 603 2287
rect 599 2281 603 2282
rect 615 2286 619 2287
rect 615 2281 619 2282
rect 679 2286 683 2287
rect 679 2281 683 2282
rect 687 2286 691 2287
rect 687 2281 691 2282
rect 751 2286 755 2287
rect 751 2281 755 2282
rect 759 2286 763 2287
rect 759 2281 763 2282
rect 174 2280 180 2281
rect 174 2276 175 2280
rect 179 2276 180 2280
rect 174 2275 180 2276
rect 230 2280 236 2281
rect 230 2276 231 2280
rect 235 2276 236 2280
rect 230 2275 236 2276
rect 302 2280 308 2281
rect 302 2276 303 2280
rect 307 2276 308 2280
rect 302 2275 308 2276
rect 374 2280 380 2281
rect 374 2276 375 2280
rect 379 2276 380 2280
rect 374 2275 380 2276
rect 454 2280 460 2281
rect 454 2276 455 2280
rect 459 2276 460 2280
rect 454 2275 460 2276
rect 534 2280 540 2281
rect 534 2276 535 2280
rect 539 2276 540 2280
rect 534 2275 540 2276
rect 614 2280 620 2281
rect 614 2276 615 2280
rect 619 2276 620 2280
rect 614 2275 620 2276
rect 686 2280 692 2281
rect 686 2276 687 2280
rect 691 2276 692 2280
rect 686 2275 692 2276
rect 758 2280 764 2281
rect 758 2276 759 2280
rect 763 2276 764 2280
rect 758 2275 764 2276
rect 784 2260 786 2346
rect 824 2344 826 2353
rect 850 2351 856 2352
rect 850 2347 851 2351
rect 855 2347 856 2351
rect 850 2346 856 2347
rect 822 2343 828 2344
rect 822 2339 823 2343
rect 827 2339 828 2343
rect 822 2338 828 2339
rect 852 2316 854 2346
rect 888 2344 890 2353
rect 914 2351 920 2352
rect 914 2347 915 2351
rect 919 2347 920 2351
rect 914 2346 920 2347
rect 886 2343 892 2344
rect 886 2339 887 2343
rect 891 2339 892 2343
rect 886 2338 892 2339
rect 916 2316 918 2346
rect 960 2344 962 2353
rect 1032 2344 1034 2353
rect 958 2343 964 2344
rect 958 2339 959 2343
rect 963 2339 964 2343
rect 958 2338 964 2339
rect 1030 2343 1036 2344
rect 1030 2339 1031 2343
rect 1035 2339 1036 2343
rect 1030 2338 1036 2339
rect 1240 2321 1242 2353
rect 1380 2352 1382 2434
rect 1388 2404 1390 2434
rect 1400 2432 1402 2441
rect 1426 2439 1432 2440
rect 1426 2435 1427 2439
rect 1431 2435 1432 2439
rect 1426 2434 1432 2435
rect 1398 2431 1404 2432
rect 1398 2427 1399 2431
rect 1403 2427 1404 2431
rect 1398 2426 1404 2427
rect 1428 2404 1430 2434
rect 1456 2432 1458 2441
rect 1482 2439 1488 2440
rect 1482 2435 1483 2439
rect 1487 2435 1488 2439
rect 1482 2434 1488 2435
rect 1454 2431 1460 2432
rect 1454 2427 1455 2431
rect 1459 2427 1460 2431
rect 1454 2426 1460 2427
rect 1484 2404 1486 2434
rect 1520 2432 1522 2441
rect 1546 2439 1552 2440
rect 1546 2435 1547 2439
rect 1551 2435 1552 2439
rect 1546 2434 1552 2435
rect 1518 2431 1524 2432
rect 1518 2427 1519 2431
rect 1523 2427 1524 2431
rect 1518 2426 1524 2427
rect 1548 2404 1550 2434
rect 1556 2412 1558 2446
rect 1575 2441 1579 2442
rect 1599 2446 1603 2447
rect 1599 2441 1603 2442
rect 1615 2446 1619 2447
rect 1642 2446 1648 2447
rect 1655 2446 1659 2447
rect 1615 2441 1619 2442
rect 1655 2441 1659 2442
rect 1679 2446 1683 2447
rect 1679 2441 1683 2442
rect 1695 2446 1699 2447
rect 1722 2446 1728 2447
rect 1735 2446 1739 2447
rect 1695 2441 1699 2442
rect 1735 2441 1739 2442
rect 1759 2446 1763 2447
rect 1759 2441 1763 2442
rect 1775 2446 1779 2447
rect 1802 2446 1808 2447
rect 1815 2446 1819 2447
rect 1775 2441 1779 2442
rect 1815 2441 1819 2442
rect 1600 2432 1602 2441
rect 1626 2439 1632 2440
rect 1626 2435 1627 2439
rect 1631 2435 1632 2439
rect 1626 2434 1632 2435
rect 1598 2431 1604 2432
rect 1598 2427 1599 2431
rect 1603 2427 1604 2431
rect 1598 2426 1604 2427
rect 1554 2411 1560 2412
rect 1554 2407 1555 2411
rect 1559 2407 1560 2411
rect 1554 2406 1560 2407
rect 1628 2404 1630 2434
rect 1680 2432 1682 2441
rect 1706 2439 1712 2440
rect 1706 2435 1707 2439
rect 1711 2435 1712 2439
rect 1706 2434 1712 2435
rect 1678 2431 1684 2432
rect 1678 2427 1679 2431
rect 1683 2427 1684 2431
rect 1678 2426 1684 2427
rect 1708 2404 1710 2434
rect 1760 2432 1762 2441
rect 1832 2440 1834 2474
rect 1844 2456 1846 2482
rect 1854 2461 1860 2462
rect 1854 2457 1855 2461
rect 1859 2457 1860 2461
rect 1854 2456 1860 2457
rect 1842 2455 1848 2456
rect 1842 2451 1843 2455
rect 1847 2451 1848 2455
rect 1842 2450 1848 2451
rect 1856 2447 1858 2456
rect 1884 2452 1886 2482
rect 1894 2461 1900 2462
rect 1894 2457 1895 2461
rect 1899 2457 1900 2461
rect 1894 2456 1900 2457
rect 1924 2456 1926 2482
rect 1934 2461 1940 2462
rect 1934 2457 1935 2461
rect 1939 2457 1940 2461
rect 1934 2456 1940 2457
rect 1882 2451 1888 2452
rect 1882 2447 1883 2451
rect 1887 2447 1888 2451
rect 1896 2447 1898 2456
rect 1922 2455 1928 2456
rect 1922 2451 1923 2455
rect 1927 2451 1928 2455
rect 1922 2450 1928 2451
rect 1936 2447 1938 2456
rect 1964 2452 1966 2482
rect 2406 2480 2407 2484
rect 2411 2480 2412 2484
rect 2406 2479 2412 2480
rect 1974 2461 1980 2462
rect 1974 2457 1975 2461
rect 1979 2457 1980 2461
rect 1974 2456 1980 2457
rect 1962 2451 1968 2452
rect 1962 2447 1963 2451
rect 1967 2447 1968 2451
rect 1976 2447 1978 2456
rect 2408 2447 2410 2479
rect 1839 2446 1843 2447
rect 1839 2441 1843 2442
rect 1855 2446 1859 2447
rect 1882 2446 1888 2447
rect 1895 2446 1899 2447
rect 1855 2441 1859 2442
rect 1895 2441 1899 2442
rect 1919 2446 1923 2447
rect 1919 2441 1923 2442
rect 1935 2446 1939 2447
rect 1962 2446 1968 2447
rect 1975 2446 1979 2447
rect 1935 2441 1939 2442
rect 1975 2441 1979 2442
rect 1999 2446 2003 2447
rect 1999 2441 2003 2442
rect 2079 2446 2083 2447
rect 2079 2441 2083 2442
rect 2159 2446 2163 2447
rect 2159 2441 2163 2442
rect 2247 2446 2251 2447
rect 2247 2441 2251 2442
rect 2335 2446 2339 2447
rect 2335 2441 2339 2442
rect 2407 2446 2411 2447
rect 2407 2441 2411 2442
rect 1830 2439 1836 2440
rect 1830 2435 1831 2439
rect 1835 2435 1836 2439
rect 1830 2434 1836 2435
rect 1840 2432 1842 2441
rect 1866 2439 1872 2440
rect 1866 2435 1867 2439
rect 1871 2435 1872 2439
rect 1866 2434 1872 2435
rect 1758 2431 1764 2432
rect 1758 2427 1759 2431
rect 1763 2427 1764 2431
rect 1758 2426 1764 2427
rect 1838 2431 1844 2432
rect 1838 2427 1839 2431
rect 1843 2427 1844 2431
rect 1838 2426 1844 2427
rect 1868 2404 1870 2434
rect 1920 2432 1922 2441
rect 1946 2439 1952 2440
rect 1946 2435 1947 2439
rect 1951 2435 1952 2439
rect 1946 2434 1952 2435
rect 1918 2431 1924 2432
rect 1918 2427 1919 2431
rect 1923 2427 1924 2431
rect 1918 2426 1924 2427
rect 1948 2404 1950 2434
rect 2000 2432 2002 2441
rect 2026 2439 2032 2440
rect 2026 2435 2027 2439
rect 2031 2435 2032 2439
rect 2026 2434 2032 2435
rect 1998 2431 2004 2432
rect 1998 2427 1999 2431
rect 2003 2427 2004 2431
rect 1998 2426 2004 2427
rect 2028 2404 2030 2434
rect 2080 2432 2082 2441
rect 2106 2439 2112 2440
rect 2106 2435 2107 2439
rect 2111 2435 2112 2439
rect 2106 2434 2112 2435
rect 2078 2431 2084 2432
rect 2078 2427 2079 2431
rect 2083 2427 2084 2431
rect 2078 2426 2084 2427
rect 2108 2404 2110 2434
rect 2160 2432 2162 2441
rect 2182 2439 2188 2440
rect 2182 2435 2183 2439
rect 2187 2435 2188 2439
rect 2182 2434 2188 2435
rect 2158 2431 2164 2432
rect 2158 2427 2159 2431
rect 2163 2427 2164 2431
rect 2158 2426 2164 2427
rect 2184 2404 2186 2434
rect 2248 2432 2250 2441
rect 2290 2439 2296 2440
rect 2290 2435 2291 2439
rect 2295 2435 2296 2439
rect 2290 2434 2296 2435
rect 2246 2431 2252 2432
rect 2246 2427 2247 2431
rect 2251 2427 2252 2431
rect 2246 2426 2252 2427
rect 1386 2403 1392 2404
rect 1386 2399 1387 2403
rect 1391 2399 1392 2403
rect 1386 2398 1392 2399
rect 1426 2403 1432 2404
rect 1426 2399 1427 2403
rect 1431 2399 1432 2403
rect 1426 2398 1432 2399
rect 1482 2403 1488 2404
rect 1482 2399 1483 2403
rect 1487 2399 1488 2403
rect 1482 2398 1488 2399
rect 1546 2403 1552 2404
rect 1546 2399 1547 2403
rect 1551 2399 1552 2403
rect 1546 2398 1552 2399
rect 1626 2403 1632 2404
rect 1626 2399 1627 2403
rect 1631 2399 1632 2403
rect 1626 2398 1632 2399
rect 1706 2403 1712 2404
rect 1706 2399 1707 2403
rect 1711 2399 1712 2403
rect 1706 2398 1712 2399
rect 1866 2403 1872 2404
rect 1866 2399 1867 2403
rect 1871 2399 1872 2403
rect 1866 2398 1872 2399
rect 1946 2403 1952 2404
rect 1946 2399 1947 2403
rect 1951 2399 1952 2403
rect 1946 2398 1952 2399
rect 2026 2403 2032 2404
rect 2026 2399 2027 2403
rect 2031 2399 2032 2403
rect 2026 2398 2032 2399
rect 2106 2403 2112 2404
rect 2106 2399 2107 2403
rect 2111 2399 2112 2403
rect 2106 2398 2112 2399
rect 2182 2403 2188 2404
rect 2182 2399 2183 2403
rect 2187 2399 2188 2403
rect 2182 2398 2188 2399
rect 1398 2384 1404 2385
rect 1398 2380 1399 2384
rect 1403 2380 1404 2384
rect 1398 2379 1404 2380
rect 1454 2384 1460 2385
rect 1454 2380 1455 2384
rect 1459 2380 1460 2384
rect 1454 2379 1460 2380
rect 1518 2384 1524 2385
rect 1518 2380 1519 2384
rect 1523 2380 1524 2384
rect 1518 2379 1524 2380
rect 1598 2384 1604 2385
rect 1598 2380 1599 2384
rect 1603 2380 1604 2384
rect 1598 2379 1604 2380
rect 1678 2384 1684 2385
rect 1678 2380 1679 2384
rect 1683 2380 1684 2384
rect 1678 2379 1684 2380
rect 1758 2384 1764 2385
rect 1758 2380 1759 2384
rect 1763 2380 1764 2384
rect 1758 2379 1764 2380
rect 1838 2384 1844 2385
rect 1838 2380 1839 2384
rect 1843 2380 1844 2384
rect 1838 2379 1844 2380
rect 1918 2384 1924 2385
rect 1918 2380 1919 2384
rect 1923 2380 1924 2384
rect 1918 2379 1924 2380
rect 1998 2384 2004 2385
rect 1998 2380 1999 2384
rect 2003 2380 2004 2384
rect 1998 2379 2004 2380
rect 2078 2384 2084 2385
rect 2078 2380 2079 2384
rect 2083 2380 2084 2384
rect 2078 2379 2084 2380
rect 2158 2384 2164 2385
rect 2158 2380 2159 2384
rect 2163 2380 2164 2384
rect 2158 2379 2164 2380
rect 2246 2384 2252 2385
rect 2246 2380 2247 2384
rect 2251 2380 2252 2384
rect 2246 2379 2252 2380
rect 1399 2378 1403 2379
rect 1399 2373 1403 2374
rect 1407 2378 1411 2379
rect 1407 2373 1411 2374
rect 1455 2378 1459 2379
rect 1455 2373 1459 2374
rect 1471 2378 1475 2379
rect 1471 2373 1475 2374
rect 1519 2378 1523 2379
rect 1519 2373 1523 2374
rect 1543 2378 1547 2379
rect 1543 2373 1547 2374
rect 1599 2378 1603 2379
rect 1599 2373 1603 2374
rect 1615 2378 1619 2379
rect 1615 2373 1619 2374
rect 1679 2378 1683 2379
rect 1679 2373 1683 2374
rect 1695 2378 1699 2379
rect 1695 2373 1699 2374
rect 1759 2378 1763 2379
rect 1759 2373 1763 2374
rect 1775 2378 1779 2379
rect 1775 2373 1779 2374
rect 1839 2378 1843 2379
rect 1839 2373 1843 2374
rect 1855 2378 1859 2379
rect 1855 2373 1859 2374
rect 1919 2378 1923 2379
rect 1919 2373 1923 2374
rect 1927 2378 1931 2379
rect 1927 2373 1931 2374
rect 1999 2378 2003 2379
rect 1999 2373 2003 2374
rect 2071 2378 2075 2379
rect 2071 2373 2075 2374
rect 2079 2378 2083 2379
rect 2079 2373 2083 2374
rect 2143 2378 2147 2379
rect 2143 2373 2147 2374
rect 2159 2378 2163 2379
rect 2159 2373 2163 2374
rect 2223 2378 2227 2379
rect 2223 2373 2227 2374
rect 2247 2378 2251 2379
rect 2247 2373 2251 2374
rect 1406 2372 1412 2373
rect 1406 2368 1407 2372
rect 1411 2368 1412 2372
rect 1406 2367 1412 2368
rect 1470 2372 1476 2373
rect 1470 2368 1471 2372
rect 1475 2368 1476 2372
rect 1470 2367 1476 2368
rect 1542 2372 1548 2373
rect 1542 2368 1543 2372
rect 1547 2368 1548 2372
rect 1542 2367 1548 2368
rect 1614 2372 1620 2373
rect 1614 2368 1615 2372
rect 1619 2368 1620 2372
rect 1614 2367 1620 2368
rect 1694 2372 1700 2373
rect 1694 2368 1695 2372
rect 1699 2368 1700 2372
rect 1694 2367 1700 2368
rect 1774 2372 1780 2373
rect 1774 2368 1775 2372
rect 1779 2368 1780 2372
rect 1774 2367 1780 2368
rect 1854 2372 1860 2373
rect 1854 2368 1855 2372
rect 1859 2368 1860 2372
rect 1854 2367 1860 2368
rect 1926 2372 1932 2373
rect 1926 2368 1927 2372
rect 1931 2368 1932 2372
rect 1926 2367 1932 2368
rect 1998 2372 2004 2373
rect 1998 2368 1999 2372
rect 2003 2368 2004 2372
rect 1998 2367 2004 2368
rect 2070 2372 2076 2373
rect 2070 2368 2071 2372
rect 2075 2368 2076 2372
rect 2070 2367 2076 2368
rect 2142 2372 2148 2373
rect 2142 2368 2143 2372
rect 2147 2368 2148 2372
rect 2142 2367 2148 2368
rect 2222 2372 2228 2373
rect 2222 2368 2223 2372
rect 2227 2368 2228 2372
rect 2222 2367 2228 2368
rect 2292 2356 2294 2434
rect 2336 2432 2338 2441
rect 2334 2431 2340 2432
rect 2334 2427 2335 2431
rect 2339 2427 2340 2431
rect 2334 2426 2340 2427
rect 2408 2409 2410 2441
rect 2406 2408 2412 2409
rect 2406 2404 2407 2408
rect 2411 2404 2412 2408
rect 2350 2403 2356 2404
rect 2406 2403 2412 2404
rect 2350 2399 2351 2403
rect 2355 2399 2356 2403
rect 2350 2398 2356 2399
rect 2334 2384 2340 2385
rect 2334 2380 2335 2384
rect 2339 2380 2340 2384
rect 2334 2379 2340 2380
rect 2303 2378 2307 2379
rect 2303 2373 2307 2374
rect 2335 2378 2339 2379
rect 2335 2373 2339 2374
rect 2302 2372 2308 2373
rect 2302 2368 2303 2372
rect 2307 2368 2308 2372
rect 2302 2367 2308 2368
rect 2290 2355 2296 2356
rect 1378 2351 1384 2352
rect 1278 2348 1284 2349
rect 1278 2344 1279 2348
rect 1283 2344 1284 2348
rect 1378 2347 1379 2351
rect 1383 2347 1384 2351
rect 1378 2346 1384 2347
rect 1686 2351 1692 2352
rect 1686 2347 1687 2351
rect 1691 2347 1692 2351
rect 1686 2346 1692 2347
rect 1766 2351 1772 2352
rect 1766 2347 1767 2351
rect 1771 2347 1772 2351
rect 1766 2346 1772 2347
rect 2046 2351 2052 2352
rect 2046 2347 2047 2351
rect 2051 2347 2052 2351
rect 2290 2351 2291 2355
rect 2295 2351 2296 2355
rect 2290 2350 2296 2351
rect 2310 2351 2316 2352
rect 2046 2346 2052 2347
rect 2310 2347 2311 2351
rect 2315 2347 2316 2351
rect 2310 2346 2316 2347
rect 1278 2343 1284 2344
rect 1550 2343 1556 2344
rect 1238 2320 1244 2321
rect 1238 2316 1239 2320
rect 1243 2316 1244 2320
rect 850 2315 856 2316
rect 850 2311 851 2315
rect 855 2311 856 2315
rect 850 2310 856 2311
rect 914 2315 920 2316
rect 914 2311 915 2315
rect 919 2311 920 2315
rect 914 2310 920 2311
rect 1002 2315 1008 2316
rect 1238 2315 1244 2316
rect 1002 2311 1003 2315
rect 1007 2311 1008 2315
rect 1002 2310 1008 2311
rect 822 2296 828 2297
rect 822 2292 823 2296
rect 827 2292 828 2296
rect 822 2291 828 2292
rect 886 2296 892 2297
rect 886 2292 887 2296
rect 891 2292 892 2296
rect 886 2291 892 2292
rect 958 2296 964 2297
rect 958 2292 959 2296
rect 963 2292 964 2296
rect 958 2291 964 2292
rect 824 2287 826 2291
rect 888 2287 890 2291
rect 960 2287 962 2291
rect 823 2286 827 2287
rect 823 2281 827 2282
rect 831 2286 835 2287
rect 831 2281 835 2282
rect 887 2286 891 2287
rect 887 2281 891 2282
rect 911 2286 915 2287
rect 911 2281 915 2282
rect 959 2286 963 2287
rect 959 2281 963 2282
rect 991 2286 995 2287
rect 991 2281 995 2282
rect 830 2280 836 2281
rect 830 2276 831 2280
rect 835 2276 836 2280
rect 830 2275 836 2276
rect 910 2280 916 2281
rect 910 2276 911 2280
rect 915 2276 916 2280
rect 910 2275 916 2276
rect 990 2280 996 2281
rect 990 2276 991 2280
rect 995 2276 996 2280
rect 990 2275 996 2276
rect 162 2259 168 2260
rect 162 2255 163 2259
rect 167 2255 168 2259
rect 162 2254 168 2255
rect 214 2259 220 2260
rect 214 2255 215 2259
rect 219 2255 220 2259
rect 214 2254 220 2255
rect 294 2259 300 2260
rect 294 2255 295 2259
rect 299 2255 300 2259
rect 294 2254 300 2255
rect 366 2259 372 2260
rect 366 2255 367 2259
rect 371 2255 372 2259
rect 366 2254 372 2255
rect 446 2259 452 2260
rect 446 2255 447 2259
rect 451 2255 452 2259
rect 446 2254 452 2255
rect 678 2259 684 2260
rect 678 2255 679 2259
rect 683 2255 684 2259
rect 678 2254 684 2255
rect 750 2259 756 2260
rect 750 2255 751 2259
rect 755 2255 756 2259
rect 750 2254 756 2255
rect 782 2259 788 2260
rect 782 2255 783 2259
rect 787 2255 788 2259
rect 782 2254 788 2255
rect 854 2259 860 2260
rect 854 2255 855 2259
rect 859 2255 860 2259
rect 854 2254 860 2255
rect 164 2224 166 2254
rect 174 2233 180 2234
rect 174 2229 175 2233
rect 179 2229 180 2233
rect 174 2228 180 2229
rect 142 2223 148 2224
rect 142 2219 143 2223
rect 147 2219 148 2223
rect 111 2218 115 2219
rect 111 2213 115 2214
rect 135 2218 139 2219
rect 142 2218 148 2219
rect 162 2223 168 2224
rect 162 2219 163 2223
rect 167 2219 168 2223
rect 176 2219 178 2228
rect 216 2224 218 2254
rect 254 2251 260 2252
rect 254 2247 255 2251
rect 259 2247 260 2251
rect 254 2246 260 2247
rect 230 2233 236 2234
rect 230 2229 231 2233
rect 235 2229 236 2233
rect 230 2228 236 2229
rect 214 2223 220 2224
rect 214 2219 215 2223
rect 219 2219 220 2223
rect 232 2219 234 2228
rect 162 2218 168 2219
rect 175 2218 179 2219
rect 214 2218 220 2219
rect 231 2218 235 2219
rect 135 2213 139 2214
rect 175 2213 179 2214
rect 231 2213 235 2214
rect 247 2218 251 2219
rect 247 2213 251 2214
rect 112 2181 114 2213
rect 248 2204 250 2213
rect 256 2212 258 2246
rect 296 2224 298 2254
rect 302 2233 308 2234
rect 302 2229 303 2233
rect 307 2229 308 2233
rect 302 2228 308 2229
rect 294 2223 300 2224
rect 294 2219 295 2223
rect 299 2219 300 2223
rect 304 2219 306 2228
rect 368 2224 370 2254
rect 374 2233 380 2234
rect 374 2229 375 2233
rect 379 2229 380 2233
rect 374 2228 380 2229
rect 366 2223 372 2224
rect 366 2219 367 2223
rect 371 2219 372 2223
rect 376 2219 378 2228
rect 448 2224 450 2254
rect 454 2233 460 2234
rect 454 2229 455 2233
rect 459 2229 460 2233
rect 454 2228 460 2229
rect 534 2233 540 2234
rect 534 2229 535 2233
rect 539 2229 540 2233
rect 534 2228 540 2229
rect 614 2233 620 2234
rect 614 2229 615 2233
rect 619 2229 620 2233
rect 614 2228 620 2229
rect 446 2223 452 2224
rect 446 2219 447 2223
rect 451 2219 452 2223
rect 456 2219 458 2228
rect 536 2219 538 2228
rect 616 2219 618 2228
rect 680 2224 682 2254
rect 686 2233 692 2234
rect 686 2229 687 2233
rect 691 2229 692 2233
rect 686 2228 692 2229
rect 678 2223 684 2224
rect 678 2219 679 2223
rect 683 2219 684 2223
rect 688 2219 690 2228
rect 752 2224 754 2254
rect 758 2233 764 2234
rect 758 2229 759 2233
rect 763 2229 764 2233
rect 758 2228 764 2229
rect 830 2233 836 2234
rect 830 2229 831 2233
rect 835 2229 836 2233
rect 830 2228 836 2229
rect 750 2223 756 2224
rect 750 2219 751 2223
rect 755 2219 756 2223
rect 760 2219 762 2228
rect 832 2219 834 2228
rect 287 2218 291 2219
rect 294 2218 300 2219
rect 303 2218 307 2219
rect 287 2213 291 2214
rect 303 2213 307 2214
rect 327 2218 331 2219
rect 366 2218 372 2219
rect 375 2218 379 2219
rect 327 2213 331 2214
rect 375 2213 379 2214
rect 431 2218 435 2219
rect 446 2218 452 2219
rect 455 2218 459 2219
rect 431 2213 435 2214
rect 455 2213 459 2214
rect 495 2218 499 2219
rect 495 2213 499 2214
rect 535 2218 539 2219
rect 535 2213 539 2214
rect 551 2218 555 2219
rect 551 2213 555 2214
rect 607 2218 611 2219
rect 607 2213 611 2214
rect 615 2218 619 2219
rect 615 2213 619 2214
rect 663 2218 667 2219
rect 678 2218 684 2219
rect 687 2218 691 2219
rect 663 2213 667 2214
rect 687 2213 691 2214
rect 719 2218 723 2219
rect 750 2218 756 2219
rect 759 2218 763 2219
rect 719 2213 723 2214
rect 759 2213 763 2214
rect 783 2218 787 2219
rect 783 2213 787 2214
rect 831 2218 835 2219
rect 831 2213 835 2214
rect 847 2218 851 2219
rect 847 2213 851 2214
rect 254 2211 260 2212
rect 254 2207 255 2211
rect 259 2207 260 2211
rect 254 2206 260 2207
rect 274 2211 280 2212
rect 274 2207 275 2211
rect 279 2207 280 2211
rect 274 2206 280 2207
rect 246 2203 252 2204
rect 246 2199 247 2203
rect 251 2199 252 2203
rect 246 2198 252 2199
rect 110 2180 116 2181
rect 110 2176 111 2180
rect 115 2176 116 2180
rect 276 2176 278 2206
rect 288 2204 290 2213
rect 314 2211 320 2212
rect 314 2207 315 2211
rect 319 2207 320 2211
rect 314 2206 320 2207
rect 286 2203 292 2204
rect 286 2199 287 2203
rect 291 2199 292 2203
rect 286 2198 292 2199
rect 316 2176 318 2206
rect 328 2204 330 2213
rect 350 2211 356 2212
rect 350 2207 351 2211
rect 355 2207 356 2211
rect 350 2206 356 2207
rect 326 2203 332 2204
rect 326 2199 327 2203
rect 331 2199 332 2203
rect 326 2198 332 2199
rect 352 2176 354 2206
rect 376 2204 378 2213
rect 402 2211 408 2212
rect 402 2207 403 2211
rect 407 2207 408 2211
rect 402 2206 408 2207
rect 374 2203 380 2204
rect 374 2199 375 2203
rect 379 2199 380 2203
rect 374 2198 380 2199
rect 404 2176 406 2206
rect 432 2204 434 2213
rect 462 2211 468 2212
rect 462 2207 463 2211
rect 467 2207 468 2211
rect 462 2206 468 2207
rect 430 2203 436 2204
rect 430 2199 431 2203
rect 435 2199 436 2203
rect 430 2198 436 2199
rect 464 2176 466 2206
rect 496 2204 498 2213
rect 552 2204 554 2213
rect 570 2211 576 2212
rect 570 2207 571 2211
rect 575 2207 576 2211
rect 570 2206 576 2207
rect 578 2211 584 2212
rect 578 2207 579 2211
rect 583 2207 584 2211
rect 578 2206 584 2207
rect 494 2203 500 2204
rect 494 2199 495 2203
rect 499 2199 500 2203
rect 494 2198 500 2199
rect 550 2203 556 2204
rect 550 2199 551 2203
rect 555 2199 556 2203
rect 550 2198 556 2199
rect 110 2175 116 2176
rect 274 2175 280 2176
rect 274 2171 275 2175
rect 279 2171 280 2175
rect 274 2170 280 2171
rect 314 2175 320 2176
rect 314 2171 315 2175
rect 319 2171 320 2175
rect 314 2170 320 2171
rect 350 2175 356 2176
rect 350 2171 351 2175
rect 355 2171 356 2175
rect 350 2170 356 2171
rect 402 2175 408 2176
rect 402 2171 403 2175
rect 407 2171 408 2175
rect 402 2170 408 2171
rect 458 2175 466 2176
rect 458 2171 459 2175
rect 463 2172 466 2175
rect 463 2171 464 2172
rect 458 2170 464 2171
rect 390 2167 396 2168
rect 110 2163 116 2164
rect 110 2159 111 2163
rect 115 2159 116 2163
rect 390 2163 391 2167
rect 395 2163 396 2167
rect 390 2162 396 2163
rect 110 2158 116 2159
rect 112 2143 114 2158
rect 246 2156 252 2157
rect 246 2152 247 2156
rect 251 2152 252 2156
rect 246 2151 252 2152
rect 286 2156 292 2157
rect 286 2152 287 2156
rect 291 2152 292 2156
rect 286 2151 292 2152
rect 326 2156 332 2157
rect 326 2152 327 2156
rect 331 2152 332 2156
rect 326 2151 332 2152
rect 374 2156 380 2157
rect 374 2152 375 2156
rect 379 2152 380 2156
rect 374 2151 380 2152
rect 248 2143 250 2151
rect 288 2143 290 2151
rect 328 2143 330 2151
rect 376 2143 378 2151
rect 111 2142 115 2143
rect 111 2137 115 2138
rect 247 2142 251 2143
rect 247 2137 251 2138
rect 287 2142 291 2143
rect 287 2137 291 2138
rect 327 2142 331 2143
rect 327 2137 331 2138
rect 375 2142 379 2143
rect 375 2137 379 2138
rect 383 2142 387 2143
rect 383 2137 387 2138
rect 112 2130 114 2137
rect 382 2136 388 2137
rect 382 2132 383 2136
rect 387 2132 388 2136
rect 382 2131 388 2132
rect 110 2129 116 2130
rect 110 2125 111 2129
rect 115 2125 116 2129
rect 110 2124 116 2125
rect 110 2112 116 2113
rect 110 2108 111 2112
rect 115 2108 116 2112
rect 110 2107 116 2108
rect 112 2075 114 2107
rect 382 2089 388 2090
rect 382 2085 383 2089
rect 387 2085 388 2089
rect 382 2084 388 2085
rect 384 2075 386 2084
rect 392 2080 394 2162
rect 430 2156 436 2157
rect 430 2152 431 2156
rect 435 2152 436 2156
rect 430 2151 436 2152
rect 494 2156 500 2157
rect 494 2152 495 2156
rect 499 2152 500 2156
rect 494 2151 500 2152
rect 550 2156 556 2157
rect 550 2152 551 2156
rect 555 2152 556 2156
rect 550 2151 556 2152
rect 432 2143 434 2151
rect 496 2143 498 2151
rect 552 2143 554 2151
rect 423 2142 427 2143
rect 423 2137 427 2138
rect 431 2142 435 2143
rect 431 2137 435 2138
rect 463 2142 467 2143
rect 463 2137 467 2138
rect 495 2142 499 2143
rect 495 2137 499 2138
rect 503 2142 507 2143
rect 503 2137 507 2138
rect 551 2142 555 2143
rect 551 2137 555 2138
rect 422 2136 428 2137
rect 422 2132 423 2136
rect 427 2132 428 2136
rect 422 2131 428 2132
rect 462 2136 468 2137
rect 462 2132 463 2136
rect 467 2132 468 2136
rect 462 2131 468 2132
rect 502 2136 508 2137
rect 502 2132 503 2136
rect 507 2132 508 2136
rect 502 2131 508 2132
rect 550 2136 556 2137
rect 550 2132 551 2136
rect 555 2132 556 2136
rect 550 2131 556 2132
rect 572 2116 574 2206
rect 580 2176 582 2206
rect 608 2204 610 2213
rect 634 2211 640 2212
rect 634 2207 635 2211
rect 639 2207 640 2211
rect 634 2206 640 2207
rect 606 2203 612 2204
rect 606 2199 607 2203
rect 611 2199 612 2203
rect 606 2198 612 2199
rect 636 2176 638 2206
rect 664 2204 666 2213
rect 720 2204 722 2213
rect 738 2211 744 2212
rect 738 2207 739 2211
rect 743 2207 744 2211
rect 738 2206 744 2207
rect 746 2211 752 2212
rect 746 2207 747 2211
rect 751 2207 752 2211
rect 746 2206 752 2207
rect 662 2203 668 2204
rect 662 2199 663 2203
rect 667 2199 668 2203
rect 662 2198 668 2199
rect 718 2203 724 2204
rect 718 2199 719 2203
rect 723 2199 724 2203
rect 718 2198 724 2199
rect 740 2184 742 2206
rect 738 2183 744 2184
rect 738 2179 739 2183
rect 743 2179 744 2183
rect 738 2178 744 2179
rect 748 2176 750 2206
rect 784 2204 786 2213
rect 848 2204 850 2213
rect 856 2212 858 2254
rect 910 2233 916 2234
rect 910 2229 911 2233
rect 915 2229 916 2233
rect 910 2228 916 2229
rect 990 2233 996 2234
rect 990 2229 991 2233
rect 995 2229 996 2233
rect 990 2228 996 2229
rect 912 2219 914 2228
rect 992 2219 994 2228
rect 1004 2224 1006 2310
rect 1280 2307 1282 2343
rect 1550 2339 1551 2343
rect 1555 2339 1556 2343
rect 1550 2338 1556 2339
rect 1358 2325 1364 2326
rect 1358 2321 1359 2325
rect 1363 2321 1364 2325
rect 1358 2320 1364 2321
rect 1406 2325 1412 2326
rect 1406 2321 1407 2325
rect 1411 2321 1412 2325
rect 1406 2320 1412 2321
rect 1470 2325 1476 2326
rect 1470 2321 1471 2325
rect 1475 2321 1476 2325
rect 1470 2320 1476 2321
rect 1542 2325 1548 2326
rect 1542 2321 1543 2325
rect 1547 2321 1548 2325
rect 1542 2320 1548 2321
rect 1360 2307 1362 2320
rect 1408 2307 1410 2320
rect 1472 2307 1474 2320
rect 1544 2307 1546 2320
rect 1552 2316 1554 2338
rect 1614 2325 1620 2326
rect 1614 2321 1615 2325
rect 1619 2321 1620 2325
rect 1614 2320 1620 2321
rect 1550 2315 1556 2316
rect 1550 2311 1551 2315
rect 1555 2311 1556 2315
rect 1550 2310 1556 2311
rect 1606 2315 1612 2316
rect 1606 2311 1607 2315
rect 1611 2311 1612 2315
rect 1606 2310 1612 2311
rect 1279 2306 1283 2307
rect 1238 2303 1244 2304
rect 1238 2299 1239 2303
rect 1243 2299 1244 2303
rect 1279 2301 1283 2302
rect 1359 2306 1363 2307
rect 1359 2301 1363 2302
rect 1407 2306 1411 2307
rect 1407 2301 1411 2302
rect 1471 2306 1475 2307
rect 1471 2301 1475 2302
rect 1503 2306 1507 2307
rect 1503 2301 1507 2302
rect 1543 2306 1547 2307
rect 1543 2301 1547 2302
rect 1583 2306 1587 2307
rect 1583 2301 1587 2302
rect 1238 2298 1244 2299
rect 1030 2296 1036 2297
rect 1030 2292 1031 2296
rect 1035 2292 1036 2296
rect 1030 2291 1036 2292
rect 1032 2287 1034 2291
rect 1240 2287 1242 2298
rect 1031 2286 1035 2287
rect 1031 2281 1035 2282
rect 1239 2286 1243 2287
rect 1239 2281 1243 2282
rect 1240 2274 1242 2281
rect 1238 2273 1244 2274
rect 1238 2269 1239 2273
rect 1243 2269 1244 2273
rect 1280 2269 1282 2301
rect 1504 2292 1506 2301
rect 1522 2299 1528 2300
rect 1522 2295 1523 2299
rect 1527 2295 1528 2299
rect 1522 2294 1528 2295
rect 1530 2299 1536 2300
rect 1530 2295 1531 2299
rect 1535 2295 1536 2299
rect 1530 2294 1536 2295
rect 1502 2291 1508 2292
rect 1502 2287 1503 2291
rect 1507 2287 1508 2291
rect 1502 2286 1508 2287
rect 1524 2272 1526 2294
rect 1522 2271 1528 2272
rect 1238 2268 1244 2269
rect 1278 2268 1284 2269
rect 1278 2264 1279 2268
rect 1283 2264 1284 2268
rect 1522 2267 1523 2271
rect 1527 2267 1528 2271
rect 1522 2266 1528 2267
rect 1532 2264 1534 2294
rect 1544 2292 1546 2301
rect 1566 2299 1572 2300
rect 1566 2295 1567 2299
rect 1571 2295 1572 2299
rect 1566 2294 1572 2295
rect 1542 2291 1548 2292
rect 1542 2287 1543 2291
rect 1547 2287 1548 2291
rect 1542 2286 1548 2287
rect 1568 2264 1570 2294
rect 1584 2292 1586 2301
rect 1582 2291 1588 2292
rect 1582 2287 1583 2291
rect 1587 2287 1588 2291
rect 1582 2286 1588 2287
rect 1608 2264 1610 2310
rect 1616 2307 1618 2320
rect 1688 2316 1690 2346
rect 1694 2325 1700 2326
rect 1694 2321 1695 2325
rect 1699 2321 1700 2325
rect 1694 2320 1700 2321
rect 1686 2315 1692 2316
rect 1686 2311 1687 2315
rect 1691 2311 1692 2315
rect 1686 2310 1692 2311
rect 1696 2307 1698 2320
rect 1615 2306 1619 2307
rect 1615 2301 1619 2302
rect 1623 2306 1627 2307
rect 1623 2301 1627 2302
rect 1663 2306 1667 2307
rect 1663 2301 1667 2302
rect 1695 2306 1699 2307
rect 1695 2301 1699 2302
rect 1703 2306 1707 2307
rect 1703 2301 1707 2302
rect 1759 2306 1763 2307
rect 1759 2301 1763 2302
rect 1624 2292 1626 2301
rect 1646 2299 1652 2300
rect 1646 2295 1647 2299
rect 1651 2295 1652 2299
rect 1646 2294 1652 2295
rect 1654 2299 1660 2300
rect 1654 2295 1655 2299
rect 1659 2295 1660 2299
rect 1654 2294 1660 2295
rect 1622 2291 1628 2292
rect 1622 2287 1623 2291
rect 1627 2287 1628 2291
rect 1622 2286 1628 2287
rect 1648 2272 1650 2294
rect 1646 2271 1652 2272
rect 1646 2267 1647 2271
rect 1651 2267 1652 2271
rect 1646 2266 1652 2267
rect 1278 2263 1284 2264
rect 1530 2263 1536 2264
rect 1530 2259 1531 2263
rect 1535 2259 1536 2263
rect 1530 2258 1536 2259
rect 1566 2263 1572 2264
rect 1566 2259 1567 2263
rect 1571 2259 1572 2263
rect 1566 2258 1572 2259
rect 1606 2263 1612 2264
rect 1606 2259 1607 2263
rect 1611 2259 1612 2263
rect 1606 2258 1612 2259
rect 1238 2256 1244 2257
rect 1238 2252 1239 2256
rect 1243 2252 1244 2256
rect 1238 2251 1244 2252
rect 1278 2251 1284 2252
rect 1002 2223 1008 2224
rect 1002 2219 1003 2223
rect 1007 2219 1008 2223
rect 1240 2219 1242 2251
rect 1278 2247 1279 2251
rect 1283 2247 1284 2251
rect 1278 2246 1284 2247
rect 1280 2231 1282 2246
rect 1502 2244 1508 2245
rect 1502 2240 1503 2244
rect 1507 2240 1508 2244
rect 1502 2239 1508 2240
rect 1542 2244 1548 2245
rect 1542 2240 1543 2244
rect 1547 2240 1548 2244
rect 1542 2239 1548 2240
rect 1582 2244 1588 2245
rect 1582 2240 1583 2244
rect 1587 2240 1588 2244
rect 1582 2239 1588 2240
rect 1622 2244 1628 2245
rect 1622 2240 1623 2244
rect 1627 2240 1628 2244
rect 1622 2239 1628 2240
rect 1504 2231 1506 2239
rect 1544 2231 1546 2239
rect 1584 2231 1586 2239
rect 1624 2231 1626 2239
rect 1279 2230 1283 2231
rect 1279 2225 1283 2226
rect 1303 2230 1307 2231
rect 1303 2225 1307 2226
rect 1343 2230 1347 2231
rect 1343 2225 1347 2226
rect 1383 2230 1387 2231
rect 1383 2225 1387 2226
rect 1431 2230 1435 2231
rect 1431 2225 1435 2226
rect 1495 2230 1499 2231
rect 1495 2225 1499 2226
rect 1503 2230 1507 2231
rect 1503 2225 1507 2226
rect 1543 2230 1547 2231
rect 1543 2225 1547 2226
rect 1567 2230 1571 2231
rect 1567 2225 1571 2226
rect 1583 2230 1587 2231
rect 1583 2225 1587 2226
rect 1623 2230 1627 2231
rect 1623 2225 1627 2226
rect 1639 2230 1643 2231
rect 1639 2225 1643 2226
rect 911 2218 915 2219
rect 911 2213 915 2214
rect 991 2218 995 2219
rect 1002 2218 1008 2219
rect 1239 2218 1243 2219
rect 1280 2218 1282 2225
rect 1302 2224 1308 2225
rect 1302 2220 1303 2224
rect 1307 2220 1308 2224
rect 1302 2219 1308 2220
rect 1342 2224 1348 2225
rect 1342 2220 1343 2224
rect 1347 2220 1348 2224
rect 1342 2219 1348 2220
rect 1382 2224 1388 2225
rect 1382 2220 1383 2224
rect 1387 2220 1388 2224
rect 1382 2219 1388 2220
rect 1430 2224 1436 2225
rect 1430 2220 1431 2224
rect 1435 2220 1436 2224
rect 1430 2219 1436 2220
rect 1494 2224 1500 2225
rect 1494 2220 1495 2224
rect 1499 2220 1500 2224
rect 1494 2219 1500 2220
rect 1566 2224 1572 2225
rect 1566 2220 1567 2224
rect 1571 2220 1572 2224
rect 1566 2219 1572 2220
rect 1638 2224 1644 2225
rect 1638 2220 1639 2224
rect 1643 2220 1644 2224
rect 1638 2219 1644 2220
rect 991 2213 995 2214
rect 1239 2213 1243 2214
rect 1278 2217 1284 2218
rect 1278 2213 1279 2217
rect 1283 2213 1284 2217
rect 854 2211 860 2212
rect 854 2207 855 2211
rect 859 2207 860 2211
rect 854 2206 860 2207
rect 874 2211 880 2212
rect 874 2207 875 2211
rect 879 2207 880 2211
rect 874 2206 880 2207
rect 782 2203 788 2204
rect 782 2199 783 2203
rect 787 2199 788 2203
rect 782 2198 788 2199
rect 846 2203 852 2204
rect 846 2199 847 2203
rect 851 2199 852 2203
rect 846 2198 852 2199
rect 876 2176 878 2206
rect 912 2204 914 2213
rect 910 2203 916 2204
rect 910 2199 911 2203
rect 915 2199 916 2203
rect 910 2198 916 2199
rect 1240 2181 1242 2213
rect 1278 2212 1284 2213
rect 1656 2204 1658 2294
rect 1664 2292 1666 2301
rect 1686 2299 1692 2300
rect 1686 2295 1687 2299
rect 1691 2295 1692 2299
rect 1686 2294 1692 2295
rect 1662 2291 1668 2292
rect 1662 2287 1663 2291
rect 1667 2287 1668 2291
rect 1662 2286 1668 2287
rect 1688 2264 1690 2294
rect 1704 2292 1706 2301
rect 1760 2292 1762 2301
rect 1768 2300 1770 2346
rect 1774 2325 1780 2326
rect 1774 2321 1775 2325
rect 1779 2321 1780 2325
rect 1774 2320 1780 2321
rect 1854 2325 1860 2326
rect 1854 2321 1855 2325
rect 1859 2321 1860 2325
rect 1854 2320 1860 2321
rect 1926 2325 1932 2326
rect 1926 2321 1927 2325
rect 1931 2321 1932 2325
rect 1926 2320 1932 2321
rect 1998 2325 2004 2326
rect 1998 2321 1999 2325
rect 2003 2321 2004 2325
rect 1998 2320 2004 2321
rect 1776 2307 1778 2320
rect 1856 2307 1858 2320
rect 1928 2307 1930 2320
rect 2000 2307 2002 2320
rect 2048 2316 2050 2346
rect 2070 2325 2076 2326
rect 2070 2321 2071 2325
rect 2075 2321 2076 2325
rect 2070 2320 2076 2321
rect 2142 2325 2148 2326
rect 2142 2321 2143 2325
rect 2147 2321 2148 2325
rect 2142 2320 2148 2321
rect 2222 2325 2228 2326
rect 2222 2321 2223 2325
rect 2227 2321 2228 2325
rect 2222 2320 2228 2321
rect 2302 2325 2308 2326
rect 2302 2321 2303 2325
rect 2307 2321 2308 2325
rect 2302 2320 2308 2321
rect 2046 2315 2052 2316
rect 2046 2311 2047 2315
rect 2051 2311 2052 2315
rect 2046 2310 2052 2311
rect 2072 2307 2074 2320
rect 2144 2307 2146 2320
rect 2224 2307 2226 2320
rect 2230 2315 2236 2316
rect 2230 2311 2231 2315
rect 2235 2311 2236 2315
rect 2230 2310 2236 2311
rect 1775 2306 1779 2307
rect 1775 2301 1779 2302
rect 1823 2306 1827 2307
rect 1823 2301 1827 2302
rect 1855 2306 1859 2307
rect 1855 2301 1859 2302
rect 1895 2306 1899 2307
rect 1895 2301 1899 2302
rect 1927 2306 1931 2307
rect 1927 2301 1931 2302
rect 1967 2306 1971 2307
rect 1967 2301 1971 2302
rect 1999 2306 2003 2307
rect 1999 2301 2003 2302
rect 2047 2306 2051 2307
rect 2047 2301 2051 2302
rect 2071 2306 2075 2307
rect 2071 2301 2075 2302
rect 2127 2306 2131 2307
rect 2127 2301 2131 2302
rect 2143 2306 2147 2307
rect 2143 2301 2147 2302
rect 2207 2306 2211 2307
rect 2207 2301 2211 2302
rect 2223 2306 2227 2307
rect 2223 2301 2227 2302
rect 1766 2299 1772 2300
rect 1766 2295 1767 2299
rect 1771 2295 1772 2299
rect 1766 2294 1772 2295
rect 1786 2299 1792 2300
rect 1786 2295 1787 2299
rect 1791 2295 1792 2299
rect 1786 2294 1792 2295
rect 1702 2291 1708 2292
rect 1702 2287 1703 2291
rect 1707 2287 1708 2291
rect 1702 2286 1708 2287
rect 1758 2291 1764 2292
rect 1758 2287 1759 2291
rect 1763 2287 1764 2291
rect 1758 2286 1764 2287
rect 1788 2264 1790 2294
rect 1824 2292 1826 2301
rect 1896 2292 1898 2301
rect 1968 2292 1970 2301
rect 2018 2299 2024 2300
rect 2018 2295 2019 2299
rect 2023 2295 2024 2299
rect 2018 2294 2024 2295
rect 1822 2291 1828 2292
rect 1822 2287 1823 2291
rect 1827 2287 1828 2291
rect 1822 2286 1828 2287
rect 1894 2291 1900 2292
rect 1894 2287 1895 2291
rect 1899 2287 1900 2291
rect 1894 2286 1900 2287
rect 1966 2291 1972 2292
rect 1966 2287 1967 2291
rect 1971 2287 1972 2291
rect 1966 2286 1972 2287
rect 2020 2264 2022 2294
rect 2048 2292 2050 2301
rect 2128 2292 2130 2301
rect 2134 2299 2140 2300
rect 2134 2295 2135 2299
rect 2139 2295 2140 2299
rect 2134 2294 2140 2295
rect 2154 2299 2160 2300
rect 2154 2295 2155 2299
rect 2159 2295 2160 2299
rect 2154 2294 2160 2295
rect 2046 2291 2052 2292
rect 2046 2287 2047 2291
rect 2051 2287 2052 2291
rect 2046 2286 2052 2287
rect 2126 2291 2132 2292
rect 2126 2287 2127 2291
rect 2131 2287 2132 2291
rect 2126 2286 2132 2287
rect 1686 2263 1692 2264
rect 1686 2259 1687 2263
rect 1691 2259 1692 2263
rect 1686 2258 1692 2259
rect 1786 2263 1792 2264
rect 1786 2259 1787 2263
rect 1791 2259 1792 2263
rect 1786 2258 1792 2259
rect 2018 2263 2024 2264
rect 2018 2259 2019 2263
rect 2023 2259 2024 2263
rect 2018 2258 2024 2259
rect 1790 2255 1796 2256
rect 1790 2251 1791 2255
rect 1795 2251 1796 2255
rect 1790 2250 1796 2251
rect 1662 2244 1668 2245
rect 1662 2240 1663 2244
rect 1667 2240 1668 2244
rect 1662 2239 1668 2240
rect 1702 2244 1708 2245
rect 1702 2240 1703 2244
rect 1707 2240 1708 2244
rect 1702 2239 1708 2240
rect 1758 2244 1764 2245
rect 1758 2240 1759 2244
rect 1763 2240 1764 2244
rect 1758 2239 1764 2240
rect 1664 2231 1666 2239
rect 1704 2231 1706 2239
rect 1760 2231 1762 2239
rect 1663 2230 1667 2231
rect 1663 2225 1667 2226
rect 1703 2230 1707 2231
rect 1703 2225 1707 2226
rect 1711 2230 1715 2231
rect 1711 2225 1715 2226
rect 1759 2230 1763 2231
rect 1759 2225 1763 2226
rect 1783 2230 1787 2231
rect 1783 2225 1787 2226
rect 1710 2224 1716 2225
rect 1710 2220 1711 2224
rect 1715 2220 1716 2224
rect 1710 2219 1716 2220
rect 1782 2224 1788 2225
rect 1782 2220 1783 2224
rect 1787 2220 1788 2224
rect 1782 2219 1788 2220
rect 1330 2203 1336 2204
rect 1278 2200 1284 2201
rect 1278 2196 1279 2200
rect 1283 2196 1284 2200
rect 1330 2199 1331 2203
rect 1335 2199 1336 2203
rect 1330 2198 1336 2199
rect 1370 2203 1376 2204
rect 1370 2199 1371 2203
rect 1375 2199 1376 2203
rect 1370 2198 1376 2199
rect 1422 2203 1428 2204
rect 1422 2199 1423 2203
rect 1427 2199 1428 2203
rect 1422 2198 1428 2199
rect 1486 2203 1492 2204
rect 1486 2199 1487 2203
rect 1491 2199 1492 2203
rect 1486 2198 1492 2199
rect 1558 2203 1564 2204
rect 1558 2199 1559 2203
rect 1563 2199 1564 2203
rect 1558 2198 1564 2199
rect 1622 2203 1628 2204
rect 1622 2199 1623 2203
rect 1627 2199 1628 2203
rect 1622 2198 1628 2199
rect 1654 2203 1660 2204
rect 1654 2199 1655 2203
rect 1659 2199 1660 2203
rect 1654 2198 1660 2199
rect 1278 2195 1284 2196
rect 1238 2180 1244 2181
rect 1238 2176 1239 2180
rect 1243 2176 1244 2180
rect 578 2175 584 2176
rect 578 2171 579 2175
rect 583 2171 584 2175
rect 578 2170 584 2171
rect 634 2175 640 2176
rect 634 2171 635 2175
rect 639 2171 640 2175
rect 634 2170 640 2171
rect 746 2175 752 2176
rect 746 2171 747 2175
rect 751 2171 752 2175
rect 746 2170 752 2171
rect 806 2175 812 2176
rect 806 2171 807 2175
rect 811 2171 812 2175
rect 806 2170 812 2171
rect 874 2175 880 2176
rect 1238 2175 1244 2176
rect 874 2171 875 2175
rect 879 2171 880 2175
rect 874 2170 880 2171
rect 606 2156 612 2157
rect 606 2152 607 2156
rect 611 2152 612 2156
rect 606 2151 612 2152
rect 662 2156 668 2157
rect 662 2152 663 2156
rect 667 2152 668 2156
rect 662 2151 668 2152
rect 718 2156 724 2157
rect 718 2152 719 2156
rect 723 2152 724 2156
rect 718 2151 724 2152
rect 782 2156 788 2157
rect 782 2152 783 2156
rect 787 2152 788 2156
rect 782 2151 788 2152
rect 608 2143 610 2151
rect 664 2143 666 2151
rect 720 2143 722 2151
rect 784 2143 786 2151
rect 607 2142 611 2143
rect 607 2137 611 2138
rect 663 2142 667 2143
rect 663 2137 667 2138
rect 719 2142 723 2143
rect 719 2137 723 2138
rect 727 2142 731 2143
rect 727 2137 731 2138
rect 783 2142 787 2143
rect 783 2137 787 2138
rect 791 2142 795 2143
rect 791 2137 795 2138
rect 606 2136 612 2137
rect 606 2132 607 2136
rect 611 2132 612 2136
rect 606 2131 612 2132
rect 662 2136 668 2137
rect 662 2132 663 2136
rect 667 2132 668 2136
rect 662 2131 668 2132
rect 726 2136 732 2137
rect 726 2132 727 2136
rect 731 2132 732 2136
rect 726 2131 732 2132
rect 790 2136 796 2137
rect 790 2132 791 2136
rect 795 2132 796 2136
rect 790 2131 796 2132
rect 410 2115 416 2116
rect 410 2111 411 2115
rect 415 2111 416 2115
rect 410 2110 416 2111
rect 450 2115 456 2116
rect 450 2111 451 2115
rect 455 2111 456 2115
rect 450 2110 456 2111
rect 490 2115 496 2116
rect 490 2111 491 2115
rect 495 2111 496 2115
rect 490 2110 496 2111
rect 570 2115 576 2116
rect 570 2111 571 2115
rect 575 2111 576 2115
rect 570 2110 576 2111
rect 750 2115 756 2116
rect 750 2111 751 2115
rect 755 2111 756 2115
rect 750 2110 756 2111
rect 770 2115 776 2116
rect 770 2111 771 2115
rect 775 2111 776 2115
rect 770 2110 776 2111
rect 398 2107 404 2108
rect 398 2103 399 2107
rect 403 2103 404 2107
rect 398 2102 404 2103
rect 390 2079 396 2080
rect 390 2075 391 2079
rect 395 2075 396 2079
rect 111 2074 115 2075
rect 111 2069 115 2070
rect 383 2074 387 2075
rect 390 2074 396 2075
rect 383 2069 387 2070
rect 112 2037 114 2069
rect 384 2060 386 2069
rect 400 2068 402 2102
rect 412 2080 414 2110
rect 422 2089 428 2090
rect 422 2085 423 2089
rect 427 2085 428 2089
rect 422 2084 428 2085
rect 410 2079 416 2080
rect 410 2075 411 2079
rect 415 2075 416 2079
rect 424 2075 426 2084
rect 452 2080 454 2110
rect 462 2089 468 2090
rect 462 2085 463 2089
rect 467 2085 468 2089
rect 462 2084 468 2085
rect 450 2079 456 2080
rect 450 2075 451 2079
rect 455 2075 456 2079
rect 464 2075 466 2084
rect 492 2080 494 2110
rect 502 2089 508 2090
rect 502 2085 503 2089
rect 507 2085 508 2089
rect 502 2084 508 2085
rect 550 2089 556 2090
rect 550 2085 551 2089
rect 555 2085 556 2089
rect 550 2084 556 2085
rect 606 2089 612 2090
rect 606 2085 607 2089
rect 611 2085 612 2089
rect 606 2084 612 2085
rect 662 2089 668 2090
rect 662 2085 663 2089
rect 667 2085 668 2089
rect 662 2084 668 2085
rect 726 2089 732 2090
rect 726 2085 727 2089
rect 731 2085 732 2089
rect 726 2084 732 2085
rect 490 2079 496 2080
rect 490 2075 491 2079
rect 495 2075 496 2079
rect 504 2075 506 2084
rect 552 2075 554 2084
rect 608 2075 610 2084
rect 654 2079 660 2080
rect 654 2075 655 2079
rect 659 2075 660 2079
rect 664 2075 666 2084
rect 728 2075 730 2084
rect 410 2074 416 2075
rect 423 2074 427 2075
rect 450 2074 456 2075
rect 463 2074 467 2075
rect 490 2074 496 2075
rect 503 2074 507 2075
rect 423 2069 427 2070
rect 463 2069 467 2070
rect 503 2069 507 2070
rect 543 2074 547 2075
rect 543 2069 547 2070
rect 551 2074 555 2075
rect 551 2069 555 2070
rect 583 2074 587 2075
rect 583 2069 587 2070
rect 607 2074 611 2075
rect 607 2069 611 2070
rect 631 2074 635 2075
rect 654 2074 660 2075
rect 663 2074 667 2075
rect 631 2069 635 2070
rect 398 2067 404 2068
rect 398 2063 399 2067
rect 403 2063 404 2067
rect 398 2062 404 2063
rect 410 2067 416 2068
rect 410 2063 411 2067
rect 415 2063 416 2067
rect 410 2062 416 2063
rect 382 2059 388 2060
rect 382 2055 383 2059
rect 387 2055 388 2059
rect 382 2054 388 2055
rect 110 2036 116 2037
rect 110 2032 111 2036
rect 115 2032 116 2036
rect 412 2032 414 2062
rect 424 2060 426 2069
rect 446 2067 452 2068
rect 446 2063 447 2067
rect 451 2063 452 2067
rect 446 2062 452 2063
rect 422 2059 428 2060
rect 422 2055 423 2059
rect 427 2055 428 2059
rect 422 2054 428 2055
rect 448 2032 450 2062
rect 464 2060 466 2069
rect 490 2067 496 2068
rect 490 2063 491 2067
rect 495 2063 496 2067
rect 490 2062 496 2063
rect 462 2059 468 2060
rect 462 2055 463 2059
rect 467 2055 468 2059
rect 462 2054 468 2055
rect 492 2032 494 2062
rect 504 2060 506 2069
rect 526 2067 532 2068
rect 526 2063 527 2067
rect 531 2063 532 2067
rect 526 2062 532 2063
rect 502 2059 508 2060
rect 502 2055 503 2059
rect 507 2055 508 2059
rect 502 2054 508 2055
rect 528 2032 530 2062
rect 544 2060 546 2069
rect 570 2067 576 2068
rect 570 2063 571 2067
rect 575 2063 576 2067
rect 570 2062 576 2063
rect 542 2059 548 2060
rect 542 2055 543 2059
rect 547 2055 548 2059
rect 542 2054 548 2055
rect 572 2032 574 2062
rect 584 2060 586 2069
rect 614 2067 620 2068
rect 614 2063 615 2067
rect 619 2063 620 2067
rect 614 2062 620 2063
rect 582 2059 588 2060
rect 582 2055 583 2059
rect 587 2055 588 2059
rect 582 2054 588 2055
rect 616 2032 618 2062
rect 632 2060 634 2069
rect 630 2059 636 2060
rect 630 2055 631 2059
rect 635 2055 636 2059
rect 630 2054 636 2055
rect 656 2032 658 2074
rect 663 2069 667 2070
rect 687 2074 691 2075
rect 687 2069 691 2070
rect 727 2074 731 2075
rect 727 2069 731 2070
rect 743 2074 747 2075
rect 743 2069 747 2070
rect 688 2060 690 2069
rect 744 2060 746 2069
rect 752 2068 754 2110
rect 772 2080 774 2110
rect 790 2089 796 2090
rect 790 2085 791 2089
rect 795 2085 796 2089
rect 790 2084 796 2085
rect 770 2079 776 2080
rect 770 2075 771 2079
rect 775 2075 776 2079
rect 792 2075 794 2084
rect 808 2080 810 2170
rect 1238 2163 1244 2164
rect 1280 2163 1282 2195
rect 1302 2177 1308 2178
rect 1302 2173 1303 2177
rect 1307 2173 1308 2177
rect 1302 2172 1308 2173
rect 1304 2163 1306 2172
rect 1332 2168 1334 2198
rect 1342 2177 1348 2178
rect 1342 2173 1343 2177
rect 1347 2173 1348 2177
rect 1342 2172 1348 2173
rect 1314 2167 1320 2168
rect 1314 2163 1315 2167
rect 1319 2163 1320 2167
rect 1238 2159 1239 2163
rect 1243 2159 1244 2163
rect 1238 2158 1244 2159
rect 1279 2162 1283 2163
rect 846 2156 852 2157
rect 846 2152 847 2156
rect 851 2152 852 2156
rect 846 2151 852 2152
rect 910 2156 916 2157
rect 910 2152 911 2156
rect 915 2152 916 2156
rect 910 2151 916 2152
rect 848 2143 850 2151
rect 912 2143 914 2151
rect 1240 2143 1242 2158
rect 1279 2157 1283 2158
rect 1303 2162 1307 2163
rect 1314 2162 1320 2163
rect 1330 2167 1336 2168
rect 1330 2163 1331 2167
rect 1335 2163 1336 2167
rect 1344 2163 1346 2172
rect 1372 2168 1374 2198
rect 1382 2177 1388 2178
rect 1382 2173 1383 2177
rect 1387 2173 1388 2177
rect 1382 2172 1388 2173
rect 1370 2167 1376 2168
rect 1370 2163 1371 2167
rect 1375 2163 1376 2167
rect 1384 2163 1386 2172
rect 1424 2168 1426 2198
rect 1430 2177 1436 2178
rect 1430 2173 1431 2177
rect 1435 2173 1436 2177
rect 1430 2172 1436 2173
rect 1422 2167 1428 2168
rect 1422 2163 1423 2167
rect 1427 2163 1428 2167
rect 1432 2163 1434 2172
rect 1488 2168 1490 2198
rect 1494 2177 1500 2178
rect 1494 2173 1495 2177
rect 1499 2173 1500 2177
rect 1494 2172 1500 2173
rect 1486 2167 1492 2168
rect 1486 2163 1487 2167
rect 1491 2163 1492 2167
rect 1496 2163 1498 2172
rect 1560 2168 1562 2198
rect 1566 2177 1572 2178
rect 1566 2173 1567 2177
rect 1571 2173 1572 2177
rect 1566 2172 1572 2173
rect 1558 2167 1564 2168
rect 1558 2163 1559 2167
rect 1563 2163 1564 2167
rect 1568 2163 1570 2172
rect 1330 2162 1336 2163
rect 1343 2162 1347 2163
rect 1303 2157 1307 2158
rect 847 2142 851 2143
rect 847 2137 851 2138
rect 855 2142 859 2143
rect 855 2137 859 2138
rect 911 2142 915 2143
rect 911 2137 915 2138
rect 967 2142 971 2143
rect 967 2137 971 2138
rect 1023 2142 1027 2143
rect 1023 2137 1027 2138
rect 1079 2142 1083 2143
rect 1079 2137 1083 2138
rect 1143 2142 1147 2143
rect 1143 2137 1147 2138
rect 1239 2142 1243 2143
rect 1239 2137 1243 2138
rect 854 2136 860 2137
rect 854 2132 855 2136
rect 859 2132 860 2136
rect 854 2131 860 2132
rect 910 2136 916 2137
rect 910 2132 911 2136
rect 915 2132 916 2136
rect 910 2131 916 2132
rect 966 2136 972 2137
rect 966 2132 967 2136
rect 971 2132 972 2136
rect 966 2131 972 2132
rect 1022 2136 1028 2137
rect 1022 2132 1023 2136
rect 1027 2132 1028 2136
rect 1022 2131 1028 2132
rect 1078 2136 1084 2137
rect 1078 2132 1079 2136
rect 1083 2132 1084 2136
rect 1078 2131 1084 2132
rect 1142 2136 1148 2137
rect 1142 2132 1143 2136
rect 1147 2132 1148 2136
rect 1142 2131 1148 2132
rect 1240 2130 1242 2137
rect 1238 2129 1244 2130
rect 1238 2125 1239 2129
rect 1243 2125 1244 2129
rect 1280 2125 1282 2157
rect 1304 2148 1306 2157
rect 1302 2147 1308 2148
rect 1302 2143 1303 2147
rect 1307 2143 1308 2147
rect 1302 2142 1308 2143
rect 1316 2128 1318 2162
rect 1343 2157 1347 2158
rect 1351 2162 1355 2163
rect 1370 2162 1376 2163
rect 1383 2162 1387 2163
rect 1422 2162 1428 2163
rect 1431 2162 1435 2163
rect 1351 2157 1355 2158
rect 1383 2157 1387 2158
rect 1431 2157 1435 2158
rect 1439 2162 1443 2163
rect 1486 2162 1492 2163
rect 1495 2162 1499 2163
rect 1439 2157 1443 2158
rect 1495 2157 1499 2158
rect 1535 2162 1539 2163
rect 1558 2162 1564 2163
rect 1567 2162 1571 2163
rect 1535 2157 1539 2158
rect 1567 2157 1571 2158
rect 1322 2155 1328 2156
rect 1322 2151 1323 2155
rect 1327 2151 1328 2155
rect 1322 2150 1328 2151
rect 1330 2155 1336 2156
rect 1330 2151 1331 2155
rect 1335 2151 1336 2155
rect 1330 2150 1336 2151
rect 1314 2127 1320 2128
rect 1238 2124 1244 2125
rect 1278 2124 1284 2125
rect 1278 2120 1279 2124
rect 1283 2120 1284 2124
rect 1314 2123 1315 2127
rect 1319 2123 1320 2127
rect 1314 2122 1320 2123
rect 1278 2119 1284 2120
rect 894 2115 900 2116
rect 894 2111 895 2115
rect 899 2111 900 2115
rect 894 2110 900 2111
rect 950 2115 956 2116
rect 950 2111 951 2115
rect 955 2111 956 2115
rect 950 2110 956 2111
rect 1006 2115 1012 2116
rect 1006 2111 1007 2115
rect 1011 2111 1012 2115
rect 1006 2110 1012 2111
rect 1062 2115 1068 2116
rect 1062 2111 1063 2115
rect 1067 2111 1068 2115
rect 1062 2110 1068 2111
rect 1134 2115 1140 2116
rect 1134 2111 1135 2115
rect 1139 2111 1140 2115
rect 1134 2110 1140 2111
rect 1150 2115 1156 2116
rect 1150 2111 1151 2115
rect 1155 2111 1156 2115
rect 1150 2110 1156 2111
rect 1238 2112 1244 2113
rect 854 2089 860 2090
rect 854 2085 855 2089
rect 859 2085 860 2089
rect 854 2084 860 2085
rect 806 2079 812 2080
rect 806 2075 807 2079
rect 811 2075 812 2079
rect 856 2075 858 2084
rect 896 2080 898 2110
rect 910 2089 916 2090
rect 910 2085 911 2089
rect 915 2085 916 2089
rect 910 2084 916 2085
rect 886 2079 892 2080
rect 886 2075 887 2079
rect 891 2075 892 2079
rect 770 2074 776 2075
rect 791 2074 795 2075
rect 791 2069 795 2070
rect 799 2074 803 2075
rect 806 2074 812 2075
rect 847 2074 851 2075
rect 799 2069 803 2070
rect 847 2069 851 2070
rect 855 2074 859 2075
rect 886 2074 892 2075
rect 894 2079 900 2080
rect 894 2075 895 2079
rect 899 2075 900 2079
rect 912 2075 914 2084
rect 952 2080 954 2110
rect 966 2089 972 2090
rect 966 2085 967 2089
rect 971 2085 972 2089
rect 966 2084 972 2085
rect 950 2079 956 2080
rect 950 2075 951 2079
rect 955 2075 956 2079
rect 968 2075 970 2084
rect 1008 2080 1010 2110
rect 1022 2089 1028 2090
rect 1022 2085 1023 2089
rect 1027 2085 1028 2089
rect 1022 2084 1028 2085
rect 1006 2079 1012 2080
rect 1006 2075 1007 2079
rect 1011 2075 1012 2079
rect 1024 2075 1026 2084
rect 1064 2080 1066 2110
rect 1078 2089 1084 2090
rect 1078 2085 1079 2089
rect 1083 2085 1084 2089
rect 1078 2084 1084 2085
rect 1062 2079 1068 2080
rect 1062 2075 1063 2079
rect 1067 2075 1068 2079
rect 1080 2075 1082 2084
rect 1136 2080 1138 2110
rect 1142 2089 1148 2090
rect 1142 2085 1143 2089
rect 1147 2085 1148 2089
rect 1142 2084 1148 2085
rect 1134 2079 1140 2080
rect 1134 2075 1135 2079
rect 1139 2075 1140 2079
rect 1144 2075 1146 2084
rect 894 2074 900 2075
rect 903 2074 907 2075
rect 855 2069 859 2070
rect 750 2067 756 2068
rect 750 2063 751 2067
rect 755 2063 756 2067
rect 750 2062 756 2063
rect 782 2067 788 2068
rect 782 2063 783 2067
rect 787 2063 788 2067
rect 782 2062 788 2063
rect 686 2059 692 2060
rect 686 2055 687 2059
rect 691 2055 692 2059
rect 686 2054 692 2055
rect 742 2059 748 2060
rect 742 2055 743 2059
rect 747 2055 748 2059
rect 742 2054 748 2055
rect 110 2031 116 2032
rect 410 2031 416 2032
rect 410 2027 411 2031
rect 415 2027 416 2031
rect 410 2026 416 2027
rect 446 2031 452 2032
rect 446 2027 447 2031
rect 451 2027 452 2031
rect 446 2026 452 2027
rect 490 2031 496 2032
rect 490 2027 491 2031
rect 495 2027 496 2031
rect 490 2026 496 2027
rect 526 2031 532 2032
rect 526 2027 527 2031
rect 531 2027 532 2031
rect 526 2026 532 2027
rect 570 2031 576 2032
rect 570 2027 571 2031
rect 575 2027 576 2031
rect 570 2026 576 2027
rect 610 2031 618 2032
rect 610 2027 611 2031
rect 615 2028 618 2031
rect 654 2031 660 2032
rect 615 2027 616 2028
rect 610 2026 616 2027
rect 654 2027 655 2031
rect 659 2027 660 2031
rect 654 2026 660 2027
rect 110 2019 116 2020
rect 110 2015 111 2019
rect 115 2015 116 2019
rect 110 2014 116 2015
rect 112 1999 114 2014
rect 382 2012 388 2013
rect 382 2008 383 2012
rect 387 2008 388 2012
rect 382 2007 388 2008
rect 422 2012 428 2013
rect 422 2008 423 2012
rect 427 2008 428 2012
rect 422 2007 428 2008
rect 462 2012 468 2013
rect 462 2008 463 2012
rect 467 2008 468 2012
rect 462 2007 468 2008
rect 502 2012 508 2013
rect 502 2008 503 2012
rect 507 2008 508 2012
rect 502 2007 508 2008
rect 542 2012 548 2013
rect 542 2008 543 2012
rect 547 2008 548 2012
rect 542 2007 548 2008
rect 582 2012 588 2013
rect 582 2008 583 2012
rect 587 2008 588 2012
rect 582 2007 588 2008
rect 630 2012 636 2013
rect 630 2008 631 2012
rect 635 2008 636 2012
rect 630 2007 636 2008
rect 686 2012 692 2013
rect 686 2008 687 2012
rect 691 2008 692 2012
rect 686 2007 692 2008
rect 742 2012 748 2013
rect 742 2008 743 2012
rect 747 2008 748 2012
rect 742 2007 748 2008
rect 384 1999 386 2007
rect 424 1999 426 2007
rect 464 1999 466 2007
rect 504 1999 506 2007
rect 544 1999 546 2007
rect 584 1999 586 2007
rect 632 1999 634 2007
rect 688 1999 690 2007
rect 744 1999 746 2007
rect 111 1998 115 1999
rect 111 1993 115 1994
rect 367 1998 371 1999
rect 367 1993 371 1994
rect 383 1998 387 1999
rect 383 1993 387 1994
rect 407 1998 411 1999
rect 407 1993 411 1994
rect 423 1998 427 1999
rect 423 1993 427 1994
rect 455 1998 459 1999
rect 455 1993 459 1994
rect 463 1998 467 1999
rect 463 1993 467 1994
rect 503 1998 507 1999
rect 503 1993 507 1994
rect 511 1998 515 1999
rect 511 1993 515 1994
rect 543 1998 547 1999
rect 543 1993 547 1994
rect 567 1998 571 1999
rect 567 1993 571 1994
rect 583 1998 587 1999
rect 583 1993 587 1994
rect 631 1998 635 1999
rect 631 1993 635 1994
rect 687 1998 691 1999
rect 687 1993 691 1994
rect 695 1998 699 1999
rect 695 1993 699 1994
rect 743 1998 747 1999
rect 743 1993 747 1994
rect 759 1998 763 1999
rect 759 1993 763 1994
rect 112 1986 114 1993
rect 366 1992 372 1993
rect 366 1988 367 1992
rect 371 1988 372 1992
rect 366 1987 372 1988
rect 406 1992 412 1993
rect 406 1988 407 1992
rect 411 1988 412 1992
rect 406 1987 412 1988
rect 454 1992 460 1993
rect 454 1988 455 1992
rect 459 1988 460 1992
rect 454 1987 460 1988
rect 510 1992 516 1993
rect 510 1988 511 1992
rect 515 1988 516 1992
rect 510 1987 516 1988
rect 566 1992 572 1993
rect 566 1988 567 1992
rect 571 1988 572 1992
rect 566 1987 572 1988
rect 630 1992 636 1993
rect 630 1988 631 1992
rect 635 1988 636 1992
rect 630 1987 636 1988
rect 694 1992 700 1993
rect 694 1988 695 1992
rect 699 1988 700 1992
rect 694 1987 700 1988
rect 758 1992 764 1993
rect 758 1988 759 1992
rect 763 1988 764 1992
rect 758 1987 764 1988
rect 110 1985 116 1986
rect 110 1981 111 1985
rect 115 1981 116 1985
rect 110 1980 116 1981
rect 784 1972 786 2062
rect 800 2060 802 2069
rect 826 2067 832 2068
rect 826 2063 827 2067
rect 831 2063 832 2067
rect 826 2062 832 2063
rect 798 2059 804 2060
rect 798 2055 799 2059
rect 803 2055 804 2059
rect 798 2054 804 2055
rect 828 2032 830 2062
rect 848 2060 850 2069
rect 874 2067 880 2068
rect 874 2063 875 2067
rect 879 2063 880 2067
rect 874 2062 880 2063
rect 846 2059 852 2060
rect 846 2055 847 2059
rect 851 2055 852 2059
rect 846 2054 852 2055
rect 876 2032 878 2062
rect 888 2032 890 2074
rect 903 2069 907 2070
rect 911 2074 915 2075
rect 950 2074 956 2075
rect 959 2074 963 2075
rect 911 2069 915 2070
rect 959 2069 963 2070
rect 967 2074 971 2075
rect 1006 2074 1012 2075
rect 1015 2074 1019 2075
rect 967 2069 971 2070
rect 1015 2069 1019 2070
rect 1023 2074 1027 2075
rect 1062 2074 1068 2075
rect 1071 2074 1075 2075
rect 1023 2069 1027 2070
rect 1071 2069 1075 2070
rect 1079 2074 1083 2075
rect 1134 2074 1140 2075
rect 1143 2074 1147 2075
rect 1079 2069 1083 2070
rect 1143 2069 1147 2070
rect 904 2060 906 2069
rect 960 2060 962 2069
rect 1002 2067 1008 2068
rect 1002 2063 1003 2067
rect 1007 2063 1008 2067
rect 1002 2062 1008 2063
rect 902 2059 908 2060
rect 902 2055 903 2059
rect 907 2055 908 2059
rect 902 2054 908 2055
rect 958 2059 964 2060
rect 958 2055 959 2059
rect 963 2055 964 2059
rect 958 2054 964 2055
rect 1004 2032 1006 2062
rect 1016 2060 1018 2069
rect 1058 2067 1064 2068
rect 1058 2063 1059 2067
rect 1063 2063 1064 2067
rect 1058 2062 1064 2063
rect 1014 2059 1020 2060
rect 1014 2055 1015 2059
rect 1019 2055 1020 2059
rect 1014 2054 1020 2055
rect 1060 2032 1062 2062
rect 1072 2060 1074 2069
rect 1152 2068 1154 2110
rect 1238 2108 1239 2112
rect 1243 2108 1244 2112
rect 1238 2107 1244 2108
rect 1278 2107 1284 2108
rect 1240 2075 1242 2107
rect 1278 2103 1279 2107
rect 1283 2103 1284 2107
rect 1278 2102 1284 2103
rect 1280 2091 1282 2102
rect 1302 2100 1308 2101
rect 1302 2096 1303 2100
rect 1307 2096 1308 2100
rect 1302 2095 1308 2096
rect 1304 2091 1306 2095
rect 1279 2090 1283 2091
rect 1279 2085 1283 2086
rect 1303 2090 1307 2091
rect 1303 2085 1307 2086
rect 1280 2078 1282 2085
rect 1302 2084 1308 2085
rect 1302 2080 1303 2084
rect 1307 2080 1308 2084
rect 1302 2079 1308 2080
rect 1278 2077 1284 2078
rect 1239 2074 1243 2075
rect 1278 2073 1279 2077
rect 1283 2073 1284 2077
rect 1278 2072 1284 2073
rect 1239 2069 1243 2070
rect 1150 2067 1156 2068
rect 1150 2063 1151 2067
rect 1155 2063 1156 2067
rect 1150 2062 1156 2063
rect 1070 2059 1076 2060
rect 1070 2055 1071 2059
rect 1075 2055 1076 2059
rect 1070 2054 1076 2055
rect 1240 2037 1242 2069
rect 1324 2064 1326 2150
rect 1332 2120 1334 2150
rect 1352 2148 1354 2157
rect 1440 2148 1442 2157
rect 1522 2155 1528 2156
rect 1522 2151 1523 2155
rect 1527 2151 1528 2155
rect 1522 2150 1528 2151
rect 1350 2147 1356 2148
rect 1350 2143 1351 2147
rect 1355 2143 1356 2147
rect 1350 2142 1356 2143
rect 1438 2147 1444 2148
rect 1438 2143 1439 2147
rect 1443 2143 1444 2147
rect 1438 2142 1444 2143
rect 1524 2120 1526 2150
rect 1536 2148 1538 2157
rect 1624 2156 1626 2198
rect 1638 2177 1644 2178
rect 1638 2173 1639 2177
rect 1643 2173 1644 2177
rect 1638 2172 1644 2173
rect 1710 2177 1716 2178
rect 1710 2173 1711 2177
rect 1715 2173 1716 2177
rect 1710 2172 1716 2173
rect 1782 2177 1788 2178
rect 1782 2173 1783 2177
rect 1787 2173 1788 2177
rect 1782 2172 1788 2173
rect 1640 2163 1642 2172
rect 1712 2163 1714 2172
rect 1750 2167 1756 2168
rect 1750 2163 1751 2167
rect 1755 2163 1756 2167
rect 1784 2163 1786 2172
rect 1792 2168 1794 2250
rect 1822 2244 1828 2245
rect 1822 2240 1823 2244
rect 1827 2240 1828 2244
rect 1822 2239 1828 2240
rect 1894 2244 1900 2245
rect 1894 2240 1895 2244
rect 1899 2240 1900 2244
rect 1894 2239 1900 2240
rect 1966 2244 1972 2245
rect 1966 2240 1967 2244
rect 1971 2240 1972 2244
rect 1966 2239 1972 2240
rect 2046 2244 2052 2245
rect 2046 2240 2047 2244
rect 2051 2240 2052 2244
rect 2046 2239 2052 2240
rect 2126 2244 2132 2245
rect 2126 2240 2127 2244
rect 2131 2240 2132 2244
rect 2126 2239 2132 2240
rect 1824 2231 1826 2239
rect 1896 2231 1898 2239
rect 1968 2231 1970 2239
rect 2048 2231 2050 2239
rect 2128 2231 2130 2239
rect 1823 2230 1827 2231
rect 1823 2225 1827 2226
rect 1855 2230 1859 2231
rect 1855 2225 1859 2226
rect 1895 2230 1899 2231
rect 1895 2225 1899 2226
rect 1935 2230 1939 2231
rect 1935 2225 1939 2226
rect 1967 2230 1971 2231
rect 1967 2225 1971 2226
rect 2015 2230 2019 2231
rect 2015 2225 2019 2226
rect 2047 2230 2051 2231
rect 2047 2225 2051 2226
rect 2095 2230 2099 2231
rect 2095 2225 2099 2226
rect 2127 2230 2131 2231
rect 2127 2225 2131 2226
rect 1854 2224 1860 2225
rect 1854 2220 1855 2224
rect 1859 2220 1860 2224
rect 1854 2219 1860 2220
rect 1934 2224 1940 2225
rect 1934 2220 1935 2224
rect 1939 2220 1940 2224
rect 1934 2219 1940 2220
rect 2014 2224 2020 2225
rect 2014 2220 2015 2224
rect 2019 2220 2020 2224
rect 2014 2219 2020 2220
rect 2094 2224 2100 2225
rect 2094 2220 2095 2224
rect 2099 2220 2100 2224
rect 2094 2219 2100 2220
rect 2136 2204 2138 2294
rect 2156 2264 2158 2294
rect 2208 2292 2210 2301
rect 2206 2291 2212 2292
rect 2206 2287 2207 2291
rect 2211 2287 2212 2291
rect 2206 2286 2212 2287
rect 2232 2264 2234 2310
rect 2304 2307 2306 2320
rect 2295 2306 2299 2307
rect 2295 2301 2299 2302
rect 2303 2306 2307 2307
rect 2303 2301 2307 2302
rect 2296 2292 2298 2301
rect 2312 2300 2314 2346
rect 2352 2316 2354 2398
rect 2406 2391 2412 2392
rect 2406 2387 2407 2391
rect 2411 2387 2412 2391
rect 2406 2386 2412 2387
rect 2408 2379 2410 2386
rect 2359 2378 2363 2379
rect 2359 2373 2363 2374
rect 2407 2378 2411 2379
rect 2407 2373 2411 2374
rect 2358 2372 2364 2373
rect 2358 2368 2359 2372
rect 2363 2368 2364 2372
rect 2358 2367 2364 2368
rect 2408 2366 2410 2373
rect 2406 2365 2412 2366
rect 2406 2361 2407 2365
rect 2411 2361 2412 2365
rect 2406 2360 2412 2361
rect 2406 2348 2412 2349
rect 2406 2344 2407 2348
rect 2411 2344 2412 2348
rect 2406 2343 2412 2344
rect 2358 2325 2364 2326
rect 2358 2321 2359 2325
rect 2363 2321 2364 2325
rect 2358 2320 2364 2321
rect 2350 2315 2356 2316
rect 2350 2311 2351 2315
rect 2355 2311 2356 2315
rect 2350 2310 2356 2311
rect 2360 2307 2362 2320
rect 2408 2307 2410 2343
rect 2359 2306 2363 2307
rect 2359 2301 2363 2302
rect 2407 2306 2411 2307
rect 2407 2301 2411 2302
rect 2310 2299 2316 2300
rect 2310 2295 2311 2299
rect 2315 2295 2316 2299
rect 2310 2294 2316 2295
rect 2322 2299 2328 2300
rect 2322 2295 2323 2299
rect 2327 2295 2328 2299
rect 2322 2294 2328 2295
rect 2294 2291 2300 2292
rect 2294 2287 2295 2291
rect 2299 2287 2300 2291
rect 2294 2286 2300 2287
rect 2324 2264 2326 2294
rect 2360 2292 2362 2301
rect 2358 2291 2364 2292
rect 2358 2287 2359 2291
rect 2363 2287 2364 2291
rect 2358 2286 2364 2287
rect 2408 2269 2410 2301
rect 2406 2268 2412 2269
rect 2406 2264 2407 2268
rect 2411 2264 2412 2268
rect 2154 2263 2160 2264
rect 2154 2259 2155 2263
rect 2159 2259 2160 2263
rect 2154 2258 2160 2259
rect 2230 2263 2236 2264
rect 2230 2259 2231 2263
rect 2235 2259 2236 2263
rect 2230 2258 2236 2259
rect 2322 2263 2328 2264
rect 2322 2259 2323 2263
rect 2327 2259 2328 2263
rect 2322 2258 2328 2259
rect 2366 2263 2372 2264
rect 2406 2263 2412 2264
rect 2366 2259 2367 2263
rect 2371 2259 2372 2263
rect 2366 2258 2372 2259
rect 2206 2244 2212 2245
rect 2206 2240 2207 2244
rect 2211 2240 2212 2244
rect 2206 2239 2212 2240
rect 2294 2244 2300 2245
rect 2294 2240 2295 2244
rect 2299 2240 2300 2244
rect 2294 2239 2300 2240
rect 2358 2244 2364 2245
rect 2358 2240 2359 2244
rect 2363 2240 2364 2244
rect 2358 2239 2364 2240
rect 2208 2231 2210 2239
rect 2296 2231 2298 2239
rect 2360 2231 2362 2239
rect 2183 2230 2187 2231
rect 2183 2225 2187 2226
rect 2207 2230 2211 2231
rect 2207 2225 2211 2226
rect 2279 2230 2283 2231
rect 2279 2225 2283 2226
rect 2295 2230 2299 2231
rect 2295 2225 2299 2226
rect 2359 2230 2363 2231
rect 2359 2225 2363 2226
rect 2182 2224 2188 2225
rect 2182 2220 2183 2224
rect 2187 2220 2188 2224
rect 2182 2219 2188 2220
rect 2278 2224 2284 2225
rect 2278 2220 2279 2224
rect 2283 2220 2284 2224
rect 2278 2219 2284 2220
rect 2358 2224 2364 2225
rect 2358 2220 2359 2224
rect 2363 2220 2364 2224
rect 2358 2219 2364 2220
rect 1846 2203 1852 2204
rect 1846 2199 1847 2203
rect 1851 2199 1852 2203
rect 1846 2198 1852 2199
rect 1926 2203 1932 2204
rect 1926 2199 1927 2203
rect 1931 2199 1932 2203
rect 1926 2198 1932 2199
rect 2006 2203 2012 2204
rect 2006 2199 2007 2203
rect 2011 2199 2012 2203
rect 2006 2198 2012 2199
rect 2086 2203 2092 2204
rect 2086 2199 2087 2203
rect 2091 2199 2092 2203
rect 2086 2198 2092 2199
rect 2134 2203 2140 2204
rect 2134 2199 2135 2203
rect 2139 2199 2140 2203
rect 2134 2198 2140 2199
rect 2318 2203 2324 2204
rect 2318 2199 2319 2203
rect 2323 2199 2324 2203
rect 2318 2198 2324 2199
rect 1822 2195 1828 2196
rect 1822 2191 1823 2195
rect 1827 2191 1828 2195
rect 1822 2190 1828 2191
rect 1790 2167 1796 2168
rect 1790 2163 1791 2167
rect 1795 2163 1796 2167
rect 1631 2162 1635 2163
rect 1631 2157 1635 2158
rect 1639 2162 1643 2163
rect 1639 2157 1643 2158
rect 1711 2162 1715 2163
rect 1711 2157 1715 2158
rect 1727 2162 1731 2163
rect 1750 2162 1756 2163
rect 1783 2162 1787 2163
rect 1790 2162 1796 2163
rect 1815 2162 1819 2163
rect 1727 2157 1731 2158
rect 1614 2155 1620 2156
rect 1614 2151 1615 2155
rect 1619 2151 1620 2155
rect 1614 2150 1620 2151
rect 1622 2155 1628 2156
rect 1622 2151 1623 2155
rect 1627 2151 1628 2155
rect 1622 2150 1628 2151
rect 1534 2147 1540 2148
rect 1534 2143 1535 2147
rect 1539 2143 1540 2147
rect 1534 2142 1540 2143
rect 1616 2120 1618 2150
rect 1632 2148 1634 2157
rect 1728 2148 1730 2157
rect 1630 2147 1636 2148
rect 1630 2143 1631 2147
rect 1635 2143 1636 2147
rect 1630 2142 1636 2143
rect 1726 2147 1732 2148
rect 1726 2143 1727 2147
rect 1731 2143 1732 2147
rect 1726 2142 1732 2143
rect 1752 2120 1754 2162
rect 1783 2157 1787 2158
rect 1815 2157 1819 2158
rect 1774 2155 1780 2156
rect 1774 2151 1775 2155
rect 1779 2151 1780 2155
rect 1774 2150 1780 2151
rect 1330 2119 1336 2120
rect 1330 2115 1331 2119
rect 1335 2115 1336 2119
rect 1330 2114 1336 2115
rect 1406 2119 1412 2120
rect 1406 2115 1407 2119
rect 1411 2115 1412 2119
rect 1406 2114 1412 2115
rect 1522 2119 1528 2120
rect 1522 2115 1523 2119
rect 1527 2115 1528 2119
rect 1522 2114 1528 2115
rect 1614 2119 1620 2120
rect 1614 2115 1615 2119
rect 1619 2115 1620 2119
rect 1614 2114 1620 2115
rect 1750 2119 1756 2120
rect 1750 2115 1751 2119
rect 1755 2115 1756 2119
rect 1750 2114 1756 2115
rect 1350 2100 1356 2101
rect 1350 2096 1351 2100
rect 1355 2096 1356 2100
rect 1350 2095 1356 2096
rect 1352 2091 1354 2095
rect 1343 2090 1347 2091
rect 1343 2085 1347 2086
rect 1351 2090 1355 2091
rect 1351 2085 1355 2086
rect 1399 2090 1403 2091
rect 1399 2085 1403 2086
rect 1342 2084 1348 2085
rect 1342 2080 1343 2084
rect 1347 2080 1348 2084
rect 1342 2079 1348 2080
rect 1398 2084 1404 2085
rect 1398 2080 1399 2084
rect 1403 2080 1404 2084
rect 1398 2079 1404 2080
rect 1322 2063 1328 2064
rect 1278 2060 1284 2061
rect 1278 2056 1279 2060
rect 1283 2056 1284 2060
rect 1322 2059 1323 2063
rect 1327 2059 1328 2063
rect 1338 2063 1344 2064
rect 1338 2062 1339 2063
rect 1322 2058 1328 2059
rect 1332 2060 1339 2062
rect 1278 2055 1284 2056
rect 1238 2036 1244 2037
rect 1238 2032 1239 2036
rect 1243 2032 1244 2036
rect 826 2031 832 2032
rect 826 2027 827 2031
rect 831 2027 832 2031
rect 826 2026 832 2027
rect 874 2031 880 2032
rect 874 2027 875 2031
rect 879 2027 880 2031
rect 874 2026 880 2027
rect 886 2031 892 2032
rect 886 2027 887 2031
rect 891 2027 892 2031
rect 886 2026 892 2027
rect 1002 2031 1008 2032
rect 1002 2027 1003 2031
rect 1007 2027 1008 2031
rect 1002 2026 1008 2027
rect 1058 2031 1064 2032
rect 1238 2031 1244 2032
rect 1058 2027 1059 2031
rect 1063 2027 1064 2031
rect 1058 2026 1064 2027
rect 878 2023 884 2024
rect 878 2019 879 2023
rect 883 2019 884 2023
rect 878 2018 884 2019
rect 1238 2019 1244 2020
rect 798 2012 804 2013
rect 798 2008 799 2012
rect 803 2008 804 2012
rect 798 2007 804 2008
rect 846 2012 852 2013
rect 846 2008 847 2012
rect 851 2008 852 2012
rect 846 2007 852 2008
rect 800 1999 802 2007
rect 848 1999 850 2007
rect 799 1998 803 1999
rect 799 1993 803 1994
rect 815 1998 819 1999
rect 815 1993 819 1994
rect 847 1998 851 1999
rect 847 1993 851 1994
rect 871 1998 875 1999
rect 871 1993 875 1994
rect 814 1992 820 1993
rect 814 1988 815 1992
rect 819 1988 820 1992
rect 814 1987 820 1988
rect 870 1992 876 1993
rect 870 1988 871 1992
rect 875 1988 876 1992
rect 870 1987 876 1988
rect 394 1971 400 1972
rect 110 1968 116 1969
rect 110 1964 111 1968
rect 115 1964 116 1968
rect 394 1967 395 1971
rect 399 1967 400 1971
rect 394 1966 400 1967
rect 446 1971 452 1972
rect 446 1967 447 1971
rect 451 1967 452 1971
rect 446 1966 452 1967
rect 478 1971 484 1972
rect 478 1967 479 1971
rect 483 1967 484 1971
rect 478 1966 484 1967
rect 602 1971 608 1972
rect 602 1967 603 1971
rect 607 1967 608 1971
rect 602 1966 608 1967
rect 750 1971 756 1972
rect 750 1967 751 1971
rect 755 1967 756 1971
rect 750 1966 756 1967
rect 782 1971 788 1972
rect 782 1967 783 1971
rect 787 1967 788 1971
rect 782 1966 788 1967
rect 110 1963 116 1964
rect 374 1963 380 1964
rect 112 1927 114 1963
rect 374 1959 375 1963
rect 379 1959 380 1963
rect 374 1958 380 1959
rect 366 1945 372 1946
rect 366 1941 367 1945
rect 371 1941 372 1945
rect 366 1940 372 1941
rect 368 1927 370 1940
rect 376 1936 378 1958
rect 396 1936 398 1966
rect 406 1945 412 1946
rect 406 1941 407 1945
rect 411 1941 412 1945
rect 406 1940 412 1941
rect 374 1935 380 1936
rect 374 1931 375 1935
rect 379 1931 380 1935
rect 374 1930 380 1931
rect 394 1935 400 1936
rect 394 1931 395 1935
rect 399 1931 400 1935
rect 394 1930 400 1931
rect 408 1927 410 1940
rect 448 1936 450 1966
rect 454 1945 460 1946
rect 454 1941 455 1945
rect 459 1941 460 1945
rect 454 1940 460 1941
rect 446 1935 452 1936
rect 446 1931 447 1935
rect 451 1931 452 1935
rect 446 1930 452 1931
rect 456 1927 458 1940
rect 111 1926 115 1927
rect 111 1921 115 1922
rect 175 1926 179 1927
rect 175 1921 179 1922
rect 215 1926 219 1927
rect 215 1921 219 1922
rect 263 1926 267 1927
rect 263 1921 267 1922
rect 319 1926 323 1927
rect 319 1921 323 1922
rect 367 1926 371 1927
rect 367 1921 371 1922
rect 391 1926 395 1927
rect 391 1921 395 1922
rect 407 1926 411 1927
rect 407 1921 411 1922
rect 455 1926 459 1927
rect 455 1921 459 1922
rect 471 1926 475 1927
rect 471 1921 475 1922
rect 112 1889 114 1921
rect 176 1912 178 1921
rect 190 1919 196 1920
rect 190 1915 191 1919
rect 195 1915 196 1919
rect 190 1914 196 1915
rect 198 1919 204 1920
rect 198 1915 199 1919
rect 203 1915 204 1919
rect 198 1914 204 1915
rect 174 1911 180 1912
rect 174 1907 175 1911
rect 179 1907 180 1911
rect 174 1906 180 1907
rect 192 1892 194 1914
rect 190 1891 196 1892
rect 110 1888 116 1889
rect 110 1884 111 1888
rect 115 1884 116 1888
rect 190 1887 191 1891
rect 195 1887 196 1891
rect 190 1886 196 1887
rect 200 1884 202 1914
rect 216 1912 218 1921
rect 264 1912 266 1921
rect 320 1912 322 1921
rect 378 1919 384 1920
rect 378 1915 379 1919
rect 383 1915 384 1919
rect 378 1914 384 1915
rect 214 1911 220 1912
rect 214 1907 215 1911
rect 219 1907 220 1911
rect 214 1906 220 1907
rect 262 1911 268 1912
rect 262 1907 263 1911
rect 267 1907 268 1911
rect 262 1906 268 1907
rect 318 1911 324 1912
rect 318 1907 319 1911
rect 323 1907 324 1911
rect 318 1906 324 1907
rect 380 1884 382 1914
rect 392 1912 394 1921
rect 472 1912 474 1921
rect 480 1920 482 1966
rect 510 1945 516 1946
rect 510 1941 511 1945
rect 515 1941 516 1945
rect 510 1940 516 1941
rect 566 1945 572 1946
rect 566 1941 567 1945
rect 571 1941 572 1945
rect 566 1940 572 1941
rect 512 1927 514 1940
rect 568 1927 570 1940
rect 604 1936 606 1966
rect 702 1963 708 1964
rect 702 1959 703 1963
rect 707 1959 708 1963
rect 702 1958 708 1959
rect 630 1945 636 1946
rect 630 1941 631 1945
rect 635 1941 636 1945
rect 630 1940 636 1941
rect 694 1945 700 1946
rect 694 1941 695 1945
rect 699 1941 700 1945
rect 694 1940 700 1941
rect 602 1935 608 1936
rect 602 1931 603 1935
rect 607 1931 608 1935
rect 602 1930 608 1931
rect 632 1927 634 1940
rect 696 1927 698 1940
rect 704 1936 706 1958
rect 752 1936 754 1966
rect 758 1945 764 1946
rect 758 1941 759 1945
rect 763 1941 764 1945
rect 758 1940 764 1941
rect 814 1945 820 1946
rect 814 1941 815 1945
rect 819 1941 820 1945
rect 814 1940 820 1941
rect 870 1945 876 1946
rect 870 1941 871 1945
rect 875 1941 876 1945
rect 870 1940 876 1941
rect 702 1935 708 1936
rect 702 1931 703 1935
rect 707 1931 708 1935
rect 702 1930 708 1931
rect 750 1935 756 1936
rect 750 1931 751 1935
rect 755 1931 756 1935
rect 750 1930 756 1931
rect 760 1927 762 1940
rect 816 1927 818 1940
rect 822 1935 828 1936
rect 822 1931 823 1935
rect 827 1931 828 1935
rect 822 1930 828 1931
rect 511 1926 515 1927
rect 511 1921 515 1922
rect 551 1926 555 1927
rect 551 1921 555 1922
rect 567 1926 571 1927
rect 567 1921 571 1922
rect 631 1926 635 1927
rect 631 1921 635 1922
rect 639 1926 643 1927
rect 639 1921 643 1922
rect 695 1926 699 1927
rect 695 1921 699 1922
rect 719 1926 723 1927
rect 719 1921 723 1922
rect 759 1926 763 1927
rect 759 1921 763 1922
rect 799 1926 803 1927
rect 799 1921 803 1922
rect 815 1926 819 1927
rect 815 1921 819 1922
rect 478 1919 484 1920
rect 478 1915 479 1919
rect 483 1915 484 1919
rect 478 1914 484 1915
rect 498 1919 504 1920
rect 498 1915 499 1919
rect 503 1915 504 1919
rect 498 1914 504 1915
rect 390 1911 396 1912
rect 390 1907 391 1911
rect 395 1907 396 1911
rect 390 1906 396 1907
rect 470 1911 476 1912
rect 470 1907 471 1911
rect 475 1907 476 1911
rect 470 1906 476 1907
rect 500 1884 502 1914
rect 552 1912 554 1921
rect 640 1912 642 1921
rect 654 1919 660 1920
rect 654 1915 655 1919
rect 659 1915 660 1919
rect 654 1914 660 1915
rect 550 1911 556 1912
rect 550 1907 551 1911
rect 555 1907 556 1911
rect 550 1906 556 1907
rect 638 1911 644 1912
rect 638 1907 639 1911
rect 643 1907 644 1911
rect 638 1906 644 1907
rect 110 1883 116 1884
rect 198 1883 204 1884
rect 198 1879 199 1883
rect 203 1879 204 1883
rect 198 1878 204 1879
rect 334 1883 340 1884
rect 334 1879 335 1883
rect 339 1879 340 1883
rect 334 1878 340 1879
rect 378 1883 384 1884
rect 378 1879 379 1883
rect 383 1879 384 1883
rect 378 1878 384 1879
rect 498 1883 504 1884
rect 498 1879 499 1883
rect 503 1879 504 1883
rect 498 1878 504 1879
rect 110 1871 116 1872
rect 110 1867 111 1871
rect 115 1867 116 1871
rect 110 1866 116 1867
rect 112 1851 114 1866
rect 174 1864 180 1865
rect 174 1860 175 1864
rect 179 1860 180 1864
rect 174 1859 180 1860
rect 214 1864 220 1865
rect 214 1860 215 1864
rect 219 1860 220 1864
rect 214 1859 220 1860
rect 262 1864 268 1865
rect 262 1860 263 1864
rect 267 1860 268 1864
rect 262 1859 268 1860
rect 318 1864 324 1865
rect 318 1860 319 1864
rect 323 1860 324 1864
rect 318 1859 324 1860
rect 176 1851 178 1859
rect 216 1851 218 1859
rect 264 1851 266 1859
rect 320 1851 322 1859
rect 111 1850 115 1851
rect 111 1845 115 1846
rect 135 1850 139 1851
rect 135 1845 139 1846
rect 175 1850 179 1851
rect 175 1845 179 1846
rect 215 1850 219 1851
rect 215 1845 219 1846
rect 263 1850 267 1851
rect 263 1845 267 1846
rect 271 1850 275 1851
rect 271 1845 275 1846
rect 319 1850 323 1851
rect 319 1845 323 1846
rect 112 1838 114 1845
rect 134 1844 140 1845
rect 134 1840 135 1844
rect 139 1840 140 1844
rect 134 1839 140 1840
rect 174 1844 180 1845
rect 174 1840 175 1844
rect 179 1840 180 1844
rect 174 1839 180 1840
rect 214 1844 220 1845
rect 214 1840 215 1844
rect 219 1840 220 1844
rect 214 1839 220 1840
rect 270 1844 276 1845
rect 270 1840 271 1844
rect 275 1840 276 1844
rect 270 1839 276 1840
rect 110 1837 116 1838
rect 110 1833 111 1837
rect 115 1833 116 1837
rect 110 1832 116 1833
rect 142 1823 148 1824
rect 110 1820 116 1821
rect 110 1816 111 1820
rect 115 1816 116 1820
rect 142 1819 143 1823
rect 147 1819 148 1823
rect 142 1818 148 1819
rect 110 1815 116 1816
rect 112 1783 114 1815
rect 134 1797 140 1798
rect 134 1793 135 1797
rect 139 1793 140 1797
rect 134 1792 140 1793
rect 136 1783 138 1792
rect 111 1782 115 1783
rect 111 1777 115 1778
rect 135 1782 139 1783
rect 135 1777 139 1778
rect 112 1745 114 1777
rect 136 1768 138 1777
rect 144 1776 146 1818
rect 150 1815 156 1816
rect 150 1811 151 1815
rect 155 1811 156 1815
rect 150 1810 156 1811
rect 182 1815 188 1816
rect 182 1811 183 1815
rect 187 1811 188 1815
rect 182 1810 188 1811
rect 294 1815 300 1816
rect 294 1811 295 1815
rect 299 1811 300 1815
rect 294 1810 300 1811
rect 152 1788 154 1810
rect 174 1797 180 1798
rect 174 1793 175 1797
rect 179 1793 180 1797
rect 174 1792 180 1793
rect 150 1787 156 1788
rect 150 1783 151 1787
rect 155 1783 156 1787
rect 176 1783 178 1792
rect 184 1788 186 1810
rect 214 1797 220 1798
rect 214 1793 215 1797
rect 219 1793 220 1797
rect 214 1792 220 1793
rect 270 1797 276 1798
rect 270 1793 271 1797
rect 275 1793 276 1797
rect 270 1792 276 1793
rect 182 1787 188 1788
rect 182 1783 183 1787
rect 187 1783 188 1787
rect 216 1783 218 1792
rect 272 1783 274 1792
rect 296 1788 298 1810
rect 336 1788 338 1878
rect 390 1864 396 1865
rect 390 1860 391 1864
rect 395 1860 396 1864
rect 390 1859 396 1860
rect 470 1864 476 1865
rect 470 1860 471 1864
rect 475 1860 476 1864
rect 470 1859 476 1860
rect 550 1864 556 1865
rect 550 1860 551 1864
rect 555 1860 556 1864
rect 550 1859 556 1860
rect 638 1864 644 1865
rect 638 1860 639 1864
rect 643 1860 644 1864
rect 638 1859 644 1860
rect 392 1851 394 1859
rect 472 1851 474 1859
rect 552 1851 554 1859
rect 640 1851 642 1859
rect 351 1850 355 1851
rect 351 1845 355 1846
rect 391 1850 395 1851
rect 391 1845 395 1846
rect 439 1850 443 1851
rect 439 1845 443 1846
rect 471 1850 475 1851
rect 471 1845 475 1846
rect 535 1850 539 1851
rect 535 1845 539 1846
rect 551 1850 555 1851
rect 551 1845 555 1846
rect 631 1850 635 1851
rect 631 1845 635 1846
rect 639 1850 643 1851
rect 639 1845 643 1846
rect 350 1844 356 1845
rect 350 1840 351 1844
rect 355 1840 356 1844
rect 350 1839 356 1840
rect 438 1844 444 1845
rect 438 1840 439 1844
rect 443 1840 444 1844
rect 438 1839 444 1840
rect 534 1844 540 1845
rect 534 1840 535 1844
rect 539 1840 540 1844
rect 534 1839 540 1840
rect 630 1844 636 1845
rect 630 1840 631 1844
rect 635 1840 636 1844
rect 630 1839 636 1840
rect 656 1824 658 1914
rect 720 1912 722 1921
rect 746 1919 752 1920
rect 746 1915 747 1919
rect 751 1915 752 1919
rect 746 1914 752 1915
rect 718 1911 724 1912
rect 718 1907 719 1911
rect 723 1907 724 1911
rect 718 1906 724 1907
rect 748 1884 750 1914
rect 800 1912 802 1921
rect 798 1911 804 1912
rect 798 1907 799 1911
rect 803 1907 804 1911
rect 798 1906 804 1907
rect 824 1884 826 1930
rect 872 1927 874 1940
rect 880 1936 882 2018
rect 1238 2015 1239 2019
rect 1243 2015 1244 2019
rect 1280 2015 1282 2055
rect 1302 2037 1308 2038
rect 1302 2033 1303 2037
rect 1307 2033 1308 2037
rect 1302 2032 1308 2033
rect 1304 2015 1306 2032
rect 1332 2028 1334 2060
rect 1338 2059 1339 2060
rect 1343 2059 1344 2063
rect 1338 2058 1344 2059
rect 1342 2037 1348 2038
rect 1342 2033 1343 2037
rect 1347 2033 1348 2037
rect 1342 2032 1348 2033
rect 1398 2037 1404 2038
rect 1398 2033 1399 2037
rect 1403 2033 1404 2037
rect 1398 2032 1404 2033
rect 1330 2027 1336 2028
rect 1330 2023 1331 2027
rect 1335 2023 1336 2027
rect 1330 2022 1336 2023
rect 1344 2015 1346 2032
rect 1374 2027 1380 2028
rect 1374 2023 1375 2027
rect 1379 2023 1380 2027
rect 1374 2022 1380 2023
rect 1238 2014 1244 2015
rect 1279 2014 1283 2015
rect 902 2012 908 2013
rect 902 2008 903 2012
rect 907 2008 908 2012
rect 902 2007 908 2008
rect 958 2012 964 2013
rect 958 2008 959 2012
rect 963 2008 964 2012
rect 958 2007 964 2008
rect 1014 2012 1020 2013
rect 1014 2008 1015 2012
rect 1019 2008 1020 2012
rect 1014 2007 1020 2008
rect 1070 2012 1076 2013
rect 1070 2008 1071 2012
rect 1075 2008 1076 2012
rect 1070 2007 1076 2008
rect 904 1999 906 2007
rect 960 1999 962 2007
rect 1016 1999 1018 2007
rect 1072 1999 1074 2007
rect 1240 1999 1242 2014
rect 1279 2009 1283 2010
rect 1303 2014 1307 2015
rect 1303 2009 1307 2010
rect 1343 2014 1347 2015
rect 1343 2009 1347 2010
rect 1351 2014 1355 2015
rect 1351 2009 1355 2010
rect 903 1998 907 1999
rect 903 1993 907 1994
rect 935 1998 939 1999
rect 935 1993 939 1994
rect 959 1998 963 1999
rect 959 1993 963 1994
rect 999 1998 1003 1999
rect 999 1993 1003 1994
rect 1015 1998 1019 1999
rect 1015 1993 1019 1994
rect 1063 1998 1067 1999
rect 1063 1993 1067 1994
rect 1071 1998 1075 1999
rect 1071 1993 1075 1994
rect 1239 1998 1243 1999
rect 1239 1993 1243 1994
rect 934 1992 940 1993
rect 934 1988 935 1992
rect 939 1988 940 1992
rect 934 1987 940 1988
rect 998 1992 1004 1993
rect 998 1988 999 1992
rect 1003 1988 1004 1992
rect 998 1987 1004 1988
rect 1062 1992 1068 1993
rect 1062 1988 1063 1992
rect 1067 1988 1068 1992
rect 1062 1987 1068 1988
rect 1240 1986 1242 1993
rect 1238 1985 1244 1986
rect 1238 1981 1239 1985
rect 1243 1981 1244 1985
rect 1238 1980 1244 1981
rect 1280 1977 1282 2009
rect 1304 2000 1306 2009
rect 1322 2007 1328 2008
rect 1322 2003 1323 2007
rect 1327 2003 1328 2007
rect 1322 2002 1328 2003
rect 1330 2007 1336 2008
rect 1330 2003 1331 2007
rect 1335 2003 1336 2007
rect 1330 2002 1336 2003
rect 1302 1999 1308 2000
rect 1302 1995 1303 1999
rect 1307 1995 1308 1999
rect 1302 1994 1308 1995
rect 1278 1976 1284 1977
rect 1278 1972 1279 1976
rect 1283 1972 1284 1976
rect 926 1971 932 1972
rect 926 1967 927 1971
rect 931 1967 932 1971
rect 926 1966 932 1967
rect 990 1971 996 1972
rect 990 1967 991 1971
rect 995 1967 996 1971
rect 990 1966 996 1967
rect 1054 1971 1060 1972
rect 1054 1967 1055 1971
rect 1059 1967 1060 1971
rect 1054 1966 1060 1967
rect 1070 1971 1076 1972
rect 1278 1971 1284 1972
rect 1070 1967 1071 1971
rect 1075 1967 1076 1971
rect 1070 1966 1076 1967
rect 1238 1968 1244 1969
rect 928 1936 930 1966
rect 934 1945 940 1946
rect 934 1941 935 1945
rect 939 1941 940 1945
rect 934 1940 940 1941
rect 878 1935 884 1936
rect 878 1931 879 1935
rect 883 1931 884 1935
rect 878 1930 884 1931
rect 926 1935 932 1936
rect 926 1931 927 1935
rect 931 1931 932 1935
rect 926 1930 932 1931
rect 936 1927 938 1940
rect 992 1936 994 1966
rect 998 1945 1004 1946
rect 998 1941 999 1945
rect 1003 1941 1004 1945
rect 998 1940 1004 1941
rect 990 1935 996 1936
rect 990 1931 991 1935
rect 995 1931 996 1935
rect 990 1930 996 1931
rect 1000 1927 1002 1940
rect 1056 1936 1058 1966
rect 1062 1945 1068 1946
rect 1062 1941 1063 1945
rect 1067 1941 1068 1945
rect 1062 1940 1068 1941
rect 1054 1935 1060 1936
rect 1054 1931 1055 1935
rect 1059 1931 1060 1935
rect 1054 1930 1060 1931
rect 1064 1927 1066 1940
rect 1072 1928 1074 1966
rect 1238 1964 1239 1968
rect 1243 1964 1244 1968
rect 1238 1963 1244 1964
rect 1070 1927 1076 1928
rect 1240 1927 1242 1963
rect 1278 1959 1284 1960
rect 1278 1955 1279 1959
rect 1283 1955 1284 1959
rect 1278 1954 1284 1955
rect 1280 1947 1282 1954
rect 1302 1952 1308 1953
rect 1302 1948 1303 1952
rect 1307 1948 1308 1952
rect 1302 1947 1308 1948
rect 1279 1946 1283 1947
rect 1279 1941 1283 1942
rect 1303 1946 1307 1947
rect 1303 1941 1307 1942
rect 1280 1934 1282 1941
rect 1302 1940 1308 1941
rect 1302 1936 1303 1940
rect 1307 1936 1308 1940
rect 1302 1935 1308 1936
rect 1278 1933 1284 1934
rect 1278 1929 1279 1933
rect 1283 1929 1284 1933
rect 1278 1928 1284 1929
rect 871 1926 875 1927
rect 871 1921 875 1922
rect 879 1926 883 1927
rect 879 1921 883 1922
rect 935 1926 939 1927
rect 935 1921 939 1922
rect 959 1926 963 1927
rect 959 1921 963 1922
rect 999 1926 1003 1927
rect 999 1921 1003 1922
rect 1039 1926 1043 1927
rect 1039 1921 1043 1922
rect 1063 1926 1067 1927
rect 1070 1923 1071 1927
rect 1075 1923 1076 1927
rect 1070 1922 1076 1923
rect 1119 1926 1123 1927
rect 1063 1921 1067 1922
rect 1119 1921 1123 1922
rect 1239 1926 1243 1927
rect 1239 1921 1243 1922
rect 880 1912 882 1921
rect 902 1919 908 1920
rect 902 1915 903 1919
rect 907 1915 908 1919
rect 902 1914 908 1915
rect 878 1911 884 1912
rect 878 1907 879 1911
rect 883 1907 884 1911
rect 878 1906 884 1907
rect 904 1884 906 1914
rect 960 1912 962 1921
rect 986 1919 992 1920
rect 986 1915 987 1919
rect 991 1915 992 1919
rect 986 1914 992 1915
rect 958 1911 964 1912
rect 958 1907 959 1911
rect 963 1907 964 1911
rect 958 1906 964 1907
rect 988 1884 990 1914
rect 1040 1912 1042 1921
rect 1070 1919 1076 1920
rect 1070 1915 1071 1919
rect 1075 1915 1076 1919
rect 1070 1914 1076 1915
rect 1038 1911 1044 1912
rect 1038 1907 1039 1911
rect 1043 1907 1044 1911
rect 1038 1906 1044 1907
rect 1072 1884 1074 1914
rect 1120 1912 1122 1921
rect 1118 1911 1124 1912
rect 1118 1907 1119 1911
rect 1123 1907 1124 1911
rect 1118 1906 1124 1907
rect 1240 1889 1242 1921
rect 1324 1920 1326 2002
rect 1332 1972 1334 2002
rect 1352 2000 1354 2009
rect 1350 1999 1356 2000
rect 1350 1995 1351 1999
rect 1355 1995 1356 1999
rect 1350 1994 1356 1995
rect 1376 1972 1378 2022
rect 1400 2015 1402 2032
rect 1408 2028 1410 2114
rect 1438 2100 1444 2101
rect 1438 2096 1439 2100
rect 1443 2096 1444 2100
rect 1438 2095 1444 2096
rect 1534 2100 1540 2101
rect 1534 2096 1535 2100
rect 1539 2096 1540 2100
rect 1534 2095 1540 2096
rect 1630 2100 1636 2101
rect 1630 2096 1631 2100
rect 1635 2096 1636 2100
rect 1630 2095 1636 2096
rect 1726 2100 1732 2101
rect 1726 2096 1727 2100
rect 1731 2096 1732 2100
rect 1726 2095 1732 2096
rect 1440 2091 1442 2095
rect 1536 2091 1538 2095
rect 1632 2091 1634 2095
rect 1728 2091 1730 2095
rect 1439 2090 1443 2091
rect 1439 2085 1443 2086
rect 1479 2090 1483 2091
rect 1479 2085 1483 2086
rect 1535 2090 1539 2091
rect 1535 2085 1539 2086
rect 1567 2090 1571 2091
rect 1567 2085 1571 2086
rect 1631 2090 1635 2091
rect 1631 2085 1635 2086
rect 1663 2090 1667 2091
rect 1663 2085 1667 2086
rect 1727 2090 1731 2091
rect 1727 2085 1731 2086
rect 1759 2090 1763 2091
rect 1759 2085 1763 2086
rect 1478 2084 1484 2085
rect 1478 2080 1479 2084
rect 1483 2080 1484 2084
rect 1478 2079 1484 2080
rect 1566 2084 1572 2085
rect 1566 2080 1567 2084
rect 1571 2080 1572 2084
rect 1566 2079 1572 2080
rect 1662 2084 1668 2085
rect 1662 2080 1663 2084
rect 1667 2080 1668 2084
rect 1662 2079 1668 2080
rect 1758 2084 1764 2085
rect 1758 2080 1759 2084
rect 1763 2080 1764 2084
rect 1758 2079 1764 2080
rect 1776 2064 1778 2150
rect 1816 2148 1818 2157
rect 1824 2156 1826 2190
rect 1848 2168 1850 2198
rect 1854 2177 1860 2178
rect 1854 2173 1855 2177
rect 1859 2173 1860 2177
rect 1854 2172 1860 2173
rect 1846 2167 1852 2168
rect 1846 2163 1847 2167
rect 1851 2163 1852 2167
rect 1856 2163 1858 2172
rect 1928 2168 1930 2198
rect 1934 2177 1940 2178
rect 1934 2173 1935 2177
rect 1939 2173 1940 2177
rect 1934 2172 1940 2173
rect 1926 2167 1932 2168
rect 1926 2163 1927 2167
rect 1931 2163 1932 2167
rect 1936 2163 1938 2172
rect 2008 2168 2010 2198
rect 2014 2177 2020 2178
rect 2014 2173 2015 2177
rect 2019 2173 2020 2177
rect 2014 2172 2020 2173
rect 2006 2167 2012 2168
rect 2006 2163 2007 2167
rect 2011 2163 2012 2167
rect 2016 2163 2018 2172
rect 2088 2168 2090 2198
rect 2094 2177 2100 2178
rect 2094 2173 2095 2177
rect 2099 2173 2100 2177
rect 2094 2172 2100 2173
rect 2182 2177 2188 2178
rect 2182 2173 2183 2177
rect 2187 2173 2188 2177
rect 2182 2172 2188 2173
rect 2278 2177 2284 2178
rect 2278 2173 2279 2177
rect 2283 2173 2284 2177
rect 2278 2172 2284 2173
rect 2086 2167 2092 2168
rect 2086 2163 2087 2167
rect 2091 2163 2092 2167
rect 2096 2163 2098 2172
rect 2184 2163 2186 2172
rect 2266 2167 2272 2168
rect 2266 2163 2267 2167
rect 2271 2163 2272 2167
rect 2280 2163 2282 2172
rect 1846 2162 1852 2163
rect 1855 2162 1859 2163
rect 1855 2157 1859 2158
rect 1895 2162 1899 2163
rect 1926 2162 1932 2163
rect 1935 2162 1939 2163
rect 1895 2157 1899 2158
rect 1935 2157 1939 2158
rect 1975 2162 1979 2163
rect 2006 2162 2012 2163
rect 2015 2162 2019 2163
rect 1975 2157 1979 2158
rect 2015 2157 2019 2158
rect 2047 2162 2051 2163
rect 2086 2162 2092 2163
rect 2095 2162 2099 2163
rect 2047 2157 2051 2158
rect 2095 2157 2099 2158
rect 2111 2162 2115 2163
rect 2111 2157 2115 2158
rect 2175 2162 2179 2163
rect 2175 2157 2179 2158
rect 2183 2162 2187 2163
rect 2183 2157 2187 2158
rect 2239 2162 2243 2163
rect 2266 2162 2272 2163
rect 2279 2162 2283 2163
rect 2239 2157 2243 2158
rect 1822 2155 1828 2156
rect 1822 2151 1823 2155
rect 1827 2151 1828 2155
rect 1822 2150 1828 2151
rect 1842 2155 1848 2156
rect 1842 2151 1843 2155
rect 1847 2151 1848 2155
rect 1842 2150 1848 2151
rect 1814 2147 1820 2148
rect 1814 2143 1815 2147
rect 1819 2143 1820 2147
rect 1814 2142 1820 2143
rect 1844 2120 1846 2150
rect 1896 2148 1898 2157
rect 1976 2148 1978 2157
rect 1998 2155 2004 2156
rect 1998 2151 1999 2155
rect 2003 2151 2004 2155
rect 1998 2150 2004 2151
rect 1894 2147 1900 2148
rect 1894 2143 1895 2147
rect 1899 2143 1900 2147
rect 1894 2142 1900 2143
rect 1974 2147 1980 2148
rect 1974 2143 1975 2147
rect 1979 2143 1980 2147
rect 1974 2142 1980 2143
rect 2000 2120 2002 2150
rect 2048 2148 2050 2157
rect 2054 2155 2060 2156
rect 2054 2151 2055 2155
rect 2059 2151 2060 2155
rect 2054 2150 2060 2151
rect 2046 2147 2052 2148
rect 2046 2143 2047 2147
rect 2051 2143 2052 2147
rect 2046 2142 2052 2143
rect 1842 2119 1848 2120
rect 1842 2115 1843 2119
rect 1847 2115 1848 2119
rect 1842 2114 1848 2115
rect 1998 2119 2004 2120
rect 1998 2115 1999 2119
rect 2003 2115 2004 2119
rect 1998 2114 2004 2115
rect 1942 2111 1948 2112
rect 1942 2107 1943 2111
rect 1947 2107 1948 2111
rect 1942 2106 1948 2107
rect 1814 2100 1820 2101
rect 1814 2096 1815 2100
rect 1819 2096 1820 2100
rect 1814 2095 1820 2096
rect 1894 2100 1900 2101
rect 1894 2096 1895 2100
rect 1899 2096 1900 2100
rect 1894 2095 1900 2096
rect 1816 2091 1818 2095
rect 1896 2091 1898 2095
rect 1815 2090 1819 2091
rect 1815 2085 1819 2086
rect 1847 2090 1851 2091
rect 1847 2085 1851 2086
rect 1895 2090 1899 2091
rect 1895 2085 1899 2086
rect 1935 2090 1939 2091
rect 1935 2085 1939 2086
rect 1846 2084 1852 2085
rect 1846 2080 1847 2084
rect 1851 2080 1852 2084
rect 1846 2079 1852 2080
rect 1934 2084 1940 2085
rect 1934 2080 1935 2084
rect 1939 2080 1940 2084
rect 1934 2079 1940 2080
rect 1470 2063 1476 2064
rect 1470 2059 1471 2063
rect 1475 2059 1476 2063
rect 1470 2058 1476 2059
rect 1546 2063 1552 2064
rect 1546 2059 1547 2063
rect 1551 2059 1552 2063
rect 1546 2058 1552 2059
rect 1654 2063 1660 2064
rect 1654 2059 1655 2063
rect 1659 2059 1660 2063
rect 1654 2058 1660 2059
rect 1670 2063 1676 2064
rect 1670 2059 1671 2063
rect 1675 2059 1676 2063
rect 1670 2058 1676 2059
rect 1774 2063 1780 2064
rect 1774 2059 1775 2063
rect 1779 2059 1780 2063
rect 1774 2058 1780 2059
rect 1472 2028 1474 2058
rect 1478 2037 1484 2038
rect 1478 2033 1479 2037
rect 1483 2033 1484 2037
rect 1478 2032 1484 2033
rect 1406 2027 1412 2028
rect 1406 2023 1407 2027
rect 1411 2023 1412 2027
rect 1406 2022 1412 2023
rect 1470 2027 1476 2028
rect 1470 2023 1471 2027
rect 1475 2023 1476 2027
rect 1470 2022 1476 2023
rect 1480 2015 1482 2032
rect 1548 2028 1550 2058
rect 1566 2037 1572 2038
rect 1566 2033 1567 2037
rect 1571 2033 1572 2037
rect 1566 2032 1572 2033
rect 1546 2027 1552 2028
rect 1546 2023 1547 2027
rect 1551 2023 1552 2027
rect 1546 2022 1552 2023
rect 1568 2015 1570 2032
rect 1656 2028 1658 2058
rect 1662 2037 1668 2038
rect 1662 2033 1663 2037
rect 1667 2033 1668 2037
rect 1662 2032 1668 2033
rect 1654 2027 1660 2028
rect 1654 2023 1655 2027
rect 1659 2023 1660 2027
rect 1654 2022 1660 2023
rect 1664 2015 1666 2032
rect 1672 2016 1674 2058
rect 1758 2037 1764 2038
rect 1758 2033 1759 2037
rect 1763 2033 1764 2037
rect 1758 2032 1764 2033
rect 1846 2037 1852 2038
rect 1846 2033 1847 2037
rect 1851 2033 1852 2037
rect 1846 2032 1852 2033
rect 1934 2037 1940 2038
rect 1934 2033 1935 2037
rect 1939 2033 1940 2037
rect 1934 2032 1940 2033
rect 1670 2015 1676 2016
rect 1760 2015 1762 2032
rect 1848 2015 1850 2032
rect 1862 2027 1868 2028
rect 1862 2023 1863 2027
rect 1867 2023 1868 2027
rect 1862 2022 1868 2023
rect 1399 2014 1403 2015
rect 1399 2009 1403 2010
rect 1423 2014 1427 2015
rect 1423 2009 1427 2010
rect 1479 2014 1483 2015
rect 1479 2009 1483 2010
rect 1495 2014 1499 2015
rect 1495 2009 1499 2010
rect 1567 2014 1571 2015
rect 1567 2009 1571 2010
rect 1575 2014 1579 2015
rect 1575 2009 1579 2010
rect 1663 2014 1667 2015
rect 1670 2011 1671 2015
rect 1675 2011 1676 2015
rect 1670 2010 1676 2011
rect 1751 2014 1755 2015
rect 1663 2009 1667 2010
rect 1751 2009 1755 2010
rect 1759 2014 1763 2015
rect 1759 2009 1763 2010
rect 1839 2014 1843 2015
rect 1839 2009 1843 2010
rect 1847 2014 1851 2015
rect 1847 2009 1851 2010
rect 1424 2000 1426 2009
rect 1442 2007 1448 2008
rect 1442 2003 1443 2007
rect 1447 2003 1448 2007
rect 1442 2002 1448 2003
rect 1450 2007 1456 2008
rect 1450 2003 1451 2007
rect 1455 2003 1456 2007
rect 1450 2002 1456 2003
rect 1422 1999 1428 2000
rect 1422 1995 1423 1999
rect 1427 1995 1428 1999
rect 1422 1994 1428 1995
rect 1444 1980 1446 2002
rect 1442 1979 1448 1980
rect 1442 1975 1443 1979
rect 1447 1975 1448 1979
rect 1442 1974 1448 1975
rect 1452 1972 1454 2002
rect 1496 2000 1498 2009
rect 1576 2000 1578 2009
rect 1664 2000 1666 2009
rect 1690 2007 1696 2008
rect 1690 2003 1691 2007
rect 1695 2003 1696 2007
rect 1690 2002 1696 2003
rect 1494 1999 1500 2000
rect 1494 1995 1495 1999
rect 1499 1995 1500 1999
rect 1494 1994 1500 1995
rect 1574 1999 1580 2000
rect 1574 1995 1575 1999
rect 1579 1995 1580 1999
rect 1574 1994 1580 1995
rect 1662 1999 1668 2000
rect 1662 1995 1663 1999
rect 1667 1995 1668 1999
rect 1662 1994 1668 1995
rect 1692 1972 1694 2002
rect 1752 2000 1754 2009
rect 1778 2007 1784 2008
rect 1778 2003 1779 2007
rect 1783 2003 1784 2007
rect 1778 2002 1784 2003
rect 1734 1999 1740 2000
rect 1734 1995 1735 1999
rect 1739 1995 1740 1999
rect 1734 1994 1740 1995
rect 1750 1999 1756 2000
rect 1750 1995 1751 1999
rect 1755 1995 1756 1999
rect 1750 1994 1756 1995
rect 1330 1971 1336 1972
rect 1330 1967 1331 1971
rect 1335 1967 1336 1971
rect 1330 1966 1336 1967
rect 1374 1971 1380 1972
rect 1374 1967 1375 1971
rect 1379 1967 1380 1971
rect 1374 1966 1380 1967
rect 1450 1971 1456 1972
rect 1450 1967 1451 1971
rect 1455 1967 1456 1971
rect 1450 1966 1456 1967
rect 1522 1971 1528 1972
rect 1522 1967 1523 1971
rect 1527 1967 1528 1971
rect 1522 1966 1528 1967
rect 1690 1971 1696 1972
rect 1690 1967 1691 1971
rect 1695 1967 1696 1971
rect 1690 1966 1696 1967
rect 1350 1952 1356 1953
rect 1350 1948 1351 1952
rect 1355 1948 1356 1952
rect 1350 1947 1356 1948
rect 1422 1952 1428 1953
rect 1422 1948 1423 1952
rect 1427 1948 1428 1952
rect 1422 1947 1428 1948
rect 1494 1952 1500 1953
rect 1494 1948 1495 1952
rect 1499 1948 1500 1952
rect 1494 1947 1500 1948
rect 1351 1946 1355 1947
rect 1351 1941 1355 1942
rect 1359 1946 1363 1947
rect 1359 1941 1363 1942
rect 1423 1946 1427 1947
rect 1423 1941 1427 1942
rect 1447 1946 1451 1947
rect 1447 1941 1451 1942
rect 1495 1946 1499 1947
rect 1495 1941 1499 1942
rect 1358 1940 1364 1941
rect 1358 1936 1359 1940
rect 1363 1936 1364 1940
rect 1358 1935 1364 1936
rect 1446 1940 1452 1941
rect 1446 1936 1447 1940
rect 1451 1936 1452 1940
rect 1446 1935 1452 1936
rect 1322 1919 1328 1920
rect 1278 1916 1284 1917
rect 1278 1912 1279 1916
rect 1283 1912 1284 1916
rect 1322 1915 1323 1919
rect 1327 1915 1328 1919
rect 1322 1914 1328 1915
rect 1278 1911 1284 1912
rect 746 1883 752 1884
rect 746 1879 747 1883
rect 751 1879 752 1883
rect 746 1878 752 1879
rect 822 1883 828 1884
rect 822 1879 823 1883
rect 827 1879 828 1883
rect 822 1878 828 1879
rect 902 1883 908 1884
rect 902 1879 903 1883
rect 907 1879 908 1883
rect 902 1878 908 1879
rect 986 1883 992 1884
rect 986 1879 987 1883
rect 991 1879 992 1883
rect 986 1878 992 1879
rect 1066 1883 1074 1884
rect 1238 1888 1244 1889
rect 1238 1884 1239 1888
rect 1243 1884 1244 1888
rect 1238 1883 1244 1884
rect 1066 1879 1067 1883
rect 1071 1880 1074 1883
rect 1071 1879 1072 1880
rect 1280 1879 1282 1911
rect 1302 1893 1308 1894
rect 1302 1889 1303 1893
rect 1307 1889 1308 1893
rect 1302 1888 1308 1889
rect 1358 1893 1364 1894
rect 1358 1889 1359 1893
rect 1363 1889 1364 1893
rect 1358 1888 1364 1889
rect 1446 1893 1452 1894
rect 1446 1889 1447 1893
rect 1451 1889 1452 1893
rect 1446 1888 1452 1889
rect 1304 1879 1306 1888
rect 1360 1879 1362 1888
rect 1438 1883 1444 1884
rect 1438 1879 1439 1883
rect 1443 1879 1444 1883
rect 1448 1879 1450 1888
rect 1524 1884 1526 1966
rect 1574 1952 1580 1953
rect 1574 1948 1575 1952
rect 1579 1948 1580 1952
rect 1574 1947 1580 1948
rect 1662 1952 1668 1953
rect 1662 1948 1663 1952
rect 1667 1948 1668 1952
rect 1662 1947 1668 1948
rect 1535 1946 1539 1947
rect 1535 1941 1539 1942
rect 1575 1946 1579 1947
rect 1575 1941 1579 1942
rect 1623 1946 1627 1947
rect 1623 1941 1627 1942
rect 1663 1946 1667 1947
rect 1663 1941 1667 1942
rect 1711 1946 1715 1947
rect 1711 1941 1715 1942
rect 1534 1940 1540 1941
rect 1534 1936 1535 1940
rect 1539 1936 1540 1940
rect 1534 1935 1540 1936
rect 1622 1940 1628 1941
rect 1622 1936 1623 1940
rect 1627 1936 1628 1940
rect 1622 1935 1628 1936
rect 1710 1940 1716 1941
rect 1710 1936 1711 1940
rect 1715 1936 1716 1940
rect 1710 1935 1716 1936
rect 1736 1920 1738 1994
rect 1780 1972 1782 2002
rect 1840 2000 1842 2009
rect 1838 1999 1844 2000
rect 1838 1995 1839 1999
rect 1843 1995 1844 1999
rect 1838 1994 1844 1995
rect 1864 1972 1866 2022
rect 1936 2015 1938 2032
rect 1944 2028 1946 2106
rect 1974 2100 1980 2101
rect 1974 2096 1975 2100
rect 1979 2096 1980 2100
rect 1974 2095 1980 2096
rect 2046 2100 2052 2101
rect 2046 2096 2047 2100
rect 2051 2096 2052 2100
rect 2046 2095 2052 2096
rect 1976 2091 1978 2095
rect 2048 2091 2050 2095
rect 1975 2090 1979 2091
rect 1975 2085 1979 2086
rect 2015 2090 2019 2091
rect 2015 2085 2019 2086
rect 2047 2090 2051 2091
rect 2047 2085 2051 2086
rect 2014 2084 2020 2085
rect 2014 2080 2015 2084
rect 2019 2080 2020 2084
rect 2014 2079 2020 2080
rect 2056 2064 2058 2150
rect 2112 2148 2114 2157
rect 2138 2155 2144 2156
rect 2138 2151 2139 2155
rect 2143 2151 2144 2155
rect 2138 2150 2144 2151
rect 2110 2147 2116 2148
rect 2110 2143 2111 2147
rect 2115 2143 2116 2147
rect 2110 2142 2116 2143
rect 2140 2120 2142 2150
rect 2176 2148 2178 2157
rect 2202 2155 2208 2156
rect 2202 2151 2203 2155
rect 2207 2151 2208 2155
rect 2202 2150 2208 2151
rect 2174 2147 2180 2148
rect 2174 2143 2175 2147
rect 2179 2143 2180 2147
rect 2174 2142 2180 2143
rect 2204 2120 2206 2150
rect 2240 2148 2242 2157
rect 2238 2147 2244 2148
rect 2238 2143 2239 2147
rect 2243 2143 2244 2147
rect 2238 2142 2244 2143
rect 2268 2120 2270 2162
rect 2279 2157 2283 2158
rect 2311 2162 2315 2163
rect 2311 2157 2315 2158
rect 2312 2148 2314 2157
rect 2320 2156 2322 2198
rect 2358 2177 2364 2178
rect 2358 2173 2359 2177
rect 2363 2173 2364 2177
rect 2358 2172 2364 2173
rect 2360 2163 2362 2172
rect 2368 2168 2370 2258
rect 2406 2251 2412 2252
rect 2406 2247 2407 2251
rect 2411 2247 2412 2251
rect 2406 2246 2412 2247
rect 2408 2231 2410 2246
rect 2407 2230 2411 2231
rect 2407 2225 2411 2226
rect 2408 2218 2410 2225
rect 2406 2217 2412 2218
rect 2406 2213 2407 2217
rect 2411 2213 2412 2217
rect 2406 2212 2412 2213
rect 2406 2200 2412 2201
rect 2406 2196 2407 2200
rect 2411 2196 2412 2200
rect 2406 2195 2412 2196
rect 2366 2167 2372 2168
rect 2366 2163 2367 2167
rect 2371 2163 2372 2167
rect 2408 2163 2410 2195
rect 2359 2162 2363 2163
rect 2366 2162 2372 2163
rect 2407 2162 2411 2163
rect 2359 2157 2363 2158
rect 2407 2157 2411 2158
rect 2318 2155 2324 2156
rect 2318 2151 2319 2155
rect 2323 2151 2324 2155
rect 2318 2150 2324 2151
rect 2338 2155 2344 2156
rect 2338 2151 2339 2155
rect 2343 2151 2344 2155
rect 2338 2150 2344 2151
rect 2310 2147 2316 2148
rect 2310 2143 2311 2147
rect 2315 2143 2316 2147
rect 2310 2142 2316 2143
rect 2340 2120 2342 2150
rect 2360 2148 2362 2157
rect 2358 2147 2364 2148
rect 2358 2143 2359 2147
rect 2363 2143 2364 2147
rect 2358 2142 2364 2143
rect 2408 2125 2410 2157
rect 2406 2124 2412 2125
rect 2406 2120 2407 2124
rect 2411 2120 2412 2124
rect 2138 2119 2144 2120
rect 2138 2115 2139 2119
rect 2143 2115 2144 2119
rect 2138 2114 2144 2115
rect 2202 2119 2208 2120
rect 2202 2115 2203 2119
rect 2207 2115 2208 2119
rect 2202 2114 2208 2115
rect 2266 2119 2272 2120
rect 2266 2115 2267 2119
rect 2271 2115 2272 2119
rect 2266 2114 2272 2115
rect 2338 2119 2344 2120
rect 2338 2115 2339 2119
rect 2343 2115 2344 2119
rect 2338 2114 2344 2115
rect 2366 2119 2372 2120
rect 2406 2119 2412 2120
rect 2366 2115 2367 2119
rect 2371 2115 2372 2119
rect 2366 2114 2372 2115
rect 2110 2100 2116 2101
rect 2110 2096 2111 2100
rect 2115 2096 2116 2100
rect 2110 2095 2116 2096
rect 2174 2100 2180 2101
rect 2174 2096 2175 2100
rect 2179 2096 2180 2100
rect 2174 2095 2180 2096
rect 2238 2100 2244 2101
rect 2238 2096 2239 2100
rect 2243 2096 2244 2100
rect 2238 2095 2244 2096
rect 2310 2100 2316 2101
rect 2310 2096 2311 2100
rect 2315 2096 2316 2100
rect 2310 2095 2316 2096
rect 2358 2100 2364 2101
rect 2358 2096 2359 2100
rect 2363 2096 2364 2100
rect 2358 2095 2364 2096
rect 2112 2091 2114 2095
rect 2176 2091 2178 2095
rect 2240 2091 2242 2095
rect 2312 2091 2314 2095
rect 2360 2091 2362 2095
rect 2095 2090 2099 2091
rect 2095 2085 2099 2086
rect 2111 2090 2115 2091
rect 2111 2085 2115 2086
rect 2167 2090 2171 2091
rect 2167 2085 2171 2086
rect 2175 2090 2179 2091
rect 2175 2085 2179 2086
rect 2239 2090 2243 2091
rect 2239 2085 2243 2086
rect 2311 2090 2315 2091
rect 2311 2085 2315 2086
rect 2359 2090 2363 2091
rect 2359 2085 2363 2086
rect 2094 2084 2100 2085
rect 2094 2080 2095 2084
rect 2099 2080 2100 2084
rect 2094 2079 2100 2080
rect 2166 2084 2172 2085
rect 2166 2080 2167 2084
rect 2171 2080 2172 2084
rect 2166 2079 2172 2080
rect 2238 2084 2244 2085
rect 2238 2080 2239 2084
rect 2243 2080 2244 2084
rect 2238 2079 2244 2080
rect 2310 2084 2316 2085
rect 2310 2080 2311 2084
rect 2315 2080 2316 2084
rect 2310 2079 2316 2080
rect 2358 2084 2364 2085
rect 2358 2080 2359 2084
rect 2363 2080 2364 2084
rect 2358 2079 2364 2080
rect 2006 2063 2012 2064
rect 2006 2059 2007 2063
rect 2011 2059 2012 2063
rect 2006 2058 2012 2059
rect 2054 2063 2060 2064
rect 2054 2059 2055 2063
rect 2059 2059 2060 2063
rect 2054 2058 2060 2059
rect 2158 2063 2164 2064
rect 2158 2059 2159 2063
rect 2163 2059 2164 2063
rect 2158 2058 2164 2059
rect 2182 2063 2188 2064
rect 2182 2059 2183 2063
rect 2187 2059 2188 2063
rect 2182 2058 2188 2059
rect 2274 2063 2280 2064
rect 2274 2059 2275 2063
rect 2279 2059 2280 2063
rect 2274 2058 2280 2059
rect 2008 2028 2010 2058
rect 2102 2055 2108 2056
rect 2102 2051 2103 2055
rect 2107 2051 2108 2055
rect 2102 2050 2108 2051
rect 2014 2037 2020 2038
rect 2014 2033 2015 2037
rect 2019 2033 2020 2037
rect 2014 2032 2020 2033
rect 2094 2037 2100 2038
rect 2094 2033 2095 2037
rect 2099 2033 2100 2037
rect 2094 2032 2100 2033
rect 1942 2027 1948 2028
rect 1942 2023 1943 2027
rect 1947 2023 1948 2027
rect 1942 2022 1948 2023
rect 2006 2027 2012 2028
rect 2006 2023 2007 2027
rect 2011 2023 2012 2027
rect 2006 2022 2012 2023
rect 2016 2015 2018 2032
rect 2096 2015 2098 2032
rect 2104 2028 2106 2050
rect 2160 2028 2162 2058
rect 2166 2037 2172 2038
rect 2166 2033 2167 2037
rect 2171 2033 2172 2037
rect 2166 2032 2172 2033
rect 2102 2027 2108 2028
rect 2102 2023 2103 2027
rect 2107 2023 2108 2027
rect 2102 2022 2108 2023
rect 2158 2027 2164 2028
rect 2158 2023 2159 2027
rect 2163 2023 2164 2027
rect 2158 2022 2164 2023
rect 2168 2015 2170 2032
rect 1919 2014 1923 2015
rect 1919 2009 1923 2010
rect 1935 2014 1939 2015
rect 1935 2009 1939 2010
rect 1999 2014 2003 2015
rect 1999 2009 2003 2010
rect 2015 2014 2019 2015
rect 2015 2009 2019 2010
rect 2071 2014 2075 2015
rect 2071 2009 2075 2010
rect 2095 2014 2099 2015
rect 2095 2009 2099 2010
rect 2135 2014 2139 2015
rect 2135 2009 2139 2010
rect 2167 2014 2171 2015
rect 2167 2009 2171 2010
rect 1920 2000 1922 2009
rect 1926 2007 1932 2008
rect 1926 2003 1927 2007
rect 1931 2003 1932 2007
rect 1926 2002 1932 2003
rect 1946 2007 1952 2008
rect 1946 2003 1947 2007
rect 1951 2003 1952 2007
rect 1946 2002 1952 2003
rect 1918 1999 1924 2000
rect 1918 1995 1919 1999
rect 1923 1995 1924 1999
rect 1918 1994 1924 1995
rect 1928 1980 1930 2002
rect 1926 1979 1932 1980
rect 1926 1975 1927 1979
rect 1931 1975 1932 1979
rect 1926 1974 1932 1975
rect 1948 1972 1950 2002
rect 2000 2000 2002 2009
rect 2072 2000 2074 2009
rect 2122 2007 2128 2008
rect 2122 2003 2123 2007
rect 2127 2003 2128 2007
rect 2122 2002 2128 2003
rect 1998 1999 2004 2000
rect 1998 1995 1999 1999
rect 2003 1995 2004 1999
rect 1998 1994 2004 1995
rect 2070 1999 2076 2000
rect 2070 1995 2071 1999
rect 2075 1995 2076 1999
rect 2070 1994 2076 1995
rect 2124 1972 2126 2002
rect 2136 2000 2138 2009
rect 2184 2008 2186 2058
rect 2238 2037 2244 2038
rect 2238 2033 2239 2037
rect 2243 2033 2244 2037
rect 2238 2032 2244 2033
rect 2240 2015 2242 2032
rect 2276 2028 2278 2058
rect 2310 2037 2316 2038
rect 2310 2033 2311 2037
rect 2315 2033 2316 2037
rect 2310 2032 2316 2033
rect 2358 2037 2364 2038
rect 2358 2033 2359 2037
rect 2363 2033 2364 2037
rect 2358 2032 2364 2033
rect 2274 2027 2280 2028
rect 2274 2023 2275 2027
rect 2279 2023 2280 2027
rect 2274 2022 2280 2023
rect 2312 2015 2314 2032
rect 2342 2027 2348 2028
rect 2342 2023 2343 2027
rect 2347 2023 2348 2027
rect 2342 2022 2348 2023
rect 2191 2014 2195 2015
rect 2191 2009 2195 2010
rect 2239 2014 2243 2015
rect 2239 2009 2243 2010
rect 2255 2014 2259 2015
rect 2255 2009 2259 2010
rect 2311 2014 2315 2015
rect 2311 2009 2315 2010
rect 2319 2014 2323 2015
rect 2319 2009 2323 2010
rect 2174 2007 2180 2008
rect 2174 2003 2175 2007
rect 2179 2003 2180 2007
rect 2174 2002 2180 2003
rect 2182 2007 2188 2008
rect 2182 2003 2183 2007
rect 2187 2003 2188 2007
rect 2182 2002 2188 2003
rect 2134 1999 2140 2000
rect 2134 1995 2135 1999
rect 2139 1995 2140 1999
rect 2134 1994 2140 1995
rect 2176 1972 2178 2002
rect 2192 2000 2194 2009
rect 2256 2000 2258 2009
rect 2320 2000 2322 2009
rect 2334 2007 2340 2008
rect 2334 2003 2335 2007
rect 2339 2003 2340 2007
rect 2334 2002 2340 2003
rect 2190 1999 2196 2000
rect 2190 1995 2191 1999
rect 2195 1995 2196 1999
rect 2190 1994 2196 1995
rect 2254 1999 2260 2000
rect 2254 1995 2255 1999
rect 2259 1995 2260 1999
rect 2254 1994 2260 1995
rect 2318 1999 2324 2000
rect 2318 1995 2319 1999
rect 2323 1995 2324 1999
rect 2318 1994 2324 1995
rect 2336 1980 2338 2002
rect 2334 1979 2340 1980
rect 2334 1975 2335 1979
rect 2339 1975 2340 1979
rect 2334 1974 2340 1975
rect 2344 1972 2346 2022
rect 2360 2015 2362 2032
rect 2368 2028 2370 2114
rect 2406 2107 2412 2108
rect 2406 2103 2407 2107
rect 2411 2103 2412 2107
rect 2406 2102 2412 2103
rect 2408 2091 2410 2102
rect 2407 2090 2411 2091
rect 2407 2085 2411 2086
rect 2408 2078 2410 2085
rect 2406 2077 2412 2078
rect 2406 2073 2407 2077
rect 2411 2073 2412 2077
rect 2406 2072 2412 2073
rect 2406 2060 2412 2061
rect 2406 2056 2407 2060
rect 2411 2056 2412 2060
rect 2406 2055 2412 2056
rect 2366 2027 2372 2028
rect 2366 2023 2367 2027
rect 2371 2023 2372 2027
rect 2366 2022 2372 2023
rect 2408 2015 2410 2055
rect 2359 2014 2363 2015
rect 2359 2009 2363 2010
rect 2407 2014 2411 2015
rect 2407 2009 2411 2010
rect 2360 2000 2362 2009
rect 2382 2007 2388 2008
rect 2382 2003 2383 2007
rect 2387 2003 2388 2007
rect 2382 2002 2388 2003
rect 2358 1999 2364 2000
rect 2358 1995 2359 1999
rect 2363 1995 2364 1999
rect 2358 1994 2364 1995
rect 1778 1971 1784 1972
rect 1778 1967 1779 1971
rect 1783 1967 1784 1971
rect 1778 1966 1784 1967
rect 1862 1971 1868 1972
rect 1862 1967 1863 1971
rect 1867 1967 1868 1971
rect 1862 1966 1868 1967
rect 1946 1971 1952 1972
rect 1946 1967 1947 1971
rect 1951 1967 1952 1971
rect 1946 1966 1952 1967
rect 2122 1971 2128 1972
rect 2122 1967 2123 1971
rect 2127 1967 2128 1971
rect 2122 1966 2128 1967
rect 2174 1971 2180 1972
rect 2174 1967 2175 1971
rect 2179 1967 2180 1971
rect 2174 1966 2180 1967
rect 2230 1971 2236 1972
rect 2230 1967 2231 1971
rect 2235 1967 2236 1971
rect 2230 1966 2236 1967
rect 2342 1971 2348 1972
rect 2342 1967 2343 1971
rect 2347 1967 2348 1971
rect 2342 1966 2348 1967
rect 1750 1952 1756 1953
rect 1750 1948 1751 1952
rect 1755 1948 1756 1952
rect 1750 1947 1756 1948
rect 1838 1952 1844 1953
rect 1838 1948 1839 1952
rect 1843 1948 1844 1952
rect 1838 1947 1844 1948
rect 1918 1952 1924 1953
rect 1918 1948 1919 1952
rect 1923 1948 1924 1952
rect 1918 1947 1924 1948
rect 1998 1952 2004 1953
rect 1998 1948 1999 1952
rect 2003 1948 2004 1952
rect 1998 1947 2004 1948
rect 2070 1952 2076 1953
rect 2070 1948 2071 1952
rect 2075 1948 2076 1952
rect 2070 1947 2076 1948
rect 2134 1952 2140 1953
rect 2134 1948 2135 1952
rect 2139 1948 2140 1952
rect 2134 1947 2140 1948
rect 2190 1952 2196 1953
rect 2190 1948 2191 1952
rect 2195 1948 2196 1952
rect 2190 1947 2196 1948
rect 1751 1946 1755 1947
rect 1751 1941 1755 1942
rect 1791 1946 1795 1947
rect 1791 1941 1795 1942
rect 1839 1946 1843 1947
rect 1839 1941 1843 1942
rect 1863 1946 1867 1947
rect 1863 1941 1867 1942
rect 1919 1946 1923 1947
rect 1919 1941 1923 1942
rect 1935 1946 1939 1947
rect 1935 1941 1939 1942
rect 1999 1946 2003 1947
rect 1999 1941 2003 1942
rect 2007 1946 2011 1947
rect 2007 1941 2011 1942
rect 2071 1946 2075 1947
rect 2071 1941 2075 1942
rect 2079 1946 2083 1947
rect 2079 1941 2083 1942
rect 2135 1946 2139 1947
rect 2135 1941 2139 1942
rect 2151 1946 2155 1947
rect 2151 1941 2155 1942
rect 2191 1946 2195 1947
rect 2191 1941 2195 1942
rect 2223 1946 2227 1947
rect 2223 1941 2227 1942
rect 1790 1940 1796 1941
rect 1790 1936 1791 1940
rect 1795 1936 1796 1940
rect 1790 1935 1796 1936
rect 1862 1940 1868 1941
rect 1862 1936 1863 1940
rect 1867 1936 1868 1940
rect 1862 1935 1868 1936
rect 1934 1940 1940 1941
rect 1934 1936 1935 1940
rect 1939 1936 1940 1940
rect 1934 1935 1940 1936
rect 2006 1940 2012 1941
rect 2006 1936 2007 1940
rect 2011 1936 2012 1940
rect 2006 1935 2012 1936
rect 2078 1940 2084 1941
rect 2078 1936 2079 1940
rect 2083 1936 2084 1940
rect 2078 1935 2084 1936
rect 2150 1940 2156 1941
rect 2150 1936 2151 1940
rect 2155 1936 2156 1940
rect 2150 1935 2156 1936
rect 2222 1940 2228 1941
rect 2222 1936 2223 1940
rect 2227 1936 2228 1940
rect 2222 1935 2228 1936
rect 1702 1919 1708 1920
rect 1702 1915 1703 1919
rect 1707 1915 1708 1919
rect 1702 1914 1708 1915
rect 1734 1919 1740 1920
rect 1734 1915 1735 1919
rect 1739 1915 1740 1919
rect 1734 1914 1740 1915
rect 1854 1919 1860 1920
rect 1854 1915 1855 1919
rect 1859 1915 1860 1919
rect 1854 1914 1860 1915
rect 1926 1919 1932 1920
rect 1926 1915 1927 1919
rect 1931 1915 1932 1919
rect 1926 1914 1932 1915
rect 1962 1919 1968 1920
rect 1962 1915 1963 1919
rect 1967 1915 1968 1919
rect 1962 1914 1968 1915
rect 2142 1919 2148 1920
rect 2142 1915 2143 1919
rect 2147 1915 2148 1919
rect 2142 1914 2148 1915
rect 1534 1893 1540 1894
rect 1534 1889 1535 1893
rect 1539 1889 1540 1893
rect 1534 1888 1540 1889
rect 1622 1893 1628 1894
rect 1622 1889 1623 1893
rect 1627 1889 1628 1893
rect 1622 1888 1628 1889
rect 1522 1883 1528 1884
rect 1522 1879 1523 1883
rect 1527 1879 1528 1883
rect 1536 1879 1538 1888
rect 1624 1879 1626 1888
rect 1704 1884 1706 1914
rect 1798 1911 1804 1912
rect 1798 1907 1799 1911
rect 1803 1907 1804 1911
rect 1798 1906 1804 1907
rect 1710 1893 1716 1894
rect 1710 1889 1711 1893
rect 1715 1889 1716 1893
rect 1710 1888 1716 1889
rect 1790 1893 1796 1894
rect 1790 1889 1791 1893
rect 1795 1889 1796 1893
rect 1790 1888 1796 1889
rect 1702 1883 1708 1884
rect 1702 1879 1703 1883
rect 1707 1879 1708 1883
rect 1712 1879 1714 1888
rect 1792 1879 1794 1888
rect 1800 1884 1802 1906
rect 1856 1884 1858 1914
rect 1862 1893 1868 1894
rect 1862 1889 1863 1893
rect 1867 1889 1868 1893
rect 1862 1888 1868 1889
rect 1798 1883 1804 1884
rect 1798 1879 1799 1883
rect 1803 1879 1804 1883
rect 1066 1878 1072 1879
rect 1279 1878 1283 1879
rect 918 1875 924 1876
rect 918 1871 919 1875
rect 923 1871 924 1875
rect 1279 1873 1283 1874
rect 1303 1878 1307 1879
rect 1303 1873 1307 1874
rect 1311 1878 1315 1879
rect 1311 1873 1315 1874
rect 1359 1878 1363 1879
rect 1359 1873 1363 1874
rect 1415 1878 1419 1879
rect 1438 1878 1444 1879
rect 1447 1878 1451 1879
rect 1415 1873 1419 1874
rect 918 1870 924 1871
rect 1238 1871 1244 1872
rect 718 1864 724 1865
rect 718 1860 719 1864
rect 723 1860 724 1864
rect 718 1859 724 1860
rect 798 1864 804 1865
rect 798 1860 799 1864
rect 803 1860 804 1864
rect 798 1859 804 1860
rect 878 1864 884 1865
rect 878 1860 879 1864
rect 883 1860 884 1864
rect 878 1859 884 1860
rect 720 1851 722 1859
rect 800 1851 802 1859
rect 880 1851 882 1859
rect 719 1850 723 1851
rect 719 1845 723 1846
rect 727 1850 731 1851
rect 727 1845 731 1846
rect 799 1850 803 1851
rect 799 1845 803 1846
rect 823 1850 827 1851
rect 823 1845 827 1846
rect 879 1850 883 1851
rect 879 1845 883 1846
rect 911 1850 915 1851
rect 911 1845 915 1846
rect 726 1844 732 1845
rect 726 1840 727 1844
rect 731 1840 732 1844
rect 726 1839 732 1840
rect 822 1844 828 1845
rect 822 1840 823 1844
rect 827 1840 828 1844
rect 822 1839 828 1840
rect 910 1844 916 1845
rect 910 1840 911 1844
rect 915 1840 916 1844
rect 910 1839 916 1840
rect 430 1823 436 1824
rect 430 1819 431 1823
rect 435 1819 436 1823
rect 430 1818 436 1819
rect 526 1823 532 1824
rect 526 1819 527 1823
rect 531 1819 532 1823
rect 526 1818 532 1819
rect 654 1823 660 1824
rect 654 1819 655 1823
rect 659 1819 660 1823
rect 654 1818 660 1819
rect 350 1797 356 1798
rect 350 1793 351 1797
rect 355 1793 356 1797
rect 350 1792 356 1793
rect 294 1787 300 1788
rect 294 1783 295 1787
rect 299 1783 300 1787
rect 150 1782 156 1783
rect 175 1782 179 1783
rect 182 1782 188 1783
rect 215 1782 219 1783
rect 175 1777 179 1778
rect 215 1777 219 1778
rect 271 1782 275 1783
rect 271 1777 275 1778
rect 287 1782 291 1783
rect 294 1782 300 1783
rect 334 1787 340 1788
rect 334 1783 335 1787
rect 339 1783 340 1787
rect 352 1783 354 1792
rect 432 1788 434 1818
rect 438 1797 444 1798
rect 438 1793 439 1797
rect 443 1793 444 1797
rect 438 1792 444 1793
rect 430 1787 436 1788
rect 430 1783 431 1787
rect 435 1783 436 1787
rect 440 1783 442 1792
rect 528 1788 530 1818
rect 534 1797 540 1798
rect 534 1793 535 1797
rect 539 1793 540 1797
rect 534 1792 540 1793
rect 630 1797 636 1798
rect 630 1793 631 1797
rect 635 1793 636 1797
rect 630 1792 636 1793
rect 726 1797 732 1798
rect 726 1793 727 1797
rect 731 1793 732 1797
rect 726 1792 732 1793
rect 822 1797 828 1798
rect 822 1793 823 1797
rect 827 1793 828 1797
rect 822 1792 828 1793
rect 910 1797 916 1798
rect 910 1793 911 1797
rect 915 1793 916 1797
rect 910 1792 916 1793
rect 526 1787 532 1788
rect 526 1783 527 1787
rect 531 1783 532 1787
rect 536 1783 538 1792
rect 632 1783 634 1792
rect 728 1783 730 1792
rect 778 1787 784 1788
rect 778 1783 779 1787
rect 783 1783 784 1787
rect 824 1783 826 1792
rect 912 1783 914 1792
rect 920 1788 922 1870
rect 1238 1867 1239 1871
rect 1243 1867 1244 1871
rect 1238 1866 1244 1867
rect 958 1864 964 1865
rect 958 1860 959 1864
rect 963 1860 964 1864
rect 958 1859 964 1860
rect 1038 1864 1044 1865
rect 1038 1860 1039 1864
rect 1043 1860 1044 1864
rect 1038 1859 1044 1860
rect 1118 1864 1124 1865
rect 1118 1860 1119 1864
rect 1123 1860 1124 1864
rect 1118 1859 1124 1860
rect 960 1851 962 1859
rect 1040 1851 1042 1859
rect 1120 1851 1122 1859
rect 1240 1851 1242 1866
rect 959 1850 963 1851
rect 959 1845 963 1846
rect 991 1850 995 1851
rect 991 1845 995 1846
rect 1039 1850 1043 1851
rect 1039 1845 1043 1846
rect 1063 1850 1067 1851
rect 1063 1845 1067 1846
rect 1119 1850 1123 1851
rect 1119 1845 1123 1846
rect 1135 1850 1139 1851
rect 1135 1845 1139 1846
rect 1191 1850 1195 1851
rect 1191 1845 1195 1846
rect 1239 1850 1243 1851
rect 1239 1845 1243 1846
rect 990 1844 996 1845
rect 990 1840 991 1844
rect 995 1840 996 1844
rect 990 1839 996 1840
rect 1062 1844 1068 1845
rect 1062 1840 1063 1844
rect 1067 1840 1068 1844
rect 1062 1839 1068 1840
rect 1134 1844 1140 1845
rect 1134 1840 1135 1844
rect 1139 1840 1140 1844
rect 1134 1839 1140 1840
rect 1190 1844 1196 1845
rect 1190 1840 1191 1844
rect 1195 1840 1196 1844
rect 1190 1839 1196 1840
rect 1240 1838 1242 1845
rect 1280 1841 1282 1873
rect 1312 1864 1314 1873
rect 1330 1871 1336 1872
rect 1330 1867 1331 1871
rect 1335 1867 1336 1871
rect 1330 1866 1336 1867
rect 1338 1871 1344 1872
rect 1338 1867 1339 1871
rect 1343 1867 1344 1871
rect 1338 1866 1344 1867
rect 1310 1863 1316 1864
rect 1310 1859 1311 1863
rect 1315 1859 1316 1863
rect 1310 1858 1316 1859
rect 1332 1844 1334 1866
rect 1330 1843 1336 1844
rect 1278 1840 1284 1841
rect 1238 1837 1244 1838
rect 1238 1833 1239 1837
rect 1243 1833 1244 1837
rect 1278 1836 1279 1840
rect 1283 1836 1284 1840
rect 1330 1839 1331 1843
rect 1335 1839 1336 1843
rect 1330 1838 1336 1839
rect 1340 1836 1342 1866
rect 1360 1864 1362 1873
rect 1386 1871 1392 1872
rect 1386 1867 1387 1871
rect 1391 1867 1392 1871
rect 1386 1866 1392 1867
rect 1358 1863 1364 1864
rect 1358 1859 1359 1863
rect 1363 1859 1364 1863
rect 1358 1858 1364 1859
rect 1388 1836 1390 1866
rect 1416 1864 1418 1873
rect 1414 1863 1420 1864
rect 1414 1859 1415 1863
rect 1419 1859 1420 1863
rect 1414 1858 1420 1859
rect 1440 1836 1442 1878
rect 1447 1873 1451 1874
rect 1479 1878 1483 1879
rect 1522 1878 1528 1879
rect 1535 1878 1539 1879
rect 1479 1873 1483 1874
rect 1535 1873 1539 1874
rect 1543 1878 1547 1879
rect 1543 1873 1547 1874
rect 1615 1878 1619 1879
rect 1615 1873 1619 1874
rect 1623 1878 1627 1879
rect 1623 1873 1627 1874
rect 1687 1878 1691 1879
rect 1702 1878 1708 1879
rect 1711 1878 1715 1879
rect 1687 1873 1691 1874
rect 1711 1873 1715 1874
rect 1767 1878 1771 1879
rect 1767 1873 1771 1874
rect 1791 1878 1795 1879
rect 1798 1878 1804 1879
rect 1854 1883 1860 1884
rect 1854 1879 1855 1883
rect 1859 1879 1860 1883
rect 1864 1879 1866 1888
rect 1928 1884 1930 1914
rect 1934 1893 1940 1894
rect 1934 1889 1935 1893
rect 1939 1889 1940 1893
rect 1934 1888 1940 1889
rect 1926 1883 1932 1884
rect 1926 1879 1927 1883
rect 1931 1879 1932 1883
rect 1936 1879 1938 1888
rect 1854 1878 1860 1879
rect 1863 1878 1867 1879
rect 1926 1878 1932 1879
rect 1935 1878 1939 1879
rect 1791 1873 1795 1874
rect 1863 1873 1867 1874
rect 1935 1873 1939 1874
rect 1480 1864 1482 1873
rect 1544 1864 1546 1873
rect 1598 1871 1604 1872
rect 1598 1867 1599 1871
rect 1603 1867 1604 1871
rect 1598 1866 1604 1867
rect 1606 1871 1612 1872
rect 1606 1867 1607 1871
rect 1611 1867 1612 1871
rect 1606 1866 1612 1867
rect 1478 1863 1484 1864
rect 1478 1859 1479 1863
rect 1483 1859 1484 1863
rect 1478 1858 1484 1859
rect 1542 1863 1548 1864
rect 1542 1859 1543 1863
rect 1547 1859 1548 1863
rect 1542 1858 1548 1859
rect 1600 1836 1602 1866
rect 1278 1835 1284 1836
rect 1338 1835 1344 1836
rect 1238 1832 1244 1833
rect 1338 1831 1339 1835
rect 1343 1831 1344 1835
rect 1338 1830 1344 1831
rect 1386 1835 1392 1836
rect 1386 1831 1387 1835
rect 1391 1831 1392 1835
rect 1386 1830 1392 1831
rect 1438 1835 1444 1836
rect 1438 1831 1439 1835
rect 1443 1831 1444 1835
rect 1438 1830 1444 1831
rect 1598 1835 1604 1836
rect 1598 1831 1599 1835
rect 1603 1831 1604 1835
rect 1598 1830 1604 1831
rect 982 1823 988 1824
rect 982 1819 983 1823
rect 987 1819 988 1823
rect 982 1818 988 1819
rect 1054 1823 1060 1824
rect 1054 1819 1055 1823
rect 1059 1819 1060 1823
rect 1054 1818 1060 1819
rect 1126 1823 1132 1824
rect 1126 1819 1127 1823
rect 1131 1819 1132 1823
rect 1126 1818 1132 1819
rect 1182 1823 1188 1824
rect 1182 1819 1183 1823
rect 1187 1819 1188 1823
rect 1278 1823 1284 1824
rect 1182 1818 1188 1819
rect 1238 1820 1244 1821
rect 984 1788 986 1818
rect 1038 1815 1044 1816
rect 1038 1811 1039 1815
rect 1043 1811 1044 1815
rect 1038 1810 1044 1811
rect 990 1797 996 1798
rect 990 1793 991 1797
rect 995 1793 996 1797
rect 990 1792 996 1793
rect 918 1787 924 1788
rect 918 1783 919 1787
rect 923 1783 924 1787
rect 982 1787 988 1788
rect 982 1783 983 1787
rect 987 1783 988 1787
rect 992 1783 994 1792
rect 334 1782 340 1783
rect 351 1782 355 1783
rect 287 1777 291 1778
rect 351 1777 355 1778
rect 375 1782 379 1783
rect 430 1782 436 1783
rect 439 1782 443 1783
rect 375 1777 379 1778
rect 439 1777 443 1778
rect 471 1782 475 1783
rect 526 1782 532 1783
rect 535 1782 539 1783
rect 471 1777 475 1778
rect 535 1777 539 1778
rect 567 1782 571 1783
rect 567 1777 571 1778
rect 631 1782 635 1783
rect 631 1777 635 1778
rect 663 1782 667 1783
rect 663 1777 667 1778
rect 727 1782 731 1783
rect 727 1777 731 1778
rect 751 1782 755 1783
rect 778 1782 784 1783
rect 823 1782 827 1783
rect 751 1777 755 1778
rect 142 1775 148 1776
rect 142 1771 143 1775
rect 147 1771 148 1775
rect 142 1770 148 1771
rect 158 1775 164 1776
rect 158 1771 159 1775
rect 163 1771 164 1775
rect 158 1770 164 1771
rect 134 1767 140 1768
rect 134 1763 135 1767
rect 139 1763 140 1767
rect 134 1762 140 1763
rect 110 1744 116 1745
rect 110 1740 111 1744
rect 115 1740 116 1744
rect 160 1740 162 1770
rect 176 1768 178 1777
rect 198 1775 204 1776
rect 198 1771 199 1775
rect 203 1771 204 1775
rect 198 1770 204 1771
rect 174 1767 180 1768
rect 174 1763 175 1767
rect 179 1763 180 1767
rect 174 1762 180 1763
rect 200 1740 202 1770
rect 216 1768 218 1777
rect 242 1775 248 1776
rect 242 1771 243 1775
rect 247 1771 248 1775
rect 242 1770 248 1771
rect 214 1767 220 1768
rect 214 1763 215 1767
rect 219 1763 220 1767
rect 214 1762 220 1763
rect 244 1740 246 1770
rect 288 1768 290 1777
rect 314 1775 320 1776
rect 314 1771 315 1775
rect 319 1771 320 1775
rect 314 1770 320 1771
rect 286 1767 292 1768
rect 286 1763 287 1767
rect 291 1763 292 1767
rect 286 1762 292 1763
rect 316 1740 318 1770
rect 376 1768 378 1777
rect 402 1775 408 1776
rect 402 1771 403 1775
rect 407 1771 408 1775
rect 402 1770 408 1771
rect 374 1767 380 1768
rect 374 1763 375 1767
rect 379 1763 380 1767
rect 374 1762 380 1763
rect 404 1740 406 1770
rect 472 1768 474 1777
rect 498 1775 504 1776
rect 498 1771 499 1775
rect 503 1771 504 1775
rect 498 1770 504 1771
rect 470 1767 476 1768
rect 470 1763 471 1767
rect 475 1763 476 1767
rect 470 1762 476 1763
rect 500 1740 502 1770
rect 568 1768 570 1777
rect 664 1768 666 1777
rect 682 1775 688 1776
rect 682 1771 683 1775
rect 687 1771 688 1775
rect 682 1770 688 1771
rect 690 1775 696 1776
rect 690 1771 691 1775
rect 695 1771 696 1775
rect 690 1770 696 1771
rect 566 1767 572 1768
rect 566 1763 567 1767
rect 571 1763 572 1767
rect 566 1762 572 1763
rect 662 1767 668 1768
rect 662 1763 663 1767
rect 667 1763 668 1767
rect 662 1762 668 1763
rect 684 1748 686 1770
rect 682 1747 688 1748
rect 682 1743 683 1747
rect 687 1743 688 1747
rect 682 1742 688 1743
rect 692 1740 694 1770
rect 752 1768 754 1777
rect 750 1767 756 1768
rect 750 1763 751 1767
rect 755 1763 756 1767
rect 750 1762 756 1763
rect 780 1740 782 1782
rect 823 1777 827 1778
rect 831 1782 835 1783
rect 831 1777 835 1778
rect 903 1782 907 1783
rect 903 1777 907 1778
rect 911 1782 915 1783
rect 918 1782 924 1783
rect 967 1782 971 1783
rect 982 1782 988 1783
rect 991 1782 995 1783
rect 911 1777 915 1778
rect 967 1777 971 1778
rect 991 1777 995 1778
rect 1031 1782 1035 1783
rect 1031 1777 1035 1778
rect 832 1768 834 1777
rect 890 1775 896 1776
rect 890 1771 891 1775
rect 895 1771 896 1775
rect 890 1770 896 1771
rect 830 1767 836 1768
rect 830 1763 831 1767
rect 835 1763 836 1767
rect 830 1762 836 1763
rect 892 1740 894 1770
rect 904 1768 906 1777
rect 954 1775 960 1776
rect 954 1771 955 1775
rect 959 1771 960 1775
rect 954 1770 960 1771
rect 902 1767 908 1768
rect 902 1763 903 1767
rect 907 1763 908 1767
rect 902 1762 908 1763
rect 956 1740 958 1770
rect 968 1768 970 1777
rect 1006 1775 1012 1776
rect 1006 1771 1007 1775
rect 1011 1771 1012 1775
rect 1006 1770 1012 1771
rect 966 1767 972 1768
rect 966 1763 967 1767
rect 971 1763 972 1767
rect 966 1762 972 1763
rect 110 1739 116 1740
rect 158 1739 164 1740
rect 158 1735 159 1739
rect 163 1735 164 1739
rect 158 1734 164 1735
rect 198 1739 204 1740
rect 198 1735 199 1739
rect 203 1735 204 1739
rect 198 1734 204 1735
rect 242 1739 248 1740
rect 242 1735 243 1739
rect 247 1735 248 1739
rect 242 1734 248 1735
rect 314 1739 320 1740
rect 314 1735 315 1739
rect 319 1735 320 1739
rect 314 1734 320 1735
rect 402 1739 408 1740
rect 402 1735 403 1739
rect 407 1735 408 1739
rect 402 1734 408 1735
rect 498 1739 504 1740
rect 498 1735 499 1739
rect 503 1735 504 1739
rect 498 1734 504 1735
rect 690 1739 696 1740
rect 690 1735 691 1739
rect 695 1735 696 1739
rect 690 1734 696 1735
rect 778 1739 784 1740
rect 778 1735 779 1739
rect 783 1735 784 1739
rect 778 1734 784 1735
rect 890 1739 896 1740
rect 890 1735 891 1739
rect 895 1735 896 1739
rect 890 1734 896 1735
rect 954 1739 960 1740
rect 954 1735 955 1739
rect 959 1735 960 1739
rect 954 1734 960 1735
rect 142 1731 148 1732
rect 110 1727 116 1728
rect 110 1723 111 1727
rect 115 1723 116 1727
rect 142 1727 143 1731
rect 147 1727 148 1731
rect 142 1726 148 1727
rect 110 1722 116 1723
rect 112 1711 114 1722
rect 134 1720 140 1721
rect 134 1716 135 1720
rect 139 1716 140 1720
rect 134 1715 140 1716
rect 136 1711 138 1715
rect 111 1710 115 1711
rect 111 1705 115 1706
rect 135 1710 139 1711
rect 135 1705 139 1706
rect 112 1698 114 1705
rect 134 1704 140 1705
rect 134 1700 135 1704
rect 139 1700 140 1704
rect 134 1699 140 1700
rect 110 1697 116 1698
rect 110 1693 111 1697
rect 115 1693 116 1697
rect 110 1692 116 1693
rect 110 1680 116 1681
rect 110 1676 111 1680
rect 115 1676 116 1680
rect 110 1675 116 1676
rect 112 1639 114 1675
rect 134 1657 140 1658
rect 134 1653 135 1657
rect 139 1653 140 1657
rect 134 1652 140 1653
rect 136 1639 138 1652
rect 144 1648 146 1726
rect 174 1720 180 1721
rect 174 1716 175 1720
rect 179 1716 180 1720
rect 174 1715 180 1716
rect 214 1720 220 1721
rect 214 1716 215 1720
rect 219 1716 220 1720
rect 214 1715 220 1716
rect 286 1720 292 1721
rect 286 1716 287 1720
rect 291 1716 292 1720
rect 286 1715 292 1716
rect 374 1720 380 1721
rect 374 1716 375 1720
rect 379 1716 380 1720
rect 374 1715 380 1716
rect 470 1720 476 1721
rect 470 1716 471 1720
rect 475 1716 476 1720
rect 470 1715 476 1716
rect 566 1720 572 1721
rect 566 1716 567 1720
rect 571 1716 572 1720
rect 566 1715 572 1716
rect 662 1720 668 1721
rect 662 1716 663 1720
rect 667 1716 668 1720
rect 662 1715 668 1716
rect 750 1720 756 1721
rect 750 1716 751 1720
rect 755 1716 756 1720
rect 750 1715 756 1716
rect 830 1720 836 1721
rect 830 1716 831 1720
rect 835 1716 836 1720
rect 830 1715 836 1716
rect 902 1720 908 1721
rect 902 1716 903 1720
rect 907 1716 908 1720
rect 902 1715 908 1716
rect 966 1720 972 1721
rect 966 1716 967 1720
rect 971 1716 972 1720
rect 966 1715 972 1716
rect 176 1711 178 1715
rect 216 1711 218 1715
rect 288 1711 290 1715
rect 376 1711 378 1715
rect 472 1711 474 1715
rect 568 1711 570 1715
rect 664 1711 666 1715
rect 752 1711 754 1715
rect 832 1711 834 1715
rect 904 1711 906 1715
rect 968 1711 970 1715
rect 175 1710 179 1711
rect 175 1705 179 1706
rect 215 1710 219 1711
rect 215 1705 219 1706
rect 239 1710 243 1711
rect 239 1705 243 1706
rect 287 1710 291 1711
rect 287 1705 291 1706
rect 319 1710 323 1711
rect 319 1705 323 1706
rect 375 1710 379 1711
rect 375 1705 379 1706
rect 415 1710 419 1711
rect 415 1705 419 1706
rect 471 1710 475 1711
rect 471 1705 475 1706
rect 511 1710 515 1711
rect 511 1705 515 1706
rect 567 1710 571 1711
rect 567 1705 571 1706
rect 615 1710 619 1711
rect 615 1705 619 1706
rect 663 1710 667 1711
rect 663 1705 667 1706
rect 711 1710 715 1711
rect 711 1705 715 1706
rect 751 1710 755 1711
rect 751 1705 755 1706
rect 799 1710 803 1711
rect 799 1705 803 1706
rect 831 1710 835 1711
rect 831 1705 835 1706
rect 879 1710 883 1711
rect 879 1705 883 1706
rect 903 1710 907 1711
rect 903 1705 907 1706
rect 951 1710 955 1711
rect 951 1705 955 1706
rect 967 1710 971 1711
rect 967 1705 971 1706
rect 174 1704 180 1705
rect 174 1700 175 1704
rect 179 1700 180 1704
rect 174 1699 180 1700
rect 238 1704 244 1705
rect 238 1700 239 1704
rect 243 1700 244 1704
rect 238 1699 244 1700
rect 318 1704 324 1705
rect 318 1700 319 1704
rect 323 1700 324 1704
rect 318 1699 324 1700
rect 414 1704 420 1705
rect 414 1700 415 1704
rect 419 1700 420 1704
rect 414 1699 420 1700
rect 510 1704 516 1705
rect 510 1700 511 1704
rect 515 1700 516 1704
rect 510 1699 516 1700
rect 614 1704 620 1705
rect 614 1700 615 1704
rect 619 1700 620 1704
rect 614 1699 620 1700
rect 710 1704 716 1705
rect 710 1700 711 1704
rect 715 1700 716 1704
rect 710 1699 716 1700
rect 798 1704 804 1705
rect 798 1700 799 1704
rect 803 1700 804 1704
rect 798 1699 804 1700
rect 878 1704 884 1705
rect 878 1700 879 1704
rect 883 1700 884 1704
rect 878 1699 884 1700
rect 950 1704 956 1705
rect 950 1700 951 1704
rect 955 1700 956 1704
rect 950 1699 956 1700
rect 1008 1692 1010 1770
rect 1032 1768 1034 1777
rect 1040 1776 1042 1810
rect 1056 1788 1058 1818
rect 1062 1797 1068 1798
rect 1062 1793 1063 1797
rect 1067 1793 1068 1797
rect 1062 1792 1068 1793
rect 1054 1787 1060 1788
rect 1054 1783 1055 1787
rect 1059 1783 1060 1787
rect 1064 1783 1066 1792
rect 1128 1788 1130 1818
rect 1134 1797 1140 1798
rect 1134 1793 1135 1797
rect 1139 1793 1140 1797
rect 1134 1792 1140 1793
rect 1126 1787 1132 1788
rect 1126 1783 1127 1787
rect 1131 1783 1132 1787
rect 1136 1783 1138 1792
rect 1184 1788 1186 1818
rect 1238 1816 1239 1820
rect 1243 1816 1244 1820
rect 1278 1819 1279 1823
rect 1283 1819 1284 1823
rect 1278 1818 1284 1819
rect 1238 1815 1244 1816
rect 1190 1797 1196 1798
rect 1190 1793 1191 1797
rect 1195 1793 1196 1797
rect 1190 1792 1196 1793
rect 1182 1787 1188 1788
rect 1182 1783 1183 1787
rect 1187 1783 1188 1787
rect 1192 1783 1194 1792
rect 1240 1783 1242 1815
rect 1280 1807 1282 1818
rect 1310 1816 1316 1817
rect 1310 1812 1311 1816
rect 1315 1812 1316 1816
rect 1310 1811 1316 1812
rect 1358 1816 1364 1817
rect 1358 1812 1359 1816
rect 1363 1812 1364 1816
rect 1358 1811 1364 1812
rect 1414 1816 1420 1817
rect 1414 1812 1415 1816
rect 1419 1812 1420 1816
rect 1414 1811 1420 1812
rect 1478 1816 1484 1817
rect 1478 1812 1479 1816
rect 1483 1812 1484 1816
rect 1478 1811 1484 1812
rect 1542 1816 1548 1817
rect 1542 1812 1543 1816
rect 1547 1812 1548 1816
rect 1542 1811 1548 1812
rect 1312 1807 1314 1811
rect 1360 1807 1362 1811
rect 1416 1807 1418 1811
rect 1480 1807 1482 1811
rect 1544 1807 1546 1811
rect 1279 1806 1283 1807
rect 1279 1801 1283 1802
rect 1311 1806 1315 1807
rect 1311 1801 1315 1802
rect 1359 1806 1363 1807
rect 1359 1801 1363 1802
rect 1407 1806 1411 1807
rect 1407 1801 1411 1802
rect 1415 1806 1419 1807
rect 1415 1801 1419 1802
rect 1471 1806 1475 1807
rect 1471 1801 1475 1802
rect 1479 1806 1483 1807
rect 1479 1801 1483 1802
rect 1535 1806 1539 1807
rect 1535 1801 1539 1802
rect 1543 1806 1547 1807
rect 1543 1801 1547 1802
rect 1599 1806 1603 1807
rect 1599 1801 1603 1802
rect 1280 1794 1282 1801
rect 1406 1800 1412 1801
rect 1406 1796 1407 1800
rect 1411 1796 1412 1800
rect 1406 1795 1412 1796
rect 1470 1800 1476 1801
rect 1470 1796 1471 1800
rect 1475 1796 1476 1800
rect 1470 1795 1476 1796
rect 1534 1800 1540 1801
rect 1534 1796 1535 1800
rect 1539 1796 1540 1800
rect 1534 1795 1540 1796
rect 1598 1800 1604 1801
rect 1598 1796 1599 1800
rect 1603 1796 1604 1800
rect 1598 1795 1604 1796
rect 1278 1793 1284 1794
rect 1278 1789 1279 1793
rect 1283 1789 1284 1793
rect 1278 1788 1284 1789
rect 1054 1782 1060 1783
rect 1063 1782 1067 1783
rect 1063 1777 1067 1778
rect 1087 1782 1091 1783
rect 1126 1782 1132 1783
rect 1135 1782 1139 1783
rect 1087 1777 1091 1778
rect 1135 1777 1139 1778
rect 1151 1782 1155 1783
rect 1182 1782 1188 1783
rect 1191 1782 1195 1783
rect 1151 1777 1155 1778
rect 1191 1777 1195 1778
rect 1239 1782 1243 1783
rect 1608 1780 1610 1866
rect 1616 1864 1618 1873
rect 1688 1864 1690 1873
rect 1754 1871 1760 1872
rect 1754 1867 1755 1871
rect 1759 1867 1760 1871
rect 1754 1866 1760 1867
rect 1614 1863 1620 1864
rect 1614 1859 1615 1863
rect 1619 1859 1620 1863
rect 1614 1858 1620 1859
rect 1686 1863 1692 1864
rect 1686 1859 1687 1863
rect 1691 1859 1692 1863
rect 1686 1858 1692 1859
rect 1756 1836 1758 1866
rect 1768 1864 1770 1873
rect 1850 1871 1856 1872
rect 1850 1867 1851 1871
rect 1855 1867 1856 1871
rect 1850 1866 1856 1867
rect 1766 1863 1772 1864
rect 1766 1859 1767 1863
rect 1771 1859 1772 1863
rect 1766 1858 1772 1859
rect 1852 1836 1854 1866
rect 1864 1864 1866 1873
rect 1964 1872 1966 1914
rect 2014 1911 2020 1912
rect 2014 1907 2015 1911
rect 2019 1907 2020 1911
rect 2014 1906 2020 1907
rect 2006 1893 2012 1894
rect 2006 1889 2007 1893
rect 2011 1889 2012 1893
rect 2006 1888 2012 1889
rect 2008 1879 2010 1888
rect 2016 1884 2018 1906
rect 2078 1893 2084 1894
rect 2078 1889 2079 1893
rect 2083 1889 2084 1893
rect 2078 1888 2084 1889
rect 2014 1883 2020 1884
rect 2014 1879 2015 1883
rect 2019 1879 2020 1883
rect 2080 1879 2082 1888
rect 2144 1884 2146 1914
rect 2150 1893 2156 1894
rect 2150 1889 2151 1893
rect 2155 1889 2156 1893
rect 2150 1888 2156 1889
rect 2222 1893 2228 1894
rect 2222 1889 2223 1893
rect 2227 1889 2228 1893
rect 2222 1888 2228 1889
rect 2142 1883 2148 1884
rect 2142 1879 2143 1883
rect 2147 1879 2148 1883
rect 2152 1879 2154 1888
rect 2224 1879 2226 1888
rect 2232 1884 2234 1966
rect 2254 1952 2260 1953
rect 2254 1948 2255 1952
rect 2259 1948 2260 1952
rect 2254 1947 2260 1948
rect 2318 1952 2324 1953
rect 2318 1948 2319 1952
rect 2323 1948 2324 1952
rect 2318 1947 2324 1948
rect 2358 1952 2364 1953
rect 2358 1948 2359 1952
rect 2363 1948 2364 1952
rect 2358 1947 2364 1948
rect 2255 1946 2259 1947
rect 2255 1941 2259 1942
rect 2303 1946 2307 1947
rect 2303 1941 2307 1942
rect 2319 1946 2323 1947
rect 2319 1941 2323 1942
rect 2359 1946 2363 1947
rect 2359 1941 2363 1942
rect 2302 1940 2308 1941
rect 2302 1936 2303 1940
rect 2307 1936 2308 1940
rect 2302 1935 2308 1936
rect 2358 1940 2364 1941
rect 2358 1936 2359 1940
rect 2363 1936 2364 1940
rect 2358 1935 2364 1936
rect 2384 1920 2386 2002
rect 2408 1977 2410 2009
rect 2406 1976 2412 1977
rect 2406 1972 2407 1976
rect 2411 1972 2412 1976
rect 2406 1971 2412 1972
rect 2406 1959 2412 1960
rect 2406 1955 2407 1959
rect 2411 1955 2412 1959
rect 2406 1954 2412 1955
rect 2408 1947 2410 1954
rect 2407 1946 2411 1947
rect 2407 1941 2411 1942
rect 2408 1934 2410 1941
rect 2406 1933 2412 1934
rect 2406 1929 2407 1933
rect 2411 1929 2412 1933
rect 2406 1928 2412 1929
rect 2294 1919 2300 1920
rect 2294 1915 2295 1919
rect 2299 1915 2300 1919
rect 2294 1914 2300 1915
rect 2350 1919 2356 1920
rect 2350 1915 2351 1919
rect 2355 1915 2356 1919
rect 2350 1914 2356 1915
rect 2382 1919 2388 1920
rect 2382 1915 2383 1919
rect 2387 1915 2388 1919
rect 2382 1914 2388 1915
rect 2406 1916 2412 1917
rect 2296 1884 2298 1914
rect 2302 1893 2308 1894
rect 2302 1889 2303 1893
rect 2307 1889 2308 1893
rect 2302 1888 2308 1889
rect 2230 1883 2236 1884
rect 2230 1879 2231 1883
rect 2235 1879 2236 1883
rect 1975 1878 1979 1879
rect 1975 1873 1979 1874
rect 2007 1878 2011 1879
rect 2014 1878 2020 1879
rect 2079 1878 2083 1879
rect 2007 1873 2011 1874
rect 2079 1873 2083 1874
rect 2095 1878 2099 1879
rect 2142 1878 2148 1879
rect 2151 1878 2155 1879
rect 2095 1873 2099 1874
rect 2151 1873 2155 1874
rect 2223 1878 2227 1879
rect 2230 1878 2236 1879
rect 2294 1883 2300 1884
rect 2294 1879 2295 1883
rect 2299 1879 2300 1883
rect 2304 1879 2306 1888
rect 2294 1878 2300 1879
rect 2303 1878 2307 1879
rect 2223 1873 2227 1874
rect 2303 1873 2307 1874
rect 1962 1871 1968 1872
rect 1962 1867 1963 1871
rect 1967 1867 1968 1871
rect 1962 1866 1968 1867
rect 1976 1864 1978 1873
rect 2096 1864 2098 1873
rect 2122 1871 2128 1872
rect 2122 1867 2123 1871
rect 2127 1867 2128 1871
rect 2122 1866 2128 1867
rect 1862 1863 1868 1864
rect 1862 1859 1863 1863
rect 1867 1859 1868 1863
rect 1862 1858 1868 1859
rect 1974 1863 1980 1864
rect 1974 1859 1975 1863
rect 1979 1859 1980 1863
rect 1974 1858 1980 1859
rect 2094 1863 2100 1864
rect 2094 1859 2095 1863
rect 2099 1859 2100 1863
rect 2094 1858 2100 1859
rect 2124 1836 2126 1866
rect 2224 1864 2226 1873
rect 2352 1872 2354 1914
rect 2406 1912 2407 1916
rect 2411 1912 2412 1916
rect 2406 1911 2412 1912
rect 2358 1893 2364 1894
rect 2358 1889 2359 1893
rect 2363 1889 2364 1893
rect 2358 1888 2364 1889
rect 2360 1879 2362 1888
rect 2382 1883 2388 1884
rect 2382 1879 2383 1883
rect 2387 1879 2388 1883
rect 2408 1879 2410 1911
rect 2359 1878 2363 1879
rect 2382 1878 2388 1879
rect 2407 1878 2411 1879
rect 2359 1873 2363 1874
rect 2350 1871 2356 1872
rect 2350 1867 2351 1871
rect 2355 1867 2356 1871
rect 2350 1866 2356 1867
rect 2360 1864 2362 1873
rect 2222 1863 2228 1864
rect 2222 1859 2223 1863
rect 2227 1859 2228 1863
rect 2222 1858 2228 1859
rect 2358 1863 2364 1864
rect 2358 1859 2359 1863
rect 2363 1859 2364 1863
rect 2358 1858 2364 1859
rect 2384 1836 2386 1878
rect 2407 1873 2411 1874
rect 2408 1841 2410 1873
rect 2406 1840 2412 1841
rect 2406 1836 2407 1840
rect 2411 1836 2412 1840
rect 1670 1835 1676 1836
rect 1670 1831 1671 1835
rect 1675 1831 1676 1835
rect 1670 1830 1676 1831
rect 1754 1835 1760 1836
rect 1754 1831 1755 1835
rect 1759 1831 1760 1835
rect 1754 1830 1760 1831
rect 1850 1835 1856 1836
rect 1850 1831 1851 1835
rect 1855 1831 1856 1835
rect 1850 1830 1856 1831
rect 2122 1835 2128 1836
rect 2122 1831 2123 1835
rect 2127 1831 2128 1835
rect 2122 1830 2128 1831
rect 2382 1835 2388 1836
rect 2406 1835 2412 1836
rect 2382 1831 2383 1835
rect 2387 1831 2388 1835
rect 2382 1830 2388 1831
rect 1614 1816 1620 1817
rect 1614 1812 1615 1816
rect 1619 1812 1620 1816
rect 1614 1811 1620 1812
rect 1616 1807 1618 1811
rect 1615 1806 1619 1807
rect 1615 1801 1619 1802
rect 1663 1806 1667 1807
rect 1663 1801 1667 1802
rect 1662 1800 1668 1801
rect 1662 1796 1663 1800
rect 1667 1796 1668 1800
rect 1662 1795 1668 1796
rect 1239 1777 1243 1778
rect 1462 1779 1468 1780
rect 1038 1775 1044 1776
rect 1038 1771 1039 1775
rect 1043 1771 1044 1775
rect 1038 1770 1044 1771
rect 1088 1768 1090 1777
rect 1114 1775 1120 1776
rect 1114 1771 1115 1775
rect 1119 1771 1120 1775
rect 1114 1770 1120 1771
rect 1030 1767 1036 1768
rect 1030 1763 1031 1767
rect 1035 1763 1036 1767
rect 1030 1762 1036 1763
rect 1086 1767 1092 1768
rect 1086 1763 1087 1767
rect 1091 1763 1092 1767
rect 1086 1762 1092 1763
rect 1116 1740 1118 1770
rect 1152 1768 1154 1777
rect 1174 1775 1180 1776
rect 1174 1771 1175 1775
rect 1179 1771 1180 1775
rect 1174 1770 1180 1771
rect 1150 1767 1156 1768
rect 1150 1763 1151 1767
rect 1155 1763 1156 1767
rect 1150 1762 1156 1763
rect 1176 1740 1178 1770
rect 1192 1768 1194 1777
rect 1190 1767 1196 1768
rect 1190 1763 1191 1767
rect 1195 1763 1196 1767
rect 1190 1762 1196 1763
rect 1240 1745 1242 1777
rect 1278 1776 1284 1777
rect 1278 1772 1279 1776
rect 1283 1772 1284 1776
rect 1462 1775 1463 1779
rect 1467 1775 1468 1779
rect 1462 1774 1468 1775
rect 1526 1779 1532 1780
rect 1526 1775 1527 1779
rect 1531 1775 1532 1779
rect 1526 1774 1532 1775
rect 1590 1779 1596 1780
rect 1590 1775 1591 1779
rect 1595 1775 1596 1779
rect 1590 1774 1596 1775
rect 1606 1779 1612 1780
rect 1606 1775 1607 1779
rect 1611 1775 1612 1779
rect 1606 1774 1612 1775
rect 1278 1771 1284 1772
rect 1238 1744 1244 1745
rect 1238 1740 1239 1744
rect 1243 1740 1244 1744
rect 1114 1739 1120 1740
rect 1114 1735 1115 1739
rect 1119 1735 1120 1739
rect 1114 1734 1120 1735
rect 1174 1739 1180 1740
rect 1238 1739 1244 1740
rect 1280 1739 1282 1771
rect 1406 1753 1412 1754
rect 1406 1749 1407 1753
rect 1411 1749 1412 1753
rect 1406 1748 1412 1749
rect 1408 1739 1410 1748
rect 1464 1744 1466 1774
rect 1470 1753 1476 1754
rect 1470 1749 1471 1753
rect 1475 1749 1476 1753
rect 1470 1748 1476 1749
rect 1446 1743 1452 1744
rect 1446 1739 1447 1743
rect 1451 1739 1452 1743
rect 1174 1735 1175 1739
rect 1179 1735 1180 1739
rect 1174 1734 1180 1735
rect 1279 1738 1283 1739
rect 1279 1733 1283 1734
rect 1303 1738 1307 1739
rect 1303 1733 1307 1734
rect 1351 1738 1355 1739
rect 1351 1733 1355 1734
rect 1407 1738 1411 1739
rect 1407 1733 1411 1734
rect 1423 1738 1427 1739
rect 1446 1738 1452 1739
rect 1462 1743 1468 1744
rect 1462 1739 1463 1743
rect 1467 1739 1468 1743
rect 1472 1739 1474 1748
rect 1528 1744 1530 1774
rect 1534 1753 1540 1754
rect 1534 1749 1535 1753
rect 1539 1749 1540 1753
rect 1534 1748 1540 1749
rect 1526 1743 1532 1744
rect 1526 1739 1527 1743
rect 1531 1739 1532 1743
rect 1536 1739 1538 1748
rect 1592 1744 1594 1774
rect 1598 1753 1604 1754
rect 1598 1749 1599 1753
rect 1603 1749 1604 1753
rect 1598 1748 1604 1749
rect 1662 1753 1668 1754
rect 1662 1749 1663 1753
rect 1667 1749 1668 1753
rect 1662 1748 1668 1749
rect 1590 1743 1596 1744
rect 1590 1739 1591 1743
rect 1595 1739 1596 1743
rect 1600 1739 1602 1748
rect 1664 1739 1666 1748
rect 1672 1744 1674 1830
rect 2406 1823 2412 1824
rect 2406 1819 2407 1823
rect 2411 1819 2412 1823
rect 2406 1818 2412 1819
rect 1686 1816 1692 1817
rect 1686 1812 1687 1816
rect 1691 1812 1692 1816
rect 1686 1811 1692 1812
rect 1766 1816 1772 1817
rect 1766 1812 1767 1816
rect 1771 1812 1772 1816
rect 1766 1811 1772 1812
rect 1862 1816 1868 1817
rect 1862 1812 1863 1816
rect 1867 1812 1868 1816
rect 1862 1811 1868 1812
rect 1974 1816 1980 1817
rect 1974 1812 1975 1816
rect 1979 1812 1980 1816
rect 1974 1811 1980 1812
rect 2094 1816 2100 1817
rect 2094 1812 2095 1816
rect 2099 1812 2100 1816
rect 2094 1811 2100 1812
rect 2222 1816 2228 1817
rect 2222 1812 2223 1816
rect 2227 1812 2228 1816
rect 2222 1811 2228 1812
rect 2358 1816 2364 1817
rect 2358 1812 2359 1816
rect 2363 1812 2364 1816
rect 2358 1811 2364 1812
rect 1688 1807 1690 1811
rect 1768 1807 1770 1811
rect 1864 1807 1866 1811
rect 1976 1807 1978 1811
rect 2096 1807 2098 1811
rect 2224 1807 2226 1811
rect 2360 1807 2362 1811
rect 2408 1807 2410 1818
rect 1687 1806 1691 1807
rect 1687 1801 1691 1802
rect 1727 1806 1731 1807
rect 1727 1801 1731 1802
rect 1767 1806 1771 1807
rect 1767 1801 1771 1802
rect 1783 1806 1787 1807
rect 1783 1801 1787 1802
rect 1839 1806 1843 1807
rect 1839 1801 1843 1802
rect 1863 1806 1867 1807
rect 1863 1801 1867 1802
rect 1895 1806 1899 1807
rect 1895 1801 1899 1802
rect 1959 1806 1963 1807
rect 1959 1801 1963 1802
rect 1975 1806 1979 1807
rect 1975 1801 1979 1802
rect 2095 1806 2099 1807
rect 2095 1801 2099 1802
rect 2223 1806 2227 1807
rect 2223 1801 2227 1802
rect 2359 1806 2363 1807
rect 2359 1801 2363 1802
rect 2407 1806 2411 1807
rect 2407 1801 2411 1802
rect 1726 1800 1732 1801
rect 1726 1796 1727 1800
rect 1731 1796 1732 1800
rect 1726 1795 1732 1796
rect 1782 1800 1788 1801
rect 1782 1796 1783 1800
rect 1787 1796 1788 1800
rect 1782 1795 1788 1796
rect 1838 1800 1844 1801
rect 1838 1796 1839 1800
rect 1843 1796 1844 1800
rect 1838 1795 1844 1796
rect 1894 1800 1900 1801
rect 1894 1796 1895 1800
rect 1899 1796 1900 1800
rect 1894 1795 1900 1796
rect 1958 1800 1964 1801
rect 1958 1796 1959 1800
rect 1963 1796 1964 1800
rect 1958 1795 1964 1796
rect 2408 1794 2410 1801
rect 2406 1793 2412 1794
rect 2406 1789 2407 1793
rect 2411 1789 2412 1793
rect 2406 1788 2412 1789
rect 1718 1779 1724 1780
rect 1718 1775 1719 1779
rect 1723 1775 1724 1779
rect 1718 1774 1724 1775
rect 1774 1779 1780 1780
rect 1774 1775 1775 1779
rect 1779 1775 1780 1779
rect 1774 1774 1780 1775
rect 1830 1779 1836 1780
rect 1830 1775 1831 1779
rect 1835 1775 1836 1779
rect 1830 1774 1836 1775
rect 1886 1779 1892 1780
rect 1886 1775 1887 1779
rect 1891 1775 1892 1779
rect 1886 1774 1892 1775
rect 1950 1779 1956 1780
rect 1950 1775 1951 1779
rect 1955 1775 1956 1779
rect 1950 1774 1956 1775
rect 2406 1776 2412 1777
rect 1720 1744 1722 1774
rect 1742 1771 1748 1772
rect 1742 1767 1743 1771
rect 1747 1767 1748 1771
rect 1742 1766 1748 1767
rect 1726 1753 1732 1754
rect 1726 1749 1727 1753
rect 1731 1749 1732 1753
rect 1726 1748 1732 1749
rect 1670 1743 1676 1744
rect 1670 1739 1671 1743
rect 1675 1739 1676 1743
rect 1462 1738 1468 1739
rect 1471 1738 1475 1739
rect 1423 1733 1427 1734
rect 1238 1727 1244 1728
rect 1238 1723 1239 1727
rect 1243 1723 1244 1727
rect 1238 1722 1244 1723
rect 1030 1720 1036 1721
rect 1030 1716 1031 1720
rect 1035 1716 1036 1720
rect 1030 1715 1036 1716
rect 1086 1720 1092 1721
rect 1086 1716 1087 1720
rect 1091 1716 1092 1720
rect 1086 1715 1092 1716
rect 1150 1720 1156 1721
rect 1150 1716 1151 1720
rect 1155 1716 1156 1720
rect 1150 1715 1156 1716
rect 1190 1720 1196 1721
rect 1190 1716 1191 1720
rect 1195 1716 1196 1720
rect 1190 1715 1196 1716
rect 1032 1711 1034 1715
rect 1088 1711 1090 1715
rect 1152 1711 1154 1715
rect 1192 1711 1194 1715
rect 1240 1711 1242 1722
rect 1015 1710 1019 1711
rect 1015 1705 1019 1706
rect 1031 1710 1035 1711
rect 1031 1705 1035 1706
rect 1087 1710 1091 1711
rect 1087 1705 1091 1706
rect 1151 1710 1155 1711
rect 1151 1705 1155 1706
rect 1159 1710 1163 1711
rect 1159 1705 1163 1706
rect 1191 1710 1195 1711
rect 1191 1705 1195 1706
rect 1239 1710 1243 1711
rect 1239 1705 1243 1706
rect 1014 1704 1020 1705
rect 1014 1700 1015 1704
rect 1019 1700 1020 1704
rect 1014 1699 1020 1700
rect 1086 1704 1092 1705
rect 1086 1700 1087 1704
rect 1091 1700 1092 1704
rect 1086 1699 1092 1700
rect 1158 1704 1164 1705
rect 1158 1700 1159 1704
rect 1163 1700 1164 1704
rect 1158 1699 1164 1700
rect 1240 1698 1242 1705
rect 1280 1701 1282 1733
rect 1304 1724 1306 1733
rect 1330 1731 1336 1732
rect 1330 1727 1331 1731
rect 1335 1727 1336 1731
rect 1330 1726 1336 1727
rect 1302 1723 1308 1724
rect 1302 1719 1303 1723
rect 1307 1719 1308 1723
rect 1302 1718 1308 1719
rect 1278 1700 1284 1701
rect 1238 1697 1244 1698
rect 1238 1693 1239 1697
rect 1243 1693 1244 1697
rect 1278 1696 1279 1700
rect 1283 1696 1284 1700
rect 1332 1696 1334 1726
rect 1352 1724 1354 1733
rect 1424 1724 1426 1733
rect 1350 1723 1356 1724
rect 1350 1719 1351 1723
rect 1355 1719 1356 1723
rect 1350 1718 1356 1719
rect 1422 1723 1428 1724
rect 1422 1719 1423 1723
rect 1427 1719 1428 1723
rect 1422 1718 1428 1719
rect 1448 1696 1450 1738
rect 1471 1733 1475 1734
rect 1503 1738 1507 1739
rect 1526 1738 1532 1739
rect 1535 1738 1539 1739
rect 1503 1733 1507 1734
rect 1535 1733 1539 1734
rect 1583 1738 1587 1739
rect 1590 1738 1596 1739
rect 1599 1738 1603 1739
rect 1583 1733 1587 1734
rect 1599 1733 1603 1734
rect 1663 1738 1667 1739
rect 1670 1738 1676 1739
rect 1718 1743 1724 1744
rect 1718 1739 1719 1743
rect 1723 1739 1724 1743
rect 1728 1739 1730 1748
rect 1718 1738 1724 1739
rect 1727 1738 1731 1739
rect 1663 1733 1667 1734
rect 1727 1733 1731 1734
rect 1735 1738 1739 1739
rect 1735 1733 1739 1734
rect 1486 1731 1492 1732
rect 1486 1727 1487 1731
rect 1491 1727 1492 1731
rect 1486 1726 1492 1727
rect 1488 1696 1490 1726
rect 1504 1724 1506 1733
rect 1570 1731 1576 1732
rect 1570 1727 1571 1731
rect 1575 1727 1576 1731
rect 1570 1726 1576 1727
rect 1502 1723 1508 1724
rect 1502 1719 1503 1723
rect 1507 1719 1508 1723
rect 1502 1718 1508 1719
rect 1572 1696 1574 1726
rect 1584 1724 1586 1733
rect 1650 1731 1656 1732
rect 1650 1727 1651 1731
rect 1655 1727 1656 1731
rect 1650 1726 1656 1727
rect 1582 1723 1588 1724
rect 1582 1719 1583 1723
rect 1587 1719 1588 1723
rect 1582 1718 1588 1719
rect 1652 1696 1654 1726
rect 1664 1724 1666 1733
rect 1736 1724 1738 1733
rect 1744 1732 1746 1766
rect 1776 1744 1778 1774
rect 1782 1753 1788 1754
rect 1782 1749 1783 1753
rect 1787 1749 1788 1753
rect 1782 1748 1788 1749
rect 1774 1743 1780 1744
rect 1774 1739 1775 1743
rect 1779 1739 1780 1743
rect 1784 1739 1786 1748
rect 1832 1744 1834 1774
rect 1838 1753 1844 1754
rect 1838 1749 1839 1753
rect 1843 1749 1844 1753
rect 1838 1748 1844 1749
rect 1830 1743 1836 1744
rect 1830 1739 1831 1743
rect 1835 1739 1836 1743
rect 1840 1739 1842 1748
rect 1888 1744 1890 1774
rect 1894 1753 1900 1754
rect 1894 1749 1895 1753
rect 1899 1749 1900 1753
rect 1894 1748 1900 1749
rect 1886 1743 1892 1744
rect 1886 1739 1887 1743
rect 1891 1739 1892 1743
rect 1896 1739 1898 1748
rect 1952 1744 1954 1774
rect 2406 1772 2407 1776
rect 2411 1772 2412 1776
rect 2406 1771 2412 1772
rect 1958 1753 1964 1754
rect 1958 1749 1959 1753
rect 1963 1749 1964 1753
rect 1958 1748 1964 1749
rect 1950 1743 1956 1744
rect 1950 1739 1951 1743
rect 1955 1739 1956 1743
rect 1960 1739 1962 1748
rect 2408 1739 2410 1771
rect 1774 1738 1780 1739
rect 1783 1738 1787 1739
rect 1783 1733 1787 1734
rect 1807 1738 1811 1739
rect 1830 1738 1836 1739
rect 1839 1738 1843 1739
rect 1807 1733 1811 1734
rect 1839 1733 1843 1734
rect 1871 1738 1875 1739
rect 1886 1738 1892 1739
rect 1895 1738 1899 1739
rect 1871 1733 1875 1734
rect 1895 1733 1899 1734
rect 1935 1738 1939 1739
rect 1950 1738 1956 1739
rect 1959 1738 1963 1739
rect 1935 1733 1939 1734
rect 1959 1733 1963 1734
rect 1999 1738 2003 1739
rect 1999 1733 2003 1734
rect 2063 1738 2067 1739
rect 2063 1733 2067 1734
rect 2407 1738 2411 1739
rect 2407 1733 2411 1734
rect 1742 1731 1748 1732
rect 1742 1727 1743 1731
rect 1747 1727 1748 1731
rect 1742 1726 1748 1727
rect 1762 1731 1768 1732
rect 1762 1727 1763 1731
rect 1767 1727 1768 1731
rect 1762 1726 1768 1727
rect 1662 1723 1668 1724
rect 1662 1719 1663 1723
rect 1667 1719 1668 1723
rect 1662 1718 1668 1719
rect 1734 1723 1740 1724
rect 1734 1719 1735 1723
rect 1739 1719 1740 1723
rect 1734 1718 1740 1719
rect 1764 1696 1766 1726
rect 1808 1724 1810 1733
rect 1872 1724 1874 1733
rect 1918 1731 1924 1732
rect 1918 1727 1919 1731
rect 1923 1727 1924 1731
rect 1918 1726 1924 1727
rect 1806 1723 1812 1724
rect 1806 1719 1807 1723
rect 1811 1719 1812 1723
rect 1806 1718 1812 1719
rect 1870 1723 1876 1724
rect 1870 1719 1871 1723
rect 1875 1719 1876 1723
rect 1870 1718 1876 1719
rect 1920 1700 1922 1726
rect 1936 1724 1938 1733
rect 1966 1731 1972 1732
rect 1966 1727 1967 1731
rect 1971 1727 1972 1731
rect 1966 1726 1972 1727
rect 1934 1723 1940 1724
rect 1934 1719 1935 1723
rect 1939 1719 1940 1723
rect 1934 1718 1940 1719
rect 1918 1699 1924 1700
rect 1278 1695 1284 1696
rect 1330 1695 1336 1696
rect 1238 1692 1244 1693
rect 1006 1691 1012 1692
rect 1006 1687 1007 1691
rect 1011 1687 1012 1691
rect 1330 1691 1331 1695
rect 1335 1691 1336 1695
rect 1330 1690 1336 1691
rect 1338 1695 1344 1696
rect 1338 1691 1339 1695
rect 1343 1691 1344 1695
rect 1338 1690 1344 1691
rect 1446 1695 1452 1696
rect 1446 1691 1447 1695
rect 1451 1691 1452 1695
rect 1446 1690 1452 1691
rect 1486 1695 1492 1696
rect 1486 1691 1487 1695
rect 1491 1691 1492 1695
rect 1486 1690 1492 1691
rect 1570 1695 1576 1696
rect 1570 1691 1571 1695
rect 1575 1691 1576 1695
rect 1570 1690 1576 1691
rect 1650 1695 1656 1696
rect 1650 1691 1651 1695
rect 1655 1691 1656 1695
rect 1650 1690 1656 1691
rect 1762 1695 1768 1696
rect 1762 1691 1763 1695
rect 1767 1691 1768 1695
rect 1918 1695 1919 1699
rect 1923 1695 1924 1699
rect 1968 1696 1970 1726
rect 2000 1724 2002 1733
rect 2026 1731 2032 1732
rect 2026 1727 2027 1731
rect 2031 1727 2032 1731
rect 2026 1726 2032 1727
rect 1998 1723 2004 1724
rect 1998 1719 1999 1723
rect 2003 1719 2004 1723
rect 1998 1718 2004 1719
rect 2028 1696 2030 1726
rect 2064 1724 2066 1733
rect 2062 1723 2068 1724
rect 2062 1719 2063 1723
rect 2067 1719 2068 1723
rect 2062 1718 2068 1719
rect 2408 1701 2410 1733
rect 2406 1700 2412 1701
rect 2406 1696 2407 1700
rect 2411 1696 2412 1700
rect 1918 1694 1924 1695
rect 1962 1695 1970 1696
rect 1762 1690 1768 1691
rect 1962 1691 1963 1695
rect 1967 1692 1970 1695
rect 2026 1695 2032 1696
rect 2406 1695 2412 1696
rect 1967 1691 1968 1692
rect 1962 1690 1968 1691
rect 2026 1691 2027 1695
rect 2031 1691 2032 1695
rect 2026 1690 2032 1691
rect 1006 1686 1012 1687
rect 162 1683 168 1684
rect 162 1679 163 1683
rect 167 1679 168 1683
rect 162 1678 168 1679
rect 230 1683 236 1684
rect 230 1679 231 1683
rect 235 1679 236 1683
rect 230 1678 236 1679
rect 310 1683 316 1684
rect 310 1679 311 1683
rect 315 1679 316 1683
rect 310 1678 316 1679
rect 406 1683 412 1684
rect 406 1679 407 1683
rect 411 1679 412 1683
rect 406 1678 412 1679
rect 502 1683 508 1684
rect 502 1679 503 1683
rect 507 1679 508 1683
rect 502 1678 508 1679
rect 606 1683 612 1684
rect 606 1679 607 1683
rect 611 1679 612 1683
rect 606 1678 612 1679
rect 622 1683 628 1684
rect 622 1679 623 1683
rect 627 1679 628 1683
rect 622 1678 628 1679
rect 790 1683 796 1684
rect 790 1679 791 1683
rect 795 1679 796 1683
rect 790 1678 796 1679
rect 870 1683 876 1684
rect 870 1679 871 1683
rect 875 1679 876 1683
rect 870 1678 876 1679
rect 942 1683 948 1684
rect 942 1679 943 1683
rect 947 1679 948 1683
rect 942 1678 948 1679
rect 1006 1683 1012 1684
rect 1006 1679 1007 1683
rect 1011 1679 1012 1683
rect 1006 1678 1012 1679
rect 1078 1683 1084 1684
rect 1078 1679 1079 1683
rect 1083 1679 1084 1683
rect 1078 1678 1084 1679
rect 1150 1683 1156 1684
rect 1150 1679 1151 1683
rect 1155 1679 1156 1683
rect 1278 1683 1284 1684
rect 1150 1678 1156 1679
rect 1238 1680 1244 1681
rect 164 1648 166 1678
rect 174 1657 180 1658
rect 174 1653 175 1657
rect 179 1653 180 1657
rect 174 1652 180 1653
rect 142 1647 148 1648
rect 142 1643 143 1647
rect 147 1643 148 1647
rect 142 1642 148 1643
rect 162 1647 168 1648
rect 162 1643 163 1647
rect 167 1643 168 1647
rect 162 1642 168 1643
rect 176 1639 178 1652
rect 232 1648 234 1678
rect 279 1660 283 1661
rect 238 1657 244 1658
rect 238 1653 239 1657
rect 243 1653 244 1657
rect 279 1655 283 1656
rect 238 1652 244 1653
rect 230 1647 236 1648
rect 230 1643 231 1647
rect 235 1643 236 1647
rect 230 1642 236 1643
rect 240 1639 242 1652
rect 111 1638 115 1639
rect 111 1633 115 1634
rect 135 1638 139 1639
rect 135 1633 139 1634
rect 175 1638 179 1639
rect 175 1633 179 1634
rect 239 1638 243 1639
rect 239 1633 243 1634
rect 271 1638 275 1639
rect 271 1633 275 1634
rect 112 1601 114 1633
rect 272 1624 274 1633
rect 280 1632 282 1655
rect 312 1648 314 1678
rect 318 1657 324 1658
rect 318 1653 319 1657
rect 323 1653 324 1657
rect 318 1652 324 1653
rect 310 1647 316 1648
rect 310 1643 311 1647
rect 315 1643 316 1647
rect 310 1642 316 1643
rect 320 1639 322 1652
rect 408 1648 410 1678
rect 414 1657 420 1658
rect 414 1653 415 1657
rect 419 1653 420 1657
rect 414 1652 420 1653
rect 406 1647 412 1648
rect 406 1643 407 1647
rect 411 1643 412 1647
rect 406 1642 412 1643
rect 416 1639 418 1652
rect 504 1648 506 1678
rect 510 1657 516 1658
rect 510 1653 511 1657
rect 515 1653 516 1657
rect 510 1652 516 1653
rect 502 1647 508 1648
rect 502 1643 503 1647
rect 507 1643 508 1647
rect 502 1642 508 1643
rect 512 1639 514 1652
rect 608 1648 610 1678
rect 624 1661 626 1678
rect 623 1660 627 1661
rect 614 1657 620 1658
rect 614 1653 615 1657
rect 619 1653 620 1657
rect 623 1655 627 1656
rect 710 1657 716 1658
rect 614 1652 620 1653
rect 710 1653 711 1657
rect 715 1653 716 1657
rect 710 1652 716 1653
rect 606 1647 612 1648
rect 606 1643 607 1647
rect 611 1643 612 1647
rect 606 1642 612 1643
rect 616 1639 618 1652
rect 712 1639 714 1652
rect 792 1648 794 1678
rect 798 1657 804 1658
rect 798 1653 799 1657
rect 803 1653 804 1657
rect 798 1652 804 1653
rect 790 1647 796 1648
rect 790 1643 791 1647
rect 795 1643 796 1647
rect 790 1642 796 1643
rect 766 1639 772 1640
rect 800 1639 802 1652
rect 872 1648 874 1678
rect 878 1657 884 1658
rect 878 1653 879 1657
rect 883 1653 884 1657
rect 878 1652 884 1653
rect 870 1647 876 1648
rect 870 1643 871 1647
rect 875 1643 876 1647
rect 870 1642 876 1643
rect 880 1639 882 1652
rect 944 1648 946 1678
rect 950 1657 956 1658
rect 950 1653 951 1657
rect 955 1653 956 1657
rect 950 1652 956 1653
rect 942 1647 948 1648
rect 942 1643 943 1647
rect 947 1643 948 1647
rect 942 1642 948 1643
rect 952 1639 954 1652
rect 1008 1648 1010 1678
rect 1014 1657 1020 1658
rect 1014 1653 1015 1657
rect 1019 1653 1020 1657
rect 1014 1652 1020 1653
rect 1006 1647 1012 1648
rect 1006 1643 1007 1647
rect 1011 1643 1012 1647
rect 1006 1642 1012 1643
rect 1016 1639 1018 1652
rect 1080 1648 1082 1678
rect 1086 1657 1092 1658
rect 1086 1653 1087 1657
rect 1091 1653 1092 1657
rect 1086 1652 1092 1653
rect 1078 1647 1084 1648
rect 1078 1643 1079 1647
rect 1083 1643 1084 1647
rect 1078 1642 1084 1643
rect 1022 1639 1028 1640
rect 1088 1639 1090 1652
rect 1152 1648 1154 1678
rect 1238 1676 1239 1680
rect 1243 1676 1244 1680
rect 1278 1679 1279 1683
rect 1283 1679 1284 1683
rect 1278 1678 1284 1679
rect 1238 1675 1244 1676
rect 1158 1657 1164 1658
rect 1158 1653 1159 1657
rect 1163 1653 1164 1657
rect 1158 1652 1164 1653
rect 1150 1647 1156 1648
rect 1150 1643 1151 1647
rect 1155 1643 1156 1647
rect 1150 1642 1156 1643
rect 1160 1639 1162 1652
rect 1240 1639 1242 1675
rect 1280 1671 1282 1678
rect 1302 1676 1308 1677
rect 1302 1672 1303 1676
rect 1307 1672 1308 1676
rect 1302 1671 1308 1672
rect 1279 1670 1283 1671
rect 1279 1665 1283 1666
rect 1303 1670 1307 1671
rect 1303 1665 1307 1666
rect 1280 1658 1282 1665
rect 1302 1664 1308 1665
rect 1302 1660 1303 1664
rect 1307 1660 1308 1664
rect 1302 1659 1308 1660
rect 1278 1657 1284 1658
rect 1278 1653 1279 1657
rect 1283 1653 1284 1657
rect 1278 1652 1284 1653
rect 1278 1640 1284 1641
rect 311 1638 315 1639
rect 311 1633 315 1634
rect 319 1638 323 1639
rect 319 1633 323 1634
rect 359 1638 363 1639
rect 359 1633 363 1634
rect 415 1638 419 1639
rect 415 1633 419 1634
rect 471 1638 475 1639
rect 471 1633 475 1634
rect 511 1638 515 1639
rect 511 1633 515 1634
rect 535 1638 539 1639
rect 535 1633 539 1634
rect 599 1638 603 1639
rect 599 1633 603 1634
rect 615 1638 619 1639
rect 615 1633 619 1634
rect 663 1638 667 1639
rect 663 1633 667 1634
rect 711 1638 715 1639
rect 711 1633 715 1634
rect 719 1638 723 1639
rect 766 1635 767 1639
rect 771 1635 772 1639
rect 766 1634 772 1635
rect 775 1638 779 1639
rect 719 1633 723 1634
rect 278 1631 284 1632
rect 278 1627 279 1631
rect 283 1627 284 1631
rect 278 1626 284 1627
rect 298 1631 304 1632
rect 298 1627 299 1631
rect 303 1627 304 1631
rect 298 1626 304 1627
rect 270 1623 276 1624
rect 270 1619 271 1623
rect 275 1619 276 1623
rect 270 1618 276 1619
rect 110 1600 116 1601
rect 110 1596 111 1600
rect 115 1596 116 1600
rect 300 1596 302 1626
rect 312 1624 314 1633
rect 338 1631 344 1632
rect 338 1627 339 1631
rect 343 1627 344 1631
rect 338 1626 344 1627
rect 310 1623 316 1624
rect 310 1619 311 1623
rect 315 1619 316 1623
rect 310 1618 316 1619
rect 340 1596 342 1626
rect 360 1624 362 1633
rect 394 1631 400 1632
rect 394 1627 395 1631
rect 399 1627 400 1631
rect 394 1626 400 1627
rect 358 1623 364 1624
rect 358 1619 359 1623
rect 363 1619 364 1623
rect 358 1618 364 1619
rect 396 1596 398 1626
rect 416 1624 418 1633
rect 442 1631 448 1632
rect 442 1627 443 1631
rect 447 1627 448 1631
rect 442 1626 448 1627
rect 414 1623 420 1624
rect 414 1619 415 1623
rect 419 1619 420 1623
rect 414 1618 420 1619
rect 444 1596 446 1626
rect 472 1624 474 1633
rect 498 1631 504 1632
rect 498 1627 499 1631
rect 503 1627 504 1631
rect 498 1626 504 1627
rect 470 1623 476 1624
rect 470 1619 471 1623
rect 475 1619 476 1623
rect 470 1618 476 1619
rect 500 1596 502 1626
rect 536 1624 538 1633
rect 562 1631 568 1632
rect 562 1627 563 1631
rect 567 1627 568 1631
rect 562 1626 568 1627
rect 534 1623 540 1624
rect 534 1619 535 1623
rect 539 1619 540 1623
rect 534 1618 540 1619
rect 564 1596 566 1626
rect 600 1624 602 1633
rect 664 1624 666 1633
rect 690 1631 696 1632
rect 690 1627 691 1631
rect 695 1627 696 1631
rect 690 1626 696 1627
rect 598 1623 604 1624
rect 598 1619 599 1623
rect 603 1619 604 1623
rect 598 1618 604 1619
rect 662 1623 668 1624
rect 662 1619 663 1623
rect 667 1619 668 1623
rect 662 1618 668 1619
rect 692 1596 694 1626
rect 720 1624 722 1633
rect 746 1631 752 1632
rect 746 1627 747 1631
rect 751 1627 752 1631
rect 746 1626 752 1627
rect 718 1623 724 1624
rect 718 1619 719 1623
rect 723 1619 724 1623
rect 718 1618 724 1619
rect 748 1596 750 1626
rect 110 1595 116 1596
rect 298 1595 304 1596
rect 298 1591 299 1595
rect 303 1591 304 1595
rect 298 1590 304 1591
rect 338 1595 344 1596
rect 338 1591 339 1595
rect 343 1591 344 1595
rect 338 1590 344 1591
rect 394 1595 400 1596
rect 394 1591 395 1595
rect 399 1591 400 1595
rect 394 1590 400 1591
rect 442 1595 448 1596
rect 442 1591 443 1595
rect 447 1591 448 1595
rect 442 1590 448 1591
rect 498 1595 504 1596
rect 498 1591 499 1595
rect 503 1591 504 1595
rect 498 1590 504 1591
rect 562 1595 568 1596
rect 562 1591 563 1595
rect 567 1591 568 1595
rect 562 1590 568 1591
rect 690 1595 696 1596
rect 690 1591 691 1595
rect 695 1591 696 1595
rect 690 1590 696 1591
rect 746 1595 752 1596
rect 746 1591 747 1595
rect 751 1591 752 1595
rect 746 1590 752 1591
rect 768 1588 770 1634
rect 775 1633 779 1634
rect 799 1638 803 1639
rect 799 1633 803 1634
rect 831 1638 835 1639
rect 831 1633 835 1634
rect 879 1638 883 1639
rect 879 1633 883 1634
rect 887 1638 891 1639
rect 887 1633 891 1634
rect 943 1638 947 1639
rect 943 1633 947 1634
rect 951 1638 955 1639
rect 951 1633 955 1634
rect 999 1638 1003 1639
rect 999 1633 1003 1634
rect 1015 1638 1019 1639
rect 1022 1635 1023 1639
rect 1027 1635 1028 1639
rect 1022 1634 1028 1635
rect 1087 1638 1091 1639
rect 1015 1633 1019 1634
rect 776 1624 778 1633
rect 810 1631 816 1632
rect 810 1627 811 1631
rect 815 1627 816 1631
rect 810 1626 816 1627
rect 774 1623 780 1624
rect 774 1619 775 1623
rect 779 1619 780 1623
rect 774 1618 780 1619
rect 812 1596 814 1626
rect 832 1624 834 1633
rect 858 1631 864 1632
rect 858 1627 859 1631
rect 863 1627 864 1631
rect 858 1626 864 1627
rect 830 1623 836 1624
rect 830 1619 831 1623
rect 835 1619 836 1623
rect 830 1618 836 1619
rect 860 1596 862 1626
rect 888 1624 890 1633
rect 914 1631 920 1632
rect 914 1627 915 1631
rect 919 1627 920 1631
rect 914 1626 920 1627
rect 886 1623 892 1624
rect 886 1619 887 1623
rect 891 1619 892 1623
rect 886 1618 892 1619
rect 916 1596 918 1626
rect 944 1624 946 1633
rect 970 1631 976 1632
rect 970 1627 971 1631
rect 975 1627 976 1631
rect 970 1626 976 1627
rect 942 1623 948 1624
rect 942 1619 943 1623
rect 947 1619 948 1623
rect 942 1618 948 1619
rect 972 1596 974 1626
rect 1000 1624 1002 1633
rect 998 1623 1004 1624
rect 998 1619 999 1623
rect 1003 1619 1004 1623
rect 998 1618 1004 1619
rect 1024 1596 1026 1634
rect 1087 1633 1091 1634
rect 1159 1638 1163 1639
rect 1159 1633 1163 1634
rect 1239 1638 1243 1639
rect 1278 1636 1279 1640
rect 1283 1636 1284 1640
rect 1278 1635 1284 1636
rect 1239 1633 1243 1634
rect 1240 1601 1242 1633
rect 1280 1603 1282 1635
rect 1302 1617 1308 1618
rect 1302 1613 1303 1617
rect 1307 1613 1308 1617
rect 1302 1612 1308 1613
rect 1304 1603 1306 1612
rect 1340 1608 1342 1690
rect 1822 1687 1828 1688
rect 1822 1683 1823 1687
rect 1827 1683 1828 1687
rect 1822 1682 1828 1683
rect 2406 1683 2412 1684
rect 1350 1676 1356 1677
rect 1350 1672 1351 1676
rect 1355 1672 1356 1676
rect 1350 1671 1356 1672
rect 1422 1676 1428 1677
rect 1422 1672 1423 1676
rect 1427 1672 1428 1676
rect 1422 1671 1428 1672
rect 1502 1676 1508 1677
rect 1502 1672 1503 1676
rect 1507 1672 1508 1676
rect 1502 1671 1508 1672
rect 1582 1676 1588 1677
rect 1582 1672 1583 1676
rect 1587 1672 1588 1676
rect 1582 1671 1588 1672
rect 1662 1676 1668 1677
rect 1662 1672 1663 1676
rect 1667 1672 1668 1676
rect 1662 1671 1668 1672
rect 1734 1676 1740 1677
rect 1734 1672 1735 1676
rect 1739 1672 1740 1676
rect 1734 1671 1740 1672
rect 1806 1676 1812 1677
rect 1806 1672 1807 1676
rect 1811 1672 1812 1676
rect 1806 1671 1812 1672
rect 1351 1670 1355 1671
rect 1351 1665 1355 1666
rect 1359 1670 1363 1671
rect 1359 1665 1363 1666
rect 1423 1670 1427 1671
rect 1423 1665 1427 1666
rect 1447 1670 1451 1671
rect 1447 1665 1451 1666
rect 1503 1670 1507 1671
rect 1503 1665 1507 1666
rect 1543 1670 1547 1671
rect 1543 1665 1547 1666
rect 1583 1670 1587 1671
rect 1583 1665 1587 1666
rect 1639 1670 1643 1671
rect 1639 1665 1643 1666
rect 1663 1670 1667 1671
rect 1663 1665 1667 1666
rect 1727 1670 1731 1671
rect 1727 1665 1731 1666
rect 1735 1670 1739 1671
rect 1735 1665 1739 1666
rect 1807 1670 1811 1671
rect 1807 1665 1811 1666
rect 1815 1670 1819 1671
rect 1815 1665 1819 1666
rect 1358 1664 1364 1665
rect 1358 1660 1359 1664
rect 1363 1660 1364 1664
rect 1358 1659 1364 1660
rect 1446 1664 1452 1665
rect 1446 1660 1447 1664
rect 1451 1660 1452 1664
rect 1446 1659 1452 1660
rect 1542 1664 1548 1665
rect 1542 1660 1543 1664
rect 1547 1660 1548 1664
rect 1542 1659 1548 1660
rect 1638 1664 1644 1665
rect 1638 1660 1639 1664
rect 1643 1660 1644 1664
rect 1638 1659 1644 1660
rect 1726 1664 1732 1665
rect 1726 1660 1727 1664
rect 1731 1660 1732 1664
rect 1726 1659 1732 1660
rect 1814 1664 1820 1665
rect 1814 1660 1815 1664
rect 1819 1660 1820 1664
rect 1814 1659 1820 1660
rect 1350 1643 1356 1644
rect 1350 1639 1351 1643
rect 1355 1639 1356 1643
rect 1350 1638 1356 1639
rect 1438 1643 1444 1644
rect 1438 1639 1439 1643
rect 1443 1639 1444 1643
rect 1438 1638 1444 1639
rect 1454 1643 1460 1644
rect 1454 1639 1455 1643
rect 1459 1639 1460 1643
rect 1454 1638 1460 1639
rect 1630 1643 1636 1644
rect 1630 1639 1631 1643
rect 1635 1639 1636 1643
rect 1630 1638 1636 1639
rect 1718 1643 1724 1644
rect 1718 1639 1719 1643
rect 1723 1639 1724 1643
rect 1718 1638 1724 1639
rect 1352 1608 1354 1638
rect 1358 1617 1364 1618
rect 1358 1613 1359 1617
rect 1363 1613 1364 1617
rect 1358 1612 1364 1613
rect 1338 1607 1344 1608
rect 1338 1603 1339 1607
rect 1343 1603 1344 1607
rect 1279 1602 1283 1603
rect 1238 1600 1244 1601
rect 1238 1596 1239 1600
rect 1243 1596 1244 1600
rect 1279 1597 1283 1598
rect 1303 1602 1307 1603
rect 1303 1597 1307 1598
rect 1327 1602 1331 1603
rect 1338 1602 1344 1603
rect 1350 1607 1356 1608
rect 1350 1603 1351 1607
rect 1355 1603 1356 1607
rect 1360 1603 1362 1612
rect 1440 1608 1442 1638
rect 1446 1617 1452 1618
rect 1446 1613 1447 1617
rect 1451 1613 1452 1617
rect 1446 1612 1452 1613
rect 1438 1607 1444 1608
rect 1438 1603 1439 1607
rect 1443 1603 1444 1607
rect 1448 1603 1450 1612
rect 1350 1602 1356 1603
rect 1359 1602 1363 1603
rect 1327 1597 1331 1598
rect 1359 1597 1363 1598
rect 1399 1602 1403 1603
rect 1438 1602 1444 1603
rect 1447 1602 1451 1603
rect 1399 1597 1403 1598
rect 1447 1597 1451 1598
rect 810 1595 816 1596
rect 810 1591 811 1595
rect 815 1591 816 1595
rect 810 1590 816 1591
rect 858 1595 864 1596
rect 858 1591 859 1595
rect 863 1591 864 1595
rect 858 1590 864 1591
rect 914 1595 920 1596
rect 914 1591 915 1595
rect 919 1591 920 1595
rect 914 1590 920 1591
rect 970 1595 976 1596
rect 970 1591 971 1595
rect 975 1591 976 1595
rect 970 1590 976 1591
rect 1022 1595 1028 1596
rect 1238 1595 1244 1596
rect 1022 1591 1023 1595
rect 1027 1591 1028 1595
rect 1022 1590 1028 1591
rect 346 1587 352 1588
rect 110 1583 116 1584
rect 110 1579 111 1583
rect 115 1579 116 1583
rect 346 1583 347 1587
rect 351 1583 352 1587
rect 346 1582 352 1583
rect 766 1587 772 1588
rect 766 1583 767 1587
rect 771 1583 772 1587
rect 766 1582 772 1583
rect 950 1587 956 1588
rect 950 1583 951 1587
rect 955 1583 956 1587
rect 950 1582 956 1583
rect 1238 1583 1244 1584
rect 110 1578 116 1579
rect 112 1563 114 1578
rect 270 1576 276 1577
rect 270 1572 271 1576
rect 275 1572 276 1576
rect 270 1571 276 1572
rect 310 1576 316 1577
rect 310 1572 311 1576
rect 315 1572 316 1576
rect 310 1571 316 1572
rect 272 1563 274 1571
rect 312 1563 314 1571
rect 111 1562 115 1563
rect 111 1557 115 1558
rect 271 1562 275 1563
rect 271 1557 275 1558
rect 311 1562 315 1563
rect 311 1557 315 1558
rect 327 1562 331 1563
rect 327 1557 331 1558
rect 112 1550 114 1557
rect 326 1556 332 1557
rect 326 1552 327 1556
rect 331 1552 332 1556
rect 326 1551 332 1552
rect 110 1549 116 1550
rect 110 1545 111 1549
rect 115 1545 116 1549
rect 110 1544 116 1545
rect 110 1532 116 1533
rect 110 1528 111 1532
rect 115 1528 116 1532
rect 110 1527 116 1528
rect 112 1455 114 1527
rect 326 1509 332 1510
rect 326 1505 327 1509
rect 331 1505 332 1509
rect 326 1504 332 1505
rect 328 1455 330 1504
rect 348 1500 350 1582
rect 358 1576 364 1577
rect 358 1572 359 1576
rect 363 1572 364 1576
rect 358 1571 364 1572
rect 414 1576 420 1577
rect 414 1572 415 1576
rect 419 1572 420 1576
rect 414 1571 420 1572
rect 470 1576 476 1577
rect 470 1572 471 1576
rect 475 1572 476 1576
rect 470 1571 476 1572
rect 534 1576 540 1577
rect 534 1572 535 1576
rect 539 1572 540 1576
rect 534 1571 540 1572
rect 598 1576 604 1577
rect 598 1572 599 1576
rect 603 1572 604 1576
rect 598 1571 604 1572
rect 662 1576 668 1577
rect 662 1572 663 1576
rect 667 1572 668 1576
rect 662 1571 668 1572
rect 718 1576 724 1577
rect 718 1572 719 1576
rect 723 1572 724 1576
rect 718 1571 724 1572
rect 774 1576 780 1577
rect 774 1572 775 1576
rect 779 1572 780 1576
rect 774 1571 780 1572
rect 830 1576 836 1577
rect 830 1572 831 1576
rect 835 1572 836 1576
rect 830 1571 836 1572
rect 886 1576 892 1577
rect 886 1572 887 1576
rect 891 1572 892 1576
rect 886 1571 892 1572
rect 942 1576 948 1577
rect 942 1572 943 1576
rect 947 1572 948 1576
rect 942 1571 948 1572
rect 360 1563 362 1571
rect 416 1563 418 1571
rect 472 1563 474 1571
rect 536 1563 538 1571
rect 600 1563 602 1571
rect 664 1563 666 1571
rect 720 1563 722 1571
rect 776 1563 778 1571
rect 832 1563 834 1571
rect 888 1563 890 1571
rect 944 1563 946 1571
rect 359 1562 363 1563
rect 359 1557 363 1558
rect 367 1562 371 1563
rect 367 1557 371 1558
rect 407 1562 411 1563
rect 407 1557 411 1558
rect 415 1562 419 1563
rect 415 1557 419 1558
rect 447 1562 451 1563
rect 447 1557 451 1558
rect 471 1562 475 1563
rect 471 1557 475 1558
rect 487 1562 491 1563
rect 487 1557 491 1558
rect 527 1562 531 1563
rect 527 1557 531 1558
rect 535 1562 539 1563
rect 535 1557 539 1558
rect 567 1562 571 1563
rect 567 1557 571 1558
rect 599 1562 603 1563
rect 599 1557 603 1558
rect 607 1562 611 1563
rect 607 1557 611 1558
rect 647 1562 651 1563
rect 647 1557 651 1558
rect 663 1562 667 1563
rect 663 1557 667 1558
rect 687 1562 691 1563
rect 687 1557 691 1558
rect 719 1562 723 1563
rect 719 1557 723 1558
rect 727 1562 731 1563
rect 727 1557 731 1558
rect 767 1562 771 1563
rect 767 1557 771 1558
rect 775 1562 779 1563
rect 775 1557 779 1558
rect 807 1562 811 1563
rect 807 1557 811 1558
rect 831 1562 835 1563
rect 831 1557 835 1558
rect 847 1562 851 1563
rect 847 1557 851 1558
rect 887 1562 891 1563
rect 887 1557 891 1558
rect 927 1562 931 1563
rect 927 1557 931 1558
rect 943 1562 947 1563
rect 943 1557 947 1558
rect 366 1556 372 1557
rect 366 1552 367 1556
rect 371 1552 372 1556
rect 366 1551 372 1552
rect 406 1556 412 1557
rect 406 1552 407 1556
rect 411 1552 412 1556
rect 406 1551 412 1552
rect 446 1556 452 1557
rect 446 1552 447 1556
rect 451 1552 452 1556
rect 446 1551 452 1552
rect 486 1556 492 1557
rect 486 1552 487 1556
rect 491 1552 492 1556
rect 486 1551 492 1552
rect 526 1556 532 1557
rect 526 1552 527 1556
rect 531 1552 532 1556
rect 526 1551 532 1552
rect 566 1556 572 1557
rect 566 1552 567 1556
rect 571 1552 572 1556
rect 566 1551 572 1552
rect 606 1556 612 1557
rect 606 1552 607 1556
rect 611 1552 612 1556
rect 606 1551 612 1552
rect 646 1556 652 1557
rect 646 1552 647 1556
rect 651 1552 652 1556
rect 646 1551 652 1552
rect 686 1556 692 1557
rect 686 1552 687 1556
rect 691 1552 692 1556
rect 686 1551 692 1552
rect 726 1556 732 1557
rect 726 1552 727 1556
rect 731 1552 732 1556
rect 726 1551 732 1552
rect 766 1556 772 1557
rect 766 1552 767 1556
rect 771 1552 772 1556
rect 766 1551 772 1552
rect 806 1556 812 1557
rect 806 1552 807 1556
rect 811 1552 812 1556
rect 806 1551 812 1552
rect 846 1556 852 1557
rect 846 1552 847 1556
rect 851 1552 852 1556
rect 846 1551 852 1552
rect 886 1556 892 1557
rect 886 1552 887 1556
rect 891 1552 892 1556
rect 886 1551 892 1552
rect 926 1556 932 1557
rect 926 1552 927 1556
rect 931 1552 932 1556
rect 926 1551 932 1552
rect 952 1536 954 1582
rect 1238 1579 1239 1583
rect 1243 1579 1244 1583
rect 1238 1578 1244 1579
rect 998 1576 1004 1577
rect 998 1572 999 1576
rect 1003 1572 1004 1576
rect 998 1571 1004 1572
rect 1000 1563 1002 1571
rect 1240 1563 1242 1578
rect 1280 1565 1282 1597
rect 1328 1588 1330 1597
rect 1382 1595 1388 1596
rect 1382 1591 1383 1595
rect 1387 1591 1388 1595
rect 1382 1590 1388 1591
rect 1326 1587 1332 1588
rect 1326 1583 1327 1587
rect 1331 1583 1332 1587
rect 1326 1582 1332 1583
rect 1278 1564 1284 1565
rect 999 1562 1003 1563
rect 999 1557 1003 1558
rect 1239 1562 1243 1563
rect 1278 1560 1279 1564
rect 1283 1560 1284 1564
rect 1384 1560 1386 1590
rect 1400 1588 1402 1597
rect 1456 1596 1458 1638
rect 1542 1617 1548 1618
rect 1542 1613 1543 1617
rect 1547 1613 1548 1617
rect 1542 1612 1548 1613
rect 1506 1607 1512 1608
rect 1506 1603 1507 1607
rect 1511 1603 1512 1607
rect 1544 1603 1546 1612
rect 1632 1608 1634 1638
rect 1638 1617 1644 1618
rect 1638 1613 1639 1617
rect 1643 1613 1644 1617
rect 1638 1612 1644 1613
rect 1630 1607 1636 1608
rect 1630 1603 1631 1607
rect 1635 1603 1636 1607
rect 1640 1603 1642 1612
rect 1720 1608 1722 1638
rect 1726 1617 1732 1618
rect 1726 1613 1727 1617
rect 1731 1613 1732 1617
rect 1726 1612 1732 1613
rect 1814 1617 1820 1618
rect 1814 1613 1815 1617
rect 1819 1613 1820 1617
rect 1814 1612 1820 1613
rect 1718 1607 1724 1608
rect 1718 1603 1719 1607
rect 1723 1603 1724 1607
rect 1728 1603 1730 1612
rect 1816 1603 1818 1612
rect 1824 1608 1826 1682
rect 2406 1679 2407 1683
rect 2411 1679 2412 1683
rect 2406 1678 2412 1679
rect 1870 1676 1876 1677
rect 1870 1672 1871 1676
rect 1875 1672 1876 1676
rect 1870 1671 1876 1672
rect 1934 1676 1940 1677
rect 1934 1672 1935 1676
rect 1939 1672 1940 1676
rect 1934 1671 1940 1672
rect 1998 1676 2004 1677
rect 1998 1672 1999 1676
rect 2003 1672 2004 1676
rect 1998 1671 2004 1672
rect 2062 1676 2068 1677
rect 2062 1672 2063 1676
rect 2067 1672 2068 1676
rect 2062 1671 2068 1672
rect 2408 1671 2410 1678
rect 1871 1670 1875 1671
rect 1871 1665 1875 1666
rect 1895 1670 1899 1671
rect 1895 1665 1899 1666
rect 1935 1670 1939 1671
rect 1935 1665 1939 1666
rect 1967 1670 1971 1671
rect 1967 1665 1971 1666
rect 1999 1670 2003 1671
rect 1999 1665 2003 1666
rect 2031 1670 2035 1671
rect 2031 1665 2035 1666
rect 2063 1670 2067 1671
rect 2063 1665 2067 1666
rect 2095 1670 2099 1671
rect 2095 1665 2099 1666
rect 2159 1670 2163 1671
rect 2159 1665 2163 1666
rect 2223 1670 2227 1671
rect 2223 1665 2227 1666
rect 2407 1670 2411 1671
rect 2407 1665 2411 1666
rect 1894 1664 1900 1665
rect 1894 1660 1895 1664
rect 1899 1660 1900 1664
rect 1894 1659 1900 1660
rect 1966 1664 1972 1665
rect 1966 1660 1967 1664
rect 1971 1660 1972 1664
rect 1966 1659 1972 1660
rect 2030 1664 2036 1665
rect 2030 1660 2031 1664
rect 2035 1660 2036 1664
rect 2030 1659 2036 1660
rect 2094 1664 2100 1665
rect 2094 1660 2095 1664
rect 2099 1660 2100 1664
rect 2094 1659 2100 1660
rect 2158 1664 2164 1665
rect 2158 1660 2159 1664
rect 2163 1660 2164 1664
rect 2158 1659 2164 1660
rect 2222 1664 2228 1665
rect 2222 1660 2223 1664
rect 2227 1660 2228 1664
rect 2222 1659 2228 1660
rect 2408 1658 2410 1665
rect 2406 1657 2412 1658
rect 2406 1653 2407 1657
rect 2411 1653 2412 1657
rect 2406 1652 2412 1653
rect 1886 1643 1892 1644
rect 1886 1639 1887 1643
rect 1891 1639 1892 1643
rect 1886 1638 1892 1639
rect 1958 1643 1964 1644
rect 1958 1639 1959 1643
rect 1963 1639 1964 1643
rect 1958 1638 1964 1639
rect 2022 1643 2028 1644
rect 2022 1639 2023 1643
rect 2027 1639 2028 1643
rect 2022 1638 2028 1639
rect 2086 1643 2092 1644
rect 2086 1639 2087 1643
rect 2091 1639 2092 1643
rect 2086 1638 2092 1639
rect 2150 1643 2156 1644
rect 2150 1639 2151 1643
rect 2155 1639 2156 1643
rect 2150 1638 2156 1639
rect 2206 1643 2212 1644
rect 2206 1639 2207 1643
rect 2211 1639 2212 1643
rect 2206 1638 2212 1639
rect 2406 1640 2412 1641
rect 1888 1608 1890 1638
rect 1918 1635 1924 1636
rect 1918 1631 1919 1635
rect 1923 1631 1924 1635
rect 1918 1630 1924 1631
rect 1894 1617 1900 1618
rect 1894 1613 1895 1617
rect 1899 1613 1900 1617
rect 1894 1612 1900 1613
rect 1822 1607 1828 1608
rect 1822 1603 1823 1607
rect 1827 1603 1828 1607
rect 1886 1607 1892 1608
rect 1886 1603 1887 1607
rect 1891 1603 1892 1607
rect 1896 1603 1898 1612
rect 1479 1602 1483 1603
rect 1506 1602 1512 1603
rect 1543 1602 1547 1603
rect 1479 1597 1483 1598
rect 1454 1595 1460 1596
rect 1454 1591 1455 1595
rect 1459 1591 1460 1595
rect 1454 1590 1460 1591
rect 1480 1588 1482 1597
rect 1398 1587 1404 1588
rect 1398 1583 1399 1587
rect 1403 1583 1404 1587
rect 1398 1582 1404 1583
rect 1478 1587 1484 1588
rect 1478 1583 1479 1587
rect 1483 1583 1484 1587
rect 1478 1582 1484 1583
rect 1508 1560 1510 1602
rect 1543 1597 1547 1598
rect 1567 1602 1571 1603
rect 1630 1602 1636 1603
rect 1639 1602 1643 1603
rect 1567 1597 1571 1598
rect 1639 1597 1643 1598
rect 1655 1602 1659 1603
rect 1718 1602 1724 1603
rect 1727 1602 1731 1603
rect 1655 1597 1659 1598
rect 1727 1597 1731 1598
rect 1743 1602 1747 1603
rect 1743 1597 1747 1598
rect 1815 1602 1819 1603
rect 1822 1602 1828 1603
rect 1831 1602 1835 1603
rect 1886 1602 1892 1603
rect 1895 1602 1899 1603
rect 1815 1597 1819 1598
rect 1831 1597 1835 1598
rect 1895 1597 1899 1598
rect 1911 1602 1915 1603
rect 1911 1597 1915 1598
rect 1554 1595 1560 1596
rect 1554 1591 1555 1595
rect 1559 1591 1560 1595
rect 1554 1590 1560 1591
rect 1556 1560 1558 1590
rect 1568 1588 1570 1597
rect 1656 1588 1658 1597
rect 1718 1595 1724 1596
rect 1718 1591 1719 1595
rect 1723 1591 1724 1595
rect 1718 1590 1724 1591
rect 1566 1587 1572 1588
rect 1566 1583 1567 1587
rect 1571 1583 1572 1587
rect 1566 1582 1572 1583
rect 1654 1587 1660 1588
rect 1654 1583 1655 1587
rect 1659 1583 1660 1587
rect 1654 1582 1660 1583
rect 1720 1560 1722 1590
rect 1744 1588 1746 1597
rect 1832 1588 1834 1597
rect 1912 1588 1914 1597
rect 1920 1596 1922 1630
rect 1960 1608 1962 1638
rect 1966 1617 1972 1618
rect 1966 1613 1967 1617
rect 1971 1613 1972 1617
rect 1966 1612 1972 1613
rect 1958 1607 1964 1608
rect 1958 1603 1959 1607
rect 1963 1603 1964 1607
rect 1968 1603 1970 1612
rect 2024 1608 2026 1638
rect 2030 1617 2036 1618
rect 2030 1613 2031 1617
rect 2035 1613 2036 1617
rect 2030 1612 2036 1613
rect 2022 1607 2028 1608
rect 2022 1603 2023 1607
rect 2027 1603 2028 1607
rect 2032 1603 2034 1612
rect 2088 1608 2090 1638
rect 2094 1617 2100 1618
rect 2094 1613 2095 1617
rect 2099 1613 2100 1617
rect 2094 1612 2100 1613
rect 2086 1607 2092 1608
rect 2086 1603 2087 1607
rect 2091 1603 2092 1607
rect 2096 1603 2098 1612
rect 2152 1608 2154 1638
rect 2158 1617 2164 1618
rect 2158 1613 2159 1617
rect 2163 1613 2164 1617
rect 2158 1612 2164 1613
rect 2150 1607 2156 1608
rect 2150 1603 2151 1607
rect 2155 1603 2156 1607
rect 2160 1603 2162 1612
rect 2208 1608 2210 1638
rect 2406 1636 2407 1640
rect 2411 1636 2412 1640
rect 2406 1635 2412 1636
rect 2222 1617 2228 1618
rect 2222 1613 2223 1617
rect 2227 1613 2228 1617
rect 2222 1612 2228 1613
rect 2206 1607 2212 1608
rect 2206 1603 2207 1607
rect 2211 1603 2212 1607
rect 2224 1603 2226 1612
rect 2408 1603 2410 1635
rect 1958 1602 1964 1603
rect 1967 1602 1971 1603
rect 1967 1597 1971 1598
rect 1983 1602 1987 1603
rect 2022 1602 2028 1603
rect 2031 1602 2035 1603
rect 1983 1597 1987 1598
rect 2031 1597 2035 1598
rect 2047 1602 2051 1603
rect 2086 1602 2092 1603
rect 2095 1602 2099 1603
rect 2047 1597 2051 1598
rect 2095 1597 2099 1598
rect 2111 1602 2115 1603
rect 2150 1602 2156 1603
rect 2159 1602 2163 1603
rect 2111 1597 2115 1598
rect 2159 1597 2163 1598
rect 2167 1602 2171 1603
rect 2206 1602 2212 1603
rect 2215 1602 2219 1603
rect 2167 1597 2171 1598
rect 2215 1597 2219 1598
rect 2223 1602 2227 1603
rect 2223 1597 2227 1598
rect 2271 1602 2275 1603
rect 2271 1597 2275 1598
rect 2319 1602 2323 1603
rect 2319 1597 2323 1598
rect 2359 1602 2363 1603
rect 2359 1597 2363 1598
rect 2407 1602 2411 1603
rect 2407 1597 2411 1598
rect 1918 1595 1924 1596
rect 1918 1591 1919 1595
rect 1923 1591 1924 1595
rect 1918 1590 1924 1591
rect 1938 1595 1944 1596
rect 1938 1591 1939 1595
rect 1943 1591 1944 1595
rect 1938 1590 1944 1591
rect 1742 1587 1748 1588
rect 1742 1583 1743 1587
rect 1747 1583 1748 1587
rect 1742 1582 1748 1583
rect 1830 1587 1836 1588
rect 1830 1583 1831 1587
rect 1835 1583 1836 1587
rect 1830 1582 1836 1583
rect 1910 1587 1916 1588
rect 1910 1583 1911 1587
rect 1915 1583 1916 1587
rect 1910 1582 1916 1583
rect 1940 1560 1942 1590
rect 1984 1588 1986 1597
rect 2010 1595 2016 1596
rect 2010 1591 2011 1595
rect 2015 1591 2016 1595
rect 2010 1590 2016 1591
rect 1982 1587 1988 1588
rect 1982 1583 1983 1587
rect 1987 1583 1988 1587
rect 1982 1582 1988 1583
rect 2012 1560 2014 1590
rect 2048 1588 2050 1597
rect 2074 1595 2080 1596
rect 2074 1591 2075 1595
rect 2079 1591 2080 1595
rect 2074 1590 2080 1591
rect 2046 1587 2052 1588
rect 2046 1583 2047 1587
rect 2051 1583 2052 1587
rect 2046 1582 2052 1583
rect 2076 1560 2078 1590
rect 2112 1588 2114 1597
rect 2150 1595 2156 1596
rect 2150 1591 2151 1595
rect 2155 1591 2156 1595
rect 2150 1590 2156 1591
rect 2110 1587 2116 1588
rect 2110 1583 2111 1587
rect 2115 1583 2116 1587
rect 2110 1582 2116 1583
rect 2152 1560 2154 1590
rect 2168 1588 2170 1597
rect 2194 1595 2200 1596
rect 2194 1591 2195 1595
rect 2199 1591 2200 1595
rect 2194 1590 2200 1591
rect 2166 1587 2172 1588
rect 2166 1583 2167 1587
rect 2171 1583 2172 1587
rect 2166 1582 2172 1583
rect 2196 1560 2198 1590
rect 2216 1588 2218 1597
rect 2242 1595 2248 1596
rect 2242 1591 2243 1595
rect 2247 1591 2248 1595
rect 2242 1590 2248 1591
rect 2214 1587 2220 1588
rect 2214 1583 2215 1587
rect 2219 1583 2220 1587
rect 2214 1582 2220 1583
rect 2244 1560 2246 1590
rect 2272 1588 2274 1597
rect 2298 1595 2304 1596
rect 2298 1591 2299 1595
rect 2303 1591 2304 1595
rect 2298 1590 2304 1591
rect 2270 1587 2276 1588
rect 2270 1583 2271 1587
rect 2275 1583 2276 1587
rect 2270 1582 2276 1583
rect 2300 1560 2302 1590
rect 2320 1588 2322 1597
rect 2346 1595 2352 1596
rect 2346 1591 2347 1595
rect 2351 1591 2352 1595
rect 2346 1590 2352 1591
rect 2318 1587 2324 1588
rect 2318 1583 2319 1587
rect 2323 1583 2324 1587
rect 2318 1582 2324 1583
rect 2348 1560 2350 1590
rect 2360 1588 2362 1597
rect 2358 1587 2364 1588
rect 2358 1583 2359 1587
rect 2363 1583 2364 1587
rect 2358 1582 2364 1583
rect 2408 1565 2410 1597
rect 2406 1564 2412 1565
rect 2406 1560 2407 1564
rect 2411 1560 2412 1564
rect 1278 1559 1284 1560
rect 1342 1559 1348 1560
rect 1239 1557 1243 1558
rect 1240 1550 1242 1557
rect 1342 1555 1343 1559
rect 1347 1555 1348 1559
rect 1342 1554 1348 1555
rect 1382 1559 1388 1560
rect 1382 1555 1383 1559
rect 1387 1555 1388 1559
rect 1382 1554 1388 1555
rect 1506 1559 1512 1560
rect 1506 1555 1507 1559
rect 1511 1555 1512 1559
rect 1506 1554 1512 1555
rect 1554 1559 1560 1560
rect 1554 1555 1555 1559
rect 1559 1555 1560 1559
rect 1554 1554 1560 1555
rect 1718 1559 1724 1560
rect 1718 1555 1719 1559
rect 1723 1555 1724 1559
rect 1718 1554 1724 1555
rect 1938 1559 1944 1560
rect 1938 1555 1939 1559
rect 1943 1555 1944 1559
rect 1938 1554 1944 1555
rect 2010 1559 2016 1560
rect 2010 1555 2011 1559
rect 2015 1555 2016 1559
rect 2010 1554 2016 1555
rect 2074 1559 2080 1560
rect 2074 1555 2075 1559
rect 2079 1555 2080 1559
rect 2074 1554 2080 1555
rect 2150 1559 2156 1560
rect 2150 1555 2151 1559
rect 2155 1555 2156 1559
rect 2150 1554 2156 1555
rect 2194 1559 2200 1560
rect 2194 1555 2195 1559
rect 2199 1555 2200 1559
rect 2194 1554 2200 1555
rect 2242 1559 2248 1560
rect 2242 1555 2243 1559
rect 2247 1555 2248 1559
rect 2242 1554 2248 1555
rect 2298 1559 2304 1560
rect 2298 1555 2299 1559
rect 2303 1555 2304 1559
rect 2298 1554 2304 1555
rect 2346 1559 2352 1560
rect 2406 1559 2412 1560
rect 2346 1555 2347 1559
rect 2351 1555 2352 1559
rect 2346 1554 2352 1555
rect 1238 1549 1244 1550
rect 1238 1545 1239 1549
rect 1243 1545 1244 1549
rect 1238 1544 1244 1545
rect 1278 1547 1284 1548
rect 1278 1543 1279 1547
rect 1283 1543 1284 1547
rect 1278 1542 1284 1543
rect 354 1535 360 1536
rect 354 1531 355 1535
rect 359 1531 360 1535
rect 354 1530 360 1531
rect 394 1535 400 1536
rect 394 1531 395 1535
rect 399 1531 400 1535
rect 394 1530 400 1531
rect 434 1535 440 1536
rect 434 1531 435 1535
rect 439 1531 440 1535
rect 434 1530 440 1531
rect 474 1535 480 1536
rect 474 1531 475 1535
rect 479 1531 480 1535
rect 474 1530 480 1531
rect 514 1535 520 1536
rect 514 1531 515 1535
rect 519 1531 520 1535
rect 514 1530 520 1531
rect 554 1535 560 1536
rect 554 1531 555 1535
rect 559 1531 560 1535
rect 554 1530 560 1531
rect 594 1535 600 1536
rect 594 1531 595 1535
rect 599 1531 600 1535
rect 594 1530 600 1531
rect 634 1535 640 1536
rect 634 1531 635 1535
rect 639 1531 640 1535
rect 634 1530 640 1531
rect 674 1535 680 1536
rect 674 1531 675 1535
rect 679 1531 680 1535
rect 674 1530 680 1531
rect 714 1535 720 1536
rect 714 1531 715 1535
rect 719 1531 720 1535
rect 714 1530 720 1531
rect 754 1535 760 1536
rect 754 1531 755 1535
rect 759 1531 760 1535
rect 754 1530 760 1531
rect 794 1535 800 1536
rect 794 1531 795 1535
rect 799 1531 800 1535
rect 794 1530 800 1531
rect 834 1535 840 1536
rect 834 1531 835 1535
rect 839 1531 840 1535
rect 834 1530 840 1531
rect 874 1535 880 1536
rect 874 1531 875 1535
rect 879 1531 880 1535
rect 874 1530 880 1531
rect 914 1535 920 1536
rect 914 1531 915 1535
rect 919 1531 920 1535
rect 914 1530 920 1531
rect 950 1535 956 1536
rect 950 1531 951 1535
rect 955 1531 956 1535
rect 950 1530 956 1531
rect 1238 1532 1244 1533
rect 356 1500 358 1530
rect 366 1509 372 1510
rect 366 1505 367 1509
rect 371 1505 372 1509
rect 366 1504 372 1505
rect 346 1499 352 1500
rect 346 1495 347 1499
rect 351 1495 352 1499
rect 346 1494 352 1495
rect 354 1499 360 1500
rect 354 1495 355 1499
rect 359 1495 360 1499
rect 354 1494 360 1495
rect 368 1455 370 1504
rect 396 1500 398 1530
rect 406 1509 412 1510
rect 406 1505 407 1509
rect 411 1505 412 1509
rect 406 1504 412 1505
rect 394 1499 400 1500
rect 394 1495 395 1499
rect 399 1495 400 1499
rect 394 1494 400 1495
rect 408 1455 410 1504
rect 436 1500 438 1530
rect 446 1509 452 1510
rect 446 1505 447 1509
rect 451 1505 452 1509
rect 446 1504 452 1505
rect 434 1499 440 1500
rect 434 1495 435 1499
rect 439 1495 440 1499
rect 434 1494 440 1495
rect 448 1455 450 1504
rect 476 1500 478 1530
rect 486 1509 492 1510
rect 486 1505 487 1509
rect 491 1505 492 1509
rect 486 1504 492 1505
rect 474 1499 480 1500
rect 474 1495 475 1499
rect 479 1495 480 1499
rect 474 1494 480 1495
rect 488 1455 490 1504
rect 516 1500 518 1530
rect 526 1509 532 1510
rect 526 1505 527 1509
rect 531 1505 532 1509
rect 526 1504 532 1505
rect 514 1499 520 1500
rect 514 1495 515 1499
rect 519 1495 520 1499
rect 514 1494 520 1495
rect 528 1455 530 1504
rect 556 1500 558 1530
rect 566 1509 572 1510
rect 566 1505 567 1509
rect 571 1505 572 1509
rect 566 1504 572 1505
rect 554 1499 560 1500
rect 554 1495 555 1499
rect 559 1495 560 1499
rect 554 1494 560 1495
rect 568 1455 570 1504
rect 596 1500 598 1530
rect 606 1509 612 1510
rect 606 1505 607 1509
rect 611 1505 612 1509
rect 606 1504 612 1505
rect 594 1499 600 1500
rect 594 1495 595 1499
rect 599 1495 600 1499
rect 594 1494 600 1495
rect 608 1455 610 1504
rect 636 1500 638 1530
rect 646 1509 652 1510
rect 646 1505 647 1509
rect 651 1505 652 1509
rect 646 1504 652 1505
rect 634 1499 640 1500
rect 634 1495 635 1499
rect 639 1495 640 1499
rect 634 1494 640 1495
rect 648 1455 650 1504
rect 676 1500 678 1530
rect 686 1509 692 1510
rect 686 1505 687 1509
rect 691 1505 692 1509
rect 686 1504 692 1505
rect 674 1499 680 1500
rect 674 1495 675 1499
rect 679 1495 680 1499
rect 674 1494 680 1495
rect 688 1455 690 1504
rect 716 1500 718 1530
rect 726 1509 732 1510
rect 726 1505 727 1509
rect 731 1505 732 1509
rect 726 1504 732 1505
rect 714 1499 720 1500
rect 714 1495 715 1499
rect 719 1495 720 1499
rect 714 1494 720 1495
rect 728 1455 730 1504
rect 756 1500 758 1530
rect 766 1509 772 1510
rect 766 1505 767 1509
rect 771 1505 772 1509
rect 766 1504 772 1505
rect 754 1499 760 1500
rect 754 1495 755 1499
rect 759 1495 760 1499
rect 754 1494 760 1495
rect 768 1455 770 1504
rect 796 1500 798 1530
rect 806 1509 812 1510
rect 806 1505 807 1509
rect 811 1505 812 1509
rect 806 1504 812 1505
rect 794 1499 800 1500
rect 794 1495 795 1499
rect 799 1495 800 1499
rect 794 1494 800 1495
rect 808 1455 810 1504
rect 836 1500 838 1530
rect 846 1509 852 1510
rect 846 1505 847 1509
rect 851 1505 852 1509
rect 846 1504 852 1505
rect 834 1499 840 1500
rect 834 1495 835 1499
rect 839 1495 840 1499
rect 834 1494 840 1495
rect 848 1455 850 1504
rect 876 1500 878 1530
rect 886 1509 892 1510
rect 886 1505 887 1509
rect 891 1505 892 1509
rect 886 1504 892 1505
rect 874 1499 880 1500
rect 874 1495 875 1499
rect 879 1495 880 1499
rect 874 1494 880 1495
rect 888 1455 890 1504
rect 916 1500 918 1530
rect 1238 1528 1239 1532
rect 1243 1528 1244 1532
rect 1280 1531 1282 1542
rect 1326 1540 1332 1541
rect 1326 1536 1327 1540
rect 1331 1536 1332 1540
rect 1326 1535 1332 1536
rect 1328 1531 1330 1535
rect 1238 1527 1244 1528
rect 1279 1530 1283 1531
rect 926 1509 932 1510
rect 926 1505 927 1509
rect 931 1505 932 1509
rect 926 1504 932 1505
rect 914 1499 920 1500
rect 914 1495 915 1499
rect 919 1495 920 1499
rect 914 1494 920 1495
rect 928 1455 930 1504
rect 1240 1455 1242 1527
rect 1279 1525 1283 1526
rect 1327 1530 1331 1531
rect 1327 1525 1331 1526
rect 1335 1530 1339 1531
rect 1335 1525 1339 1526
rect 1280 1518 1282 1525
rect 1334 1524 1340 1525
rect 1334 1520 1335 1524
rect 1339 1520 1340 1524
rect 1334 1519 1340 1520
rect 1278 1517 1284 1518
rect 1278 1513 1279 1517
rect 1283 1513 1284 1517
rect 1278 1512 1284 1513
rect 1278 1500 1284 1501
rect 1278 1496 1279 1500
rect 1283 1496 1284 1500
rect 1278 1495 1284 1496
rect 1280 1463 1282 1495
rect 1334 1477 1340 1478
rect 1334 1473 1335 1477
rect 1339 1473 1340 1477
rect 1334 1472 1340 1473
rect 1336 1463 1338 1472
rect 1344 1468 1346 1554
rect 2222 1551 2228 1552
rect 2222 1547 2223 1551
rect 2227 1547 2228 1551
rect 2222 1546 2228 1547
rect 2406 1547 2412 1548
rect 1398 1540 1404 1541
rect 1398 1536 1399 1540
rect 1403 1536 1404 1540
rect 1398 1535 1404 1536
rect 1478 1540 1484 1541
rect 1478 1536 1479 1540
rect 1483 1536 1484 1540
rect 1478 1535 1484 1536
rect 1566 1540 1572 1541
rect 1566 1536 1567 1540
rect 1571 1536 1572 1540
rect 1566 1535 1572 1536
rect 1654 1540 1660 1541
rect 1654 1536 1655 1540
rect 1659 1536 1660 1540
rect 1654 1535 1660 1536
rect 1742 1540 1748 1541
rect 1742 1536 1743 1540
rect 1747 1536 1748 1540
rect 1742 1535 1748 1536
rect 1830 1540 1836 1541
rect 1830 1536 1831 1540
rect 1835 1536 1836 1540
rect 1830 1535 1836 1536
rect 1910 1540 1916 1541
rect 1910 1536 1911 1540
rect 1915 1536 1916 1540
rect 1910 1535 1916 1536
rect 1982 1540 1988 1541
rect 1982 1536 1983 1540
rect 1987 1536 1988 1540
rect 1982 1535 1988 1536
rect 2046 1540 2052 1541
rect 2046 1536 2047 1540
rect 2051 1536 2052 1540
rect 2046 1535 2052 1536
rect 2110 1540 2116 1541
rect 2110 1536 2111 1540
rect 2115 1536 2116 1540
rect 2110 1535 2116 1536
rect 2166 1540 2172 1541
rect 2166 1536 2167 1540
rect 2171 1536 2172 1540
rect 2166 1535 2172 1536
rect 2214 1540 2220 1541
rect 2214 1536 2215 1540
rect 2219 1536 2220 1540
rect 2214 1535 2220 1536
rect 1400 1531 1402 1535
rect 1480 1531 1482 1535
rect 1568 1531 1570 1535
rect 1656 1531 1658 1535
rect 1744 1531 1746 1535
rect 1832 1531 1834 1535
rect 1912 1531 1914 1535
rect 1984 1531 1986 1535
rect 2048 1531 2050 1535
rect 2112 1531 2114 1535
rect 2168 1531 2170 1535
rect 2216 1531 2218 1535
rect 1399 1530 1403 1531
rect 1399 1525 1403 1526
rect 1415 1530 1419 1531
rect 1415 1525 1419 1526
rect 1479 1530 1483 1531
rect 1479 1525 1483 1526
rect 1503 1530 1507 1531
rect 1503 1525 1507 1526
rect 1567 1530 1571 1531
rect 1567 1525 1571 1526
rect 1615 1530 1619 1531
rect 1615 1525 1619 1526
rect 1655 1530 1659 1531
rect 1655 1525 1659 1526
rect 1743 1530 1747 1531
rect 1743 1525 1747 1526
rect 1831 1530 1835 1531
rect 1831 1525 1835 1526
rect 1887 1530 1891 1531
rect 1887 1525 1891 1526
rect 1911 1530 1915 1531
rect 1911 1525 1915 1526
rect 1983 1530 1987 1531
rect 1983 1525 1987 1526
rect 2047 1530 2051 1531
rect 2047 1525 2051 1526
rect 2111 1530 2115 1531
rect 2111 1525 2115 1526
rect 2167 1530 2171 1531
rect 2167 1525 2171 1526
rect 2215 1530 2219 1531
rect 2215 1525 2219 1526
rect 1414 1524 1420 1525
rect 1414 1520 1415 1524
rect 1419 1520 1420 1524
rect 1414 1519 1420 1520
rect 1502 1524 1508 1525
rect 1502 1520 1503 1524
rect 1507 1520 1508 1524
rect 1502 1519 1508 1520
rect 1614 1524 1620 1525
rect 1614 1520 1615 1524
rect 1619 1520 1620 1524
rect 1614 1519 1620 1520
rect 1742 1524 1748 1525
rect 1742 1520 1743 1524
rect 1747 1520 1748 1524
rect 1742 1519 1748 1520
rect 1886 1524 1892 1525
rect 1886 1520 1887 1524
rect 1891 1520 1892 1524
rect 1886 1519 1892 1520
rect 2046 1524 2052 1525
rect 2046 1520 2047 1524
rect 2051 1520 2052 1524
rect 2046 1519 2052 1520
rect 2214 1524 2220 1525
rect 2214 1520 2215 1524
rect 2219 1520 2220 1524
rect 2214 1519 2220 1520
rect 1406 1503 1412 1504
rect 1406 1499 1407 1503
rect 1411 1499 1412 1503
rect 1406 1498 1412 1499
rect 1486 1503 1492 1504
rect 1486 1499 1487 1503
rect 1491 1499 1492 1503
rect 1486 1498 1492 1499
rect 1494 1503 1500 1504
rect 1494 1499 1495 1503
rect 1499 1499 1500 1503
rect 1494 1498 1500 1499
rect 1734 1503 1740 1504
rect 1734 1499 1735 1503
rect 1739 1499 1740 1503
rect 1734 1498 1740 1499
rect 2038 1503 2044 1504
rect 2038 1499 2039 1503
rect 2043 1499 2044 1503
rect 2038 1498 2044 1499
rect 1408 1468 1410 1498
rect 1414 1477 1420 1478
rect 1414 1473 1415 1477
rect 1419 1473 1420 1477
rect 1414 1472 1420 1473
rect 1342 1467 1348 1468
rect 1342 1463 1343 1467
rect 1347 1463 1348 1467
rect 1406 1467 1412 1468
rect 1406 1463 1407 1467
rect 1411 1463 1412 1467
rect 1416 1463 1418 1472
rect 1488 1468 1490 1498
rect 1486 1467 1492 1468
rect 1486 1463 1487 1467
rect 1491 1463 1492 1467
rect 1279 1462 1283 1463
rect 1279 1457 1283 1458
rect 1335 1462 1339 1463
rect 1342 1462 1348 1463
rect 1375 1462 1379 1463
rect 1406 1462 1412 1463
rect 1415 1462 1419 1463
rect 1335 1457 1339 1458
rect 1375 1457 1379 1458
rect 1415 1457 1419 1458
rect 1463 1462 1467 1463
rect 1486 1462 1492 1463
rect 1463 1457 1467 1458
rect 111 1454 115 1455
rect 111 1449 115 1450
rect 143 1454 147 1455
rect 143 1449 147 1450
rect 183 1454 187 1455
rect 183 1449 187 1450
rect 223 1454 227 1455
rect 223 1449 227 1450
rect 263 1454 267 1455
rect 263 1449 267 1450
rect 319 1454 323 1455
rect 319 1449 323 1450
rect 327 1454 331 1455
rect 327 1449 331 1450
rect 367 1454 371 1455
rect 367 1449 371 1450
rect 391 1454 395 1455
rect 391 1449 395 1450
rect 407 1454 411 1455
rect 407 1449 411 1450
rect 447 1454 451 1455
rect 447 1449 451 1450
rect 471 1454 475 1455
rect 471 1449 475 1450
rect 487 1454 491 1455
rect 487 1449 491 1450
rect 527 1454 531 1455
rect 527 1449 531 1450
rect 559 1454 563 1455
rect 559 1449 563 1450
rect 567 1454 571 1455
rect 567 1449 571 1450
rect 607 1454 611 1455
rect 607 1449 611 1450
rect 647 1454 651 1455
rect 647 1449 651 1450
rect 687 1454 691 1455
rect 687 1449 691 1450
rect 727 1454 731 1455
rect 727 1449 731 1450
rect 767 1454 771 1455
rect 767 1449 771 1450
rect 807 1454 811 1455
rect 807 1449 811 1450
rect 847 1454 851 1455
rect 847 1449 851 1450
rect 879 1454 883 1455
rect 879 1449 883 1450
rect 887 1454 891 1455
rect 887 1449 891 1450
rect 927 1454 931 1455
rect 927 1449 931 1450
rect 943 1454 947 1455
rect 943 1449 947 1450
rect 999 1454 1003 1455
rect 999 1449 1003 1450
rect 1047 1454 1051 1455
rect 1047 1449 1051 1450
rect 1103 1454 1107 1455
rect 1103 1449 1107 1450
rect 1151 1454 1155 1455
rect 1151 1449 1155 1450
rect 1191 1454 1195 1455
rect 1191 1449 1195 1450
rect 1239 1454 1243 1455
rect 1239 1449 1243 1450
rect 112 1417 114 1449
rect 144 1440 146 1449
rect 158 1447 164 1448
rect 158 1443 159 1447
rect 163 1443 164 1447
rect 158 1442 164 1443
rect 166 1447 172 1448
rect 166 1443 167 1447
rect 171 1443 172 1447
rect 166 1442 172 1443
rect 142 1439 148 1440
rect 142 1435 143 1439
rect 147 1435 148 1439
rect 142 1434 148 1435
rect 110 1416 116 1417
rect 110 1412 111 1416
rect 115 1412 116 1416
rect 110 1411 116 1412
rect 110 1399 116 1400
rect 110 1395 111 1399
rect 115 1395 116 1399
rect 110 1394 116 1395
rect 112 1387 114 1394
rect 142 1392 148 1393
rect 142 1388 143 1392
rect 147 1388 148 1392
rect 142 1387 148 1388
rect 111 1386 115 1387
rect 111 1381 115 1382
rect 143 1386 147 1387
rect 143 1381 147 1382
rect 112 1374 114 1381
rect 110 1373 116 1374
rect 110 1369 111 1373
rect 115 1369 116 1373
rect 110 1368 116 1369
rect 160 1368 162 1442
rect 168 1412 170 1442
rect 184 1440 186 1449
rect 206 1447 212 1448
rect 206 1443 207 1447
rect 211 1443 212 1447
rect 206 1442 212 1443
rect 182 1439 188 1440
rect 182 1435 183 1439
rect 187 1435 188 1439
rect 182 1434 188 1435
rect 208 1412 210 1442
rect 224 1440 226 1449
rect 250 1447 256 1448
rect 250 1443 251 1447
rect 255 1443 256 1447
rect 250 1442 256 1443
rect 222 1439 228 1440
rect 222 1435 223 1439
rect 227 1435 228 1439
rect 222 1434 228 1435
rect 252 1412 254 1442
rect 264 1440 266 1449
rect 320 1440 322 1449
rect 346 1447 352 1448
rect 346 1443 347 1447
rect 351 1443 352 1447
rect 346 1442 352 1443
rect 262 1439 268 1440
rect 262 1435 263 1439
rect 267 1435 268 1439
rect 262 1434 268 1435
rect 318 1439 324 1440
rect 318 1435 319 1439
rect 323 1435 324 1439
rect 318 1434 324 1435
rect 348 1412 350 1442
rect 392 1440 394 1449
rect 418 1447 424 1448
rect 418 1443 419 1447
rect 423 1443 424 1447
rect 418 1442 424 1443
rect 390 1439 396 1440
rect 390 1435 391 1439
rect 395 1435 396 1439
rect 390 1434 396 1435
rect 420 1412 422 1442
rect 472 1440 474 1449
rect 498 1447 504 1448
rect 498 1443 499 1447
rect 503 1443 504 1447
rect 498 1442 504 1443
rect 470 1439 476 1440
rect 470 1435 471 1439
rect 475 1435 476 1439
rect 470 1434 476 1435
rect 500 1412 502 1442
rect 560 1440 562 1449
rect 586 1447 592 1448
rect 586 1443 587 1447
rect 591 1443 592 1447
rect 586 1442 592 1443
rect 558 1439 564 1440
rect 558 1435 559 1439
rect 563 1435 564 1439
rect 558 1434 564 1435
rect 588 1412 590 1442
rect 648 1440 650 1449
rect 728 1440 730 1449
rect 742 1447 748 1448
rect 742 1443 743 1447
rect 747 1443 748 1447
rect 742 1442 748 1443
rect 754 1447 760 1448
rect 754 1443 755 1447
rect 759 1443 760 1447
rect 754 1442 760 1443
rect 646 1439 652 1440
rect 646 1435 647 1439
rect 651 1435 652 1439
rect 646 1434 652 1435
rect 726 1439 732 1440
rect 726 1435 727 1439
rect 731 1435 732 1439
rect 726 1434 732 1435
rect 166 1411 172 1412
rect 166 1407 167 1411
rect 171 1407 172 1411
rect 166 1406 172 1407
rect 206 1411 212 1412
rect 206 1407 207 1411
rect 211 1407 212 1411
rect 206 1406 212 1407
rect 250 1411 256 1412
rect 250 1407 251 1411
rect 255 1407 256 1411
rect 250 1406 256 1407
rect 346 1411 352 1412
rect 346 1407 347 1411
rect 351 1407 352 1411
rect 346 1406 352 1407
rect 418 1411 424 1412
rect 418 1407 419 1411
rect 423 1407 424 1411
rect 418 1406 424 1407
rect 498 1411 504 1412
rect 498 1407 499 1411
rect 503 1407 504 1411
rect 498 1406 504 1407
rect 586 1411 592 1412
rect 586 1407 587 1411
rect 591 1407 592 1411
rect 586 1406 592 1407
rect 374 1403 380 1404
rect 374 1399 375 1403
rect 379 1399 380 1403
rect 374 1398 380 1399
rect 182 1392 188 1393
rect 182 1388 183 1392
rect 187 1388 188 1392
rect 182 1387 188 1388
rect 222 1392 228 1393
rect 222 1388 223 1392
rect 227 1388 228 1392
rect 222 1387 228 1388
rect 262 1392 268 1393
rect 262 1388 263 1392
rect 267 1388 268 1392
rect 262 1387 268 1388
rect 318 1392 324 1393
rect 318 1388 319 1392
rect 323 1388 324 1392
rect 318 1387 324 1388
rect 167 1386 171 1387
rect 167 1381 171 1382
rect 183 1386 187 1387
rect 183 1381 187 1382
rect 207 1386 211 1387
rect 207 1381 211 1382
rect 223 1386 227 1387
rect 223 1381 227 1382
rect 247 1386 251 1387
rect 247 1381 251 1382
rect 263 1386 267 1387
rect 263 1381 267 1382
rect 303 1386 307 1387
rect 303 1381 307 1382
rect 319 1386 323 1387
rect 319 1381 323 1382
rect 367 1386 371 1387
rect 367 1381 371 1382
rect 166 1380 172 1381
rect 166 1376 167 1380
rect 171 1376 172 1380
rect 166 1375 172 1376
rect 206 1380 212 1381
rect 206 1376 207 1380
rect 211 1376 212 1380
rect 206 1375 212 1376
rect 246 1380 252 1381
rect 246 1376 247 1380
rect 251 1376 252 1380
rect 246 1375 252 1376
rect 302 1380 308 1381
rect 302 1376 303 1380
rect 307 1376 308 1380
rect 302 1375 308 1376
rect 366 1380 372 1381
rect 366 1376 367 1380
rect 371 1376 372 1380
rect 366 1375 372 1376
rect 158 1367 164 1368
rect 158 1363 159 1367
rect 163 1363 164 1367
rect 158 1362 164 1363
rect 194 1359 200 1360
rect 110 1356 116 1357
rect 110 1352 111 1356
rect 115 1352 116 1356
rect 194 1355 195 1359
rect 199 1355 200 1359
rect 194 1354 200 1355
rect 234 1359 240 1360
rect 234 1355 235 1359
rect 239 1355 240 1359
rect 234 1354 240 1355
rect 294 1359 300 1360
rect 294 1355 295 1359
rect 299 1355 300 1359
rect 294 1354 300 1355
rect 110 1351 116 1352
rect 112 1315 114 1351
rect 166 1333 172 1334
rect 166 1329 167 1333
rect 171 1329 172 1333
rect 166 1328 172 1329
rect 168 1315 170 1328
rect 196 1324 198 1354
rect 206 1333 212 1334
rect 206 1329 207 1333
rect 211 1329 212 1333
rect 206 1328 212 1329
rect 174 1323 180 1324
rect 174 1319 175 1323
rect 179 1319 180 1323
rect 174 1318 180 1319
rect 194 1323 200 1324
rect 194 1319 195 1323
rect 199 1319 200 1323
rect 194 1318 200 1319
rect 111 1314 115 1315
rect 111 1309 115 1310
rect 167 1314 171 1315
rect 167 1309 171 1310
rect 112 1277 114 1309
rect 110 1276 116 1277
rect 110 1272 111 1276
rect 115 1272 116 1276
rect 176 1272 178 1318
rect 208 1315 210 1328
rect 236 1324 238 1354
rect 246 1333 252 1334
rect 246 1329 247 1333
rect 251 1329 252 1333
rect 246 1328 252 1329
rect 234 1323 240 1324
rect 234 1319 235 1323
rect 239 1319 240 1323
rect 234 1318 240 1319
rect 248 1315 250 1328
rect 279 1324 283 1325
rect 296 1324 298 1354
rect 302 1333 308 1334
rect 302 1329 303 1333
rect 307 1329 308 1333
rect 302 1328 308 1329
rect 366 1333 372 1334
rect 366 1329 367 1333
rect 371 1329 372 1333
rect 366 1328 372 1329
rect 279 1319 283 1320
rect 294 1323 300 1324
rect 294 1319 295 1323
rect 299 1319 300 1323
rect 183 1314 187 1315
rect 183 1309 187 1310
rect 207 1314 211 1315
rect 207 1309 211 1310
rect 231 1314 235 1315
rect 231 1309 235 1310
rect 247 1314 251 1315
rect 247 1309 251 1310
rect 184 1300 186 1309
rect 218 1307 224 1308
rect 218 1303 219 1307
rect 223 1303 224 1307
rect 218 1302 224 1303
rect 182 1299 188 1300
rect 182 1295 183 1299
rect 187 1295 188 1299
rect 182 1294 188 1295
rect 220 1272 222 1302
rect 232 1300 234 1309
rect 280 1308 282 1319
rect 294 1318 300 1319
rect 304 1315 306 1328
rect 368 1315 370 1328
rect 376 1324 378 1398
rect 390 1392 396 1393
rect 390 1388 391 1392
rect 395 1388 396 1392
rect 390 1387 396 1388
rect 470 1392 476 1393
rect 470 1388 471 1392
rect 475 1388 476 1392
rect 470 1387 476 1388
rect 558 1392 564 1393
rect 558 1388 559 1392
rect 563 1388 564 1392
rect 558 1387 564 1388
rect 646 1392 652 1393
rect 646 1388 647 1392
rect 651 1388 652 1392
rect 646 1387 652 1388
rect 726 1392 732 1393
rect 726 1388 727 1392
rect 731 1388 732 1392
rect 726 1387 732 1388
rect 391 1386 395 1387
rect 391 1381 395 1382
rect 439 1386 443 1387
rect 439 1381 443 1382
rect 471 1386 475 1387
rect 471 1381 475 1382
rect 519 1386 523 1387
rect 519 1381 523 1382
rect 559 1386 563 1387
rect 559 1381 563 1382
rect 599 1386 603 1387
rect 599 1381 603 1382
rect 647 1386 651 1387
rect 647 1381 651 1382
rect 679 1386 683 1387
rect 679 1381 683 1382
rect 727 1386 731 1387
rect 727 1381 731 1382
rect 438 1380 444 1381
rect 438 1376 439 1380
rect 443 1376 444 1380
rect 438 1375 444 1376
rect 518 1380 524 1381
rect 518 1376 519 1380
rect 523 1376 524 1380
rect 518 1375 524 1376
rect 598 1380 604 1381
rect 598 1376 599 1380
rect 603 1376 604 1380
rect 598 1375 604 1376
rect 678 1380 684 1381
rect 678 1376 679 1380
rect 683 1376 684 1380
rect 678 1375 684 1376
rect 744 1368 746 1442
rect 756 1412 758 1442
rect 808 1440 810 1449
rect 834 1447 840 1448
rect 834 1443 835 1447
rect 839 1443 840 1447
rect 834 1442 840 1443
rect 806 1439 812 1440
rect 806 1435 807 1439
rect 811 1435 812 1439
rect 806 1434 812 1435
rect 836 1412 838 1442
rect 880 1440 882 1449
rect 906 1447 912 1448
rect 906 1443 907 1447
rect 911 1443 912 1447
rect 906 1442 912 1443
rect 878 1439 884 1440
rect 878 1435 879 1439
rect 883 1435 884 1439
rect 878 1434 884 1435
rect 908 1412 910 1442
rect 944 1440 946 1449
rect 970 1447 976 1448
rect 970 1443 971 1447
rect 975 1443 976 1447
rect 970 1442 976 1443
rect 942 1439 948 1440
rect 942 1435 943 1439
rect 947 1435 948 1439
rect 942 1434 948 1435
rect 972 1412 974 1442
rect 1000 1440 1002 1449
rect 1026 1447 1032 1448
rect 1026 1443 1027 1447
rect 1031 1443 1032 1447
rect 1026 1442 1032 1443
rect 998 1439 1004 1440
rect 998 1435 999 1439
rect 1003 1435 1004 1439
rect 998 1434 1004 1435
rect 1028 1412 1030 1442
rect 1048 1440 1050 1449
rect 1074 1447 1080 1448
rect 1074 1443 1075 1447
rect 1079 1443 1080 1447
rect 1074 1442 1080 1443
rect 1046 1439 1052 1440
rect 1046 1435 1047 1439
rect 1051 1435 1052 1439
rect 1046 1434 1052 1435
rect 1076 1412 1078 1442
rect 1104 1440 1106 1449
rect 1138 1447 1144 1448
rect 1138 1443 1139 1447
rect 1143 1443 1144 1447
rect 1138 1442 1144 1443
rect 1102 1439 1108 1440
rect 1102 1435 1103 1439
rect 1107 1435 1108 1439
rect 1102 1434 1108 1435
rect 1140 1412 1142 1442
rect 1152 1440 1154 1449
rect 1174 1447 1180 1448
rect 1174 1443 1175 1447
rect 1179 1443 1180 1447
rect 1174 1442 1180 1443
rect 1150 1439 1156 1440
rect 1150 1435 1151 1439
rect 1155 1435 1156 1439
rect 1150 1434 1156 1435
rect 1176 1412 1178 1442
rect 1192 1440 1194 1449
rect 1190 1439 1196 1440
rect 1190 1435 1191 1439
rect 1195 1435 1196 1439
rect 1190 1434 1196 1435
rect 1240 1417 1242 1449
rect 1280 1425 1282 1457
rect 1376 1448 1378 1457
rect 1450 1455 1456 1456
rect 1450 1451 1451 1455
rect 1455 1451 1456 1455
rect 1450 1450 1456 1451
rect 1374 1447 1380 1448
rect 1374 1443 1375 1447
rect 1379 1443 1380 1447
rect 1374 1442 1380 1443
rect 1278 1424 1284 1425
rect 1278 1420 1279 1424
rect 1283 1420 1284 1424
rect 1452 1420 1454 1450
rect 1464 1448 1466 1457
rect 1496 1456 1498 1498
rect 1502 1477 1508 1478
rect 1502 1473 1503 1477
rect 1507 1473 1508 1477
rect 1502 1472 1508 1473
rect 1614 1477 1620 1478
rect 1614 1473 1615 1477
rect 1619 1473 1620 1477
rect 1614 1472 1620 1473
rect 1504 1463 1506 1472
rect 1616 1463 1618 1472
rect 1736 1468 1738 1498
rect 1742 1477 1748 1478
rect 1742 1473 1743 1477
rect 1747 1473 1748 1477
rect 1742 1472 1748 1473
rect 1886 1477 1892 1478
rect 1886 1473 1887 1477
rect 1891 1473 1892 1477
rect 1886 1472 1892 1473
rect 1718 1467 1724 1468
rect 1718 1463 1719 1467
rect 1723 1463 1724 1467
rect 1734 1467 1740 1468
rect 1734 1463 1735 1467
rect 1739 1463 1740 1467
rect 1744 1463 1746 1472
rect 1888 1463 1890 1472
rect 2040 1468 2042 1498
rect 2046 1477 2052 1478
rect 2046 1473 2047 1477
rect 2051 1473 2052 1477
rect 2046 1472 2052 1473
rect 2214 1477 2220 1478
rect 2214 1473 2215 1477
rect 2219 1473 2220 1477
rect 2214 1472 2220 1473
rect 2038 1467 2044 1468
rect 2038 1463 2039 1467
rect 2043 1463 2044 1467
rect 2048 1463 2050 1472
rect 2216 1463 2218 1472
rect 2224 1468 2226 1546
rect 2406 1543 2407 1547
rect 2411 1543 2412 1547
rect 2406 1542 2412 1543
rect 2270 1540 2276 1541
rect 2270 1536 2271 1540
rect 2275 1536 2276 1540
rect 2270 1535 2276 1536
rect 2318 1540 2324 1541
rect 2318 1536 2319 1540
rect 2323 1536 2324 1540
rect 2318 1535 2324 1536
rect 2358 1540 2364 1541
rect 2358 1536 2359 1540
rect 2363 1536 2364 1540
rect 2358 1535 2364 1536
rect 2272 1531 2274 1535
rect 2320 1531 2322 1535
rect 2360 1531 2362 1535
rect 2408 1531 2410 1542
rect 2271 1530 2275 1531
rect 2271 1525 2275 1526
rect 2319 1530 2323 1531
rect 2319 1525 2323 1526
rect 2359 1530 2363 1531
rect 2359 1525 2363 1526
rect 2407 1530 2411 1531
rect 2407 1525 2411 1526
rect 2358 1524 2364 1525
rect 2358 1520 2359 1524
rect 2363 1520 2364 1524
rect 2358 1519 2364 1520
rect 2408 1518 2410 1525
rect 2406 1517 2412 1518
rect 2406 1513 2407 1517
rect 2411 1513 2412 1517
rect 2406 1512 2412 1513
rect 2350 1503 2356 1504
rect 2350 1499 2351 1503
rect 2355 1499 2356 1503
rect 2350 1498 2356 1499
rect 2366 1503 2372 1504
rect 2366 1499 2367 1503
rect 2371 1499 2372 1503
rect 2366 1498 2372 1499
rect 2406 1500 2412 1501
rect 2352 1468 2354 1498
rect 2358 1477 2364 1478
rect 2358 1473 2359 1477
rect 2363 1473 2364 1477
rect 2358 1472 2364 1473
rect 2222 1467 2228 1468
rect 2222 1463 2223 1467
rect 2227 1463 2228 1467
rect 2350 1467 2356 1468
rect 2350 1463 2351 1467
rect 2355 1463 2356 1467
rect 2360 1463 2362 1472
rect 1503 1462 1507 1463
rect 1503 1457 1507 1458
rect 1551 1462 1555 1463
rect 1551 1457 1555 1458
rect 1615 1462 1619 1463
rect 1615 1457 1619 1458
rect 1639 1462 1643 1463
rect 1718 1462 1724 1463
rect 1727 1462 1731 1463
rect 1734 1462 1740 1463
rect 1743 1462 1747 1463
rect 1639 1457 1643 1458
rect 1494 1455 1500 1456
rect 1494 1451 1495 1455
rect 1499 1451 1500 1455
rect 1494 1450 1500 1451
rect 1552 1448 1554 1457
rect 1558 1455 1564 1456
rect 1558 1451 1559 1455
rect 1563 1451 1564 1455
rect 1558 1450 1564 1451
rect 1578 1455 1584 1456
rect 1578 1451 1579 1455
rect 1583 1451 1584 1455
rect 1578 1450 1584 1451
rect 1462 1447 1468 1448
rect 1462 1443 1463 1447
rect 1467 1443 1468 1447
rect 1462 1442 1468 1443
rect 1550 1447 1556 1448
rect 1550 1443 1551 1447
rect 1555 1443 1556 1447
rect 1550 1442 1556 1443
rect 1278 1419 1284 1420
rect 1350 1419 1356 1420
rect 1238 1416 1244 1417
rect 1238 1412 1239 1416
rect 1243 1412 1244 1416
rect 1350 1415 1351 1419
rect 1355 1415 1356 1419
rect 1350 1414 1356 1415
rect 1450 1419 1456 1420
rect 1450 1415 1451 1419
rect 1455 1415 1456 1419
rect 1450 1414 1456 1415
rect 754 1411 760 1412
rect 754 1407 755 1411
rect 759 1407 760 1411
rect 754 1406 760 1407
rect 834 1411 840 1412
rect 834 1407 835 1411
rect 839 1407 840 1411
rect 834 1406 840 1407
rect 906 1411 912 1412
rect 906 1407 907 1411
rect 911 1407 912 1411
rect 906 1406 912 1407
rect 970 1411 976 1412
rect 970 1407 971 1411
rect 975 1407 976 1411
rect 970 1406 976 1407
rect 1026 1411 1032 1412
rect 1026 1407 1027 1411
rect 1031 1407 1032 1411
rect 1026 1406 1032 1407
rect 1074 1411 1080 1412
rect 1074 1407 1075 1411
rect 1079 1407 1080 1411
rect 1074 1406 1080 1407
rect 1138 1411 1144 1412
rect 1138 1407 1139 1411
rect 1143 1407 1144 1411
rect 1138 1406 1144 1407
rect 1174 1411 1180 1412
rect 1238 1411 1244 1412
rect 1174 1407 1175 1411
rect 1179 1407 1180 1411
rect 1174 1406 1180 1407
rect 1278 1407 1284 1408
rect 1086 1403 1092 1404
rect 1086 1399 1087 1403
rect 1091 1399 1092 1403
rect 1278 1403 1279 1407
rect 1283 1403 1284 1407
rect 1278 1402 1284 1403
rect 1086 1398 1092 1399
rect 1238 1399 1244 1400
rect 806 1392 812 1393
rect 806 1388 807 1392
rect 811 1388 812 1392
rect 806 1387 812 1388
rect 878 1392 884 1393
rect 878 1388 879 1392
rect 883 1388 884 1392
rect 878 1387 884 1388
rect 942 1392 948 1393
rect 942 1388 943 1392
rect 947 1388 948 1392
rect 942 1387 948 1388
rect 998 1392 1004 1393
rect 998 1388 999 1392
rect 1003 1388 1004 1392
rect 998 1387 1004 1388
rect 1046 1392 1052 1393
rect 1046 1388 1047 1392
rect 1051 1388 1052 1392
rect 1046 1387 1052 1388
rect 751 1386 755 1387
rect 751 1381 755 1382
rect 807 1386 811 1387
rect 807 1381 811 1382
rect 823 1386 827 1387
rect 823 1381 827 1382
rect 879 1386 883 1387
rect 879 1381 883 1382
rect 887 1386 891 1387
rect 887 1381 891 1382
rect 943 1386 947 1387
rect 943 1381 947 1382
rect 951 1386 955 1387
rect 951 1381 955 1382
rect 999 1386 1003 1387
rect 999 1381 1003 1382
rect 1015 1386 1019 1387
rect 1015 1381 1019 1382
rect 1047 1386 1051 1387
rect 1047 1381 1051 1382
rect 1079 1386 1083 1387
rect 1079 1381 1083 1382
rect 750 1380 756 1381
rect 750 1376 751 1380
rect 755 1376 756 1380
rect 750 1375 756 1376
rect 822 1380 828 1381
rect 822 1376 823 1380
rect 827 1376 828 1380
rect 822 1375 828 1376
rect 886 1380 892 1381
rect 886 1376 887 1380
rect 891 1376 892 1380
rect 886 1375 892 1376
rect 950 1380 956 1381
rect 950 1376 951 1380
rect 955 1376 956 1380
rect 950 1375 956 1376
rect 1014 1380 1020 1381
rect 1014 1376 1015 1380
rect 1019 1376 1020 1380
rect 1014 1375 1020 1376
rect 1078 1380 1084 1381
rect 1078 1376 1079 1380
rect 1083 1376 1084 1380
rect 1078 1375 1084 1376
rect 742 1367 748 1368
rect 742 1363 743 1367
rect 747 1363 748 1367
rect 742 1362 748 1363
rect 430 1359 436 1360
rect 430 1355 431 1359
rect 435 1355 436 1359
rect 430 1354 436 1355
rect 510 1359 516 1360
rect 510 1355 511 1359
rect 515 1355 516 1359
rect 510 1354 516 1355
rect 590 1359 596 1360
rect 590 1355 591 1359
rect 595 1355 596 1359
rect 590 1354 596 1355
rect 606 1359 612 1360
rect 606 1355 607 1359
rect 611 1355 612 1359
rect 606 1354 612 1355
rect 742 1359 748 1360
rect 742 1355 743 1359
rect 747 1355 748 1359
rect 742 1354 748 1355
rect 814 1359 820 1360
rect 814 1355 815 1359
rect 819 1355 820 1359
rect 814 1354 820 1355
rect 878 1359 884 1360
rect 878 1355 879 1359
rect 883 1355 884 1359
rect 878 1354 884 1355
rect 942 1359 948 1360
rect 942 1355 943 1359
rect 947 1355 948 1359
rect 942 1354 948 1355
rect 1006 1359 1012 1360
rect 1006 1355 1007 1359
rect 1011 1355 1012 1359
rect 1006 1354 1012 1355
rect 432 1324 434 1354
rect 438 1333 444 1334
rect 438 1329 439 1333
rect 443 1329 444 1333
rect 438 1328 444 1329
rect 374 1323 380 1324
rect 374 1319 375 1323
rect 379 1319 380 1323
rect 374 1318 380 1319
rect 430 1323 436 1324
rect 430 1319 431 1323
rect 435 1319 436 1323
rect 430 1318 436 1319
rect 440 1315 442 1328
rect 512 1324 514 1354
rect 518 1333 524 1334
rect 518 1329 519 1333
rect 523 1329 524 1333
rect 518 1328 524 1329
rect 510 1323 516 1324
rect 510 1319 511 1323
rect 515 1319 516 1323
rect 510 1318 516 1319
rect 520 1315 522 1328
rect 592 1324 594 1354
rect 598 1333 604 1334
rect 598 1329 599 1333
rect 603 1329 604 1333
rect 598 1328 604 1329
rect 590 1323 596 1324
rect 590 1319 591 1323
rect 595 1319 596 1323
rect 590 1318 596 1319
rect 600 1315 602 1328
rect 608 1325 610 1354
rect 678 1333 684 1334
rect 678 1329 679 1333
rect 683 1329 684 1333
rect 678 1328 684 1329
rect 607 1324 611 1325
rect 607 1319 611 1320
rect 680 1315 682 1328
rect 744 1324 746 1354
rect 750 1333 756 1334
rect 750 1329 751 1333
rect 755 1329 756 1333
rect 750 1328 756 1329
rect 742 1323 748 1324
rect 742 1319 743 1323
rect 747 1319 748 1323
rect 742 1318 748 1319
rect 752 1315 754 1328
rect 816 1324 818 1354
rect 822 1333 828 1334
rect 822 1329 823 1333
rect 827 1329 828 1333
rect 822 1328 828 1329
rect 814 1323 820 1324
rect 814 1319 815 1323
rect 819 1319 820 1323
rect 814 1318 820 1319
rect 824 1315 826 1328
rect 880 1324 882 1354
rect 886 1333 892 1334
rect 886 1329 887 1333
rect 891 1329 892 1333
rect 886 1328 892 1329
rect 878 1323 884 1324
rect 878 1319 879 1323
rect 883 1319 884 1323
rect 878 1318 884 1319
rect 888 1315 890 1328
rect 944 1324 946 1354
rect 950 1333 956 1334
rect 950 1329 951 1333
rect 955 1329 956 1333
rect 950 1328 956 1329
rect 942 1323 948 1324
rect 942 1319 943 1323
rect 947 1319 948 1323
rect 942 1318 948 1319
rect 952 1315 954 1328
rect 1008 1324 1010 1354
rect 1014 1333 1020 1334
rect 1014 1329 1015 1333
rect 1019 1329 1020 1333
rect 1014 1328 1020 1329
rect 1078 1333 1084 1334
rect 1078 1329 1079 1333
rect 1083 1329 1084 1333
rect 1078 1328 1084 1329
rect 1006 1323 1012 1324
rect 1006 1319 1007 1323
rect 1011 1319 1012 1323
rect 1006 1318 1012 1319
rect 1016 1315 1018 1328
rect 1022 1315 1028 1316
rect 1080 1315 1082 1328
rect 1088 1324 1090 1398
rect 1238 1395 1239 1399
rect 1243 1395 1244 1399
rect 1238 1394 1244 1395
rect 1102 1392 1108 1393
rect 1102 1388 1103 1392
rect 1107 1388 1108 1392
rect 1102 1387 1108 1388
rect 1150 1392 1156 1393
rect 1150 1388 1151 1392
rect 1155 1388 1156 1392
rect 1150 1387 1156 1388
rect 1190 1392 1196 1393
rect 1190 1388 1191 1392
rect 1195 1388 1196 1392
rect 1190 1387 1196 1388
rect 1240 1387 1242 1394
rect 1280 1387 1282 1402
rect 1103 1386 1107 1387
rect 1103 1381 1107 1382
rect 1143 1386 1147 1387
rect 1143 1381 1147 1382
rect 1151 1386 1155 1387
rect 1151 1381 1155 1382
rect 1191 1386 1195 1387
rect 1191 1381 1195 1382
rect 1239 1386 1243 1387
rect 1239 1381 1243 1382
rect 1279 1386 1283 1387
rect 1279 1381 1283 1382
rect 1303 1386 1307 1387
rect 1303 1381 1307 1382
rect 1343 1386 1347 1387
rect 1343 1381 1347 1382
rect 1142 1380 1148 1381
rect 1142 1376 1143 1380
rect 1147 1376 1148 1380
rect 1142 1375 1148 1376
rect 1190 1380 1196 1381
rect 1190 1376 1191 1380
rect 1195 1376 1196 1380
rect 1190 1375 1196 1376
rect 1240 1374 1242 1381
rect 1280 1374 1282 1381
rect 1302 1380 1308 1381
rect 1302 1376 1303 1380
rect 1307 1376 1308 1380
rect 1302 1375 1308 1376
rect 1342 1380 1348 1381
rect 1342 1376 1343 1380
rect 1347 1376 1348 1380
rect 1342 1375 1348 1376
rect 1238 1373 1244 1374
rect 1238 1369 1239 1373
rect 1243 1369 1244 1373
rect 1238 1368 1244 1369
rect 1278 1373 1284 1374
rect 1278 1369 1279 1373
rect 1283 1369 1284 1373
rect 1278 1368 1284 1369
rect 1134 1359 1140 1360
rect 1134 1355 1135 1359
rect 1139 1355 1140 1359
rect 1134 1354 1140 1355
rect 1182 1359 1188 1360
rect 1182 1355 1183 1359
rect 1187 1355 1188 1359
rect 1182 1354 1188 1355
rect 1230 1359 1236 1360
rect 1230 1355 1231 1359
rect 1235 1355 1236 1359
rect 1310 1359 1316 1360
rect 1230 1354 1236 1355
rect 1238 1356 1244 1357
rect 1136 1324 1138 1354
rect 1142 1333 1148 1334
rect 1142 1329 1143 1333
rect 1147 1329 1148 1333
rect 1142 1328 1148 1329
rect 1086 1323 1092 1324
rect 1086 1319 1087 1323
rect 1091 1319 1092 1323
rect 1086 1318 1092 1319
rect 1134 1323 1140 1324
rect 1134 1319 1135 1323
rect 1139 1319 1140 1323
rect 1134 1318 1140 1319
rect 1144 1315 1146 1328
rect 1184 1324 1186 1354
rect 1190 1333 1196 1334
rect 1190 1329 1191 1333
rect 1195 1329 1196 1333
rect 1190 1328 1196 1329
rect 1182 1323 1188 1324
rect 1182 1319 1183 1323
rect 1187 1319 1188 1323
rect 1182 1318 1188 1319
rect 1192 1315 1194 1328
rect 1232 1324 1234 1354
rect 1238 1352 1239 1356
rect 1243 1352 1244 1356
rect 1238 1351 1244 1352
rect 1278 1356 1284 1357
rect 1278 1352 1279 1356
rect 1283 1352 1284 1356
rect 1310 1355 1311 1359
rect 1315 1355 1316 1359
rect 1310 1354 1316 1355
rect 1278 1351 1284 1352
rect 1230 1323 1236 1324
rect 1230 1319 1231 1323
rect 1235 1319 1236 1323
rect 1230 1318 1236 1319
rect 1240 1315 1242 1351
rect 1280 1319 1282 1351
rect 1302 1333 1308 1334
rect 1302 1329 1303 1333
rect 1307 1329 1308 1333
rect 1302 1328 1308 1329
rect 1304 1319 1306 1328
rect 1279 1318 1283 1319
rect 287 1314 291 1315
rect 287 1309 291 1310
rect 303 1314 307 1315
rect 303 1309 307 1310
rect 351 1314 355 1315
rect 351 1309 355 1310
rect 367 1314 371 1315
rect 367 1309 371 1310
rect 423 1314 427 1315
rect 423 1309 427 1310
rect 439 1314 443 1315
rect 439 1309 443 1310
rect 495 1314 499 1315
rect 495 1309 499 1310
rect 519 1314 523 1315
rect 519 1309 523 1310
rect 567 1314 571 1315
rect 567 1309 571 1310
rect 599 1314 603 1315
rect 599 1309 603 1310
rect 639 1314 643 1315
rect 639 1309 643 1310
rect 679 1314 683 1315
rect 679 1309 683 1310
rect 703 1314 707 1315
rect 703 1309 707 1310
rect 751 1314 755 1315
rect 751 1309 755 1310
rect 767 1314 771 1315
rect 767 1309 771 1310
rect 823 1314 827 1315
rect 823 1309 827 1310
rect 879 1314 883 1315
rect 879 1309 883 1310
rect 887 1314 891 1315
rect 887 1309 891 1310
rect 935 1314 939 1315
rect 935 1309 939 1310
rect 951 1314 955 1315
rect 951 1309 955 1310
rect 999 1314 1003 1315
rect 999 1309 1003 1310
rect 1015 1314 1019 1315
rect 1022 1311 1023 1315
rect 1027 1311 1028 1315
rect 1022 1310 1028 1311
rect 1079 1314 1083 1315
rect 1015 1309 1019 1310
rect 254 1307 260 1308
rect 254 1303 255 1307
rect 259 1303 260 1307
rect 254 1302 260 1303
rect 278 1307 284 1308
rect 278 1303 279 1307
rect 283 1303 284 1307
rect 278 1302 284 1303
rect 230 1299 236 1300
rect 230 1295 231 1299
rect 235 1295 236 1299
rect 230 1294 236 1295
rect 110 1271 116 1272
rect 174 1271 180 1272
rect 174 1267 175 1271
rect 179 1267 180 1271
rect 174 1266 180 1267
rect 218 1271 224 1272
rect 218 1267 219 1271
rect 223 1267 224 1271
rect 218 1266 224 1267
rect 110 1259 116 1260
rect 110 1255 111 1259
rect 115 1255 116 1259
rect 110 1254 116 1255
rect 112 1243 114 1254
rect 182 1252 188 1253
rect 182 1248 183 1252
rect 187 1248 188 1252
rect 182 1247 188 1248
rect 230 1252 236 1253
rect 230 1248 231 1252
rect 235 1248 236 1252
rect 230 1247 236 1248
rect 184 1243 186 1247
rect 232 1243 234 1247
rect 111 1242 115 1243
rect 111 1237 115 1238
rect 135 1242 139 1243
rect 135 1237 139 1238
rect 175 1242 179 1243
rect 175 1237 179 1238
rect 183 1242 187 1243
rect 183 1237 187 1238
rect 231 1242 235 1243
rect 231 1237 235 1238
rect 112 1230 114 1237
rect 134 1236 140 1237
rect 134 1232 135 1236
rect 139 1232 140 1236
rect 134 1231 140 1232
rect 174 1236 180 1237
rect 174 1232 175 1236
rect 179 1232 180 1236
rect 174 1231 180 1232
rect 230 1236 236 1237
rect 230 1232 231 1236
rect 235 1232 236 1236
rect 230 1231 236 1232
rect 110 1229 116 1230
rect 110 1225 111 1229
rect 115 1225 116 1229
rect 110 1224 116 1225
rect 256 1216 258 1302
rect 288 1300 290 1309
rect 314 1307 320 1308
rect 314 1303 315 1307
rect 319 1303 320 1307
rect 314 1302 320 1303
rect 286 1299 292 1300
rect 286 1295 287 1299
rect 291 1295 292 1299
rect 286 1294 292 1295
rect 316 1272 318 1302
rect 352 1300 354 1309
rect 378 1307 384 1308
rect 378 1303 379 1307
rect 383 1303 384 1307
rect 378 1302 384 1303
rect 350 1299 356 1300
rect 350 1295 351 1299
rect 355 1295 356 1299
rect 350 1294 356 1295
rect 380 1272 382 1302
rect 424 1300 426 1309
rect 450 1307 456 1308
rect 450 1303 451 1307
rect 455 1303 456 1307
rect 450 1302 456 1303
rect 422 1299 428 1300
rect 422 1295 423 1299
rect 427 1295 428 1299
rect 422 1294 428 1295
rect 452 1272 454 1302
rect 496 1300 498 1309
rect 568 1300 570 1309
rect 640 1300 642 1309
rect 654 1307 660 1308
rect 654 1303 655 1307
rect 659 1303 660 1307
rect 654 1302 660 1303
rect 666 1307 672 1308
rect 666 1303 667 1307
rect 671 1303 672 1307
rect 666 1302 672 1303
rect 494 1299 500 1300
rect 494 1295 495 1299
rect 499 1295 500 1299
rect 494 1294 500 1295
rect 566 1299 572 1300
rect 566 1295 567 1299
rect 571 1295 572 1299
rect 566 1294 572 1295
rect 638 1299 644 1300
rect 638 1295 639 1299
rect 643 1295 644 1299
rect 638 1294 644 1295
rect 314 1271 320 1272
rect 314 1267 315 1271
rect 319 1267 320 1271
rect 314 1266 320 1267
rect 378 1271 384 1272
rect 378 1267 379 1271
rect 383 1267 384 1271
rect 378 1266 384 1267
rect 450 1271 456 1272
rect 450 1267 451 1271
rect 455 1267 456 1271
rect 450 1266 456 1267
rect 582 1271 588 1272
rect 582 1267 583 1271
rect 587 1267 588 1271
rect 582 1266 588 1267
rect 286 1252 292 1253
rect 286 1248 287 1252
rect 291 1248 292 1252
rect 286 1247 292 1248
rect 350 1252 356 1253
rect 350 1248 351 1252
rect 355 1248 356 1252
rect 350 1247 356 1248
rect 422 1252 428 1253
rect 422 1248 423 1252
rect 427 1248 428 1252
rect 422 1247 428 1248
rect 494 1252 500 1253
rect 494 1248 495 1252
rect 499 1248 500 1252
rect 494 1247 500 1248
rect 566 1252 572 1253
rect 566 1248 567 1252
rect 571 1248 572 1252
rect 566 1247 572 1248
rect 288 1243 290 1247
rect 352 1243 354 1247
rect 424 1243 426 1247
rect 496 1243 498 1247
rect 568 1243 570 1247
rect 287 1242 291 1243
rect 287 1237 291 1238
rect 311 1242 315 1243
rect 311 1237 315 1238
rect 351 1242 355 1243
rect 351 1237 355 1238
rect 399 1242 403 1243
rect 399 1237 403 1238
rect 423 1242 427 1243
rect 423 1237 427 1238
rect 487 1242 491 1243
rect 487 1237 491 1238
rect 495 1242 499 1243
rect 495 1237 499 1238
rect 567 1242 571 1243
rect 567 1237 571 1238
rect 575 1242 579 1243
rect 575 1237 579 1238
rect 310 1236 316 1237
rect 310 1232 311 1236
rect 315 1232 316 1236
rect 310 1231 316 1232
rect 398 1236 404 1237
rect 398 1232 399 1236
rect 403 1232 404 1236
rect 398 1231 404 1232
rect 486 1236 492 1237
rect 486 1232 487 1236
rect 491 1232 492 1236
rect 486 1231 492 1232
rect 574 1236 580 1237
rect 574 1232 575 1236
rect 579 1232 580 1236
rect 574 1231 580 1232
rect 162 1215 168 1216
rect 110 1212 116 1213
rect 110 1208 111 1212
rect 115 1208 116 1212
rect 162 1211 163 1215
rect 167 1211 168 1215
rect 162 1210 168 1211
rect 222 1215 228 1216
rect 222 1211 223 1215
rect 227 1211 228 1215
rect 222 1210 228 1211
rect 254 1215 260 1216
rect 254 1211 255 1215
rect 259 1211 260 1215
rect 254 1210 260 1211
rect 110 1207 116 1208
rect 112 1175 114 1207
rect 134 1189 140 1190
rect 134 1185 135 1189
rect 139 1185 140 1189
rect 134 1184 140 1185
rect 136 1175 138 1184
rect 164 1180 166 1210
rect 174 1189 180 1190
rect 174 1185 175 1189
rect 179 1185 180 1189
rect 174 1184 180 1185
rect 154 1179 160 1180
rect 154 1175 155 1179
rect 159 1175 160 1179
rect 111 1174 115 1175
rect 111 1169 115 1170
rect 135 1174 139 1175
rect 154 1174 160 1175
rect 162 1179 168 1180
rect 162 1175 163 1179
rect 167 1175 168 1179
rect 176 1175 178 1184
rect 224 1180 226 1210
rect 230 1189 236 1190
rect 230 1185 231 1189
rect 235 1185 236 1189
rect 230 1184 236 1185
rect 310 1189 316 1190
rect 310 1185 311 1189
rect 315 1185 316 1189
rect 310 1184 316 1185
rect 398 1189 404 1190
rect 398 1185 399 1189
rect 403 1185 404 1189
rect 398 1184 404 1185
rect 486 1189 492 1190
rect 486 1185 487 1189
rect 491 1185 492 1189
rect 486 1184 492 1185
rect 574 1189 580 1190
rect 574 1185 575 1189
rect 579 1185 580 1189
rect 574 1184 580 1185
rect 222 1179 228 1180
rect 222 1175 223 1179
rect 227 1175 228 1179
rect 232 1175 234 1184
rect 312 1175 314 1184
rect 400 1175 402 1184
rect 488 1175 490 1184
rect 576 1175 578 1184
rect 584 1180 586 1266
rect 638 1252 644 1253
rect 638 1248 639 1252
rect 643 1248 644 1252
rect 638 1247 644 1248
rect 640 1243 642 1247
rect 639 1242 643 1243
rect 639 1237 643 1238
rect 656 1216 658 1302
rect 668 1272 670 1302
rect 704 1300 706 1309
rect 730 1307 736 1308
rect 730 1303 731 1307
rect 735 1303 736 1307
rect 730 1302 736 1303
rect 702 1299 708 1300
rect 702 1295 703 1299
rect 707 1295 708 1299
rect 702 1294 708 1295
rect 732 1272 734 1302
rect 768 1300 770 1309
rect 794 1307 800 1308
rect 794 1303 795 1307
rect 799 1303 800 1307
rect 794 1302 800 1303
rect 766 1299 772 1300
rect 766 1295 767 1299
rect 771 1295 772 1299
rect 766 1294 772 1295
rect 796 1272 798 1302
rect 824 1300 826 1309
rect 850 1307 856 1308
rect 850 1303 851 1307
rect 855 1303 856 1307
rect 850 1302 856 1303
rect 822 1299 828 1300
rect 822 1295 823 1299
rect 827 1295 828 1299
rect 822 1294 828 1295
rect 852 1272 854 1302
rect 880 1300 882 1309
rect 906 1307 912 1308
rect 906 1303 907 1307
rect 911 1303 912 1307
rect 906 1302 912 1303
rect 878 1299 884 1300
rect 878 1295 879 1299
rect 883 1295 884 1299
rect 878 1294 884 1295
rect 908 1272 910 1302
rect 936 1300 938 1309
rect 962 1307 968 1308
rect 962 1303 963 1307
rect 967 1303 968 1307
rect 962 1302 968 1303
rect 934 1299 940 1300
rect 934 1295 935 1299
rect 939 1295 940 1299
rect 934 1294 940 1295
rect 964 1272 966 1302
rect 1000 1300 1002 1309
rect 998 1299 1004 1300
rect 998 1295 999 1299
rect 1003 1295 1004 1299
rect 998 1294 1004 1295
rect 1024 1272 1026 1310
rect 1079 1309 1083 1310
rect 1143 1314 1147 1315
rect 1143 1309 1147 1310
rect 1191 1314 1195 1315
rect 1191 1309 1195 1310
rect 1239 1314 1243 1315
rect 1279 1313 1283 1314
rect 1303 1318 1307 1319
rect 1303 1313 1307 1314
rect 1239 1309 1243 1310
rect 1240 1277 1242 1309
rect 1280 1281 1282 1313
rect 1304 1304 1306 1313
rect 1312 1312 1314 1354
rect 1342 1333 1348 1334
rect 1342 1329 1343 1333
rect 1347 1329 1348 1333
rect 1342 1328 1348 1329
rect 1344 1319 1346 1328
rect 1352 1324 1354 1414
rect 1374 1400 1380 1401
rect 1374 1396 1375 1400
rect 1379 1396 1380 1400
rect 1374 1395 1380 1396
rect 1462 1400 1468 1401
rect 1462 1396 1463 1400
rect 1467 1396 1468 1400
rect 1462 1395 1468 1396
rect 1550 1400 1556 1401
rect 1550 1396 1551 1400
rect 1555 1396 1556 1400
rect 1550 1395 1556 1396
rect 1376 1387 1378 1395
rect 1464 1387 1466 1395
rect 1552 1387 1554 1395
rect 1375 1386 1379 1387
rect 1375 1381 1379 1382
rect 1399 1386 1403 1387
rect 1399 1381 1403 1382
rect 1463 1386 1467 1387
rect 1463 1381 1467 1382
rect 1535 1386 1539 1387
rect 1535 1381 1539 1382
rect 1551 1386 1555 1387
rect 1551 1381 1555 1382
rect 1398 1380 1404 1381
rect 1398 1376 1399 1380
rect 1403 1376 1404 1380
rect 1398 1375 1404 1376
rect 1462 1380 1468 1381
rect 1462 1376 1463 1380
rect 1467 1376 1468 1380
rect 1462 1375 1468 1376
rect 1534 1380 1540 1381
rect 1534 1376 1535 1380
rect 1539 1376 1540 1380
rect 1534 1375 1540 1376
rect 1560 1360 1562 1450
rect 1580 1420 1582 1450
rect 1640 1448 1642 1457
rect 1666 1455 1672 1456
rect 1666 1451 1667 1455
rect 1671 1451 1672 1455
rect 1666 1450 1672 1451
rect 1638 1447 1644 1448
rect 1638 1443 1639 1447
rect 1643 1443 1644 1447
rect 1638 1442 1644 1443
rect 1668 1420 1670 1450
rect 1720 1420 1722 1462
rect 1727 1457 1731 1458
rect 1743 1457 1747 1458
rect 1807 1462 1811 1463
rect 1807 1457 1811 1458
rect 1879 1462 1883 1463
rect 1879 1457 1883 1458
rect 1887 1462 1891 1463
rect 1887 1457 1891 1458
rect 1943 1462 1947 1463
rect 1943 1457 1947 1458
rect 1999 1462 2003 1463
rect 2038 1462 2044 1463
rect 2047 1462 2051 1463
rect 1999 1457 2003 1458
rect 2047 1457 2051 1458
rect 2095 1462 2099 1463
rect 2095 1457 2099 1458
rect 2143 1462 2147 1463
rect 2143 1457 2147 1458
rect 2191 1462 2195 1463
rect 2191 1457 2195 1458
rect 2215 1462 2219 1463
rect 2222 1462 2228 1463
rect 2239 1462 2243 1463
rect 2215 1457 2219 1458
rect 2239 1457 2243 1458
rect 2279 1462 2283 1463
rect 2279 1457 2283 1458
rect 2319 1462 2323 1463
rect 2350 1462 2356 1463
rect 2359 1462 2363 1463
rect 2319 1457 2323 1458
rect 2359 1457 2363 1458
rect 1728 1448 1730 1457
rect 1808 1448 1810 1457
rect 1826 1455 1832 1456
rect 1826 1451 1827 1455
rect 1831 1451 1832 1455
rect 1826 1450 1832 1451
rect 1834 1455 1840 1456
rect 1834 1451 1835 1455
rect 1839 1451 1840 1455
rect 1834 1450 1840 1451
rect 1726 1447 1732 1448
rect 1726 1443 1727 1447
rect 1731 1443 1732 1447
rect 1726 1442 1732 1443
rect 1806 1447 1812 1448
rect 1806 1443 1807 1447
rect 1811 1443 1812 1447
rect 1806 1442 1812 1443
rect 1828 1428 1830 1450
rect 1826 1427 1832 1428
rect 1826 1423 1827 1427
rect 1831 1423 1832 1427
rect 1826 1422 1832 1423
rect 1836 1420 1838 1450
rect 1880 1448 1882 1457
rect 1906 1455 1912 1456
rect 1906 1451 1907 1455
rect 1911 1451 1912 1455
rect 1906 1450 1912 1451
rect 1878 1447 1884 1448
rect 1878 1443 1879 1447
rect 1883 1443 1884 1447
rect 1878 1442 1884 1443
rect 1908 1420 1910 1450
rect 1944 1448 1946 1457
rect 2000 1448 2002 1457
rect 2034 1455 2040 1456
rect 2034 1451 2035 1455
rect 2039 1451 2040 1455
rect 2034 1450 2040 1451
rect 1942 1447 1948 1448
rect 1942 1443 1943 1447
rect 1947 1443 1948 1447
rect 1942 1442 1948 1443
rect 1998 1447 2004 1448
rect 1998 1443 1999 1447
rect 2003 1443 2004 1447
rect 1998 1442 2004 1443
rect 2036 1420 2038 1450
rect 2048 1448 2050 1457
rect 2082 1455 2088 1456
rect 2082 1451 2083 1455
rect 2087 1451 2088 1455
rect 2082 1450 2088 1451
rect 2046 1447 2052 1448
rect 2046 1443 2047 1447
rect 2051 1443 2052 1447
rect 2046 1442 2052 1443
rect 2084 1420 2086 1450
rect 2096 1448 2098 1457
rect 2130 1455 2136 1456
rect 2130 1451 2131 1455
rect 2135 1451 2136 1455
rect 2130 1450 2136 1451
rect 2094 1447 2100 1448
rect 2094 1443 2095 1447
rect 2099 1443 2100 1447
rect 2094 1442 2100 1443
rect 2132 1420 2134 1450
rect 2144 1448 2146 1457
rect 2178 1455 2184 1456
rect 2178 1451 2179 1455
rect 2183 1451 2184 1455
rect 2178 1450 2184 1451
rect 2142 1447 2148 1448
rect 2142 1443 2143 1447
rect 2147 1443 2148 1447
rect 2142 1442 2148 1443
rect 2180 1420 2182 1450
rect 2192 1448 2194 1457
rect 2226 1455 2232 1456
rect 2226 1451 2227 1455
rect 2231 1451 2232 1455
rect 2226 1450 2232 1451
rect 2190 1447 2196 1448
rect 2190 1443 2191 1447
rect 2195 1443 2196 1447
rect 2190 1442 2196 1443
rect 2228 1420 2230 1450
rect 2240 1448 2242 1457
rect 2266 1455 2272 1456
rect 2266 1451 2267 1455
rect 2271 1451 2272 1455
rect 2266 1450 2272 1451
rect 2238 1447 2244 1448
rect 2238 1443 2239 1447
rect 2243 1443 2244 1447
rect 2238 1442 2244 1443
rect 2268 1428 2270 1450
rect 2280 1448 2282 1457
rect 2302 1455 2308 1456
rect 2302 1451 2303 1455
rect 2307 1451 2308 1455
rect 2302 1450 2308 1451
rect 2310 1455 2316 1456
rect 2310 1451 2311 1455
rect 2315 1451 2316 1455
rect 2310 1450 2316 1451
rect 2278 1447 2284 1448
rect 2278 1443 2279 1447
rect 2283 1443 2284 1447
rect 2278 1442 2284 1443
rect 2304 1428 2306 1450
rect 2266 1427 2272 1428
rect 2266 1423 2267 1427
rect 2271 1423 2272 1427
rect 2266 1422 2272 1423
rect 2302 1427 2308 1428
rect 2302 1423 2303 1427
rect 2307 1423 2308 1427
rect 2302 1422 2308 1423
rect 1578 1419 1584 1420
rect 1578 1415 1579 1419
rect 1583 1415 1584 1419
rect 1578 1414 1584 1415
rect 1666 1419 1672 1420
rect 1666 1415 1667 1419
rect 1671 1415 1672 1419
rect 1666 1414 1672 1415
rect 1718 1419 1724 1420
rect 1718 1415 1719 1419
rect 1723 1415 1724 1419
rect 1718 1414 1724 1415
rect 1834 1419 1840 1420
rect 1834 1415 1835 1419
rect 1839 1415 1840 1419
rect 1834 1414 1840 1415
rect 1906 1419 1912 1420
rect 1906 1415 1907 1419
rect 1911 1415 1912 1419
rect 1906 1414 1912 1415
rect 2034 1419 2040 1420
rect 2034 1415 2035 1419
rect 2039 1415 2040 1419
rect 2034 1414 2040 1415
rect 2082 1419 2088 1420
rect 2082 1415 2083 1419
rect 2087 1415 2088 1419
rect 2082 1414 2088 1415
rect 2130 1419 2136 1420
rect 2130 1415 2131 1419
rect 2135 1415 2136 1419
rect 2130 1414 2136 1415
rect 2178 1419 2184 1420
rect 2178 1415 2179 1419
rect 2183 1415 2184 1419
rect 2178 1414 2184 1415
rect 2226 1419 2232 1420
rect 2226 1415 2227 1419
rect 2231 1415 2232 1419
rect 2226 1414 2232 1415
rect 2014 1411 2020 1412
rect 2014 1407 2015 1411
rect 2019 1407 2020 1411
rect 2014 1406 2020 1407
rect 1638 1400 1644 1401
rect 1638 1396 1639 1400
rect 1643 1396 1644 1400
rect 1638 1395 1644 1396
rect 1726 1400 1732 1401
rect 1726 1396 1727 1400
rect 1731 1396 1732 1400
rect 1726 1395 1732 1396
rect 1806 1400 1812 1401
rect 1806 1396 1807 1400
rect 1811 1396 1812 1400
rect 1806 1395 1812 1396
rect 1878 1400 1884 1401
rect 1878 1396 1879 1400
rect 1883 1396 1884 1400
rect 1878 1395 1884 1396
rect 1942 1400 1948 1401
rect 1942 1396 1943 1400
rect 1947 1396 1948 1400
rect 1942 1395 1948 1396
rect 1998 1400 2004 1401
rect 1998 1396 1999 1400
rect 2003 1396 2004 1400
rect 1998 1395 2004 1396
rect 1640 1387 1642 1395
rect 1728 1387 1730 1395
rect 1808 1387 1810 1395
rect 1880 1387 1882 1395
rect 1944 1387 1946 1395
rect 2000 1387 2002 1395
rect 1607 1386 1611 1387
rect 1607 1381 1611 1382
rect 1639 1386 1643 1387
rect 1639 1381 1643 1382
rect 1687 1386 1691 1387
rect 1687 1381 1691 1382
rect 1727 1386 1731 1387
rect 1727 1381 1731 1382
rect 1767 1386 1771 1387
rect 1767 1381 1771 1382
rect 1807 1386 1811 1387
rect 1807 1381 1811 1382
rect 1847 1386 1851 1387
rect 1847 1381 1851 1382
rect 1879 1386 1883 1387
rect 1879 1381 1883 1382
rect 1935 1386 1939 1387
rect 1935 1381 1939 1382
rect 1943 1386 1947 1387
rect 1943 1381 1947 1382
rect 1999 1386 2003 1387
rect 1999 1381 2003 1382
rect 1606 1380 1612 1381
rect 1606 1376 1607 1380
rect 1611 1376 1612 1380
rect 1606 1375 1612 1376
rect 1686 1380 1692 1381
rect 1686 1376 1687 1380
rect 1691 1376 1692 1380
rect 1686 1375 1692 1376
rect 1766 1380 1772 1381
rect 1766 1376 1767 1380
rect 1771 1376 1772 1380
rect 1766 1375 1772 1376
rect 1846 1380 1852 1381
rect 1846 1376 1847 1380
rect 1851 1376 1852 1380
rect 1846 1375 1852 1376
rect 1934 1380 1940 1381
rect 1934 1376 1935 1380
rect 1939 1376 1940 1380
rect 1934 1375 1940 1376
rect 1390 1359 1396 1360
rect 1390 1355 1391 1359
rect 1395 1355 1396 1359
rect 1390 1354 1396 1355
rect 1454 1359 1460 1360
rect 1454 1355 1455 1359
rect 1459 1355 1460 1359
rect 1454 1354 1460 1355
rect 1490 1359 1496 1360
rect 1490 1355 1491 1359
rect 1495 1355 1496 1359
rect 1490 1354 1496 1355
rect 1558 1359 1564 1360
rect 1558 1355 1559 1359
rect 1563 1355 1564 1359
rect 1558 1354 1564 1355
rect 1782 1359 1788 1360
rect 1782 1355 1783 1359
rect 1787 1355 1788 1359
rect 1782 1354 1788 1355
rect 1392 1324 1394 1354
rect 1398 1333 1404 1334
rect 1398 1329 1399 1333
rect 1403 1329 1404 1333
rect 1398 1328 1404 1329
rect 1350 1323 1356 1324
rect 1350 1319 1351 1323
rect 1355 1319 1356 1323
rect 1390 1323 1396 1324
rect 1390 1319 1391 1323
rect 1395 1319 1396 1323
rect 1400 1319 1402 1328
rect 1456 1324 1458 1354
rect 1462 1333 1468 1334
rect 1462 1329 1463 1333
rect 1467 1329 1468 1333
rect 1462 1328 1468 1329
rect 1454 1323 1460 1324
rect 1454 1319 1455 1323
rect 1459 1319 1460 1323
rect 1464 1319 1466 1328
rect 1343 1318 1347 1319
rect 1350 1318 1356 1319
rect 1383 1318 1387 1319
rect 1390 1318 1396 1319
rect 1399 1318 1403 1319
rect 1343 1313 1347 1314
rect 1383 1313 1387 1314
rect 1399 1313 1403 1314
rect 1423 1318 1427 1319
rect 1454 1318 1460 1319
rect 1463 1318 1467 1319
rect 1423 1313 1427 1314
rect 1463 1313 1467 1314
rect 1310 1311 1316 1312
rect 1310 1307 1311 1311
rect 1315 1307 1316 1311
rect 1310 1306 1316 1307
rect 1330 1311 1336 1312
rect 1330 1307 1331 1311
rect 1335 1307 1336 1311
rect 1330 1306 1336 1307
rect 1302 1303 1308 1304
rect 1302 1299 1303 1303
rect 1307 1299 1308 1303
rect 1302 1298 1308 1299
rect 1278 1280 1284 1281
rect 1238 1276 1244 1277
rect 1238 1272 1239 1276
rect 1243 1272 1244 1276
rect 1278 1276 1279 1280
rect 1283 1276 1284 1280
rect 1332 1276 1334 1306
rect 1344 1304 1346 1313
rect 1370 1311 1376 1312
rect 1370 1307 1371 1311
rect 1375 1307 1376 1311
rect 1370 1306 1376 1307
rect 1342 1303 1348 1304
rect 1342 1299 1343 1303
rect 1347 1299 1348 1303
rect 1342 1298 1348 1299
rect 1372 1276 1374 1306
rect 1384 1304 1386 1313
rect 1410 1311 1416 1312
rect 1410 1307 1411 1311
rect 1415 1307 1416 1311
rect 1410 1306 1416 1307
rect 1382 1303 1388 1304
rect 1382 1299 1383 1303
rect 1387 1299 1388 1303
rect 1382 1298 1388 1299
rect 1412 1276 1414 1306
rect 1424 1304 1426 1313
rect 1446 1311 1452 1312
rect 1446 1307 1447 1311
rect 1451 1307 1452 1311
rect 1446 1306 1452 1307
rect 1422 1303 1428 1304
rect 1422 1299 1423 1303
rect 1427 1299 1428 1303
rect 1422 1298 1428 1299
rect 1448 1276 1450 1306
rect 1464 1304 1466 1313
rect 1492 1312 1494 1354
rect 1534 1333 1540 1334
rect 1534 1329 1535 1333
rect 1539 1329 1540 1333
rect 1534 1328 1540 1329
rect 1606 1333 1612 1334
rect 1606 1329 1607 1333
rect 1611 1329 1612 1333
rect 1606 1328 1612 1329
rect 1686 1333 1692 1334
rect 1686 1329 1687 1333
rect 1691 1329 1692 1333
rect 1686 1328 1692 1329
rect 1766 1333 1772 1334
rect 1766 1329 1767 1333
rect 1771 1329 1772 1333
rect 1766 1328 1772 1329
rect 1536 1319 1538 1328
rect 1608 1319 1610 1328
rect 1688 1319 1690 1328
rect 1754 1323 1760 1324
rect 1754 1319 1755 1323
rect 1759 1319 1760 1323
rect 1768 1319 1770 1328
rect 1503 1318 1507 1319
rect 1503 1313 1507 1314
rect 1535 1318 1539 1319
rect 1535 1313 1539 1314
rect 1543 1318 1547 1319
rect 1543 1313 1547 1314
rect 1583 1318 1587 1319
rect 1583 1313 1587 1314
rect 1607 1318 1611 1319
rect 1607 1313 1611 1314
rect 1623 1318 1627 1319
rect 1623 1313 1627 1314
rect 1679 1318 1683 1319
rect 1679 1313 1683 1314
rect 1687 1318 1691 1319
rect 1687 1313 1691 1314
rect 1735 1318 1739 1319
rect 1754 1318 1760 1319
rect 1767 1318 1771 1319
rect 1735 1313 1739 1314
rect 1490 1311 1496 1312
rect 1490 1307 1491 1311
rect 1495 1307 1496 1311
rect 1490 1306 1496 1307
rect 1504 1304 1506 1313
rect 1526 1311 1532 1312
rect 1526 1307 1527 1311
rect 1531 1307 1532 1311
rect 1526 1306 1532 1307
rect 1462 1303 1468 1304
rect 1462 1299 1463 1303
rect 1467 1299 1468 1303
rect 1462 1298 1468 1299
rect 1502 1303 1508 1304
rect 1502 1299 1503 1303
rect 1507 1299 1508 1303
rect 1502 1298 1508 1299
rect 1528 1276 1530 1306
rect 1544 1304 1546 1313
rect 1550 1311 1556 1312
rect 1550 1307 1551 1311
rect 1555 1307 1556 1311
rect 1550 1306 1556 1307
rect 1542 1303 1548 1304
rect 1542 1299 1543 1303
rect 1547 1299 1548 1303
rect 1542 1298 1548 1299
rect 1552 1284 1554 1306
rect 1584 1304 1586 1313
rect 1614 1311 1620 1312
rect 1614 1307 1615 1311
rect 1619 1307 1620 1311
rect 1614 1306 1620 1307
rect 1582 1303 1588 1304
rect 1582 1299 1583 1303
rect 1587 1299 1588 1303
rect 1582 1298 1588 1299
rect 1550 1283 1556 1284
rect 1550 1279 1551 1283
rect 1555 1279 1556 1283
rect 1550 1278 1556 1279
rect 1616 1276 1618 1306
rect 1624 1304 1626 1313
rect 1650 1311 1656 1312
rect 1650 1307 1651 1311
rect 1655 1307 1656 1311
rect 1650 1306 1656 1307
rect 1622 1303 1628 1304
rect 1622 1299 1623 1303
rect 1627 1299 1628 1303
rect 1622 1298 1628 1299
rect 1652 1276 1654 1306
rect 1680 1304 1682 1313
rect 1736 1304 1738 1313
rect 1678 1303 1684 1304
rect 1678 1299 1679 1303
rect 1683 1299 1684 1303
rect 1678 1298 1684 1299
rect 1734 1303 1740 1304
rect 1734 1299 1735 1303
rect 1739 1299 1740 1303
rect 1734 1298 1740 1299
rect 1756 1276 1758 1318
rect 1767 1313 1771 1314
rect 1784 1312 1786 1354
rect 1942 1351 1948 1352
rect 1942 1347 1943 1351
rect 1947 1347 1948 1351
rect 1942 1346 1948 1347
rect 1846 1333 1852 1334
rect 1846 1329 1847 1333
rect 1851 1329 1852 1333
rect 1846 1328 1852 1329
rect 1934 1333 1940 1334
rect 1934 1329 1935 1333
rect 1939 1329 1940 1333
rect 1934 1328 1940 1329
rect 1848 1319 1850 1328
rect 1936 1319 1938 1328
rect 1944 1324 1946 1346
rect 2016 1324 2018 1406
rect 2046 1400 2052 1401
rect 2046 1396 2047 1400
rect 2051 1396 2052 1400
rect 2046 1395 2052 1396
rect 2094 1400 2100 1401
rect 2094 1396 2095 1400
rect 2099 1396 2100 1400
rect 2094 1395 2100 1396
rect 2142 1400 2148 1401
rect 2142 1396 2143 1400
rect 2147 1396 2148 1400
rect 2142 1395 2148 1396
rect 2190 1400 2196 1401
rect 2190 1396 2191 1400
rect 2195 1396 2196 1400
rect 2190 1395 2196 1396
rect 2238 1400 2244 1401
rect 2238 1396 2239 1400
rect 2243 1396 2244 1400
rect 2238 1395 2244 1396
rect 2278 1400 2284 1401
rect 2278 1396 2279 1400
rect 2283 1396 2284 1400
rect 2278 1395 2284 1396
rect 2048 1387 2050 1395
rect 2096 1387 2098 1395
rect 2144 1387 2146 1395
rect 2192 1387 2194 1395
rect 2240 1387 2242 1395
rect 2280 1387 2282 1395
rect 2023 1386 2027 1387
rect 2023 1381 2027 1382
rect 2047 1386 2051 1387
rect 2047 1381 2051 1382
rect 2095 1386 2099 1387
rect 2095 1381 2099 1382
rect 2111 1386 2115 1387
rect 2111 1381 2115 1382
rect 2143 1386 2147 1387
rect 2143 1381 2147 1382
rect 2191 1386 2195 1387
rect 2191 1381 2195 1382
rect 2199 1386 2203 1387
rect 2199 1381 2203 1382
rect 2239 1386 2243 1387
rect 2239 1381 2243 1382
rect 2279 1386 2283 1387
rect 2279 1381 2283 1382
rect 2287 1386 2291 1387
rect 2287 1381 2291 1382
rect 2022 1380 2028 1381
rect 2022 1376 2023 1380
rect 2027 1376 2028 1380
rect 2022 1375 2028 1376
rect 2110 1380 2116 1381
rect 2110 1376 2111 1380
rect 2115 1376 2116 1380
rect 2110 1375 2116 1376
rect 2198 1380 2204 1381
rect 2198 1376 2199 1380
rect 2203 1376 2204 1380
rect 2198 1375 2204 1376
rect 2286 1380 2292 1381
rect 2286 1376 2287 1380
rect 2291 1376 2292 1380
rect 2286 1375 2292 1376
rect 2312 1360 2314 1450
rect 2320 1448 2322 1457
rect 2360 1448 2362 1457
rect 2368 1456 2370 1498
rect 2406 1496 2407 1500
rect 2411 1496 2412 1500
rect 2406 1495 2412 1496
rect 2408 1463 2410 1495
rect 2407 1462 2411 1463
rect 2407 1457 2411 1458
rect 2366 1455 2372 1456
rect 2366 1451 2367 1455
rect 2371 1451 2372 1455
rect 2366 1450 2372 1451
rect 2318 1447 2324 1448
rect 2318 1443 2319 1447
rect 2323 1443 2324 1447
rect 2318 1442 2324 1443
rect 2358 1447 2364 1448
rect 2358 1443 2359 1447
rect 2363 1443 2364 1447
rect 2358 1442 2364 1443
rect 2408 1425 2410 1457
rect 2406 1424 2412 1425
rect 2406 1420 2407 1424
rect 2411 1420 2412 1424
rect 2374 1419 2380 1420
rect 2406 1419 2412 1420
rect 2374 1415 2375 1419
rect 2379 1415 2380 1419
rect 2374 1414 2380 1415
rect 2318 1400 2324 1401
rect 2318 1396 2319 1400
rect 2323 1396 2324 1400
rect 2318 1395 2324 1396
rect 2358 1400 2364 1401
rect 2358 1396 2359 1400
rect 2363 1396 2364 1400
rect 2358 1395 2364 1396
rect 2320 1387 2322 1395
rect 2360 1387 2362 1395
rect 2319 1386 2323 1387
rect 2319 1381 2323 1382
rect 2359 1386 2363 1387
rect 2359 1381 2363 1382
rect 2358 1380 2364 1381
rect 2358 1376 2359 1380
rect 2363 1376 2364 1380
rect 2358 1375 2364 1376
rect 2102 1359 2108 1360
rect 2102 1355 2103 1359
rect 2107 1355 2108 1359
rect 2102 1354 2108 1355
rect 2270 1359 2276 1360
rect 2270 1355 2271 1359
rect 2275 1355 2276 1359
rect 2270 1354 2276 1355
rect 2310 1359 2316 1360
rect 2310 1355 2311 1359
rect 2315 1355 2316 1359
rect 2310 1354 2316 1355
rect 2366 1359 2372 1360
rect 2366 1355 2367 1359
rect 2371 1355 2372 1359
rect 2366 1354 2372 1355
rect 2022 1333 2028 1334
rect 2022 1329 2023 1333
rect 2027 1329 2028 1333
rect 2022 1328 2028 1329
rect 1942 1323 1948 1324
rect 1942 1319 1943 1323
rect 1947 1319 1948 1323
rect 2014 1323 2020 1324
rect 2014 1319 2015 1323
rect 2019 1319 2020 1323
rect 2024 1319 2026 1328
rect 2104 1324 2106 1354
rect 2110 1333 2116 1334
rect 2110 1329 2111 1333
rect 2115 1329 2116 1333
rect 2110 1328 2116 1329
rect 2198 1333 2204 1334
rect 2198 1329 2199 1333
rect 2203 1329 2204 1333
rect 2198 1328 2204 1329
rect 2102 1323 2108 1324
rect 2102 1319 2103 1323
rect 2107 1319 2108 1323
rect 2112 1319 2114 1328
rect 2200 1319 2202 1328
rect 2272 1324 2274 1354
rect 2286 1333 2292 1334
rect 2286 1329 2287 1333
rect 2291 1329 2292 1333
rect 2286 1328 2292 1329
rect 2358 1333 2364 1334
rect 2358 1329 2359 1333
rect 2363 1329 2364 1333
rect 2358 1328 2364 1329
rect 2262 1323 2268 1324
rect 2262 1319 2263 1323
rect 2267 1319 2268 1323
rect 1791 1318 1795 1319
rect 1791 1313 1795 1314
rect 1847 1318 1851 1319
rect 1847 1313 1851 1314
rect 1903 1318 1907 1319
rect 1903 1313 1907 1314
rect 1935 1318 1939 1319
rect 1942 1318 1948 1319
rect 1967 1318 1971 1319
rect 2014 1318 2020 1319
rect 2023 1318 2027 1319
rect 1935 1313 1939 1314
rect 1967 1313 1971 1314
rect 2023 1313 2027 1314
rect 2039 1318 2043 1319
rect 2102 1318 2108 1319
rect 2111 1318 2115 1319
rect 2039 1313 2043 1314
rect 2111 1313 2115 1314
rect 2119 1318 2123 1319
rect 2119 1313 2123 1314
rect 2199 1318 2203 1319
rect 2262 1318 2268 1319
rect 2270 1323 2276 1324
rect 2270 1319 2271 1323
rect 2275 1319 2276 1323
rect 2288 1319 2290 1328
rect 2360 1319 2362 1328
rect 2270 1318 2276 1319
rect 2287 1318 2291 1319
rect 2199 1313 2203 1314
rect 1782 1311 1788 1312
rect 1782 1307 1783 1311
rect 1787 1307 1788 1311
rect 1782 1306 1788 1307
rect 1792 1304 1794 1313
rect 1818 1311 1824 1312
rect 1818 1307 1819 1311
rect 1823 1307 1824 1311
rect 1818 1306 1824 1307
rect 1790 1303 1796 1304
rect 1790 1299 1791 1303
rect 1795 1299 1796 1303
rect 1790 1298 1796 1299
rect 1820 1276 1822 1306
rect 1848 1304 1850 1313
rect 1874 1311 1880 1312
rect 1874 1307 1875 1311
rect 1879 1307 1880 1311
rect 1874 1306 1880 1307
rect 1846 1303 1852 1304
rect 1846 1299 1847 1303
rect 1851 1299 1852 1303
rect 1846 1298 1852 1299
rect 1876 1276 1878 1306
rect 1904 1304 1906 1313
rect 1968 1304 1970 1313
rect 1994 1311 2000 1312
rect 1994 1307 1995 1311
rect 1999 1307 2000 1311
rect 1994 1306 2000 1307
rect 1902 1303 1908 1304
rect 1902 1299 1903 1303
rect 1907 1299 1908 1303
rect 1902 1298 1908 1299
rect 1966 1303 1972 1304
rect 1966 1299 1967 1303
rect 1971 1299 1972 1303
rect 1966 1298 1972 1299
rect 1996 1276 1998 1306
rect 2040 1304 2042 1313
rect 2066 1311 2072 1312
rect 2066 1307 2067 1311
rect 2071 1307 2072 1311
rect 2066 1306 2072 1307
rect 2038 1303 2044 1304
rect 2038 1299 2039 1303
rect 2043 1299 2044 1303
rect 2038 1298 2044 1299
rect 2068 1276 2070 1306
rect 2120 1304 2122 1313
rect 2146 1311 2152 1312
rect 2146 1307 2147 1311
rect 2151 1307 2152 1311
rect 2146 1306 2152 1307
rect 2118 1303 2124 1304
rect 2118 1299 2119 1303
rect 2123 1299 2124 1303
rect 2118 1298 2124 1299
rect 2148 1276 2150 1306
rect 2200 1304 2202 1313
rect 2250 1311 2256 1312
rect 2250 1307 2251 1311
rect 2255 1307 2256 1311
rect 2250 1306 2256 1307
rect 2198 1303 2204 1304
rect 2198 1299 2199 1303
rect 2203 1299 2204 1303
rect 2198 1298 2204 1299
rect 1278 1275 1284 1276
rect 1330 1275 1336 1276
rect 666 1271 672 1272
rect 666 1267 667 1271
rect 671 1267 672 1271
rect 666 1266 672 1267
rect 730 1271 736 1272
rect 730 1267 731 1271
rect 735 1267 736 1271
rect 730 1266 736 1267
rect 794 1271 800 1272
rect 794 1267 795 1271
rect 799 1267 800 1271
rect 794 1266 800 1267
rect 850 1271 856 1272
rect 850 1267 851 1271
rect 855 1267 856 1271
rect 850 1266 856 1267
rect 906 1271 912 1272
rect 906 1267 907 1271
rect 911 1267 912 1271
rect 906 1266 912 1267
rect 962 1271 968 1272
rect 962 1267 963 1271
rect 967 1267 968 1271
rect 962 1266 968 1267
rect 1022 1271 1028 1272
rect 1238 1271 1244 1272
rect 1330 1271 1331 1275
rect 1335 1271 1336 1275
rect 1022 1267 1023 1271
rect 1027 1267 1028 1271
rect 1330 1270 1336 1271
rect 1370 1275 1376 1276
rect 1370 1271 1371 1275
rect 1375 1271 1376 1275
rect 1370 1270 1376 1271
rect 1410 1275 1416 1276
rect 1410 1271 1411 1275
rect 1415 1271 1416 1275
rect 1410 1270 1416 1271
rect 1446 1275 1452 1276
rect 1446 1271 1447 1275
rect 1451 1271 1452 1275
rect 1446 1270 1452 1271
rect 1526 1275 1532 1276
rect 1526 1271 1527 1275
rect 1531 1271 1532 1275
rect 1526 1270 1532 1271
rect 1570 1275 1576 1276
rect 1570 1271 1571 1275
rect 1575 1271 1576 1275
rect 1570 1270 1576 1271
rect 1610 1275 1618 1276
rect 1610 1271 1611 1275
rect 1615 1272 1618 1275
rect 1650 1275 1656 1276
rect 1615 1271 1616 1272
rect 1610 1270 1616 1271
rect 1650 1271 1651 1275
rect 1655 1271 1656 1275
rect 1650 1270 1656 1271
rect 1754 1275 1760 1276
rect 1754 1271 1755 1275
rect 1759 1271 1760 1275
rect 1754 1270 1760 1271
rect 1818 1275 1824 1276
rect 1818 1271 1819 1275
rect 1823 1271 1824 1275
rect 1818 1270 1824 1271
rect 1874 1275 1880 1276
rect 1874 1271 1875 1275
rect 1879 1271 1880 1275
rect 1874 1270 1880 1271
rect 1994 1275 2000 1276
rect 1994 1271 1995 1275
rect 1999 1271 2000 1275
rect 1994 1270 2000 1271
rect 2066 1275 2072 1276
rect 2066 1271 2067 1275
rect 2071 1271 2072 1275
rect 2066 1270 2072 1271
rect 2146 1275 2152 1276
rect 2146 1271 2147 1275
rect 2151 1271 2152 1275
rect 2146 1270 2152 1271
rect 1022 1266 1028 1267
rect 1278 1263 1284 1264
rect 1238 1259 1244 1260
rect 1238 1255 1239 1259
rect 1243 1255 1244 1259
rect 1278 1259 1279 1263
rect 1283 1259 1284 1263
rect 1278 1258 1284 1259
rect 1238 1254 1244 1255
rect 702 1252 708 1253
rect 702 1248 703 1252
rect 707 1248 708 1252
rect 702 1247 708 1248
rect 766 1252 772 1253
rect 766 1248 767 1252
rect 771 1248 772 1252
rect 766 1247 772 1248
rect 822 1252 828 1253
rect 822 1248 823 1252
rect 827 1248 828 1252
rect 822 1247 828 1248
rect 878 1252 884 1253
rect 878 1248 879 1252
rect 883 1248 884 1252
rect 878 1247 884 1248
rect 934 1252 940 1253
rect 934 1248 935 1252
rect 939 1248 940 1252
rect 934 1247 940 1248
rect 998 1252 1004 1253
rect 998 1248 999 1252
rect 1003 1248 1004 1252
rect 998 1247 1004 1248
rect 704 1243 706 1247
rect 768 1243 770 1247
rect 824 1243 826 1247
rect 880 1243 882 1247
rect 936 1243 938 1247
rect 1000 1243 1002 1247
rect 1240 1243 1242 1254
rect 1280 1243 1282 1258
rect 1302 1256 1308 1257
rect 1302 1252 1303 1256
rect 1307 1252 1308 1256
rect 1302 1251 1308 1252
rect 1342 1256 1348 1257
rect 1342 1252 1343 1256
rect 1347 1252 1348 1256
rect 1342 1251 1348 1252
rect 1382 1256 1388 1257
rect 1382 1252 1383 1256
rect 1387 1252 1388 1256
rect 1382 1251 1388 1252
rect 1422 1256 1428 1257
rect 1422 1252 1423 1256
rect 1427 1252 1428 1256
rect 1422 1251 1428 1252
rect 1462 1256 1468 1257
rect 1462 1252 1463 1256
rect 1467 1252 1468 1256
rect 1462 1251 1468 1252
rect 1502 1256 1508 1257
rect 1502 1252 1503 1256
rect 1507 1252 1508 1256
rect 1502 1251 1508 1252
rect 1542 1256 1548 1257
rect 1542 1252 1543 1256
rect 1547 1252 1548 1256
rect 1542 1251 1548 1252
rect 1304 1243 1306 1251
rect 1344 1243 1346 1251
rect 1384 1243 1386 1251
rect 1424 1243 1426 1251
rect 1464 1243 1466 1251
rect 1504 1243 1506 1251
rect 1544 1243 1546 1251
rect 663 1242 667 1243
rect 663 1237 667 1238
rect 703 1242 707 1243
rect 703 1237 707 1238
rect 743 1242 747 1243
rect 743 1237 747 1238
rect 767 1242 771 1243
rect 767 1237 771 1238
rect 815 1242 819 1243
rect 815 1237 819 1238
rect 823 1242 827 1243
rect 823 1237 827 1238
rect 879 1242 883 1243
rect 879 1237 883 1238
rect 935 1242 939 1243
rect 935 1237 939 1238
rect 943 1242 947 1243
rect 943 1237 947 1238
rect 999 1242 1003 1243
rect 999 1237 1003 1238
rect 1007 1242 1011 1243
rect 1007 1237 1011 1238
rect 1071 1242 1075 1243
rect 1071 1237 1075 1238
rect 1239 1242 1243 1243
rect 1239 1237 1243 1238
rect 1279 1242 1283 1243
rect 1279 1237 1283 1238
rect 1303 1242 1307 1243
rect 1303 1237 1307 1238
rect 1343 1242 1347 1243
rect 1343 1237 1347 1238
rect 1375 1242 1379 1243
rect 1375 1237 1379 1238
rect 1383 1242 1387 1243
rect 1383 1237 1387 1238
rect 1423 1242 1427 1243
rect 1423 1237 1427 1238
rect 1463 1242 1467 1243
rect 1463 1237 1467 1238
rect 1479 1242 1483 1243
rect 1479 1237 1483 1238
rect 1503 1242 1507 1243
rect 1503 1237 1507 1238
rect 1543 1242 1547 1243
rect 1543 1237 1547 1238
rect 662 1236 668 1237
rect 662 1232 663 1236
rect 667 1232 668 1236
rect 662 1231 668 1232
rect 742 1236 748 1237
rect 742 1232 743 1236
rect 747 1232 748 1236
rect 742 1231 748 1232
rect 814 1236 820 1237
rect 814 1232 815 1236
rect 819 1232 820 1236
rect 814 1231 820 1232
rect 878 1236 884 1237
rect 878 1232 879 1236
rect 883 1232 884 1236
rect 878 1231 884 1232
rect 942 1236 948 1237
rect 942 1232 943 1236
rect 947 1232 948 1236
rect 942 1231 948 1232
rect 1006 1236 1012 1237
rect 1006 1232 1007 1236
rect 1011 1232 1012 1236
rect 1006 1231 1012 1232
rect 1070 1236 1076 1237
rect 1070 1232 1071 1236
rect 1075 1232 1076 1236
rect 1070 1231 1076 1232
rect 1240 1230 1242 1237
rect 1280 1230 1282 1237
rect 1302 1236 1308 1237
rect 1302 1232 1303 1236
rect 1307 1232 1308 1236
rect 1302 1231 1308 1232
rect 1374 1236 1380 1237
rect 1374 1232 1375 1236
rect 1379 1232 1380 1236
rect 1374 1231 1380 1232
rect 1478 1236 1484 1237
rect 1478 1232 1479 1236
rect 1483 1232 1484 1236
rect 1478 1231 1484 1232
rect 1238 1229 1244 1230
rect 1238 1225 1239 1229
rect 1243 1225 1244 1229
rect 1238 1224 1244 1225
rect 1278 1229 1284 1230
rect 1278 1225 1279 1229
rect 1283 1225 1284 1229
rect 1278 1224 1284 1225
rect 654 1215 660 1216
rect 654 1211 655 1215
rect 659 1211 660 1215
rect 654 1210 660 1211
rect 710 1215 716 1216
rect 710 1211 711 1215
rect 715 1211 716 1215
rect 1310 1215 1316 1216
rect 710 1210 716 1211
rect 1238 1212 1244 1213
rect 662 1189 668 1190
rect 662 1185 663 1189
rect 667 1185 668 1189
rect 662 1184 668 1185
rect 582 1179 588 1180
rect 582 1175 583 1179
rect 587 1175 588 1179
rect 664 1175 666 1184
rect 712 1180 714 1210
rect 1238 1208 1239 1212
rect 1243 1208 1244 1212
rect 1238 1207 1244 1208
rect 1278 1212 1284 1213
rect 1278 1208 1279 1212
rect 1283 1208 1284 1212
rect 1310 1211 1311 1215
rect 1315 1211 1316 1215
rect 1310 1210 1316 1211
rect 1278 1207 1284 1208
rect 742 1189 748 1190
rect 742 1185 743 1189
rect 747 1185 748 1189
rect 742 1184 748 1185
rect 814 1189 820 1190
rect 814 1185 815 1189
rect 819 1185 820 1189
rect 814 1184 820 1185
rect 878 1189 884 1190
rect 878 1185 879 1189
rect 883 1185 884 1189
rect 878 1184 884 1185
rect 942 1189 948 1190
rect 942 1185 943 1189
rect 947 1185 948 1189
rect 942 1184 948 1185
rect 1006 1189 1012 1190
rect 1006 1185 1007 1189
rect 1011 1185 1012 1189
rect 1006 1184 1012 1185
rect 1070 1189 1076 1190
rect 1070 1185 1071 1189
rect 1075 1185 1076 1189
rect 1070 1184 1076 1185
rect 710 1179 716 1180
rect 710 1175 711 1179
rect 715 1175 716 1179
rect 744 1175 746 1184
rect 816 1175 818 1184
rect 880 1175 882 1184
rect 944 1175 946 1184
rect 1008 1175 1010 1184
rect 1072 1175 1074 1184
rect 1214 1179 1220 1180
rect 1214 1175 1215 1179
rect 1219 1175 1220 1179
rect 1240 1175 1242 1207
rect 1280 1175 1282 1207
rect 1302 1189 1308 1190
rect 1302 1185 1303 1189
rect 1307 1185 1308 1189
rect 1302 1184 1308 1185
rect 1304 1175 1306 1184
rect 162 1174 168 1175
rect 175 1174 179 1175
rect 222 1174 228 1175
rect 231 1174 235 1175
rect 135 1169 139 1170
rect 112 1137 114 1169
rect 136 1160 138 1169
rect 146 1167 152 1168
rect 146 1163 147 1167
rect 151 1163 152 1167
rect 146 1162 152 1163
rect 134 1159 140 1160
rect 134 1155 135 1159
rect 139 1155 140 1159
rect 134 1154 140 1155
rect 148 1140 150 1162
rect 146 1139 152 1140
rect 110 1136 116 1137
rect 110 1132 111 1136
rect 115 1132 116 1136
rect 146 1135 147 1139
rect 151 1135 152 1139
rect 146 1134 152 1135
rect 156 1132 158 1174
rect 175 1169 179 1170
rect 231 1169 235 1170
rect 239 1174 243 1175
rect 239 1169 243 1170
rect 311 1174 315 1175
rect 311 1169 315 1170
rect 327 1174 331 1175
rect 327 1169 331 1170
rect 399 1174 403 1175
rect 399 1169 403 1170
rect 431 1174 435 1175
rect 431 1169 435 1170
rect 487 1174 491 1175
rect 487 1169 491 1170
rect 535 1174 539 1175
rect 535 1169 539 1170
rect 575 1174 579 1175
rect 582 1174 588 1175
rect 639 1174 643 1175
rect 575 1169 579 1170
rect 639 1169 643 1170
rect 663 1174 667 1175
rect 710 1174 716 1175
rect 743 1174 747 1175
rect 663 1169 667 1170
rect 743 1169 747 1170
rect 815 1174 819 1175
rect 815 1169 819 1170
rect 839 1174 843 1175
rect 839 1169 843 1170
rect 879 1174 883 1175
rect 879 1169 883 1170
rect 919 1174 923 1175
rect 919 1169 923 1170
rect 943 1174 947 1175
rect 943 1169 947 1170
rect 999 1174 1003 1175
rect 999 1169 1003 1170
rect 1007 1174 1011 1175
rect 1007 1169 1011 1170
rect 1071 1174 1075 1175
rect 1071 1169 1075 1170
rect 1143 1174 1147 1175
rect 1143 1169 1147 1170
rect 1191 1174 1195 1175
rect 1214 1174 1220 1175
rect 1239 1174 1243 1175
rect 1191 1169 1195 1170
rect 162 1167 168 1168
rect 162 1163 163 1167
rect 167 1163 168 1167
rect 162 1162 168 1163
rect 110 1131 116 1132
rect 154 1131 160 1132
rect 154 1127 155 1131
rect 159 1127 160 1131
rect 154 1126 160 1127
rect 110 1119 116 1120
rect 110 1115 111 1119
rect 115 1115 116 1119
rect 110 1114 116 1115
rect 112 1103 114 1114
rect 134 1112 140 1113
rect 134 1108 135 1112
rect 139 1108 140 1112
rect 134 1107 140 1108
rect 136 1103 138 1107
rect 111 1102 115 1103
rect 111 1097 115 1098
rect 135 1102 139 1103
rect 135 1097 139 1098
rect 112 1090 114 1097
rect 134 1096 140 1097
rect 134 1092 135 1096
rect 139 1092 140 1096
rect 134 1091 140 1092
rect 110 1089 116 1090
rect 110 1085 111 1089
rect 115 1085 116 1089
rect 110 1084 116 1085
rect 164 1076 166 1162
rect 176 1160 178 1169
rect 240 1160 242 1169
rect 328 1160 330 1169
rect 354 1167 360 1168
rect 354 1163 355 1167
rect 359 1163 360 1167
rect 354 1162 360 1163
rect 174 1159 180 1160
rect 174 1155 175 1159
rect 179 1155 180 1159
rect 174 1154 180 1155
rect 238 1159 244 1160
rect 238 1155 239 1159
rect 243 1155 244 1159
rect 238 1154 244 1155
rect 326 1159 332 1160
rect 326 1155 327 1159
rect 331 1155 332 1159
rect 326 1154 332 1155
rect 356 1132 358 1162
rect 432 1160 434 1169
rect 458 1167 464 1168
rect 458 1163 459 1167
rect 463 1163 464 1167
rect 458 1162 464 1163
rect 430 1159 436 1160
rect 430 1155 431 1159
rect 435 1155 436 1159
rect 430 1154 436 1155
rect 460 1132 462 1162
rect 536 1160 538 1169
rect 562 1167 568 1168
rect 562 1163 563 1167
rect 567 1163 568 1167
rect 562 1162 568 1163
rect 534 1159 540 1160
rect 534 1155 535 1159
rect 539 1155 540 1159
rect 534 1154 540 1155
rect 564 1132 566 1162
rect 640 1160 642 1169
rect 744 1160 746 1169
rect 762 1167 768 1168
rect 762 1163 763 1167
rect 767 1163 768 1167
rect 762 1162 768 1163
rect 770 1167 776 1168
rect 770 1163 771 1167
rect 775 1163 776 1167
rect 770 1162 776 1163
rect 638 1159 644 1160
rect 638 1155 639 1159
rect 643 1155 644 1159
rect 638 1154 644 1155
rect 742 1159 748 1160
rect 742 1155 743 1159
rect 747 1155 748 1159
rect 742 1154 748 1155
rect 354 1131 360 1132
rect 354 1127 355 1131
rect 359 1127 360 1131
rect 354 1126 360 1127
rect 458 1131 464 1132
rect 458 1127 459 1131
rect 463 1127 464 1131
rect 458 1126 464 1127
rect 562 1131 568 1132
rect 562 1127 563 1131
rect 567 1127 568 1131
rect 562 1126 568 1127
rect 346 1123 352 1124
rect 346 1119 347 1123
rect 351 1119 352 1123
rect 346 1118 352 1119
rect 174 1112 180 1113
rect 174 1108 175 1112
rect 179 1108 180 1112
rect 174 1107 180 1108
rect 238 1112 244 1113
rect 238 1108 239 1112
rect 243 1108 244 1112
rect 238 1107 244 1108
rect 326 1112 332 1113
rect 326 1108 327 1112
rect 331 1108 332 1112
rect 326 1107 332 1108
rect 176 1103 178 1107
rect 240 1103 242 1107
rect 328 1103 330 1107
rect 175 1102 179 1103
rect 175 1097 179 1098
rect 239 1102 243 1103
rect 239 1097 243 1098
rect 247 1102 251 1103
rect 247 1097 251 1098
rect 327 1102 331 1103
rect 327 1097 331 1098
rect 174 1096 180 1097
rect 174 1092 175 1096
rect 179 1092 180 1096
rect 174 1091 180 1092
rect 246 1096 252 1097
rect 246 1092 247 1096
rect 251 1092 252 1096
rect 246 1091 252 1092
rect 326 1096 332 1097
rect 326 1092 327 1096
rect 331 1092 332 1096
rect 326 1091 332 1092
rect 162 1075 168 1076
rect 110 1072 116 1073
rect 110 1068 111 1072
rect 115 1068 116 1072
rect 162 1071 163 1075
rect 167 1071 168 1075
rect 162 1070 168 1071
rect 238 1075 244 1076
rect 238 1071 239 1075
rect 243 1071 244 1075
rect 238 1070 244 1071
rect 110 1067 116 1068
rect 142 1067 148 1068
rect 112 1035 114 1067
rect 142 1063 143 1067
rect 147 1063 148 1067
rect 142 1062 148 1063
rect 134 1049 140 1050
rect 134 1045 135 1049
rect 139 1045 140 1049
rect 134 1044 140 1045
rect 136 1035 138 1044
rect 144 1040 146 1062
rect 174 1049 180 1050
rect 174 1045 175 1049
rect 179 1045 180 1049
rect 174 1044 180 1045
rect 142 1039 148 1040
rect 142 1035 143 1039
rect 147 1035 148 1039
rect 176 1035 178 1044
rect 240 1040 242 1070
rect 334 1067 340 1068
rect 334 1063 335 1067
rect 339 1063 340 1067
rect 334 1062 340 1063
rect 246 1049 252 1050
rect 246 1045 247 1049
rect 251 1045 252 1049
rect 246 1044 252 1045
rect 326 1049 332 1050
rect 326 1045 327 1049
rect 331 1045 332 1049
rect 326 1044 332 1045
rect 198 1039 204 1040
rect 198 1035 199 1039
rect 203 1035 204 1039
rect 111 1034 115 1035
rect 111 1029 115 1030
rect 135 1034 139 1035
rect 142 1034 148 1035
rect 175 1034 179 1035
rect 198 1034 204 1035
rect 238 1039 244 1040
rect 238 1035 239 1039
rect 243 1035 244 1039
rect 248 1035 250 1044
rect 328 1035 330 1044
rect 238 1034 244 1035
rect 247 1034 251 1035
rect 135 1029 139 1030
rect 175 1029 179 1030
rect 112 997 114 1029
rect 176 1020 178 1029
rect 174 1019 180 1020
rect 174 1015 175 1019
rect 179 1015 180 1019
rect 174 1014 180 1015
rect 110 996 116 997
rect 110 992 111 996
rect 115 992 116 996
rect 200 992 202 1034
rect 247 1029 251 1030
rect 255 1034 259 1035
rect 255 1029 259 1030
rect 327 1034 331 1035
rect 327 1029 331 1030
rect 238 1027 244 1028
rect 238 1023 239 1027
rect 243 1023 244 1027
rect 238 1022 244 1023
rect 240 992 242 1022
rect 256 1020 258 1029
rect 278 1027 284 1028
rect 278 1023 279 1027
rect 283 1023 284 1027
rect 278 1022 284 1023
rect 254 1019 260 1020
rect 254 1015 255 1019
rect 259 1015 260 1019
rect 254 1014 260 1015
rect 110 991 116 992
rect 198 991 204 992
rect 198 987 199 991
rect 203 987 204 991
rect 198 986 204 987
rect 238 991 244 992
rect 238 987 239 991
rect 243 987 244 991
rect 238 986 244 987
rect 110 979 116 980
rect 110 975 111 979
rect 115 975 116 979
rect 110 974 116 975
rect 112 967 114 974
rect 174 972 180 973
rect 174 968 175 972
rect 179 968 180 972
rect 174 967 180 968
rect 254 972 260 973
rect 254 968 255 972
rect 259 968 260 972
rect 254 967 260 968
rect 111 966 115 967
rect 111 961 115 962
rect 175 966 179 967
rect 175 961 179 962
rect 215 966 219 967
rect 215 961 219 962
rect 255 966 259 967
rect 255 961 259 962
rect 112 954 114 961
rect 214 960 220 961
rect 214 956 215 960
rect 219 956 220 960
rect 214 955 220 956
rect 254 960 260 961
rect 254 956 255 960
rect 259 956 260 960
rect 254 955 260 956
rect 110 953 116 954
rect 110 949 111 953
rect 115 949 116 953
rect 110 948 116 949
rect 280 940 282 1022
rect 328 1020 330 1029
rect 336 1028 338 1062
rect 348 1040 350 1118
rect 430 1112 436 1113
rect 430 1108 431 1112
rect 435 1108 436 1112
rect 430 1107 436 1108
rect 534 1112 540 1113
rect 534 1108 535 1112
rect 539 1108 540 1112
rect 534 1107 540 1108
rect 638 1112 644 1113
rect 638 1108 639 1112
rect 643 1108 644 1112
rect 638 1107 644 1108
rect 742 1112 748 1113
rect 742 1108 743 1112
rect 747 1108 748 1112
rect 742 1107 748 1108
rect 432 1103 434 1107
rect 536 1103 538 1107
rect 640 1103 642 1107
rect 744 1103 746 1107
rect 415 1102 419 1103
rect 415 1097 419 1098
rect 431 1102 435 1103
rect 431 1097 435 1098
rect 503 1102 507 1103
rect 503 1097 507 1098
rect 535 1102 539 1103
rect 535 1097 539 1098
rect 583 1102 587 1103
rect 583 1097 587 1098
rect 639 1102 643 1103
rect 639 1097 643 1098
rect 663 1102 667 1103
rect 663 1097 667 1098
rect 735 1102 739 1103
rect 735 1097 739 1098
rect 743 1102 747 1103
rect 743 1097 747 1098
rect 414 1096 420 1097
rect 414 1092 415 1096
rect 419 1092 420 1096
rect 414 1091 420 1092
rect 502 1096 508 1097
rect 502 1092 503 1096
rect 507 1092 508 1096
rect 502 1091 508 1092
rect 582 1096 588 1097
rect 582 1092 583 1096
rect 587 1092 588 1096
rect 582 1091 588 1092
rect 662 1096 668 1097
rect 662 1092 663 1096
rect 667 1092 668 1096
rect 662 1091 668 1092
rect 734 1096 740 1097
rect 734 1092 735 1096
rect 739 1092 740 1096
rect 734 1091 740 1092
rect 764 1085 766 1162
rect 772 1132 774 1162
rect 840 1160 842 1169
rect 866 1167 872 1168
rect 866 1163 867 1167
rect 871 1163 872 1167
rect 866 1162 872 1163
rect 838 1159 844 1160
rect 838 1155 839 1159
rect 843 1155 844 1159
rect 838 1154 844 1155
rect 868 1132 870 1162
rect 920 1160 922 1169
rect 970 1167 976 1168
rect 970 1163 971 1167
rect 975 1163 976 1167
rect 970 1162 976 1163
rect 918 1159 924 1160
rect 918 1155 919 1159
rect 923 1155 924 1159
rect 918 1154 924 1155
rect 972 1132 974 1162
rect 1000 1160 1002 1169
rect 1026 1167 1032 1168
rect 1026 1163 1027 1167
rect 1031 1163 1032 1167
rect 1026 1162 1032 1163
rect 998 1159 1004 1160
rect 998 1155 999 1159
rect 1003 1155 1004 1159
rect 998 1154 1004 1155
rect 1028 1132 1030 1162
rect 1072 1160 1074 1169
rect 1098 1167 1104 1168
rect 1098 1163 1099 1167
rect 1103 1163 1104 1167
rect 1098 1162 1104 1163
rect 1070 1159 1076 1160
rect 1070 1155 1071 1159
rect 1075 1155 1076 1159
rect 1070 1154 1076 1155
rect 1100 1132 1102 1162
rect 1144 1160 1146 1169
rect 1170 1167 1176 1168
rect 1170 1163 1171 1167
rect 1175 1163 1176 1167
rect 1170 1162 1176 1163
rect 1142 1159 1148 1160
rect 1142 1155 1143 1159
rect 1147 1155 1148 1159
rect 1142 1154 1148 1155
rect 1172 1132 1174 1162
rect 1192 1160 1194 1169
rect 1190 1159 1196 1160
rect 1190 1155 1191 1159
rect 1195 1155 1196 1159
rect 1190 1154 1196 1155
rect 1216 1132 1218 1174
rect 1239 1169 1243 1170
rect 1279 1174 1283 1175
rect 1279 1169 1283 1170
rect 1303 1174 1307 1175
rect 1303 1169 1307 1170
rect 1240 1137 1242 1169
rect 1280 1137 1282 1169
rect 1304 1160 1306 1169
rect 1312 1168 1314 1210
rect 1494 1207 1500 1208
rect 1494 1203 1495 1207
rect 1499 1203 1500 1207
rect 1494 1202 1500 1203
rect 1374 1189 1380 1190
rect 1374 1185 1375 1189
rect 1379 1185 1380 1189
rect 1374 1184 1380 1185
rect 1478 1189 1484 1190
rect 1478 1185 1479 1189
rect 1483 1185 1484 1189
rect 1478 1184 1484 1185
rect 1376 1175 1378 1184
rect 1480 1175 1482 1184
rect 1496 1180 1498 1202
rect 1572 1180 1574 1270
rect 1806 1267 1812 1268
rect 1806 1263 1807 1267
rect 1811 1263 1812 1267
rect 1806 1262 1812 1263
rect 1582 1256 1588 1257
rect 1582 1252 1583 1256
rect 1587 1252 1588 1256
rect 1582 1251 1588 1252
rect 1622 1256 1628 1257
rect 1622 1252 1623 1256
rect 1627 1252 1628 1256
rect 1622 1251 1628 1252
rect 1678 1256 1684 1257
rect 1678 1252 1679 1256
rect 1683 1252 1684 1256
rect 1678 1251 1684 1252
rect 1734 1256 1740 1257
rect 1734 1252 1735 1256
rect 1739 1252 1740 1256
rect 1734 1251 1740 1252
rect 1790 1256 1796 1257
rect 1790 1252 1791 1256
rect 1795 1252 1796 1256
rect 1790 1251 1796 1252
rect 1584 1243 1586 1251
rect 1624 1243 1626 1251
rect 1680 1243 1682 1251
rect 1736 1243 1738 1251
rect 1792 1243 1794 1251
rect 1583 1242 1587 1243
rect 1583 1237 1587 1238
rect 1623 1242 1627 1243
rect 1623 1237 1627 1238
rect 1679 1242 1683 1243
rect 1679 1237 1683 1238
rect 1687 1242 1691 1243
rect 1687 1237 1691 1238
rect 1735 1242 1739 1243
rect 1735 1237 1739 1238
rect 1791 1242 1795 1243
rect 1791 1237 1795 1238
rect 1582 1236 1588 1237
rect 1582 1232 1583 1236
rect 1587 1232 1588 1236
rect 1582 1231 1588 1232
rect 1686 1236 1692 1237
rect 1686 1232 1687 1236
rect 1691 1232 1692 1236
rect 1686 1231 1692 1232
rect 1790 1236 1796 1237
rect 1790 1232 1791 1236
rect 1795 1232 1796 1236
rect 1790 1231 1796 1232
rect 1678 1215 1684 1216
rect 1678 1211 1679 1215
rect 1683 1211 1684 1215
rect 1678 1210 1684 1211
rect 1582 1189 1588 1190
rect 1582 1185 1583 1189
rect 1587 1185 1588 1189
rect 1582 1184 1588 1185
rect 1494 1179 1500 1180
rect 1494 1175 1495 1179
rect 1499 1175 1500 1179
rect 1343 1174 1347 1175
rect 1343 1169 1347 1170
rect 1375 1174 1379 1175
rect 1375 1169 1379 1170
rect 1407 1174 1411 1175
rect 1407 1169 1411 1170
rect 1479 1174 1483 1175
rect 1479 1169 1483 1170
rect 1487 1174 1491 1175
rect 1494 1174 1500 1175
rect 1570 1179 1576 1180
rect 1570 1175 1571 1179
rect 1575 1175 1576 1179
rect 1584 1175 1586 1184
rect 1680 1180 1682 1210
rect 1686 1189 1692 1190
rect 1686 1185 1687 1189
rect 1691 1185 1692 1189
rect 1686 1184 1692 1185
rect 1790 1189 1796 1190
rect 1790 1185 1791 1189
rect 1795 1185 1796 1189
rect 1790 1184 1796 1185
rect 1678 1179 1684 1180
rect 1678 1175 1679 1179
rect 1683 1175 1684 1179
rect 1688 1175 1690 1184
rect 1792 1175 1794 1184
rect 1808 1180 1810 1262
rect 1846 1256 1852 1257
rect 1846 1252 1847 1256
rect 1851 1252 1852 1256
rect 1846 1251 1852 1252
rect 1902 1256 1908 1257
rect 1902 1252 1903 1256
rect 1907 1252 1908 1256
rect 1902 1251 1908 1252
rect 1966 1256 1972 1257
rect 1966 1252 1967 1256
rect 1971 1252 1972 1256
rect 1966 1251 1972 1252
rect 2038 1256 2044 1257
rect 2038 1252 2039 1256
rect 2043 1252 2044 1256
rect 2038 1251 2044 1252
rect 2118 1256 2124 1257
rect 2118 1252 2119 1256
rect 2123 1252 2124 1256
rect 2118 1251 2124 1252
rect 2198 1256 2204 1257
rect 2198 1252 2199 1256
rect 2203 1252 2204 1256
rect 2198 1251 2204 1252
rect 1848 1243 1850 1251
rect 1904 1243 1906 1251
rect 1968 1243 1970 1251
rect 2040 1243 2042 1251
rect 2120 1243 2122 1251
rect 2200 1243 2202 1251
rect 1847 1242 1851 1243
rect 1847 1237 1851 1238
rect 1887 1242 1891 1243
rect 1887 1237 1891 1238
rect 1903 1242 1907 1243
rect 1903 1237 1907 1238
rect 1967 1242 1971 1243
rect 1967 1237 1971 1238
rect 1983 1242 1987 1243
rect 1983 1237 1987 1238
rect 2039 1242 2043 1243
rect 2039 1237 2043 1238
rect 2071 1242 2075 1243
rect 2071 1237 2075 1238
rect 2119 1242 2123 1243
rect 2119 1237 2123 1238
rect 2151 1242 2155 1243
rect 2151 1237 2155 1238
rect 2199 1242 2203 1243
rect 2199 1237 2203 1238
rect 2223 1242 2227 1243
rect 2223 1237 2227 1238
rect 1886 1236 1892 1237
rect 1886 1232 1887 1236
rect 1891 1232 1892 1236
rect 1886 1231 1892 1232
rect 1982 1236 1988 1237
rect 1982 1232 1983 1236
rect 1987 1232 1988 1236
rect 1982 1231 1988 1232
rect 2070 1236 2076 1237
rect 2070 1232 2071 1236
rect 2075 1232 2076 1236
rect 2070 1231 2076 1232
rect 2150 1236 2156 1237
rect 2150 1232 2151 1236
rect 2155 1232 2156 1236
rect 2150 1231 2156 1232
rect 2222 1236 2228 1237
rect 2222 1232 2223 1236
rect 2227 1232 2228 1236
rect 2222 1231 2228 1232
rect 2252 1216 2254 1306
rect 2264 1276 2266 1318
rect 2287 1313 2291 1314
rect 2359 1318 2363 1319
rect 2359 1313 2363 1314
rect 2288 1304 2290 1313
rect 2360 1304 2362 1313
rect 2368 1312 2370 1354
rect 2376 1324 2378 1414
rect 2406 1407 2412 1408
rect 2406 1403 2407 1407
rect 2411 1403 2412 1407
rect 2406 1402 2412 1403
rect 2408 1387 2410 1402
rect 2407 1386 2411 1387
rect 2407 1381 2411 1382
rect 2408 1374 2410 1381
rect 2406 1373 2412 1374
rect 2406 1369 2407 1373
rect 2411 1369 2412 1373
rect 2406 1368 2412 1369
rect 2406 1356 2412 1357
rect 2406 1352 2407 1356
rect 2411 1352 2412 1356
rect 2406 1351 2412 1352
rect 2374 1323 2380 1324
rect 2374 1319 2375 1323
rect 2379 1319 2380 1323
rect 2408 1319 2410 1351
rect 2374 1318 2380 1319
rect 2407 1318 2411 1319
rect 2407 1313 2411 1314
rect 2366 1311 2372 1312
rect 2366 1307 2367 1311
rect 2371 1307 2372 1311
rect 2366 1306 2372 1307
rect 2286 1303 2292 1304
rect 2286 1299 2287 1303
rect 2291 1299 2292 1303
rect 2286 1298 2292 1299
rect 2358 1303 2364 1304
rect 2358 1299 2359 1303
rect 2363 1299 2364 1303
rect 2358 1298 2364 1299
rect 2408 1281 2410 1313
rect 2406 1280 2412 1281
rect 2406 1276 2407 1280
rect 2411 1276 2412 1280
rect 2262 1275 2268 1276
rect 2262 1271 2263 1275
rect 2267 1271 2268 1275
rect 2262 1270 2268 1271
rect 2366 1275 2372 1276
rect 2406 1275 2412 1276
rect 2366 1271 2367 1275
rect 2371 1271 2372 1275
rect 2366 1270 2372 1271
rect 2286 1256 2292 1257
rect 2286 1252 2287 1256
rect 2291 1252 2292 1256
rect 2286 1251 2292 1252
rect 2358 1256 2364 1257
rect 2358 1252 2359 1256
rect 2363 1252 2364 1256
rect 2358 1251 2364 1252
rect 2288 1243 2290 1251
rect 2360 1243 2362 1251
rect 2287 1242 2291 1243
rect 2287 1237 2291 1238
rect 2303 1242 2307 1243
rect 2303 1237 2307 1238
rect 2359 1242 2363 1243
rect 2359 1237 2363 1238
rect 2302 1236 2308 1237
rect 2302 1232 2303 1236
rect 2307 1232 2308 1236
rect 2302 1231 2308 1232
rect 2358 1236 2364 1237
rect 2358 1232 2359 1236
rect 2363 1232 2364 1236
rect 2358 1231 2364 1232
rect 1878 1215 1884 1216
rect 1878 1211 1879 1215
rect 1883 1211 1884 1215
rect 1878 1210 1884 1211
rect 1974 1215 1980 1216
rect 1974 1211 1975 1215
rect 1979 1211 1980 1215
rect 1974 1210 1980 1211
rect 2062 1215 2068 1216
rect 2062 1211 2063 1215
rect 2067 1211 2068 1215
rect 2062 1210 2068 1211
rect 2142 1215 2148 1216
rect 2142 1211 2143 1215
rect 2147 1211 2148 1215
rect 2142 1210 2148 1211
rect 2250 1215 2256 1216
rect 2250 1211 2251 1215
rect 2255 1211 2256 1215
rect 2250 1210 2256 1211
rect 2350 1215 2356 1216
rect 2350 1211 2351 1215
rect 2355 1211 2356 1215
rect 2350 1210 2356 1211
rect 1880 1180 1882 1210
rect 1910 1207 1916 1208
rect 1910 1203 1911 1207
rect 1915 1203 1916 1207
rect 1910 1202 1916 1203
rect 1886 1189 1892 1190
rect 1886 1185 1887 1189
rect 1891 1185 1892 1189
rect 1886 1184 1892 1185
rect 1806 1179 1812 1180
rect 1806 1175 1807 1179
rect 1811 1175 1812 1179
rect 1570 1174 1576 1175
rect 1583 1174 1587 1175
rect 1678 1174 1684 1175
rect 1687 1174 1691 1175
rect 1487 1169 1491 1170
rect 1583 1169 1587 1170
rect 1687 1169 1691 1170
rect 1791 1174 1795 1175
rect 1791 1169 1795 1170
rect 1799 1174 1803 1175
rect 1806 1174 1812 1175
rect 1878 1179 1884 1180
rect 1878 1175 1879 1179
rect 1883 1175 1884 1179
rect 1888 1175 1890 1184
rect 1878 1174 1884 1175
rect 1887 1174 1891 1175
rect 1799 1169 1803 1170
rect 1887 1169 1891 1170
rect 1903 1174 1907 1175
rect 1903 1169 1907 1170
rect 1310 1167 1316 1168
rect 1310 1163 1311 1167
rect 1315 1163 1316 1167
rect 1310 1162 1316 1163
rect 1330 1167 1336 1168
rect 1330 1163 1331 1167
rect 1335 1163 1336 1167
rect 1330 1162 1336 1163
rect 1302 1159 1308 1160
rect 1302 1155 1303 1159
rect 1307 1155 1308 1159
rect 1302 1154 1308 1155
rect 1238 1136 1244 1137
rect 1238 1132 1239 1136
rect 1243 1132 1244 1136
rect 770 1131 776 1132
rect 770 1127 771 1131
rect 775 1127 776 1131
rect 770 1126 776 1127
rect 866 1131 872 1132
rect 866 1127 867 1131
rect 871 1127 872 1131
rect 866 1126 872 1127
rect 970 1131 976 1132
rect 970 1127 971 1131
rect 975 1127 976 1131
rect 970 1126 976 1127
rect 1026 1131 1032 1132
rect 1026 1127 1027 1131
rect 1031 1127 1032 1131
rect 1026 1126 1032 1127
rect 1098 1131 1104 1132
rect 1098 1127 1099 1131
rect 1103 1127 1104 1131
rect 1098 1126 1104 1127
rect 1170 1131 1176 1132
rect 1170 1127 1171 1131
rect 1175 1127 1176 1131
rect 1170 1126 1176 1127
rect 1214 1131 1220 1132
rect 1238 1131 1244 1132
rect 1278 1136 1284 1137
rect 1278 1132 1279 1136
rect 1283 1132 1284 1136
rect 1332 1132 1334 1162
rect 1344 1160 1346 1169
rect 1408 1160 1410 1169
rect 1434 1167 1440 1168
rect 1434 1163 1435 1167
rect 1439 1163 1440 1167
rect 1434 1162 1440 1163
rect 1342 1159 1348 1160
rect 1342 1155 1343 1159
rect 1347 1155 1348 1159
rect 1342 1154 1348 1155
rect 1406 1159 1412 1160
rect 1406 1155 1407 1159
rect 1411 1155 1412 1159
rect 1406 1154 1412 1155
rect 1436 1132 1438 1162
rect 1488 1160 1490 1169
rect 1514 1167 1520 1168
rect 1514 1163 1515 1167
rect 1519 1163 1520 1167
rect 1514 1162 1520 1163
rect 1486 1159 1492 1160
rect 1486 1155 1487 1159
rect 1491 1155 1492 1159
rect 1486 1154 1492 1155
rect 1516 1132 1518 1162
rect 1584 1160 1586 1169
rect 1610 1167 1616 1168
rect 1610 1163 1611 1167
rect 1615 1163 1616 1167
rect 1610 1162 1616 1163
rect 1582 1159 1588 1160
rect 1582 1155 1583 1159
rect 1587 1155 1588 1159
rect 1582 1154 1588 1155
rect 1612 1132 1614 1162
rect 1688 1160 1690 1169
rect 1714 1167 1720 1168
rect 1714 1163 1715 1167
rect 1719 1163 1720 1167
rect 1714 1162 1720 1163
rect 1686 1159 1692 1160
rect 1686 1155 1687 1159
rect 1691 1155 1692 1159
rect 1686 1154 1692 1155
rect 1716 1132 1718 1162
rect 1800 1160 1802 1169
rect 1904 1160 1906 1169
rect 1912 1168 1914 1202
rect 1976 1180 1978 1210
rect 1982 1189 1988 1190
rect 1982 1185 1983 1189
rect 1987 1185 1988 1189
rect 1982 1184 1988 1185
rect 1974 1179 1980 1180
rect 1974 1175 1975 1179
rect 1979 1175 1980 1179
rect 1984 1175 1986 1184
rect 2064 1180 2066 1210
rect 2070 1189 2076 1190
rect 2070 1185 2071 1189
rect 2075 1185 2076 1189
rect 2070 1184 2076 1185
rect 2062 1179 2068 1180
rect 2062 1175 2063 1179
rect 2067 1175 2068 1179
rect 2072 1175 2074 1184
rect 2144 1180 2146 1210
rect 2310 1207 2316 1208
rect 2310 1203 2311 1207
rect 2315 1203 2316 1207
rect 2310 1202 2316 1203
rect 2150 1189 2156 1190
rect 2150 1185 2151 1189
rect 2155 1185 2156 1189
rect 2150 1184 2156 1185
rect 2222 1189 2228 1190
rect 2222 1185 2223 1189
rect 2227 1185 2228 1189
rect 2222 1184 2228 1185
rect 2302 1189 2308 1190
rect 2302 1185 2303 1189
rect 2307 1185 2308 1189
rect 2302 1184 2308 1185
rect 2142 1179 2148 1180
rect 2142 1175 2143 1179
rect 2147 1175 2148 1179
rect 2152 1175 2154 1184
rect 2186 1179 2192 1180
rect 2186 1175 2187 1179
rect 2191 1175 2192 1179
rect 2224 1175 2226 1184
rect 2304 1175 2306 1184
rect 2312 1180 2314 1202
rect 2310 1179 2316 1180
rect 2310 1175 2311 1179
rect 2315 1175 2316 1179
rect 1974 1174 1980 1175
rect 1983 1174 1987 1175
rect 1983 1169 1987 1170
rect 1999 1174 2003 1175
rect 2062 1174 2068 1175
rect 2071 1174 2075 1175
rect 1999 1169 2003 1170
rect 2071 1169 2075 1170
rect 2079 1174 2083 1175
rect 2142 1174 2148 1175
rect 2151 1174 2155 1175
rect 2079 1169 2083 1170
rect 2151 1169 2155 1170
rect 2159 1174 2163 1175
rect 2186 1174 2192 1175
rect 2223 1174 2227 1175
rect 2159 1169 2163 1170
rect 1910 1167 1916 1168
rect 1910 1163 1911 1167
rect 1915 1163 1916 1167
rect 1910 1162 1916 1163
rect 1930 1167 1936 1168
rect 1930 1163 1931 1167
rect 1935 1163 1936 1167
rect 1930 1162 1936 1163
rect 1798 1159 1804 1160
rect 1798 1155 1799 1159
rect 1803 1155 1804 1159
rect 1798 1154 1804 1155
rect 1902 1159 1908 1160
rect 1902 1155 1903 1159
rect 1907 1155 1908 1159
rect 1902 1154 1908 1155
rect 1932 1132 1934 1162
rect 2000 1160 2002 1169
rect 2026 1167 2032 1168
rect 2026 1163 2027 1167
rect 2031 1163 2032 1167
rect 2026 1162 2032 1163
rect 1998 1159 2004 1160
rect 1998 1155 1999 1159
rect 2003 1155 2004 1159
rect 1998 1154 2004 1155
rect 2028 1132 2030 1162
rect 2080 1160 2082 1169
rect 2160 1160 2162 1169
rect 2078 1159 2084 1160
rect 2078 1155 2079 1159
rect 2083 1155 2084 1159
rect 2078 1154 2084 1155
rect 2158 1159 2164 1160
rect 2158 1155 2159 1159
rect 2163 1155 2164 1159
rect 2158 1154 2164 1155
rect 2188 1132 2190 1174
rect 2223 1169 2227 1170
rect 2231 1174 2235 1175
rect 2231 1169 2235 1170
rect 2303 1174 2307 1175
rect 2310 1174 2316 1175
rect 2303 1169 2307 1170
rect 2232 1160 2234 1169
rect 2290 1167 2296 1168
rect 2290 1163 2291 1167
rect 2295 1163 2296 1167
rect 2290 1162 2296 1163
rect 2230 1159 2236 1160
rect 2230 1155 2231 1159
rect 2235 1155 2236 1159
rect 2230 1154 2236 1155
rect 2292 1132 2294 1162
rect 2304 1160 2306 1169
rect 2352 1168 2354 1210
rect 2358 1189 2364 1190
rect 2358 1185 2359 1189
rect 2363 1185 2364 1189
rect 2358 1184 2364 1185
rect 2360 1175 2362 1184
rect 2368 1180 2370 1270
rect 2406 1263 2412 1264
rect 2406 1259 2407 1263
rect 2411 1259 2412 1263
rect 2406 1258 2412 1259
rect 2408 1243 2410 1258
rect 2407 1242 2411 1243
rect 2407 1237 2411 1238
rect 2408 1230 2410 1237
rect 2406 1229 2412 1230
rect 2406 1225 2407 1229
rect 2411 1225 2412 1229
rect 2406 1224 2412 1225
rect 2406 1212 2412 1213
rect 2406 1208 2407 1212
rect 2411 1208 2412 1212
rect 2406 1207 2412 1208
rect 2366 1179 2372 1180
rect 2366 1175 2367 1179
rect 2371 1175 2372 1179
rect 2408 1175 2410 1207
rect 2359 1174 2363 1175
rect 2366 1174 2372 1175
rect 2407 1174 2411 1175
rect 2359 1169 2363 1170
rect 2407 1169 2411 1170
rect 2342 1167 2348 1168
rect 2342 1163 2343 1167
rect 2347 1163 2348 1167
rect 2342 1162 2348 1163
rect 2350 1167 2356 1168
rect 2350 1163 2351 1167
rect 2355 1163 2356 1167
rect 2350 1162 2356 1163
rect 2302 1159 2308 1160
rect 2302 1155 2303 1159
rect 2307 1155 2308 1159
rect 2302 1154 2308 1155
rect 2344 1132 2346 1162
rect 2360 1160 2362 1169
rect 2358 1159 2364 1160
rect 2358 1155 2359 1159
rect 2363 1155 2364 1159
rect 2358 1154 2364 1155
rect 2408 1137 2410 1169
rect 2406 1136 2412 1137
rect 2406 1132 2407 1136
rect 2411 1132 2412 1136
rect 1278 1131 1284 1132
rect 1330 1131 1336 1132
rect 1214 1127 1215 1131
rect 1219 1127 1220 1131
rect 1214 1126 1220 1127
rect 1330 1127 1331 1131
rect 1335 1127 1336 1131
rect 1330 1126 1336 1127
rect 1434 1131 1440 1132
rect 1434 1127 1435 1131
rect 1439 1127 1440 1131
rect 1434 1126 1440 1127
rect 1514 1131 1520 1132
rect 1514 1127 1515 1131
rect 1519 1127 1520 1131
rect 1514 1126 1520 1127
rect 1610 1131 1616 1132
rect 1610 1127 1611 1131
rect 1615 1127 1616 1131
rect 1610 1126 1616 1127
rect 1714 1131 1720 1132
rect 1714 1127 1715 1131
rect 1719 1127 1720 1131
rect 1714 1126 1720 1127
rect 1734 1131 1740 1132
rect 1734 1127 1735 1131
rect 1739 1127 1740 1131
rect 1734 1126 1740 1127
rect 1930 1131 1936 1132
rect 1930 1127 1931 1131
rect 1935 1127 1936 1131
rect 1930 1126 1936 1127
rect 2026 1131 2032 1132
rect 2026 1127 2027 1131
rect 2031 1127 2032 1131
rect 2026 1126 2032 1127
rect 2166 1131 2172 1132
rect 2166 1127 2167 1131
rect 2171 1127 2172 1131
rect 2166 1126 2172 1127
rect 2186 1131 2192 1132
rect 2186 1127 2187 1131
rect 2191 1127 2192 1131
rect 2186 1126 2192 1127
rect 2290 1131 2296 1132
rect 2290 1127 2291 1131
rect 2295 1127 2296 1131
rect 2290 1126 2296 1127
rect 2342 1131 2348 1132
rect 2406 1131 2412 1132
rect 2342 1127 2343 1131
rect 2347 1127 2348 1131
rect 2342 1126 2348 1127
rect 1238 1119 1244 1120
rect 1238 1115 1239 1119
rect 1243 1115 1244 1119
rect 1238 1114 1244 1115
rect 1278 1119 1284 1120
rect 1278 1115 1279 1119
rect 1283 1115 1284 1119
rect 1278 1114 1284 1115
rect 838 1112 844 1113
rect 838 1108 839 1112
rect 843 1108 844 1112
rect 838 1107 844 1108
rect 918 1112 924 1113
rect 918 1108 919 1112
rect 923 1108 924 1112
rect 918 1107 924 1108
rect 998 1112 1004 1113
rect 998 1108 999 1112
rect 1003 1108 1004 1112
rect 998 1107 1004 1108
rect 1070 1112 1076 1113
rect 1070 1108 1071 1112
rect 1075 1108 1076 1112
rect 1070 1107 1076 1108
rect 1142 1112 1148 1113
rect 1142 1108 1143 1112
rect 1147 1108 1148 1112
rect 1142 1107 1148 1108
rect 1190 1112 1196 1113
rect 1190 1108 1191 1112
rect 1195 1108 1196 1112
rect 1190 1107 1196 1108
rect 840 1103 842 1107
rect 920 1103 922 1107
rect 1000 1103 1002 1107
rect 1072 1103 1074 1107
rect 1144 1103 1146 1107
rect 1192 1103 1194 1107
rect 1240 1103 1242 1114
rect 1280 1107 1282 1114
rect 1302 1112 1308 1113
rect 1302 1108 1303 1112
rect 1307 1108 1308 1112
rect 1302 1107 1308 1108
rect 1342 1112 1348 1113
rect 1342 1108 1343 1112
rect 1347 1108 1348 1112
rect 1342 1107 1348 1108
rect 1406 1112 1412 1113
rect 1406 1108 1407 1112
rect 1411 1108 1412 1112
rect 1406 1107 1412 1108
rect 1486 1112 1492 1113
rect 1486 1108 1487 1112
rect 1491 1108 1492 1112
rect 1486 1107 1492 1108
rect 1582 1112 1588 1113
rect 1582 1108 1583 1112
rect 1587 1108 1588 1112
rect 1582 1107 1588 1108
rect 1686 1112 1692 1113
rect 1686 1108 1687 1112
rect 1691 1108 1692 1112
rect 1686 1107 1692 1108
rect 1279 1106 1283 1107
rect 799 1102 803 1103
rect 799 1097 803 1098
rect 839 1102 843 1103
rect 839 1097 843 1098
rect 863 1102 867 1103
rect 863 1097 867 1098
rect 919 1102 923 1103
rect 919 1097 923 1098
rect 983 1102 987 1103
rect 983 1097 987 1098
rect 999 1102 1003 1103
rect 999 1097 1003 1098
rect 1047 1102 1051 1103
rect 1047 1097 1051 1098
rect 1071 1102 1075 1103
rect 1071 1097 1075 1098
rect 1143 1102 1147 1103
rect 1143 1097 1147 1098
rect 1191 1102 1195 1103
rect 1191 1097 1195 1098
rect 1239 1102 1243 1103
rect 1279 1101 1283 1102
rect 1303 1106 1307 1107
rect 1303 1101 1307 1102
rect 1343 1106 1347 1107
rect 1343 1101 1347 1102
rect 1407 1106 1411 1107
rect 1407 1101 1411 1102
rect 1431 1106 1435 1107
rect 1431 1101 1435 1102
rect 1471 1106 1475 1107
rect 1471 1101 1475 1102
rect 1487 1106 1491 1107
rect 1487 1101 1491 1102
rect 1511 1106 1515 1107
rect 1511 1101 1515 1102
rect 1559 1106 1563 1107
rect 1559 1101 1563 1102
rect 1583 1106 1587 1107
rect 1583 1101 1587 1102
rect 1615 1106 1619 1107
rect 1615 1101 1619 1102
rect 1671 1106 1675 1107
rect 1671 1101 1675 1102
rect 1687 1106 1691 1107
rect 1687 1101 1691 1102
rect 1727 1106 1731 1107
rect 1727 1101 1731 1102
rect 1239 1097 1243 1098
rect 798 1096 804 1097
rect 798 1092 799 1096
rect 803 1092 804 1096
rect 798 1091 804 1092
rect 862 1096 868 1097
rect 862 1092 863 1096
rect 867 1092 868 1096
rect 862 1091 868 1092
rect 918 1096 924 1097
rect 918 1092 919 1096
rect 923 1092 924 1096
rect 918 1091 924 1092
rect 982 1096 988 1097
rect 982 1092 983 1096
rect 987 1092 988 1096
rect 982 1091 988 1092
rect 1046 1096 1052 1097
rect 1046 1092 1047 1096
rect 1051 1092 1052 1096
rect 1046 1091 1052 1092
rect 1240 1090 1242 1097
rect 1280 1094 1282 1101
rect 1430 1100 1436 1101
rect 1430 1096 1431 1100
rect 1435 1096 1436 1100
rect 1430 1095 1436 1096
rect 1470 1100 1476 1101
rect 1470 1096 1471 1100
rect 1475 1096 1476 1100
rect 1470 1095 1476 1096
rect 1510 1100 1516 1101
rect 1510 1096 1511 1100
rect 1515 1096 1516 1100
rect 1510 1095 1516 1096
rect 1558 1100 1564 1101
rect 1558 1096 1559 1100
rect 1563 1096 1564 1100
rect 1558 1095 1564 1096
rect 1614 1100 1620 1101
rect 1614 1096 1615 1100
rect 1619 1096 1620 1100
rect 1614 1095 1620 1096
rect 1670 1100 1676 1101
rect 1670 1096 1671 1100
rect 1675 1096 1676 1100
rect 1670 1095 1676 1096
rect 1726 1100 1732 1101
rect 1726 1096 1727 1100
rect 1731 1096 1732 1100
rect 1726 1095 1732 1096
rect 1278 1093 1284 1094
rect 1238 1089 1244 1090
rect 1238 1085 1239 1089
rect 1243 1085 1244 1089
rect 1278 1089 1279 1093
rect 1283 1089 1284 1093
rect 1278 1088 1284 1089
rect 763 1084 767 1085
rect 763 1079 767 1080
rect 1071 1084 1075 1085
rect 1238 1084 1244 1085
rect 1071 1079 1075 1080
rect 1458 1079 1464 1080
rect 1072 1076 1074 1079
rect 1278 1076 1284 1077
rect 406 1075 412 1076
rect 406 1071 407 1075
rect 411 1071 412 1075
rect 406 1070 412 1071
rect 494 1075 500 1076
rect 494 1071 495 1075
rect 499 1071 500 1075
rect 494 1070 500 1071
rect 726 1075 732 1076
rect 726 1071 727 1075
rect 731 1071 732 1075
rect 726 1070 732 1071
rect 790 1075 796 1076
rect 790 1071 791 1075
rect 795 1071 796 1075
rect 790 1070 796 1071
rect 854 1075 860 1076
rect 854 1071 855 1075
rect 859 1071 860 1075
rect 854 1070 860 1071
rect 910 1075 916 1076
rect 910 1071 911 1075
rect 915 1071 916 1075
rect 910 1070 916 1071
rect 974 1075 980 1076
rect 974 1071 975 1075
rect 979 1071 980 1075
rect 974 1070 980 1071
rect 1038 1075 1044 1076
rect 1038 1071 1039 1075
rect 1043 1071 1044 1075
rect 1038 1070 1044 1071
rect 1070 1075 1076 1076
rect 1070 1071 1071 1075
rect 1075 1071 1076 1075
rect 1070 1070 1076 1071
rect 1238 1072 1244 1073
rect 408 1040 410 1070
rect 414 1049 420 1050
rect 414 1045 415 1049
rect 419 1045 420 1049
rect 414 1044 420 1045
rect 346 1039 352 1040
rect 346 1035 347 1039
rect 351 1035 352 1039
rect 406 1039 412 1040
rect 406 1035 407 1039
rect 411 1035 412 1039
rect 416 1035 418 1044
rect 496 1040 498 1070
rect 502 1049 508 1050
rect 502 1045 503 1049
rect 507 1045 508 1049
rect 502 1044 508 1045
rect 582 1049 588 1050
rect 582 1045 583 1049
rect 587 1045 588 1049
rect 582 1044 588 1045
rect 662 1049 668 1050
rect 662 1045 663 1049
rect 667 1045 668 1049
rect 662 1044 668 1045
rect 494 1039 500 1040
rect 494 1035 495 1039
rect 499 1035 500 1039
rect 504 1035 506 1044
rect 584 1035 586 1044
rect 664 1035 666 1044
rect 728 1040 730 1070
rect 734 1049 740 1050
rect 734 1045 735 1049
rect 739 1045 740 1049
rect 734 1044 740 1045
rect 718 1039 724 1040
rect 718 1035 719 1039
rect 723 1035 724 1039
rect 346 1034 352 1035
rect 399 1034 403 1035
rect 406 1034 412 1035
rect 415 1034 419 1035
rect 399 1029 403 1030
rect 415 1029 419 1030
rect 463 1034 467 1035
rect 494 1034 500 1035
rect 503 1034 507 1035
rect 463 1029 467 1030
rect 503 1029 507 1030
rect 519 1034 523 1035
rect 519 1029 523 1030
rect 575 1034 579 1035
rect 575 1029 579 1030
rect 583 1034 587 1035
rect 583 1029 587 1030
rect 623 1034 627 1035
rect 623 1029 627 1030
rect 663 1034 667 1035
rect 663 1029 667 1030
rect 671 1034 675 1035
rect 718 1034 724 1035
rect 726 1039 732 1040
rect 726 1035 727 1039
rect 731 1035 732 1039
rect 736 1035 738 1044
rect 792 1040 794 1070
rect 798 1049 804 1050
rect 798 1045 799 1049
rect 803 1045 804 1049
rect 798 1044 804 1045
rect 790 1039 796 1040
rect 790 1035 791 1039
rect 795 1035 796 1039
rect 800 1035 802 1044
rect 856 1040 858 1070
rect 862 1049 868 1050
rect 862 1045 863 1049
rect 867 1045 868 1049
rect 862 1044 868 1045
rect 854 1039 860 1040
rect 854 1035 855 1039
rect 859 1035 860 1039
rect 864 1035 866 1044
rect 912 1040 914 1070
rect 918 1049 924 1050
rect 918 1045 919 1049
rect 923 1045 924 1049
rect 918 1044 924 1045
rect 910 1039 916 1040
rect 910 1035 911 1039
rect 915 1035 916 1039
rect 920 1035 922 1044
rect 976 1040 978 1070
rect 982 1049 988 1050
rect 982 1045 983 1049
rect 987 1045 988 1049
rect 982 1044 988 1045
rect 974 1039 980 1040
rect 974 1035 975 1039
rect 979 1035 980 1039
rect 984 1035 986 1044
rect 1040 1040 1042 1070
rect 1238 1068 1239 1072
rect 1243 1068 1244 1072
rect 1278 1072 1279 1076
rect 1283 1072 1284 1076
rect 1458 1075 1459 1079
rect 1463 1075 1464 1079
rect 1458 1074 1464 1075
rect 1498 1079 1504 1080
rect 1498 1075 1499 1079
rect 1503 1075 1504 1079
rect 1498 1074 1504 1075
rect 1550 1079 1556 1080
rect 1550 1075 1551 1079
rect 1555 1075 1556 1079
rect 1550 1074 1556 1075
rect 1606 1079 1612 1080
rect 1606 1075 1607 1079
rect 1611 1075 1612 1079
rect 1606 1074 1612 1075
rect 1662 1079 1668 1080
rect 1662 1075 1663 1079
rect 1667 1075 1668 1079
rect 1662 1074 1668 1075
rect 1714 1079 1720 1080
rect 1714 1075 1715 1079
rect 1719 1075 1720 1079
rect 1714 1074 1720 1075
rect 1278 1071 1284 1072
rect 1238 1067 1244 1068
rect 1046 1049 1052 1050
rect 1046 1045 1047 1049
rect 1051 1045 1052 1049
rect 1046 1044 1052 1045
rect 1038 1039 1044 1040
rect 1038 1035 1039 1039
rect 1043 1035 1044 1039
rect 1048 1035 1050 1044
rect 1240 1035 1242 1067
rect 1280 1039 1282 1071
rect 1439 1068 1443 1069
rect 1439 1063 1443 1064
rect 1430 1053 1436 1054
rect 1430 1049 1431 1053
rect 1435 1049 1436 1053
rect 1430 1048 1436 1049
rect 1432 1039 1434 1048
rect 1440 1044 1442 1063
rect 1460 1044 1462 1074
rect 1470 1053 1476 1054
rect 1470 1049 1471 1053
rect 1475 1049 1476 1053
rect 1470 1048 1476 1049
rect 1438 1043 1444 1044
rect 1438 1039 1439 1043
rect 1443 1039 1444 1043
rect 1279 1038 1283 1039
rect 726 1034 732 1035
rect 735 1034 739 1035
rect 790 1034 796 1035
rect 799 1034 803 1035
rect 671 1029 675 1030
rect 334 1027 340 1028
rect 334 1023 335 1027
rect 339 1023 340 1027
rect 334 1022 340 1023
rect 354 1027 360 1028
rect 354 1023 355 1027
rect 359 1023 360 1027
rect 354 1022 360 1023
rect 326 1019 332 1020
rect 326 1015 327 1019
rect 331 1015 332 1019
rect 326 1014 332 1015
rect 356 992 358 1022
rect 400 1020 402 1029
rect 426 1027 432 1028
rect 426 1023 427 1027
rect 431 1023 432 1027
rect 426 1022 432 1023
rect 398 1019 404 1020
rect 398 1015 399 1019
rect 403 1015 404 1019
rect 398 1014 404 1015
rect 428 992 430 1022
rect 464 1020 466 1029
rect 490 1027 496 1028
rect 490 1023 491 1027
rect 495 1023 496 1027
rect 490 1022 496 1023
rect 462 1019 468 1020
rect 462 1015 463 1019
rect 467 1015 468 1019
rect 462 1014 468 1015
rect 492 992 494 1022
rect 520 1020 522 1029
rect 546 1027 552 1028
rect 546 1023 547 1027
rect 551 1023 552 1027
rect 546 1022 552 1023
rect 518 1019 524 1020
rect 518 1015 519 1019
rect 523 1015 524 1019
rect 518 1014 524 1015
rect 548 992 550 1022
rect 576 1020 578 1029
rect 624 1020 626 1029
rect 630 1027 636 1028
rect 630 1023 631 1027
rect 635 1023 636 1027
rect 630 1022 636 1023
rect 650 1027 656 1028
rect 650 1023 651 1027
rect 655 1023 656 1027
rect 650 1022 656 1023
rect 574 1019 580 1020
rect 574 1015 575 1019
rect 579 1015 580 1019
rect 574 1014 580 1015
rect 622 1019 628 1020
rect 622 1015 623 1019
rect 627 1015 628 1019
rect 622 1014 628 1015
rect 354 991 360 992
rect 354 987 355 991
rect 359 987 360 991
rect 354 986 360 987
rect 426 991 432 992
rect 426 987 427 991
rect 431 987 432 991
rect 426 986 432 987
rect 490 991 496 992
rect 490 987 491 991
rect 495 987 496 991
rect 490 986 496 987
rect 546 991 552 992
rect 546 987 547 991
rect 551 987 552 991
rect 546 986 552 987
rect 470 983 476 984
rect 470 979 471 983
rect 475 979 476 983
rect 470 978 476 979
rect 326 972 332 973
rect 326 968 327 972
rect 331 968 332 972
rect 326 967 332 968
rect 398 972 404 973
rect 398 968 399 972
rect 403 968 404 972
rect 398 967 404 968
rect 462 972 468 973
rect 462 968 463 972
rect 467 968 468 972
rect 462 967 468 968
rect 303 966 307 967
rect 303 961 307 962
rect 327 966 331 967
rect 327 961 331 962
rect 359 966 363 967
rect 359 961 363 962
rect 399 966 403 967
rect 399 961 403 962
rect 415 966 419 967
rect 415 961 419 962
rect 463 966 467 967
rect 463 961 467 962
rect 302 960 308 961
rect 302 956 303 960
rect 307 956 308 960
rect 302 955 308 956
rect 358 960 364 961
rect 358 956 359 960
rect 363 956 364 960
rect 358 955 364 956
rect 414 960 420 961
rect 414 956 415 960
rect 419 956 420 960
rect 414 955 420 956
rect 462 960 468 961
rect 462 956 463 960
rect 467 956 468 960
rect 462 955 468 956
rect 242 939 248 940
rect 110 936 116 937
rect 110 932 111 936
rect 115 932 116 936
rect 242 935 243 939
rect 247 935 248 939
rect 242 934 248 935
rect 278 939 284 940
rect 278 935 279 939
rect 283 935 284 939
rect 278 934 284 935
rect 346 939 352 940
rect 346 935 347 939
rect 351 935 352 939
rect 346 934 352 935
rect 110 931 116 932
rect 222 931 228 932
rect 112 891 114 931
rect 222 927 223 931
rect 227 927 228 931
rect 222 926 228 927
rect 214 913 220 914
rect 214 909 215 913
rect 219 909 220 913
rect 214 908 220 909
rect 216 891 218 908
rect 224 904 226 926
rect 244 904 246 934
rect 254 913 260 914
rect 254 909 255 913
rect 259 909 260 913
rect 254 908 260 909
rect 302 913 308 914
rect 302 909 303 913
rect 307 909 308 913
rect 302 908 308 909
rect 222 903 228 904
rect 222 899 223 903
rect 227 899 228 903
rect 222 898 228 899
rect 242 903 248 904
rect 242 899 243 903
rect 247 899 248 903
rect 242 898 248 899
rect 256 891 258 908
rect 274 891 280 892
rect 304 891 306 908
rect 348 904 350 934
rect 358 913 364 914
rect 358 909 359 913
rect 363 909 364 913
rect 358 908 364 909
rect 414 913 420 914
rect 414 909 415 913
rect 419 909 420 913
rect 414 908 420 909
rect 462 913 468 914
rect 462 909 463 913
rect 467 909 468 913
rect 462 908 468 909
rect 346 903 352 904
rect 346 899 347 903
rect 351 899 352 903
rect 346 898 352 899
rect 360 891 362 908
rect 416 891 418 908
rect 464 891 466 908
rect 472 904 474 978
rect 518 972 524 973
rect 518 968 519 972
rect 523 968 524 972
rect 518 967 524 968
rect 574 972 580 973
rect 574 968 575 972
rect 579 968 580 972
rect 574 967 580 968
rect 622 972 628 973
rect 622 968 623 972
rect 627 968 628 972
rect 622 967 628 968
rect 519 966 523 967
rect 519 961 523 962
rect 575 966 579 967
rect 575 961 579 962
rect 623 966 627 967
rect 623 961 627 962
rect 518 960 524 961
rect 518 956 519 960
rect 523 956 524 960
rect 518 955 524 956
rect 574 960 580 961
rect 574 956 575 960
rect 579 956 580 960
rect 574 955 580 956
rect 632 948 634 1022
rect 652 992 654 1022
rect 672 1020 674 1029
rect 698 1027 704 1028
rect 698 1023 699 1027
rect 703 1023 704 1027
rect 698 1022 704 1023
rect 670 1019 676 1020
rect 670 1015 671 1019
rect 675 1015 676 1019
rect 670 1014 676 1015
rect 700 992 702 1022
rect 720 997 722 1034
rect 735 1029 739 1030
rect 799 1029 803 1030
rect 807 1034 811 1035
rect 854 1034 860 1035
rect 863 1034 867 1035
rect 807 1029 811 1030
rect 863 1029 867 1030
rect 895 1034 899 1035
rect 910 1034 916 1035
rect 919 1034 923 1035
rect 974 1034 980 1035
rect 983 1034 987 1035
rect 895 1029 899 1030
rect 919 1029 923 1030
rect 983 1029 987 1030
rect 999 1034 1003 1035
rect 1038 1034 1044 1035
rect 1047 1034 1051 1035
rect 999 1029 1003 1030
rect 1047 1029 1051 1030
rect 1103 1034 1107 1035
rect 1103 1029 1107 1030
rect 1191 1034 1195 1035
rect 1191 1029 1195 1030
rect 1239 1034 1243 1035
rect 1279 1033 1283 1034
rect 1431 1038 1435 1039
rect 1438 1038 1444 1039
rect 1458 1043 1464 1044
rect 1458 1039 1459 1043
rect 1463 1039 1464 1043
rect 1472 1039 1474 1048
rect 1500 1044 1502 1074
rect 1510 1053 1516 1054
rect 1510 1049 1511 1053
rect 1515 1049 1516 1053
rect 1510 1048 1516 1049
rect 1498 1043 1504 1044
rect 1498 1039 1499 1043
rect 1503 1039 1504 1043
rect 1512 1039 1514 1048
rect 1552 1044 1554 1074
rect 1582 1071 1588 1072
rect 1582 1067 1583 1071
rect 1587 1067 1588 1071
rect 1582 1066 1588 1067
rect 1558 1053 1564 1054
rect 1558 1049 1559 1053
rect 1563 1049 1564 1053
rect 1558 1048 1564 1049
rect 1550 1043 1556 1044
rect 1550 1039 1551 1043
rect 1555 1039 1556 1043
rect 1560 1039 1562 1048
rect 1458 1038 1464 1039
rect 1471 1038 1475 1039
rect 1498 1038 1504 1039
rect 1511 1038 1515 1039
rect 1550 1038 1556 1039
rect 1559 1038 1563 1039
rect 1431 1033 1435 1034
rect 1471 1033 1475 1034
rect 1511 1033 1515 1034
rect 1559 1033 1563 1034
rect 1575 1038 1579 1039
rect 1575 1033 1579 1034
rect 1239 1029 1243 1030
rect 736 1020 738 1029
rect 762 1027 768 1028
rect 762 1023 763 1027
rect 767 1023 768 1027
rect 762 1022 768 1023
rect 734 1019 740 1020
rect 734 1015 735 1019
rect 739 1015 740 1019
rect 734 1014 740 1015
rect 719 996 723 997
rect 764 992 766 1022
rect 808 1020 810 1029
rect 834 1027 840 1028
rect 834 1023 835 1027
rect 839 1023 840 1027
rect 834 1022 840 1023
rect 806 1019 812 1020
rect 806 1015 807 1019
rect 811 1015 812 1019
rect 806 1014 812 1015
rect 836 992 838 1022
rect 896 1020 898 1029
rect 926 1027 932 1028
rect 926 1023 927 1027
rect 931 1023 932 1027
rect 926 1022 932 1023
rect 894 1019 900 1020
rect 894 1015 895 1019
rect 899 1015 900 1019
rect 894 1014 900 1015
rect 928 992 930 1022
rect 1000 1020 1002 1029
rect 1026 1027 1032 1028
rect 1026 1023 1027 1027
rect 1031 1023 1032 1027
rect 1026 1022 1032 1023
rect 998 1019 1004 1020
rect 998 1015 999 1019
rect 1003 1015 1004 1019
rect 998 1014 1004 1015
rect 1028 992 1030 1022
rect 1104 1020 1106 1029
rect 1192 1020 1194 1029
rect 1214 1027 1220 1028
rect 1214 1023 1215 1027
rect 1219 1023 1220 1027
rect 1214 1022 1220 1023
rect 1102 1019 1108 1020
rect 1102 1015 1103 1019
rect 1107 1015 1108 1019
rect 1102 1014 1108 1015
rect 1190 1019 1196 1020
rect 1190 1015 1191 1019
rect 1195 1015 1196 1019
rect 1190 1014 1196 1015
rect 1127 996 1131 997
rect 650 991 656 992
rect 650 987 651 991
rect 655 987 656 991
rect 650 986 656 987
rect 698 991 704 992
rect 719 991 723 992
rect 762 991 768 992
rect 698 987 699 991
rect 703 987 704 991
rect 698 986 704 987
rect 762 987 763 991
rect 767 987 768 991
rect 762 986 768 987
rect 834 991 840 992
rect 834 987 835 991
rect 839 987 840 991
rect 834 986 840 987
rect 922 991 930 992
rect 922 987 923 991
rect 927 988 930 991
rect 1026 991 1032 992
rect 927 987 928 988
rect 922 986 928 987
rect 1026 987 1027 991
rect 1031 987 1032 991
rect 1026 986 1032 987
rect 1126 991 1132 992
rect 1126 987 1127 991
rect 1131 987 1132 991
rect 1126 986 1132 987
rect 1150 991 1156 992
rect 1150 987 1151 991
rect 1155 987 1156 991
rect 1150 986 1156 987
rect 670 972 676 973
rect 670 968 671 972
rect 675 968 676 972
rect 670 967 676 968
rect 734 972 740 973
rect 734 968 735 972
rect 739 968 740 972
rect 734 967 740 968
rect 806 972 812 973
rect 806 968 807 972
rect 811 968 812 972
rect 806 967 812 968
rect 894 972 900 973
rect 894 968 895 972
rect 899 968 900 972
rect 894 967 900 968
rect 998 972 1004 973
rect 998 968 999 972
rect 1003 968 1004 972
rect 998 967 1004 968
rect 1102 972 1108 973
rect 1102 968 1103 972
rect 1107 968 1108 972
rect 1102 967 1108 968
rect 639 966 643 967
rect 639 961 643 962
rect 671 966 675 967
rect 671 961 675 962
rect 711 966 715 967
rect 711 961 715 962
rect 735 966 739 967
rect 735 961 739 962
rect 783 966 787 967
rect 783 961 787 962
rect 807 966 811 967
rect 807 961 811 962
rect 855 966 859 967
rect 855 961 859 962
rect 895 966 899 967
rect 895 961 899 962
rect 927 966 931 967
rect 927 961 931 962
rect 999 966 1003 967
rect 999 961 1003 962
rect 1071 966 1075 967
rect 1071 961 1075 962
rect 1103 966 1107 967
rect 1103 961 1107 962
rect 1143 966 1147 967
rect 1143 961 1147 962
rect 638 960 644 961
rect 638 956 639 960
rect 643 956 644 960
rect 638 955 644 956
rect 710 960 716 961
rect 710 956 711 960
rect 715 956 716 960
rect 710 955 716 956
rect 782 960 788 961
rect 782 956 783 960
rect 787 956 788 960
rect 782 955 788 956
rect 854 960 860 961
rect 854 956 855 960
rect 859 956 860 960
rect 854 955 860 956
rect 926 960 932 961
rect 926 956 927 960
rect 931 956 932 960
rect 926 955 932 956
rect 998 960 1004 961
rect 998 956 999 960
rect 1003 956 1004 960
rect 998 955 1004 956
rect 1070 960 1076 961
rect 1070 956 1071 960
rect 1075 956 1076 960
rect 1070 955 1076 956
rect 1142 960 1148 961
rect 1142 956 1143 960
rect 1147 956 1148 960
rect 1142 955 1148 956
rect 630 947 636 948
rect 630 943 631 947
rect 635 943 636 947
rect 630 942 636 943
rect 502 939 508 940
rect 502 935 503 939
rect 507 935 508 939
rect 502 934 508 935
rect 558 939 564 940
rect 558 935 559 939
rect 563 935 564 939
rect 558 934 564 935
rect 630 939 636 940
rect 630 935 631 939
rect 635 935 636 939
rect 630 934 636 935
rect 702 939 708 940
rect 702 935 703 939
rect 707 935 708 939
rect 702 934 708 935
rect 774 939 780 940
rect 774 935 775 939
rect 779 935 780 939
rect 774 934 780 935
rect 846 939 852 940
rect 846 935 847 939
rect 851 935 852 939
rect 846 934 852 935
rect 990 939 996 940
rect 990 935 991 939
rect 995 935 996 939
rect 990 934 996 935
rect 1014 939 1020 940
rect 1014 935 1015 939
rect 1019 935 1020 939
rect 1014 934 1020 935
rect 504 904 506 934
rect 518 913 524 914
rect 518 909 519 913
rect 523 909 524 913
rect 518 908 524 909
rect 470 903 476 904
rect 470 899 471 903
rect 475 899 476 903
rect 470 898 476 899
rect 502 903 508 904
rect 502 899 503 903
rect 507 899 508 903
rect 502 898 508 899
rect 520 891 522 908
rect 560 904 562 934
rect 574 913 580 914
rect 574 909 575 913
rect 579 909 580 913
rect 574 908 580 909
rect 558 903 564 904
rect 558 899 559 903
rect 563 899 564 903
rect 558 898 564 899
rect 576 891 578 908
rect 632 904 634 934
rect 638 913 644 914
rect 638 909 639 913
rect 643 909 644 913
rect 638 908 644 909
rect 630 903 636 904
rect 630 899 631 903
rect 635 899 636 903
rect 630 898 636 899
rect 640 891 642 908
rect 704 904 706 934
rect 710 913 716 914
rect 710 909 711 913
rect 715 909 716 913
rect 710 908 716 909
rect 702 903 708 904
rect 702 899 703 903
rect 707 899 708 903
rect 702 898 708 899
rect 662 895 668 896
rect 662 891 663 895
rect 667 891 668 895
rect 712 891 714 908
rect 776 904 778 934
rect 782 913 788 914
rect 782 909 783 913
rect 787 909 788 913
rect 782 908 788 909
rect 774 903 780 904
rect 774 899 775 903
rect 779 899 780 903
rect 774 898 780 899
rect 784 891 786 908
rect 848 904 850 934
rect 938 931 944 932
rect 938 927 939 931
rect 943 927 944 931
rect 938 926 944 927
rect 854 913 860 914
rect 854 909 855 913
rect 859 909 860 913
rect 854 908 860 909
rect 926 913 932 914
rect 926 909 927 913
rect 931 909 932 913
rect 926 908 932 909
rect 846 903 852 904
rect 846 899 847 903
rect 851 899 852 903
rect 846 898 852 899
rect 856 891 858 908
rect 928 891 930 908
rect 940 904 942 926
rect 992 904 994 934
rect 998 913 1004 914
rect 998 909 999 913
rect 1003 909 1004 913
rect 998 908 1004 909
rect 938 903 944 904
rect 938 899 939 903
rect 943 899 944 903
rect 938 898 944 899
rect 990 903 996 904
rect 990 899 991 903
rect 995 899 996 903
rect 990 898 996 899
rect 1000 891 1002 908
rect 111 890 115 891
rect 111 885 115 886
rect 191 890 195 891
rect 191 885 195 886
rect 215 890 219 891
rect 215 885 219 886
rect 231 890 235 891
rect 231 885 235 886
rect 255 890 259 891
rect 274 887 275 891
rect 279 887 280 891
rect 274 886 280 887
rect 287 890 291 891
rect 255 885 259 886
rect 112 853 114 885
rect 192 876 194 885
rect 214 879 220 880
rect 190 875 196 876
rect 190 871 191 875
rect 195 871 196 875
rect 214 875 215 879
rect 219 875 220 879
rect 232 876 234 885
rect 254 879 260 880
rect 214 874 220 875
rect 230 875 236 876
rect 190 870 196 871
rect 110 852 116 853
rect 110 848 111 852
rect 115 848 116 852
rect 216 848 218 874
rect 230 871 231 875
rect 235 871 236 875
rect 254 875 255 879
rect 259 875 260 879
rect 254 874 260 875
rect 230 870 236 871
rect 256 848 258 874
rect 110 847 116 848
rect 214 847 220 848
rect 214 843 215 847
rect 219 843 220 847
rect 214 842 220 843
rect 254 847 260 848
rect 254 843 255 847
rect 259 843 260 847
rect 254 842 260 843
rect 110 835 116 836
rect 110 831 111 835
rect 115 831 116 835
rect 110 830 116 831
rect 112 823 114 830
rect 190 828 196 829
rect 190 824 191 828
rect 195 824 196 828
rect 190 823 196 824
rect 230 828 236 829
rect 230 824 231 828
rect 235 824 236 828
rect 230 823 236 824
rect 111 822 115 823
rect 111 817 115 818
rect 135 822 139 823
rect 135 817 139 818
rect 175 822 179 823
rect 175 817 179 818
rect 191 822 195 823
rect 191 817 195 818
rect 231 822 235 823
rect 231 817 235 818
rect 239 822 243 823
rect 239 817 243 818
rect 112 810 114 817
rect 134 816 140 817
rect 134 812 135 816
rect 139 812 140 816
rect 134 811 140 812
rect 174 816 180 817
rect 174 812 175 816
rect 179 812 180 816
rect 174 811 180 812
rect 238 816 244 817
rect 238 812 239 816
rect 243 812 244 816
rect 238 811 244 812
rect 110 809 116 810
rect 110 805 111 809
rect 115 805 116 809
rect 110 804 116 805
rect 276 804 278 886
rect 287 885 291 886
rect 303 890 307 891
rect 303 885 307 886
rect 359 890 363 891
rect 359 885 363 886
rect 415 890 419 891
rect 415 885 419 886
rect 447 890 451 891
rect 447 885 451 886
rect 463 890 467 891
rect 463 885 467 886
rect 519 890 523 891
rect 519 885 523 886
rect 543 890 547 891
rect 543 885 547 886
rect 575 890 579 891
rect 575 885 579 886
rect 639 890 643 891
rect 662 890 668 891
rect 711 890 715 891
rect 639 885 643 886
rect 288 876 290 885
rect 360 876 362 885
rect 386 883 392 884
rect 386 879 387 883
rect 391 879 392 883
rect 386 878 392 879
rect 286 875 292 876
rect 286 871 287 875
rect 291 871 292 875
rect 286 870 292 871
rect 358 875 364 876
rect 358 871 359 875
rect 363 871 364 875
rect 358 870 364 871
rect 388 848 390 878
rect 448 876 450 885
rect 498 883 504 884
rect 498 879 499 883
rect 503 879 504 883
rect 498 878 504 879
rect 446 875 452 876
rect 446 871 447 875
rect 451 871 452 875
rect 446 870 452 871
rect 500 848 502 878
rect 544 876 546 885
rect 602 883 608 884
rect 602 879 603 883
rect 607 879 608 883
rect 602 878 608 879
rect 542 875 548 876
rect 542 871 543 875
rect 547 871 548 875
rect 542 870 548 871
rect 604 848 606 878
rect 640 876 642 885
rect 638 875 644 876
rect 638 871 639 875
rect 643 871 644 875
rect 638 870 644 871
rect 664 848 666 890
rect 711 885 715 886
rect 727 890 731 891
rect 727 885 731 886
rect 783 890 787 891
rect 783 885 787 886
rect 807 890 811 891
rect 807 885 811 886
rect 855 890 859 891
rect 855 885 859 886
rect 887 890 891 891
rect 887 885 891 886
rect 927 890 931 891
rect 927 885 931 886
rect 959 890 963 891
rect 959 885 963 886
rect 999 890 1003 891
rect 999 885 1003 886
rect 728 876 730 885
rect 746 883 752 884
rect 746 879 747 883
rect 751 879 752 883
rect 746 878 752 879
rect 754 883 760 884
rect 754 879 755 883
rect 759 879 760 883
rect 754 878 760 879
rect 726 875 732 876
rect 726 871 727 875
rect 731 871 732 875
rect 726 870 732 871
rect 748 856 750 878
rect 746 855 752 856
rect 746 851 747 855
rect 751 851 752 855
rect 746 850 752 851
rect 756 848 758 878
rect 808 876 810 885
rect 888 876 890 885
rect 946 883 952 884
rect 946 879 947 883
rect 951 879 952 883
rect 946 878 952 879
rect 806 875 812 876
rect 806 871 807 875
rect 811 871 812 875
rect 806 870 812 871
rect 886 875 892 876
rect 886 871 887 875
rect 891 871 892 875
rect 886 870 892 871
rect 948 848 950 878
rect 960 876 962 885
rect 1016 884 1018 934
rect 1070 913 1076 914
rect 1070 909 1071 913
rect 1075 909 1076 913
rect 1070 908 1076 909
rect 1142 913 1148 914
rect 1142 909 1143 913
rect 1147 909 1148 913
rect 1142 908 1148 909
rect 1072 891 1074 908
rect 1144 891 1146 908
rect 1152 904 1154 986
rect 1190 972 1196 973
rect 1190 968 1191 972
rect 1195 968 1196 972
rect 1190 967 1196 968
rect 1191 966 1195 967
rect 1191 961 1195 962
rect 1190 960 1196 961
rect 1190 956 1191 960
rect 1195 956 1196 960
rect 1190 955 1196 956
rect 1216 940 1218 1022
rect 1240 997 1242 1029
rect 1280 1001 1282 1033
rect 1576 1024 1578 1033
rect 1584 1032 1586 1066
rect 1608 1044 1610 1074
rect 1614 1053 1620 1054
rect 1614 1049 1615 1053
rect 1619 1049 1620 1053
rect 1614 1048 1620 1049
rect 1606 1043 1612 1044
rect 1606 1039 1607 1043
rect 1611 1039 1612 1043
rect 1616 1039 1618 1048
rect 1664 1044 1666 1074
rect 1670 1053 1676 1054
rect 1670 1049 1671 1053
rect 1675 1049 1676 1053
rect 1670 1048 1676 1049
rect 1662 1043 1668 1044
rect 1662 1039 1663 1043
rect 1667 1039 1668 1043
rect 1672 1039 1674 1048
rect 1716 1044 1718 1074
rect 1736 1069 1738 1126
rect 1798 1112 1804 1113
rect 1798 1108 1799 1112
rect 1803 1108 1804 1112
rect 1798 1107 1804 1108
rect 1902 1112 1908 1113
rect 1902 1108 1903 1112
rect 1907 1108 1908 1112
rect 1902 1107 1908 1108
rect 1998 1112 2004 1113
rect 1998 1108 1999 1112
rect 2003 1108 2004 1112
rect 1998 1107 2004 1108
rect 2078 1112 2084 1113
rect 2078 1108 2079 1112
rect 2083 1108 2084 1112
rect 2078 1107 2084 1108
rect 2158 1112 2164 1113
rect 2158 1108 2159 1112
rect 2163 1108 2164 1112
rect 2158 1107 2164 1108
rect 1775 1106 1779 1107
rect 1775 1101 1779 1102
rect 1799 1106 1803 1107
rect 1799 1101 1803 1102
rect 1823 1106 1827 1107
rect 1823 1101 1827 1102
rect 1871 1106 1875 1107
rect 1871 1101 1875 1102
rect 1903 1106 1907 1107
rect 1903 1101 1907 1102
rect 1919 1106 1923 1107
rect 1919 1101 1923 1102
rect 1967 1106 1971 1107
rect 1967 1101 1971 1102
rect 1999 1106 2003 1107
rect 1999 1101 2003 1102
rect 2015 1106 2019 1107
rect 2015 1101 2019 1102
rect 2063 1106 2067 1107
rect 2063 1101 2067 1102
rect 2079 1106 2083 1107
rect 2079 1101 2083 1102
rect 2119 1106 2123 1107
rect 2119 1101 2123 1102
rect 2159 1106 2163 1107
rect 2159 1101 2163 1102
rect 1774 1100 1780 1101
rect 1774 1096 1775 1100
rect 1779 1096 1780 1100
rect 1774 1095 1780 1096
rect 1822 1100 1828 1101
rect 1822 1096 1823 1100
rect 1827 1096 1828 1100
rect 1822 1095 1828 1096
rect 1870 1100 1876 1101
rect 1870 1096 1871 1100
rect 1875 1096 1876 1100
rect 1870 1095 1876 1096
rect 1918 1100 1924 1101
rect 1918 1096 1919 1100
rect 1923 1096 1924 1100
rect 1918 1095 1924 1096
rect 1966 1100 1972 1101
rect 1966 1096 1967 1100
rect 1971 1096 1972 1100
rect 1966 1095 1972 1096
rect 2014 1100 2020 1101
rect 2014 1096 2015 1100
rect 2019 1096 2020 1100
rect 2014 1095 2020 1096
rect 2062 1100 2068 1101
rect 2062 1096 2063 1100
rect 2067 1096 2068 1100
rect 2062 1095 2068 1096
rect 2118 1100 2124 1101
rect 2118 1096 2119 1100
rect 2123 1096 2124 1100
rect 2118 1095 2124 1096
rect 1814 1079 1820 1080
rect 1814 1075 1815 1079
rect 1819 1075 1820 1079
rect 1814 1074 1820 1075
rect 2002 1079 2008 1080
rect 2002 1075 2003 1079
rect 2007 1075 2008 1079
rect 2002 1074 2008 1075
rect 1782 1071 1788 1072
rect 1735 1068 1739 1069
rect 1782 1067 1783 1071
rect 1787 1067 1788 1071
rect 1782 1066 1788 1067
rect 1735 1063 1739 1064
rect 1726 1053 1732 1054
rect 1726 1049 1727 1053
rect 1731 1049 1732 1053
rect 1726 1048 1732 1049
rect 1774 1053 1780 1054
rect 1774 1049 1775 1053
rect 1779 1049 1780 1053
rect 1774 1048 1780 1049
rect 1714 1043 1720 1044
rect 1714 1039 1715 1043
rect 1719 1039 1720 1043
rect 1728 1039 1730 1048
rect 1776 1039 1778 1048
rect 1784 1044 1786 1066
rect 1782 1043 1788 1044
rect 1782 1039 1783 1043
rect 1787 1039 1788 1043
rect 1606 1038 1612 1039
rect 1615 1038 1619 1039
rect 1615 1033 1619 1034
rect 1655 1038 1659 1039
rect 1662 1038 1668 1039
rect 1671 1038 1675 1039
rect 1655 1033 1659 1034
rect 1671 1033 1675 1034
rect 1695 1038 1699 1039
rect 1714 1038 1720 1039
rect 1727 1038 1731 1039
rect 1695 1033 1699 1034
rect 1727 1033 1731 1034
rect 1735 1038 1739 1039
rect 1735 1033 1739 1034
rect 1775 1038 1779 1039
rect 1782 1038 1788 1039
rect 1775 1033 1779 1034
rect 1582 1031 1588 1032
rect 1582 1027 1583 1031
rect 1587 1027 1588 1031
rect 1582 1026 1588 1027
rect 1602 1031 1608 1032
rect 1602 1027 1603 1031
rect 1607 1027 1608 1031
rect 1602 1026 1608 1027
rect 1574 1023 1580 1024
rect 1574 1019 1575 1023
rect 1579 1019 1580 1023
rect 1574 1018 1580 1019
rect 1278 1000 1284 1001
rect 1238 996 1244 997
rect 1238 992 1239 996
rect 1243 992 1244 996
rect 1278 996 1279 1000
rect 1283 996 1284 1000
rect 1604 996 1606 1026
rect 1616 1024 1618 1033
rect 1642 1031 1648 1032
rect 1642 1027 1643 1031
rect 1647 1027 1648 1031
rect 1642 1026 1648 1027
rect 1614 1023 1620 1024
rect 1614 1019 1615 1023
rect 1619 1019 1620 1023
rect 1614 1018 1620 1019
rect 1644 996 1646 1026
rect 1656 1024 1658 1033
rect 1682 1031 1688 1032
rect 1682 1027 1683 1031
rect 1687 1027 1688 1031
rect 1682 1026 1688 1027
rect 1654 1023 1660 1024
rect 1654 1019 1655 1023
rect 1659 1019 1660 1023
rect 1654 1018 1660 1019
rect 1684 996 1686 1026
rect 1696 1024 1698 1033
rect 1718 1031 1724 1032
rect 1718 1027 1719 1031
rect 1723 1027 1724 1031
rect 1718 1026 1724 1027
rect 1694 1023 1700 1024
rect 1694 1019 1695 1023
rect 1699 1019 1700 1023
rect 1694 1018 1700 1019
rect 1720 996 1722 1026
rect 1736 1024 1738 1033
rect 1762 1031 1768 1032
rect 1762 1027 1763 1031
rect 1767 1027 1768 1031
rect 1762 1026 1768 1027
rect 1734 1023 1740 1024
rect 1734 1019 1735 1023
rect 1739 1019 1740 1023
rect 1734 1018 1740 1019
rect 1764 996 1766 1026
rect 1776 1024 1778 1033
rect 1816 1032 1818 1074
rect 1822 1053 1828 1054
rect 1822 1049 1823 1053
rect 1827 1049 1828 1053
rect 1822 1048 1828 1049
rect 1870 1053 1876 1054
rect 1870 1049 1871 1053
rect 1875 1049 1876 1053
rect 1870 1048 1876 1049
rect 1918 1053 1924 1054
rect 1918 1049 1919 1053
rect 1923 1049 1924 1053
rect 1918 1048 1924 1049
rect 1966 1053 1972 1054
rect 1966 1049 1967 1053
rect 1971 1049 1972 1053
rect 1966 1048 1972 1049
rect 1824 1039 1826 1048
rect 1872 1039 1874 1048
rect 1920 1039 1922 1048
rect 1968 1039 1970 1048
rect 2004 1044 2006 1074
rect 2014 1053 2020 1054
rect 2014 1049 2015 1053
rect 2019 1049 2020 1053
rect 2014 1048 2020 1049
rect 2062 1053 2068 1054
rect 2062 1049 2063 1053
rect 2067 1049 2068 1053
rect 2062 1048 2068 1049
rect 2118 1053 2124 1054
rect 2118 1049 2119 1053
rect 2123 1049 2124 1053
rect 2118 1048 2124 1049
rect 2002 1043 2008 1044
rect 2002 1039 2003 1043
rect 2007 1039 2008 1043
rect 2016 1039 2018 1048
rect 2064 1039 2066 1048
rect 2110 1043 2116 1044
rect 2110 1039 2111 1043
rect 2115 1039 2116 1043
rect 2120 1039 2122 1048
rect 2168 1044 2170 1126
rect 2406 1119 2412 1120
rect 2406 1115 2407 1119
rect 2411 1115 2412 1119
rect 2406 1114 2412 1115
rect 2230 1112 2236 1113
rect 2230 1108 2231 1112
rect 2235 1108 2236 1112
rect 2230 1107 2236 1108
rect 2302 1112 2308 1113
rect 2302 1108 2303 1112
rect 2307 1108 2308 1112
rect 2302 1107 2308 1108
rect 2358 1112 2364 1113
rect 2358 1108 2359 1112
rect 2363 1108 2364 1112
rect 2358 1107 2364 1108
rect 2408 1107 2410 1114
rect 2175 1106 2179 1107
rect 2175 1101 2179 1102
rect 2231 1106 2235 1107
rect 2231 1101 2235 1102
rect 2303 1106 2307 1107
rect 2303 1101 2307 1102
rect 2359 1106 2363 1107
rect 2359 1101 2363 1102
rect 2407 1106 2411 1107
rect 2407 1101 2411 1102
rect 2174 1100 2180 1101
rect 2174 1096 2175 1100
rect 2179 1096 2180 1100
rect 2174 1095 2180 1096
rect 2230 1100 2236 1101
rect 2230 1096 2231 1100
rect 2235 1096 2236 1100
rect 2230 1095 2236 1096
rect 2408 1094 2410 1101
rect 2406 1093 2412 1094
rect 2406 1089 2407 1093
rect 2411 1089 2412 1093
rect 2406 1088 2412 1089
rect 2222 1079 2228 1080
rect 2222 1075 2223 1079
rect 2227 1075 2228 1079
rect 2222 1074 2228 1075
rect 2246 1079 2252 1080
rect 2246 1075 2247 1079
rect 2251 1075 2252 1079
rect 2246 1074 2252 1075
rect 2406 1076 2412 1077
rect 2174 1053 2180 1054
rect 2174 1049 2175 1053
rect 2179 1049 2180 1053
rect 2174 1048 2180 1049
rect 2166 1043 2172 1044
rect 2166 1039 2167 1043
rect 2171 1039 2172 1043
rect 2176 1039 2178 1048
rect 2224 1044 2226 1074
rect 2230 1053 2236 1054
rect 2230 1049 2231 1053
rect 2235 1049 2236 1053
rect 2230 1048 2236 1049
rect 2222 1043 2228 1044
rect 2222 1039 2223 1043
rect 2227 1039 2228 1043
rect 2232 1039 2234 1048
rect 1823 1038 1827 1039
rect 1823 1033 1827 1034
rect 1871 1038 1875 1039
rect 1871 1033 1875 1034
rect 1879 1038 1883 1039
rect 1879 1033 1883 1034
rect 1919 1038 1923 1039
rect 1919 1033 1923 1034
rect 1943 1038 1947 1039
rect 1943 1033 1947 1034
rect 1967 1038 1971 1039
rect 2002 1038 2008 1039
rect 2015 1038 2019 1039
rect 1967 1033 1971 1034
rect 2015 1033 2019 1034
rect 2063 1038 2067 1039
rect 2063 1033 2067 1034
rect 2095 1038 2099 1039
rect 2110 1038 2116 1039
rect 2119 1038 2123 1039
rect 2166 1038 2172 1039
rect 2175 1038 2179 1039
rect 2222 1038 2228 1039
rect 2231 1038 2235 1039
rect 2095 1033 2099 1034
rect 1814 1031 1820 1032
rect 1814 1027 1815 1031
rect 1819 1027 1820 1031
rect 1814 1026 1820 1027
rect 1824 1024 1826 1033
rect 1850 1031 1856 1032
rect 1850 1027 1851 1031
rect 1855 1027 1856 1031
rect 1850 1026 1856 1027
rect 1774 1023 1780 1024
rect 1774 1019 1775 1023
rect 1779 1019 1780 1023
rect 1774 1018 1780 1019
rect 1822 1023 1828 1024
rect 1822 1019 1823 1023
rect 1827 1019 1828 1023
rect 1822 1018 1828 1019
rect 1852 996 1854 1026
rect 1880 1024 1882 1033
rect 1906 1031 1912 1032
rect 1906 1027 1907 1031
rect 1911 1027 1912 1031
rect 1906 1026 1912 1027
rect 1878 1023 1884 1024
rect 1878 1019 1879 1023
rect 1883 1019 1884 1023
rect 1878 1018 1884 1019
rect 1908 996 1910 1026
rect 1944 1024 1946 1033
rect 2016 1024 2018 1033
rect 2096 1024 2098 1033
rect 1942 1023 1948 1024
rect 1942 1019 1943 1023
rect 1947 1019 1948 1023
rect 1942 1018 1948 1019
rect 2014 1023 2020 1024
rect 2014 1019 2015 1023
rect 2019 1019 2020 1023
rect 2014 1018 2020 1019
rect 2094 1023 2100 1024
rect 2094 1019 2095 1023
rect 2099 1019 2100 1023
rect 2094 1018 2100 1019
rect 2112 996 2114 1038
rect 2119 1033 2123 1034
rect 2175 1033 2179 1034
rect 2231 1033 2235 1034
rect 2126 1031 2132 1032
rect 2126 1027 2127 1031
rect 2131 1027 2132 1031
rect 2126 1026 2132 1027
rect 1278 995 1284 996
rect 1602 995 1608 996
rect 1238 991 1244 992
rect 1602 991 1603 995
rect 1607 991 1608 995
rect 1602 990 1608 991
rect 1642 995 1648 996
rect 1642 991 1643 995
rect 1647 991 1648 995
rect 1642 990 1648 991
rect 1682 995 1688 996
rect 1682 991 1683 995
rect 1687 991 1688 995
rect 1682 990 1688 991
rect 1718 995 1724 996
rect 1718 991 1719 995
rect 1723 991 1724 995
rect 1718 990 1724 991
rect 1762 995 1768 996
rect 1762 991 1763 995
rect 1767 991 1768 995
rect 1762 990 1768 991
rect 1850 995 1856 996
rect 1850 991 1851 995
rect 1855 991 1856 995
rect 1850 990 1856 991
rect 1906 995 1912 996
rect 1906 991 1907 995
rect 1911 991 1912 995
rect 1906 990 1912 991
rect 2110 995 2116 996
rect 2110 991 2111 995
rect 2115 991 2116 995
rect 2110 990 2116 991
rect 1686 987 1692 988
rect 1278 983 1284 984
rect 1238 979 1244 980
rect 1238 975 1239 979
rect 1243 975 1244 979
rect 1278 979 1279 983
rect 1283 979 1284 983
rect 1686 983 1687 987
rect 1691 983 1692 987
rect 1686 982 1692 983
rect 1278 978 1284 979
rect 1238 974 1244 975
rect 1240 967 1242 974
rect 1239 966 1243 967
rect 1280 963 1282 978
rect 1574 976 1580 977
rect 1574 972 1575 976
rect 1579 972 1580 976
rect 1574 971 1580 972
rect 1614 976 1620 977
rect 1614 972 1615 976
rect 1619 972 1620 976
rect 1614 971 1620 972
rect 1654 976 1660 977
rect 1654 972 1655 976
rect 1659 972 1660 976
rect 1654 971 1660 972
rect 1576 963 1578 971
rect 1616 963 1618 971
rect 1656 963 1658 971
rect 1239 961 1243 962
rect 1279 962 1283 963
rect 1240 954 1242 961
rect 1279 957 1283 958
rect 1303 962 1307 963
rect 1303 957 1307 958
rect 1351 962 1355 963
rect 1351 957 1355 958
rect 1431 962 1435 963
rect 1431 957 1435 958
rect 1511 962 1515 963
rect 1511 957 1515 958
rect 1575 962 1579 963
rect 1575 957 1579 958
rect 1591 962 1595 963
rect 1591 957 1595 958
rect 1615 962 1619 963
rect 1615 957 1619 958
rect 1655 962 1659 963
rect 1655 957 1659 958
rect 1679 962 1683 963
rect 1679 957 1683 958
rect 1238 953 1244 954
rect 1238 949 1239 953
rect 1243 949 1244 953
rect 1280 950 1282 957
rect 1302 956 1308 957
rect 1302 952 1303 956
rect 1307 952 1308 956
rect 1302 951 1308 952
rect 1350 956 1356 957
rect 1350 952 1351 956
rect 1355 952 1356 956
rect 1350 951 1356 952
rect 1430 956 1436 957
rect 1430 952 1431 956
rect 1435 952 1436 956
rect 1430 951 1436 952
rect 1510 956 1516 957
rect 1510 952 1511 956
rect 1515 952 1516 956
rect 1510 951 1516 952
rect 1590 956 1596 957
rect 1590 952 1591 956
rect 1595 952 1596 956
rect 1590 951 1596 952
rect 1678 956 1684 957
rect 1678 952 1679 956
rect 1683 952 1684 956
rect 1678 951 1684 952
rect 1238 948 1244 949
rect 1278 949 1284 950
rect 1278 945 1279 949
rect 1283 945 1284 949
rect 1278 944 1284 945
rect 1214 939 1220 940
rect 1214 935 1215 939
rect 1219 935 1220 939
rect 1214 934 1220 935
rect 1238 936 1244 937
rect 1238 932 1239 936
rect 1243 932 1244 936
rect 1286 935 1292 936
rect 1238 931 1244 932
rect 1278 932 1284 933
rect 1190 913 1196 914
rect 1190 909 1191 913
rect 1195 909 1196 913
rect 1190 908 1196 909
rect 1150 903 1156 904
rect 1150 899 1151 903
rect 1155 899 1156 903
rect 1150 898 1156 899
rect 1192 891 1194 908
rect 1240 891 1242 931
rect 1278 928 1279 932
rect 1283 928 1284 932
rect 1286 931 1287 935
rect 1291 931 1292 935
rect 1286 930 1292 931
rect 1646 935 1652 936
rect 1646 931 1647 935
rect 1651 931 1652 935
rect 1646 930 1652 931
rect 1278 927 1284 928
rect 1280 895 1282 927
rect 1288 904 1290 930
rect 1302 909 1308 910
rect 1302 905 1303 909
rect 1307 905 1308 909
rect 1302 904 1308 905
rect 1350 909 1356 910
rect 1350 905 1351 909
rect 1355 905 1356 909
rect 1350 904 1356 905
rect 1430 909 1436 910
rect 1430 905 1431 909
rect 1435 905 1436 909
rect 1430 904 1436 905
rect 1510 909 1516 910
rect 1510 905 1511 909
rect 1515 905 1516 909
rect 1510 904 1516 905
rect 1590 909 1596 910
rect 1590 905 1591 909
rect 1595 905 1596 909
rect 1590 904 1596 905
rect 1286 903 1292 904
rect 1286 899 1287 903
rect 1291 899 1292 903
rect 1286 898 1292 899
rect 1304 895 1306 904
rect 1352 895 1354 904
rect 1432 895 1434 904
rect 1512 895 1514 904
rect 1570 899 1576 900
rect 1570 895 1571 899
rect 1575 895 1576 899
rect 1592 895 1594 904
rect 1279 894 1283 895
rect 1023 890 1027 891
rect 1023 885 1027 886
rect 1071 890 1075 891
rect 1071 885 1075 886
rect 1087 890 1091 891
rect 1087 885 1091 886
rect 1143 890 1147 891
rect 1143 885 1147 886
rect 1159 890 1163 891
rect 1159 885 1163 886
rect 1191 890 1195 891
rect 1191 885 1195 886
rect 1239 890 1243 891
rect 1279 889 1283 890
rect 1303 894 1307 895
rect 1303 889 1307 890
rect 1351 894 1355 895
rect 1351 889 1355 890
rect 1431 894 1435 895
rect 1431 889 1435 890
rect 1439 894 1443 895
rect 1439 889 1443 890
rect 1479 894 1483 895
rect 1479 889 1483 890
rect 1511 894 1515 895
rect 1511 889 1515 890
rect 1519 894 1523 895
rect 1519 889 1523 890
rect 1559 894 1563 895
rect 1570 894 1576 895
rect 1591 894 1595 895
rect 1559 889 1563 890
rect 1239 885 1243 886
rect 1006 883 1012 884
rect 1006 879 1007 883
rect 1011 879 1012 883
rect 1006 878 1012 879
rect 1014 883 1020 884
rect 1014 879 1015 883
rect 1019 879 1020 883
rect 1014 878 1020 879
rect 958 875 964 876
rect 958 871 959 875
rect 963 871 964 875
rect 958 870 964 871
rect 1008 856 1010 878
rect 1024 876 1026 885
rect 1050 883 1056 884
rect 1050 879 1051 883
rect 1055 879 1056 883
rect 1050 878 1056 879
rect 1022 875 1028 876
rect 1022 871 1023 875
rect 1027 871 1028 875
rect 1022 870 1028 871
rect 1006 855 1012 856
rect 1006 851 1007 855
rect 1011 851 1012 855
rect 1006 850 1012 851
rect 1052 848 1054 878
rect 1088 876 1090 885
rect 1114 883 1120 884
rect 1114 879 1115 883
rect 1119 879 1120 883
rect 1114 878 1120 879
rect 1086 875 1092 876
rect 1086 871 1087 875
rect 1091 871 1092 875
rect 1086 870 1092 871
rect 1116 848 1118 878
rect 1160 876 1162 885
rect 1158 875 1164 876
rect 1158 871 1159 875
rect 1163 871 1164 875
rect 1158 870 1164 871
rect 1240 853 1242 885
rect 1280 857 1282 889
rect 1440 880 1442 889
rect 1454 887 1460 888
rect 1454 883 1455 887
rect 1459 883 1460 887
rect 1454 882 1460 883
rect 1462 887 1468 888
rect 1462 883 1463 887
rect 1467 883 1468 887
rect 1462 882 1468 883
rect 1438 879 1444 880
rect 1438 875 1439 879
rect 1443 875 1444 879
rect 1438 874 1444 875
rect 1278 856 1284 857
rect 1238 852 1244 853
rect 1238 848 1239 852
rect 1243 848 1244 852
rect 1278 852 1279 856
rect 1283 852 1284 856
rect 1278 851 1284 852
rect 386 847 392 848
rect 386 843 387 847
rect 391 843 392 847
rect 386 842 392 843
rect 498 847 504 848
rect 498 843 499 847
rect 503 843 504 847
rect 498 842 504 843
rect 602 847 608 848
rect 602 843 603 847
rect 607 843 608 847
rect 602 842 608 843
rect 662 847 668 848
rect 662 843 663 847
rect 667 843 668 847
rect 662 842 668 843
rect 754 847 760 848
rect 754 843 755 847
rect 759 843 760 847
rect 754 842 760 843
rect 870 847 876 848
rect 870 843 871 847
rect 875 843 876 847
rect 870 842 876 843
rect 946 847 952 848
rect 946 843 947 847
rect 951 843 952 847
rect 946 842 952 843
rect 1050 847 1056 848
rect 1050 843 1051 847
rect 1055 843 1056 847
rect 1050 842 1056 843
rect 1114 847 1120 848
rect 1238 847 1244 848
rect 1114 843 1115 847
rect 1119 843 1120 847
rect 1114 842 1120 843
rect 286 828 292 829
rect 286 824 287 828
rect 291 824 292 828
rect 286 823 292 824
rect 358 828 364 829
rect 358 824 359 828
rect 363 824 364 828
rect 358 823 364 824
rect 446 828 452 829
rect 446 824 447 828
rect 451 824 452 828
rect 446 823 452 824
rect 542 828 548 829
rect 542 824 543 828
rect 547 824 548 828
rect 542 823 548 824
rect 638 828 644 829
rect 638 824 639 828
rect 643 824 644 828
rect 638 823 644 824
rect 726 828 732 829
rect 726 824 727 828
rect 731 824 732 828
rect 726 823 732 824
rect 806 828 812 829
rect 806 824 807 828
rect 811 824 812 828
rect 806 823 812 824
rect 287 822 291 823
rect 287 817 291 818
rect 327 822 331 823
rect 327 817 331 818
rect 359 822 363 823
rect 359 817 363 818
rect 415 822 419 823
rect 415 817 419 818
rect 447 822 451 823
rect 447 817 451 818
rect 503 822 507 823
rect 503 817 507 818
rect 543 822 547 823
rect 543 817 547 818
rect 591 822 595 823
rect 591 817 595 818
rect 639 822 643 823
rect 639 817 643 818
rect 671 822 675 823
rect 671 817 675 818
rect 727 822 731 823
rect 727 817 731 818
rect 743 822 747 823
rect 743 817 747 818
rect 807 822 811 823
rect 807 817 811 818
rect 815 822 819 823
rect 815 817 819 818
rect 326 816 332 817
rect 326 812 327 816
rect 331 812 332 816
rect 326 811 332 812
rect 414 816 420 817
rect 414 812 415 816
rect 419 812 420 816
rect 414 811 420 812
rect 502 816 508 817
rect 502 812 503 816
rect 507 812 508 816
rect 502 811 508 812
rect 590 816 596 817
rect 590 812 591 816
rect 595 812 596 816
rect 590 811 596 812
rect 670 816 676 817
rect 670 812 671 816
rect 675 812 676 816
rect 670 811 676 812
rect 742 816 748 817
rect 742 812 743 816
rect 747 812 748 816
rect 742 811 748 812
rect 814 816 820 817
rect 814 812 815 816
rect 819 812 820 816
rect 814 811 820 812
rect 274 803 280 804
rect 274 799 275 803
rect 279 799 280 803
rect 274 798 280 799
rect 162 795 168 796
rect 110 792 116 793
rect 110 788 111 792
rect 115 788 116 792
rect 162 791 163 795
rect 167 791 168 795
rect 162 790 168 791
rect 230 795 236 796
rect 230 791 231 795
rect 235 791 236 795
rect 230 790 236 791
rect 318 795 324 796
rect 318 791 319 795
rect 323 791 324 795
rect 318 790 324 791
rect 406 795 412 796
rect 406 791 407 795
rect 411 791 412 795
rect 406 790 412 791
rect 494 795 500 796
rect 494 791 495 795
rect 499 791 500 795
rect 494 790 500 791
rect 662 795 668 796
rect 662 791 663 795
rect 667 791 668 795
rect 662 790 668 791
rect 734 795 740 796
rect 734 791 735 795
rect 739 791 740 795
rect 734 790 740 791
rect 806 795 812 796
rect 806 791 807 795
rect 811 791 812 795
rect 806 790 812 791
rect 110 787 116 788
rect 112 751 114 787
rect 134 769 140 770
rect 134 765 135 769
rect 139 765 140 769
rect 134 764 140 765
rect 136 751 138 764
rect 164 760 166 790
rect 174 769 180 770
rect 174 765 175 769
rect 179 765 180 769
rect 174 764 180 765
rect 154 759 160 760
rect 154 755 155 759
rect 159 755 160 759
rect 154 754 160 755
rect 162 759 168 760
rect 162 755 163 759
rect 167 755 168 759
rect 162 754 168 755
rect 111 750 115 751
rect 111 745 115 746
rect 135 750 139 751
rect 135 745 139 746
rect 112 713 114 745
rect 136 736 138 745
rect 134 735 140 736
rect 134 731 135 735
rect 139 731 140 735
rect 134 730 140 731
rect 110 712 116 713
rect 110 708 111 712
rect 115 708 116 712
rect 156 708 158 754
rect 176 751 178 764
rect 232 760 234 790
rect 238 769 244 770
rect 238 765 239 769
rect 243 765 244 769
rect 238 764 244 765
rect 230 759 236 760
rect 230 755 231 759
rect 235 755 236 759
rect 230 754 236 755
rect 240 751 242 764
rect 320 760 322 790
rect 326 769 332 770
rect 326 765 327 769
rect 331 765 332 769
rect 326 764 332 765
rect 318 759 324 760
rect 318 755 319 759
rect 323 755 324 759
rect 318 754 324 755
rect 328 751 330 764
rect 408 760 410 790
rect 414 769 420 770
rect 414 765 415 769
rect 419 765 420 769
rect 414 764 420 765
rect 406 759 412 760
rect 406 755 407 759
rect 411 755 412 759
rect 406 754 412 755
rect 416 751 418 764
rect 496 760 498 790
rect 606 787 612 788
rect 606 783 607 787
rect 611 783 612 787
rect 606 782 612 783
rect 502 769 508 770
rect 502 765 503 769
rect 507 765 508 769
rect 502 764 508 765
rect 590 769 596 770
rect 590 765 591 769
rect 595 765 596 769
rect 590 764 596 765
rect 494 759 500 760
rect 494 755 495 759
rect 499 755 500 759
rect 494 754 500 755
rect 504 751 506 764
rect 592 751 594 764
rect 608 760 610 782
rect 664 760 666 790
rect 670 769 676 770
rect 670 765 671 769
rect 675 765 676 769
rect 670 764 676 765
rect 606 759 612 760
rect 606 755 607 759
rect 611 755 612 759
rect 606 754 612 755
rect 662 759 668 760
rect 662 755 663 759
rect 667 755 668 759
rect 662 754 668 755
rect 672 751 674 764
rect 736 760 738 790
rect 742 769 748 770
rect 742 765 743 769
rect 747 765 748 769
rect 742 764 748 765
rect 734 759 740 760
rect 734 755 735 759
rect 739 755 740 759
rect 734 754 740 755
rect 744 751 746 764
rect 175 750 179 751
rect 175 745 179 746
rect 191 750 195 751
rect 191 745 195 746
rect 239 750 243 751
rect 239 745 243 746
rect 263 750 267 751
rect 263 745 267 746
rect 327 750 331 751
rect 327 745 331 746
rect 335 750 339 751
rect 335 745 339 746
rect 399 750 403 751
rect 399 745 403 746
rect 415 750 419 751
rect 415 745 419 746
rect 455 750 459 751
rect 455 745 459 746
rect 503 750 507 751
rect 503 745 507 746
rect 543 750 547 751
rect 543 745 547 746
rect 583 750 587 751
rect 583 745 587 746
rect 591 750 595 751
rect 591 745 595 746
rect 623 750 627 751
rect 623 745 627 746
rect 671 750 675 751
rect 671 745 675 746
rect 719 750 723 751
rect 719 745 723 746
rect 743 750 747 751
rect 743 745 747 746
rect 767 750 771 751
rect 767 745 771 746
rect 192 736 194 745
rect 222 743 228 744
rect 222 739 223 743
rect 227 739 228 743
rect 222 738 228 739
rect 190 735 196 736
rect 190 731 191 735
rect 195 731 196 735
rect 190 730 196 731
rect 110 707 116 708
rect 154 707 160 708
rect 154 703 155 707
rect 159 703 160 707
rect 154 702 160 703
rect 110 695 116 696
rect 110 691 111 695
rect 115 691 116 695
rect 110 690 116 691
rect 112 679 114 690
rect 134 688 140 689
rect 134 684 135 688
rect 139 684 140 688
rect 134 683 140 684
rect 190 688 196 689
rect 190 684 191 688
rect 195 684 196 688
rect 190 683 196 684
rect 136 679 138 683
rect 192 679 194 683
rect 111 678 115 679
rect 111 673 115 674
rect 135 678 139 679
rect 135 673 139 674
rect 191 678 195 679
rect 191 673 195 674
rect 199 678 203 679
rect 199 673 203 674
rect 112 666 114 673
rect 134 672 140 673
rect 134 668 135 672
rect 139 668 140 672
rect 134 667 140 668
rect 198 672 204 673
rect 198 668 199 672
rect 203 668 204 672
rect 198 667 204 668
rect 110 665 116 666
rect 110 661 111 665
rect 115 661 116 665
rect 110 660 116 661
rect 224 652 226 738
rect 264 736 266 745
rect 336 736 338 745
rect 386 743 392 744
rect 386 739 387 743
rect 391 739 392 743
rect 386 738 392 739
rect 262 735 268 736
rect 262 731 263 735
rect 267 731 268 735
rect 262 730 268 731
rect 334 735 340 736
rect 334 731 335 735
rect 339 731 340 735
rect 334 730 340 731
rect 388 708 390 738
rect 400 736 402 745
rect 442 743 448 744
rect 442 739 443 743
rect 447 739 448 743
rect 442 738 448 739
rect 398 735 404 736
rect 398 731 399 735
rect 403 731 404 735
rect 398 730 404 731
rect 444 708 446 738
rect 456 736 458 745
rect 490 743 496 744
rect 490 739 491 743
rect 495 739 496 743
rect 490 738 496 739
rect 454 735 460 736
rect 454 731 455 735
rect 459 731 460 735
rect 454 730 460 731
rect 492 708 494 738
rect 504 736 506 745
rect 530 743 536 744
rect 530 739 531 743
rect 535 739 536 743
rect 530 738 536 739
rect 502 735 508 736
rect 502 731 503 735
rect 507 731 508 735
rect 502 730 508 731
rect 532 715 534 738
rect 544 736 546 745
rect 570 743 576 744
rect 570 739 571 743
rect 575 739 576 743
rect 570 738 576 739
rect 542 735 548 736
rect 542 731 543 735
rect 547 731 548 735
rect 542 730 548 731
rect 572 715 574 738
rect 584 736 586 745
rect 610 743 616 744
rect 610 739 611 743
rect 615 739 616 743
rect 610 738 616 739
rect 582 735 588 736
rect 582 731 583 735
rect 587 731 588 735
rect 582 730 588 731
rect 612 715 614 738
rect 624 736 626 745
rect 658 743 664 744
rect 658 739 659 743
rect 663 739 664 743
rect 658 738 664 739
rect 622 735 628 736
rect 622 731 623 735
rect 627 731 628 735
rect 622 730 628 731
rect 532 713 542 715
rect 572 713 582 715
rect 612 713 622 715
rect 540 708 542 713
rect 580 708 582 713
rect 620 708 622 713
rect 286 707 292 708
rect 286 703 287 707
rect 291 703 292 707
rect 286 702 292 703
rect 386 707 392 708
rect 386 703 387 707
rect 391 703 392 707
rect 386 702 392 703
rect 442 707 448 708
rect 442 703 443 707
rect 447 703 448 707
rect 442 702 448 703
rect 490 707 496 708
rect 490 703 491 707
rect 495 703 496 707
rect 490 702 496 703
rect 538 707 544 708
rect 538 703 539 707
rect 543 703 544 707
rect 538 702 544 703
rect 578 707 584 708
rect 578 703 579 707
rect 583 703 584 707
rect 578 702 584 703
rect 618 707 624 708
rect 618 703 619 707
rect 623 703 624 707
rect 618 702 624 703
rect 262 688 268 689
rect 262 684 263 688
rect 267 684 268 688
rect 262 683 268 684
rect 264 679 266 683
rect 263 678 267 679
rect 263 673 267 674
rect 279 678 283 679
rect 279 673 283 674
rect 278 672 284 673
rect 278 668 279 672
rect 283 668 284 672
rect 278 667 284 668
rect 190 651 196 652
rect 110 648 116 649
rect 110 644 111 648
rect 115 644 116 648
rect 190 647 191 651
rect 195 647 196 651
rect 190 646 196 647
rect 222 651 228 652
rect 222 647 223 651
rect 227 647 228 651
rect 222 646 228 647
rect 110 643 116 644
rect 112 603 114 643
rect 134 625 140 626
rect 134 621 135 625
rect 139 621 140 625
rect 134 620 140 621
rect 136 603 138 620
rect 192 616 194 646
rect 198 625 204 626
rect 198 621 199 625
rect 203 621 204 625
rect 198 620 204 621
rect 278 625 284 626
rect 278 621 279 625
rect 283 621 284 625
rect 278 620 284 621
rect 158 615 164 616
rect 158 611 159 615
rect 163 611 164 615
rect 158 610 164 611
rect 190 615 196 616
rect 190 611 191 615
rect 195 611 196 615
rect 190 610 196 611
rect 111 602 115 603
rect 111 597 115 598
rect 135 602 139 603
rect 135 597 139 598
rect 112 565 114 597
rect 136 588 138 597
rect 134 587 140 588
rect 134 583 135 587
rect 139 583 140 587
rect 134 582 140 583
rect 110 564 116 565
rect 110 560 111 564
rect 115 560 116 564
rect 160 560 162 610
rect 200 603 202 620
rect 280 603 282 620
rect 288 616 290 702
rect 334 688 340 689
rect 334 684 335 688
rect 339 684 340 688
rect 334 683 340 684
rect 398 688 404 689
rect 398 684 399 688
rect 403 684 404 688
rect 398 683 404 684
rect 454 688 460 689
rect 454 684 455 688
rect 459 684 460 688
rect 454 683 460 684
rect 502 688 508 689
rect 502 684 503 688
rect 507 684 508 688
rect 502 683 508 684
rect 542 688 548 689
rect 542 684 543 688
rect 547 684 548 688
rect 542 683 548 684
rect 582 688 588 689
rect 582 684 583 688
rect 587 684 588 688
rect 582 683 588 684
rect 622 688 628 689
rect 622 684 623 688
rect 627 684 628 688
rect 622 683 628 684
rect 336 679 338 683
rect 400 679 402 683
rect 456 679 458 683
rect 504 679 506 683
rect 544 679 546 683
rect 584 679 586 683
rect 624 679 626 683
rect 335 678 339 679
rect 335 673 339 674
rect 351 678 355 679
rect 351 673 355 674
rect 399 678 403 679
rect 399 673 403 674
rect 415 678 419 679
rect 415 673 419 674
rect 455 678 459 679
rect 455 673 459 674
rect 487 678 491 679
rect 487 673 491 674
rect 503 678 507 679
rect 503 673 507 674
rect 543 678 547 679
rect 543 673 547 674
rect 559 678 563 679
rect 559 673 563 674
rect 583 678 587 679
rect 583 673 587 674
rect 623 678 627 679
rect 623 673 627 674
rect 639 678 643 679
rect 639 673 643 674
rect 350 672 356 673
rect 350 668 351 672
rect 355 668 356 672
rect 350 667 356 668
rect 414 672 420 673
rect 414 668 415 672
rect 419 668 420 672
rect 414 667 420 668
rect 486 672 492 673
rect 486 668 487 672
rect 491 668 492 672
rect 486 667 492 668
rect 558 672 564 673
rect 558 668 559 672
rect 563 668 564 672
rect 558 667 564 668
rect 638 672 644 673
rect 638 668 639 672
rect 643 668 644 672
rect 638 667 644 668
rect 660 652 662 738
rect 672 736 674 745
rect 698 743 704 744
rect 698 739 699 743
rect 703 739 704 743
rect 698 738 704 739
rect 706 743 712 744
rect 706 739 707 743
rect 711 739 712 743
rect 706 738 712 739
rect 670 735 676 736
rect 670 731 671 735
rect 675 731 676 735
rect 670 730 676 731
rect 700 720 702 738
rect 698 719 704 720
rect 698 715 699 719
rect 703 715 704 719
rect 698 714 704 715
rect 708 708 710 738
rect 720 736 722 745
rect 754 743 760 744
rect 754 739 755 743
rect 759 739 760 743
rect 754 738 760 739
rect 718 735 724 736
rect 718 731 719 735
rect 723 731 724 735
rect 718 730 724 731
rect 756 712 758 738
rect 768 736 770 745
rect 808 744 810 790
rect 822 787 828 788
rect 822 783 823 787
rect 827 783 828 787
rect 822 782 828 783
rect 814 769 820 770
rect 814 765 815 769
rect 819 765 820 769
rect 814 764 820 765
rect 816 751 818 764
rect 824 760 826 782
rect 872 760 874 842
rect 1278 839 1284 840
rect 1238 835 1244 836
rect 1238 831 1239 835
rect 1243 831 1244 835
rect 1278 835 1279 839
rect 1283 835 1284 839
rect 1278 834 1284 835
rect 1238 830 1244 831
rect 886 828 892 829
rect 886 824 887 828
rect 891 824 892 828
rect 886 823 892 824
rect 958 828 964 829
rect 958 824 959 828
rect 963 824 964 828
rect 958 823 964 824
rect 1022 828 1028 829
rect 1022 824 1023 828
rect 1027 824 1028 828
rect 1022 823 1028 824
rect 1086 828 1092 829
rect 1086 824 1087 828
rect 1091 824 1092 828
rect 1086 823 1092 824
rect 1158 828 1164 829
rect 1158 824 1159 828
rect 1163 824 1164 828
rect 1158 823 1164 824
rect 1240 823 1242 830
rect 879 822 883 823
rect 879 817 883 818
rect 887 822 891 823
rect 887 817 891 818
rect 943 822 947 823
rect 943 817 947 818
rect 959 822 963 823
rect 959 817 963 818
rect 1015 822 1019 823
rect 1015 817 1019 818
rect 1023 822 1027 823
rect 1023 817 1027 818
rect 1087 822 1091 823
rect 1087 817 1091 818
rect 1159 822 1163 823
rect 1159 817 1163 818
rect 1239 822 1243 823
rect 1239 817 1243 818
rect 878 816 884 817
rect 878 812 879 816
rect 883 812 884 816
rect 878 811 884 812
rect 942 816 948 817
rect 942 812 943 816
rect 947 812 948 816
rect 942 811 948 812
rect 1014 816 1020 817
rect 1014 812 1015 816
rect 1019 812 1020 816
rect 1014 811 1020 812
rect 1240 810 1242 817
rect 1280 815 1282 834
rect 1438 832 1444 833
rect 1438 828 1439 832
rect 1443 828 1444 832
rect 1438 827 1444 828
rect 1440 815 1442 827
rect 1279 814 1283 815
rect 1238 809 1244 810
rect 1279 809 1283 810
rect 1359 814 1363 815
rect 1359 809 1363 810
rect 1415 814 1419 815
rect 1415 809 1419 810
rect 1439 814 1443 815
rect 1439 809 1443 810
rect 1238 805 1239 809
rect 1243 805 1244 809
rect 1238 804 1244 805
rect 1280 802 1282 809
rect 1358 808 1364 809
rect 1358 804 1359 808
rect 1363 804 1364 808
rect 1358 803 1364 804
rect 1414 808 1420 809
rect 1414 804 1415 808
rect 1419 804 1420 808
rect 1414 803 1420 804
rect 1278 801 1284 802
rect 1278 797 1279 801
rect 1283 797 1284 801
rect 1278 796 1284 797
rect 1456 796 1458 882
rect 1464 852 1466 882
rect 1480 880 1482 889
rect 1502 887 1508 888
rect 1502 883 1503 887
rect 1507 883 1508 887
rect 1502 882 1508 883
rect 1478 879 1484 880
rect 1478 875 1479 879
rect 1483 875 1484 879
rect 1478 874 1484 875
rect 1504 852 1506 882
rect 1520 880 1522 889
rect 1546 887 1552 888
rect 1546 883 1547 887
rect 1551 883 1552 887
rect 1546 882 1552 883
rect 1518 879 1524 880
rect 1518 875 1519 879
rect 1523 875 1524 879
rect 1518 874 1524 875
rect 1548 852 1550 882
rect 1560 880 1562 889
rect 1558 879 1564 880
rect 1558 875 1559 879
rect 1563 875 1564 879
rect 1558 874 1564 875
rect 1572 860 1574 894
rect 1591 889 1595 890
rect 1607 894 1611 895
rect 1607 889 1611 890
rect 1608 880 1610 889
rect 1648 888 1650 930
rect 1678 909 1684 910
rect 1678 905 1679 909
rect 1683 905 1684 909
rect 1678 904 1684 905
rect 1680 895 1682 904
rect 1688 900 1690 982
rect 1694 976 1700 977
rect 1694 972 1695 976
rect 1699 972 1700 976
rect 1694 971 1700 972
rect 1734 976 1740 977
rect 1734 972 1735 976
rect 1739 972 1740 976
rect 1734 971 1740 972
rect 1774 976 1780 977
rect 1774 972 1775 976
rect 1779 972 1780 976
rect 1774 971 1780 972
rect 1822 976 1828 977
rect 1822 972 1823 976
rect 1827 972 1828 976
rect 1822 971 1828 972
rect 1878 976 1884 977
rect 1878 972 1879 976
rect 1883 972 1884 976
rect 1878 971 1884 972
rect 1942 976 1948 977
rect 1942 972 1943 976
rect 1947 972 1948 976
rect 1942 971 1948 972
rect 2014 976 2020 977
rect 2014 972 2015 976
rect 2019 972 2020 976
rect 2014 971 2020 972
rect 2094 976 2100 977
rect 2094 972 2095 976
rect 2099 972 2100 976
rect 2094 971 2100 972
rect 1696 963 1698 971
rect 1736 963 1738 971
rect 1776 963 1778 971
rect 1824 963 1826 971
rect 1880 963 1882 971
rect 1944 963 1946 971
rect 2016 963 2018 971
rect 2096 963 2098 971
rect 1695 962 1699 963
rect 1695 957 1699 958
rect 1735 962 1739 963
rect 1735 957 1739 958
rect 1767 962 1771 963
rect 1767 957 1771 958
rect 1775 962 1779 963
rect 1775 957 1779 958
rect 1823 962 1827 963
rect 1823 957 1827 958
rect 1855 962 1859 963
rect 1855 957 1859 958
rect 1879 962 1883 963
rect 1879 957 1883 958
rect 1943 962 1947 963
rect 1943 957 1947 958
rect 2015 962 2019 963
rect 2015 957 2019 958
rect 2023 962 2027 963
rect 2023 957 2027 958
rect 2095 962 2099 963
rect 2095 957 2099 958
rect 2103 962 2107 963
rect 2103 957 2107 958
rect 1766 956 1772 957
rect 1766 952 1767 956
rect 1771 952 1772 956
rect 1766 951 1772 952
rect 1854 956 1860 957
rect 1854 952 1855 956
rect 1859 952 1860 956
rect 1854 951 1860 952
rect 1942 956 1948 957
rect 1942 952 1943 956
rect 1947 952 1948 956
rect 1942 951 1948 952
rect 2022 956 2028 957
rect 2022 952 2023 956
rect 2027 952 2028 956
rect 2022 951 2028 952
rect 2102 956 2108 957
rect 2102 952 2103 956
rect 2107 952 2108 956
rect 2102 951 2108 952
rect 2128 936 2130 1026
rect 2176 1024 2178 1033
rect 2248 1032 2250 1074
rect 2406 1072 2407 1076
rect 2411 1072 2412 1076
rect 2406 1071 2412 1072
rect 2408 1039 2410 1071
rect 2255 1038 2259 1039
rect 2255 1033 2259 1034
rect 2407 1038 2411 1039
rect 2407 1033 2411 1034
rect 2238 1031 2244 1032
rect 2238 1027 2239 1031
rect 2243 1027 2244 1031
rect 2238 1026 2244 1027
rect 2246 1031 2252 1032
rect 2246 1027 2247 1031
rect 2251 1027 2252 1031
rect 2246 1026 2252 1027
rect 2174 1023 2180 1024
rect 2174 1019 2175 1023
rect 2179 1019 2180 1023
rect 2174 1018 2180 1019
rect 2240 996 2242 1026
rect 2256 1024 2258 1033
rect 2254 1023 2260 1024
rect 2254 1019 2255 1023
rect 2259 1019 2260 1023
rect 2254 1018 2260 1019
rect 2408 1001 2410 1033
rect 2406 1000 2412 1001
rect 2406 996 2407 1000
rect 2411 996 2412 1000
rect 2190 995 2196 996
rect 2190 991 2191 995
rect 2195 991 2196 995
rect 2190 990 2196 991
rect 2238 995 2244 996
rect 2406 995 2412 996
rect 2238 991 2239 995
rect 2243 991 2244 995
rect 2238 990 2244 991
rect 2174 976 2180 977
rect 2174 972 2175 976
rect 2179 972 2180 976
rect 2174 971 2180 972
rect 2176 963 2178 971
rect 2175 962 2179 963
rect 2175 957 2179 958
rect 2183 962 2187 963
rect 2183 957 2187 958
rect 2182 956 2188 957
rect 2182 952 2183 956
rect 2187 952 2188 956
rect 2182 951 2188 952
rect 1782 935 1788 936
rect 1782 931 1783 935
rect 1787 931 1788 935
rect 1782 930 1788 931
rect 2094 935 2100 936
rect 2094 931 2095 935
rect 2099 931 2100 935
rect 2094 930 2100 931
rect 2126 935 2132 936
rect 2126 931 2127 935
rect 2131 931 2132 935
rect 2126 930 2132 931
rect 1766 909 1772 910
rect 1766 905 1767 909
rect 1771 905 1772 909
rect 1766 904 1772 905
rect 1686 899 1692 900
rect 1686 895 1687 899
rect 1691 895 1692 899
rect 1768 895 1770 904
rect 1655 894 1659 895
rect 1655 889 1659 890
rect 1679 894 1683 895
rect 1686 894 1692 895
rect 1711 894 1715 895
rect 1679 889 1683 890
rect 1711 889 1715 890
rect 1767 894 1771 895
rect 1767 889 1771 890
rect 1775 894 1779 895
rect 1775 889 1779 890
rect 1646 887 1652 888
rect 1646 883 1647 887
rect 1651 883 1652 887
rect 1646 882 1652 883
rect 1656 880 1658 889
rect 1712 880 1714 889
rect 1776 880 1778 889
rect 1784 888 1786 930
rect 1854 909 1860 910
rect 1854 905 1855 909
rect 1859 905 1860 909
rect 1854 904 1860 905
rect 1942 909 1948 910
rect 1942 905 1943 909
rect 1947 905 1948 909
rect 1942 904 1948 905
rect 2022 909 2028 910
rect 2022 905 2023 909
rect 2027 905 2028 909
rect 2022 904 2028 905
rect 1856 895 1858 904
rect 1944 895 1946 904
rect 2024 895 2026 904
rect 2096 900 2098 930
rect 2102 909 2108 910
rect 2102 905 2103 909
rect 2107 905 2108 909
rect 2102 904 2108 905
rect 2182 909 2188 910
rect 2182 905 2183 909
rect 2187 905 2188 909
rect 2182 904 2188 905
rect 2086 899 2092 900
rect 2086 895 2087 899
rect 2091 895 2092 899
rect 1847 894 1851 895
rect 1847 889 1851 890
rect 1855 894 1859 895
rect 1855 889 1859 890
rect 1919 894 1923 895
rect 1919 889 1923 890
rect 1943 894 1947 895
rect 1943 889 1947 890
rect 1991 894 1995 895
rect 1991 889 1995 890
rect 2023 894 2027 895
rect 2023 889 2027 890
rect 2063 894 2067 895
rect 2086 894 2092 895
rect 2094 899 2100 900
rect 2094 895 2095 899
rect 2099 895 2100 899
rect 2104 895 2106 904
rect 2184 895 2186 904
rect 2192 900 2194 990
rect 2406 983 2412 984
rect 2406 979 2407 983
rect 2411 979 2412 983
rect 2406 978 2412 979
rect 2254 976 2260 977
rect 2254 972 2255 976
rect 2259 972 2260 976
rect 2254 971 2260 972
rect 2256 963 2258 971
rect 2408 963 2410 978
rect 2255 962 2259 963
rect 2255 957 2259 958
rect 2271 962 2275 963
rect 2271 957 2275 958
rect 2407 962 2411 963
rect 2407 957 2411 958
rect 2270 956 2276 957
rect 2270 952 2271 956
rect 2275 952 2276 956
rect 2270 951 2276 952
rect 2408 950 2410 957
rect 2406 949 2412 950
rect 2406 945 2407 949
rect 2411 945 2412 949
rect 2406 944 2412 945
rect 2262 935 2268 936
rect 2262 931 2263 935
rect 2267 931 2268 935
rect 2262 930 2268 931
rect 2286 935 2292 936
rect 2286 931 2287 935
rect 2291 931 2292 935
rect 2286 930 2292 931
rect 2406 932 2412 933
rect 2264 900 2266 930
rect 2270 909 2276 910
rect 2270 905 2271 909
rect 2275 905 2276 909
rect 2270 904 2276 905
rect 2190 899 2196 900
rect 2190 895 2191 899
rect 2195 895 2196 899
rect 2262 899 2268 900
rect 2262 895 2263 899
rect 2267 895 2268 899
rect 2272 895 2274 904
rect 2094 894 2100 895
rect 2103 894 2107 895
rect 2063 889 2067 890
rect 1782 887 1788 888
rect 1782 883 1783 887
rect 1787 883 1788 887
rect 1782 882 1788 883
rect 1802 887 1808 888
rect 1802 883 1803 887
rect 1807 883 1808 887
rect 1802 882 1808 883
rect 1606 879 1612 880
rect 1606 875 1607 879
rect 1611 875 1612 879
rect 1606 874 1612 875
rect 1654 879 1660 880
rect 1654 875 1655 879
rect 1659 875 1660 879
rect 1654 874 1660 875
rect 1710 879 1716 880
rect 1710 875 1711 879
rect 1715 875 1716 879
rect 1710 874 1716 875
rect 1774 879 1780 880
rect 1774 875 1775 879
rect 1779 875 1780 879
rect 1774 874 1780 875
rect 1570 859 1576 860
rect 1570 855 1571 859
rect 1575 855 1576 859
rect 1570 854 1576 855
rect 1804 852 1806 882
rect 1848 880 1850 889
rect 1874 887 1880 888
rect 1874 883 1875 887
rect 1879 883 1880 887
rect 1874 882 1880 883
rect 1846 879 1852 880
rect 1846 875 1847 879
rect 1851 875 1852 879
rect 1846 874 1852 875
rect 1876 852 1878 882
rect 1920 880 1922 889
rect 1992 880 1994 889
rect 2064 880 2066 889
rect 1918 879 1924 880
rect 1918 875 1919 879
rect 1923 875 1924 879
rect 1918 874 1924 875
rect 1990 879 1996 880
rect 1990 875 1991 879
rect 1995 875 1996 879
rect 1990 874 1996 875
rect 2062 879 2068 880
rect 2062 875 2063 879
rect 2067 875 2068 879
rect 2062 874 2068 875
rect 2088 852 2090 894
rect 2103 889 2107 890
rect 2135 894 2139 895
rect 2135 889 2139 890
rect 2183 894 2187 895
rect 2190 894 2196 895
rect 2215 894 2219 895
rect 2262 894 2268 895
rect 2271 894 2275 895
rect 2183 889 2187 890
rect 2215 889 2219 890
rect 2271 889 2275 890
rect 2110 887 2116 888
rect 2110 883 2111 887
rect 2115 883 2116 887
rect 2110 882 2116 883
rect 2112 852 2114 882
rect 2136 880 2138 889
rect 2202 887 2208 888
rect 2202 883 2203 887
rect 2207 883 2208 887
rect 2202 882 2208 883
rect 2134 879 2140 880
rect 2134 875 2135 879
rect 2139 875 2140 879
rect 2134 874 2140 875
rect 2204 852 2206 882
rect 2216 880 2218 889
rect 2288 888 2290 930
rect 2406 928 2407 932
rect 2411 928 2412 932
rect 2406 927 2412 928
rect 2408 895 2410 927
rect 2295 894 2299 895
rect 2295 889 2299 890
rect 2407 894 2411 895
rect 2407 889 2411 890
rect 2278 887 2284 888
rect 2278 883 2279 887
rect 2283 883 2284 887
rect 2278 882 2284 883
rect 2286 887 2292 888
rect 2286 883 2287 887
rect 2291 883 2292 887
rect 2286 882 2292 883
rect 2214 879 2220 880
rect 2214 875 2215 879
rect 2219 875 2220 879
rect 2214 874 2220 875
rect 2280 852 2282 882
rect 2296 880 2298 889
rect 2294 879 2300 880
rect 2294 875 2295 879
rect 2299 875 2300 879
rect 2294 874 2300 875
rect 2408 857 2410 889
rect 2406 856 2412 857
rect 2406 852 2407 856
rect 2411 852 2412 856
rect 1462 851 1468 852
rect 1462 847 1463 851
rect 1467 847 1468 851
rect 1462 846 1468 847
rect 1502 851 1508 852
rect 1502 847 1503 851
rect 1507 847 1508 851
rect 1502 846 1508 847
rect 1546 851 1552 852
rect 1546 847 1547 851
rect 1551 847 1552 851
rect 1546 846 1552 847
rect 1718 851 1724 852
rect 1718 847 1719 851
rect 1723 847 1724 851
rect 1718 846 1724 847
rect 1802 851 1808 852
rect 1802 847 1803 851
rect 1807 847 1808 851
rect 1802 846 1808 847
rect 1874 851 1880 852
rect 1874 847 1875 851
rect 1879 847 1880 851
rect 1874 846 1880 847
rect 2086 851 2092 852
rect 2086 847 2087 851
rect 2091 847 2092 851
rect 2086 846 2092 847
rect 2110 851 2116 852
rect 2110 847 2111 851
rect 2115 847 2116 851
rect 2110 846 2116 847
rect 2202 851 2208 852
rect 2202 847 2203 851
rect 2207 847 2208 851
rect 2202 846 2208 847
rect 2278 851 2284 852
rect 2406 851 2412 852
rect 2278 847 2279 851
rect 2283 847 2284 851
rect 2278 846 2284 847
rect 1478 832 1484 833
rect 1478 828 1479 832
rect 1483 828 1484 832
rect 1478 827 1484 828
rect 1518 832 1524 833
rect 1518 828 1519 832
rect 1523 828 1524 832
rect 1518 827 1524 828
rect 1558 832 1564 833
rect 1558 828 1559 832
rect 1563 828 1564 832
rect 1558 827 1564 828
rect 1606 832 1612 833
rect 1606 828 1607 832
rect 1611 828 1612 832
rect 1606 827 1612 828
rect 1654 832 1660 833
rect 1654 828 1655 832
rect 1659 828 1660 832
rect 1654 827 1660 828
rect 1710 832 1716 833
rect 1710 828 1711 832
rect 1715 828 1716 832
rect 1710 827 1716 828
rect 1480 815 1482 827
rect 1520 815 1522 827
rect 1560 815 1562 827
rect 1608 815 1610 827
rect 1656 815 1658 827
rect 1712 815 1714 827
rect 1471 814 1475 815
rect 1471 809 1475 810
rect 1479 814 1483 815
rect 1479 809 1483 810
rect 1519 814 1523 815
rect 1519 809 1523 810
rect 1535 814 1539 815
rect 1535 809 1539 810
rect 1559 814 1563 815
rect 1559 809 1563 810
rect 1591 814 1595 815
rect 1591 809 1595 810
rect 1607 814 1611 815
rect 1607 809 1611 810
rect 1647 814 1651 815
rect 1647 809 1651 810
rect 1655 814 1659 815
rect 1655 809 1659 810
rect 1703 814 1707 815
rect 1703 809 1707 810
rect 1711 814 1715 815
rect 1711 809 1715 810
rect 1470 808 1476 809
rect 1470 804 1471 808
rect 1475 804 1476 808
rect 1470 803 1476 804
rect 1534 808 1540 809
rect 1534 804 1535 808
rect 1539 804 1540 808
rect 1534 803 1540 804
rect 1590 808 1596 809
rect 1590 804 1591 808
rect 1595 804 1596 808
rect 1590 803 1596 804
rect 1646 808 1652 809
rect 1646 804 1647 808
rect 1651 804 1652 808
rect 1646 803 1652 804
rect 1702 808 1708 809
rect 1702 804 1703 808
rect 1707 804 1708 808
rect 1702 803 1708 804
rect 934 795 940 796
rect 934 791 935 795
rect 939 791 940 795
rect 934 790 940 791
rect 1006 795 1012 796
rect 1006 791 1007 795
rect 1011 791 1012 795
rect 1454 795 1460 796
rect 1006 790 1012 791
rect 1238 792 1244 793
rect 878 769 884 770
rect 878 765 879 769
rect 883 765 884 769
rect 878 764 884 765
rect 822 759 828 760
rect 822 755 823 759
rect 827 755 828 759
rect 822 754 828 755
rect 870 759 876 760
rect 870 755 871 759
rect 875 755 876 759
rect 870 754 876 755
rect 880 751 882 764
rect 936 760 938 790
rect 942 769 948 770
rect 942 765 943 769
rect 947 765 948 769
rect 942 764 948 765
rect 934 759 940 760
rect 934 755 935 759
rect 939 755 940 759
rect 934 754 940 755
rect 944 751 946 764
rect 1008 760 1010 790
rect 1238 788 1239 792
rect 1243 788 1244 792
rect 1454 791 1455 795
rect 1459 791 1460 795
rect 1454 790 1460 791
rect 1238 787 1244 788
rect 1398 787 1404 788
rect 1014 769 1020 770
rect 1014 765 1015 769
rect 1019 765 1020 769
rect 1014 764 1020 765
rect 1006 759 1012 760
rect 1006 755 1007 759
rect 1011 755 1012 759
rect 1006 754 1012 755
rect 1016 751 1018 764
rect 1240 751 1242 787
rect 1278 784 1284 785
rect 1278 780 1279 784
rect 1283 780 1284 784
rect 1398 783 1399 787
rect 1403 783 1404 787
rect 1398 782 1404 783
rect 1462 787 1468 788
rect 1462 783 1463 787
rect 1467 783 1468 787
rect 1462 782 1468 783
rect 1526 787 1532 788
rect 1526 783 1527 787
rect 1531 783 1532 787
rect 1526 782 1532 783
rect 1638 787 1644 788
rect 1638 783 1639 787
rect 1643 783 1644 787
rect 1638 782 1644 783
rect 1670 787 1676 788
rect 1670 783 1671 787
rect 1675 783 1676 787
rect 1670 782 1676 783
rect 1278 779 1284 780
rect 815 750 819 751
rect 815 745 819 746
rect 863 750 867 751
rect 863 745 867 746
rect 879 750 883 751
rect 879 745 883 746
rect 911 750 915 751
rect 911 745 915 746
rect 943 750 947 751
rect 943 745 947 746
rect 1015 750 1019 751
rect 1015 745 1019 746
rect 1239 750 1243 751
rect 1280 747 1282 779
rect 1358 761 1364 762
rect 1358 757 1359 761
rect 1363 757 1364 761
rect 1358 756 1364 757
rect 1360 747 1362 756
rect 1400 752 1402 782
rect 1414 761 1420 762
rect 1414 757 1415 761
rect 1419 757 1420 761
rect 1414 756 1420 757
rect 1390 751 1396 752
rect 1390 747 1391 751
rect 1395 747 1396 751
rect 1239 745 1243 746
rect 1279 746 1283 747
rect 806 743 812 744
rect 806 739 807 743
rect 811 739 812 743
rect 806 738 812 739
rect 816 736 818 745
rect 850 743 856 744
rect 850 739 851 743
rect 855 739 856 743
rect 850 738 856 739
rect 766 735 772 736
rect 766 731 767 735
rect 771 731 772 735
rect 766 730 772 731
rect 814 735 820 736
rect 814 731 815 735
rect 819 731 820 735
rect 814 730 820 731
rect 754 711 760 712
rect 706 707 712 708
rect 706 703 707 707
rect 711 703 712 707
rect 754 707 755 711
rect 759 707 760 711
rect 852 708 854 738
rect 864 736 866 745
rect 898 743 904 744
rect 898 739 899 743
rect 903 739 904 743
rect 898 738 904 739
rect 862 735 868 736
rect 862 731 863 735
rect 867 731 868 735
rect 862 730 868 731
rect 900 708 902 738
rect 912 736 914 745
rect 910 735 916 736
rect 910 731 911 735
rect 915 731 916 735
rect 910 730 916 731
rect 1240 713 1242 745
rect 1279 741 1283 742
rect 1303 746 1307 747
rect 1303 741 1307 742
rect 1343 746 1347 747
rect 1343 741 1347 742
rect 1359 746 1363 747
rect 1390 746 1396 747
rect 1398 751 1404 752
rect 1398 747 1399 751
rect 1403 747 1404 751
rect 1416 747 1418 756
rect 1464 752 1466 782
rect 1470 761 1476 762
rect 1470 757 1471 761
rect 1475 757 1476 761
rect 1470 756 1476 757
rect 1462 751 1468 752
rect 1462 747 1463 751
rect 1467 747 1468 751
rect 1472 747 1474 756
rect 1528 752 1530 782
rect 1598 779 1604 780
rect 1598 775 1599 779
rect 1603 775 1604 779
rect 1598 774 1604 775
rect 1534 761 1540 762
rect 1534 757 1535 761
rect 1539 757 1540 761
rect 1534 756 1540 757
rect 1590 761 1596 762
rect 1590 757 1591 761
rect 1595 757 1596 761
rect 1590 756 1596 757
rect 1526 751 1532 752
rect 1526 747 1527 751
rect 1531 747 1532 751
rect 1536 747 1538 756
rect 1592 747 1594 756
rect 1600 752 1602 774
rect 1640 752 1642 782
rect 1646 761 1652 762
rect 1646 757 1647 761
rect 1651 757 1652 761
rect 1646 756 1652 757
rect 1598 751 1604 752
rect 1598 747 1599 751
rect 1603 747 1604 751
rect 1398 746 1404 747
rect 1407 746 1411 747
rect 1359 741 1363 742
rect 1238 712 1244 713
rect 1238 708 1239 712
rect 1243 708 1244 712
rect 1280 709 1282 741
rect 1304 732 1306 741
rect 1322 739 1328 740
rect 1322 735 1323 739
rect 1327 735 1328 739
rect 1322 734 1328 735
rect 1330 739 1336 740
rect 1330 735 1331 739
rect 1335 735 1336 739
rect 1330 734 1336 735
rect 1302 731 1308 732
rect 1302 727 1303 731
rect 1307 727 1308 731
rect 1302 726 1308 727
rect 754 706 760 707
rect 790 707 796 708
rect 706 702 712 703
rect 790 703 791 707
rect 795 703 796 707
rect 790 702 796 703
rect 850 707 856 708
rect 850 703 851 707
rect 855 703 856 707
rect 850 702 856 703
rect 898 707 904 708
rect 1238 707 1244 708
rect 1278 708 1284 709
rect 898 703 899 707
rect 903 703 904 707
rect 1278 704 1279 708
rect 1283 704 1284 708
rect 1278 703 1284 704
rect 898 702 904 703
rect 670 688 676 689
rect 670 684 671 688
rect 675 684 676 688
rect 670 683 676 684
rect 718 688 724 689
rect 718 684 719 688
rect 723 684 724 688
rect 718 683 724 684
rect 766 688 772 689
rect 766 684 767 688
rect 771 684 772 688
rect 766 683 772 684
rect 672 679 674 683
rect 720 679 722 683
rect 768 679 770 683
rect 671 678 675 679
rect 671 673 675 674
rect 711 678 715 679
rect 711 673 715 674
rect 719 678 723 679
rect 719 673 723 674
rect 767 678 771 679
rect 767 673 771 674
rect 783 678 787 679
rect 783 673 787 674
rect 710 672 716 673
rect 710 668 711 672
rect 715 668 716 672
rect 710 667 716 668
rect 782 672 788 673
rect 782 668 783 672
rect 787 668 788 672
rect 782 667 788 668
rect 342 651 348 652
rect 342 647 343 651
rect 347 647 348 651
rect 342 646 348 647
rect 406 651 412 652
rect 406 647 407 651
rect 411 647 412 651
rect 406 646 412 647
rect 478 651 484 652
rect 478 647 479 651
rect 483 647 484 651
rect 478 646 484 647
rect 550 651 556 652
rect 550 647 551 651
rect 555 647 556 651
rect 550 646 556 647
rect 614 651 620 652
rect 614 647 615 651
rect 619 647 620 651
rect 614 646 620 647
rect 658 651 664 652
rect 658 647 659 651
rect 663 647 664 651
rect 658 646 664 647
rect 344 616 346 646
rect 350 625 356 626
rect 350 621 351 625
rect 355 621 356 625
rect 350 620 356 621
rect 286 615 292 616
rect 286 611 287 615
rect 291 611 292 615
rect 286 610 292 611
rect 342 615 348 616
rect 342 611 343 615
rect 347 611 348 615
rect 342 610 348 611
rect 352 603 354 620
rect 408 616 410 646
rect 414 625 420 626
rect 414 621 415 625
rect 419 621 420 625
rect 414 620 420 621
rect 406 615 412 616
rect 406 611 407 615
rect 411 611 412 615
rect 406 610 412 611
rect 416 603 418 620
rect 480 616 482 646
rect 486 625 492 626
rect 486 621 487 625
rect 491 621 492 625
rect 486 620 492 621
rect 478 615 484 616
rect 478 611 479 615
rect 483 611 484 615
rect 478 610 484 611
rect 488 603 490 620
rect 552 616 554 646
rect 558 625 564 626
rect 558 621 559 625
rect 563 621 564 625
rect 558 620 564 621
rect 550 615 556 616
rect 550 611 551 615
rect 555 611 556 615
rect 550 610 556 611
rect 560 603 562 620
rect 191 602 195 603
rect 191 597 195 598
rect 199 602 203 603
rect 199 597 203 598
rect 271 602 275 603
rect 271 597 275 598
rect 279 602 283 603
rect 279 597 283 598
rect 351 602 355 603
rect 351 597 355 598
rect 359 602 363 603
rect 359 597 363 598
rect 415 602 419 603
rect 415 597 419 598
rect 447 602 451 603
rect 447 597 451 598
rect 487 602 491 603
rect 487 597 491 598
rect 535 602 539 603
rect 535 597 539 598
rect 559 602 563 603
rect 559 597 563 598
rect 178 595 184 596
rect 178 591 179 595
rect 183 591 184 595
rect 178 590 184 591
rect 180 560 182 590
rect 192 588 194 597
rect 258 595 264 596
rect 258 591 259 595
rect 263 591 264 595
rect 258 590 264 591
rect 190 587 196 588
rect 190 583 191 587
rect 195 583 196 587
rect 190 582 196 583
rect 260 560 262 590
rect 272 588 274 597
rect 286 595 292 596
rect 286 591 287 595
rect 291 591 292 595
rect 286 590 292 591
rect 270 587 276 588
rect 270 583 271 587
rect 275 583 276 587
rect 270 582 276 583
rect 110 559 116 560
rect 158 559 164 560
rect 158 555 159 559
rect 163 555 164 559
rect 158 554 164 555
rect 178 559 184 560
rect 178 555 179 559
rect 183 555 184 559
rect 178 554 184 555
rect 258 559 264 560
rect 258 555 259 559
rect 263 555 264 559
rect 258 554 264 555
rect 110 547 116 548
rect 110 543 111 547
rect 115 543 116 547
rect 110 542 116 543
rect 112 527 114 542
rect 134 540 140 541
rect 134 536 135 540
rect 139 536 140 540
rect 134 535 140 536
rect 190 540 196 541
rect 190 536 191 540
rect 195 536 196 540
rect 190 535 196 536
rect 270 540 276 541
rect 270 536 271 540
rect 275 536 276 540
rect 270 535 276 536
rect 136 527 138 535
rect 192 527 194 535
rect 272 527 274 535
rect 111 526 115 527
rect 111 521 115 522
rect 135 526 139 527
rect 135 521 139 522
rect 191 526 195 527
rect 191 521 195 522
rect 263 526 267 527
rect 263 521 267 522
rect 271 526 275 527
rect 271 521 275 522
rect 112 514 114 521
rect 134 520 140 521
rect 134 516 135 520
rect 139 516 140 520
rect 134 515 140 516
rect 190 520 196 521
rect 190 516 191 520
rect 195 516 196 520
rect 190 515 196 516
rect 262 520 268 521
rect 262 516 263 520
rect 267 516 268 520
rect 262 515 268 516
rect 110 513 116 514
rect 110 509 111 513
rect 115 509 116 513
rect 110 508 116 509
rect 288 500 290 590
rect 360 588 362 597
rect 378 595 384 596
rect 378 591 379 595
rect 383 591 384 595
rect 378 590 384 591
rect 386 595 392 596
rect 386 591 387 595
rect 391 591 392 595
rect 386 590 392 591
rect 358 587 364 588
rect 358 583 359 587
rect 363 583 364 587
rect 358 582 364 583
rect 380 568 382 590
rect 378 567 384 568
rect 378 563 379 567
rect 383 563 384 567
rect 378 562 384 563
rect 388 560 390 590
rect 448 588 450 597
rect 474 595 480 596
rect 474 591 475 595
rect 479 591 480 595
rect 474 590 480 591
rect 446 587 452 588
rect 446 583 447 587
rect 451 583 452 587
rect 446 582 452 583
rect 476 560 478 590
rect 536 588 538 597
rect 616 596 618 646
rect 638 625 644 626
rect 638 621 639 625
rect 643 621 644 625
rect 638 620 644 621
rect 710 625 716 626
rect 710 621 711 625
rect 715 621 716 625
rect 710 620 716 621
rect 782 625 788 626
rect 782 621 783 625
rect 787 621 788 625
rect 782 620 788 621
rect 640 603 642 620
rect 712 603 714 620
rect 784 603 786 620
rect 792 616 794 702
rect 1238 695 1244 696
rect 1238 691 1239 695
rect 1243 691 1244 695
rect 1238 690 1244 691
rect 1278 691 1284 692
rect 814 688 820 689
rect 814 684 815 688
rect 819 684 820 688
rect 814 683 820 684
rect 862 688 868 689
rect 862 684 863 688
rect 867 684 868 688
rect 862 683 868 684
rect 910 688 916 689
rect 910 684 911 688
rect 915 684 916 688
rect 910 683 916 684
rect 816 679 818 683
rect 864 679 866 683
rect 912 679 914 683
rect 1240 679 1242 690
rect 1278 687 1279 691
rect 1283 687 1284 691
rect 1278 686 1284 687
rect 815 678 819 679
rect 815 673 819 674
rect 855 678 859 679
rect 855 673 859 674
rect 863 678 867 679
rect 863 673 867 674
rect 911 678 915 679
rect 911 673 915 674
rect 919 678 923 679
rect 919 673 923 674
rect 983 678 987 679
rect 983 673 987 674
rect 1039 678 1043 679
rect 1039 673 1043 674
rect 1095 678 1099 679
rect 1095 673 1099 674
rect 1151 678 1155 679
rect 1151 673 1155 674
rect 1191 678 1195 679
rect 1191 673 1195 674
rect 1239 678 1243 679
rect 1280 675 1282 686
rect 1302 684 1308 685
rect 1302 680 1303 684
rect 1307 680 1308 684
rect 1302 679 1308 680
rect 1304 675 1306 679
rect 1239 673 1243 674
rect 1279 674 1283 675
rect 854 672 860 673
rect 854 668 855 672
rect 859 668 860 672
rect 854 667 860 668
rect 918 672 924 673
rect 918 668 919 672
rect 923 668 924 672
rect 918 667 924 668
rect 982 672 988 673
rect 982 668 983 672
rect 987 668 988 672
rect 982 667 988 668
rect 1038 672 1044 673
rect 1038 668 1039 672
rect 1043 668 1044 672
rect 1038 667 1044 668
rect 1094 672 1100 673
rect 1094 668 1095 672
rect 1099 668 1100 672
rect 1094 667 1100 668
rect 1150 672 1156 673
rect 1150 668 1151 672
rect 1155 668 1156 672
rect 1150 667 1156 668
rect 1190 672 1196 673
rect 1190 668 1191 672
rect 1195 668 1196 672
rect 1190 667 1196 668
rect 1240 666 1242 673
rect 1279 669 1283 670
rect 1303 674 1307 675
rect 1303 669 1307 670
rect 1238 665 1244 666
rect 1238 661 1239 665
rect 1243 661 1244 665
rect 1280 662 1282 669
rect 1302 668 1308 669
rect 1302 664 1303 668
rect 1307 664 1308 668
rect 1302 663 1308 664
rect 1238 660 1244 661
rect 1278 661 1284 662
rect 1278 657 1279 661
rect 1283 657 1284 661
rect 1278 656 1284 657
rect 910 651 916 652
rect 910 647 911 651
rect 915 647 916 651
rect 910 646 916 647
rect 974 651 980 652
rect 974 647 975 651
rect 979 647 980 651
rect 974 646 980 647
rect 1022 651 1028 652
rect 1022 647 1023 651
rect 1027 647 1028 651
rect 1022 646 1028 647
rect 1086 651 1092 652
rect 1086 647 1087 651
rect 1091 647 1092 651
rect 1086 646 1092 647
rect 1142 651 1148 652
rect 1142 647 1143 651
rect 1147 647 1148 651
rect 1142 646 1148 647
rect 1178 651 1184 652
rect 1178 647 1179 651
rect 1183 647 1184 651
rect 1178 646 1184 647
rect 1230 651 1236 652
rect 1230 647 1231 651
rect 1235 647 1236 651
rect 1230 646 1236 647
rect 1238 648 1244 649
rect 1324 648 1326 734
rect 1332 704 1334 734
rect 1344 732 1346 741
rect 1370 739 1376 740
rect 1370 735 1371 739
rect 1375 735 1376 739
rect 1370 734 1376 735
rect 1342 731 1348 732
rect 1342 727 1343 731
rect 1347 727 1348 731
rect 1342 726 1348 727
rect 1372 704 1374 734
rect 1392 712 1394 746
rect 1407 741 1411 742
rect 1415 746 1419 747
rect 1462 746 1468 747
rect 1471 746 1475 747
rect 1415 741 1419 742
rect 1471 741 1475 742
rect 1487 746 1491 747
rect 1526 746 1532 747
rect 1535 746 1539 747
rect 1487 741 1491 742
rect 1535 741 1539 742
rect 1575 746 1579 747
rect 1575 741 1579 742
rect 1591 746 1595 747
rect 1598 746 1604 747
rect 1638 751 1644 752
rect 1638 747 1639 751
rect 1643 747 1644 751
rect 1648 747 1650 756
rect 1638 746 1644 747
rect 1647 746 1651 747
rect 1591 741 1595 742
rect 1647 741 1651 742
rect 1663 746 1667 747
rect 1663 741 1667 742
rect 1408 732 1410 741
rect 1434 739 1440 740
rect 1434 735 1435 739
rect 1439 735 1440 739
rect 1434 734 1440 735
rect 1406 731 1412 732
rect 1406 727 1407 731
rect 1411 727 1412 731
rect 1406 726 1412 727
rect 1390 711 1396 712
rect 1390 707 1391 711
rect 1395 707 1396 711
rect 1390 706 1396 707
rect 1436 704 1438 734
rect 1488 732 1490 741
rect 1514 739 1520 740
rect 1514 735 1515 739
rect 1519 735 1520 739
rect 1514 734 1520 735
rect 1486 731 1492 732
rect 1486 727 1487 731
rect 1491 727 1492 731
rect 1486 726 1492 727
rect 1516 704 1518 734
rect 1576 732 1578 741
rect 1664 732 1666 741
rect 1672 740 1674 782
rect 1702 761 1708 762
rect 1702 757 1703 761
rect 1707 757 1708 761
rect 1702 756 1708 757
rect 1704 747 1706 756
rect 1720 752 1722 846
rect 1766 843 1772 844
rect 1766 839 1767 843
rect 1771 839 1772 843
rect 1766 838 1772 839
rect 2406 839 2412 840
rect 1759 814 1763 815
rect 1759 809 1763 810
rect 1758 808 1764 809
rect 1758 804 1759 808
rect 1763 804 1764 808
rect 1758 803 1764 804
rect 1758 761 1764 762
rect 1758 757 1759 761
rect 1763 757 1764 761
rect 1758 756 1764 757
rect 1718 751 1724 752
rect 1718 747 1719 751
rect 1723 747 1724 751
rect 1760 747 1762 756
rect 1768 752 1770 838
rect 2406 835 2407 839
rect 2411 835 2412 839
rect 2406 834 2412 835
rect 1774 832 1780 833
rect 1774 828 1775 832
rect 1779 828 1780 832
rect 1774 827 1780 828
rect 1846 832 1852 833
rect 1846 828 1847 832
rect 1851 828 1852 832
rect 1846 827 1852 828
rect 1918 832 1924 833
rect 1918 828 1919 832
rect 1923 828 1924 832
rect 1918 827 1924 828
rect 1990 832 1996 833
rect 1990 828 1991 832
rect 1995 828 1996 832
rect 1990 827 1996 828
rect 2062 832 2068 833
rect 2062 828 2063 832
rect 2067 828 2068 832
rect 2062 827 2068 828
rect 2134 832 2140 833
rect 2134 828 2135 832
rect 2139 828 2140 832
rect 2134 827 2140 828
rect 2214 832 2220 833
rect 2214 828 2215 832
rect 2219 828 2220 832
rect 2214 827 2220 828
rect 2294 832 2300 833
rect 2294 828 2295 832
rect 2299 828 2300 832
rect 2294 827 2300 828
rect 1776 815 1778 827
rect 1848 815 1850 827
rect 1920 815 1922 827
rect 1992 815 1994 827
rect 2064 815 2066 827
rect 2136 815 2138 827
rect 2216 815 2218 827
rect 2296 815 2298 827
rect 2408 815 2410 834
rect 1775 814 1779 815
rect 1775 809 1779 810
rect 1815 814 1819 815
rect 1815 809 1819 810
rect 1847 814 1851 815
rect 1847 809 1851 810
rect 1871 814 1875 815
rect 1871 809 1875 810
rect 1919 814 1923 815
rect 1919 809 1923 810
rect 1935 814 1939 815
rect 1935 809 1939 810
rect 1991 814 1995 815
rect 1991 809 1995 810
rect 1999 814 2003 815
rect 1999 809 2003 810
rect 2063 814 2067 815
rect 2063 809 2067 810
rect 2071 814 2075 815
rect 2071 809 2075 810
rect 2135 814 2139 815
rect 2135 809 2139 810
rect 2143 814 2147 815
rect 2143 809 2147 810
rect 2215 814 2219 815
rect 2215 809 2219 810
rect 2223 814 2227 815
rect 2223 809 2227 810
rect 2295 814 2299 815
rect 2295 809 2299 810
rect 2303 814 2307 815
rect 2303 809 2307 810
rect 2359 814 2363 815
rect 2359 809 2363 810
rect 2407 814 2411 815
rect 2407 809 2411 810
rect 1814 808 1820 809
rect 1814 804 1815 808
rect 1819 804 1820 808
rect 1814 803 1820 804
rect 1870 808 1876 809
rect 1870 804 1871 808
rect 1875 804 1876 808
rect 1870 803 1876 804
rect 1934 808 1940 809
rect 1934 804 1935 808
rect 1939 804 1940 808
rect 1934 803 1940 804
rect 1998 808 2004 809
rect 1998 804 1999 808
rect 2003 804 2004 808
rect 1998 803 2004 804
rect 2070 808 2076 809
rect 2070 804 2071 808
rect 2075 804 2076 808
rect 2070 803 2076 804
rect 2142 808 2148 809
rect 2142 804 2143 808
rect 2147 804 2148 808
rect 2142 803 2148 804
rect 2222 808 2228 809
rect 2222 804 2223 808
rect 2227 804 2228 808
rect 2222 803 2228 804
rect 2302 808 2308 809
rect 2302 804 2303 808
rect 2307 804 2308 808
rect 2302 803 2308 804
rect 2358 808 2364 809
rect 2358 804 2359 808
rect 2363 804 2364 808
rect 2358 803 2364 804
rect 2408 802 2410 809
rect 2406 801 2412 802
rect 2406 797 2407 801
rect 2411 797 2412 801
rect 2406 796 2412 797
rect 1798 787 1804 788
rect 1798 783 1799 787
rect 1803 783 1804 787
rect 1798 782 1804 783
rect 1862 787 1868 788
rect 1862 783 1863 787
rect 1867 783 1868 787
rect 1862 782 1868 783
rect 1926 787 1932 788
rect 1926 783 1927 787
rect 1931 783 1932 787
rect 1926 782 1932 783
rect 1982 787 1988 788
rect 1982 783 1983 787
rect 1987 783 1988 787
rect 1982 782 1988 783
rect 2062 787 2068 788
rect 2062 783 2063 787
rect 2067 783 2068 787
rect 2062 782 2068 783
rect 2134 787 2140 788
rect 2134 783 2135 787
rect 2139 783 2140 787
rect 2134 782 2140 783
rect 2150 787 2156 788
rect 2150 783 2151 787
rect 2155 783 2156 787
rect 2150 782 2156 783
rect 2294 787 2300 788
rect 2294 783 2295 787
rect 2299 783 2300 787
rect 2294 782 2300 783
rect 2350 787 2356 788
rect 2350 783 2351 787
rect 2355 783 2356 787
rect 2350 782 2356 783
rect 2370 787 2376 788
rect 2370 783 2371 787
rect 2375 783 2376 787
rect 2370 782 2376 783
rect 2406 784 2412 785
rect 1800 752 1802 782
rect 1839 764 1843 765
rect 1814 761 1820 762
rect 1814 757 1815 761
rect 1819 757 1820 761
rect 1839 759 1843 760
rect 1814 756 1820 757
rect 1766 751 1772 752
rect 1766 747 1767 751
rect 1771 747 1772 751
rect 1703 746 1707 747
rect 1718 746 1724 747
rect 1751 746 1755 747
rect 1703 741 1707 742
rect 1751 741 1755 742
rect 1759 746 1763 747
rect 1766 746 1772 747
rect 1798 751 1804 752
rect 1798 747 1799 751
rect 1803 747 1804 751
rect 1816 747 1818 756
rect 1798 746 1804 747
rect 1815 746 1819 747
rect 1759 741 1763 742
rect 1815 741 1819 742
rect 1831 746 1835 747
rect 1831 741 1835 742
rect 1670 739 1676 740
rect 1670 735 1671 739
rect 1675 735 1676 739
rect 1670 734 1676 735
rect 1690 739 1696 740
rect 1690 735 1691 739
rect 1695 735 1696 739
rect 1690 734 1696 735
rect 1574 731 1580 732
rect 1574 727 1575 731
rect 1579 727 1580 731
rect 1574 726 1580 727
rect 1662 731 1668 732
rect 1662 727 1663 731
rect 1667 727 1668 731
rect 1662 726 1668 727
rect 1692 704 1694 734
rect 1752 732 1754 741
rect 1832 732 1834 741
rect 1840 740 1842 759
rect 1864 752 1866 782
rect 1870 761 1876 762
rect 1870 757 1871 761
rect 1875 757 1876 761
rect 1870 756 1876 757
rect 1862 751 1868 752
rect 1862 747 1863 751
rect 1867 747 1868 751
rect 1872 747 1874 756
rect 1928 752 1930 782
rect 1934 761 1940 762
rect 1934 757 1935 761
rect 1939 757 1940 761
rect 1934 756 1940 757
rect 1926 751 1932 752
rect 1926 747 1927 751
rect 1931 747 1932 751
rect 1936 747 1938 756
rect 1984 752 1986 782
rect 1998 761 2004 762
rect 1998 757 1999 761
rect 2003 757 2004 761
rect 1998 756 2004 757
rect 1982 751 1988 752
rect 1982 747 1983 751
rect 1987 747 1988 751
rect 2000 747 2002 756
rect 2064 752 2066 782
rect 2070 761 2076 762
rect 2070 757 2071 761
rect 2075 757 2076 761
rect 2070 756 2076 757
rect 2062 751 2068 752
rect 2062 747 2063 751
rect 2067 747 2068 751
rect 2072 747 2074 756
rect 2136 752 2138 782
rect 2152 765 2154 782
rect 2151 764 2155 765
rect 2142 761 2148 762
rect 2142 757 2143 761
rect 2147 757 2148 761
rect 2151 759 2155 760
rect 2222 761 2228 762
rect 2142 756 2148 757
rect 2222 757 2223 761
rect 2227 757 2228 761
rect 2222 756 2228 757
rect 2134 751 2140 752
rect 2134 747 2135 751
rect 2139 747 2140 751
rect 2144 747 2146 756
rect 2224 747 2226 756
rect 2296 752 2298 782
rect 2302 761 2308 762
rect 2302 757 2303 761
rect 2307 757 2308 761
rect 2302 756 2308 757
rect 2286 751 2292 752
rect 2286 747 2287 751
rect 2291 747 2292 751
rect 1862 746 1868 747
rect 1871 746 1875 747
rect 1871 741 1875 742
rect 1911 746 1915 747
rect 1926 746 1932 747
rect 1935 746 1939 747
rect 1982 746 1988 747
rect 1991 746 1995 747
rect 1911 741 1915 742
rect 1935 741 1939 742
rect 1991 741 1995 742
rect 1999 746 2003 747
rect 2062 746 2068 747
rect 2071 746 2075 747
rect 1999 741 2003 742
rect 2071 741 2075 742
rect 2079 746 2083 747
rect 2134 746 2140 747
rect 2143 746 2147 747
rect 2079 741 2083 742
rect 2143 741 2147 742
rect 2175 746 2179 747
rect 2175 741 2179 742
rect 2223 746 2227 747
rect 2223 741 2227 742
rect 2279 746 2283 747
rect 2286 746 2292 747
rect 2294 751 2300 752
rect 2294 747 2295 751
rect 2299 747 2300 751
rect 2304 747 2306 756
rect 2352 752 2354 782
rect 2358 761 2364 762
rect 2358 757 2359 761
rect 2363 757 2364 761
rect 2358 756 2364 757
rect 2350 751 2356 752
rect 2350 747 2351 751
rect 2355 747 2356 751
rect 2360 747 2362 756
rect 2294 746 2300 747
rect 2303 746 2307 747
rect 2350 746 2356 747
rect 2359 746 2363 747
rect 2279 741 2283 742
rect 1838 739 1844 740
rect 1838 735 1839 739
rect 1843 735 1844 739
rect 1838 734 1844 735
rect 1858 739 1864 740
rect 1858 735 1859 739
rect 1863 735 1864 739
rect 1858 734 1864 735
rect 1750 731 1756 732
rect 1750 727 1751 731
rect 1755 727 1756 731
rect 1750 726 1756 727
rect 1830 731 1836 732
rect 1830 727 1831 731
rect 1835 727 1836 731
rect 1830 726 1836 727
rect 1860 704 1862 734
rect 1912 732 1914 741
rect 1934 735 1940 736
rect 1910 731 1916 732
rect 1910 727 1911 731
rect 1915 727 1916 731
rect 1934 731 1935 735
rect 1939 731 1940 735
rect 1992 732 1994 741
rect 2018 739 2024 740
rect 2018 735 2019 739
rect 2023 735 2024 739
rect 2018 734 2024 735
rect 1934 730 1940 731
rect 1990 731 1996 732
rect 1910 726 1916 727
rect 1936 704 1938 730
rect 1990 727 1991 731
rect 1995 727 1996 731
rect 1990 726 1996 727
rect 2020 704 2022 734
rect 2080 732 2082 741
rect 2106 739 2112 740
rect 2106 735 2107 739
rect 2111 735 2112 739
rect 2106 734 2112 735
rect 2078 731 2084 732
rect 2078 727 2079 731
rect 2083 727 2084 731
rect 2078 726 2084 727
rect 2108 704 2110 734
rect 2176 732 2178 741
rect 2202 739 2208 740
rect 2202 735 2203 739
rect 2207 735 2208 739
rect 2202 734 2208 735
rect 2174 731 2180 732
rect 2174 727 2175 731
rect 2179 727 2180 731
rect 2174 726 2180 727
rect 2204 704 2206 734
rect 2280 732 2282 741
rect 2278 731 2284 732
rect 2278 727 2279 731
rect 2283 727 2284 731
rect 2278 726 2284 727
rect 1330 703 1336 704
rect 1330 699 1331 703
rect 1335 699 1336 703
rect 1330 698 1336 699
rect 1370 703 1376 704
rect 1370 699 1371 703
rect 1375 699 1376 703
rect 1370 698 1376 699
rect 1434 703 1440 704
rect 1434 699 1435 703
rect 1439 699 1440 703
rect 1434 698 1440 699
rect 1514 703 1520 704
rect 1514 699 1515 703
rect 1519 699 1520 703
rect 1514 698 1520 699
rect 1690 703 1696 704
rect 1690 699 1691 703
rect 1695 699 1696 703
rect 1690 698 1696 699
rect 1734 703 1740 704
rect 1734 699 1735 703
rect 1739 699 1740 703
rect 1734 698 1740 699
rect 1858 703 1864 704
rect 1858 699 1859 703
rect 1863 699 1864 703
rect 1858 698 1864 699
rect 1934 703 1940 704
rect 1934 699 1935 703
rect 1939 699 1940 703
rect 1934 698 1940 699
rect 2018 703 2024 704
rect 2018 699 2019 703
rect 2023 699 2024 703
rect 2018 698 2024 699
rect 2106 703 2112 704
rect 2106 699 2107 703
rect 2111 699 2112 703
rect 2106 698 2112 699
rect 2202 703 2208 704
rect 2202 699 2203 703
rect 2207 699 2208 703
rect 2202 698 2208 699
rect 2246 703 2252 704
rect 2246 699 2247 703
rect 2251 699 2252 703
rect 2246 698 2252 699
rect 1342 684 1348 685
rect 1342 680 1343 684
rect 1347 680 1348 684
rect 1342 679 1348 680
rect 1406 684 1412 685
rect 1406 680 1407 684
rect 1411 680 1412 684
rect 1406 679 1412 680
rect 1486 684 1492 685
rect 1486 680 1487 684
rect 1491 680 1492 684
rect 1486 679 1492 680
rect 1574 684 1580 685
rect 1574 680 1575 684
rect 1579 680 1580 684
rect 1574 679 1580 680
rect 1662 684 1668 685
rect 1662 680 1663 684
rect 1667 680 1668 684
rect 1662 679 1668 680
rect 1344 675 1346 679
rect 1408 675 1410 679
rect 1488 675 1490 679
rect 1576 675 1578 679
rect 1664 675 1666 679
rect 1343 674 1347 675
rect 1343 669 1347 670
rect 1399 674 1403 675
rect 1399 669 1403 670
rect 1407 674 1411 675
rect 1407 669 1411 670
rect 1487 674 1491 675
rect 1487 669 1491 670
rect 1511 674 1515 675
rect 1511 669 1515 670
rect 1575 674 1579 675
rect 1575 669 1579 670
rect 1623 674 1627 675
rect 1623 669 1627 670
rect 1663 674 1667 675
rect 1663 669 1667 670
rect 1727 674 1731 675
rect 1727 669 1731 670
rect 1398 668 1404 669
rect 1398 664 1399 668
rect 1403 664 1404 668
rect 1398 663 1404 664
rect 1510 668 1516 669
rect 1510 664 1511 668
rect 1515 664 1516 668
rect 1510 663 1516 664
rect 1622 668 1628 669
rect 1622 664 1623 668
rect 1627 664 1628 668
rect 1622 663 1628 664
rect 1726 668 1732 669
rect 1726 664 1727 668
rect 1731 664 1732 668
rect 1726 663 1732 664
rect 854 625 860 626
rect 854 621 855 625
rect 859 621 860 625
rect 854 620 860 621
rect 790 615 796 616
rect 790 611 791 615
rect 795 611 796 615
rect 790 610 796 611
rect 856 603 858 620
rect 912 616 914 646
rect 918 625 924 626
rect 918 621 919 625
rect 923 621 924 625
rect 918 620 924 621
rect 902 615 908 616
rect 902 611 903 615
rect 907 611 908 615
rect 902 610 908 611
rect 910 615 916 616
rect 910 611 911 615
rect 915 611 916 615
rect 910 610 916 611
rect 623 602 627 603
rect 623 597 627 598
rect 639 602 643 603
rect 639 597 643 598
rect 703 602 707 603
rect 703 597 707 598
rect 711 602 715 603
rect 711 597 715 598
rect 783 602 787 603
rect 783 597 787 598
rect 855 602 859 603
rect 855 597 859 598
rect 614 595 620 596
rect 614 591 615 595
rect 619 591 620 595
rect 614 590 620 591
rect 624 588 626 597
rect 650 595 656 596
rect 650 591 651 595
rect 655 591 656 595
rect 650 590 656 591
rect 534 587 540 588
rect 534 583 535 587
rect 539 583 540 587
rect 534 582 540 583
rect 622 587 628 588
rect 622 583 623 587
rect 627 583 628 587
rect 622 582 628 583
rect 652 560 654 590
rect 704 588 706 597
rect 784 588 786 597
rect 802 595 808 596
rect 802 591 803 595
rect 807 591 808 595
rect 802 590 808 591
rect 810 595 816 596
rect 810 591 811 595
rect 815 591 816 595
rect 810 590 816 591
rect 702 587 708 588
rect 702 583 703 587
rect 707 583 708 587
rect 702 582 708 583
rect 782 587 788 588
rect 782 583 783 587
rect 787 583 788 587
rect 782 582 788 583
rect 386 559 392 560
rect 386 555 387 559
rect 391 555 392 559
rect 386 554 392 555
rect 474 559 480 560
rect 474 555 475 559
rect 479 555 480 559
rect 474 554 480 555
rect 562 559 568 560
rect 562 555 563 559
rect 567 555 568 559
rect 562 554 568 555
rect 650 559 656 560
rect 650 555 651 559
rect 655 555 656 559
rect 650 554 656 555
rect 358 540 364 541
rect 358 536 359 540
rect 363 536 364 540
rect 358 535 364 536
rect 446 540 452 541
rect 446 536 447 540
rect 451 536 452 540
rect 446 535 452 536
rect 534 540 540 541
rect 534 536 535 540
rect 539 536 540 540
rect 534 535 540 536
rect 360 527 362 535
rect 448 527 450 535
rect 536 527 538 535
rect 335 526 339 527
rect 335 521 339 522
rect 359 526 363 527
rect 359 521 363 522
rect 415 526 419 527
rect 415 521 419 522
rect 447 526 451 527
rect 447 521 451 522
rect 495 526 499 527
rect 495 521 499 522
rect 535 526 539 527
rect 535 521 539 522
rect 334 520 340 521
rect 334 516 335 520
rect 339 516 340 520
rect 334 515 340 516
rect 414 520 420 521
rect 414 516 415 520
rect 419 516 420 520
rect 414 515 420 516
rect 494 520 500 521
rect 494 516 495 520
rect 499 516 500 520
rect 494 515 500 516
rect 254 499 260 500
rect 110 496 116 497
rect 110 492 111 496
rect 115 492 116 496
rect 254 495 255 499
rect 259 495 260 499
rect 254 494 260 495
rect 286 499 292 500
rect 286 495 287 499
rect 291 495 292 499
rect 286 494 292 495
rect 342 499 348 500
rect 342 495 343 499
rect 347 495 348 499
rect 342 494 348 495
rect 110 491 116 492
rect 112 459 114 491
rect 134 473 140 474
rect 134 469 135 473
rect 139 469 140 473
rect 134 468 140 469
rect 190 473 196 474
rect 190 469 191 473
rect 195 469 196 473
rect 190 468 196 469
rect 136 459 138 468
rect 192 459 194 468
rect 256 464 258 494
rect 262 473 268 474
rect 262 469 263 473
rect 267 469 268 473
rect 262 468 268 469
rect 334 473 340 474
rect 334 469 335 473
rect 339 469 340 473
rect 334 468 340 469
rect 254 463 260 464
rect 254 459 255 463
rect 259 459 260 463
rect 264 459 266 468
rect 336 459 338 468
rect 111 458 115 459
rect 111 453 115 454
rect 135 458 139 459
rect 135 453 139 454
rect 183 458 187 459
rect 183 453 187 454
rect 191 458 195 459
rect 191 453 195 454
rect 223 458 227 459
rect 254 458 260 459
rect 263 458 267 459
rect 223 453 227 454
rect 263 453 267 454
rect 311 458 315 459
rect 311 453 315 454
rect 335 458 339 459
rect 335 453 339 454
rect 112 421 114 453
rect 184 444 186 453
rect 210 451 216 452
rect 210 447 211 451
rect 215 447 216 451
rect 210 446 216 447
rect 182 443 188 444
rect 182 439 183 443
rect 187 439 188 443
rect 182 438 188 439
rect 110 420 116 421
rect 110 416 111 420
rect 115 416 116 420
rect 110 415 116 416
rect 212 414 214 446
rect 224 444 226 453
rect 250 451 256 452
rect 250 447 251 451
rect 255 447 256 451
rect 250 446 256 447
rect 222 443 228 444
rect 222 439 223 443
rect 227 439 228 443
rect 222 438 228 439
rect 218 415 224 416
rect 218 414 219 415
rect 212 412 219 414
rect 218 411 219 412
rect 223 411 224 415
rect 252 414 254 446
rect 264 444 266 453
rect 298 451 304 452
rect 298 447 299 451
rect 303 447 304 451
rect 298 446 304 447
rect 262 443 268 444
rect 262 439 263 443
rect 267 439 268 443
rect 262 438 268 439
rect 258 415 264 416
rect 258 414 259 415
rect 252 412 259 414
rect 218 410 224 411
rect 258 411 259 412
rect 263 411 264 415
rect 258 410 264 411
rect 110 403 116 404
rect 110 399 111 403
rect 115 399 116 403
rect 110 398 116 399
rect 112 391 114 398
rect 182 396 188 397
rect 182 392 183 396
rect 187 392 188 396
rect 182 391 188 392
rect 222 396 228 397
rect 222 392 223 396
rect 227 392 228 396
rect 222 391 228 392
rect 262 396 268 397
rect 262 392 263 396
rect 267 392 268 396
rect 262 391 268 392
rect 111 390 115 391
rect 111 385 115 386
rect 135 390 139 391
rect 135 385 139 386
rect 175 390 179 391
rect 175 385 179 386
rect 183 390 187 391
rect 183 385 187 386
rect 223 390 227 391
rect 223 385 227 386
rect 231 390 235 391
rect 231 385 235 386
rect 263 390 267 391
rect 263 385 267 386
rect 287 390 291 391
rect 287 385 291 386
rect 112 378 114 385
rect 134 384 140 385
rect 134 380 135 384
rect 139 380 140 384
rect 134 379 140 380
rect 174 384 180 385
rect 174 380 175 384
rect 179 380 180 384
rect 174 379 180 380
rect 230 384 236 385
rect 230 380 231 384
rect 235 380 236 384
rect 230 379 236 380
rect 286 384 292 385
rect 286 380 287 384
rect 291 380 292 384
rect 286 379 292 380
rect 110 377 116 378
rect 110 373 111 377
rect 115 373 116 377
rect 110 372 116 373
rect 300 364 302 446
rect 312 444 314 453
rect 344 452 346 494
rect 414 473 420 474
rect 414 469 415 473
rect 419 469 420 473
rect 414 468 420 469
rect 494 473 500 474
rect 494 469 495 473
rect 499 469 500 473
rect 494 468 500 469
rect 564 468 566 554
rect 622 540 628 541
rect 622 536 623 540
rect 627 536 628 540
rect 622 535 628 536
rect 702 540 708 541
rect 702 536 703 540
rect 707 536 708 540
rect 702 535 708 536
rect 782 540 788 541
rect 782 536 783 540
rect 787 536 788 540
rect 782 535 788 536
rect 624 527 626 535
rect 704 527 706 535
rect 784 527 786 535
rect 575 526 579 527
rect 575 521 579 522
rect 623 526 627 527
rect 623 521 627 522
rect 647 526 651 527
rect 647 521 651 522
rect 703 526 707 527
rect 703 521 707 522
rect 719 526 723 527
rect 719 521 723 522
rect 783 526 787 527
rect 783 521 787 522
rect 574 520 580 521
rect 574 516 575 520
rect 579 516 580 520
rect 574 515 580 516
rect 646 520 652 521
rect 646 516 647 520
rect 651 516 652 520
rect 646 515 652 516
rect 718 520 724 521
rect 718 516 719 520
rect 723 516 724 520
rect 718 515 724 516
rect 782 520 788 521
rect 782 516 783 520
rect 787 516 788 520
rect 782 515 788 516
rect 804 508 806 590
rect 812 560 814 590
rect 856 588 858 597
rect 882 595 888 596
rect 882 591 883 595
rect 887 591 888 595
rect 882 590 888 591
rect 854 587 860 588
rect 854 583 855 587
rect 859 583 860 587
rect 854 582 860 583
rect 884 560 886 590
rect 904 565 906 610
rect 920 603 922 620
rect 976 616 978 646
rect 982 625 988 626
rect 982 621 983 625
rect 987 621 988 625
rect 982 620 988 621
rect 974 615 980 616
rect 974 611 975 615
rect 979 611 980 615
rect 974 610 980 611
rect 984 603 986 620
rect 1024 616 1026 646
rect 1038 625 1044 626
rect 1038 621 1039 625
rect 1043 621 1044 625
rect 1038 620 1044 621
rect 1022 615 1028 616
rect 1022 611 1023 615
rect 1027 611 1028 615
rect 1022 610 1028 611
rect 1040 603 1042 620
rect 1088 616 1090 646
rect 1094 625 1100 626
rect 1094 621 1095 625
rect 1099 621 1100 625
rect 1094 620 1100 621
rect 1086 615 1092 616
rect 1086 611 1087 615
rect 1091 611 1092 615
rect 1086 610 1092 611
rect 1096 603 1098 620
rect 1144 616 1146 646
rect 1150 625 1156 626
rect 1150 621 1151 625
rect 1155 621 1156 625
rect 1150 620 1156 621
rect 1142 615 1148 616
rect 1142 611 1143 615
rect 1147 611 1148 615
rect 1142 610 1148 611
rect 1152 603 1154 620
rect 1180 616 1182 646
rect 1190 625 1196 626
rect 1190 621 1191 625
rect 1195 621 1196 625
rect 1190 620 1196 621
rect 1178 615 1184 616
rect 1178 611 1179 615
rect 1183 611 1184 615
rect 1178 610 1184 611
rect 1192 603 1194 620
rect 1232 612 1234 646
rect 1238 644 1239 648
rect 1243 644 1244 648
rect 1322 647 1328 648
rect 1238 643 1244 644
rect 1278 644 1284 645
rect 1230 611 1236 612
rect 1230 607 1231 611
rect 1235 607 1236 611
rect 1230 606 1236 607
rect 1240 603 1242 643
rect 1278 640 1279 644
rect 1283 640 1284 644
rect 1322 643 1323 647
rect 1327 643 1328 647
rect 1322 642 1328 643
rect 1502 647 1508 648
rect 1502 643 1503 647
rect 1507 643 1508 647
rect 1502 642 1508 643
rect 1590 647 1596 648
rect 1590 643 1591 647
rect 1595 643 1596 647
rect 1590 642 1596 643
rect 1278 639 1284 640
rect 1406 639 1412 640
rect 1280 603 1282 639
rect 1406 635 1407 639
rect 1411 635 1412 639
rect 1406 634 1412 635
rect 1302 621 1308 622
rect 1302 617 1303 621
rect 1307 617 1308 621
rect 1302 616 1308 617
rect 1398 621 1404 622
rect 1398 617 1399 621
rect 1403 617 1404 621
rect 1398 616 1404 617
rect 1304 603 1306 616
rect 1400 603 1402 616
rect 1408 612 1410 634
rect 1504 612 1506 642
rect 1510 621 1516 622
rect 1510 617 1511 621
rect 1515 617 1516 621
rect 1510 616 1516 617
rect 1406 611 1412 612
rect 1406 607 1407 611
rect 1411 607 1412 611
rect 1406 606 1412 607
rect 1502 611 1508 612
rect 1502 607 1503 611
rect 1507 607 1508 611
rect 1502 606 1508 607
rect 1512 603 1514 616
rect 919 602 923 603
rect 919 597 923 598
rect 975 602 979 603
rect 975 597 979 598
rect 983 602 987 603
rect 983 597 987 598
rect 1023 602 1027 603
rect 1023 597 1027 598
rect 1039 602 1043 603
rect 1039 597 1043 598
rect 1079 602 1083 603
rect 1079 597 1083 598
rect 1095 602 1099 603
rect 1095 597 1099 598
rect 1135 602 1139 603
rect 1135 597 1139 598
rect 1151 602 1155 603
rect 1151 597 1155 598
rect 1191 602 1195 603
rect 1191 597 1195 598
rect 1239 602 1243 603
rect 1239 597 1243 598
rect 1279 602 1283 603
rect 1279 597 1283 598
rect 1303 602 1307 603
rect 1303 597 1307 598
rect 1399 602 1403 603
rect 1399 597 1403 598
rect 1415 602 1419 603
rect 1415 597 1419 598
rect 1455 602 1459 603
rect 1455 597 1459 598
rect 1495 602 1499 603
rect 1495 597 1499 598
rect 1511 602 1515 603
rect 1511 597 1515 598
rect 1543 602 1547 603
rect 1543 597 1547 598
rect 920 588 922 597
rect 946 595 952 596
rect 946 591 947 595
rect 951 591 952 595
rect 946 590 952 591
rect 918 587 924 588
rect 918 583 919 587
rect 923 583 924 587
rect 918 582 924 583
rect 903 564 907 565
rect 948 560 950 590
rect 976 588 978 597
rect 1002 595 1008 596
rect 1002 591 1003 595
rect 1007 591 1008 595
rect 1002 590 1008 591
rect 974 587 980 588
rect 974 583 975 587
rect 979 583 980 587
rect 974 582 980 583
rect 1004 560 1006 590
rect 1024 588 1026 597
rect 1050 595 1056 596
rect 1050 591 1051 595
rect 1055 591 1056 595
rect 1050 590 1056 591
rect 1022 587 1028 588
rect 1022 583 1023 587
rect 1027 583 1028 587
rect 1022 582 1028 583
rect 1052 560 1054 590
rect 1080 588 1082 597
rect 1106 595 1112 596
rect 1106 591 1107 595
rect 1111 591 1112 595
rect 1106 590 1112 591
rect 1078 587 1084 588
rect 1078 583 1079 587
rect 1083 583 1084 587
rect 1078 582 1084 583
rect 1108 560 1110 590
rect 1136 588 1138 597
rect 1162 595 1168 596
rect 1162 591 1163 595
rect 1167 591 1168 595
rect 1162 590 1168 591
rect 1134 587 1140 588
rect 1134 583 1135 587
rect 1139 583 1140 587
rect 1134 582 1140 583
rect 1164 560 1166 590
rect 1192 588 1194 597
rect 1190 587 1196 588
rect 1190 583 1191 587
rect 1195 583 1196 587
rect 1190 582 1196 583
rect 1240 565 1242 597
rect 1280 565 1282 597
rect 1416 588 1418 597
rect 1434 595 1440 596
rect 1434 591 1435 595
rect 1439 591 1440 595
rect 1434 590 1440 591
rect 1442 595 1448 596
rect 1442 591 1443 595
rect 1447 591 1448 595
rect 1442 590 1448 591
rect 1414 587 1420 588
rect 1414 583 1415 587
rect 1419 583 1420 587
rect 1414 582 1420 583
rect 1436 568 1438 590
rect 1434 567 1440 568
rect 1215 564 1219 565
rect 1238 564 1244 565
rect 1238 560 1239 564
rect 1243 560 1244 564
rect 810 559 816 560
rect 810 555 811 559
rect 815 555 816 559
rect 810 554 816 555
rect 882 559 888 560
rect 903 559 907 560
rect 946 559 952 560
rect 882 555 883 559
rect 887 555 888 559
rect 882 554 888 555
rect 946 555 947 559
rect 951 555 952 559
rect 946 554 952 555
rect 1002 559 1008 560
rect 1002 555 1003 559
rect 1007 555 1008 559
rect 1002 554 1008 555
rect 1050 559 1056 560
rect 1050 555 1051 559
rect 1055 555 1056 559
rect 1050 554 1056 555
rect 1106 559 1112 560
rect 1106 555 1107 559
rect 1111 555 1112 559
rect 1106 554 1112 555
rect 1162 559 1168 560
rect 1162 555 1163 559
rect 1167 555 1168 559
rect 1162 554 1168 555
rect 1214 559 1220 560
rect 1238 559 1244 560
rect 1278 564 1284 565
rect 1278 560 1279 564
rect 1283 560 1284 564
rect 1434 563 1435 567
rect 1439 563 1440 567
rect 1434 562 1440 563
rect 1444 560 1446 590
rect 1456 588 1458 597
rect 1482 595 1488 596
rect 1482 591 1483 595
rect 1487 591 1488 595
rect 1482 590 1488 591
rect 1454 587 1460 588
rect 1454 583 1455 587
rect 1459 583 1460 587
rect 1454 582 1460 583
rect 1484 560 1486 590
rect 1496 588 1498 597
rect 1544 588 1546 597
rect 1592 596 1594 642
rect 1622 621 1628 622
rect 1622 617 1623 621
rect 1627 617 1628 621
rect 1622 616 1628 617
rect 1726 621 1732 622
rect 1726 617 1727 621
rect 1731 617 1732 621
rect 1726 616 1732 617
rect 1624 603 1626 616
rect 1728 603 1730 616
rect 1736 612 1738 698
rect 1750 684 1756 685
rect 1750 680 1751 684
rect 1755 680 1756 684
rect 1750 679 1756 680
rect 1830 684 1836 685
rect 1830 680 1831 684
rect 1835 680 1836 684
rect 1830 679 1836 680
rect 1910 684 1916 685
rect 1910 680 1911 684
rect 1915 680 1916 684
rect 1910 679 1916 680
rect 1990 684 1996 685
rect 1990 680 1991 684
rect 1995 680 1996 684
rect 1990 679 1996 680
rect 2078 684 2084 685
rect 2078 680 2079 684
rect 2083 680 2084 684
rect 2078 679 2084 680
rect 2174 684 2180 685
rect 2174 680 2175 684
rect 2179 680 2180 684
rect 2174 679 2180 680
rect 1752 675 1754 679
rect 1832 675 1834 679
rect 1912 675 1914 679
rect 1992 675 1994 679
rect 2080 675 2082 679
rect 2176 675 2178 679
rect 1751 674 1755 675
rect 1751 669 1755 670
rect 1815 674 1819 675
rect 1815 669 1819 670
rect 1831 674 1835 675
rect 1831 669 1835 670
rect 1895 674 1899 675
rect 1895 669 1899 670
rect 1911 674 1915 675
rect 1911 669 1915 670
rect 1975 674 1979 675
rect 1975 669 1979 670
rect 1991 674 1995 675
rect 1991 669 1995 670
rect 2047 674 2051 675
rect 2047 669 2051 670
rect 2079 674 2083 675
rect 2079 669 2083 670
rect 2111 674 2115 675
rect 2111 669 2115 670
rect 2175 674 2179 675
rect 2175 669 2179 670
rect 2239 674 2243 675
rect 2239 669 2243 670
rect 1814 668 1820 669
rect 1814 664 1815 668
rect 1819 664 1820 668
rect 1814 663 1820 664
rect 1894 668 1900 669
rect 1894 664 1895 668
rect 1899 664 1900 668
rect 1894 663 1900 664
rect 1974 668 1980 669
rect 1974 664 1975 668
rect 1979 664 1980 668
rect 1974 663 1980 664
rect 2046 668 2052 669
rect 2046 664 2047 668
rect 2051 664 2052 668
rect 2046 663 2052 664
rect 2110 668 2116 669
rect 2110 664 2111 668
rect 2115 664 2116 668
rect 2110 663 2116 664
rect 2174 668 2180 669
rect 2174 664 2175 668
rect 2179 664 2180 668
rect 2174 663 2180 664
rect 2238 668 2244 669
rect 2238 664 2239 668
rect 2243 664 2244 668
rect 2238 663 2244 664
rect 1886 647 1892 648
rect 1886 643 1887 647
rect 1891 643 1892 647
rect 1886 642 1892 643
rect 1966 647 1972 648
rect 1966 643 1967 647
rect 1971 643 1972 647
rect 1966 642 1972 643
rect 2022 647 2028 648
rect 2022 643 2023 647
rect 2027 643 2028 647
rect 2022 642 2028 643
rect 1822 639 1828 640
rect 1822 635 1823 639
rect 1827 635 1828 639
rect 1822 634 1828 635
rect 1814 621 1820 622
rect 1814 617 1815 621
rect 1819 617 1820 621
rect 1814 616 1820 617
rect 1734 611 1740 612
rect 1734 607 1735 611
rect 1739 607 1740 611
rect 1734 606 1740 607
rect 1816 603 1818 616
rect 1824 612 1826 634
rect 1888 612 1890 642
rect 1894 621 1900 622
rect 1894 617 1895 621
rect 1899 617 1900 621
rect 1894 616 1900 617
rect 1822 611 1828 612
rect 1822 607 1823 611
rect 1827 607 1828 611
rect 1822 606 1828 607
rect 1886 611 1892 612
rect 1886 607 1887 611
rect 1891 607 1892 611
rect 1886 606 1892 607
rect 1896 603 1898 616
rect 1968 612 1970 642
rect 1974 621 1980 622
rect 1974 617 1975 621
rect 1979 617 1980 621
rect 1974 616 1980 617
rect 1966 611 1972 612
rect 1966 607 1967 611
rect 1971 607 1972 611
rect 1966 606 1972 607
rect 1976 603 1978 616
rect 1599 602 1603 603
rect 1599 597 1603 598
rect 1623 602 1627 603
rect 1623 597 1627 598
rect 1663 602 1667 603
rect 1663 597 1667 598
rect 1727 602 1731 603
rect 1727 597 1731 598
rect 1791 602 1795 603
rect 1791 597 1795 598
rect 1815 602 1819 603
rect 1815 597 1819 598
rect 1847 602 1851 603
rect 1847 597 1851 598
rect 1895 602 1899 603
rect 1895 597 1899 598
rect 1911 602 1915 603
rect 1911 597 1915 598
rect 1975 602 1979 603
rect 1975 597 1979 598
rect 1582 595 1588 596
rect 1582 591 1583 595
rect 1587 591 1588 595
rect 1582 590 1588 591
rect 1590 595 1596 596
rect 1590 591 1591 595
rect 1595 591 1596 595
rect 1590 590 1596 591
rect 1494 587 1500 588
rect 1494 583 1495 587
rect 1499 583 1500 587
rect 1494 582 1500 583
rect 1542 587 1548 588
rect 1542 583 1543 587
rect 1547 583 1548 587
rect 1542 582 1548 583
rect 1584 572 1586 590
rect 1600 588 1602 597
rect 1634 595 1640 596
rect 1634 591 1635 595
rect 1639 591 1640 595
rect 1634 590 1640 591
rect 1598 587 1604 588
rect 1598 583 1599 587
rect 1603 583 1604 587
rect 1598 582 1604 583
rect 1582 571 1588 572
rect 1582 567 1583 571
rect 1587 567 1588 571
rect 1582 566 1588 567
rect 1636 564 1638 590
rect 1664 588 1666 597
rect 1690 595 1696 596
rect 1690 591 1691 595
rect 1695 591 1696 595
rect 1690 590 1696 591
rect 1662 587 1668 588
rect 1662 583 1663 587
rect 1667 583 1668 587
rect 1662 582 1668 583
rect 1634 563 1640 564
rect 1278 559 1284 560
rect 1442 559 1448 560
rect 1214 555 1215 559
rect 1219 555 1220 559
rect 1214 554 1220 555
rect 1442 555 1443 559
rect 1447 555 1448 559
rect 1442 554 1448 555
rect 1482 559 1488 560
rect 1482 555 1483 559
rect 1487 555 1488 559
rect 1482 554 1488 555
rect 1558 559 1564 560
rect 1558 555 1559 559
rect 1563 555 1564 559
rect 1634 559 1635 563
rect 1639 559 1640 563
rect 1692 560 1694 590
rect 1728 588 1730 597
rect 1792 588 1794 597
rect 1848 588 1850 597
rect 1912 588 1914 597
rect 1976 588 1978 597
rect 2024 596 2026 642
rect 2046 621 2052 622
rect 2046 617 2047 621
rect 2051 617 2052 621
rect 2046 616 2052 617
rect 2110 621 2116 622
rect 2110 617 2111 621
rect 2115 617 2116 621
rect 2110 616 2116 617
rect 2174 621 2180 622
rect 2174 617 2175 621
rect 2179 617 2180 621
rect 2174 616 2180 617
rect 2238 621 2244 622
rect 2238 617 2239 621
rect 2243 617 2244 621
rect 2238 616 2244 617
rect 2048 603 2050 616
rect 2112 603 2114 616
rect 2176 603 2178 616
rect 2240 603 2242 616
rect 2248 612 2250 698
rect 2278 684 2284 685
rect 2278 680 2279 684
rect 2283 680 2284 684
rect 2278 679 2284 680
rect 2280 675 2282 679
rect 2279 674 2283 675
rect 2279 669 2283 670
rect 2288 648 2290 746
rect 2303 741 2307 742
rect 2359 741 2363 742
rect 2360 732 2362 741
rect 2372 740 2374 782
rect 2406 780 2407 784
rect 2411 780 2412 784
rect 2406 779 2412 780
rect 2408 747 2410 779
rect 2407 746 2411 747
rect 2407 741 2411 742
rect 2370 739 2376 740
rect 2370 735 2371 739
rect 2375 735 2376 739
rect 2370 734 2376 735
rect 2358 731 2364 732
rect 2358 727 2359 731
rect 2363 727 2364 731
rect 2358 726 2364 727
rect 2408 709 2410 741
rect 2406 708 2412 709
rect 2406 704 2407 708
rect 2411 704 2412 708
rect 2378 703 2384 704
rect 2406 703 2412 704
rect 2378 699 2379 703
rect 2383 699 2384 703
rect 2378 698 2384 699
rect 2358 684 2364 685
rect 2358 680 2359 684
rect 2363 680 2364 684
rect 2358 679 2364 680
rect 2360 675 2362 679
rect 2311 674 2315 675
rect 2311 669 2315 670
rect 2359 674 2363 675
rect 2359 669 2363 670
rect 2310 668 2316 669
rect 2310 664 2311 668
rect 2315 664 2316 668
rect 2310 663 2316 664
rect 2358 668 2364 669
rect 2358 664 2359 668
rect 2363 664 2364 668
rect 2358 663 2364 664
rect 2286 647 2292 648
rect 2286 643 2287 647
rect 2291 643 2292 647
rect 2286 642 2292 643
rect 2370 647 2376 648
rect 2370 643 2371 647
rect 2375 643 2376 647
rect 2370 642 2376 643
rect 2310 621 2316 622
rect 2310 617 2311 621
rect 2315 617 2316 621
rect 2310 616 2316 617
rect 2358 621 2364 622
rect 2358 617 2359 621
rect 2363 617 2364 621
rect 2358 616 2364 617
rect 2246 611 2252 612
rect 2246 607 2247 611
rect 2251 607 2252 611
rect 2246 606 2252 607
rect 2302 611 2308 612
rect 2302 607 2303 611
rect 2307 607 2308 611
rect 2302 606 2308 607
rect 2047 602 2051 603
rect 2047 597 2051 598
rect 2111 602 2115 603
rect 2111 597 2115 598
rect 2119 602 2123 603
rect 2119 597 2123 598
rect 2175 602 2179 603
rect 2175 597 2179 598
rect 2199 602 2203 603
rect 2199 597 2203 598
rect 2239 602 2243 603
rect 2239 597 2243 598
rect 2287 602 2291 603
rect 2287 597 2291 598
rect 2014 595 2020 596
rect 2014 591 2015 595
rect 2019 591 2020 595
rect 2014 590 2020 591
rect 2022 595 2028 596
rect 2022 591 2023 595
rect 2027 591 2028 595
rect 2022 590 2028 591
rect 1726 587 1732 588
rect 1726 583 1727 587
rect 1731 583 1732 587
rect 1726 582 1732 583
rect 1790 587 1796 588
rect 1790 583 1791 587
rect 1795 583 1796 587
rect 1790 582 1796 583
rect 1846 587 1852 588
rect 1846 583 1847 587
rect 1851 583 1852 587
rect 1846 582 1852 583
rect 1910 587 1916 588
rect 1910 583 1911 587
rect 1915 583 1916 587
rect 1910 582 1916 583
rect 1974 587 1980 588
rect 1974 583 1975 587
rect 1979 583 1980 587
rect 1974 582 1980 583
rect 2016 568 2018 590
rect 2048 588 2050 597
rect 2074 595 2080 596
rect 2074 591 2075 595
rect 2079 591 2080 595
rect 2074 590 2080 591
rect 2046 587 2052 588
rect 2046 583 2047 587
rect 2051 583 2052 587
rect 2046 582 2052 583
rect 2014 567 2020 568
rect 2014 563 2015 567
rect 2019 563 2020 567
rect 2014 562 2020 563
rect 2076 560 2078 590
rect 2120 588 2122 597
rect 2146 595 2152 596
rect 2146 591 2147 595
rect 2151 591 2152 595
rect 2146 590 2152 591
rect 2118 587 2124 588
rect 2118 583 2119 587
rect 2123 583 2124 587
rect 2118 582 2124 583
rect 2148 560 2150 590
rect 2200 588 2202 597
rect 2288 588 2290 597
rect 2294 595 2300 596
rect 2294 591 2295 595
rect 2299 591 2300 595
rect 2294 590 2300 591
rect 2198 587 2204 588
rect 2198 583 2199 587
rect 2203 583 2204 587
rect 2198 582 2204 583
rect 2286 587 2292 588
rect 2286 583 2287 587
rect 2291 583 2292 587
rect 2286 582 2292 583
rect 1634 558 1640 559
rect 1690 559 1696 560
rect 1558 554 1564 555
rect 1690 555 1691 559
rect 1695 555 1696 559
rect 1690 554 1696 555
rect 1894 559 1900 560
rect 1894 555 1895 559
rect 1899 555 1900 559
rect 1894 554 1900 555
rect 2074 559 2080 560
rect 2074 555 2075 559
rect 2079 555 2080 559
rect 2074 554 2080 555
rect 2146 559 2152 560
rect 2146 555 2147 559
rect 2151 555 2152 559
rect 2146 554 2152 555
rect 1238 547 1244 548
rect 1238 543 1239 547
rect 1243 543 1244 547
rect 1238 542 1244 543
rect 1278 547 1284 548
rect 1278 543 1279 547
rect 1283 543 1284 547
rect 1278 542 1284 543
rect 854 540 860 541
rect 854 536 855 540
rect 859 536 860 540
rect 854 535 860 536
rect 918 540 924 541
rect 918 536 919 540
rect 923 536 924 540
rect 918 535 924 536
rect 974 540 980 541
rect 974 536 975 540
rect 979 536 980 540
rect 974 535 980 536
rect 1022 540 1028 541
rect 1022 536 1023 540
rect 1027 536 1028 540
rect 1022 535 1028 536
rect 1078 540 1084 541
rect 1078 536 1079 540
rect 1083 536 1084 540
rect 1078 535 1084 536
rect 1134 540 1140 541
rect 1134 536 1135 540
rect 1139 536 1140 540
rect 1134 535 1140 536
rect 1190 540 1196 541
rect 1190 536 1191 540
rect 1195 536 1196 540
rect 1190 535 1196 536
rect 856 527 858 535
rect 920 527 922 535
rect 976 527 978 535
rect 1024 527 1026 535
rect 1080 527 1082 535
rect 1136 527 1138 535
rect 1192 527 1194 535
rect 1240 527 1242 542
rect 1280 535 1282 542
rect 1414 540 1420 541
rect 1414 536 1415 540
rect 1419 536 1420 540
rect 1414 535 1420 536
rect 1454 540 1460 541
rect 1454 536 1455 540
rect 1459 536 1460 540
rect 1454 535 1460 536
rect 1494 540 1500 541
rect 1494 536 1495 540
rect 1499 536 1500 540
rect 1494 535 1500 536
rect 1542 540 1548 541
rect 1542 536 1543 540
rect 1547 536 1548 540
rect 1542 535 1548 536
rect 1279 534 1283 535
rect 1279 529 1283 530
rect 1303 534 1307 535
rect 1303 529 1307 530
rect 1375 534 1379 535
rect 1375 529 1379 530
rect 1415 534 1419 535
rect 1415 529 1419 530
rect 1455 534 1459 535
rect 1455 529 1459 530
rect 1479 534 1483 535
rect 1479 529 1483 530
rect 1495 534 1499 535
rect 1495 529 1499 530
rect 1543 534 1547 535
rect 1543 529 1547 530
rect 847 526 851 527
rect 847 521 851 522
rect 855 526 859 527
rect 855 521 859 522
rect 903 526 907 527
rect 903 521 907 522
rect 919 526 923 527
rect 919 521 923 522
rect 959 526 963 527
rect 959 521 963 522
rect 975 526 979 527
rect 975 521 979 522
rect 1023 526 1027 527
rect 1023 521 1027 522
rect 1079 526 1083 527
rect 1079 521 1083 522
rect 1087 526 1091 527
rect 1087 521 1091 522
rect 1135 526 1139 527
rect 1135 521 1139 522
rect 1151 526 1155 527
rect 1151 521 1155 522
rect 1191 526 1195 527
rect 1191 521 1195 522
rect 1239 526 1243 527
rect 1280 522 1282 529
rect 1302 528 1308 529
rect 1302 524 1303 528
rect 1307 524 1308 528
rect 1302 523 1308 524
rect 1374 528 1380 529
rect 1374 524 1375 528
rect 1379 524 1380 528
rect 1374 523 1380 524
rect 1478 528 1484 529
rect 1478 524 1479 528
rect 1483 524 1484 528
rect 1478 523 1484 524
rect 1239 521 1243 522
rect 1278 521 1284 522
rect 846 520 852 521
rect 846 516 847 520
rect 851 516 852 520
rect 846 515 852 516
rect 902 520 908 521
rect 902 516 903 520
rect 907 516 908 520
rect 902 515 908 516
rect 958 520 964 521
rect 958 516 959 520
rect 963 516 964 520
rect 958 515 964 516
rect 1022 520 1028 521
rect 1022 516 1023 520
rect 1027 516 1028 520
rect 1022 515 1028 516
rect 1086 520 1092 521
rect 1086 516 1087 520
rect 1091 516 1092 520
rect 1086 515 1092 516
rect 1150 520 1156 521
rect 1150 516 1151 520
rect 1155 516 1156 520
rect 1150 515 1156 516
rect 1190 520 1196 521
rect 1190 516 1191 520
rect 1195 516 1196 520
rect 1190 515 1196 516
rect 1240 514 1242 521
rect 1278 517 1279 521
rect 1283 517 1284 521
rect 1278 516 1284 517
rect 1238 513 1244 514
rect 1238 509 1239 513
rect 1243 509 1244 513
rect 1238 508 1244 509
rect 802 507 808 508
rect 802 503 803 507
rect 807 503 808 507
rect 1310 507 1316 508
rect 802 502 808 503
rect 1278 504 1284 505
rect 1278 500 1279 504
rect 1283 500 1284 504
rect 1310 503 1311 507
rect 1315 503 1316 507
rect 1310 502 1316 503
rect 710 499 716 500
rect 710 495 711 499
rect 715 495 716 499
rect 710 494 716 495
rect 838 499 844 500
rect 838 495 839 499
rect 843 495 844 499
rect 838 494 844 495
rect 894 499 900 500
rect 894 495 895 499
rect 899 495 900 499
rect 894 494 900 495
rect 950 499 956 500
rect 950 495 951 499
rect 955 495 956 499
rect 950 494 956 495
rect 1014 499 1020 500
rect 1014 495 1015 499
rect 1019 495 1020 499
rect 1014 494 1020 495
rect 1142 499 1148 500
rect 1142 495 1143 499
rect 1147 495 1148 499
rect 1142 494 1148 495
rect 1178 499 1184 500
rect 1178 495 1179 499
rect 1183 495 1184 499
rect 1178 494 1184 495
rect 1230 499 1236 500
rect 1278 499 1284 500
rect 1230 495 1231 499
rect 1235 495 1236 499
rect 1230 494 1236 495
rect 1238 496 1244 497
rect 574 473 580 474
rect 574 469 575 473
rect 579 469 580 473
rect 574 468 580 469
rect 646 473 652 474
rect 646 469 647 473
rect 651 469 652 473
rect 646 468 652 469
rect 416 459 418 468
rect 496 459 498 468
rect 562 467 568 468
rect 562 463 563 467
rect 567 463 568 467
rect 562 462 568 463
rect 576 459 578 468
rect 648 459 650 468
rect 712 464 714 494
rect 718 473 724 474
rect 718 469 719 473
rect 723 469 724 473
rect 718 468 724 469
rect 782 473 788 474
rect 782 469 783 473
rect 787 469 788 473
rect 782 468 788 469
rect 690 463 696 464
rect 690 459 691 463
rect 695 459 696 463
rect 367 458 371 459
rect 367 453 371 454
rect 415 458 419 459
rect 415 453 419 454
rect 431 458 435 459
rect 431 453 435 454
rect 495 458 499 459
rect 495 453 499 454
rect 559 458 563 459
rect 559 453 563 454
rect 575 458 579 459
rect 575 453 579 454
rect 615 458 619 459
rect 615 453 619 454
rect 647 458 651 459
rect 647 453 651 454
rect 671 458 675 459
rect 690 458 696 459
rect 710 463 716 464
rect 710 459 711 463
rect 715 459 716 463
rect 720 459 722 468
rect 784 459 786 468
rect 840 464 842 494
rect 846 473 852 474
rect 846 469 847 473
rect 851 469 852 473
rect 846 468 852 469
rect 838 463 844 464
rect 838 459 839 463
rect 843 459 844 463
rect 848 459 850 468
rect 896 464 898 494
rect 902 473 908 474
rect 902 469 903 473
rect 907 469 908 473
rect 902 468 908 469
rect 894 463 900 464
rect 894 459 895 463
rect 899 459 900 463
rect 904 459 906 468
rect 952 464 954 494
rect 958 473 964 474
rect 958 469 959 473
rect 963 469 964 473
rect 958 468 964 469
rect 950 463 956 464
rect 950 459 951 463
rect 955 459 956 463
rect 960 459 962 468
rect 1016 464 1018 494
rect 1094 487 1100 488
rect 1094 483 1095 487
rect 1099 483 1100 487
rect 1094 482 1100 483
rect 1022 473 1028 474
rect 1022 469 1023 473
rect 1027 469 1028 473
rect 1022 468 1028 469
rect 1086 473 1092 474
rect 1086 469 1087 473
rect 1091 469 1092 473
rect 1086 468 1092 469
rect 1014 463 1020 464
rect 1014 459 1015 463
rect 1019 459 1020 463
rect 1024 459 1026 468
rect 1088 459 1090 468
rect 1096 464 1098 482
rect 1144 464 1146 494
rect 1150 473 1156 474
rect 1150 469 1151 473
rect 1155 469 1156 473
rect 1150 468 1156 469
rect 1094 463 1100 464
rect 1094 459 1095 463
rect 1099 459 1100 463
rect 710 458 716 459
rect 719 458 723 459
rect 671 453 675 454
rect 342 451 348 452
rect 342 447 343 451
rect 347 447 348 451
rect 342 446 348 447
rect 350 451 356 452
rect 350 447 351 451
rect 355 447 356 451
rect 350 446 356 447
rect 310 443 316 444
rect 310 439 311 443
rect 315 439 316 443
rect 310 438 316 439
rect 352 416 354 446
rect 368 444 370 453
rect 394 451 400 452
rect 394 447 395 451
rect 399 447 400 451
rect 394 446 400 447
rect 366 443 372 444
rect 366 439 367 443
rect 371 439 372 443
rect 366 438 372 439
rect 396 416 398 446
rect 432 444 434 453
rect 458 451 464 452
rect 458 447 459 451
rect 463 447 464 451
rect 458 446 464 447
rect 430 443 436 444
rect 430 439 431 443
rect 435 439 436 443
rect 430 438 436 439
rect 460 416 462 446
rect 496 444 498 453
rect 560 444 562 453
rect 566 451 572 452
rect 566 447 567 451
rect 571 447 572 451
rect 566 446 572 447
rect 586 451 592 452
rect 586 447 587 451
rect 591 447 592 451
rect 586 446 592 447
rect 494 443 500 444
rect 494 439 495 443
rect 499 439 500 443
rect 494 438 500 439
rect 558 443 564 444
rect 558 439 559 443
rect 563 439 564 443
rect 558 438 564 439
rect 350 415 356 416
rect 350 411 351 415
rect 355 411 356 415
rect 350 410 356 411
rect 394 415 400 416
rect 394 411 395 415
rect 399 411 400 415
rect 394 410 400 411
rect 458 415 464 416
rect 458 411 459 415
rect 463 411 464 415
rect 458 410 464 411
rect 466 415 472 416
rect 466 411 467 415
rect 471 411 472 415
rect 466 410 472 411
rect 310 396 316 397
rect 310 392 311 396
rect 315 392 316 396
rect 310 391 316 392
rect 366 396 372 397
rect 366 392 367 396
rect 371 392 372 396
rect 366 391 372 392
rect 430 396 436 397
rect 430 392 431 396
rect 435 392 436 396
rect 430 391 436 392
rect 311 390 315 391
rect 311 385 315 386
rect 343 390 347 391
rect 343 385 347 386
rect 367 390 371 391
rect 367 385 371 386
rect 391 390 395 391
rect 391 385 395 386
rect 431 390 435 391
rect 431 385 435 386
rect 439 390 443 391
rect 439 385 443 386
rect 342 384 348 385
rect 342 380 343 384
rect 347 380 348 384
rect 342 379 348 380
rect 390 384 396 385
rect 390 380 391 384
rect 395 380 396 384
rect 390 379 396 380
rect 438 384 444 385
rect 438 380 439 384
rect 443 380 444 384
rect 438 379 444 380
rect 162 363 168 364
rect 110 360 116 361
rect 110 356 111 360
rect 115 356 116 360
rect 162 359 163 363
rect 167 359 168 363
rect 162 358 168 359
rect 222 363 228 364
rect 222 359 223 363
rect 227 359 228 363
rect 222 358 228 359
rect 278 363 284 364
rect 278 359 279 363
rect 283 359 284 363
rect 278 358 284 359
rect 298 363 304 364
rect 298 359 299 363
rect 303 359 304 363
rect 298 358 304 359
rect 334 363 340 364
rect 334 359 335 363
rect 339 359 340 363
rect 334 358 340 359
rect 110 355 116 356
rect 112 319 114 355
rect 134 337 140 338
rect 134 333 135 337
rect 139 333 140 337
rect 134 332 140 333
rect 136 319 138 332
rect 164 328 166 358
rect 174 337 180 338
rect 174 333 175 337
rect 179 333 180 337
rect 174 332 180 333
rect 162 327 168 328
rect 162 323 163 327
rect 167 323 168 327
rect 162 322 168 323
rect 176 319 178 332
rect 224 328 226 358
rect 230 337 236 338
rect 230 333 231 337
rect 235 333 236 337
rect 230 332 236 333
rect 222 327 228 328
rect 222 323 223 327
rect 227 323 228 327
rect 222 322 228 323
rect 232 319 234 332
rect 280 328 282 358
rect 286 337 292 338
rect 286 333 287 337
rect 291 333 292 337
rect 286 332 292 333
rect 278 327 284 328
rect 278 323 279 327
rect 283 323 284 327
rect 278 322 284 323
rect 278 319 284 320
rect 288 319 290 332
rect 111 318 115 319
rect 111 313 115 314
rect 135 318 139 319
rect 135 313 139 314
rect 175 318 179 319
rect 175 313 179 314
rect 183 318 187 319
rect 183 313 187 314
rect 231 318 235 319
rect 231 313 235 314
rect 255 318 259 319
rect 278 315 279 319
rect 283 315 284 319
rect 278 314 284 315
rect 287 318 291 319
rect 255 313 259 314
rect 112 281 114 313
rect 136 304 138 313
rect 154 311 160 312
rect 154 307 155 311
rect 159 307 160 311
rect 154 306 160 307
rect 162 311 168 312
rect 162 307 163 311
rect 167 307 168 311
rect 162 306 168 307
rect 134 303 140 304
rect 134 299 135 303
rect 139 299 140 303
rect 134 298 140 299
rect 110 280 116 281
rect 110 276 111 280
rect 115 276 116 280
rect 110 275 116 276
rect 110 263 116 264
rect 110 259 111 263
rect 115 259 116 263
rect 110 258 116 259
rect 112 243 114 258
rect 134 256 140 257
rect 134 252 135 256
rect 139 252 140 256
rect 134 251 140 252
rect 136 243 138 251
rect 111 242 115 243
rect 111 237 115 238
rect 135 242 139 243
rect 135 237 139 238
rect 112 230 114 237
rect 134 236 140 237
rect 134 232 135 236
rect 139 232 140 236
rect 134 231 140 232
rect 110 229 116 230
rect 110 225 111 229
rect 115 225 116 229
rect 110 224 116 225
rect 156 216 158 306
rect 164 276 166 306
rect 184 304 186 313
rect 210 311 216 312
rect 210 307 211 311
rect 215 307 216 311
rect 210 306 216 307
rect 182 303 188 304
rect 182 299 183 303
rect 187 299 188 303
rect 182 298 188 299
rect 212 276 214 306
rect 256 304 258 313
rect 254 303 260 304
rect 254 299 255 303
rect 259 299 260 303
rect 254 298 260 299
rect 280 276 282 314
rect 287 313 291 314
rect 327 318 331 319
rect 327 313 331 314
rect 328 304 330 313
rect 336 312 338 358
rect 342 337 348 338
rect 342 333 343 337
rect 347 333 348 337
rect 342 332 348 333
rect 390 337 396 338
rect 390 333 391 337
rect 395 333 396 337
rect 390 332 396 333
rect 438 337 444 338
rect 438 333 439 337
rect 443 333 444 337
rect 438 332 444 333
rect 344 319 346 332
rect 392 319 394 332
rect 440 319 442 332
rect 468 328 470 410
rect 494 396 500 397
rect 494 392 495 396
rect 499 392 500 396
rect 494 391 500 392
rect 558 396 564 397
rect 558 392 559 396
rect 563 392 564 396
rect 558 391 564 392
rect 487 390 491 391
rect 487 385 491 386
rect 495 390 499 391
rect 495 385 499 386
rect 535 390 539 391
rect 535 385 539 386
rect 559 390 563 391
rect 559 385 563 386
rect 486 384 492 385
rect 486 380 487 384
rect 491 380 492 384
rect 486 379 492 380
rect 534 384 540 385
rect 534 380 535 384
rect 539 380 540 384
rect 534 379 540 380
rect 568 376 570 446
rect 588 416 590 446
rect 616 444 618 453
rect 672 444 674 453
rect 614 443 620 444
rect 614 439 615 443
rect 619 439 620 443
rect 614 438 620 439
rect 670 443 676 444
rect 670 439 671 443
rect 675 439 676 443
rect 670 438 676 439
rect 692 424 694 458
rect 719 453 723 454
rect 775 458 779 459
rect 775 453 779 454
rect 783 458 787 459
rect 783 453 787 454
rect 831 458 835 459
rect 838 458 844 459
rect 847 458 851 459
rect 831 453 835 454
rect 847 453 851 454
rect 887 458 891 459
rect 894 458 900 459
rect 903 458 907 459
rect 950 458 956 459
rect 959 458 963 459
rect 1014 458 1020 459
rect 1023 458 1027 459
rect 887 453 891 454
rect 903 453 907 454
rect 959 453 963 454
rect 1023 453 1027 454
rect 1087 458 1091 459
rect 1094 458 1100 459
rect 1142 463 1148 464
rect 1142 459 1143 463
rect 1147 459 1148 463
rect 1152 459 1154 468
rect 1180 464 1182 494
rect 1190 473 1196 474
rect 1190 469 1191 473
rect 1195 469 1196 473
rect 1232 472 1234 494
rect 1238 492 1239 496
rect 1243 492 1244 496
rect 1238 491 1244 492
rect 1190 468 1196 469
rect 1230 471 1236 472
rect 1178 463 1184 464
rect 1178 459 1179 463
rect 1183 459 1184 463
rect 1192 459 1194 468
rect 1230 467 1231 471
rect 1235 467 1236 471
rect 1230 466 1236 467
rect 1240 459 1242 491
rect 1280 463 1282 499
rect 1302 481 1308 482
rect 1302 477 1303 481
rect 1307 477 1308 481
rect 1302 476 1308 477
rect 1304 463 1306 476
rect 1279 462 1283 463
rect 1142 458 1148 459
rect 1151 458 1155 459
rect 1178 458 1184 459
rect 1191 458 1195 459
rect 1087 453 1091 454
rect 1151 453 1155 454
rect 1191 453 1195 454
rect 1239 458 1243 459
rect 1279 457 1283 458
rect 1303 462 1307 463
rect 1303 457 1307 458
rect 1239 453 1243 454
rect 698 451 704 452
rect 698 447 699 451
rect 703 447 704 451
rect 698 446 704 447
rect 690 423 696 424
rect 690 419 691 423
rect 695 419 696 423
rect 690 418 696 419
rect 700 416 702 446
rect 720 444 722 453
rect 776 444 778 453
rect 802 451 808 452
rect 802 447 803 451
rect 807 447 808 451
rect 802 446 808 447
rect 718 443 724 444
rect 718 439 719 443
rect 723 439 724 443
rect 718 438 724 439
rect 774 443 780 444
rect 774 439 775 443
rect 779 439 780 443
rect 774 438 780 439
rect 804 416 806 446
rect 832 444 834 453
rect 858 451 864 452
rect 858 447 859 451
rect 863 447 864 451
rect 858 446 864 447
rect 830 443 836 444
rect 830 439 831 443
rect 835 439 836 443
rect 830 438 836 439
rect 860 416 862 446
rect 888 444 890 453
rect 886 443 892 444
rect 886 439 887 443
rect 891 439 892 443
rect 886 438 892 439
rect 1240 421 1242 453
rect 1280 425 1282 457
rect 1304 448 1306 457
rect 1312 456 1314 502
rect 1374 481 1380 482
rect 1374 477 1375 481
rect 1379 477 1380 481
rect 1374 476 1380 477
rect 1478 481 1484 482
rect 1478 477 1479 481
rect 1483 477 1484 481
rect 1478 476 1484 477
rect 1376 463 1378 476
rect 1480 463 1482 476
rect 1560 472 1562 554
rect 1598 540 1604 541
rect 1598 536 1599 540
rect 1603 536 1604 540
rect 1598 535 1604 536
rect 1662 540 1668 541
rect 1662 536 1663 540
rect 1667 536 1668 540
rect 1662 535 1668 536
rect 1726 540 1732 541
rect 1726 536 1727 540
rect 1731 536 1732 540
rect 1726 535 1732 536
rect 1790 540 1796 541
rect 1790 536 1791 540
rect 1795 536 1796 540
rect 1790 535 1796 536
rect 1846 540 1852 541
rect 1846 536 1847 540
rect 1851 536 1852 540
rect 1846 535 1852 536
rect 1583 534 1587 535
rect 1583 529 1587 530
rect 1599 534 1603 535
rect 1599 529 1603 530
rect 1663 534 1667 535
rect 1663 529 1667 530
rect 1695 534 1699 535
rect 1695 529 1699 530
rect 1727 534 1731 535
rect 1727 529 1731 530
rect 1791 534 1795 535
rect 1791 529 1795 530
rect 1799 534 1803 535
rect 1799 529 1803 530
rect 1847 534 1851 535
rect 1847 529 1851 530
rect 1582 528 1588 529
rect 1582 524 1583 528
rect 1587 524 1588 528
rect 1582 523 1588 524
rect 1694 528 1700 529
rect 1694 524 1695 528
rect 1699 524 1700 528
rect 1694 523 1700 524
rect 1798 528 1804 529
rect 1798 524 1799 528
rect 1803 524 1804 528
rect 1798 523 1804 524
rect 1722 507 1728 508
rect 1722 503 1723 507
rect 1727 503 1728 507
rect 1722 502 1728 503
rect 1730 507 1736 508
rect 1730 503 1731 507
rect 1735 503 1736 507
rect 1730 502 1736 503
rect 1582 481 1588 482
rect 1582 477 1583 481
rect 1587 477 1588 481
rect 1582 476 1588 477
rect 1694 481 1700 482
rect 1694 477 1695 481
rect 1699 477 1700 481
rect 1694 476 1700 477
rect 1558 471 1564 472
rect 1558 467 1559 471
rect 1563 467 1564 471
rect 1558 466 1564 467
rect 1584 463 1586 476
rect 1696 463 1698 476
rect 1343 462 1347 463
rect 1343 457 1347 458
rect 1375 462 1379 463
rect 1375 457 1379 458
rect 1399 462 1403 463
rect 1399 457 1403 458
rect 1463 462 1467 463
rect 1463 457 1467 458
rect 1479 462 1483 463
rect 1479 457 1483 458
rect 1527 462 1531 463
rect 1527 457 1531 458
rect 1583 462 1587 463
rect 1583 457 1587 458
rect 1591 462 1595 463
rect 1591 457 1595 458
rect 1663 462 1667 463
rect 1663 457 1667 458
rect 1695 462 1699 463
rect 1695 457 1699 458
rect 1310 455 1316 456
rect 1310 451 1311 455
rect 1315 451 1316 455
rect 1310 450 1316 451
rect 1330 455 1336 456
rect 1330 451 1331 455
rect 1335 451 1336 455
rect 1330 450 1336 451
rect 1302 447 1308 448
rect 1302 443 1303 447
rect 1307 443 1308 447
rect 1302 442 1308 443
rect 1278 424 1284 425
rect 1238 420 1244 421
rect 1238 416 1239 420
rect 1243 416 1244 420
rect 1278 420 1279 424
rect 1283 420 1284 424
rect 1332 420 1334 450
rect 1344 448 1346 457
rect 1400 448 1402 457
rect 1426 455 1432 456
rect 1426 451 1427 455
rect 1431 451 1432 455
rect 1426 450 1432 451
rect 1342 447 1348 448
rect 1342 443 1343 447
rect 1347 443 1348 447
rect 1342 442 1348 443
rect 1398 447 1404 448
rect 1398 443 1399 447
rect 1403 443 1404 447
rect 1398 442 1404 443
rect 1428 420 1430 450
rect 1464 448 1466 457
rect 1490 455 1496 456
rect 1490 451 1491 455
rect 1495 451 1496 455
rect 1490 450 1496 451
rect 1462 447 1468 448
rect 1462 443 1463 447
rect 1467 443 1468 447
rect 1462 442 1468 443
rect 1492 420 1494 450
rect 1528 448 1530 457
rect 1592 448 1594 457
rect 1634 455 1640 456
rect 1634 451 1635 455
rect 1639 451 1640 455
rect 1634 450 1640 451
rect 1526 447 1532 448
rect 1526 443 1527 447
rect 1531 443 1532 447
rect 1526 442 1532 443
rect 1590 447 1596 448
rect 1590 443 1591 447
rect 1595 443 1596 447
rect 1590 442 1596 443
rect 1636 428 1638 450
rect 1664 448 1666 457
rect 1724 456 1726 502
rect 1732 472 1734 502
rect 1806 499 1812 500
rect 1806 495 1807 499
rect 1811 495 1812 499
rect 1806 494 1812 495
rect 1798 481 1804 482
rect 1798 477 1799 481
rect 1803 477 1804 481
rect 1798 476 1804 477
rect 1730 471 1736 472
rect 1730 467 1731 471
rect 1735 467 1736 471
rect 1730 466 1736 467
rect 1800 463 1802 476
rect 1808 472 1810 494
rect 1896 472 1898 554
rect 1910 540 1916 541
rect 1910 536 1911 540
rect 1915 536 1916 540
rect 1910 535 1916 536
rect 1974 540 1980 541
rect 1974 536 1975 540
rect 1979 536 1980 540
rect 1974 535 1980 536
rect 2046 540 2052 541
rect 2046 536 2047 540
rect 2051 536 2052 540
rect 2046 535 2052 536
rect 2118 540 2124 541
rect 2118 536 2119 540
rect 2123 536 2124 540
rect 2118 535 2124 536
rect 2198 540 2204 541
rect 2198 536 2199 540
rect 2203 536 2204 540
rect 2198 535 2204 536
rect 2286 540 2292 541
rect 2286 536 2287 540
rect 2291 536 2292 540
rect 2286 535 2292 536
rect 1903 534 1907 535
rect 1903 529 1907 530
rect 1911 534 1915 535
rect 1911 529 1915 530
rect 1975 534 1979 535
rect 1975 529 1979 530
rect 2007 534 2011 535
rect 2007 529 2011 530
rect 2047 534 2051 535
rect 2047 529 2051 530
rect 2103 534 2107 535
rect 2103 529 2107 530
rect 2119 534 2123 535
rect 2119 529 2123 530
rect 2191 534 2195 535
rect 2191 529 2195 530
rect 2199 534 2203 535
rect 2199 529 2203 530
rect 2287 534 2291 535
rect 2287 529 2291 530
rect 1902 528 1908 529
rect 1902 524 1903 528
rect 1907 524 1908 528
rect 1902 523 1908 524
rect 2006 528 2012 529
rect 2006 524 2007 528
rect 2011 524 2012 528
rect 2006 523 2012 524
rect 2102 528 2108 529
rect 2102 524 2103 528
rect 2107 524 2108 528
rect 2102 523 2108 524
rect 2190 528 2196 529
rect 2190 524 2191 528
rect 2195 524 2196 528
rect 2190 523 2196 524
rect 2286 528 2292 529
rect 2286 524 2287 528
rect 2291 524 2292 528
rect 2286 523 2292 524
rect 2296 508 2298 590
rect 2304 560 2306 606
rect 2312 603 2314 616
rect 2360 603 2362 616
rect 2311 602 2315 603
rect 2311 597 2315 598
rect 2359 602 2363 603
rect 2359 597 2363 598
rect 2360 588 2362 597
rect 2372 596 2374 642
rect 2380 612 2382 698
rect 2406 691 2412 692
rect 2406 687 2407 691
rect 2411 687 2412 691
rect 2406 686 2412 687
rect 2408 675 2410 686
rect 2407 674 2411 675
rect 2407 669 2411 670
rect 2408 662 2410 669
rect 2406 661 2412 662
rect 2406 657 2407 661
rect 2411 657 2412 661
rect 2406 656 2412 657
rect 2406 644 2412 645
rect 2406 640 2407 644
rect 2411 640 2412 644
rect 2406 639 2412 640
rect 2378 611 2384 612
rect 2378 607 2379 611
rect 2383 607 2384 611
rect 2378 606 2384 607
rect 2408 603 2410 639
rect 2407 602 2411 603
rect 2407 597 2411 598
rect 2370 595 2376 596
rect 2370 591 2371 595
rect 2375 591 2376 595
rect 2370 590 2376 591
rect 2358 587 2364 588
rect 2358 583 2359 587
rect 2363 583 2364 587
rect 2358 582 2364 583
rect 2408 565 2410 597
rect 2406 564 2412 565
rect 2406 560 2407 564
rect 2411 560 2412 564
rect 2302 559 2308 560
rect 2302 555 2303 559
rect 2307 555 2308 559
rect 2302 554 2308 555
rect 2374 559 2380 560
rect 2406 559 2412 560
rect 2374 555 2375 559
rect 2379 555 2380 559
rect 2374 554 2380 555
rect 2358 540 2364 541
rect 2358 536 2359 540
rect 2363 536 2364 540
rect 2358 535 2364 536
rect 2359 534 2363 535
rect 2359 529 2363 530
rect 2358 528 2364 529
rect 2358 524 2359 528
rect 2363 524 2364 528
rect 2358 523 2364 524
rect 1998 507 2004 508
rect 1998 503 1999 507
rect 2003 503 2004 507
rect 1998 502 2004 503
rect 2182 507 2188 508
rect 2182 503 2183 507
rect 2187 503 2188 507
rect 2182 502 2188 503
rect 2278 507 2284 508
rect 2278 503 2279 507
rect 2283 503 2284 507
rect 2278 502 2284 503
rect 2294 507 2300 508
rect 2294 503 2295 507
rect 2299 503 2300 507
rect 2294 502 2300 503
rect 2366 507 2372 508
rect 2366 503 2367 507
rect 2371 503 2372 507
rect 2366 502 2372 503
rect 1902 481 1908 482
rect 1902 477 1903 481
rect 1907 477 1908 481
rect 1902 476 1908 477
rect 1806 471 1812 472
rect 1806 467 1807 471
rect 1811 467 1812 471
rect 1806 466 1812 467
rect 1894 471 1900 472
rect 1894 467 1895 471
rect 1899 467 1900 471
rect 1894 466 1900 467
rect 1904 463 1906 476
rect 2000 472 2002 502
rect 2006 481 2012 482
rect 2006 477 2007 481
rect 2011 477 2012 481
rect 2006 476 2012 477
rect 2102 481 2108 482
rect 2102 477 2103 481
rect 2107 477 2108 481
rect 2102 476 2108 477
rect 1998 471 2004 472
rect 1998 467 1999 471
rect 2003 467 2004 471
rect 1998 466 2004 467
rect 2008 463 2010 476
rect 2104 463 2106 476
rect 2184 472 2186 502
rect 2190 481 2196 482
rect 2190 477 2191 481
rect 2195 477 2196 481
rect 2190 476 2196 477
rect 2174 471 2180 472
rect 2174 467 2175 471
rect 2179 467 2180 471
rect 2174 466 2180 467
rect 2182 471 2188 472
rect 2182 467 2183 471
rect 2187 467 2188 471
rect 2182 466 2188 467
rect 1735 462 1739 463
rect 1735 457 1739 458
rect 1799 462 1803 463
rect 1799 457 1803 458
rect 1815 462 1819 463
rect 1815 457 1819 458
rect 1895 462 1899 463
rect 1895 457 1899 458
rect 1903 462 1907 463
rect 1903 457 1907 458
rect 1975 462 1979 463
rect 1975 457 1979 458
rect 2007 462 2011 463
rect 2007 457 2011 458
rect 2055 462 2059 463
rect 2055 457 2059 458
rect 2103 462 2107 463
rect 2103 457 2107 458
rect 2135 462 2139 463
rect 2135 457 2139 458
rect 1714 455 1720 456
rect 1714 451 1715 455
rect 1719 451 1720 455
rect 1714 450 1720 451
rect 1722 455 1728 456
rect 1722 451 1723 455
rect 1727 451 1728 455
rect 1722 450 1728 451
rect 1662 447 1668 448
rect 1662 443 1663 447
rect 1667 443 1668 447
rect 1662 442 1668 443
rect 1634 427 1640 428
rect 1634 423 1635 427
rect 1639 423 1640 427
rect 1634 422 1640 423
rect 1278 419 1284 420
rect 1330 419 1336 420
rect 586 415 592 416
rect 586 411 587 415
rect 591 411 592 415
rect 586 410 592 411
rect 698 415 704 416
rect 698 411 699 415
rect 703 411 704 415
rect 698 410 704 411
rect 802 415 808 416
rect 802 411 803 415
rect 807 411 808 415
rect 802 410 808 411
rect 858 415 864 416
rect 1238 415 1244 416
rect 1330 415 1331 419
rect 1335 415 1336 419
rect 858 411 859 415
rect 863 411 864 415
rect 1330 414 1336 415
rect 1426 419 1432 420
rect 1426 415 1427 419
rect 1431 415 1432 419
rect 1426 414 1432 415
rect 1490 419 1496 420
rect 1490 415 1491 419
rect 1495 415 1496 419
rect 1490 414 1496 415
rect 1654 419 1660 420
rect 1654 415 1655 419
rect 1659 415 1660 419
rect 1654 414 1660 415
rect 858 410 864 411
rect 1454 411 1460 412
rect 1278 407 1284 408
rect 1238 403 1244 404
rect 1238 399 1239 403
rect 1243 399 1244 403
rect 1278 403 1279 407
rect 1283 403 1284 407
rect 1454 407 1455 411
rect 1459 407 1460 411
rect 1454 406 1460 407
rect 1278 402 1284 403
rect 1238 398 1244 399
rect 614 396 620 397
rect 614 392 615 396
rect 619 392 620 396
rect 614 391 620 392
rect 670 396 676 397
rect 670 392 671 396
rect 675 392 676 396
rect 670 391 676 392
rect 718 396 724 397
rect 718 392 719 396
rect 723 392 724 396
rect 718 391 724 392
rect 774 396 780 397
rect 774 392 775 396
rect 779 392 780 396
rect 774 391 780 392
rect 830 396 836 397
rect 830 392 831 396
rect 835 392 836 396
rect 830 391 836 392
rect 886 396 892 397
rect 886 392 887 396
rect 891 392 892 396
rect 886 391 892 392
rect 1240 391 1242 398
rect 1280 391 1282 402
rect 1302 400 1308 401
rect 1302 396 1303 400
rect 1307 396 1308 400
rect 1302 395 1308 396
rect 1342 400 1348 401
rect 1342 396 1343 400
rect 1347 396 1348 400
rect 1342 395 1348 396
rect 1398 400 1404 401
rect 1398 396 1399 400
rect 1403 396 1404 400
rect 1398 395 1404 396
rect 1304 391 1306 395
rect 1344 391 1346 395
rect 1400 391 1402 395
rect 583 390 587 391
rect 583 385 587 386
rect 615 390 619 391
rect 615 385 619 386
rect 631 390 635 391
rect 631 385 635 386
rect 671 390 675 391
rect 671 385 675 386
rect 679 390 683 391
rect 679 385 683 386
rect 719 390 723 391
rect 719 385 723 386
rect 727 390 731 391
rect 727 385 731 386
rect 775 390 779 391
rect 775 385 779 386
rect 831 390 835 391
rect 831 385 835 386
rect 887 390 891 391
rect 887 385 891 386
rect 1239 390 1243 391
rect 1239 385 1243 386
rect 1279 390 1283 391
rect 1279 385 1283 386
rect 1303 390 1307 391
rect 1303 385 1307 386
rect 1343 390 1347 391
rect 1343 385 1347 386
rect 1399 390 1403 391
rect 1399 385 1403 386
rect 1447 390 1451 391
rect 1447 385 1451 386
rect 582 384 588 385
rect 582 380 583 384
rect 587 380 588 384
rect 582 379 588 380
rect 630 384 636 385
rect 630 380 631 384
rect 635 380 636 384
rect 630 379 636 380
rect 678 384 684 385
rect 678 380 679 384
rect 683 380 684 384
rect 678 379 684 380
rect 726 384 732 385
rect 726 380 727 384
rect 731 380 732 384
rect 726 379 732 380
rect 774 384 780 385
rect 774 380 775 384
rect 779 380 780 384
rect 774 379 780 380
rect 1240 378 1242 385
rect 1280 378 1282 385
rect 1446 384 1452 385
rect 1446 380 1447 384
rect 1451 380 1452 384
rect 1446 379 1452 380
rect 1238 377 1244 378
rect 566 375 572 376
rect 566 371 567 375
rect 571 371 572 375
rect 1238 373 1239 377
rect 1243 373 1244 377
rect 1238 372 1244 373
rect 1278 377 1284 378
rect 1278 373 1279 377
rect 1283 373 1284 377
rect 1278 372 1284 373
rect 566 370 572 371
rect 526 363 532 364
rect 526 359 527 363
rect 531 359 532 363
rect 526 358 532 359
rect 574 363 580 364
rect 574 359 575 363
rect 579 359 580 363
rect 574 358 580 359
rect 622 363 628 364
rect 622 359 623 363
rect 627 359 628 363
rect 622 358 628 359
rect 670 363 676 364
rect 670 359 671 363
rect 675 359 676 363
rect 670 358 676 359
rect 718 363 724 364
rect 718 359 719 363
rect 723 359 724 363
rect 718 358 724 359
rect 766 363 772 364
rect 766 359 767 363
rect 771 359 772 363
rect 766 358 772 359
rect 1238 360 1244 361
rect 486 337 492 338
rect 486 333 487 337
rect 491 333 492 337
rect 486 332 492 333
rect 466 327 472 328
rect 466 323 467 327
rect 471 323 472 327
rect 466 322 472 323
rect 488 319 490 332
rect 528 328 530 358
rect 534 337 540 338
rect 534 333 535 337
rect 539 333 540 337
rect 534 332 540 333
rect 526 327 532 328
rect 526 323 527 327
rect 531 323 532 327
rect 526 322 532 323
rect 536 319 538 332
rect 576 328 578 358
rect 582 337 588 338
rect 582 333 583 337
rect 587 333 588 337
rect 582 332 588 333
rect 574 327 580 328
rect 574 323 575 327
rect 579 323 580 327
rect 574 322 580 323
rect 584 319 586 332
rect 624 328 626 358
rect 630 337 636 338
rect 630 333 631 337
rect 635 333 636 337
rect 630 332 636 333
rect 622 327 628 328
rect 622 323 623 327
rect 627 323 628 327
rect 622 322 628 323
rect 610 319 616 320
rect 632 319 634 332
rect 672 328 674 358
rect 678 337 684 338
rect 678 333 679 337
rect 683 333 684 337
rect 678 332 684 333
rect 670 327 676 328
rect 670 323 671 327
rect 675 323 676 327
rect 670 322 676 323
rect 680 319 682 332
rect 720 328 722 358
rect 726 337 732 338
rect 726 333 727 337
rect 731 333 732 337
rect 726 332 732 333
rect 718 327 724 328
rect 718 323 719 327
rect 723 323 724 327
rect 718 322 724 323
rect 728 319 730 332
rect 768 328 770 358
rect 1238 356 1239 360
rect 1243 356 1244 360
rect 1238 355 1244 356
rect 1278 360 1284 361
rect 1278 356 1279 360
rect 1283 356 1284 360
rect 1278 355 1284 356
rect 774 337 780 338
rect 774 333 775 337
rect 779 333 780 337
rect 774 332 780 333
rect 766 327 772 328
rect 766 323 767 327
rect 771 323 772 327
rect 766 322 772 323
rect 776 319 778 332
rect 1240 319 1242 355
rect 1280 319 1282 355
rect 1446 337 1452 338
rect 1446 333 1447 337
rect 1451 333 1452 337
rect 1446 332 1452 333
rect 1448 319 1450 332
rect 1456 328 1458 406
rect 1462 400 1468 401
rect 1462 396 1463 400
rect 1467 396 1468 400
rect 1462 395 1468 396
rect 1526 400 1532 401
rect 1526 396 1527 400
rect 1531 396 1532 400
rect 1526 395 1532 396
rect 1590 400 1596 401
rect 1590 396 1591 400
rect 1595 396 1596 400
rect 1590 395 1596 396
rect 1464 391 1466 395
rect 1528 391 1530 395
rect 1592 391 1594 395
rect 1463 390 1467 391
rect 1463 385 1467 386
rect 1487 390 1491 391
rect 1487 385 1491 386
rect 1527 390 1531 391
rect 1527 385 1531 386
rect 1535 390 1539 391
rect 1535 385 1539 386
rect 1591 390 1595 391
rect 1591 385 1595 386
rect 1486 384 1492 385
rect 1486 380 1487 384
rect 1491 380 1492 384
rect 1486 379 1492 380
rect 1534 384 1540 385
rect 1534 380 1535 384
rect 1539 380 1540 384
rect 1534 379 1540 380
rect 1590 384 1596 385
rect 1590 380 1591 384
rect 1595 380 1596 384
rect 1590 379 1596 380
rect 1474 363 1480 364
rect 1474 359 1475 363
rect 1479 359 1480 363
rect 1474 358 1480 359
rect 1526 363 1532 364
rect 1526 359 1527 363
rect 1531 359 1532 363
rect 1526 358 1532 359
rect 1582 363 1588 364
rect 1582 359 1583 363
rect 1587 359 1588 363
rect 1582 358 1588 359
rect 1598 363 1604 364
rect 1598 359 1599 363
rect 1603 359 1604 363
rect 1598 358 1604 359
rect 1476 328 1478 358
rect 1486 337 1492 338
rect 1486 333 1487 337
rect 1491 333 1492 337
rect 1486 332 1492 333
rect 1454 327 1460 328
rect 1454 323 1455 327
rect 1459 323 1460 327
rect 1454 322 1460 323
rect 1474 327 1480 328
rect 1474 323 1475 327
rect 1479 323 1480 327
rect 1474 322 1480 323
rect 1488 319 1490 332
rect 1528 328 1530 358
rect 1534 337 1540 338
rect 1534 333 1535 337
rect 1539 333 1540 337
rect 1534 332 1540 333
rect 1526 327 1532 328
rect 1526 323 1527 327
rect 1531 323 1532 327
rect 1526 322 1532 323
rect 1536 319 1538 332
rect 1584 328 1586 358
rect 1590 337 1596 338
rect 1590 333 1591 337
rect 1595 333 1596 337
rect 1590 332 1596 333
rect 1582 327 1588 328
rect 1582 323 1583 327
rect 1587 323 1588 327
rect 1582 322 1588 323
rect 1592 319 1594 332
rect 1600 320 1602 358
rect 1656 328 1658 414
rect 1662 400 1668 401
rect 1662 396 1663 400
rect 1667 396 1668 400
rect 1662 395 1668 396
rect 1664 391 1666 395
rect 1663 390 1667 391
rect 1663 385 1667 386
rect 1662 384 1668 385
rect 1662 380 1663 384
rect 1667 380 1668 384
rect 1662 379 1668 380
rect 1716 372 1718 450
rect 1736 448 1738 457
rect 1762 455 1768 456
rect 1762 451 1763 455
rect 1767 451 1768 455
rect 1762 450 1768 451
rect 1734 447 1740 448
rect 1734 443 1735 447
rect 1739 443 1740 447
rect 1734 442 1740 443
rect 1764 420 1766 450
rect 1816 448 1818 457
rect 1842 455 1848 456
rect 1842 451 1843 455
rect 1847 451 1848 455
rect 1842 450 1848 451
rect 1814 447 1820 448
rect 1814 443 1815 447
rect 1819 443 1820 447
rect 1814 442 1820 443
rect 1844 420 1846 450
rect 1896 448 1898 457
rect 1922 455 1928 456
rect 1922 451 1923 455
rect 1927 451 1928 455
rect 1922 450 1928 451
rect 1894 447 1900 448
rect 1894 443 1895 447
rect 1899 443 1900 447
rect 1894 442 1900 443
rect 1924 420 1926 450
rect 1976 448 1978 457
rect 2056 448 2058 457
rect 2062 455 2068 456
rect 2062 451 2063 455
rect 2067 451 2068 455
rect 2062 450 2068 451
rect 2082 455 2088 456
rect 2082 451 2083 455
rect 2087 451 2088 455
rect 2082 450 2088 451
rect 1974 447 1980 448
rect 1974 443 1975 447
rect 1979 443 1980 447
rect 1974 442 1980 443
rect 2054 447 2060 448
rect 2054 443 2055 447
rect 2059 443 2060 447
rect 2054 442 2060 443
rect 1762 419 1768 420
rect 1762 415 1763 419
rect 1767 415 1768 419
rect 1762 414 1768 415
rect 1842 419 1848 420
rect 1842 415 1843 419
rect 1847 415 1848 419
rect 1842 414 1848 415
rect 1922 419 1928 420
rect 1922 415 1923 419
rect 1927 415 1928 419
rect 1922 414 1928 415
rect 1930 419 1936 420
rect 1930 415 1931 419
rect 1935 415 1936 419
rect 1930 414 1936 415
rect 1734 400 1740 401
rect 1734 396 1735 400
rect 1739 396 1740 400
rect 1734 395 1740 396
rect 1814 400 1820 401
rect 1814 396 1815 400
rect 1819 396 1820 400
rect 1814 395 1820 396
rect 1894 400 1900 401
rect 1894 396 1895 400
rect 1899 396 1900 400
rect 1894 395 1900 396
rect 1736 391 1738 395
rect 1816 391 1818 395
rect 1896 391 1898 395
rect 1735 390 1739 391
rect 1735 385 1739 386
rect 1815 390 1819 391
rect 1815 385 1819 386
rect 1895 390 1899 391
rect 1895 385 1899 386
rect 1734 384 1740 385
rect 1734 380 1735 384
rect 1739 380 1740 384
rect 1734 379 1740 380
rect 1814 384 1820 385
rect 1814 380 1815 384
rect 1819 380 1820 384
rect 1814 379 1820 380
rect 1894 384 1900 385
rect 1894 380 1895 384
rect 1899 380 1900 384
rect 1894 379 1900 380
rect 1714 371 1720 372
rect 1714 367 1715 371
rect 1719 367 1720 371
rect 1714 366 1720 367
rect 1726 363 1732 364
rect 1726 359 1727 363
rect 1731 359 1732 363
rect 1726 358 1732 359
rect 1806 363 1812 364
rect 1806 359 1807 363
rect 1811 359 1812 363
rect 1806 358 1812 359
rect 1822 363 1828 364
rect 1822 359 1823 363
rect 1827 359 1828 363
rect 1822 358 1828 359
rect 1662 337 1668 338
rect 1662 333 1663 337
rect 1667 333 1668 337
rect 1662 332 1668 333
rect 1654 327 1660 328
rect 1654 323 1655 327
rect 1659 323 1660 327
rect 1654 322 1660 323
rect 1598 319 1604 320
rect 1664 319 1666 332
rect 1728 328 1730 358
rect 1734 337 1740 338
rect 1734 333 1735 337
rect 1739 333 1740 337
rect 1734 332 1740 333
rect 1726 327 1732 328
rect 1726 323 1727 327
rect 1731 323 1732 327
rect 1726 322 1732 323
rect 1736 319 1738 332
rect 1808 328 1810 358
rect 1814 337 1820 338
rect 1814 333 1815 337
rect 1819 333 1820 337
rect 1814 332 1820 333
rect 1806 327 1812 328
rect 1806 323 1807 327
rect 1811 323 1812 327
rect 1806 322 1812 323
rect 1816 319 1818 332
rect 1824 320 1826 358
rect 1894 337 1900 338
rect 1894 333 1895 337
rect 1899 333 1900 337
rect 1894 332 1900 333
rect 1822 319 1828 320
rect 1896 319 1898 332
rect 1932 328 1934 414
rect 1974 400 1980 401
rect 1974 396 1975 400
rect 1979 396 1980 400
rect 1974 395 1980 396
rect 2054 400 2060 401
rect 2054 396 2055 400
rect 2059 396 2060 400
rect 2054 395 2060 396
rect 1976 391 1978 395
rect 2056 391 2058 395
rect 1967 390 1971 391
rect 1967 385 1971 386
rect 1975 390 1979 391
rect 1975 385 1979 386
rect 2039 390 2043 391
rect 2039 385 2043 386
rect 2055 390 2059 391
rect 2055 385 2059 386
rect 1966 384 1972 385
rect 1966 380 1967 384
rect 1971 380 1972 384
rect 1966 379 1972 380
rect 2038 384 2044 385
rect 2038 380 2039 384
rect 2043 380 2044 384
rect 2038 379 2044 380
rect 2064 364 2066 450
rect 2084 420 2086 450
rect 2136 448 2138 457
rect 2162 455 2168 456
rect 2162 451 2163 455
rect 2167 451 2168 455
rect 2162 450 2168 451
rect 2134 447 2140 448
rect 2134 443 2135 447
rect 2139 443 2140 447
rect 2134 442 2140 443
rect 2164 420 2166 450
rect 2176 420 2178 466
rect 2192 463 2194 476
rect 2280 472 2282 502
rect 2286 481 2292 482
rect 2286 477 2287 481
rect 2291 477 2292 481
rect 2286 476 2292 477
rect 2358 481 2364 482
rect 2358 477 2359 481
rect 2363 477 2364 481
rect 2358 476 2364 477
rect 2278 471 2284 472
rect 2278 467 2279 471
rect 2283 467 2284 471
rect 2278 466 2284 467
rect 2288 463 2290 476
rect 2360 463 2362 476
rect 2191 462 2195 463
rect 2191 457 2195 458
rect 2215 462 2219 463
rect 2215 457 2219 458
rect 2287 462 2291 463
rect 2287 457 2291 458
rect 2295 462 2299 463
rect 2295 457 2299 458
rect 2359 462 2363 463
rect 2359 457 2363 458
rect 2216 448 2218 457
rect 2296 448 2298 457
rect 2360 448 2362 457
rect 2368 456 2370 502
rect 2376 472 2378 554
rect 2406 547 2412 548
rect 2406 543 2407 547
rect 2411 543 2412 547
rect 2406 542 2412 543
rect 2408 535 2410 542
rect 2407 534 2411 535
rect 2407 529 2411 530
rect 2408 522 2410 529
rect 2406 521 2412 522
rect 2406 517 2407 521
rect 2411 517 2412 521
rect 2406 516 2412 517
rect 2406 504 2412 505
rect 2406 500 2407 504
rect 2411 500 2412 504
rect 2406 499 2412 500
rect 2374 471 2380 472
rect 2374 467 2375 471
rect 2379 467 2380 471
rect 2374 466 2380 467
rect 2408 463 2410 499
rect 2407 462 2411 463
rect 2407 457 2411 458
rect 2366 455 2372 456
rect 2366 451 2367 455
rect 2371 451 2372 455
rect 2366 450 2372 451
rect 2214 447 2220 448
rect 2214 443 2215 447
rect 2219 443 2220 447
rect 2214 442 2220 443
rect 2294 447 2300 448
rect 2294 443 2295 447
rect 2299 443 2300 447
rect 2294 442 2300 443
rect 2358 447 2364 448
rect 2358 443 2359 447
rect 2363 443 2364 447
rect 2358 442 2364 443
rect 2408 425 2410 457
rect 2406 424 2412 425
rect 2406 420 2407 424
rect 2411 420 2412 424
rect 2082 419 2088 420
rect 2082 415 2083 419
rect 2087 415 2088 419
rect 2082 414 2088 415
rect 2162 419 2168 420
rect 2162 415 2163 419
rect 2167 415 2168 419
rect 2162 414 2168 415
rect 2174 419 2180 420
rect 2174 415 2175 419
rect 2179 415 2180 419
rect 2174 414 2180 415
rect 2350 419 2356 420
rect 2406 419 2412 420
rect 2350 415 2351 419
rect 2355 415 2356 419
rect 2350 414 2356 415
rect 2134 400 2140 401
rect 2134 396 2135 400
rect 2139 396 2140 400
rect 2134 395 2140 396
rect 2214 400 2220 401
rect 2214 396 2215 400
rect 2219 396 2220 400
rect 2214 395 2220 396
rect 2294 400 2300 401
rect 2294 396 2295 400
rect 2299 396 2300 400
rect 2294 395 2300 396
rect 2136 391 2138 395
rect 2216 391 2218 395
rect 2296 391 2298 395
rect 2111 390 2115 391
rect 2111 385 2115 386
rect 2135 390 2139 391
rect 2135 385 2139 386
rect 2175 390 2179 391
rect 2175 385 2179 386
rect 2215 390 2219 391
rect 2215 385 2219 386
rect 2239 390 2243 391
rect 2239 385 2243 386
rect 2295 390 2299 391
rect 2295 385 2299 386
rect 2303 390 2307 391
rect 2303 385 2307 386
rect 2110 384 2116 385
rect 2110 380 2111 384
rect 2115 380 2116 384
rect 2110 379 2116 380
rect 2174 384 2180 385
rect 2174 380 2175 384
rect 2179 380 2180 384
rect 2174 379 2180 380
rect 2238 384 2244 385
rect 2238 380 2239 384
rect 2243 380 2244 384
rect 2238 379 2244 380
rect 2302 384 2308 385
rect 2302 380 2303 384
rect 2307 380 2308 384
rect 2302 379 2308 380
rect 2030 363 2036 364
rect 2030 359 2031 363
rect 2035 359 2036 363
rect 2030 358 2036 359
rect 2062 363 2068 364
rect 2062 359 2063 363
rect 2067 359 2068 363
rect 2062 358 2068 359
rect 2338 363 2344 364
rect 2338 359 2339 363
rect 2343 359 2344 363
rect 2338 358 2344 359
rect 1974 355 1980 356
rect 1974 351 1975 355
rect 1979 351 1980 355
rect 1974 350 1980 351
rect 1966 337 1972 338
rect 1966 333 1967 337
rect 1971 333 1972 337
rect 1966 332 1972 333
rect 1930 327 1936 328
rect 1930 323 1931 327
rect 1935 323 1936 327
rect 1930 322 1936 323
rect 1968 319 1970 332
rect 1976 328 1978 350
rect 2032 328 2034 358
rect 2038 337 2044 338
rect 2038 333 2039 337
rect 2043 333 2044 337
rect 2038 332 2044 333
rect 2110 337 2116 338
rect 2110 333 2111 337
rect 2115 333 2116 337
rect 2110 332 2116 333
rect 2174 337 2180 338
rect 2174 333 2175 337
rect 2179 333 2180 337
rect 2174 332 2180 333
rect 2238 337 2244 338
rect 2238 333 2239 337
rect 2243 333 2244 337
rect 2238 332 2244 333
rect 2302 337 2308 338
rect 2302 333 2303 337
rect 2307 333 2308 337
rect 2302 332 2308 333
rect 1974 327 1980 328
rect 1974 323 1975 327
rect 1979 323 1980 327
rect 1974 322 1980 323
rect 2030 327 2036 328
rect 2030 323 2031 327
rect 2035 323 2036 327
rect 2030 322 2036 323
rect 2040 319 2042 332
rect 2112 319 2114 332
rect 2176 319 2178 332
rect 2240 319 2242 332
rect 2282 327 2288 328
rect 2282 323 2283 327
rect 2287 323 2288 327
rect 2282 322 2288 323
rect 343 318 347 319
rect 343 313 347 314
rect 391 318 395 319
rect 391 313 395 314
rect 439 318 443 319
rect 439 313 443 314
rect 447 318 451 319
rect 447 313 451 314
rect 487 318 491 319
rect 487 313 491 314
rect 503 318 507 319
rect 503 313 507 314
rect 535 318 539 319
rect 535 313 539 314
rect 551 318 555 319
rect 551 313 555 314
rect 583 318 587 319
rect 583 313 587 314
rect 591 318 595 319
rect 610 315 611 319
rect 615 315 616 319
rect 610 314 616 315
rect 631 318 635 319
rect 591 313 595 314
rect 334 311 340 312
rect 334 307 335 311
rect 339 307 340 311
rect 334 306 340 307
rect 354 311 360 312
rect 354 307 355 311
rect 359 307 360 311
rect 354 306 360 307
rect 326 303 332 304
rect 326 299 327 303
rect 331 299 332 303
rect 326 298 332 299
rect 356 276 358 306
rect 392 304 394 313
rect 418 311 424 312
rect 418 307 419 311
rect 423 307 424 311
rect 418 306 424 307
rect 390 303 396 304
rect 390 299 391 303
rect 395 299 396 303
rect 390 298 396 299
rect 420 276 422 306
rect 448 304 450 313
rect 474 311 480 312
rect 474 307 475 311
rect 479 307 480 311
rect 474 306 480 307
rect 446 303 452 304
rect 446 299 447 303
rect 451 299 452 303
rect 446 298 452 299
rect 476 276 478 306
rect 504 304 506 313
rect 552 304 554 313
rect 592 304 594 313
rect 502 303 508 304
rect 502 299 503 303
rect 507 299 508 303
rect 502 298 508 299
rect 550 303 556 304
rect 550 299 551 303
rect 555 299 556 303
rect 550 298 556 299
rect 590 303 596 304
rect 590 299 591 303
rect 595 299 596 303
rect 590 298 596 299
rect 612 276 614 314
rect 631 313 635 314
rect 679 318 683 319
rect 679 313 683 314
rect 727 318 731 319
rect 727 313 731 314
rect 775 318 779 319
rect 775 313 779 314
rect 823 318 827 319
rect 823 313 827 314
rect 871 318 875 319
rect 871 313 875 314
rect 919 318 923 319
rect 919 313 923 314
rect 1239 318 1243 319
rect 1239 313 1243 314
rect 1279 318 1283 319
rect 1279 313 1283 314
rect 1447 318 1451 319
rect 1447 313 1451 314
rect 1487 318 1491 319
rect 1487 313 1491 314
rect 1495 318 1499 319
rect 1495 313 1499 314
rect 1535 318 1539 319
rect 1535 313 1539 314
rect 1575 318 1579 319
rect 1575 313 1579 314
rect 1591 318 1595 319
rect 1598 315 1599 319
rect 1603 315 1604 319
rect 1598 314 1604 315
rect 1615 318 1619 319
rect 1591 313 1595 314
rect 1615 313 1619 314
rect 1655 318 1659 319
rect 1655 313 1659 314
rect 1663 318 1667 319
rect 1663 313 1667 314
rect 1695 318 1699 319
rect 1695 313 1699 314
rect 1735 318 1739 319
rect 1735 313 1739 314
rect 1743 318 1747 319
rect 1743 313 1747 314
rect 1799 318 1803 319
rect 1799 313 1803 314
rect 1815 318 1819 319
rect 1822 315 1823 319
rect 1827 315 1828 319
rect 1822 314 1828 315
rect 1863 318 1867 319
rect 1815 313 1819 314
rect 1863 313 1867 314
rect 1895 318 1899 319
rect 1895 313 1899 314
rect 1935 318 1939 319
rect 1935 313 1939 314
rect 1967 318 1971 319
rect 1967 313 1971 314
rect 2007 318 2011 319
rect 2007 313 2011 314
rect 2039 318 2043 319
rect 2039 313 2043 314
rect 2071 318 2075 319
rect 2071 313 2075 314
rect 2111 318 2115 319
rect 2111 313 2115 314
rect 2135 318 2139 319
rect 2135 313 2139 314
rect 2175 318 2179 319
rect 2175 313 2179 314
rect 2191 318 2195 319
rect 2191 313 2195 314
rect 2239 318 2243 319
rect 2239 313 2243 314
rect 2255 318 2259 319
rect 2255 313 2259 314
rect 618 311 624 312
rect 618 307 619 311
rect 623 307 624 311
rect 618 306 624 307
rect 162 275 168 276
rect 162 271 163 275
rect 167 271 168 275
rect 162 270 168 271
rect 210 275 216 276
rect 210 271 211 275
rect 215 271 216 275
rect 210 270 216 271
rect 278 275 284 276
rect 278 271 279 275
rect 283 271 284 275
rect 278 270 284 271
rect 354 275 360 276
rect 354 271 355 275
rect 359 271 360 275
rect 354 270 360 271
rect 418 275 424 276
rect 418 271 419 275
rect 423 271 424 275
rect 418 270 424 271
rect 474 275 480 276
rect 474 271 475 275
rect 479 271 480 275
rect 474 270 480 271
rect 566 275 572 276
rect 566 271 567 275
rect 571 271 572 275
rect 566 270 572 271
rect 610 275 616 276
rect 610 271 611 275
rect 615 271 616 275
rect 620 275 622 306
rect 632 304 634 313
rect 666 311 672 312
rect 666 307 667 311
rect 671 307 672 311
rect 666 306 672 307
rect 630 303 636 304
rect 630 299 631 303
rect 635 299 636 303
rect 630 298 636 299
rect 668 276 670 306
rect 680 304 682 313
rect 714 311 720 312
rect 714 307 715 311
rect 719 307 720 311
rect 714 306 720 307
rect 678 303 684 304
rect 678 299 679 303
rect 683 299 684 303
rect 678 298 684 299
rect 716 276 718 306
rect 728 304 730 313
rect 762 311 768 312
rect 762 307 763 311
rect 767 307 768 311
rect 762 306 768 307
rect 726 303 732 304
rect 726 299 727 303
rect 731 299 732 303
rect 726 298 732 299
rect 764 276 766 306
rect 776 304 778 313
rect 806 311 812 312
rect 806 307 807 311
rect 811 307 812 311
rect 806 306 812 307
rect 814 311 820 312
rect 814 307 815 311
rect 819 307 820 311
rect 814 306 820 307
rect 774 303 780 304
rect 774 299 775 303
rect 779 299 780 303
rect 774 298 780 299
rect 808 284 810 306
rect 806 283 812 284
rect 806 279 807 283
rect 811 279 812 283
rect 806 278 812 279
rect 626 275 632 276
rect 620 273 627 275
rect 610 270 616 271
rect 626 271 627 273
rect 631 271 632 275
rect 626 270 632 271
rect 666 275 672 276
rect 666 271 667 275
rect 671 271 672 275
rect 666 270 672 271
rect 714 275 720 276
rect 714 271 715 275
rect 719 271 720 275
rect 714 270 720 271
rect 762 275 768 276
rect 762 271 763 275
rect 767 271 768 275
rect 762 270 768 271
rect 182 256 188 257
rect 182 252 183 256
rect 187 252 188 256
rect 182 251 188 252
rect 254 256 260 257
rect 254 252 255 256
rect 259 252 260 256
rect 254 251 260 252
rect 326 256 332 257
rect 326 252 327 256
rect 331 252 332 256
rect 326 251 332 252
rect 390 256 396 257
rect 390 252 391 256
rect 395 252 396 256
rect 390 251 396 252
rect 446 256 452 257
rect 446 252 447 256
rect 451 252 452 256
rect 446 251 452 252
rect 502 256 508 257
rect 502 252 503 256
rect 507 252 508 256
rect 502 251 508 252
rect 550 256 556 257
rect 550 252 551 256
rect 555 252 556 256
rect 550 251 556 252
rect 184 243 186 251
rect 256 243 258 251
rect 328 243 330 251
rect 392 243 394 251
rect 448 243 450 251
rect 504 243 506 251
rect 552 243 554 251
rect 175 242 179 243
rect 175 237 179 238
rect 183 242 187 243
rect 183 237 187 238
rect 247 242 251 243
rect 247 237 251 238
rect 255 242 259 243
rect 255 237 259 238
rect 327 242 331 243
rect 327 237 331 238
rect 391 242 395 243
rect 391 237 395 238
rect 415 242 419 243
rect 415 237 419 238
rect 447 242 451 243
rect 447 237 451 238
rect 495 242 499 243
rect 495 237 499 238
rect 503 242 507 243
rect 503 237 507 238
rect 551 242 555 243
rect 551 237 555 238
rect 174 236 180 237
rect 174 232 175 236
rect 179 232 180 236
rect 174 231 180 232
rect 246 236 252 237
rect 246 232 247 236
rect 251 232 252 236
rect 246 231 252 232
rect 326 236 332 237
rect 326 232 327 236
rect 331 232 332 236
rect 326 231 332 232
rect 414 236 420 237
rect 414 232 415 236
rect 419 232 420 236
rect 414 231 420 232
rect 494 236 500 237
rect 494 232 495 236
rect 499 232 500 236
rect 494 231 500 232
rect 154 215 160 216
rect 110 212 116 213
rect 110 208 111 212
rect 115 208 116 212
rect 154 211 155 215
rect 159 211 160 215
rect 170 215 176 216
rect 170 214 171 215
rect 154 210 160 211
rect 164 212 171 214
rect 110 207 116 208
rect 112 155 114 207
rect 134 189 140 190
rect 134 185 135 189
rect 139 185 140 189
rect 134 184 140 185
rect 136 155 138 184
rect 164 180 166 212
rect 170 211 171 212
rect 175 211 176 215
rect 170 210 176 211
rect 318 215 324 216
rect 318 211 319 215
rect 323 211 324 215
rect 318 210 324 211
rect 486 215 492 216
rect 486 211 487 215
rect 491 211 492 215
rect 486 210 492 211
rect 518 215 524 216
rect 518 211 519 215
rect 523 211 524 215
rect 518 210 524 211
rect 182 207 188 208
rect 182 203 183 207
rect 187 203 188 207
rect 182 202 188 203
rect 174 189 180 190
rect 174 185 175 189
rect 179 185 180 189
rect 174 184 180 185
rect 162 179 168 180
rect 162 175 163 179
rect 167 175 168 179
rect 162 174 168 175
rect 176 155 178 184
rect 184 180 186 202
rect 246 189 252 190
rect 246 185 247 189
rect 251 185 252 189
rect 246 184 252 185
rect 182 179 188 180
rect 182 175 183 179
rect 187 175 188 179
rect 182 174 188 175
rect 238 179 244 180
rect 238 175 239 179
rect 243 175 244 179
rect 238 174 244 175
rect 111 154 115 155
rect 111 149 115 150
rect 135 154 139 155
rect 135 149 139 150
rect 175 154 179 155
rect 175 149 179 150
rect 215 154 219 155
rect 215 149 219 150
rect 112 117 114 149
rect 136 140 138 149
rect 150 147 156 148
rect 150 143 151 147
rect 155 143 156 147
rect 150 142 156 143
rect 158 147 164 148
rect 158 143 159 147
rect 163 143 164 147
rect 158 142 164 143
rect 134 139 140 140
rect 134 135 135 139
rect 139 135 140 139
rect 134 134 140 135
rect 152 120 154 142
rect 150 119 156 120
rect 110 116 116 117
rect 110 112 111 116
rect 115 112 116 116
rect 150 115 151 119
rect 155 115 156 119
rect 150 114 156 115
rect 160 112 162 142
rect 176 140 178 149
rect 202 147 208 148
rect 202 143 203 147
rect 207 143 208 147
rect 202 142 208 143
rect 174 139 180 140
rect 174 135 175 139
rect 179 135 180 139
rect 174 134 180 135
rect 204 112 206 142
rect 216 140 218 149
rect 214 139 220 140
rect 214 135 215 139
rect 219 135 220 139
rect 214 134 220 135
rect 240 112 242 174
rect 248 155 250 184
rect 320 180 322 210
rect 422 207 428 208
rect 422 203 423 207
rect 427 203 428 207
rect 422 202 428 203
rect 326 189 332 190
rect 326 185 327 189
rect 331 185 332 189
rect 326 184 332 185
rect 414 189 420 190
rect 414 185 415 189
rect 419 185 420 189
rect 414 184 420 185
rect 318 179 324 180
rect 318 175 319 179
rect 323 175 324 179
rect 318 174 324 175
rect 328 155 330 184
rect 416 155 418 184
rect 424 180 426 202
rect 488 180 490 210
rect 494 189 500 190
rect 494 185 495 189
rect 499 185 500 189
rect 494 184 500 185
rect 422 179 428 180
rect 422 175 423 179
rect 427 175 428 179
rect 422 174 428 175
rect 486 179 492 180
rect 486 175 487 179
rect 491 175 492 179
rect 486 174 492 175
rect 496 155 498 184
rect 247 154 251 155
rect 247 149 251 150
rect 255 154 259 155
rect 255 149 259 150
rect 295 154 299 155
rect 295 149 299 150
rect 327 154 331 155
rect 327 149 331 150
rect 335 154 339 155
rect 335 149 339 150
rect 375 154 379 155
rect 375 149 379 150
rect 415 154 419 155
rect 415 149 419 150
rect 423 154 427 155
rect 423 149 427 150
rect 471 154 475 155
rect 471 149 475 150
rect 495 154 499 155
rect 495 149 499 150
rect 256 140 258 149
rect 282 147 288 148
rect 282 143 283 147
rect 287 143 288 147
rect 282 142 288 143
rect 254 139 260 140
rect 254 135 255 139
rect 259 135 260 139
rect 254 134 260 135
rect 284 120 286 142
rect 296 140 298 149
rect 318 147 324 148
rect 318 143 319 147
rect 323 143 324 147
rect 318 142 324 143
rect 294 139 300 140
rect 294 135 295 139
rect 299 135 300 139
rect 294 134 300 135
rect 320 120 322 142
rect 336 140 338 149
rect 362 147 368 148
rect 362 143 363 147
rect 367 143 368 147
rect 362 142 368 143
rect 334 139 340 140
rect 334 135 335 139
rect 339 135 340 139
rect 334 134 340 135
rect 364 120 366 142
rect 376 140 378 149
rect 424 140 426 149
rect 458 147 464 148
rect 458 143 459 147
rect 463 143 464 147
rect 458 142 464 143
rect 374 139 380 140
rect 374 135 375 139
rect 379 135 380 139
rect 374 134 380 135
rect 422 139 428 140
rect 422 135 423 139
rect 427 135 428 139
rect 422 134 428 135
rect 282 119 288 120
rect 282 115 283 119
rect 287 115 288 119
rect 282 114 288 115
rect 318 119 324 120
rect 318 115 319 119
rect 323 115 324 119
rect 318 114 324 115
rect 362 119 368 120
rect 362 115 363 119
rect 367 115 368 119
rect 362 114 368 115
rect 460 112 462 142
rect 472 140 474 149
rect 520 148 522 210
rect 568 180 570 270
rect 590 256 596 257
rect 590 252 591 256
rect 595 252 596 256
rect 590 251 596 252
rect 630 256 636 257
rect 630 252 631 256
rect 635 252 636 256
rect 630 251 636 252
rect 678 256 684 257
rect 678 252 679 256
rect 683 252 684 256
rect 678 251 684 252
rect 726 256 732 257
rect 726 252 727 256
rect 731 252 732 256
rect 726 251 732 252
rect 774 256 780 257
rect 774 252 775 256
rect 779 252 780 256
rect 774 251 780 252
rect 592 243 594 251
rect 632 243 634 251
rect 680 243 682 251
rect 728 243 730 251
rect 776 243 778 251
rect 575 242 579 243
rect 575 237 579 238
rect 591 242 595 243
rect 591 237 595 238
rect 631 242 635 243
rect 631 237 635 238
rect 655 242 659 243
rect 655 237 659 238
rect 679 242 683 243
rect 679 237 683 238
rect 727 242 731 243
rect 727 237 731 238
rect 775 242 779 243
rect 775 237 779 238
rect 791 242 795 243
rect 791 237 795 238
rect 574 236 580 237
rect 574 232 575 236
rect 579 232 580 236
rect 574 231 580 232
rect 654 236 660 237
rect 654 232 655 236
rect 659 232 660 236
rect 654 231 660 232
rect 726 236 732 237
rect 726 232 727 236
rect 731 232 732 236
rect 726 231 732 232
rect 790 236 796 237
rect 790 232 791 236
rect 795 232 796 236
rect 790 231 796 232
rect 816 216 818 306
rect 824 304 826 313
rect 858 311 864 312
rect 858 307 859 311
rect 863 307 864 311
rect 858 306 864 307
rect 822 303 828 304
rect 822 299 823 303
rect 827 299 828 303
rect 822 298 828 299
rect 860 276 862 306
rect 872 304 874 313
rect 906 311 912 312
rect 906 307 907 311
rect 911 307 912 311
rect 906 306 912 307
rect 870 303 876 304
rect 870 299 871 303
rect 875 299 876 303
rect 870 298 876 299
rect 908 276 910 306
rect 920 304 922 313
rect 918 303 924 304
rect 918 299 919 303
rect 923 299 924 303
rect 918 298 924 299
rect 1240 281 1242 313
rect 1280 281 1282 313
rect 1496 304 1498 313
rect 1522 311 1528 312
rect 1522 307 1523 311
rect 1527 307 1528 311
rect 1522 306 1528 307
rect 1494 303 1500 304
rect 1494 299 1495 303
rect 1499 299 1500 303
rect 1494 298 1500 299
rect 1238 280 1244 281
rect 1238 276 1239 280
rect 1243 276 1244 280
rect 858 275 864 276
rect 858 271 859 275
rect 863 271 864 275
rect 858 270 864 271
rect 906 275 912 276
rect 1238 275 1244 276
rect 1278 280 1284 281
rect 1278 276 1279 280
rect 1283 276 1284 280
rect 1524 276 1526 306
rect 1536 304 1538 313
rect 1562 311 1568 312
rect 1562 307 1563 311
rect 1567 307 1568 311
rect 1562 306 1568 307
rect 1534 303 1540 304
rect 1534 299 1535 303
rect 1539 299 1540 303
rect 1534 298 1540 299
rect 1564 276 1566 306
rect 1576 304 1578 313
rect 1602 311 1608 312
rect 1602 307 1603 311
rect 1607 307 1608 311
rect 1602 306 1608 307
rect 1574 303 1580 304
rect 1574 299 1575 303
rect 1579 299 1580 303
rect 1574 298 1580 299
rect 1604 276 1606 306
rect 1616 304 1618 313
rect 1642 311 1648 312
rect 1642 307 1643 311
rect 1647 307 1648 311
rect 1642 306 1648 307
rect 1614 303 1620 304
rect 1614 299 1615 303
rect 1619 299 1620 303
rect 1614 298 1620 299
rect 1644 276 1646 306
rect 1656 304 1658 313
rect 1682 311 1688 312
rect 1682 307 1683 311
rect 1687 307 1688 311
rect 1682 306 1688 307
rect 1654 303 1660 304
rect 1654 299 1655 303
rect 1659 299 1660 303
rect 1654 298 1660 299
rect 1684 276 1686 306
rect 1696 304 1698 313
rect 1722 311 1728 312
rect 1722 307 1723 311
rect 1727 307 1728 311
rect 1722 306 1728 307
rect 1694 303 1700 304
rect 1694 299 1695 303
rect 1699 299 1700 303
rect 1694 298 1700 299
rect 1724 276 1726 306
rect 1744 304 1746 313
rect 1800 304 1802 313
rect 1826 311 1832 312
rect 1826 307 1827 311
rect 1831 307 1832 311
rect 1826 306 1832 307
rect 1742 303 1748 304
rect 1742 299 1743 303
rect 1747 299 1748 303
rect 1742 298 1748 299
rect 1798 303 1804 304
rect 1798 299 1799 303
rect 1803 299 1804 303
rect 1798 298 1804 299
rect 1828 276 1830 306
rect 1864 304 1866 313
rect 1936 304 1938 313
rect 1974 311 1980 312
rect 1974 307 1975 311
rect 1979 307 1980 311
rect 1974 306 1980 307
rect 1862 303 1868 304
rect 1862 299 1863 303
rect 1867 299 1868 303
rect 1862 298 1868 299
rect 1934 303 1940 304
rect 1934 299 1935 303
rect 1939 299 1940 303
rect 1934 298 1940 299
rect 1976 276 1978 306
rect 2008 304 2010 313
rect 2072 304 2074 313
rect 2090 311 2096 312
rect 2090 307 2091 311
rect 2095 307 2096 311
rect 2090 306 2096 307
rect 2098 311 2104 312
rect 2098 307 2099 311
rect 2103 307 2104 311
rect 2098 306 2104 307
rect 2006 303 2012 304
rect 2006 299 2007 303
rect 2011 299 2012 303
rect 2006 298 2012 299
rect 2070 303 2076 304
rect 2070 299 2071 303
rect 2075 299 2076 303
rect 2070 298 2076 299
rect 1278 275 1284 276
rect 1522 275 1528 276
rect 906 271 907 275
rect 911 271 912 275
rect 906 270 912 271
rect 1522 271 1523 275
rect 1527 271 1528 275
rect 1522 270 1528 271
rect 1562 275 1568 276
rect 1562 271 1563 275
rect 1567 271 1568 275
rect 1562 270 1568 271
rect 1602 275 1608 276
rect 1602 271 1603 275
rect 1607 271 1608 275
rect 1602 270 1608 271
rect 1642 275 1648 276
rect 1642 271 1643 275
rect 1647 271 1648 275
rect 1642 270 1648 271
rect 1682 275 1688 276
rect 1682 271 1683 275
rect 1687 271 1688 275
rect 1682 270 1688 271
rect 1722 275 1728 276
rect 1722 271 1723 275
rect 1727 271 1728 275
rect 1722 270 1728 271
rect 1826 275 1832 276
rect 1826 271 1827 275
rect 1831 271 1832 275
rect 1826 270 1832 271
rect 1974 275 1980 276
rect 1974 271 1975 275
rect 1979 271 1980 275
rect 1974 270 1980 271
rect 1982 275 1988 276
rect 1982 271 1983 275
rect 1987 271 1988 275
rect 1982 270 1988 271
rect 1710 267 1716 268
rect 1238 263 1244 264
rect 1238 259 1239 263
rect 1243 259 1244 263
rect 1238 258 1244 259
rect 1278 263 1284 264
rect 1278 259 1279 263
rect 1283 259 1284 263
rect 1710 263 1711 267
rect 1715 263 1716 267
rect 1710 262 1716 263
rect 1278 258 1284 259
rect 822 256 828 257
rect 822 252 823 256
rect 827 252 828 256
rect 822 251 828 252
rect 870 256 876 257
rect 870 252 871 256
rect 875 252 876 256
rect 870 251 876 252
rect 918 256 924 257
rect 918 252 919 256
rect 923 252 924 256
rect 918 251 924 252
rect 824 243 826 251
rect 872 243 874 251
rect 920 243 922 251
rect 1240 243 1242 258
rect 1280 247 1282 258
rect 1494 256 1500 257
rect 1494 252 1495 256
rect 1499 252 1500 256
rect 1494 251 1500 252
rect 1534 256 1540 257
rect 1534 252 1535 256
rect 1539 252 1540 256
rect 1534 251 1540 252
rect 1574 256 1580 257
rect 1574 252 1575 256
rect 1579 252 1580 256
rect 1574 251 1580 252
rect 1614 256 1620 257
rect 1614 252 1615 256
rect 1619 252 1620 256
rect 1614 251 1620 252
rect 1654 256 1660 257
rect 1654 252 1655 256
rect 1659 252 1660 256
rect 1654 251 1660 252
rect 1694 256 1700 257
rect 1694 252 1695 256
rect 1699 252 1700 256
rect 1694 251 1700 252
rect 1496 247 1498 251
rect 1536 247 1538 251
rect 1576 247 1578 251
rect 1616 247 1618 251
rect 1656 247 1658 251
rect 1696 247 1698 251
rect 1279 246 1283 247
rect 823 242 827 243
rect 823 237 827 238
rect 847 242 851 243
rect 847 237 851 238
rect 871 242 875 243
rect 871 237 875 238
rect 903 242 907 243
rect 903 237 907 238
rect 919 242 923 243
rect 919 237 923 238
rect 959 242 963 243
rect 959 237 963 238
rect 1023 242 1027 243
rect 1023 237 1027 238
rect 1239 242 1243 243
rect 1279 241 1283 242
rect 1367 246 1371 247
rect 1367 241 1371 242
rect 1407 246 1411 247
rect 1407 241 1411 242
rect 1447 246 1451 247
rect 1447 241 1451 242
rect 1495 246 1499 247
rect 1495 241 1499 242
rect 1535 246 1539 247
rect 1535 241 1539 242
rect 1551 246 1555 247
rect 1551 241 1555 242
rect 1575 246 1579 247
rect 1575 241 1579 242
rect 1607 246 1611 247
rect 1607 241 1611 242
rect 1615 246 1619 247
rect 1615 241 1619 242
rect 1655 246 1659 247
rect 1655 241 1659 242
rect 1671 246 1675 247
rect 1671 241 1675 242
rect 1695 246 1699 247
rect 1695 241 1699 242
rect 1239 237 1243 238
rect 846 236 852 237
rect 846 232 847 236
rect 851 232 852 236
rect 846 231 852 232
rect 902 236 908 237
rect 902 232 903 236
rect 907 232 908 236
rect 902 231 908 232
rect 958 236 964 237
rect 958 232 959 236
rect 963 232 964 236
rect 958 231 964 232
rect 1022 236 1028 237
rect 1022 232 1023 236
rect 1027 232 1028 236
rect 1022 231 1028 232
rect 1240 230 1242 237
rect 1280 234 1282 241
rect 1366 240 1372 241
rect 1366 236 1367 240
rect 1371 236 1372 240
rect 1366 235 1372 236
rect 1406 240 1412 241
rect 1406 236 1407 240
rect 1411 236 1412 240
rect 1406 235 1412 236
rect 1446 240 1452 241
rect 1446 236 1447 240
rect 1451 236 1452 240
rect 1446 235 1452 236
rect 1494 240 1500 241
rect 1494 236 1495 240
rect 1499 236 1500 240
rect 1494 235 1500 236
rect 1550 240 1556 241
rect 1550 236 1551 240
rect 1555 236 1556 240
rect 1550 235 1556 236
rect 1606 240 1612 241
rect 1606 236 1607 240
rect 1611 236 1612 240
rect 1606 235 1612 236
rect 1670 240 1676 241
rect 1670 236 1671 240
rect 1675 236 1676 240
rect 1670 235 1676 236
rect 1278 233 1284 234
rect 1238 229 1244 230
rect 1238 225 1239 229
rect 1243 225 1244 229
rect 1278 229 1279 233
rect 1283 229 1284 233
rect 1278 228 1284 229
rect 1238 224 1244 225
rect 1394 219 1400 220
rect 1278 216 1284 217
rect 718 215 724 216
rect 718 211 719 215
rect 723 211 724 215
rect 718 210 724 211
rect 782 215 788 216
rect 782 211 783 215
rect 787 211 788 215
rect 782 210 788 211
rect 814 215 820 216
rect 814 211 815 215
rect 819 211 820 215
rect 814 210 820 211
rect 942 215 948 216
rect 942 211 943 215
rect 947 211 948 215
rect 942 210 948 211
rect 1014 215 1020 216
rect 1014 211 1015 215
rect 1019 211 1020 215
rect 1014 210 1020 211
rect 1238 212 1244 213
rect 662 207 668 208
rect 662 203 663 207
rect 667 203 668 207
rect 662 202 668 203
rect 574 189 580 190
rect 574 185 575 189
rect 579 185 580 189
rect 574 184 580 185
rect 654 189 660 190
rect 654 185 655 189
rect 659 185 660 189
rect 654 184 660 185
rect 566 179 572 180
rect 566 175 567 179
rect 571 175 572 179
rect 566 174 572 175
rect 576 155 578 184
rect 656 155 658 184
rect 664 180 666 202
rect 720 180 722 210
rect 726 189 732 190
rect 726 185 727 189
rect 731 185 732 189
rect 726 184 732 185
rect 662 179 668 180
rect 662 175 663 179
rect 667 175 668 179
rect 662 174 668 175
rect 718 179 724 180
rect 718 175 719 179
rect 723 175 724 179
rect 718 174 724 175
rect 728 155 730 184
rect 784 180 786 210
rect 854 207 860 208
rect 854 203 855 207
rect 859 203 860 207
rect 854 202 860 203
rect 790 189 796 190
rect 790 185 791 189
rect 795 185 796 189
rect 790 184 796 185
rect 846 189 852 190
rect 846 185 847 189
rect 851 185 852 189
rect 846 184 852 185
rect 782 179 788 180
rect 782 175 783 179
rect 787 175 788 179
rect 782 174 788 175
rect 750 171 756 172
rect 750 167 751 171
rect 755 167 756 171
rect 750 166 756 167
rect 527 154 531 155
rect 527 149 531 150
rect 575 154 579 155
rect 575 149 579 150
rect 583 154 587 155
rect 583 149 587 150
rect 631 154 635 155
rect 631 149 635 150
rect 655 154 659 155
rect 655 149 659 150
rect 679 154 683 155
rect 679 149 683 150
rect 727 154 731 155
rect 727 149 731 150
rect 510 147 516 148
rect 510 143 511 147
rect 515 143 516 147
rect 510 142 516 143
rect 518 147 524 148
rect 518 143 519 147
rect 523 143 524 147
rect 518 142 524 143
rect 470 139 476 140
rect 470 135 471 139
rect 475 135 476 139
rect 470 134 476 135
rect 512 120 514 142
rect 528 140 530 149
rect 554 147 560 148
rect 554 143 555 147
rect 559 143 560 147
rect 554 142 560 143
rect 526 139 532 140
rect 526 135 527 139
rect 531 135 532 139
rect 526 134 532 135
rect 510 119 516 120
rect 510 115 511 119
rect 515 115 516 119
rect 510 114 516 115
rect 556 112 558 142
rect 584 140 586 149
rect 632 140 634 149
rect 646 147 652 148
rect 646 143 647 147
rect 651 143 652 147
rect 646 142 652 143
rect 582 139 588 140
rect 582 135 583 139
rect 587 135 588 139
rect 582 134 588 135
rect 630 139 636 140
rect 630 135 631 139
rect 635 135 636 139
rect 630 134 636 135
rect 648 124 650 142
rect 680 140 682 149
rect 706 147 712 148
rect 706 143 707 147
rect 711 143 712 147
rect 706 142 712 143
rect 678 139 684 140
rect 678 135 679 139
rect 683 135 684 139
rect 678 134 684 135
rect 646 123 652 124
rect 646 119 647 123
rect 651 119 652 123
rect 646 118 652 119
rect 708 112 710 142
rect 728 140 730 149
rect 726 139 732 140
rect 726 135 727 139
rect 731 135 732 139
rect 726 134 732 135
rect 752 112 754 166
rect 792 155 794 184
rect 848 155 850 184
rect 856 180 858 202
rect 902 189 908 190
rect 902 185 903 189
rect 907 185 908 189
rect 902 184 908 185
rect 854 179 860 180
rect 854 175 855 179
rect 859 175 860 179
rect 854 174 860 175
rect 904 155 906 184
rect 944 180 946 210
rect 958 189 964 190
rect 958 185 959 189
rect 963 185 964 189
rect 958 184 964 185
rect 942 179 948 180
rect 942 175 943 179
rect 947 175 948 179
rect 942 174 948 175
rect 960 155 962 184
rect 1016 180 1018 210
rect 1238 208 1239 212
rect 1243 208 1244 212
rect 1278 212 1279 216
rect 1283 212 1284 216
rect 1394 215 1395 219
rect 1399 215 1400 219
rect 1394 214 1400 215
rect 1434 219 1440 220
rect 1434 215 1435 219
rect 1439 215 1440 219
rect 1434 214 1440 215
rect 1510 219 1516 220
rect 1510 215 1511 219
rect 1515 215 1516 219
rect 1510 214 1516 215
rect 1642 219 1648 220
rect 1642 215 1643 219
rect 1647 215 1648 219
rect 1642 214 1648 215
rect 1278 211 1284 212
rect 1374 211 1380 212
rect 1238 207 1244 208
rect 1022 189 1028 190
rect 1022 185 1023 189
rect 1027 185 1028 189
rect 1022 184 1028 185
rect 1014 179 1020 180
rect 1014 175 1015 179
rect 1019 175 1020 179
rect 1014 174 1020 175
rect 1024 155 1026 184
rect 1240 155 1242 207
rect 1280 163 1282 211
rect 1374 207 1375 211
rect 1379 207 1380 211
rect 1374 206 1380 207
rect 1366 193 1372 194
rect 1366 189 1367 193
rect 1371 189 1372 193
rect 1366 188 1372 189
rect 1368 163 1370 188
rect 1376 184 1378 206
rect 1396 184 1398 214
rect 1406 193 1412 194
rect 1406 189 1407 193
rect 1411 189 1412 193
rect 1406 188 1412 189
rect 1374 183 1380 184
rect 1374 179 1375 183
rect 1379 179 1380 183
rect 1374 178 1380 179
rect 1394 183 1400 184
rect 1394 179 1395 183
rect 1399 179 1400 183
rect 1394 178 1400 179
rect 1408 163 1410 188
rect 1436 184 1438 214
rect 1446 193 1452 194
rect 1446 189 1447 193
rect 1451 189 1452 193
rect 1446 188 1452 189
rect 1494 193 1500 194
rect 1494 189 1495 193
rect 1499 189 1500 193
rect 1494 188 1500 189
rect 1434 183 1440 184
rect 1434 179 1435 183
rect 1439 179 1440 183
rect 1434 178 1440 179
rect 1448 163 1450 188
rect 1496 163 1498 188
rect 1279 162 1283 163
rect 1279 157 1283 158
rect 1303 162 1307 163
rect 1303 157 1307 158
rect 1343 162 1347 163
rect 1343 157 1347 158
rect 1367 162 1371 163
rect 1367 157 1371 158
rect 1383 162 1387 163
rect 1383 157 1387 158
rect 1407 162 1411 163
rect 1407 157 1411 158
rect 1423 162 1427 163
rect 1423 157 1427 158
rect 1447 162 1451 163
rect 1447 157 1451 158
rect 1463 162 1467 163
rect 1463 157 1467 158
rect 1495 162 1499 163
rect 1495 157 1499 158
rect 767 154 771 155
rect 767 149 771 150
rect 791 154 795 155
rect 791 149 795 150
rect 807 154 811 155
rect 807 149 811 150
rect 847 154 851 155
rect 847 149 851 150
rect 887 154 891 155
rect 887 149 891 150
rect 903 154 907 155
rect 903 149 907 150
rect 927 154 931 155
rect 927 149 931 150
rect 959 154 963 155
rect 959 149 963 150
rect 975 154 979 155
rect 975 149 979 150
rect 1023 154 1027 155
rect 1023 149 1027 150
rect 1071 154 1075 155
rect 1071 149 1075 150
rect 1111 154 1115 155
rect 1111 149 1115 150
rect 1151 154 1155 155
rect 1151 149 1155 150
rect 1191 154 1195 155
rect 1191 149 1195 150
rect 1239 154 1243 155
rect 1239 149 1243 150
rect 768 140 770 149
rect 782 147 788 148
rect 782 143 783 147
rect 787 143 788 147
rect 782 142 788 143
rect 766 139 772 140
rect 766 135 767 139
rect 771 135 772 139
rect 766 134 772 135
rect 784 120 786 142
rect 808 140 810 149
rect 834 147 840 148
rect 834 143 835 147
rect 839 143 840 147
rect 834 142 840 143
rect 806 139 812 140
rect 806 135 807 139
rect 811 135 812 139
rect 806 134 812 135
rect 836 120 838 142
rect 848 140 850 149
rect 874 147 880 148
rect 874 143 875 147
rect 879 143 880 147
rect 874 142 880 143
rect 846 139 852 140
rect 846 135 847 139
rect 851 135 852 139
rect 846 134 852 135
rect 876 120 878 142
rect 888 140 890 149
rect 914 147 920 148
rect 914 143 915 147
rect 919 143 920 147
rect 914 142 920 143
rect 886 139 892 140
rect 886 135 887 139
rect 891 135 892 139
rect 886 134 892 135
rect 916 120 918 142
rect 928 140 930 149
rect 976 140 978 149
rect 1010 147 1016 148
rect 1010 143 1011 147
rect 1015 143 1016 147
rect 1010 142 1016 143
rect 926 139 932 140
rect 926 135 927 139
rect 931 135 932 139
rect 926 134 932 135
rect 974 139 980 140
rect 974 135 975 139
rect 979 135 980 139
rect 974 134 980 135
rect 782 119 788 120
rect 782 115 783 119
rect 787 115 788 119
rect 782 114 788 115
rect 834 119 840 120
rect 834 115 835 119
rect 839 115 840 119
rect 834 114 840 115
rect 874 119 880 120
rect 874 115 875 119
rect 879 115 880 119
rect 874 114 880 115
rect 914 119 920 120
rect 914 115 915 119
rect 919 115 920 119
rect 914 114 920 115
rect 1012 112 1014 142
rect 1024 140 1026 149
rect 1058 147 1064 148
rect 1058 143 1059 147
rect 1063 143 1064 147
rect 1058 142 1064 143
rect 1022 139 1028 140
rect 1022 135 1023 139
rect 1027 135 1028 139
rect 1022 134 1028 135
rect 1060 112 1062 142
rect 1072 140 1074 149
rect 1098 147 1104 148
rect 1098 143 1099 147
rect 1103 143 1104 147
rect 1098 142 1104 143
rect 1070 139 1076 140
rect 1070 135 1071 139
rect 1075 135 1076 139
rect 1070 134 1076 135
rect 1100 120 1102 142
rect 1112 140 1114 149
rect 1134 147 1140 148
rect 1134 143 1135 147
rect 1139 143 1140 147
rect 1134 142 1140 143
rect 1110 139 1116 140
rect 1110 135 1111 139
rect 1115 135 1116 139
rect 1110 134 1116 135
rect 1136 120 1138 142
rect 1152 140 1154 149
rect 1178 147 1184 148
rect 1178 143 1179 147
rect 1183 143 1184 147
rect 1178 142 1184 143
rect 1150 139 1156 140
rect 1150 135 1151 139
rect 1155 135 1156 139
rect 1150 134 1156 135
rect 1180 120 1182 142
rect 1192 140 1194 149
rect 1190 139 1196 140
rect 1190 135 1191 139
rect 1195 135 1196 139
rect 1190 134 1196 135
rect 1098 119 1104 120
rect 1098 115 1099 119
rect 1103 115 1104 119
rect 1098 114 1104 115
rect 1134 119 1140 120
rect 1134 115 1135 119
rect 1139 115 1140 119
rect 1134 114 1140 115
rect 1178 119 1184 120
rect 1178 115 1179 119
rect 1183 115 1184 119
rect 1240 117 1242 149
rect 1280 125 1282 157
rect 1304 148 1306 157
rect 1330 155 1336 156
rect 1330 151 1331 155
rect 1335 151 1336 155
rect 1330 150 1336 151
rect 1294 147 1300 148
rect 1294 143 1295 147
rect 1299 143 1300 147
rect 1294 142 1300 143
rect 1302 147 1308 148
rect 1302 143 1303 147
rect 1307 143 1308 147
rect 1302 142 1308 143
rect 1278 124 1284 125
rect 1278 120 1279 124
rect 1283 120 1284 124
rect 1296 120 1298 142
rect 1278 119 1284 120
rect 1294 119 1300 120
rect 1178 114 1184 115
rect 1238 116 1244 117
rect 1238 112 1239 116
rect 1243 112 1244 116
rect 1294 115 1295 119
rect 1299 115 1300 119
rect 1332 118 1334 150
rect 1344 148 1346 157
rect 1358 155 1364 156
rect 1358 151 1359 155
rect 1363 151 1364 155
rect 1358 150 1364 151
rect 1342 147 1348 148
rect 1342 143 1343 147
rect 1347 143 1348 147
rect 1342 142 1348 143
rect 1360 128 1362 150
rect 1384 148 1386 157
rect 1398 155 1404 156
rect 1398 151 1399 155
rect 1403 151 1404 155
rect 1398 150 1404 151
rect 1382 147 1388 148
rect 1382 143 1383 147
rect 1387 143 1388 147
rect 1382 142 1388 143
rect 1400 128 1402 150
rect 1424 148 1426 157
rect 1438 155 1444 156
rect 1438 151 1439 155
rect 1443 151 1444 155
rect 1438 150 1444 151
rect 1422 147 1428 148
rect 1422 143 1423 147
rect 1427 143 1428 147
rect 1422 142 1428 143
rect 1440 128 1442 150
rect 1464 148 1466 157
rect 1512 156 1514 214
rect 1550 193 1556 194
rect 1550 189 1551 193
rect 1555 189 1556 193
rect 1550 188 1556 189
rect 1606 193 1612 194
rect 1606 189 1607 193
rect 1611 189 1612 193
rect 1606 188 1612 189
rect 1552 163 1554 188
rect 1608 163 1610 188
rect 1644 184 1646 214
rect 1670 193 1676 194
rect 1670 189 1671 193
rect 1675 189 1676 193
rect 1670 188 1676 189
rect 1642 183 1648 184
rect 1642 179 1643 183
rect 1647 179 1648 183
rect 1642 178 1648 179
rect 1672 163 1674 188
rect 1712 184 1714 262
rect 1742 256 1748 257
rect 1742 252 1743 256
rect 1747 252 1748 256
rect 1742 251 1748 252
rect 1798 256 1804 257
rect 1798 252 1799 256
rect 1803 252 1804 256
rect 1798 251 1804 252
rect 1862 256 1868 257
rect 1862 252 1863 256
rect 1867 252 1868 256
rect 1862 251 1868 252
rect 1934 256 1940 257
rect 1934 252 1935 256
rect 1939 252 1940 256
rect 1934 251 1940 252
rect 1744 247 1746 251
rect 1800 247 1802 251
rect 1864 247 1866 251
rect 1936 247 1938 251
rect 1735 246 1739 247
rect 1735 241 1739 242
rect 1743 246 1747 247
rect 1743 241 1747 242
rect 1799 246 1803 247
rect 1799 241 1803 242
rect 1807 246 1811 247
rect 1807 241 1811 242
rect 1863 246 1867 247
rect 1863 241 1867 242
rect 1887 246 1891 247
rect 1887 241 1891 242
rect 1935 246 1939 247
rect 1935 241 1939 242
rect 1975 246 1979 247
rect 1975 241 1979 242
rect 1734 240 1740 241
rect 1734 236 1735 240
rect 1739 236 1740 240
rect 1734 235 1740 236
rect 1806 240 1812 241
rect 1806 236 1807 240
rect 1811 236 1812 240
rect 1806 235 1812 236
rect 1886 240 1892 241
rect 1886 236 1887 240
rect 1891 236 1892 240
rect 1886 235 1892 236
rect 1974 240 1980 241
rect 1974 236 1975 240
rect 1979 236 1980 240
rect 1974 235 1980 236
rect 1798 219 1804 220
rect 1798 215 1799 219
rect 1803 215 1804 219
rect 1798 214 1804 215
rect 1878 219 1884 220
rect 1878 215 1879 219
rect 1883 215 1884 219
rect 1878 214 1884 215
rect 1966 219 1972 220
rect 1966 215 1967 219
rect 1971 215 1972 219
rect 1966 214 1972 215
rect 1734 193 1740 194
rect 1734 189 1735 193
rect 1739 189 1740 193
rect 1734 188 1740 189
rect 1743 188 1747 189
rect 1710 183 1716 184
rect 1710 179 1711 183
rect 1715 179 1716 183
rect 1710 178 1716 179
rect 1736 163 1738 188
rect 1800 184 1802 214
rect 1806 193 1812 194
rect 1806 189 1807 193
rect 1811 189 1812 193
rect 1806 188 1812 189
rect 1742 183 1748 184
rect 1742 179 1743 183
rect 1747 179 1748 183
rect 1742 178 1748 179
rect 1798 183 1804 184
rect 1798 179 1799 183
rect 1803 179 1804 183
rect 1798 178 1804 179
rect 1808 163 1810 188
rect 1880 184 1882 214
rect 1886 193 1892 194
rect 1886 189 1887 193
rect 1891 189 1892 193
rect 1886 188 1892 189
rect 1878 183 1884 184
rect 1878 179 1879 183
rect 1883 179 1884 183
rect 1878 178 1884 179
rect 1888 163 1890 188
rect 1968 184 1970 214
rect 1974 193 1980 194
rect 1974 189 1975 193
rect 1979 189 1980 193
rect 1984 189 1986 270
rect 2006 256 2012 257
rect 2006 252 2007 256
rect 2011 252 2012 256
rect 2006 251 2012 252
rect 2070 256 2076 257
rect 2070 252 2071 256
rect 2075 252 2076 256
rect 2070 251 2076 252
rect 2008 247 2010 251
rect 2072 247 2074 251
rect 2007 246 2011 247
rect 2007 241 2011 242
rect 2071 246 2075 247
rect 2071 241 2075 242
rect 2070 240 2076 241
rect 2070 236 2071 240
rect 2075 236 2076 240
rect 2070 235 2076 236
rect 2092 220 2094 306
rect 2100 276 2102 306
rect 2136 304 2138 313
rect 2162 311 2168 312
rect 2162 307 2163 311
rect 2167 307 2168 311
rect 2162 306 2168 307
rect 2134 303 2140 304
rect 2134 299 2135 303
rect 2139 299 2140 303
rect 2134 298 2140 299
rect 2164 276 2166 306
rect 2192 304 2194 313
rect 2218 311 2224 312
rect 2218 307 2219 311
rect 2223 307 2224 311
rect 2218 306 2224 307
rect 2190 303 2196 304
rect 2190 299 2191 303
rect 2195 299 2196 303
rect 2190 298 2196 299
rect 2220 276 2222 306
rect 2256 304 2258 313
rect 2254 303 2260 304
rect 2254 299 2255 303
rect 2259 299 2260 303
rect 2254 298 2260 299
rect 2284 276 2286 322
rect 2304 319 2306 332
rect 2303 318 2307 319
rect 2303 313 2307 314
rect 2319 318 2323 319
rect 2319 313 2323 314
rect 2320 304 2322 313
rect 2340 312 2342 358
rect 2352 328 2354 414
rect 2406 407 2412 408
rect 2406 403 2407 407
rect 2411 403 2412 407
rect 2406 402 2412 403
rect 2358 400 2364 401
rect 2358 396 2359 400
rect 2363 396 2364 400
rect 2358 395 2364 396
rect 2360 391 2362 395
rect 2408 391 2410 402
rect 2359 390 2363 391
rect 2359 385 2363 386
rect 2407 390 2411 391
rect 2407 385 2411 386
rect 2358 384 2364 385
rect 2358 380 2359 384
rect 2363 380 2364 384
rect 2358 379 2364 380
rect 2408 378 2410 385
rect 2406 377 2412 378
rect 2406 373 2407 377
rect 2411 373 2412 377
rect 2406 372 2412 373
rect 2406 360 2412 361
rect 2406 356 2407 360
rect 2411 356 2412 360
rect 2406 355 2412 356
rect 2358 337 2364 338
rect 2358 333 2359 337
rect 2363 333 2364 337
rect 2358 332 2364 333
rect 2350 327 2356 328
rect 2350 323 2351 327
rect 2355 323 2356 327
rect 2350 322 2356 323
rect 2360 319 2362 332
rect 2408 319 2410 355
rect 2359 318 2363 319
rect 2359 313 2363 314
rect 2407 318 2411 319
rect 2407 313 2411 314
rect 2338 311 2344 312
rect 2338 307 2339 311
rect 2343 307 2344 311
rect 2338 306 2344 307
rect 2346 311 2352 312
rect 2346 307 2347 311
rect 2351 307 2352 311
rect 2346 306 2352 307
rect 2318 303 2324 304
rect 2318 299 2319 303
rect 2323 299 2324 303
rect 2318 298 2324 299
rect 2348 276 2350 306
rect 2360 304 2362 313
rect 2358 303 2364 304
rect 2358 299 2359 303
rect 2363 299 2364 303
rect 2358 298 2364 299
rect 2408 281 2410 313
rect 2406 280 2412 281
rect 2406 276 2407 280
rect 2411 276 2412 280
rect 2098 275 2104 276
rect 2098 271 2099 275
rect 2103 271 2104 275
rect 2098 270 2104 271
rect 2162 275 2168 276
rect 2162 271 2163 275
rect 2167 271 2168 275
rect 2162 270 2168 271
rect 2218 275 2224 276
rect 2218 271 2219 275
rect 2223 271 2224 275
rect 2218 270 2224 271
rect 2282 275 2288 276
rect 2282 271 2283 275
rect 2287 271 2288 275
rect 2282 270 2288 271
rect 2346 275 2352 276
rect 2346 271 2347 275
rect 2351 271 2352 275
rect 2346 270 2352 271
rect 2374 275 2380 276
rect 2406 275 2412 276
rect 2374 271 2375 275
rect 2379 271 2380 275
rect 2374 270 2380 271
rect 2134 256 2140 257
rect 2134 252 2135 256
rect 2139 252 2140 256
rect 2134 251 2140 252
rect 2190 256 2196 257
rect 2190 252 2191 256
rect 2195 252 2196 256
rect 2190 251 2196 252
rect 2254 256 2260 257
rect 2254 252 2255 256
rect 2259 252 2260 256
rect 2254 251 2260 252
rect 2318 256 2324 257
rect 2318 252 2319 256
rect 2323 252 2324 256
rect 2318 251 2324 252
rect 2358 256 2364 257
rect 2358 252 2359 256
rect 2363 252 2364 256
rect 2358 251 2364 252
rect 2136 247 2138 251
rect 2192 247 2194 251
rect 2256 247 2258 251
rect 2320 247 2322 251
rect 2360 247 2362 251
rect 2135 246 2139 247
rect 2135 241 2139 242
rect 2167 246 2171 247
rect 2167 241 2171 242
rect 2191 246 2195 247
rect 2191 241 2195 242
rect 2255 246 2259 247
rect 2255 241 2259 242
rect 2271 246 2275 247
rect 2271 241 2275 242
rect 2319 246 2323 247
rect 2319 241 2323 242
rect 2359 246 2363 247
rect 2359 241 2363 242
rect 2166 240 2172 241
rect 2166 236 2167 240
rect 2171 236 2172 240
rect 2166 235 2172 236
rect 2270 240 2276 241
rect 2270 236 2271 240
rect 2275 236 2276 240
rect 2270 235 2276 236
rect 2358 240 2364 241
rect 2358 236 2359 240
rect 2363 236 2364 240
rect 2358 235 2364 236
rect 1990 219 1996 220
rect 1990 215 1991 219
rect 1995 215 1996 219
rect 1990 214 1996 215
rect 2090 219 2096 220
rect 2090 215 2091 219
rect 2095 215 2096 219
rect 2090 214 2096 215
rect 2366 219 2372 220
rect 2366 215 2367 219
rect 2371 215 2372 219
rect 2366 214 2372 215
rect 1974 188 1980 189
rect 1983 188 1987 189
rect 1966 183 1972 184
rect 1966 179 1967 183
rect 1971 179 1972 183
rect 1966 178 1972 179
rect 1976 163 1978 188
rect 1983 183 1987 184
rect 1992 164 1994 214
rect 2070 193 2076 194
rect 2070 189 2071 193
rect 2075 189 2076 193
rect 2070 188 2076 189
rect 2166 193 2172 194
rect 2166 189 2167 193
rect 2171 189 2172 193
rect 2166 188 2172 189
rect 2270 193 2276 194
rect 2270 189 2271 193
rect 2275 189 2276 193
rect 2270 188 2276 189
rect 2358 193 2364 194
rect 2358 189 2359 193
rect 2363 189 2364 193
rect 2358 188 2364 189
rect 1990 163 1996 164
rect 2072 163 2074 188
rect 2168 163 2170 188
rect 2242 183 2248 184
rect 2242 179 2243 183
rect 2247 179 2248 183
rect 2242 178 2248 179
rect 1519 162 1523 163
rect 1519 157 1523 158
rect 1551 162 1555 163
rect 1551 157 1555 158
rect 1583 162 1587 163
rect 1583 157 1587 158
rect 1607 162 1611 163
rect 1607 157 1611 158
rect 1647 162 1651 163
rect 1647 157 1651 158
rect 1671 162 1675 163
rect 1671 157 1675 158
rect 1711 162 1715 163
rect 1711 157 1715 158
rect 1735 162 1739 163
rect 1735 157 1739 158
rect 1767 162 1771 163
rect 1767 157 1771 158
rect 1807 162 1811 163
rect 1807 157 1811 158
rect 1823 162 1827 163
rect 1823 157 1827 158
rect 1871 162 1875 163
rect 1871 157 1875 158
rect 1887 162 1891 163
rect 1887 157 1891 158
rect 1919 162 1923 163
rect 1919 157 1923 158
rect 1967 162 1971 163
rect 1967 157 1971 158
rect 1975 162 1979 163
rect 1990 159 1991 163
rect 1995 159 1996 163
rect 1990 158 1996 159
rect 2015 162 2019 163
rect 1975 157 1979 158
rect 2015 157 2019 158
rect 2063 162 2067 163
rect 2063 157 2067 158
rect 2071 162 2075 163
rect 2071 157 2075 158
rect 2111 162 2115 163
rect 2111 157 2115 158
rect 2159 162 2163 163
rect 2159 157 2163 158
rect 2167 162 2171 163
rect 2167 157 2171 158
rect 2215 162 2219 163
rect 2215 157 2219 158
rect 1502 155 1508 156
rect 1502 151 1503 155
rect 1507 151 1508 155
rect 1502 150 1508 151
rect 1510 155 1516 156
rect 1510 151 1511 155
rect 1515 151 1516 155
rect 1510 150 1516 151
rect 1462 147 1468 148
rect 1462 143 1463 147
rect 1467 143 1468 147
rect 1462 142 1468 143
rect 1504 132 1506 150
rect 1520 148 1522 157
rect 1584 148 1586 157
rect 1648 148 1650 157
rect 1712 148 1714 157
rect 1768 148 1770 157
rect 1824 148 1826 157
rect 1850 155 1856 156
rect 1850 151 1851 155
rect 1855 151 1856 155
rect 1850 150 1856 151
rect 1518 147 1524 148
rect 1518 143 1519 147
rect 1523 143 1524 147
rect 1518 142 1524 143
rect 1582 147 1588 148
rect 1582 143 1583 147
rect 1587 143 1588 147
rect 1582 142 1588 143
rect 1646 147 1652 148
rect 1646 143 1647 147
rect 1651 143 1652 147
rect 1646 142 1652 143
rect 1710 147 1716 148
rect 1710 143 1711 147
rect 1715 143 1716 147
rect 1710 142 1716 143
rect 1766 147 1772 148
rect 1766 143 1767 147
rect 1771 143 1772 147
rect 1766 142 1772 143
rect 1822 147 1828 148
rect 1822 143 1823 147
rect 1827 143 1828 147
rect 1822 142 1828 143
rect 1502 131 1508 132
rect 1358 127 1364 128
rect 1358 123 1359 127
rect 1363 123 1364 127
rect 1358 122 1364 123
rect 1398 127 1404 128
rect 1398 123 1399 127
rect 1403 123 1404 127
rect 1398 122 1404 123
rect 1438 127 1444 128
rect 1438 123 1439 127
rect 1443 123 1444 127
rect 1502 127 1503 131
rect 1507 127 1508 131
rect 1502 126 1508 127
rect 1438 122 1444 123
rect 1852 120 1854 150
rect 1872 148 1874 157
rect 1898 155 1904 156
rect 1898 151 1899 155
rect 1903 151 1904 155
rect 1898 150 1904 151
rect 1870 147 1876 148
rect 1870 143 1871 147
rect 1875 143 1876 147
rect 1870 142 1876 143
rect 1900 120 1902 150
rect 1920 148 1922 157
rect 1946 155 1952 156
rect 1946 151 1947 155
rect 1951 151 1952 155
rect 1946 150 1952 151
rect 1918 147 1924 148
rect 1918 143 1919 147
rect 1923 143 1924 147
rect 1918 142 1924 143
rect 1948 120 1950 150
rect 1968 148 1970 157
rect 1994 155 2000 156
rect 1994 151 1995 155
rect 1999 151 2000 155
rect 1994 150 2000 151
rect 1966 147 1972 148
rect 1966 143 1967 147
rect 1971 143 1972 147
rect 1966 142 1972 143
rect 1996 120 1998 150
rect 2016 148 2018 157
rect 2042 155 2048 156
rect 2042 151 2043 155
rect 2047 151 2048 155
rect 2042 150 2048 151
rect 2014 147 2020 148
rect 2014 143 2015 147
rect 2019 143 2020 147
rect 2014 142 2020 143
rect 2044 120 2046 150
rect 2064 148 2066 157
rect 2090 155 2096 156
rect 2090 151 2091 155
rect 2095 151 2096 155
rect 2090 150 2096 151
rect 2062 147 2068 148
rect 2062 143 2063 147
rect 2067 143 2068 147
rect 2062 142 2068 143
rect 2092 120 2094 150
rect 2112 148 2114 157
rect 2138 155 2144 156
rect 2138 151 2139 155
rect 2143 151 2144 155
rect 2138 150 2144 151
rect 2110 147 2116 148
rect 2110 143 2111 147
rect 2115 143 2116 147
rect 2110 142 2116 143
rect 2140 120 2142 150
rect 2160 148 2162 157
rect 2186 155 2192 156
rect 2186 151 2187 155
rect 2191 151 2192 155
rect 2186 150 2192 151
rect 2158 147 2164 148
rect 2158 143 2159 147
rect 2163 143 2164 147
rect 2158 142 2164 143
rect 2188 120 2190 150
rect 2216 148 2218 157
rect 2214 147 2220 148
rect 2214 143 2215 147
rect 2219 143 2220 147
rect 2214 142 2220 143
rect 2244 120 2246 178
rect 2272 163 2274 188
rect 2360 163 2362 188
rect 2271 162 2275 163
rect 2271 157 2275 158
rect 2319 162 2323 163
rect 2319 157 2323 158
rect 2359 162 2363 163
rect 2359 157 2363 158
rect 2272 148 2274 157
rect 2306 155 2312 156
rect 2306 151 2307 155
rect 2311 151 2312 155
rect 2306 150 2312 151
rect 2270 147 2276 148
rect 2270 143 2271 147
rect 2275 143 2276 147
rect 2270 142 2276 143
rect 2308 120 2310 150
rect 2320 148 2322 157
rect 2346 155 2352 156
rect 2346 151 2347 155
rect 2351 151 2352 155
rect 2346 150 2352 151
rect 2318 147 2324 148
rect 2318 143 2319 147
rect 2323 143 2324 147
rect 2318 142 2324 143
rect 2348 128 2350 150
rect 2360 148 2362 157
rect 2368 156 2370 214
rect 2376 184 2378 270
rect 2406 263 2412 264
rect 2406 259 2407 263
rect 2411 259 2412 263
rect 2406 258 2412 259
rect 2408 247 2410 258
rect 2407 246 2411 247
rect 2407 241 2411 242
rect 2408 234 2410 241
rect 2406 233 2412 234
rect 2406 229 2407 233
rect 2411 229 2412 233
rect 2406 228 2412 229
rect 2406 216 2412 217
rect 2406 212 2407 216
rect 2411 212 2412 216
rect 2406 211 2412 212
rect 2374 183 2380 184
rect 2374 179 2375 183
rect 2379 179 2380 183
rect 2374 178 2380 179
rect 2408 163 2410 211
rect 2407 162 2411 163
rect 2407 157 2411 158
rect 2366 155 2372 156
rect 2366 151 2367 155
rect 2371 151 2372 155
rect 2366 150 2372 151
rect 2358 147 2364 148
rect 2358 143 2359 147
rect 2363 143 2364 147
rect 2358 142 2364 143
rect 2346 127 2352 128
rect 2346 123 2347 127
rect 2351 123 2352 127
rect 2408 125 2410 157
rect 2346 122 2352 123
rect 2406 124 2412 125
rect 2406 120 2407 124
rect 2411 120 2412 124
rect 1338 119 1344 120
rect 1338 118 1339 119
rect 1332 116 1339 118
rect 1294 114 1300 115
rect 1338 115 1339 116
rect 1343 115 1344 119
rect 1338 114 1344 115
rect 1850 119 1856 120
rect 1850 115 1851 119
rect 1855 115 1856 119
rect 1850 114 1856 115
rect 1898 119 1904 120
rect 1898 115 1899 119
rect 1903 115 1904 119
rect 1898 114 1904 115
rect 1946 119 1952 120
rect 1946 115 1947 119
rect 1951 115 1952 119
rect 1946 114 1952 115
rect 1994 119 2000 120
rect 1994 115 1995 119
rect 1999 115 2000 119
rect 1994 114 2000 115
rect 2042 119 2048 120
rect 2042 115 2043 119
rect 2047 115 2048 119
rect 2042 114 2048 115
rect 2090 119 2096 120
rect 2090 115 2091 119
rect 2095 115 2096 119
rect 2090 114 2096 115
rect 2138 119 2144 120
rect 2138 115 2139 119
rect 2143 115 2144 119
rect 2138 114 2144 115
rect 2186 119 2192 120
rect 2186 115 2187 119
rect 2191 115 2192 119
rect 2186 114 2192 115
rect 2242 119 2248 120
rect 2242 115 2243 119
rect 2247 115 2248 119
rect 2242 114 2248 115
rect 2306 119 2312 120
rect 2406 119 2412 120
rect 2306 115 2307 119
rect 2311 115 2312 119
rect 2306 114 2312 115
rect 110 111 116 112
rect 158 111 164 112
rect 158 107 159 111
rect 163 107 164 111
rect 158 106 164 107
rect 202 111 208 112
rect 202 107 203 111
rect 207 107 208 111
rect 202 106 208 107
rect 238 111 244 112
rect 238 107 239 111
rect 243 107 244 111
rect 238 106 244 107
rect 458 111 464 112
rect 458 107 459 111
rect 463 107 464 111
rect 458 106 464 107
rect 554 111 560 112
rect 554 107 555 111
rect 559 107 560 111
rect 554 106 560 107
rect 706 111 712 112
rect 706 107 707 111
rect 711 107 712 111
rect 706 106 712 107
rect 750 111 756 112
rect 750 107 751 111
rect 755 107 756 111
rect 750 106 756 107
rect 1010 111 1016 112
rect 1010 107 1011 111
rect 1015 107 1016 111
rect 1010 106 1016 107
rect 1058 111 1064 112
rect 1238 111 1244 112
rect 1058 107 1059 111
rect 1063 107 1064 111
rect 1058 106 1064 107
rect 1278 107 1284 108
rect 1278 103 1279 107
rect 1283 103 1284 107
rect 1278 102 1284 103
rect 2406 107 2412 108
rect 2406 103 2407 107
rect 2411 103 2412 107
rect 2406 102 2412 103
rect 110 99 116 100
rect 110 95 111 99
rect 115 95 116 99
rect 110 94 116 95
rect 1238 99 1244 100
rect 1238 95 1239 99
rect 1243 95 1244 99
rect 1280 95 1282 102
rect 1302 100 1308 101
rect 1302 96 1303 100
rect 1307 96 1308 100
rect 1302 95 1308 96
rect 1342 100 1348 101
rect 1342 96 1343 100
rect 1347 96 1348 100
rect 1342 95 1348 96
rect 1382 100 1388 101
rect 1382 96 1383 100
rect 1387 96 1388 100
rect 1382 95 1388 96
rect 1422 100 1428 101
rect 1422 96 1423 100
rect 1427 96 1428 100
rect 1422 95 1428 96
rect 1462 100 1468 101
rect 1462 96 1463 100
rect 1467 96 1468 100
rect 1462 95 1468 96
rect 1518 100 1524 101
rect 1518 96 1519 100
rect 1523 96 1524 100
rect 1518 95 1524 96
rect 1582 100 1588 101
rect 1582 96 1583 100
rect 1587 96 1588 100
rect 1582 95 1588 96
rect 1646 100 1652 101
rect 1646 96 1647 100
rect 1651 96 1652 100
rect 1646 95 1652 96
rect 1710 100 1716 101
rect 1710 96 1711 100
rect 1715 96 1716 100
rect 1710 95 1716 96
rect 1766 100 1772 101
rect 1766 96 1767 100
rect 1771 96 1772 100
rect 1766 95 1772 96
rect 1822 100 1828 101
rect 1822 96 1823 100
rect 1827 96 1828 100
rect 1822 95 1828 96
rect 1870 100 1876 101
rect 1870 96 1871 100
rect 1875 96 1876 100
rect 1870 95 1876 96
rect 1918 100 1924 101
rect 1918 96 1919 100
rect 1923 96 1924 100
rect 1918 95 1924 96
rect 1966 100 1972 101
rect 1966 96 1967 100
rect 1971 96 1972 100
rect 1966 95 1972 96
rect 2014 100 2020 101
rect 2014 96 2015 100
rect 2019 96 2020 100
rect 2014 95 2020 96
rect 2062 100 2068 101
rect 2062 96 2063 100
rect 2067 96 2068 100
rect 2062 95 2068 96
rect 2110 100 2116 101
rect 2110 96 2111 100
rect 2115 96 2116 100
rect 2110 95 2116 96
rect 2158 100 2164 101
rect 2158 96 2159 100
rect 2163 96 2164 100
rect 2158 95 2164 96
rect 2214 100 2220 101
rect 2214 96 2215 100
rect 2219 96 2220 100
rect 2214 95 2220 96
rect 2270 100 2276 101
rect 2270 96 2271 100
rect 2275 96 2276 100
rect 2270 95 2276 96
rect 2318 100 2324 101
rect 2318 96 2319 100
rect 2323 96 2324 100
rect 2318 95 2324 96
rect 2358 100 2364 101
rect 2358 96 2359 100
rect 2363 96 2364 100
rect 2358 95 2364 96
rect 2408 95 2410 102
rect 1238 94 1244 95
rect 1279 94 1283 95
rect 112 87 114 94
rect 134 92 140 93
rect 134 88 135 92
rect 139 88 140 92
rect 134 87 140 88
rect 174 92 180 93
rect 174 88 175 92
rect 179 88 180 92
rect 174 87 180 88
rect 214 92 220 93
rect 214 88 215 92
rect 219 88 220 92
rect 214 87 220 88
rect 254 92 260 93
rect 254 88 255 92
rect 259 88 260 92
rect 254 87 260 88
rect 294 92 300 93
rect 294 88 295 92
rect 299 88 300 92
rect 294 87 300 88
rect 334 92 340 93
rect 334 88 335 92
rect 339 88 340 92
rect 334 87 340 88
rect 374 92 380 93
rect 374 88 375 92
rect 379 88 380 92
rect 374 87 380 88
rect 422 92 428 93
rect 422 88 423 92
rect 427 88 428 92
rect 422 87 428 88
rect 470 92 476 93
rect 470 88 471 92
rect 475 88 476 92
rect 470 87 476 88
rect 526 92 532 93
rect 526 88 527 92
rect 531 88 532 92
rect 526 87 532 88
rect 582 92 588 93
rect 582 88 583 92
rect 587 88 588 92
rect 582 87 588 88
rect 630 92 636 93
rect 630 88 631 92
rect 635 88 636 92
rect 630 87 636 88
rect 678 92 684 93
rect 678 88 679 92
rect 683 88 684 92
rect 678 87 684 88
rect 726 92 732 93
rect 726 88 727 92
rect 731 88 732 92
rect 726 87 732 88
rect 766 92 772 93
rect 766 88 767 92
rect 771 88 772 92
rect 766 87 772 88
rect 806 92 812 93
rect 806 88 807 92
rect 811 88 812 92
rect 806 87 812 88
rect 846 92 852 93
rect 846 88 847 92
rect 851 88 852 92
rect 846 87 852 88
rect 886 92 892 93
rect 886 88 887 92
rect 891 88 892 92
rect 886 87 892 88
rect 926 92 932 93
rect 926 88 927 92
rect 931 88 932 92
rect 926 87 932 88
rect 974 92 980 93
rect 974 88 975 92
rect 979 88 980 92
rect 974 87 980 88
rect 1022 92 1028 93
rect 1022 88 1023 92
rect 1027 88 1028 92
rect 1022 87 1028 88
rect 1070 92 1076 93
rect 1070 88 1071 92
rect 1075 88 1076 92
rect 1070 87 1076 88
rect 1110 92 1116 93
rect 1110 88 1111 92
rect 1115 88 1116 92
rect 1110 87 1116 88
rect 1150 92 1156 93
rect 1150 88 1151 92
rect 1155 88 1156 92
rect 1150 87 1156 88
rect 1190 92 1196 93
rect 1190 88 1191 92
rect 1195 88 1196 92
rect 1190 87 1196 88
rect 1240 87 1242 94
rect 1279 89 1283 90
rect 1303 94 1307 95
rect 1303 89 1307 90
rect 1343 94 1347 95
rect 1343 89 1347 90
rect 1383 94 1387 95
rect 1383 89 1387 90
rect 1423 94 1427 95
rect 1423 89 1427 90
rect 1463 94 1467 95
rect 1463 89 1467 90
rect 1519 94 1523 95
rect 1519 89 1523 90
rect 1583 94 1587 95
rect 1583 89 1587 90
rect 1647 94 1651 95
rect 1647 89 1651 90
rect 1711 94 1715 95
rect 1711 89 1715 90
rect 1767 94 1771 95
rect 1767 89 1771 90
rect 1823 94 1827 95
rect 1823 89 1827 90
rect 1871 94 1875 95
rect 1871 89 1875 90
rect 1919 94 1923 95
rect 1919 89 1923 90
rect 1967 94 1971 95
rect 1967 89 1971 90
rect 2015 94 2019 95
rect 2015 89 2019 90
rect 2063 94 2067 95
rect 2063 89 2067 90
rect 2111 94 2115 95
rect 2111 89 2115 90
rect 2159 94 2163 95
rect 2159 89 2163 90
rect 2215 94 2219 95
rect 2215 89 2219 90
rect 2271 94 2275 95
rect 2271 89 2275 90
rect 2319 94 2323 95
rect 2319 89 2323 90
rect 2359 94 2363 95
rect 2359 89 2363 90
rect 2407 94 2411 95
rect 2407 89 2411 90
rect 111 86 115 87
rect 111 81 115 82
rect 135 86 139 87
rect 135 81 139 82
rect 175 86 179 87
rect 175 81 179 82
rect 215 86 219 87
rect 215 81 219 82
rect 255 86 259 87
rect 255 81 259 82
rect 295 86 299 87
rect 295 81 299 82
rect 335 86 339 87
rect 335 81 339 82
rect 375 86 379 87
rect 375 81 379 82
rect 423 86 427 87
rect 423 81 427 82
rect 471 86 475 87
rect 471 81 475 82
rect 527 86 531 87
rect 527 81 531 82
rect 583 86 587 87
rect 583 81 587 82
rect 631 86 635 87
rect 631 81 635 82
rect 679 86 683 87
rect 679 81 683 82
rect 727 86 731 87
rect 727 81 731 82
rect 767 86 771 87
rect 767 81 771 82
rect 807 86 811 87
rect 807 81 811 82
rect 847 86 851 87
rect 847 81 851 82
rect 887 86 891 87
rect 887 81 891 82
rect 927 86 931 87
rect 927 81 931 82
rect 975 86 979 87
rect 975 81 979 82
rect 1023 86 1027 87
rect 1023 81 1027 82
rect 1071 86 1075 87
rect 1071 81 1075 82
rect 1111 86 1115 87
rect 1111 81 1115 82
rect 1151 86 1155 87
rect 1151 81 1155 82
rect 1191 86 1195 87
rect 1191 81 1195 82
rect 1239 86 1243 87
rect 1239 81 1243 82
<< m4c >>
rect 1279 2510 1283 2514
rect 1535 2510 1539 2514
rect 1575 2510 1579 2514
rect 1615 2510 1619 2514
rect 1655 2510 1659 2514
rect 1695 2510 1699 2514
rect 1735 2510 1739 2514
rect 1775 2510 1779 2514
rect 1815 2510 1819 2514
rect 1855 2510 1859 2514
rect 1895 2510 1899 2514
rect 1935 2510 1939 2514
rect 1975 2510 1979 2514
rect 2407 2510 2411 2514
rect 111 2498 115 2502
rect 135 2498 139 2502
rect 175 2498 179 2502
rect 215 2498 219 2502
rect 255 2498 259 2502
rect 311 2498 315 2502
rect 391 2498 395 2502
rect 479 2498 483 2502
rect 567 2498 571 2502
rect 655 2498 659 2502
rect 743 2498 747 2502
rect 831 2498 835 2502
rect 927 2498 931 2502
rect 1239 2498 1243 2502
rect 111 2430 115 2434
rect 135 2430 139 2434
rect 175 2430 179 2434
rect 183 2430 187 2434
rect 215 2430 219 2434
rect 247 2430 251 2434
rect 255 2430 259 2434
rect 311 2430 315 2434
rect 319 2430 323 2434
rect 391 2430 395 2434
rect 471 2430 475 2434
rect 479 2430 483 2434
rect 543 2430 547 2434
rect 567 2430 571 2434
rect 615 2430 619 2434
rect 655 2430 659 2434
rect 679 2430 683 2434
rect 735 2430 739 2434
rect 743 2430 747 2434
rect 791 2430 795 2434
rect 831 2430 835 2434
rect 839 2430 843 2434
rect 111 2354 115 2358
rect 135 2354 139 2358
rect 175 2354 179 2358
rect 183 2354 187 2358
rect 215 2354 219 2358
rect 247 2354 251 2358
rect 271 2354 275 2358
rect 319 2354 323 2358
rect 351 2354 355 2358
rect 391 2354 395 2358
rect 431 2354 435 2358
rect 471 2354 475 2358
rect 519 2354 523 2358
rect 543 2354 547 2358
rect 1279 2442 1283 2446
rect 1359 2442 1363 2446
rect 1399 2442 1403 2446
rect 1455 2442 1459 2446
rect 1519 2442 1523 2446
rect 1535 2442 1539 2446
rect 887 2430 891 2434
rect 927 2430 931 2434
rect 935 2430 939 2434
rect 991 2430 995 2434
rect 1047 2430 1051 2434
rect 1239 2430 1243 2434
rect 1279 2374 1283 2378
rect 1359 2374 1363 2378
rect 599 2354 603 2358
rect 615 2354 619 2358
rect 679 2354 683 2358
rect 735 2354 739 2358
rect 751 2354 755 2358
rect 791 2354 795 2358
rect 823 2354 827 2358
rect 839 2354 843 2358
rect 887 2354 891 2358
rect 935 2354 939 2358
rect 959 2354 963 2358
rect 991 2354 995 2358
rect 1031 2354 1035 2358
rect 1047 2354 1051 2358
rect 1239 2354 1243 2358
rect 111 2282 115 2286
rect 135 2282 139 2286
rect 175 2282 179 2286
rect 215 2282 219 2286
rect 231 2282 235 2286
rect 271 2282 275 2286
rect 303 2282 307 2286
rect 351 2282 355 2286
rect 375 2282 379 2286
rect 431 2282 435 2286
rect 455 2282 459 2286
rect 519 2282 523 2286
rect 535 2282 539 2286
rect 599 2282 603 2286
rect 615 2282 619 2286
rect 679 2282 683 2286
rect 687 2282 691 2286
rect 751 2282 755 2286
rect 759 2282 763 2286
rect 1575 2442 1579 2446
rect 1599 2442 1603 2446
rect 1615 2442 1619 2446
rect 1655 2442 1659 2446
rect 1679 2442 1683 2446
rect 1695 2442 1699 2446
rect 1735 2442 1739 2446
rect 1759 2442 1763 2446
rect 1775 2442 1779 2446
rect 1815 2442 1819 2446
rect 1839 2442 1843 2446
rect 1855 2442 1859 2446
rect 1895 2442 1899 2446
rect 1919 2442 1923 2446
rect 1935 2442 1939 2446
rect 1975 2442 1979 2446
rect 1999 2442 2003 2446
rect 2079 2442 2083 2446
rect 2159 2442 2163 2446
rect 2247 2442 2251 2446
rect 2335 2442 2339 2446
rect 2407 2442 2411 2446
rect 1399 2374 1403 2378
rect 1407 2374 1411 2378
rect 1455 2374 1459 2378
rect 1471 2374 1475 2378
rect 1519 2374 1523 2378
rect 1543 2374 1547 2378
rect 1599 2374 1603 2378
rect 1615 2374 1619 2378
rect 1679 2374 1683 2378
rect 1695 2374 1699 2378
rect 1759 2374 1763 2378
rect 1775 2374 1779 2378
rect 1839 2374 1843 2378
rect 1855 2374 1859 2378
rect 1919 2374 1923 2378
rect 1927 2374 1931 2378
rect 1999 2374 2003 2378
rect 2071 2374 2075 2378
rect 2079 2374 2083 2378
rect 2143 2374 2147 2378
rect 2159 2374 2163 2378
rect 2223 2374 2227 2378
rect 2247 2374 2251 2378
rect 2303 2374 2307 2378
rect 2335 2374 2339 2378
rect 823 2282 827 2286
rect 831 2282 835 2286
rect 887 2282 891 2286
rect 911 2282 915 2286
rect 959 2282 963 2286
rect 991 2282 995 2286
rect 111 2214 115 2218
rect 135 2214 139 2218
rect 175 2214 179 2218
rect 231 2214 235 2218
rect 247 2214 251 2218
rect 287 2214 291 2218
rect 303 2214 307 2218
rect 327 2214 331 2218
rect 375 2214 379 2218
rect 431 2214 435 2218
rect 455 2214 459 2218
rect 495 2214 499 2218
rect 535 2214 539 2218
rect 551 2214 555 2218
rect 607 2214 611 2218
rect 615 2214 619 2218
rect 663 2214 667 2218
rect 687 2214 691 2218
rect 719 2214 723 2218
rect 759 2214 763 2218
rect 783 2214 787 2218
rect 831 2214 835 2218
rect 847 2214 851 2218
rect 111 2138 115 2142
rect 247 2138 251 2142
rect 287 2138 291 2142
rect 327 2138 331 2142
rect 375 2138 379 2142
rect 383 2138 387 2142
rect 423 2138 427 2142
rect 431 2138 435 2142
rect 463 2138 467 2142
rect 495 2138 499 2142
rect 503 2138 507 2142
rect 551 2138 555 2142
rect 1279 2302 1283 2306
rect 1359 2302 1363 2306
rect 1407 2302 1411 2306
rect 1471 2302 1475 2306
rect 1503 2302 1507 2306
rect 1543 2302 1547 2306
rect 1583 2302 1587 2306
rect 1031 2282 1035 2286
rect 1239 2282 1243 2286
rect 1615 2302 1619 2306
rect 1623 2302 1627 2306
rect 1663 2302 1667 2306
rect 1695 2302 1699 2306
rect 1703 2302 1707 2306
rect 1759 2302 1763 2306
rect 1279 2226 1283 2230
rect 1303 2226 1307 2230
rect 1343 2226 1347 2230
rect 1383 2226 1387 2230
rect 1431 2226 1435 2230
rect 1495 2226 1499 2230
rect 1503 2226 1507 2230
rect 1543 2226 1547 2230
rect 1567 2226 1571 2230
rect 1583 2226 1587 2230
rect 1623 2226 1627 2230
rect 1639 2226 1643 2230
rect 911 2214 915 2218
rect 991 2214 995 2218
rect 1239 2214 1243 2218
rect 1775 2302 1779 2306
rect 1823 2302 1827 2306
rect 1855 2302 1859 2306
rect 1895 2302 1899 2306
rect 1927 2302 1931 2306
rect 1967 2302 1971 2306
rect 1999 2302 2003 2306
rect 2047 2302 2051 2306
rect 2071 2302 2075 2306
rect 2127 2302 2131 2306
rect 2143 2302 2147 2306
rect 2207 2302 2211 2306
rect 2223 2302 2227 2306
rect 1663 2226 1667 2230
rect 1703 2226 1707 2230
rect 1711 2226 1715 2230
rect 1759 2226 1763 2230
rect 1783 2226 1787 2230
rect 607 2138 611 2142
rect 663 2138 667 2142
rect 719 2138 723 2142
rect 727 2138 731 2142
rect 783 2138 787 2142
rect 791 2138 795 2142
rect 111 2070 115 2074
rect 383 2070 387 2074
rect 423 2070 427 2074
rect 463 2070 467 2074
rect 503 2070 507 2074
rect 543 2070 547 2074
rect 551 2070 555 2074
rect 583 2070 587 2074
rect 607 2070 611 2074
rect 631 2070 635 2074
rect 663 2070 667 2074
rect 687 2070 691 2074
rect 727 2070 731 2074
rect 743 2070 747 2074
rect 1279 2158 1283 2162
rect 1303 2158 1307 2162
rect 847 2138 851 2142
rect 855 2138 859 2142
rect 911 2138 915 2142
rect 967 2138 971 2142
rect 1023 2138 1027 2142
rect 1079 2138 1083 2142
rect 1143 2138 1147 2142
rect 1239 2138 1243 2142
rect 1343 2158 1347 2162
rect 1351 2158 1355 2162
rect 1383 2158 1387 2162
rect 1431 2158 1435 2162
rect 1439 2158 1443 2162
rect 1495 2158 1499 2162
rect 1535 2158 1539 2162
rect 1567 2158 1571 2162
rect 791 2070 795 2074
rect 799 2070 803 2074
rect 847 2070 851 2074
rect 855 2070 859 2074
rect 111 1994 115 1998
rect 367 1994 371 1998
rect 383 1994 387 1998
rect 407 1994 411 1998
rect 423 1994 427 1998
rect 455 1994 459 1998
rect 463 1994 467 1998
rect 503 1994 507 1998
rect 511 1994 515 1998
rect 543 1994 547 1998
rect 567 1994 571 1998
rect 583 1994 587 1998
rect 631 1994 635 1998
rect 687 1994 691 1998
rect 695 1994 699 1998
rect 743 1994 747 1998
rect 759 1994 763 1998
rect 903 2070 907 2074
rect 911 2070 915 2074
rect 959 2070 963 2074
rect 967 2070 971 2074
rect 1015 2070 1019 2074
rect 1023 2070 1027 2074
rect 1071 2070 1075 2074
rect 1079 2070 1083 2074
rect 1143 2070 1147 2074
rect 1279 2086 1283 2090
rect 1303 2086 1307 2090
rect 1239 2070 1243 2074
rect 1823 2226 1827 2230
rect 1855 2226 1859 2230
rect 1895 2226 1899 2230
rect 1935 2226 1939 2230
rect 1967 2226 1971 2230
rect 2015 2226 2019 2230
rect 2047 2226 2051 2230
rect 2095 2226 2099 2230
rect 2127 2226 2131 2230
rect 2295 2302 2299 2306
rect 2303 2302 2307 2306
rect 2359 2374 2363 2378
rect 2407 2374 2411 2378
rect 2359 2302 2363 2306
rect 2407 2302 2411 2306
rect 2183 2226 2187 2230
rect 2207 2226 2211 2230
rect 2279 2226 2283 2230
rect 2295 2226 2299 2230
rect 2359 2226 2363 2230
rect 1631 2158 1635 2162
rect 1639 2158 1643 2162
rect 1711 2158 1715 2162
rect 1727 2158 1731 2162
rect 1783 2158 1787 2162
rect 1815 2158 1819 2162
rect 1343 2086 1347 2090
rect 1351 2086 1355 2090
rect 1399 2086 1403 2090
rect 799 1994 803 1998
rect 815 1994 819 1998
rect 847 1994 851 1998
rect 871 1994 875 1998
rect 111 1922 115 1926
rect 175 1922 179 1926
rect 215 1922 219 1926
rect 263 1922 267 1926
rect 319 1922 323 1926
rect 367 1922 371 1926
rect 391 1922 395 1926
rect 407 1922 411 1926
rect 455 1922 459 1926
rect 471 1922 475 1926
rect 511 1922 515 1926
rect 551 1922 555 1926
rect 567 1922 571 1926
rect 631 1922 635 1926
rect 639 1922 643 1926
rect 695 1922 699 1926
rect 719 1922 723 1926
rect 759 1922 763 1926
rect 799 1922 803 1926
rect 815 1922 819 1926
rect 111 1846 115 1850
rect 135 1846 139 1850
rect 175 1846 179 1850
rect 215 1846 219 1850
rect 263 1846 267 1850
rect 271 1846 275 1850
rect 319 1846 323 1850
rect 111 1778 115 1782
rect 135 1778 139 1782
rect 351 1846 355 1850
rect 391 1846 395 1850
rect 439 1846 443 1850
rect 471 1846 475 1850
rect 535 1846 539 1850
rect 551 1846 555 1850
rect 631 1846 635 1850
rect 639 1846 643 1850
rect 1279 2010 1283 2014
rect 1303 2010 1307 2014
rect 1343 2010 1347 2014
rect 1351 2010 1355 2014
rect 903 1994 907 1998
rect 935 1994 939 1998
rect 959 1994 963 1998
rect 999 1994 1003 1998
rect 1015 1994 1019 1998
rect 1063 1994 1067 1998
rect 1071 1994 1075 1998
rect 1239 1994 1243 1998
rect 1279 1942 1283 1946
rect 1303 1942 1307 1946
rect 871 1922 875 1926
rect 879 1922 883 1926
rect 935 1922 939 1926
rect 959 1922 963 1926
rect 999 1922 1003 1926
rect 1039 1922 1043 1926
rect 1063 1922 1067 1926
rect 1119 1922 1123 1926
rect 1239 1922 1243 1926
rect 1439 2086 1443 2090
rect 1479 2086 1483 2090
rect 1535 2086 1539 2090
rect 1567 2086 1571 2090
rect 1631 2086 1635 2090
rect 1663 2086 1667 2090
rect 1727 2086 1731 2090
rect 1759 2086 1763 2090
rect 1855 2158 1859 2162
rect 1895 2158 1899 2162
rect 1935 2158 1939 2162
rect 1975 2158 1979 2162
rect 2015 2158 2019 2162
rect 2047 2158 2051 2162
rect 2095 2158 2099 2162
rect 2111 2158 2115 2162
rect 2175 2158 2179 2162
rect 2183 2158 2187 2162
rect 2239 2158 2243 2162
rect 1815 2086 1819 2090
rect 1847 2086 1851 2090
rect 1895 2086 1899 2090
rect 1935 2086 1939 2090
rect 1399 2010 1403 2014
rect 1423 2010 1427 2014
rect 1479 2010 1483 2014
rect 1495 2010 1499 2014
rect 1567 2010 1571 2014
rect 1575 2010 1579 2014
rect 1663 2010 1667 2014
rect 1751 2010 1755 2014
rect 1759 2010 1763 2014
rect 1839 2010 1843 2014
rect 1847 2010 1851 2014
rect 1351 1942 1355 1946
rect 1359 1942 1363 1946
rect 1423 1942 1427 1946
rect 1447 1942 1451 1946
rect 1495 1942 1499 1946
rect 1535 1942 1539 1946
rect 1575 1942 1579 1946
rect 1623 1942 1627 1946
rect 1663 1942 1667 1946
rect 1711 1942 1715 1946
rect 1975 2086 1979 2090
rect 2015 2086 2019 2090
rect 2047 2086 2051 2090
rect 2279 2158 2283 2162
rect 2311 2158 2315 2162
rect 2407 2226 2411 2230
rect 2359 2158 2363 2162
rect 2407 2158 2411 2162
rect 2095 2086 2099 2090
rect 2111 2086 2115 2090
rect 2167 2086 2171 2090
rect 2175 2086 2179 2090
rect 2239 2086 2243 2090
rect 2311 2086 2315 2090
rect 2359 2086 2363 2090
rect 1919 2010 1923 2014
rect 1935 2010 1939 2014
rect 1999 2010 2003 2014
rect 2015 2010 2019 2014
rect 2071 2010 2075 2014
rect 2095 2010 2099 2014
rect 2135 2010 2139 2014
rect 2167 2010 2171 2014
rect 2191 2010 2195 2014
rect 2239 2010 2243 2014
rect 2255 2010 2259 2014
rect 2311 2010 2315 2014
rect 2319 2010 2323 2014
rect 2407 2086 2411 2090
rect 2359 2010 2363 2014
rect 2407 2010 2411 2014
rect 1751 1942 1755 1946
rect 1791 1942 1795 1946
rect 1839 1942 1843 1946
rect 1863 1942 1867 1946
rect 1919 1942 1923 1946
rect 1935 1942 1939 1946
rect 1999 1942 2003 1946
rect 2007 1942 2011 1946
rect 2071 1942 2075 1946
rect 2079 1942 2083 1946
rect 2135 1942 2139 1946
rect 2151 1942 2155 1946
rect 2191 1942 2195 1946
rect 2223 1942 2227 1946
rect 1279 1874 1283 1878
rect 1303 1874 1307 1878
rect 1311 1874 1315 1878
rect 1359 1874 1363 1878
rect 1415 1874 1419 1878
rect 719 1846 723 1850
rect 727 1846 731 1850
rect 799 1846 803 1850
rect 823 1846 827 1850
rect 879 1846 883 1850
rect 911 1846 915 1850
rect 175 1778 179 1782
rect 215 1778 219 1782
rect 271 1778 275 1782
rect 959 1846 963 1850
rect 991 1846 995 1850
rect 1039 1846 1043 1850
rect 1063 1846 1067 1850
rect 1119 1846 1123 1850
rect 1135 1846 1139 1850
rect 1191 1846 1195 1850
rect 1239 1846 1243 1850
rect 1447 1874 1451 1878
rect 1479 1874 1483 1878
rect 1535 1874 1539 1878
rect 1543 1874 1547 1878
rect 1615 1874 1619 1878
rect 1623 1874 1627 1878
rect 1687 1874 1691 1878
rect 1711 1874 1715 1878
rect 1767 1874 1771 1878
rect 1791 1874 1795 1878
rect 1863 1874 1867 1878
rect 1935 1874 1939 1878
rect 287 1778 291 1782
rect 351 1778 355 1782
rect 375 1778 379 1782
rect 439 1778 443 1782
rect 471 1778 475 1782
rect 535 1778 539 1782
rect 567 1778 571 1782
rect 631 1778 635 1782
rect 663 1778 667 1782
rect 727 1778 731 1782
rect 751 1778 755 1782
rect 823 1778 827 1782
rect 831 1778 835 1782
rect 903 1778 907 1782
rect 911 1778 915 1782
rect 967 1778 971 1782
rect 991 1778 995 1782
rect 1031 1778 1035 1782
rect 111 1706 115 1710
rect 135 1706 139 1710
rect 175 1706 179 1710
rect 215 1706 219 1710
rect 239 1706 243 1710
rect 287 1706 291 1710
rect 319 1706 323 1710
rect 375 1706 379 1710
rect 415 1706 419 1710
rect 471 1706 475 1710
rect 511 1706 515 1710
rect 567 1706 571 1710
rect 615 1706 619 1710
rect 663 1706 667 1710
rect 711 1706 715 1710
rect 751 1706 755 1710
rect 799 1706 803 1710
rect 831 1706 835 1710
rect 879 1706 883 1710
rect 903 1706 907 1710
rect 951 1706 955 1710
rect 967 1706 971 1710
rect 1279 1802 1283 1806
rect 1311 1802 1315 1806
rect 1359 1802 1363 1806
rect 1407 1802 1411 1806
rect 1415 1802 1419 1806
rect 1471 1802 1475 1806
rect 1479 1802 1483 1806
rect 1535 1802 1539 1806
rect 1543 1802 1547 1806
rect 1599 1802 1603 1806
rect 1063 1778 1067 1782
rect 1087 1778 1091 1782
rect 1135 1778 1139 1782
rect 1151 1778 1155 1782
rect 1191 1778 1195 1782
rect 1239 1778 1243 1782
rect 2255 1942 2259 1946
rect 2303 1942 2307 1946
rect 2319 1942 2323 1946
rect 2359 1942 2363 1946
rect 2407 1942 2411 1946
rect 1975 1874 1979 1878
rect 2007 1874 2011 1878
rect 2079 1874 2083 1878
rect 2095 1874 2099 1878
rect 2151 1874 2155 1878
rect 2223 1874 2227 1878
rect 2303 1874 2307 1878
rect 2359 1874 2363 1878
rect 2407 1874 2411 1878
rect 1615 1802 1619 1806
rect 1663 1802 1667 1806
rect 1279 1734 1283 1738
rect 1303 1734 1307 1738
rect 1351 1734 1355 1738
rect 1407 1734 1411 1738
rect 1687 1802 1691 1806
rect 1727 1802 1731 1806
rect 1767 1802 1771 1806
rect 1783 1802 1787 1806
rect 1839 1802 1843 1806
rect 1863 1802 1867 1806
rect 1895 1802 1899 1806
rect 1959 1802 1963 1806
rect 1975 1802 1979 1806
rect 2095 1802 2099 1806
rect 2223 1802 2227 1806
rect 2359 1802 2363 1806
rect 2407 1802 2411 1806
rect 1423 1734 1427 1738
rect 1015 1706 1019 1710
rect 1031 1706 1035 1710
rect 1087 1706 1091 1710
rect 1151 1706 1155 1710
rect 1159 1706 1163 1710
rect 1191 1706 1195 1710
rect 1239 1706 1243 1710
rect 1471 1734 1475 1738
rect 1503 1734 1507 1738
rect 1535 1734 1539 1738
rect 1583 1734 1587 1738
rect 1599 1734 1603 1738
rect 1663 1734 1667 1738
rect 1727 1734 1731 1738
rect 1735 1734 1739 1738
rect 1783 1734 1787 1738
rect 1807 1734 1811 1738
rect 1839 1734 1843 1738
rect 1871 1734 1875 1738
rect 1895 1734 1899 1738
rect 1935 1734 1939 1738
rect 1959 1734 1963 1738
rect 1999 1734 2003 1738
rect 2063 1734 2067 1738
rect 2407 1734 2411 1738
rect 279 1656 283 1660
rect 111 1634 115 1638
rect 135 1634 139 1638
rect 175 1634 179 1638
rect 239 1634 243 1638
rect 271 1634 275 1638
rect 623 1656 627 1660
rect 1279 1666 1283 1670
rect 1303 1666 1307 1670
rect 311 1634 315 1638
rect 319 1634 323 1638
rect 359 1634 363 1638
rect 415 1634 419 1638
rect 471 1634 475 1638
rect 511 1634 515 1638
rect 535 1634 539 1638
rect 599 1634 603 1638
rect 615 1634 619 1638
rect 663 1634 667 1638
rect 711 1634 715 1638
rect 719 1634 723 1638
rect 775 1634 779 1638
rect 799 1634 803 1638
rect 831 1634 835 1638
rect 879 1634 883 1638
rect 887 1634 891 1638
rect 943 1634 947 1638
rect 951 1634 955 1638
rect 999 1634 1003 1638
rect 1015 1634 1019 1638
rect 1087 1634 1091 1638
rect 1159 1634 1163 1638
rect 1239 1634 1243 1638
rect 1351 1666 1355 1670
rect 1359 1666 1363 1670
rect 1423 1666 1427 1670
rect 1447 1666 1451 1670
rect 1503 1666 1507 1670
rect 1543 1666 1547 1670
rect 1583 1666 1587 1670
rect 1639 1666 1643 1670
rect 1663 1666 1667 1670
rect 1727 1666 1731 1670
rect 1735 1666 1739 1670
rect 1807 1666 1811 1670
rect 1815 1666 1819 1670
rect 1279 1598 1283 1602
rect 1303 1598 1307 1602
rect 1327 1598 1331 1602
rect 1359 1598 1363 1602
rect 1399 1598 1403 1602
rect 1447 1598 1451 1602
rect 111 1558 115 1562
rect 271 1558 275 1562
rect 311 1558 315 1562
rect 327 1558 331 1562
rect 359 1558 363 1562
rect 367 1558 371 1562
rect 407 1558 411 1562
rect 415 1558 419 1562
rect 447 1558 451 1562
rect 471 1558 475 1562
rect 487 1558 491 1562
rect 527 1558 531 1562
rect 535 1558 539 1562
rect 567 1558 571 1562
rect 599 1558 603 1562
rect 607 1558 611 1562
rect 647 1558 651 1562
rect 663 1558 667 1562
rect 687 1558 691 1562
rect 719 1558 723 1562
rect 727 1558 731 1562
rect 767 1558 771 1562
rect 775 1558 779 1562
rect 807 1558 811 1562
rect 831 1558 835 1562
rect 847 1558 851 1562
rect 887 1558 891 1562
rect 927 1558 931 1562
rect 943 1558 947 1562
rect 999 1558 1003 1562
rect 1239 1558 1243 1562
rect 1871 1666 1875 1670
rect 1895 1666 1899 1670
rect 1935 1666 1939 1670
rect 1967 1666 1971 1670
rect 1999 1666 2003 1670
rect 2031 1666 2035 1670
rect 2063 1666 2067 1670
rect 2095 1666 2099 1670
rect 2159 1666 2163 1670
rect 2223 1666 2227 1670
rect 2407 1666 2411 1670
rect 1479 1598 1483 1602
rect 1543 1598 1547 1602
rect 1567 1598 1571 1602
rect 1639 1598 1643 1602
rect 1655 1598 1659 1602
rect 1727 1598 1731 1602
rect 1743 1598 1747 1602
rect 1815 1598 1819 1602
rect 1831 1598 1835 1602
rect 1895 1598 1899 1602
rect 1911 1598 1915 1602
rect 1967 1598 1971 1602
rect 1983 1598 1987 1602
rect 2031 1598 2035 1602
rect 2047 1598 2051 1602
rect 2095 1598 2099 1602
rect 2111 1598 2115 1602
rect 2159 1598 2163 1602
rect 2167 1598 2171 1602
rect 2215 1598 2219 1602
rect 2223 1598 2227 1602
rect 2271 1598 2275 1602
rect 2319 1598 2323 1602
rect 2359 1598 2363 1602
rect 2407 1598 2411 1602
rect 1279 1526 1283 1530
rect 1327 1526 1331 1530
rect 1335 1526 1339 1530
rect 1399 1526 1403 1530
rect 1415 1526 1419 1530
rect 1479 1526 1483 1530
rect 1503 1526 1507 1530
rect 1567 1526 1571 1530
rect 1615 1526 1619 1530
rect 1655 1526 1659 1530
rect 1743 1526 1747 1530
rect 1831 1526 1835 1530
rect 1887 1526 1891 1530
rect 1911 1526 1915 1530
rect 1983 1526 1987 1530
rect 2047 1526 2051 1530
rect 2111 1526 2115 1530
rect 2167 1526 2171 1530
rect 2215 1526 2219 1530
rect 1279 1458 1283 1462
rect 1335 1458 1339 1462
rect 1375 1458 1379 1462
rect 1415 1458 1419 1462
rect 1463 1458 1467 1462
rect 111 1450 115 1454
rect 143 1450 147 1454
rect 183 1450 187 1454
rect 223 1450 227 1454
rect 263 1450 267 1454
rect 319 1450 323 1454
rect 327 1450 331 1454
rect 367 1450 371 1454
rect 391 1450 395 1454
rect 407 1450 411 1454
rect 447 1450 451 1454
rect 471 1450 475 1454
rect 487 1450 491 1454
rect 527 1450 531 1454
rect 559 1450 563 1454
rect 567 1450 571 1454
rect 607 1450 611 1454
rect 647 1450 651 1454
rect 687 1450 691 1454
rect 727 1450 731 1454
rect 767 1450 771 1454
rect 807 1450 811 1454
rect 847 1450 851 1454
rect 879 1450 883 1454
rect 887 1450 891 1454
rect 927 1450 931 1454
rect 943 1450 947 1454
rect 999 1450 1003 1454
rect 1047 1450 1051 1454
rect 1103 1450 1107 1454
rect 1151 1450 1155 1454
rect 1191 1450 1195 1454
rect 1239 1450 1243 1454
rect 111 1382 115 1386
rect 143 1382 147 1386
rect 167 1382 171 1386
rect 183 1382 187 1386
rect 207 1382 211 1386
rect 223 1382 227 1386
rect 247 1382 251 1386
rect 263 1382 267 1386
rect 303 1382 307 1386
rect 319 1382 323 1386
rect 367 1382 371 1386
rect 111 1310 115 1314
rect 167 1310 171 1314
rect 279 1320 283 1324
rect 183 1310 187 1314
rect 207 1310 211 1314
rect 231 1310 235 1314
rect 247 1310 251 1314
rect 391 1382 395 1386
rect 439 1382 443 1386
rect 471 1382 475 1386
rect 519 1382 523 1386
rect 559 1382 563 1386
rect 599 1382 603 1386
rect 647 1382 651 1386
rect 679 1382 683 1386
rect 727 1382 731 1386
rect 2271 1526 2275 1530
rect 2319 1526 2323 1530
rect 2359 1526 2363 1530
rect 2407 1526 2411 1530
rect 1503 1458 1507 1462
rect 1551 1458 1555 1462
rect 1615 1458 1619 1462
rect 1639 1458 1643 1462
rect 751 1382 755 1386
rect 807 1382 811 1386
rect 823 1382 827 1386
rect 879 1382 883 1386
rect 887 1382 891 1386
rect 943 1382 947 1386
rect 951 1382 955 1386
rect 999 1382 1003 1386
rect 1015 1382 1019 1386
rect 1047 1382 1051 1386
rect 1079 1382 1083 1386
rect 607 1320 611 1324
rect 1103 1382 1107 1386
rect 1143 1382 1147 1386
rect 1151 1382 1155 1386
rect 1191 1382 1195 1386
rect 1239 1382 1243 1386
rect 1279 1382 1283 1386
rect 1303 1382 1307 1386
rect 1343 1382 1347 1386
rect 287 1310 291 1314
rect 303 1310 307 1314
rect 351 1310 355 1314
rect 367 1310 371 1314
rect 423 1310 427 1314
rect 439 1310 443 1314
rect 495 1310 499 1314
rect 519 1310 523 1314
rect 567 1310 571 1314
rect 599 1310 603 1314
rect 639 1310 643 1314
rect 679 1310 683 1314
rect 703 1310 707 1314
rect 751 1310 755 1314
rect 767 1310 771 1314
rect 823 1310 827 1314
rect 879 1310 883 1314
rect 887 1310 891 1314
rect 935 1310 939 1314
rect 951 1310 955 1314
rect 999 1310 1003 1314
rect 1015 1310 1019 1314
rect 1079 1310 1083 1314
rect 111 1238 115 1242
rect 135 1238 139 1242
rect 175 1238 179 1242
rect 183 1238 187 1242
rect 231 1238 235 1242
rect 287 1238 291 1242
rect 311 1238 315 1242
rect 351 1238 355 1242
rect 399 1238 403 1242
rect 423 1238 427 1242
rect 487 1238 491 1242
rect 495 1238 499 1242
rect 567 1238 571 1242
rect 575 1238 579 1242
rect 111 1170 115 1174
rect 639 1238 643 1242
rect 1143 1310 1147 1314
rect 1191 1310 1195 1314
rect 1239 1310 1243 1314
rect 1279 1314 1283 1318
rect 1303 1314 1307 1318
rect 1375 1382 1379 1386
rect 1399 1382 1403 1386
rect 1463 1382 1467 1386
rect 1535 1382 1539 1386
rect 1551 1382 1555 1386
rect 1727 1458 1731 1462
rect 1743 1458 1747 1462
rect 1807 1458 1811 1462
rect 1879 1458 1883 1462
rect 1887 1458 1891 1462
rect 1943 1458 1947 1462
rect 1999 1458 2003 1462
rect 2047 1458 2051 1462
rect 2095 1458 2099 1462
rect 2143 1458 2147 1462
rect 2191 1458 2195 1462
rect 2215 1458 2219 1462
rect 2239 1458 2243 1462
rect 2279 1458 2283 1462
rect 2319 1458 2323 1462
rect 2359 1458 2363 1462
rect 1607 1382 1611 1386
rect 1639 1382 1643 1386
rect 1687 1382 1691 1386
rect 1727 1382 1731 1386
rect 1767 1382 1771 1386
rect 1807 1382 1811 1386
rect 1847 1382 1851 1386
rect 1879 1382 1883 1386
rect 1935 1382 1939 1386
rect 1943 1382 1947 1386
rect 1999 1382 2003 1386
rect 1343 1314 1347 1318
rect 1383 1314 1387 1318
rect 1399 1314 1403 1318
rect 1423 1314 1427 1318
rect 1463 1314 1467 1318
rect 1503 1314 1507 1318
rect 1535 1314 1539 1318
rect 1543 1314 1547 1318
rect 1583 1314 1587 1318
rect 1607 1314 1611 1318
rect 1623 1314 1627 1318
rect 1679 1314 1683 1318
rect 1687 1314 1691 1318
rect 1735 1314 1739 1318
rect 1767 1314 1771 1318
rect 2023 1382 2027 1386
rect 2047 1382 2051 1386
rect 2095 1382 2099 1386
rect 2111 1382 2115 1386
rect 2143 1382 2147 1386
rect 2191 1382 2195 1386
rect 2199 1382 2203 1386
rect 2239 1382 2243 1386
rect 2279 1382 2283 1386
rect 2287 1382 2291 1386
rect 2407 1458 2411 1462
rect 2319 1382 2323 1386
rect 2359 1382 2363 1386
rect 1791 1314 1795 1318
rect 1847 1314 1851 1318
rect 1903 1314 1907 1318
rect 1935 1314 1939 1318
rect 1967 1314 1971 1318
rect 2023 1314 2027 1318
rect 2039 1314 2043 1318
rect 2111 1314 2115 1318
rect 2119 1314 2123 1318
rect 2199 1314 2203 1318
rect 663 1238 667 1242
rect 703 1238 707 1242
rect 743 1238 747 1242
rect 767 1238 771 1242
rect 815 1238 819 1242
rect 823 1238 827 1242
rect 879 1238 883 1242
rect 935 1238 939 1242
rect 943 1238 947 1242
rect 999 1238 1003 1242
rect 1007 1238 1011 1242
rect 1071 1238 1075 1242
rect 1239 1238 1243 1242
rect 1279 1238 1283 1242
rect 1303 1238 1307 1242
rect 1343 1238 1347 1242
rect 1375 1238 1379 1242
rect 1383 1238 1387 1242
rect 1423 1238 1427 1242
rect 1463 1238 1467 1242
rect 1479 1238 1483 1242
rect 1503 1238 1507 1242
rect 1543 1238 1547 1242
rect 135 1170 139 1174
rect 175 1170 179 1174
rect 231 1170 235 1174
rect 239 1170 243 1174
rect 311 1170 315 1174
rect 327 1170 331 1174
rect 399 1170 403 1174
rect 431 1170 435 1174
rect 487 1170 491 1174
rect 535 1170 539 1174
rect 575 1170 579 1174
rect 639 1170 643 1174
rect 663 1170 667 1174
rect 743 1170 747 1174
rect 815 1170 819 1174
rect 839 1170 843 1174
rect 879 1170 883 1174
rect 919 1170 923 1174
rect 943 1170 947 1174
rect 999 1170 1003 1174
rect 1007 1170 1011 1174
rect 1071 1170 1075 1174
rect 1143 1170 1147 1174
rect 1191 1170 1195 1174
rect 111 1098 115 1102
rect 135 1098 139 1102
rect 175 1098 179 1102
rect 239 1098 243 1102
rect 247 1098 251 1102
rect 327 1098 331 1102
rect 111 1030 115 1034
rect 135 1030 139 1034
rect 175 1030 179 1034
rect 247 1030 251 1034
rect 255 1030 259 1034
rect 327 1030 331 1034
rect 111 962 115 966
rect 175 962 179 966
rect 215 962 219 966
rect 255 962 259 966
rect 415 1098 419 1102
rect 431 1098 435 1102
rect 503 1098 507 1102
rect 535 1098 539 1102
rect 583 1098 587 1102
rect 639 1098 643 1102
rect 663 1098 667 1102
rect 735 1098 739 1102
rect 743 1098 747 1102
rect 1239 1170 1243 1174
rect 1279 1170 1283 1174
rect 1303 1170 1307 1174
rect 1583 1238 1587 1242
rect 1623 1238 1627 1242
rect 1679 1238 1683 1242
rect 1687 1238 1691 1242
rect 1735 1238 1739 1242
rect 1791 1238 1795 1242
rect 1343 1170 1347 1174
rect 1375 1170 1379 1174
rect 1407 1170 1411 1174
rect 1479 1170 1483 1174
rect 1847 1238 1851 1242
rect 1887 1238 1891 1242
rect 1903 1238 1907 1242
rect 1967 1238 1971 1242
rect 1983 1238 1987 1242
rect 2039 1238 2043 1242
rect 2071 1238 2075 1242
rect 2119 1238 2123 1242
rect 2151 1238 2155 1242
rect 2199 1238 2203 1242
rect 2223 1238 2227 1242
rect 2287 1314 2291 1318
rect 2359 1314 2363 1318
rect 2407 1382 2411 1386
rect 2407 1314 2411 1318
rect 2287 1238 2291 1242
rect 2303 1238 2307 1242
rect 2359 1238 2363 1242
rect 1487 1170 1491 1174
rect 1583 1170 1587 1174
rect 1687 1170 1691 1174
rect 1791 1170 1795 1174
rect 1799 1170 1803 1174
rect 1887 1170 1891 1174
rect 1903 1170 1907 1174
rect 1983 1170 1987 1174
rect 1999 1170 2003 1174
rect 2071 1170 2075 1174
rect 2079 1170 2083 1174
rect 2151 1170 2155 1174
rect 2159 1170 2163 1174
rect 2223 1170 2227 1174
rect 2231 1170 2235 1174
rect 2303 1170 2307 1174
rect 2407 1238 2411 1242
rect 2359 1170 2363 1174
rect 2407 1170 2411 1174
rect 799 1098 803 1102
rect 839 1098 843 1102
rect 863 1098 867 1102
rect 919 1098 923 1102
rect 983 1098 987 1102
rect 999 1098 1003 1102
rect 1047 1098 1051 1102
rect 1071 1098 1075 1102
rect 1143 1098 1147 1102
rect 1191 1098 1195 1102
rect 1239 1098 1243 1102
rect 1279 1102 1283 1106
rect 1303 1102 1307 1106
rect 1343 1102 1347 1106
rect 1407 1102 1411 1106
rect 1431 1102 1435 1106
rect 1471 1102 1475 1106
rect 1487 1102 1491 1106
rect 1511 1102 1515 1106
rect 1559 1102 1563 1106
rect 1583 1102 1587 1106
rect 1615 1102 1619 1106
rect 1671 1102 1675 1106
rect 1687 1102 1691 1106
rect 1727 1102 1731 1106
rect 763 1080 767 1084
rect 1071 1080 1075 1084
rect 399 1030 403 1034
rect 415 1030 419 1034
rect 463 1030 467 1034
rect 503 1030 507 1034
rect 519 1030 523 1034
rect 575 1030 579 1034
rect 583 1030 587 1034
rect 623 1030 627 1034
rect 663 1030 667 1034
rect 1439 1064 1443 1068
rect 671 1030 675 1034
rect 303 962 307 966
rect 327 962 331 966
rect 359 962 363 966
rect 399 962 403 966
rect 415 962 419 966
rect 463 962 467 966
rect 519 962 523 966
rect 575 962 579 966
rect 623 962 627 966
rect 735 1030 739 1034
rect 799 1030 803 1034
rect 807 1030 811 1034
rect 863 1030 867 1034
rect 895 1030 899 1034
rect 919 1030 923 1034
rect 983 1030 987 1034
rect 999 1030 1003 1034
rect 1047 1030 1051 1034
rect 1103 1030 1107 1034
rect 1191 1030 1195 1034
rect 1239 1030 1243 1034
rect 1279 1034 1283 1038
rect 1431 1034 1435 1038
rect 1471 1034 1475 1038
rect 1511 1034 1515 1038
rect 1559 1034 1563 1038
rect 1575 1034 1579 1038
rect 719 992 723 996
rect 1127 992 1131 996
rect 639 962 643 966
rect 671 962 675 966
rect 711 962 715 966
rect 735 962 739 966
rect 783 962 787 966
rect 807 962 811 966
rect 855 962 859 966
rect 895 962 899 966
rect 927 962 931 966
rect 999 962 1003 966
rect 1071 962 1075 966
rect 1103 962 1107 966
rect 1143 962 1147 966
rect 111 886 115 890
rect 191 886 195 890
rect 215 886 219 890
rect 231 886 235 890
rect 255 886 259 890
rect 287 886 291 890
rect 111 818 115 822
rect 135 818 139 822
rect 175 818 179 822
rect 191 818 195 822
rect 231 818 235 822
rect 239 818 243 822
rect 303 886 307 890
rect 359 886 363 890
rect 415 886 419 890
rect 447 886 451 890
rect 463 886 467 890
rect 519 886 523 890
rect 543 886 547 890
rect 575 886 579 890
rect 639 886 643 890
rect 711 886 715 890
rect 727 886 731 890
rect 783 886 787 890
rect 807 886 811 890
rect 855 886 859 890
rect 887 886 891 890
rect 927 886 931 890
rect 959 886 963 890
rect 999 886 1003 890
rect 1191 962 1195 966
rect 1775 1102 1779 1106
rect 1799 1102 1803 1106
rect 1823 1102 1827 1106
rect 1871 1102 1875 1106
rect 1903 1102 1907 1106
rect 1919 1102 1923 1106
rect 1967 1102 1971 1106
rect 1999 1102 2003 1106
rect 2015 1102 2019 1106
rect 2063 1102 2067 1106
rect 2079 1102 2083 1106
rect 2119 1102 2123 1106
rect 2159 1102 2163 1106
rect 1735 1064 1739 1068
rect 1615 1034 1619 1038
rect 1655 1034 1659 1038
rect 1671 1034 1675 1038
rect 1695 1034 1699 1038
rect 1727 1034 1731 1038
rect 1735 1034 1739 1038
rect 1775 1034 1779 1038
rect 2175 1102 2179 1106
rect 2231 1102 2235 1106
rect 2303 1102 2307 1106
rect 2359 1102 2363 1106
rect 2407 1102 2411 1106
rect 1823 1034 1827 1038
rect 1871 1034 1875 1038
rect 1879 1034 1883 1038
rect 1919 1034 1923 1038
rect 1943 1034 1947 1038
rect 1967 1034 1971 1038
rect 2015 1034 2019 1038
rect 2063 1034 2067 1038
rect 2095 1034 2099 1038
rect 2119 1034 2123 1038
rect 2175 1034 2179 1038
rect 2231 1034 2235 1038
rect 1239 962 1243 966
rect 1279 958 1283 962
rect 1303 958 1307 962
rect 1351 958 1355 962
rect 1431 958 1435 962
rect 1511 958 1515 962
rect 1575 958 1579 962
rect 1591 958 1595 962
rect 1615 958 1619 962
rect 1655 958 1659 962
rect 1679 958 1683 962
rect 1023 886 1027 890
rect 1071 886 1075 890
rect 1087 886 1091 890
rect 1143 886 1147 890
rect 1159 886 1163 890
rect 1191 886 1195 890
rect 1239 886 1243 890
rect 1279 890 1283 894
rect 1303 890 1307 894
rect 1351 890 1355 894
rect 1431 890 1435 894
rect 1439 890 1443 894
rect 1479 890 1483 894
rect 1511 890 1515 894
rect 1519 890 1523 894
rect 1559 890 1563 894
rect 287 818 291 822
rect 327 818 331 822
rect 359 818 363 822
rect 415 818 419 822
rect 447 818 451 822
rect 503 818 507 822
rect 543 818 547 822
rect 591 818 595 822
rect 639 818 643 822
rect 671 818 675 822
rect 727 818 731 822
rect 743 818 747 822
rect 807 818 811 822
rect 815 818 819 822
rect 111 746 115 750
rect 135 746 139 750
rect 175 746 179 750
rect 191 746 195 750
rect 239 746 243 750
rect 263 746 267 750
rect 327 746 331 750
rect 335 746 339 750
rect 399 746 403 750
rect 415 746 419 750
rect 455 746 459 750
rect 503 746 507 750
rect 543 746 547 750
rect 583 746 587 750
rect 591 746 595 750
rect 623 746 627 750
rect 671 746 675 750
rect 719 746 723 750
rect 743 746 747 750
rect 767 746 771 750
rect 111 674 115 678
rect 135 674 139 678
rect 191 674 195 678
rect 199 674 203 678
rect 263 674 267 678
rect 279 674 283 678
rect 111 598 115 602
rect 135 598 139 602
rect 335 674 339 678
rect 351 674 355 678
rect 399 674 403 678
rect 415 674 419 678
rect 455 674 459 678
rect 487 674 491 678
rect 503 674 507 678
rect 543 674 547 678
rect 559 674 563 678
rect 583 674 587 678
rect 623 674 627 678
rect 639 674 643 678
rect 879 818 883 822
rect 887 818 891 822
rect 943 818 947 822
rect 959 818 963 822
rect 1015 818 1019 822
rect 1023 818 1027 822
rect 1087 818 1091 822
rect 1159 818 1163 822
rect 1239 818 1243 822
rect 1279 810 1283 814
rect 1359 810 1363 814
rect 1415 810 1419 814
rect 1439 810 1443 814
rect 1591 890 1595 894
rect 1607 890 1611 894
rect 1695 958 1699 962
rect 1735 958 1739 962
rect 1767 958 1771 962
rect 1775 958 1779 962
rect 1823 958 1827 962
rect 1855 958 1859 962
rect 1879 958 1883 962
rect 1943 958 1947 962
rect 2015 958 2019 962
rect 2023 958 2027 962
rect 2095 958 2099 962
rect 2103 958 2107 962
rect 2255 1034 2259 1038
rect 2407 1034 2411 1038
rect 2175 958 2179 962
rect 2183 958 2187 962
rect 1655 890 1659 894
rect 1679 890 1683 894
rect 1711 890 1715 894
rect 1767 890 1771 894
rect 1775 890 1779 894
rect 1847 890 1851 894
rect 1855 890 1859 894
rect 1919 890 1923 894
rect 1943 890 1947 894
rect 1991 890 1995 894
rect 2023 890 2027 894
rect 2255 958 2259 962
rect 2271 958 2275 962
rect 2407 958 2411 962
rect 2063 890 2067 894
rect 2103 890 2107 894
rect 2135 890 2139 894
rect 2183 890 2187 894
rect 2215 890 2219 894
rect 2271 890 2275 894
rect 2295 890 2299 894
rect 2407 890 2411 894
rect 1471 810 1475 814
rect 1479 810 1483 814
rect 1519 810 1523 814
rect 1535 810 1539 814
rect 1559 810 1563 814
rect 1591 810 1595 814
rect 1607 810 1611 814
rect 1647 810 1651 814
rect 1655 810 1659 814
rect 1703 810 1707 814
rect 1711 810 1715 814
rect 815 746 819 750
rect 863 746 867 750
rect 879 746 883 750
rect 911 746 915 750
rect 943 746 947 750
rect 1015 746 1019 750
rect 1239 746 1243 750
rect 1279 742 1283 746
rect 1303 742 1307 746
rect 1343 742 1347 746
rect 1359 742 1363 746
rect 671 674 675 678
rect 711 674 715 678
rect 719 674 723 678
rect 767 674 771 678
rect 783 674 787 678
rect 191 598 195 602
rect 199 598 203 602
rect 271 598 275 602
rect 279 598 283 602
rect 351 598 355 602
rect 359 598 363 602
rect 415 598 419 602
rect 447 598 451 602
rect 487 598 491 602
rect 535 598 539 602
rect 559 598 563 602
rect 111 522 115 526
rect 135 522 139 526
rect 191 522 195 526
rect 263 522 267 526
rect 271 522 275 526
rect 815 674 819 678
rect 855 674 859 678
rect 863 674 867 678
rect 911 674 915 678
rect 919 674 923 678
rect 983 674 987 678
rect 1039 674 1043 678
rect 1095 674 1099 678
rect 1151 674 1155 678
rect 1191 674 1195 678
rect 1239 674 1243 678
rect 1279 670 1283 674
rect 1303 670 1307 674
rect 1407 742 1411 746
rect 1415 742 1419 746
rect 1471 742 1475 746
rect 1487 742 1491 746
rect 1535 742 1539 746
rect 1575 742 1579 746
rect 1591 742 1595 746
rect 1647 742 1651 746
rect 1663 742 1667 746
rect 1759 810 1763 814
rect 1775 810 1779 814
rect 1815 810 1819 814
rect 1847 810 1851 814
rect 1871 810 1875 814
rect 1919 810 1923 814
rect 1935 810 1939 814
rect 1991 810 1995 814
rect 1999 810 2003 814
rect 2063 810 2067 814
rect 2071 810 2075 814
rect 2135 810 2139 814
rect 2143 810 2147 814
rect 2215 810 2219 814
rect 2223 810 2227 814
rect 2295 810 2299 814
rect 2303 810 2307 814
rect 2359 810 2363 814
rect 2407 810 2411 814
rect 1839 760 1843 764
rect 1703 742 1707 746
rect 1751 742 1755 746
rect 1759 742 1763 746
rect 1815 742 1819 746
rect 1831 742 1835 746
rect 2151 760 2155 764
rect 1871 742 1875 746
rect 1911 742 1915 746
rect 1935 742 1939 746
rect 1991 742 1995 746
rect 1999 742 2003 746
rect 2071 742 2075 746
rect 2079 742 2083 746
rect 2143 742 2147 746
rect 2175 742 2179 746
rect 2223 742 2227 746
rect 2279 742 2283 746
rect 1343 670 1347 674
rect 1399 670 1403 674
rect 1407 670 1411 674
rect 1487 670 1491 674
rect 1511 670 1515 674
rect 1575 670 1579 674
rect 1623 670 1627 674
rect 1663 670 1667 674
rect 1727 670 1731 674
rect 623 598 627 602
rect 639 598 643 602
rect 703 598 707 602
rect 711 598 715 602
rect 783 598 787 602
rect 855 598 859 602
rect 335 522 339 526
rect 359 522 363 526
rect 415 522 419 526
rect 447 522 451 526
rect 495 522 499 526
rect 535 522 539 526
rect 111 454 115 458
rect 135 454 139 458
rect 183 454 187 458
rect 191 454 195 458
rect 223 454 227 458
rect 263 454 267 458
rect 311 454 315 458
rect 335 454 339 458
rect 111 386 115 390
rect 135 386 139 390
rect 175 386 179 390
rect 183 386 187 390
rect 223 386 227 390
rect 231 386 235 390
rect 263 386 267 390
rect 287 386 291 390
rect 575 522 579 526
rect 623 522 627 526
rect 647 522 651 526
rect 703 522 707 526
rect 719 522 723 526
rect 783 522 787 526
rect 919 598 923 602
rect 975 598 979 602
rect 983 598 987 602
rect 1023 598 1027 602
rect 1039 598 1043 602
rect 1079 598 1083 602
rect 1095 598 1099 602
rect 1135 598 1139 602
rect 1151 598 1155 602
rect 1191 598 1195 602
rect 1239 598 1243 602
rect 1279 598 1283 602
rect 1303 598 1307 602
rect 1399 598 1403 602
rect 1415 598 1419 602
rect 1455 598 1459 602
rect 1495 598 1499 602
rect 1511 598 1515 602
rect 1543 598 1547 602
rect 903 560 907 564
rect 1215 560 1219 564
rect 1751 670 1755 674
rect 1815 670 1819 674
rect 1831 670 1835 674
rect 1895 670 1899 674
rect 1911 670 1915 674
rect 1975 670 1979 674
rect 1991 670 1995 674
rect 2047 670 2051 674
rect 2079 670 2083 674
rect 2111 670 2115 674
rect 2175 670 2179 674
rect 2239 670 2243 674
rect 1599 598 1603 602
rect 1623 598 1627 602
rect 1663 598 1667 602
rect 1727 598 1731 602
rect 1791 598 1795 602
rect 1815 598 1819 602
rect 1847 598 1851 602
rect 1895 598 1899 602
rect 1911 598 1915 602
rect 1975 598 1979 602
rect 2279 670 2283 674
rect 2303 742 2307 746
rect 2359 742 2363 746
rect 2407 742 2411 746
rect 2311 670 2315 674
rect 2359 670 2363 674
rect 2047 598 2051 602
rect 2111 598 2115 602
rect 2119 598 2123 602
rect 2175 598 2179 602
rect 2199 598 2203 602
rect 2239 598 2243 602
rect 2287 598 2291 602
rect 1279 530 1283 534
rect 1303 530 1307 534
rect 1375 530 1379 534
rect 1415 530 1419 534
rect 1455 530 1459 534
rect 1479 530 1483 534
rect 1495 530 1499 534
rect 1543 530 1547 534
rect 847 522 851 526
rect 855 522 859 526
rect 903 522 907 526
rect 919 522 923 526
rect 959 522 963 526
rect 975 522 979 526
rect 1023 522 1027 526
rect 1079 522 1083 526
rect 1087 522 1091 526
rect 1135 522 1139 526
rect 1151 522 1155 526
rect 1191 522 1195 526
rect 1239 522 1243 526
rect 367 454 371 458
rect 415 454 419 458
rect 431 454 435 458
rect 495 454 499 458
rect 559 454 563 458
rect 575 454 579 458
rect 615 454 619 458
rect 647 454 651 458
rect 671 454 675 458
rect 311 386 315 390
rect 343 386 347 390
rect 367 386 371 390
rect 391 386 395 390
rect 431 386 435 390
rect 439 386 443 390
rect 111 314 115 318
rect 135 314 139 318
rect 175 314 179 318
rect 183 314 187 318
rect 231 314 235 318
rect 255 314 259 318
rect 287 314 291 318
rect 111 238 115 242
rect 135 238 139 242
rect 327 314 331 318
rect 487 386 491 390
rect 495 386 499 390
rect 535 386 539 390
rect 559 386 563 390
rect 719 454 723 458
rect 775 454 779 458
rect 783 454 787 458
rect 831 454 835 458
rect 847 454 851 458
rect 887 454 891 458
rect 903 454 907 458
rect 959 454 963 458
rect 1023 454 1027 458
rect 1087 454 1091 458
rect 1151 454 1155 458
rect 1191 454 1195 458
rect 1239 454 1243 458
rect 1279 458 1283 462
rect 1303 458 1307 462
rect 1583 530 1587 534
rect 1599 530 1603 534
rect 1663 530 1667 534
rect 1695 530 1699 534
rect 1727 530 1731 534
rect 1791 530 1795 534
rect 1799 530 1803 534
rect 1847 530 1851 534
rect 1343 458 1347 462
rect 1375 458 1379 462
rect 1399 458 1403 462
rect 1463 458 1467 462
rect 1479 458 1483 462
rect 1527 458 1531 462
rect 1583 458 1587 462
rect 1591 458 1595 462
rect 1663 458 1667 462
rect 1695 458 1699 462
rect 1903 530 1907 534
rect 1911 530 1915 534
rect 1975 530 1979 534
rect 2007 530 2011 534
rect 2047 530 2051 534
rect 2103 530 2107 534
rect 2119 530 2123 534
rect 2191 530 2195 534
rect 2199 530 2203 534
rect 2287 530 2291 534
rect 2311 598 2315 602
rect 2359 598 2363 602
rect 2407 670 2411 674
rect 2407 598 2411 602
rect 2359 530 2363 534
rect 1735 458 1739 462
rect 1799 458 1803 462
rect 1815 458 1819 462
rect 1895 458 1899 462
rect 1903 458 1907 462
rect 1975 458 1979 462
rect 2007 458 2011 462
rect 2055 458 2059 462
rect 2103 458 2107 462
rect 2135 458 2139 462
rect 583 386 587 390
rect 615 386 619 390
rect 631 386 635 390
rect 671 386 675 390
rect 679 386 683 390
rect 719 386 723 390
rect 727 386 731 390
rect 775 386 779 390
rect 831 386 835 390
rect 887 386 891 390
rect 1239 386 1243 390
rect 1279 386 1283 390
rect 1303 386 1307 390
rect 1343 386 1347 390
rect 1399 386 1403 390
rect 1447 386 1451 390
rect 1463 386 1467 390
rect 1487 386 1491 390
rect 1527 386 1531 390
rect 1535 386 1539 390
rect 1591 386 1595 390
rect 1663 386 1667 390
rect 1735 386 1739 390
rect 1815 386 1819 390
rect 1895 386 1899 390
rect 1967 386 1971 390
rect 1975 386 1979 390
rect 2039 386 2043 390
rect 2055 386 2059 390
rect 2191 458 2195 462
rect 2215 458 2219 462
rect 2287 458 2291 462
rect 2295 458 2299 462
rect 2359 458 2363 462
rect 2407 530 2411 534
rect 2407 458 2411 462
rect 2111 386 2115 390
rect 2135 386 2139 390
rect 2175 386 2179 390
rect 2215 386 2219 390
rect 2239 386 2243 390
rect 2295 386 2299 390
rect 2303 386 2307 390
rect 343 314 347 318
rect 391 314 395 318
rect 439 314 443 318
rect 447 314 451 318
rect 487 314 491 318
rect 503 314 507 318
rect 535 314 539 318
rect 551 314 555 318
rect 583 314 587 318
rect 591 314 595 318
rect 631 314 635 318
rect 679 314 683 318
rect 727 314 731 318
rect 775 314 779 318
rect 823 314 827 318
rect 871 314 875 318
rect 919 314 923 318
rect 1239 314 1243 318
rect 1279 314 1283 318
rect 1447 314 1451 318
rect 1487 314 1491 318
rect 1495 314 1499 318
rect 1535 314 1539 318
rect 1575 314 1579 318
rect 1591 314 1595 318
rect 1615 314 1619 318
rect 1655 314 1659 318
rect 1663 314 1667 318
rect 1695 314 1699 318
rect 1735 314 1739 318
rect 1743 314 1747 318
rect 1799 314 1803 318
rect 1815 314 1819 318
rect 1863 314 1867 318
rect 1895 314 1899 318
rect 1935 314 1939 318
rect 1967 314 1971 318
rect 2007 314 2011 318
rect 2039 314 2043 318
rect 2071 314 2075 318
rect 2111 314 2115 318
rect 2135 314 2139 318
rect 2175 314 2179 318
rect 2191 314 2195 318
rect 2239 314 2243 318
rect 2255 314 2259 318
rect 175 238 179 242
rect 183 238 187 242
rect 247 238 251 242
rect 255 238 259 242
rect 327 238 331 242
rect 391 238 395 242
rect 415 238 419 242
rect 447 238 451 242
rect 495 238 499 242
rect 503 238 507 242
rect 551 238 555 242
rect 111 150 115 154
rect 135 150 139 154
rect 175 150 179 154
rect 215 150 219 154
rect 247 150 251 154
rect 255 150 259 154
rect 295 150 299 154
rect 327 150 331 154
rect 335 150 339 154
rect 375 150 379 154
rect 415 150 419 154
rect 423 150 427 154
rect 471 150 475 154
rect 495 150 499 154
rect 575 238 579 242
rect 591 238 595 242
rect 631 238 635 242
rect 655 238 659 242
rect 679 238 683 242
rect 727 238 731 242
rect 775 238 779 242
rect 791 238 795 242
rect 823 238 827 242
rect 847 238 851 242
rect 871 238 875 242
rect 903 238 907 242
rect 919 238 923 242
rect 959 238 963 242
rect 1023 238 1027 242
rect 1239 238 1243 242
rect 1279 242 1283 246
rect 1367 242 1371 246
rect 1407 242 1411 246
rect 1447 242 1451 246
rect 1495 242 1499 246
rect 1535 242 1539 246
rect 1551 242 1555 246
rect 1575 242 1579 246
rect 1607 242 1611 246
rect 1615 242 1619 246
rect 1655 242 1659 246
rect 1671 242 1675 246
rect 1695 242 1699 246
rect 527 150 531 154
rect 575 150 579 154
rect 583 150 587 154
rect 631 150 635 154
rect 655 150 659 154
rect 679 150 683 154
rect 727 150 731 154
rect 1279 158 1283 162
rect 1303 158 1307 162
rect 1343 158 1347 162
rect 1367 158 1371 162
rect 1383 158 1387 162
rect 1407 158 1411 162
rect 1423 158 1427 162
rect 1447 158 1451 162
rect 1463 158 1467 162
rect 1495 158 1499 162
rect 767 150 771 154
rect 791 150 795 154
rect 807 150 811 154
rect 847 150 851 154
rect 887 150 891 154
rect 903 150 907 154
rect 927 150 931 154
rect 959 150 963 154
rect 975 150 979 154
rect 1023 150 1027 154
rect 1071 150 1075 154
rect 1111 150 1115 154
rect 1151 150 1155 154
rect 1191 150 1195 154
rect 1239 150 1243 154
rect 1735 242 1739 246
rect 1743 242 1747 246
rect 1799 242 1803 246
rect 1807 242 1811 246
rect 1863 242 1867 246
rect 1887 242 1891 246
rect 1935 242 1939 246
rect 1975 242 1979 246
rect 1743 184 1747 188
rect 2007 242 2011 246
rect 2071 242 2075 246
rect 2303 314 2307 318
rect 2319 314 2323 318
rect 2359 386 2363 390
rect 2407 386 2411 390
rect 2359 314 2363 318
rect 2407 314 2411 318
rect 2135 242 2139 246
rect 2167 242 2171 246
rect 2191 242 2195 246
rect 2255 242 2259 246
rect 2271 242 2275 246
rect 2319 242 2323 246
rect 2359 242 2363 246
rect 1983 184 1987 188
rect 1519 158 1523 162
rect 1551 158 1555 162
rect 1583 158 1587 162
rect 1607 158 1611 162
rect 1647 158 1651 162
rect 1671 158 1675 162
rect 1711 158 1715 162
rect 1735 158 1739 162
rect 1767 158 1771 162
rect 1807 158 1811 162
rect 1823 158 1827 162
rect 1871 158 1875 162
rect 1887 158 1891 162
rect 1919 158 1923 162
rect 1967 158 1971 162
rect 1975 158 1979 162
rect 2015 158 2019 162
rect 2063 158 2067 162
rect 2071 158 2075 162
rect 2111 158 2115 162
rect 2159 158 2163 162
rect 2167 158 2171 162
rect 2215 158 2219 162
rect 2271 158 2275 162
rect 2319 158 2323 162
rect 2359 158 2363 162
rect 2407 242 2411 246
rect 2407 158 2411 162
rect 1279 90 1283 94
rect 1303 90 1307 94
rect 1343 90 1347 94
rect 1383 90 1387 94
rect 1423 90 1427 94
rect 1463 90 1467 94
rect 1519 90 1523 94
rect 1583 90 1587 94
rect 1647 90 1651 94
rect 1711 90 1715 94
rect 1767 90 1771 94
rect 1823 90 1827 94
rect 1871 90 1875 94
rect 1919 90 1923 94
rect 1967 90 1971 94
rect 2015 90 2019 94
rect 2063 90 2067 94
rect 2111 90 2115 94
rect 2159 90 2163 94
rect 2215 90 2219 94
rect 2271 90 2275 94
rect 2319 90 2323 94
rect 2359 90 2363 94
rect 2407 90 2411 94
rect 111 82 115 86
rect 135 82 139 86
rect 175 82 179 86
rect 215 82 219 86
rect 255 82 259 86
rect 295 82 299 86
rect 335 82 339 86
rect 375 82 379 86
rect 423 82 427 86
rect 471 82 475 86
rect 527 82 531 86
rect 583 82 587 86
rect 631 82 635 86
rect 679 82 683 86
rect 727 82 731 86
rect 767 82 771 86
rect 807 82 811 86
rect 847 82 851 86
rect 887 82 891 86
rect 927 82 931 86
rect 975 82 979 86
rect 1023 82 1027 86
rect 1071 82 1075 86
rect 1111 82 1115 86
rect 1151 82 1155 86
rect 1191 82 1195 86
rect 1239 82 1243 86
<< m4 >>
rect 1250 2509 1251 2515
rect 1257 2514 2435 2515
rect 1257 2510 1279 2514
rect 1283 2510 1535 2514
rect 1539 2510 1575 2514
rect 1579 2510 1615 2514
rect 1619 2510 1655 2514
rect 1659 2510 1695 2514
rect 1699 2510 1735 2514
rect 1739 2510 1775 2514
rect 1779 2510 1815 2514
rect 1819 2510 1855 2514
rect 1859 2510 1895 2514
rect 1899 2510 1935 2514
rect 1939 2510 1975 2514
rect 1979 2510 2407 2514
rect 2411 2510 2435 2514
rect 1257 2509 2435 2510
rect 2441 2509 2442 2515
rect 96 2497 97 2503
rect 103 2502 1263 2503
rect 103 2498 111 2502
rect 115 2498 135 2502
rect 139 2498 175 2502
rect 179 2498 215 2502
rect 219 2498 255 2502
rect 259 2498 311 2502
rect 315 2498 391 2502
rect 395 2498 479 2502
rect 483 2498 567 2502
rect 571 2498 655 2502
rect 659 2498 743 2502
rect 747 2498 831 2502
rect 835 2498 927 2502
rect 931 2498 1239 2502
rect 1243 2498 1263 2502
rect 103 2497 1263 2498
rect 1269 2497 1270 2503
rect 1262 2441 1263 2447
rect 1269 2446 2447 2447
rect 1269 2442 1279 2446
rect 1283 2442 1359 2446
rect 1363 2442 1399 2446
rect 1403 2442 1455 2446
rect 1459 2442 1519 2446
rect 1523 2442 1535 2446
rect 1539 2442 1575 2446
rect 1579 2442 1599 2446
rect 1603 2442 1615 2446
rect 1619 2442 1655 2446
rect 1659 2442 1679 2446
rect 1683 2442 1695 2446
rect 1699 2442 1735 2446
rect 1739 2442 1759 2446
rect 1763 2442 1775 2446
rect 1779 2442 1815 2446
rect 1819 2442 1839 2446
rect 1843 2442 1855 2446
rect 1859 2442 1895 2446
rect 1899 2442 1919 2446
rect 1923 2442 1935 2446
rect 1939 2442 1975 2446
rect 1979 2442 1999 2446
rect 2003 2442 2079 2446
rect 2083 2442 2159 2446
rect 2163 2442 2247 2446
rect 2251 2442 2335 2446
rect 2339 2442 2407 2446
rect 2411 2442 2447 2446
rect 1269 2441 2447 2442
rect 2453 2441 2454 2447
rect 84 2429 85 2435
rect 91 2434 1251 2435
rect 91 2430 111 2434
rect 115 2430 135 2434
rect 139 2430 175 2434
rect 179 2430 183 2434
rect 187 2430 215 2434
rect 219 2430 247 2434
rect 251 2430 255 2434
rect 259 2430 311 2434
rect 315 2430 319 2434
rect 323 2430 391 2434
rect 395 2430 471 2434
rect 475 2430 479 2434
rect 483 2430 543 2434
rect 547 2430 567 2434
rect 571 2430 615 2434
rect 619 2430 655 2434
rect 659 2430 679 2434
rect 683 2430 735 2434
rect 739 2430 743 2434
rect 747 2430 791 2434
rect 795 2430 831 2434
rect 835 2430 839 2434
rect 843 2430 887 2434
rect 891 2430 927 2434
rect 931 2430 935 2434
rect 939 2430 991 2434
rect 995 2430 1047 2434
rect 1051 2430 1239 2434
rect 1243 2430 1251 2434
rect 91 2429 1251 2430
rect 1257 2429 1258 2435
rect 1250 2373 1251 2379
rect 1257 2378 2435 2379
rect 1257 2374 1279 2378
rect 1283 2374 1359 2378
rect 1363 2374 1399 2378
rect 1403 2374 1407 2378
rect 1411 2374 1455 2378
rect 1459 2374 1471 2378
rect 1475 2374 1519 2378
rect 1523 2374 1543 2378
rect 1547 2374 1599 2378
rect 1603 2374 1615 2378
rect 1619 2374 1679 2378
rect 1683 2374 1695 2378
rect 1699 2374 1759 2378
rect 1763 2374 1775 2378
rect 1779 2374 1839 2378
rect 1843 2374 1855 2378
rect 1859 2374 1919 2378
rect 1923 2374 1927 2378
rect 1931 2374 1999 2378
rect 2003 2374 2071 2378
rect 2075 2374 2079 2378
rect 2083 2374 2143 2378
rect 2147 2374 2159 2378
rect 2163 2374 2223 2378
rect 2227 2374 2247 2378
rect 2251 2374 2303 2378
rect 2307 2374 2335 2378
rect 2339 2374 2359 2378
rect 2363 2374 2407 2378
rect 2411 2374 2435 2378
rect 1257 2373 2435 2374
rect 2441 2373 2442 2379
rect 96 2353 97 2359
rect 103 2358 1263 2359
rect 103 2354 111 2358
rect 115 2354 135 2358
rect 139 2354 175 2358
rect 179 2354 183 2358
rect 187 2354 215 2358
rect 219 2354 247 2358
rect 251 2354 271 2358
rect 275 2354 319 2358
rect 323 2354 351 2358
rect 355 2354 391 2358
rect 395 2354 431 2358
rect 435 2354 471 2358
rect 475 2354 519 2358
rect 523 2354 543 2358
rect 547 2354 599 2358
rect 603 2354 615 2358
rect 619 2354 679 2358
rect 683 2354 735 2358
rect 739 2354 751 2358
rect 755 2354 791 2358
rect 795 2354 823 2358
rect 827 2354 839 2358
rect 843 2354 887 2358
rect 891 2354 935 2358
rect 939 2354 959 2358
rect 963 2354 991 2358
rect 995 2354 1031 2358
rect 1035 2354 1047 2358
rect 1051 2354 1239 2358
rect 1243 2354 1263 2358
rect 103 2353 1263 2354
rect 1269 2353 1270 2359
rect 1262 2301 1263 2307
rect 1269 2306 2447 2307
rect 1269 2302 1279 2306
rect 1283 2302 1359 2306
rect 1363 2302 1407 2306
rect 1411 2302 1471 2306
rect 1475 2302 1503 2306
rect 1507 2302 1543 2306
rect 1547 2302 1583 2306
rect 1587 2302 1615 2306
rect 1619 2302 1623 2306
rect 1627 2302 1663 2306
rect 1667 2302 1695 2306
rect 1699 2302 1703 2306
rect 1707 2302 1759 2306
rect 1763 2302 1775 2306
rect 1779 2302 1823 2306
rect 1827 2302 1855 2306
rect 1859 2302 1895 2306
rect 1899 2302 1927 2306
rect 1931 2302 1967 2306
rect 1971 2302 1999 2306
rect 2003 2302 2047 2306
rect 2051 2302 2071 2306
rect 2075 2302 2127 2306
rect 2131 2302 2143 2306
rect 2147 2302 2207 2306
rect 2211 2302 2223 2306
rect 2227 2302 2295 2306
rect 2299 2302 2303 2306
rect 2307 2302 2359 2306
rect 2363 2302 2407 2306
rect 2411 2302 2447 2306
rect 1269 2301 2447 2302
rect 2453 2301 2454 2307
rect 84 2281 85 2287
rect 91 2286 1251 2287
rect 91 2282 111 2286
rect 115 2282 135 2286
rect 139 2282 175 2286
rect 179 2282 215 2286
rect 219 2282 231 2286
rect 235 2282 271 2286
rect 275 2282 303 2286
rect 307 2282 351 2286
rect 355 2282 375 2286
rect 379 2282 431 2286
rect 435 2282 455 2286
rect 459 2282 519 2286
rect 523 2282 535 2286
rect 539 2282 599 2286
rect 603 2282 615 2286
rect 619 2282 679 2286
rect 683 2282 687 2286
rect 691 2282 751 2286
rect 755 2282 759 2286
rect 763 2282 823 2286
rect 827 2282 831 2286
rect 835 2282 887 2286
rect 891 2282 911 2286
rect 915 2282 959 2286
rect 963 2282 991 2286
rect 995 2282 1031 2286
rect 1035 2282 1239 2286
rect 1243 2282 1251 2286
rect 91 2281 1251 2282
rect 1257 2281 1258 2287
rect 1250 2225 1251 2231
rect 1257 2230 2435 2231
rect 1257 2226 1279 2230
rect 1283 2226 1303 2230
rect 1307 2226 1343 2230
rect 1347 2226 1383 2230
rect 1387 2226 1431 2230
rect 1435 2226 1495 2230
rect 1499 2226 1503 2230
rect 1507 2226 1543 2230
rect 1547 2226 1567 2230
rect 1571 2226 1583 2230
rect 1587 2226 1623 2230
rect 1627 2226 1639 2230
rect 1643 2226 1663 2230
rect 1667 2226 1703 2230
rect 1707 2226 1711 2230
rect 1715 2226 1759 2230
rect 1763 2226 1783 2230
rect 1787 2226 1823 2230
rect 1827 2226 1855 2230
rect 1859 2226 1895 2230
rect 1899 2226 1935 2230
rect 1939 2226 1967 2230
rect 1971 2226 2015 2230
rect 2019 2226 2047 2230
rect 2051 2226 2095 2230
rect 2099 2226 2127 2230
rect 2131 2226 2183 2230
rect 2187 2226 2207 2230
rect 2211 2226 2279 2230
rect 2283 2226 2295 2230
rect 2299 2226 2359 2230
rect 2363 2226 2407 2230
rect 2411 2226 2435 2230
rect 1257 2225 2435 2226
rect 2441 2225 2442 2231
rect 96 2213 97 2219
rect 103 2218 1263 2219
rect 103 2214 111 2218
rect 115 2214 135 2218
rect 139 2214 175 2218
rect 179 2214 231 2218
rect 235 2214 247 2218
rect 251 2214 287 2218
rect 291 2214 303 2218
rect 307 2214 327 2218
rect 331 2214 375 2218
rect 379 2214 431 2218
rect 435 2214 455 2218
rect 459 2214 495 2218
rect 499 2214 535 2218
rect 539 2214 551 2218
rect 555 2214 607 2218
rect 611 2214 615 2218
rect 619 2214 663 2218
rect 667 2214 687 2218
rect 691 2214 719 2218
rect 723 2214 759 2218
rect 763 2214 783 2218
rect 787 2214 831 2218
rect 835 2214 847 2218
rect 851 2214 911 2218
rect 915 2214 991 2218
rect 995 2214 1239 2218
rect 1243 2214 1263 2218
rect 103 2213 1263 2214
rect 1269 2213 1270 2219
rect 1262 2157 1263 2163
rect 1269 2162 2447 2163
rect 1269 2158 1279 2162
rect 1283 2158 1303 2162
rect 1307 2158 1343 2162
rect 1347 2158 1351 2162
rect 1355 2158 1383 2162
rect 1387 2158 1431 2162
rect 1435 2158 1439 2162
rect 1443 2158 1495 2162
rect 1499 2158 1535 2162
rect 1539 2158 1567 2162
rect 1571 2158 1631 2162
rect 1635 2158 1639 2162
rect 1643 2158 1711 2162
rect 1715 2158 1727 2162
rect 1731 2158 1783 2162
rect 1787 2158 1815 2162
rect 1819 2158 1855 2162
rect 1859 2158 1895 2162
rect 1899 2158 1935 2162
rect 1939 2158 1975 2162
rect 1979 2158 2015 2162
rect 2019 2158 2047 2162
rect 2051 2158 2095 2162
rect 2099 2158 2111 2162
rect 2115 2158 2175 2162
rect 2179 2158 2183 2162
rect 2187 2158 2239 2162
rect 2243 2158 2279 2162
rect 2283 2158 2311 2162
rect 2315 2158 2359 2162
rect 2363 2158 2407 2162
rect 2411 2158 2447 2162
rect 1269 2157 2447 2158
rect 2453 2157 2454 2163
rect 84 2137 85 2143
rect 91 2142 1251 2143
rect 91 2138 111 2142
rect 115 2138 247 2142
rect 251 2138 287 2142
rect 291 2138 327 2142
rect 331 2138 375 2142
rect 379 2138 383 2142
rect 387 2138 423 2142
rect 427 2138 431 2142
rect 435 2138 463 2142
rect 467 2138 495 2142
rect 499 2138 503 2142
rect 507 2138 551 2142
rect 555 2138 607 2142
rect 611 2138 663 2142
rect 667 2138 719 2142
rect 723 2138 727 2142
rect 731 2138 783 2142
rect 787 2138 791 2142
rect 795 2138 847 2142
rect 851 2138 855 2142
rect 859 2138 911 2142
rect 915 2138 967 2142
rect 971 2138 1023 2142
rect 1027 2138 1079 2142
rect 1083 2138 1143 2142
rect 1147 2138 1239 2142
rect 1243 2138 1251 2142
rect 91 2137 1251 2138
rect 1257 2137 1258 2143
rect 1250 2085 1251 2091
rect 1257 2090 2435 2091
rect 1257 2086 1279 2090
rect 1283 2086 1303 2090
rect 1307 2086 1343 2090
rect 1347 2086 1351 2090
rect 1355 2086 1399 2090
rect 1403 2086 1439 2090
rect 1443 2086 1479 2090
rect 1483 2086 1535 2090
rect 1539 2086 1567 2090
rect 1571 2086 1631 2090
rect 1635 2086 1663 2090
rect 1667 2086 1727 2090
rect 1731 2086 1759 2090
rect 1763 2086 1815 2090
rect 1819 2086 1847 2090
rect 1851 2086 1895 2090
rect 1899 2086 1935 2090
rect 1939 2086 1975 2090
rect 1979 2086 2015 2090
rect 2019 2086 2047 2090
rect 2051 2086 2095 2090
rect 2099 2086 2111 2090
rect 2115 2086 2167 2090
rect 2171 2086 2175 2090
rect 2179 2086 2239 2090
rect 2243 2086 2311 2090
rect 2315 2086 2359 2090
rect 2363 2086 2407 2090
rect 2411 2086 2435 2090
rect 1257 2085 2435 2086
rect 2441 2085 2442 2091
rect 96 2069 97 2075
rect 103 2074 1263 2075
rect 103 2070 111 2074
rect 115 2070 383 2074
rect 387 2070 423 2074
rect 427 2070 463 2074
rect 467 2070 503 2074
rect 507 2070 543 2074
rect 547 2070 551 2074
rect 555 2070 583 2074
rect 587 2070 607 2074
rect 611 2070 631 2074
rect 635 2070 663 2074
rect 667 2070 687 2074
rect 691 2070 727 2074
rect 731 2070 743 2074
rect 747 2070 791 2074
rect 795 2070 799 2074
rect 803 2070 847 2074
rect 851 2070 855 2074
rect 859 2070 903 2074
rect 907 2070 911 2074
rect 915 2070 959 2074
rect 963 2070 967 2074
rect 971 2070 1015 2074
rect 1019 2070 1023 2074
rect 1027 2070 1071 2074
rect 1075 2070 1079 2074
rect 1083 2070 1143 2074
rect 1147 2070 1239 2074
rect 1243 2070 1263 2074
rect 103 2069 1263 2070
rect 1269 2069 1270 2075
rect 1262 2009 1263 2015
rect 1269 2014 2447 2015
rect 1269 2010 1279 2014
rect 1283 2010 1303 2014
rect 1307 2010 1343 2014
rect 1347 2010 1351 2014
rect 1355 2010 1399 2014
rect 1403 2010 1423 2014
rect 1427 2010 1479 2014
rect 1483 2010 1495 2014
rect 1499 2010 1567 2014
rect 1571 2010 1575 2014
rect 1579 2010 1663 2014
rect 1667 2010 1751 2014
rect 1755 2010 1759 2014
rect 1763 2010 1839 2014
rect 1843 2010 1847 2014
rect 1851 2010 1919 2014
rect 1923 2010 1935 2014
rect 1939 2010 1999 2014
rect 2003 2010 2015 2014
rect 2019 2010 2071 2014
rect 2075 2010 2095 2014
rect 2099 2010 2135 2014
rect 2139 2010 2167 2014
rect 2171 2010 2191 2014
rect 2195 2010 2239 2014
rect 2243 2010 2255 2014
rect 2259 2010 2311 2014
rect 2315 2010 2319 2014
rect 2323 2010 2359 2014
rect 2363 2010 2407 2014
rect 2411 2010 2447 2014
rect 1269 2009 2447 2010
rect 2453 2009 2454 2015
rect 84 1993 85 1999
rect 91 1998 1251 1999
rect 91 1994 111 1998
rect 115 1994 367 1998
rect 371 1994 383 1998
rect 387 1994 407 1998
rect 411 1994 423 1998
rect 427 1994 455 1998
rect 459 1994 463 1998
rect 467 1994 503 1998
rect 507 1994 511 1998
rect 515 1994 543 1998
rect 547 1994 567 1998
rect 571 1994 583 1998
rect 587 1994 631 1998
rect 635 1994 687 1998
rect 691 1994 695 1998
rect 699 1994 743 1998
rect 747 1994 759 1998
rect 763 1994 799 1998
rect 803 1994 815 1998
rect 819 1994 847 1998
rect 851 1994 871 1998
rect 875 1994 903 1998
rect 907 1994 935 1998
rect 939 1994 959 1998
rect 963 1994 999 1998
rect 1003 1994 1015 1998
rect 1019 1994 1063 1998
rect 1067 1994 1071 1998
rect 1075 1994 1239 1998
rect 1243 1994 1251 1998
rect 91 1993 1251 1994
rect 1257 1993 1258 1999
rect 1250 1941 1251 1947
rect 1257 1946 2435 1947
rect 1257 1942 1279 1946
rect 1283 1942 1303 1946
rect 1307 1942 1351 1946
rect 1355 1942 1359 1946
rect 1363 1942 1423 1946
rect 1427 1942 1447 1946
rect 1451 1942 1495 1946
rect 1499 1942 1535 1946
rect 1539 1942 1575 1946
rect 1579 1942 1623 1946
rect 1627 1942 1663 1946
rect 1667 1942 1711 1946
rect 1715 1942 1751 1946
rect 1755 1942 1791 1946
rect 1795 1942 1839 1946
rect 1843 1942 1863 1946
rect 1867 1942 1919 1946
rect 1923 1942 1935 1946
rect 1939 1942 1999 1946
rect 2003 1942 2007 1946
rect 2011 1942 2071 1946
rect 2075 1942 2079 1946
rect 2083 1942 2135 1946
rect 2139 1942 2151 1946
rect 2155 1942 2191 1946
rect 2195 1942 2223 1946
rect 2227 1942 2255 1946
rect 2259 1942 2303 1946
rect 2307 1942 2319 1946
rect 2323 1942 2359 1946
rect 2363 1942 2407 1946
rect 2411 1942 2435 1946
rect 1257 1941 2435 1942
rect 2441 1941 2442 1947
rect 96 1921 97 1927
rect 103 1926 1263 1927
rect 103 1922 111 1926
rect 115 1922 175 1926
rect 179 1922 215 1926
rect 219 1922 263 1926
rect 267 1922 319 1926
rect 323 1922 367 1926
rect 371 1922 391 1926
rect 395 1922 407 1926
rect 411 1922 455 1926
rect 459 1922 471 1926
rect 475 1922 511 1926
rect 515 1922 551 1926
rect 555 1922 567 1926
rect 571 1922 631 1926
rect 635 1922 639 1926
rect 643 1922 695 1926
rect 699 1922 719 1926
rect 723 1922 759 1926
rect 763 1922 799 1926
rect 803 1922 815 1926
rect 819 1922 871 1926
rect 875 1922 879 1926
rect 883 1922 935 1926
rect 939 1922 959 1926
rect 963 1922 999 1926
rect 1003 1922 1039 1926
rect 1043 1922 1063 1926
rect 1067 1922 1119 1926
rect 1123 1922 1239 1926
rect 1243 1922 1263 1926
rect 103 1921 1263 1922
rect 1269 1921 1270 1927
rect 1262 1873 1263 1879
rect 1269 1878 2447 1879
rect 1269 1874 1279 1878
rect 1283 1874 1303 1878
rect 1307 1874 1311 1878
rect 1315 1874 1359 1878
rect 1363 1874 1415 1878
rect 1419 1874 1447 1878
rect 1451 1874 1479 1878
rect 1483 1874 1535 1878
rect 1539 1874 1543 1878
rect 1547 1874 1615 1878
rect 1619 1874 1623 1878
rect 1627 1874 1687 1878
rect 1691 1874 1711 1878
rect 1715 1874 1767 1878
rect 1771 1874 1791 1878
rect 1795 1874 1863 1878
rect 1867 1874 1935 1878
rect 1939 1874 1975 1878
rect 1979 1874 2007 1878
rect 2011 1874 2079 1878
rect 2083 1874 2095 1878
rect 2099 1874 2151 1878
rect 2155 1874 2223 1878
rect 2227 1874 2303 1878
rect 2307 1874 2359 1878
rect 2363 1874 2407 1878
rect 2411 1874 2447 1878
rect 1269 1873 2447 1874
rect 2453 1873 2454 1879
rect 84 1845 85 1851
rect 91 1850 1251 1851
rect 91 1846 111 1850
rect 115 1846 135 1850
rect 139 1846 175 1850
rect 179 1846 215 1850
rect 219 1846 263 1850
rect 267 1846 271 1850
rect 275 1846 319 1850
rect 323 1846 351 1850
rect 355 1846 391 1850
rect 395 1846 439 1850
rect 443 1846 471 1850
rect 475 1846 535 1850
rect 539 1846 551 1850
rect 555 1846 631 1850
rect 635 1846 639 1850
rect 643 1846 719 1850
rect 723 1846 727 1850
rect 731 1846 799 1850
rect 803 1846 823 1850
rect 827 1846 879 1850
rect 883 1846 911 1850
rect 915 1846 959 1850
rect 963 1846 991 1850
rect 995 1846 1039 1850
rect 1043 1846 1063 1850
rect 1067 1846 1119 1850
rect 1123 1846 1135 1850
rect 1139 1846 1191 1850
rect 1195 1846 1239 1850
rect 1243 1846 1251 1850
rect 91 1845 1251 1846
rect 1257 1845 1258 1851
rect 1250 1801 1251 1807
rect 1257 1806 2435 1807
rect 1257 1802 1279 1806
rect 1283 1802 1311 1806
rect 1315 1802 1359 1806
rect 1363 1802 1407 1806
rect 1411 1802 1415 1806
rect 1419 1802 1471 1806
rect 1475 1802 1479 1806
rect 1483 1802 1535 1806
rect 1539 1802 1543 1806
rect 1547 1802 1599 1806
rect 1603 1802 1615 1806
rect 1619 1802 1663 1806
rect 1667 1802 1687 1806
rect 1691 1802 1727 1806
rect 1731 1802 1767 1806
rect 1771 1802 1783 1806
rect 1787 1802 1839 1806
rect 1843 1802 1863 1806
rect 1867 1802 1895 1806
rect 1899 1802 1959 1806
rect 1963 1802 1975 1806
rect 1979 1802 2095 1806
rect 2099 1802 2223 1806
rect 2227 1802 2359 1806
rect 2363 1802 2407 1806
rect 2411 1802 2435 1806
rect 1257 1801 2435 1802
rect 2441 1801 2442 1807
rect 96 1777 97 1783
rect 103 1782 1263 1783
rect 103 1778 111 1782
rect 115 1778 135 1782
rect 139 1778 175 1782
rect 179 1778 215 1782
rect 219 1778 271 1782
rect 275 1778 287 1782
rect 291 1778 351 1782
rect 355 1778 375 1782
rect 379 1778 439 1782
rect 443 1778 471 1782
rect 475 1778 535 1782
rect 539 1778 567 1782
rect 571 1778 631 1782
rect 635 1778 663 1782
rect 667 1778 727 1782
rect 731 1778 751 1782
rect 755 1778 823 1782
rect 827 1778 831 1782
rect 835 1778 903 1782
rect 907 1778 911 1782
rect 915 1778 967 1782
rect 971 1778 991 1782
rect 995 1778 1031 1782
rect 1035 1778 1063 1782
rect 1067 1778 1087 1782
rect 1091 1778 1135 1782
rect 1139 1778 1151 1782
rect 1155 1778 1191 1782
rect 1195 1778 1239 1782
rect 1243 1778 1263 1782
rect 103 1777 1263 1778
rect 1269 1777 1270 1783
rect 1262 1733 1263 1739
rect 1269 1738 2447 1739
rect 1269 1734 1279 1738
rect 1283 1734 1303 1738
rect 1307 1734 1351 1738
rect 1355 1734 1407 1738
rect 1411 1734 1423 1738
rect 1427 1734 1471 1738
rect 1475 1734 1503 1738
rect 1507 1734 1535 1738
rect 1539 1734 1583 1738
rect 1587 1734 1599 1738
rect 1603 1734 1663 1738
rect 1667 1734 1727 1738
rect 1731 1734 1735 1738
rect 1739 1734 1783 1738
rect 1787 1734 1807 1738
rect 1811 1734 1839 1738
rect 1843 1734 1871 1738
rect 1875 1734 1895 1738
rect 1899 1734 1935 1738
rect 1939 1734 1959 1738
rect 1963 1734 1999 1738
rect 2003 1734 2063 1738
rect 2067 1734 2407 1738
rect 2411 1734 2447 1738
rect 1269 1733 2447 1734
rect 2453 1733 2454 1739
rect 84 1705 85 1711
rect 91 1710 1251 1711
rect 91 1706 111 1710
rect 115 1706 135 1710
rect 139 1706 175 1710
rect 179 1706 215 1710
rect 219 1706 239 1710
rect 243 1706 287 1710
rect 291 1706 319 1710
rect 323 1706 375 1710
rect 379 1706 415 1710
rect 419 1706 471 1710
rect 475 1706 511 1710
rect 515 1706 567 1710
rect 571 1706 615 1710
rect 619 1706 663 1710
rect 667 1706 711 1710
rect 715 1706 751 1710
rect 755 1706 799 1710
rect 803 1706 831 1710
rect 835 1706 879 1710
rect 883 1706 903 1710
rect 907 1706 951 1710
rect 955 1706 967 1710
rect 971 1706 1015 1710
rect 1019 1706 1031 1710
rect 1035 1706 1087 1710
rect 1091 1706 1151 1710
rect 1155 1706 1159 1710
rect 1163 1706 1191 1710
rect 1195 1706 1239 1710
rect 1243 1706 1251 1710
rect 91 1705 1251 1706
rect 1257 1705 1258 1711
rect 1250 1665 1251 1671
rect 1257 1670 2435 1671
rect 1257 1666 1279 1670
rect 1283 1666 1303 1670
rect 1307 1666 1351 1670
rect 1355 1666 1359 1670
rect 1363 1666 1423 1670
rect 1427 1666 1447 1670
rect 1451 1666 1503 1670
rect 1507 1666 1543 1670
rect 1547 1666 1583 1670
rect 1587 1666 1639 1670
rect 1643 1666 1663 1670
rect 1667 1666 1727 1670
rect 1731 1666 1735 1670
rect 1739 1666 1807 1670
rect 1811 1666 1815 1670
rect 1819 1666 1871 1670
rect 1875 1666 1895 1670
rect 1899 1666 1935 1670
rect 1939 1666 1967 1670
rect 1971 1666 1999 1670
rect 2003 1666 2031 1670
rect 2035 1666 2063 1670
rect 2067 1666 2095 1670
rect 2099 1666 2159 1670
rect 2163 1666 2223 1670
rect 2227 1666 2407 1670
rect 2411 1666 2435 1670
rect 1257 1665 2435 1666
rect 2441 1665 2442 1671
rect 278 1660 284 1661
rect 622 1660 628 1661
rect 278 1656 279 1660
rect 283 1656 623 1660
rect 627 1656 628 1660
rect 278 1655 284 1656
rect 622 1655 628 1656
rect 96 1633 97 1639
rect 103 1638 1263 1639
rect 103 1634 111 1638
rect 115 1634 135 1638
rect 139 1634 175 1638
rect 179 1634 239 1638
rect 243 1634 271 1638
rect 275 1634 311 1638
rect 315 1634 319 1638
rect 323 1634 359 1638
rect 363 1634 415 1638
rect 419 1634 471 1638
rect 475 1634 511 1638
rect 515 1634 535 1638
rect 539 1634 599 1638
rect 603 1634 615 1638
rect 619 1634 663 1638
rect 667 1634 711 1638
rect 715 1634 719 1638
rect 723 1634 775 1638
rect 779 1634 799 1638
rect 803 1634 831 1638
rect 835 1634 879 1638
rect 883 1634 887 1638
rect 891 1634 943 1638
rect 947 1634 951 1638
rect 955 1634 999 1638
rect 1003 1634 1015 1638
rect 1019 1634 1087 1638
rect 1091 1634 1159 1638
rect 1163 1634 1239 1638
rect 1243 1634 1263 1638
rect 103 1633 1263 1634
rect 1269 1633 1270 1639
rect 1262 1597 1263 1603
rect 1269 1602 2447 1603
rect 1269 1598 1279 1602
rect 1283 1598 1303 1602
rect 1307 1598 1327 1602
rect 1331 1598 1359 1602
rect 1363 1598 1399 1602
rect 1403 1598 1447 1602
rect 1451 1598 1479 1602
rect 1483 1598 1543 1602
rect 1547 1598 1567 1602
rect 1571 1598 1639 1602
rect 1643 1598 1655 1602
rect 1659 1598 1727 1602
rect 1731 1598 1743 1602
rect 1747 1598 1815 1602
rect 1819 1598 1831 1602
rect 1835 1598 1895 1602
rect 1899 1598 1911 1602
rect 1915 1598 1967 1602
rect 1971 1598 1983 1602
rect 1987 1598 2031 1602
rect 2035 1598 2047 1602
rect 2051 1598 2095 1602
rect 2099 1598 2111 1602
rect 2115 1598 2159 1602
rect 2163 1598 2167 1602
rect 2171 1598 2215 1602
rect 2219 1598 2223 1602
rect 2227 1598 2271 1602
rect 2275 1598 2319 1602
rect 2323 1598 2359 1602
rect 2363 1598 2407 1602
rect 2411 1598 2447 1602
rect 1269 1597 2447 1598
rect 2453 1597 2454 1603
rect 84 1557 85 1563
rect 91 1562 1251 1563
rect 91 1558 111 1562
rect 115 1558 271 1562
rect 275 1558 311 1562
rect 315 1558 327 1562
rect 331 1558 359 1562
rect 363 1558 367 1562
rect 371 1558 407 1562
rect 411 1558 415 1562
rect 419 1558 447 1562
rect 451 1558 471 1562
rect 475 1558 487 1562
rect 491 1558 527 1562
rect 531 1558 535 1562
rect 539 1558 567 1562
rect 571 1558 599 1562
rect 603 1558 607 1562
rect 611 1558 647 1562
rect 651 1558 663 1562
rect 667 1558 687 1562
rect 691 1558 719 1562
rect 723 1558 727 1562
rect 731 1558 767 1562
rect 771 1558 775 1562
rect 779 1558 807 1562
rect 811 1558 831 1562
rect 835 1558 847 1562
rect 851 1558 887 1562
rect 891 1558 927 1562
rect 931 1558 943 1562
rect 947 1558 999 1562
rect 1003 1558 1239 1562
rect 1243 1558 1251 1562
rect 91 1557 1251 1558
rect 1257 1557 1258 1563
rect 1250 1525 1251 1531
rect 1257 1530 2435 1531
rect 1257 1526 1279 1530
rect 1283 1526 1327 1530
rect 1331 1526 1335 1530
rect 1339 1526 1399 1530
rect 1403 1526 1415 1530
rect 1419 1526 1479 1530
rect 1483 1526 1503 1530
rect 1507 1526 1567 1530
rect 1571 1526 1615 1530
rect 1619 1526 1655 1530
rect 1659 1526 1743 1530
rect 1747 1526 1831 1530
rect 1835 1526 1887 1530
rect 1891 1526 1911 1530
rect 1915 1526 1983 1530
rect 1987 1526 2047 1530
rect 2051 1526 2111 1530
rect 2115 1526 2167 1530
rect 2171 1526 2215 1530
rect 2219 1526 2271 1530
rect 2275 1526 2319 1530
rect 2323 1526 2359 1530
rect 2363 1526 2407 1530
rect 2411 1526 2435 1530
rect 1257 1525 2435 1526
rect 2441 1525 2442 1531
rect 1262 1457 1263 1463
rect 1269 1462 2447 1463
rect 1269 1458 1279 1462
rect 1283 1458 1335 1462
rect 1339 1458 1375 1462
rect 1379 1458 1415 1462
rect 1419 1458 1463 1462
rect 1467 1458 1503 1462
rect 1507 1458 1551 1462
rect 1555 1458 1615 1462
rect 1619 1458 1639 1462
rect 1643 1458 1727 1462
rect 1731 1458 1743 1462
rect 1747 1458 1807 1462
rect 1811 1458 1879 1462
rect 1883 1458 1887 1462
rect 1891 1458 1943 1462
rect 1947 1458 1999 1462
rect 2003 1458 2047 1462
rect 2051 1458 2095 1462
rect 2099 1458 2143 1462
rect 2147 1458 2191 1462
rect 2195 1458 2215 1462
rect 2219 1458 2239 1462
rect 2243 1458 2279 1462
rect 2283 1458 2319 1462
rect 2323 1458 2359 1462
rect 2363 1458 2407 1462
rect 2411 1458 2447 1462
rect 1269 1457 2447 1458
rect 2453 1457 2454 1463
rect 1262 1455 1270 1457
rect 96 1449 97 1455
rect 103 1454 1263 1455
rect 103 1450 111 1454
rect 115 1450 143 1454
rect 147 1450 183 1454
rect 187 1450 223 1454
rect 227 1450 263 1454
rect 267 1450 319 1454
rect 323 1450 327 1454
rect 331 1450 367 1454
rect 371 1450 391 1454
rect 395 1450 407 1454
rect 411 1450 447 1454
rect 451 1450 471 1454
rect 475 1450 487 1454
rect 491 1450 527 1454
rect 531 1450 559 1454
rect 563 1450 567 1454
rect 571 1450 607 1454
rect 611 1450 647 1454
rect 651 1450 687 1454
rect 691 1450 727 1454
rect 731 1450 767 1454
rect 771 1450 807 1454
rect 811 1450 847 1454
rect 851 1450 879 1454
rect 883 1450 887 1454
rect 891 1450 927 1454
rect 931 1450 943 1454
rect 947 1450 999 1454
rect 1003 1450 1047 1454
rect 1051 1450 1103 1454
rect 1107 1450 1151 1454
rect 1155 1450 1191 1454
rect 1195 1450 1239 1454
rect 1243 1450 1263 1454
rect 103 1449 1263 1450
rect 1269 1449 1270 1455
rect 84 1381 85 1387
rect 91 1386 1251 1387
rect 91 1382 111 1386
rect 115 1382 143 1386
rect 147 1382 167 1386
rect 171 1382 183 1386
rect 187 1382 207 1386
rect 211 1382 223 1386
rect 227 1382 247 1386
rect 251 1382 263 1386
rect 267 1382 303 1386
rect 307 1382 319 1386
rect 323 1382 367 1386
rect 371 1382 391 1386
rect 395 1382 439 1386
rect 443 1382 471 1386
rect 475 1382 519 1386
rect 523 1382 559 1386
rect 563 1382 599 1386
rect 603 1382 647 1386
rect 651 1382 679 1386
rect 683 1382 727 1386
rect 731 1382 751 1386
rect 755 1382 807 1386
rect 811 1382 823 1386
rect 827 1382 879 1386
rect 883 1382 887 1386
rect 891 1382 943 1386
rect 947 1382 951 1386
rect 955 1382 999 1386
rect 1003 1382 1015 1386
rect 1019 1382 1047 1386
rect 1051 1382 1079 1386
rect 1083 1382 1103 1386
rect 1107 1382 1143 1386
rect 1147 1382 1151 1386
rect 1155 1382 1191 1386
rect 1195 1382 1239 1386
rect 1243 1382 1251 1386
rect 91 1381 1251 1382
rect 1257 1386 2442 1387
rect 1257 1382 1279 1386
rect 1283 1382 1303 1386
rect 1307 1382 1343 1386
rect 1347 1382 1375 1386
rect 1379 1382 1399 1386
rect 1403 1382 1463 1386
rect 1467 1382 1535 1386
rect 1539 1382 1551 1386
rect 1555 1382 1607 1386
rect 1611 1382 1639 1386
rect 1643 1382 1687 1386
rect 1691 1382 1727 1386
rect 1731 1382 1767 1386
rect 1771 1382 1807 1386
rect 1811 1382 1847 1386
rect 1851 1382 1879 1386
rect 1883 1382 1935 1386
rect 1939 1382 1943 1386
rect 1947 1382 1999 1386
rect 2003 1382 2023 1386
rect 2027 1382 2047 1386
rect 2051 1382 2095 1386
rect 2099 1382 2111 1386
rect 2115 1382 2143 1386
rect 2147 1382 2191 1386
rect 2195 1382 2199 1386
rect 2203 1382 2239 1386
rect 2243 1382 2279 1386
rect 2283 1382 2287 1386
rect 2291 1382 2319 1386
rect 2323 1382 2359 1386
rect 2363 1382 2407 1386
rect 2411 1382 2442 1386
rect 1257 1381 2442 1382
rect 278 1324 284 1325
rect 606 1324 612 1325
rect 278 1320 279 1324
rect 283 1320 607 1324
rect 611 1320 612 1324
rect 278 1319 284 1320
rect 606 1319 612 1320
rect 1262 1318 2454 1319
rect 1262 1315 1279 1318
rect 96 1309 97 1315
rect 103 1314 1263 1315
rect 103 1310 111 1314
rect 115 1310 167 1314
rect 171 1310 183 1314
rect 187 1310 207 1314
rect 211 1310 231 1314
rect 235 1310 247 1314
rect 251 1310 287 1314
rect 291 1310 303 1314
rect 307 1310 351 1314
rect 355 1310 367 1314
rect 371 1310 423 1314
rect 427 1310 439 1314
rect 443 1310 495 1314
rect 499 1310 519 1314
rect 523 1310 567 1314
rect 571 1310 599 1314
rect 603 1310 639 1314
rect 643 1310 679 1314
rect 683 1310 703 1314
rect 707 1310 751 1314
rect 755 1310 767 1314
rect 771 1310 823 1314
rect 827 1310 879 1314
rect 883 1310 887 1314
rect 891 1310 935 1314
rect 939 1310 951 1314
rect 955 1310 999 1314
rect 1003 1310 1015 1314
rect 1019 1310 1079 1314
rect 1083 1310 1143 1314
rect 1147 1310 1191 1314
rect 1195 1310 1239 1314
rect 1243 1310 1263 1314
rect 103 1309 1263 1310
rect 1269 1314 1279 1315
rect 1283 1314 1303 1318
rect 1307 1314 1343 1318
rect 1347 1314 1383 1318
rect 1387 1314 1399 1318
rect 1403 1314 1423 1318
rect 1427 1314 1463 1318
rect 1467 1314 1503 1318
rect 1507 1314 1535 1318
rect 1539 1314 1543 1318
rect 1547 1314 1583 1318
rect 1587 1314 1607 1318
rect 1611 1314 1623 1318
rect 1627 1314 1679 1318
rect 1683 1314 1687 1318
rect 1691 1314 1735 1318
rect 1739 1314 1767 1318
rect 1771 1314 1791 1318
rect 1795 1314 1847 1318
rect 1851 1314 1903 1318
rect 1907 1314 1935 1318
rect 1939 1314 1967 1318
rect 1971 1314 2023 1318
rect 2027 1314 2039 1318
rect 2043 1314 2111 1318
rect 2115 1314 2119 1318
rect 2123 1314 2199 1318
rect 2203 1314 2287 1318
rect 2291 1314 2359 1318
rect 2363 1314 2407 1318
rect 2411 1314 2454 1318
rect 1269 1313 2454 1314
rect 1269 1309 1270 1313
rect 84 1237 85 1243
rect 91 1242 1251 1243
rect 91 1238 111 1242
rect 115 1238 135 1242
rect 139 1238 175 1242
rect 179 1238 183 1242
rect 187 1238 231 1242
rect 235 1238 287 1242
rect 291 1238 311 1242
rect 315 1238 351 1242
rect 355 1238 399 1242
rect 403 1238 423 1242
rect 427 1238 487 1242
rect 491 1238 495 1242
rect 499 1238 567 1242
rect 571 1238 575 1242
rect 579 1238 639 1242
rect 643 1238 663 1242
rect 667 1238 703 1242
rect 707 1238 743 1242
rect 747 1238 767 1242
rect 771 1238 815 1242
rect 819 1238 823 1242
rect 827 1238 879 1242
rect 883 1238 935 1242
rect 939 1238 943 1242
rect 947 1238 999 1242
rect 1003 1238 1007 1242
rect 1011 1238 1071 1242
rect 1075 1238 1239 1242
rect 1243 1238 1251 1242
rect 91 1237 1251 1238
rect 1257 1242 2442 1243
rect 1257 1238 1279 1242
rect 1283 1238 1303 1242
rect 1307 1238 1343 1242
rect 1347 1238 1375 1242
rect 1379 1238 1383 1242
rect 1387 1238 1423 1242
rect 1427 1238 1463 1242
rect 1467 1238 1479 1242
rect 1483 1238 1503 1242
rect 1507 1238 1543 1242
rect 1547 1238 1583 1242
rect 1587 1238 1623 1242
rect 1627 1238 1679 1242
rect 1683 1238 1687 1242
rect 1691 1238 1735 1242
rect 1739 1238 1791 1242
rect 1795 1238 1847 1242
rect 1851 1238 1887 1242
rect 1891 1238 1903 1242
rect 1907 1238 1967 1242
rect 1971 1238 1983 1242
rect 1987 1238 2039 1242
rect 2043 1238 2071 1242
rect 2075 1238 2119 1242
rect 2123 1238 2151 1242
rect 2155 1238 2199 1242
rect 2203 1238 2223 1242
rect 2227 1238 2287 1242
rect 2291 1238 2303 1242
rect 2307 1238 2359 1242
rect 2363 1238 2407 1242
rect 2411 1238 2442 1242
rect 1257 1237 2442 1238
rect 96 1169 97 1175
rect 103 1174 1263 1175
rect 103 1170 111 1174
rect 115 1170 135 1174
rect 139 1170 175 1174
rect 179 1170 231 1174
rect 235 1170 239 1174
rect 243 1170 311 1174
rect 315 1170 327 1174
rect 331 1170 399 1174
rect 403 1170 431 1174
rect 435 1170 487 1174
rect 491 1170 535 1174
rect 539 1170 575 1174
rect 579 1170 639 1174
rect 643 1170 663 1174
rect 667 1170 743 1174
rect 747 1170 815 1174
rect 819 1170 839 1174
rect 843 1170 879 1174
rect 883 1170 919 1174
rect 923 1170 943 1174
rect 947 1170 999 1174
rect 1003 1170 1007 1174
rect 1011 1170 1071 1174
rect 1075 1170 1143 1174
rect 1147 1170 1191 1174
rect 1195 1170 1239 1174
rect 1243 1170 1263 1174
rect 103 1169 1263 1170
rect 1269 1174 2454 1175
rect 1269 1170 1279 1174
rect 1283 1170 1303 1174
rect 1307 1170 1343 1174
rect 1347 1170 1375 1174
rect 1379 1170 1407 1174
rect 1411 1170 1479 1174
rect 1483 1170 1487 1174
rect 1491 1170 1583 1174
rect 1587 1170 1687 1174
rect 1691 1170 1791 1174
rect 1795 1170 1799 1174
rect 1803 1170 1887 1174
rect 1891 1170 1903 1174
rect 1907 1170 1983 1174
rect 1987 1170 1999 1174
rect 2003 1170 2071 1174
rect 2075 1170 2079 1174
rect 2083 1170 2151 1174
rect 2155 1170 2159 1174
rect 2163 1170 2223 1174
rect 2227 1170 2231 1174
rect 2235 1170 2303 1174
rect 2307 1170 2359 1174
rect 2363 1170 2407 1174
rect 2411 1170 2454 1174
rect 1269 1169 2454 1170
rect 1250 1106 2442 1107
rect 1250 1103 1279 1106
rect 84 1097 85 1103
rect 91 1102 1251 1103
rect 91 1098 111 1102
rect 115 1098 135 1102
rect 139 1098 175 1102
rect 179 1098 239 1102
rect 243 1098 247 1102
rect 251 1098 327 1102
rect 331 1098 415 1102
rect 419 1098 431 1102
rect 435 1098 503 1102
rect 507 1098 535 1102
rect 539 1098 583 1102
rect 587 1098 639 1102
rect 643 1098 663 1102
rect 667 1098 735 1102
rect 739 1098 743 1102
rect 747 1098 799 1102
rect 803 1098 839 1102
rect 843 1098 863 1102
rect 867 1098 919 1102
rect 923 1098 983 1102
rect 987 1098 999 1102
rect 1003 1098 1047 1102
rect 1051 1098 1071 1102
rect 1075 1098 1143 1102
rect 1147 1098 1191 1102
rect 1195 1098 1239 1102
rect 1243 1098 1251 1102
rect 91 1097 1251 1098
rect 1257 1102 1279 1103
rect 1283 1102 1303 1106
rect 1307 1102 1343 1106
rect 1347 1102 1407 1106
rect 1411 1102 1431 1106
rect 1435 1102 1471 1106
rect 1475 1102 1487 1106
rect 1491 1102 1511 1106
rect 1515 1102 1559 1106
rect 1563 1102 1583 1106
rect 1587 1102 1615 1106
rect 1619 1102 1671 1106
rect 1675 1102 1687 1106
rect 1691 1102 1727 1106
rect 1731 1102 1775 1106
rect 1779 1102 1799 1106
rect 1803 1102 1823 1106
rect 1827 1102 1871 1106
rect 1875 1102 1903 1106
rect 1907 1102 1919 1106
rect 1923 1102 1967 1106
rect 1971 1102 1999 1106
rect 2003 1102 2015 1106
rect 2019 1102 2063 1106
rect 2067 1102 2079 1106
rect 2083 1102 2119 1106
rect 2123 1102 2159 1106
rect 2163 1102 2175 1106
rect 2179 1102 2231 1106
rect 2235 1102 2303 1106
rect 2307 1102 2359 1106
rect 2363 1102 2407 1106
rect 2411 1102 2442 1106
rect 1257 1101 2442 1102
rect 1257 1097 1258 1101
rect 762 1084 768 1085
rect 1070 1084 1076 1085
rect 762 1080 763 1084
rect 767 1080 1071 1084
rect 1075 1080 1076 1084
rect 762 1079 768 1080
rect 1070 1079 1076 1080
rect 1438 1068 1444 1069
rect 1734 1068 1740 1069
rect 1438 1064 1439 1068
rect 1443 1064 1735 1068
rect 1739 1064 1740 1068
rect 1438 1063 1444 1064
rect 1734 1063 1740 1064
rect 1262 1038 2454 1039
rect 1262 1035 1279 1038
rect 96 1029 97 1035
rect 103 1034 1263 1035
rect 103 1030 111 1034
rect 115 1030 135 1034
rect 139 1030 175 1034
rect 179 1030 247 1034
rect 251 1030 255 1034
rect 259 1030 327 1034
rect 331 1030 399 1034
rect 403 1030 415 1034
rect 419 1030 463 1034
rect 467 1030 503 1034
rect 507 1030 519 1034
rect 523 1030 575 1034
rect 579 1030 583 1034
rect 587 1030 623 1034
rect 627 1030 663 1034
rect 667 1030 671 1034
rect 675 1030 735 1034
rect 739 1030 799 1034
rect 803 1030 807 1034
rect 811 1030 863 1034
rect 867 1030 895 1034
rect 899 1030 919 1034
rect 923 1030 983 1034
rect 987 1030 999 1034
rect 1003 1030 1047 1034
rect 1051 1030 1103 1034
rect 1107 1030 1191 1034
rect 1195 1030 1239 1034
rect 1243 1030 1263 1034
rect 103 1029 1263 1030
rect 1269 1034 1279 1035
rect 1283 1034 1431 1038
rect 1435 1034 1471 1038
rect 1475 1034 1511 1038
rect 1515 1034 1559 1038
rect 1563 1034 1575 1038
rect 1579 1034 1615 1038
rect 1619 1034 1655 1038
rect 1659 1034 1671 1038
rect 1675 1034 1695 1038
rect 1699 1034 1727 1038
rect 1731 1034 1735 1038
rect 1739 1034 1775 1038
rect 1779 1034 1823 1038
rect 1827 1034 1871 1038
rect 1875 1034 1879 1038
rect 1883 1034 1919 1038
rect 1923 1034 1943 1038
rect 1947 1034 1967 1038
rect 1971 1034 2015 1038
rect 2019 1034 2063 1038
rect 2067 1034 2095 1038
rect 2099 1034 2119 1038
rect 2123 1034 2175 1038
rect 2179 1034 2231 1038
rect 2235 1034 2255 1038
rect 2259 1034 2407 1038
rect 2411 1034 2454 1038
rect 1269 1033 2454 1034
rect 1269 1029 1270 1033
rect 718 996 724 997
rect 1126 996 1132 997
rect 718 992 719 996
rect 723 992 1127 996
rect 1131 992 1132 996
rect 718 991 724 992
rect 1126 991 1132 992
rect 84 961 85 967
rect 91 966 1251 967
rect 91 962 111 966
rect 115 962 175 966
rect 179 962 215 966
rect 219 962 255 966
rect 259 962 303 966
rect 307 962 327 966
rect 331 962 359 966
rect 363 962 399 966
rect 403 962 415 966
rect 419 962 463 966
rect 467 962 519 966
rect 523 962 575 966
rect 579 962 623 966
rect 627 962 639 966
rect 643 962 671 966
rect 675 962 711 966
rect 715 962 735 966
rect 739 962 783 966
rect 787 962 807 966
rect 811 962 855 966
rect 859 962 895 966
rect 899 962 927 966
rect 931 962 999 966
rect 1003 962 1071 966
rect 1075 962 1103 966
rect 1107 962 1143 966
rect 1147 962 1191 966
rect 1195 962 1239 966
rect 1243 962 1251 966
rect 91 961 1251 962
rect 1257 963 1258 967
rect 1257 962 2442 963
rect 1257 961 1279 962
rect 1250 958 1279 961
rect 1283 958 1303 962
rect 1307 958 1351 962
rect 1355 958 1431 962
rect 1435 958 1511 962
rect 1515 958 1575 962
rect 1579 958 1591 962
rect 1595 958 1615 962
rect 1619 958 1655 962
rect 1659 958 1679 962
rect 1683 958 1695 962
rect 1699 958 1735 962
rect 1739 958 1767 962
rect 1771 958 1775 962
rect 1779 958 1823 962
rect 1827 958 1855 962
rect 1859 958 1879 962
rect 1883 958 1943 962
rect 1947 958 2015 962
rect 2019 958 2023 962
rect 2027 958 2095 962
rect 2099 958 2103 962
rect 2107 958 2175 962
rect 2179 958 2183 962
rect 2187 958 2255 962
rect 2259 958 2271 962
rect 2275 958 2407 962
rect 2411 958 2442 962
rect 1250 957 2442 958
rect 1262 894 2454 895
rect 1262 891 1279 894
rect 96 885 97 891
rect 103 890 1263 891
rect 103 886 111 890
rect 115 886 191 890
rect 195 886 215 890
rect 219 886 231 890
rect 235 886 255 890
rect 259 886 287 890
rect 291 886 303 890
rect 307 886 359 890
rect 363 886 415 890
rect 419 886 447 890
rect 451 886 463 890
rect 467 886 519 890
rect 523 886 543 890
rect 547 886 575 890
rect 579 886 639 890
rect 643 886 711 890
rect 715 886 727 890
rect 731 886 783 890
rect 787 886 807 890
rect 811 886 855 890
rect 859 886 887 890
rect 891 886 927 890
rect 931 886 959 890
rect 963 886 999 890
rect 1003 886 1023 890
rect 1027 886 1071 890
rect 1075 886 1087 890
rect 1091 886 1143 890
rect 1147 886 1159 890
rect 1163 886 1191 890
rect 1195 886 1239 890
rect 1243 886 1263 890
rect 103 885 1263 886
rect 1269 890 1279 891
rect 1283 890 1303 894
rect 1307 890 1351 894
rect 1355 890 1431 894
rect 1435 890 1439 894
rect 1443 890 1479 894
rect 1483 890 1511 894
rect 1515 890 1519 894
rect 1523 890 1559 894
rect 1563 890 1591 894
rect 1595 890 1607 894
rect 1611 890 1655 894
rect 1659 890 1679 894
rect 1683 890 1711 894
rect 1715 890 1767 894
rect 1771 890 1775 894
rect 1779 890 1847 894
rect 1851 890 1855 894
rect 1859 890 1919 894
rect 1923 890 1943 894
rect 1947 890 1991 894
rect 1995 890 2023 894
rect 2027 890 2063 894
rect 2067 890 2103 894
rect 2107 890 2135 894
rect 2139 890 2183 894
rect 2187 890 2215 894
rect 2219 890 2271 894
rect 2275 890 2295 894
rect 2299 890 2407 894
rect 2411 890 2454 894
rect 1269 889 2454 890
rect 1269 885 1270 889
rect 84 817 85 823
rect 91 822 1251 823
rect 91 818 111 822
rect 115 818 135 822
rect 139 818 175 822
rect 179 818 191 822
rect 195 818 231 822
rect 235 818 239 822
rect 243 818 287 822
rect 291 818 327 822
rect 331 818 359 822
rect 363 818 415 822
rect 419 818 447 822
rect 451 818 503 822
rect 507 818 543 822
rect 547 818 591 822
rect 595 818 639 822
rect 643 818 671 822
rect 675 818 727 822
rect 731 818 743 822
rect 747 818 807 822
rect 811 818 815 822
rect 819 818 879 822
rect 883 818 887 822
rect 891 818 943 822
rect 947 818 959 822
rect 963 818 1015 822
rect 1019 818 1023 822
rect 1027 818 1087 822
rect 1091 818 1159 822
rect 1163 818 1239 822
rect 1243 818 1251 822
rect 91 817 1251 818
rect 1257 817 1258 823
rect 1250 815 1258 817
rect 1250 809 1251 815
rect 1257 814 2435 815
rect 1257 810 1279 814
rect 1283 810 1359 814
rect 1363 810 1415 814
rect 1419 810 1439 814
rect 1443 810 1471 814
rect 1475 810 1479 814
rect 1483 810 1519 814
rect 1523 810 1535 814
rect 1539 810 1559 814
rect 1563 810 1591 814
rect 1595 810 1607 814
rect 1611 810 1647 814
rect 1651 810 1655 814
rect 1659 810 1703 814
rect 1707 810 1711 814
rect 1715 810 1759 814
rect 1763 810 1775 814
rect 1779 810 1815 814
rect 1819 810 1847 814
rect 1851 810 1871 814
rect 1875 810 1919 814
rect 1923 810 1935 814
rect 1939 810 1991 814
rect 1995 810 1999 814
rect 2003 810 2063 814
rect 2067 810 2071 814
rect 2075 810 2135 814
rect 2139 810 2143 814
rect 2147 810 2215 814
rect 2219 810 2223 814
rect 2227 810 2295 814
rect 2299 810 2303 814
rect 2307 810 2359 814
rect 2363 810 2407 814
rect 2411 810 2435 814
rect 1257 809 2435 810
rect 2441 809 2442 815
rect 1838 764 1844 765
rect 2150 764 2156 765
rect 1838 760 1839 764
rect 1843 760 2151 764
rect 2155 760 2156 764
rect 1838 759 1844 760
rect 2150 759 2156 760
rect 96 745 97 751
rect 103 750 1263 751
rect 103 746 111 750
rect 115 746 135 750
rect 139 746 175 750
rect 179 746 191 750
rect 195 746 239 750
rect 243 746 263 750
rect 267 746 327 750
rect 331 746 335 750
rect 339 746 399 750
rect 403 746 415 750
rect 419 746 455 750
rect 459 746 503 750
rect 507 746 543 750
rect 547 746 583 750
rect 587 746 591 750
rect 595 746 623 750
rect 627 746 671 750
rect 675 746 719 750
rect 723 746 743 750
rect 747 746 767 750
rect 771 746 815 750
rect 819 746 863 750
rect 867 746 879 750
rect 883 746 911 750
rect 915 746 943 750
rect 947 746 1015 750
rect 1019 746 1239 750
rect 1243 746 1263 750
rect 103 745 1263 746
rect 1269 747 1270 751
rect 1269 746 2454 747
rect 1269 745 1279 746
rect 1262 742 1279 745
rect 1283 742 1303 746
rect 1307 742 1343 746
rect 1347 742 1359 746
rect 1363 742 1407 746
rect 1411 742 1415 746
rect 1419 742 1471 746
rect 1475 742 1487 746
rect 1491 742 1535 746
rect 1539 742 1575 746
rect 1579 742 1591 746
rect 1595 742 1647 746
rect 1651 742 1663 746
rect 1667 742 1703 746
rect 1707 742 1751 746
rect 1755 742 1759 746
rect 1763 742 1815 746
rect 1819 742 1831 746
rect 1835 742 1871 746
rect 1875 742 1911 746
rect 1915 742 1935 746
rect 1939 742 1991 746
rect 1995 742 1999 746
rect 2003 742 2071 746
rect 2075 742 2079 746
rect 2083 742 2143 746
rect 2147 742 2175 746
rect 2179 742 2223 746
rect 2227 742 2279 746
rect 2283 742 2303 746
rect 2307 742 2359 746
rect 2363 742 2407 746
rect 2411 742 2454 746
rect 1262 741 2454 742
rect 84 673 85 679
rect 91 678 1251 679
rect 91 674 111 678
rect 115 674 135 678
rect 139 674 191 678
rect 195 674 199 678
rect 203 674 263 678
rect 267 674 279 678
rect 283 674 335 678
rect 339 674 351 678
rect 355 674 399 678
rect 403 674 415 678
rect 419 674 455 678
rect 459 674 487 678
rect 491 674 503 678
rect 507 674 543 678
rect 547 674 559 678
rect 563 674 583 678
rect 587 674 623 678
rect 627 674 639 678
rect 643 674 671 678
rect 675 674 711 678
rect 715 674 719 678
rect 723 674 767 678
rect 771 674 783 678
rect 787 674 815 678
rect 819 674 855 678
rect 859 674 863 678
rect 867 674 911 678
rect 915 674 919 678
rect 923 674 983 678
rect 987 674 1039 678
rect 1043 674 1095 678
rect 1099 674 1151 678
rect 1155 674 1191 678
rect 1195 674 1239 678
rect 1243 674 1251 678
rect 91 673 1251 674
rect 1257 675 1258 679
rect 1257 674 2442 675
rect 1257 673 1279 674
rect 1250 670 1279 673
rect 1283 670 1303 674
rect 1307 670 1343 674
rect 1347 670 1399 674
rect 1403 670 1407 674
rect 1411 670 1487 674
rect 1491 670 1511 674
rect 1515 670 1575 674
rect 1579 670 1623 674
rect 1627 670 1663 674
rect 1667 670 1727 674
rect 1731 670 1751 674
rect 1755 670 1815 674
rect 1819 670 1831 674
rect 1835 670 1895 674
rect 1899 670 1911 674
rect 1915 670 1975 674
rect 1979 670 1991 674
rect 1995 670 2047 674
rect 2051 670 2079 674
rect 2083 670 2111 674
rect 2115 670 2175 674
rect 2179 670 2239 674
rect 2243 670 2279 674
rect 2283 670 2311 674
rect 2315 670 2359 674
rect 2363 670 2407 674
rect 2411 670 2442 674
rect 1250 669 2442 670
rect 96 597 97 603
rect 103 602 1263 603
rect 103 598 111 602
rect 115 598 135 602
rect 139 598 191 602
rect 195 598 199 602
rect 203 598 271 602
rect 275 598 279 602
rect 283 598 351 602
rect 355 598 359 602
rect 363 598 415 602
rect 419 598 447 602
rect 451 598 487 602
rect 491 598 535 602
rect 539 598 559 602
rect 563 598 623 602
rect 627 598 639 602
rect 643 598 703 602
rect 707 598 711 602
rect 715 598 783 602
rect 787 598 855 602
rect 859 598 919 602
rect 923 598 975 602
rect 979 598 983 602
rect 987 598 1023 602
rect 1027 598 1039 602
rect 1043 598 1079 602
rect 1083 598 1095 602
rect 1099 598 1135 602
rect 1139 598 1151 602
rect 1155 598 1191 602
rect 1195 598 1239 602
rect 1243 598 1263 602
rect 103 597 1263 598
rect 1269 602 2454 603
rect 1269 598 1279 602
rect 1283 598 1303 602
rect 1307 598 1399 602
rect 1403 598 1415 602
rect 1419 598 1455 602
rect 1459 598 1495 602
rect 1499 598 1511 602
rect 1515 598 1543 602
rect 1547 598 1599 602
rect 1603 598 1623 602
rect 1627 598 1663 602
rect 1667 598 1727 602
rect 1731 598 1791 602
rect 1795 598 1815 602
rect 1819 598 1847 602
rect 1851 598 1895 602
rect 1899 598 1911 602
rect 1915 598 1975 602
rect 1979 598 2047 602
rect 2051 598 2111 602
rect 2115 598 2119 602
rect 2123 598 2175 602
rect 2179 598 2199 602
rect 2203 598 2239 602
rect 2243 598 2287 602
rect 2291 598 2311 602
rect 2315 598 2359 602
rect 2363 598 2407 602
rect 2411 598 2454 602
rect 1269 597 2454 598
rect 902 564 908 565
rect 1214 564 1220 565
rect 902 560 903 564
rect 907 560 1215 564
rect 1219 560 1220 564
rect 902 559 908 560
rect 1214 559 1220 560
rect 1250 529 1251 535
rect 1257 534 2435 535
rect 1257 530 1279 534
rect 1283 530 1303 534
rect 1307 530 1375 534
rect 1379 530 1415 534
rect 1419 530 1455 534
rect 1459 530 1479 534
rect 1483 530 1495 534
rect 1499 530 1543 534
rect 1547 530 1583 534
rect 1587 530 1599 534
rect 1603 530 1663 534
rect 1667 530 1695 534
rect 1699 530 1727 534
rect 1731 530 1791 534
rect 1795 530 1799 534
rect 1803 530 1847 534
rect 1851 530 1903 534
rect 1907 530 1911 534
rect 1915 530 1975 534
rect 1979 530 2007 534
rect 2011 530 2047 534
rect 2051 530 2103 534
rect 2107 530 2119 534
rect 2123 530 2191 534
rect 2195 530 2199 534
rect 2203 530 2287 534
rect 2291 530 2359 534
rect 2363 530 2407 534
rect 2411 530 2435 534
rect 1257 529 2435 530
rect 2441 529 2442 535
rect 1250 527 1258 529
rect 84 521 85 527
rect 91 526 1251 527
rect 91 522 111 526
rect 115 522 135 526
rect 139 522 191 526
rect 195 522 263 526
rect 267 522 271 526
rect 275 522 335 526
rect 339 522 359 526
rect 363 522 415 526
rect 419 522 447 526
rect 451 522 495 526
rect 499 522 535 526
rect 539 522 575 526
rect 579 522 623 526
rect 627 522 647 526
rect 651 522 703 526
rect 707 522 719 526
rect 723 522 783 526
rect 787 522 847 526
rect 851 522 855 526
rect 859 522 903 526
rect 907 522 919 526
rect 923 522 959 526
rect 963 522 975 526
rect 979 522 1023 526
rect 1027 522 1079 526
rect 1083 522 1087 526
rect 1091 522 1135 526
rect 1139 522 1151 526
rect 1155 522 1191 526
rect 1195 522 1239 526
rect 1243 522 1251 526
rect 91 521 1251 522
rect 1257 521 1258 527
rect 1262 462 2454 463
rect 1262 459 1279 462
rect 96 453 97 459
rect 103 458 1263 459
rect 103 454 111 458
rect 115 454 135 458
rect 139 454 183 458
rect 187 454 191 458
rect 195 454 223 458
rect 227 454 263 458
rect 267 454 311 458
rect 315 454 335 458
rect 339 454 367 458
rect 371 454 415 458
rect 419 454 431 458
rect 435 454 495 458
rect 499 454 559 458
rect 563 454 575 458
rect 579 454 615 458
rect 619 454 647 458
rect 651 454 671 458
rect 675 454 719 458
rect 723 454 775 458
rect 779 454 783 458
rect 787 454 831 458
rect 835 454 847 458
rect 851 454 887 458
rect 891 454 903 458
rect 907 454 959 458
rect 963 454 1023 458
rect 1027 454 1087 458
rect 1091 454 1151 458
rect 1155 454 1191 458
rect 1195 454 1239 458
rect 1243 454 1263 458
rect 103 453 1263 454
rect 1269 458 1279 459
rect 1283 458 1303 462
rect 1307 458 1343 462
rect 1347 458 1375 462
rect 1379 458 1399 462
rect 1403 458 1463 462
rect 1467 458 1479 462
rect 1483 458 1527 462
rect 1531 458 1583 462
rect 1587 458 1591 462
rect 1595 458 1663 462
rect 1667 458 1695 462
rect 1699 458 1735 462
rect 1739 458 1799 462
rect 1803 458 1815 462
rect 1819 458 1895 462
rect 1899 458 1903 462
rect 1907 458 1975 462
rect 1979 458 2007 462
rect 2011 458 2055 462
rect 2059 458 2103 462
rect 2107 458 2135 462
rect 2139 458 2191 462
rect 2195 458 2215 462
rect 2219 458 2287 462
rect 2291 458 2295 462
rect 2299 458 2359 462
rect 2363 458 2407 462
rect 2411 458 2454 462
rect 1269 457 2454 458
rect 1269 453 1270 457
rect 84 385 85 391
rect 91 390 1251 391
rect 91 386 111 390
rect 115 386 135 390
rect 139 386 175 390
rect 179 386 183 390
rect 187 386 223 390
rect 227 386 231 390
rect 235 386 263 390
rect 267 386 287 390
rect 291 386 311 390
rect 315 386 343 390
rect 347 386 367 390
rect 371 386 391 390
rect 395 386 431 390
rect 435 386 439 390
rect 443 386 487 390
rect 491 386 495 390
rect 499 386 535 390
rect 539 386 559 390
rect 563 386 583 390
rect 587 386 615 390
rect 619 386 631 390
rect 635 386 671 390
rect 675 386 679 390
rect 683 386 719 390
rect 723 386 727 390
rect 731 386 775 390
rect 779 386 831 390
rect 835 386 887 390
rect 891 386 1239 390
rect 1243 386 1251 390
rect 91 385 1251 386
rect 1257 390 2442 391
rect 1257 386 1279 390
rect 1283 386 1303 390
rect 1307 386 1343 390
rect 1347 386 1399 390
rect 1403 386 1447 390
rect 1451 386 1463 390
rect 1467 386 1487 390
rect 1491 386 1527 390
rect 1531 386 1535 390
rect 1539 386 1591 390
rect 1595 386 1663 390
rect 1667 386 1735 390
rect 1739 386 1815 390
rect 1819 386 1895 390
rect 1899 386 1967 390
rect 1971 386 1975 390
rect 1979 386 2039 390
rect 2043 386 2055 390
rect 2059 386 2111 390
rect 2115 386 2135 390
rect 2139 386 2175 390
rect 2179 386 2215 390
rect 2219 386 2239 390
rect 2243 386 2295 390
rect 2299 386 2303 390
rect 2307 386 2359 390
rect 2363 386 2407 390
rect 2411 386 2442 390
rect 1257 385 2442 386
rect 96 313 97 319
rect 103 318 1263 319
rect 103 314 111 318
rect 115 314 135 318
rect 139 314 175 318
rect 179 314 183 318
rect 187 314 231 318
rect 235 314 255 318
rect 259 314 287 318
rect 291 314 327 318
rect 331 314 343 318
rect 347 314 391 318
rect 395 314 439 318
rect 443 314 447 318
rect 451 314 487 318
rect 491 314 503 318
rect 507 314 535 318
rect 539 314 551 318
rect 555 314 583 318
rect 587 314 591 318
rect 595 314 631 318
rect 635 314 679 318
rect 683 314 727 318
rect 731 314 775 318
rect 779 314 823 318
rect 827 314 871 318
rect 875 314 919 318
rect 923 314 1239 318
rect 1243 314 1263 318
rect 103 313 1263 314
rect 1269 318 2454 319
rect 1269 314 1279 318
rect 1283 314 1447 318
rect 1451 314 1487 318
rect 1491 314 1495 318
rect 1499 314 1535 318
rect 1539 314 1575 318
rect 1579 314 1591 318
rect 1595 314 1615 318
rect 1619 314 1655 318
rect 1659 314 1663 318
rect 1667 314 1695 318
rect 1699 314 1735 318
rect 1739 314 1743 318
rect 1747 314 1799 318
rect 1803 314 1815 318
rect 1819 314 1863 318
rect 1867 314 1895 318
rect 1899 314 1935 318
rect 1939 314 1967 318
rect 1971 314 2007 318
rect 2011 314 2039 318
rect 2043 314 2071 318
rect 2075 314 2111 318
rect 2115 314 2135 318
rect 2139 314 2175 318
rect 2179 314 2191 318
rect 2195 314 2239 318
rect 2243 314 2255 318
rect 2259 314 2303 318
rect 2307 314 2319 318
rect 2323 314 2359 318
rect 2363 314 2407 318
rect 2411 314 2454 318
rect 1269 313 2454 314
rect 1250 246 2442 247
rect 1250 243 1279 246
rect 84 237 85 243
rect 91 242 1251 243
rect 91 238 111 242
rect 115 238 135 242
rect 139 238 175 242
rect 179 238 183 242
rect 187 238 247 242
rect 251 238 255 242
rect 259 238 327 242
rect 331 238 391 242
rect 395 238 415 242
rect 419 238 447 242
rect 451 238 495 242
rect 499 238 503 242
rect 507 238 551 242
rect 555 238 575 242
rect 579 238 591 242
rect 595 238 631 242
rect 635 238 655 242
rect 659 238 679 242
rect 683 238 727 242
rect 731 238 775 242
rect 779 238 791 242
rect 795 238 823 242
rect 827 238 847 242
rect 851 238 871 242
rect 875 238 903 242
rect 907 238 919 242
rect 923 238 959 242
rect 963 238 1023 242
rect 1027 238 1239 242
rect 1243 238 1251 242
rect 91 237 1251 238
rect 1257 242 1279 243
rect 1283 242 1367 246
rect 1371 242 1407 246
rect 1411 242 1447 246
rect 1451 242 1495 246
rect 1499 242 1535 246
rect 1539 242 1551 246
rect 1555 242 1575 246
rect 1579 242 1607 246
rect 1611 242 1615 246
rect 1619 242 1655 246
rect 1659 242 1671 246
rect 1675 242 1695 246
rect 1699 242 1735 246
rect 1739 242 1743 246
rect 1747 242 1799 246
rect 1803 242 1807 246
rect 1811 242 1863 246
rect 1867 242 1887 246
rect 1891 242 1935 246
rect 1939 242 1975 246
rect 1979 242 2007 246
rect 2011 242 2071 246
rect 2075 242 2135 246
rect 2139 242 2167 246
rect 2171 242 2191 246
rect 2195 242 2255 246
rect 2259 242 2271 246
rect 2275 242 2319 246
rect 2323 242 2359 246
rect 2363 242 2407 246
rect 2411 242 2442 246
rect 1257 241 2442 242
rect 1257 237 1258 241
rect 1742 188 1748 189
rect 1982 188 1988 189
rect 1742 184 1743 188
rect 1747 184 1983 188
rect 1987 184 1988 188
rect 1742 183 1748 184
rect 1982 183 1988 184
rect 1262 157 1263 163
rect 1269 162 2447 163
rect 1269 158 1279 162
rect 1283 158 1303 162
rect 1307 158 1343 162
rect 1347 158 1367 162
rect 1371 158 1383 162
rect 1387 158 1407 162
rect 1411 158 1423 162
rect 1427 158 1447 162
rect 1451 158 1463 162
rect 1467 158 1495 162
rect 1499 158 1519 162
rect 1523 158 1551 162
rect 1555 158 1583 162
rect 1587 158 1607 162
rect 1611 158 1647 162
rect 1651 158 1671 162
rect 1675 158 1711 162
rect 1715 158 1735 162
rect 1739 158 1767 162
rect 1771 158 1807 162
rect 1811 158 1823 162
rect 1827 158 1871 162
rect 1875 158 1887 162
rect 1891 158 1919 162
rect 1923 158 1967 162
rect 1971 158 1975 162
rect 1979 158 2015 162
rect 2019 158 2063 162
rect 2067 158 2071 162
rect 2075 158 2111 162
rect 2115 158 2159 162
rect 2163 158 2167 162
rect 2171 158 2215 162
rect 2219 158 2271 162
rect 2275 158 2319 162
rect 2323 158 2359 162
rect 2363 158 2407 162
rect 2411 158 2447 162
rect 1269 157 2447 158
rect 2453 157 2454 163
rect 1262 155 1270 157
rect 96 149 97 155
rect 103 154 1263 155
rect 103 150 111 154
rect 115 150 135 154
rect 139 150 175 154
rect 179 150 215 154
rect 219 150 247 154
rect 251 150 255 154
rect 259 150 295 154
rect 299 150 327 154
rect 331 150 335 154
rect 339 150 375 154
rect 379 150 415 154
rect 419 150 423 154
rect 427 150 471 154
rect 475 150 495 154
rect 499 150 527 154
rect 531 150 575 154
rect 579 150 583 154
rect 587 150 631 154
rect 635 150 655 154
rect 659 150 679 154
rect 683 150 727 154
rect 731 150 767 154
rect 771 150 791 154
rect 795 150 807 154
rect 811 150 847 154
rect 851 150 887 154
rect 891 150 903 154
rect 907 150 927 154
rect 931 150 959 154
rect 963 150 975 154
rect 979 150 1023 154
rect 1027 150 1071 154
rect 1075 150 1111 154
rect 1115 150 1151 154
rect 1155 150 1191 154
rect 1195 150 1239 154
rect 1243 150 1263 154
rect 103 149 1263 150
rect 1269 149 1270 155
rect 1250 89 1251 95
rect 1257 94 2435 95
rect 1257 90 1279 94
rect 1283 90 1303 94
rect 1307 90 1343 94
rect 1347 90 1383 94
rect 1387 90 1423 94
rect 1427 90 1463 94
rect 1467 90 1519 94
rect 1523 90 1583 94
rect 1587 90 1647 94
rect 1651 90 1711 94
rect 1715 90 1767 94
rect 1771 90 1823 94
rect 1827 90 1871 94
rect 1875 90 1919 94
rect 1923 90 1967 94
rect 1971 90 2015 94
rect 2019 90 2063 94
rect 2067 90 2111 94
rect 2115 90 2159 94
rect 2163 90 2215 94
rect 2219 90 2271 94
rect 2275 90 2319 94
rect 2323 90 2359 94
rect 2363 90 2407 94
rect 2411 90 2435 94
rect 1257 89 2435 90
rect 2441 89 2442 95
rect 1250 87 1258 89
rect 84 81 85 87
rect 91 86 1251 87
rect 91 82 111 86
rect 115 82 135 86
rect 139 82 175 86
rect 179 82 215 86
rect 219 82 255 86
rect 259 82 295 86
rect 299 82 335 86
rect 339 82 375 86
rect 379 82 423 86
rect 427 82 471 86
rect 475 82 527 86
rect 531 82 583 86
rect 587 82 631 86
rect 635 82 679 86
rect 683 82 727 86
rect 731 82 767 86
rect 771 82 807 86
rect 811 82 847 86
rect 851 82 887 86
rect 891 82 927 86
rect 931 82 975 86
rect 979 82 1023 86
rect 1027 82 1071 86
rect 1075 82 1111 86
rect 1115 82 1151 86
rect 1155 82 1191 86
rect 1195 82 1239 86
rect 1243 82 1251 86
rect 91 81 1251 82
rect 1257 81 1258 87
<< m5c >>
rect 1251 2509 1257 2515
rect 2435 2509 2441 2515
rect 97 2497 103 2503
rect 1263 2497 1269 2503
rect 1263 2441 1269 2447
rect 2447 2441 2453 2447
rect 85 2429 91 2435
rect 1251 2429 1257 2435
rect 1251 2373 1257 2379
rect 2435 2373 2441 2379
rect 97 2353 103 2359
rect 1263 2353 1269 2359
rect 1263 2301 1269 2307
rect 2447 2301 2453 2307
rect 85 2281 91 2287
rect 1251 2281 1257 2287
rect 1251 2225 1257 2231
rect 2435 2225 2441 2231
rect 97 2213 103 2219
rect 1263 2213 1269 2219
rect 1263 2157 1269 2163
rect 2447 2157 2453 2163
rect 85 2137 91 2143
rect 1251 2137 1257 2143
rect 1251 2085 1257 2091
rect 2435 2085 2441 2091
rect 97 2069 103 2075
rect 1263 2069 1269 2075
rect 1263 2009 1269 2015
rect 2447 2009 2453 2015
rect 85 1993 91 1999
rect 1251 1993 1257 1999
rect 1251 1941 1257 1947
rect 2435 1941 2441 1947
rect 97 1921 103 1927
rect 1263 1921 1269 1927
rect 1263 1873 1269 1879
rect 2447 1873 2453 1879
rect 85 1845 91 1851
rect 1251 1845 1257 1851
rect 1251 1801 1257 1807
rect 2435 1801 2441 1807
rect 97 1777 103 1783
rect 1263 1777 1269 1783
rect 1263 1733 1269 1739
rect 2447 1733 2453 1739
rect 85 1705 91 1711
rect 1251 1705 1257 1711
rect 1251 1665 1257 1671
rect 2435 1665 2441 1671
rect 97 1633 103 1639
rect 1263 1633 1269 1639
rect 1263 1597 1269 1603
rect 2447 1597 2453 1603
rect 85 1557 91 1563
rect 1251 1557 1257 1563
rect 1251 1525 1257 1531
rect 2435 1525 2441 1531
rect 1263 1457 1269 1463
rect 2447 1457 2453 1463
rect 97 1449 103 1455
rect 1263 1449 1269 1455
rect 85 1381 91 1387
rect 1251 1381 1257 1387
rect 97 1309 103 1315
rect 1263 1309 1269 1315
rect 85 1237 91 1243
rect 1251 1237 1257 1243
rect 97 1169 103 1175
rect 1263 1169 1269 1175
rect 85 1097 91 1103
rect 1251 1097 1257 1103
rect 97 1029 103 1035
rect 1263 1029 1269 1035
rect 85 961 91 967
rect 1251 961 1257 967
rect 97 885 103 891
rect 1263 885 1269 891
rect 85 817 91 823
rect 1251 817 1257 823
rect 1251 809 1257 815
rect 2435 809 2441 815
rect 97 745 103 751
rect 1263 745 1269 751
rect 85 673 91 679
rect 1251 673 1257 679
rect 97 597 103 603
rect 1263 597 1269 603
rect 1251 529 1257 535
rect 2435 529 2441 535
rect 85 521 91 527
rect 1251 521 1257 527
rect 97 453 103 459
rect 1263 453 1269 459
rect 85 385 91 391
rect 1251 385 1257 391
rect 97 313 103 319
rect 1263 313 1269 319
rect 85 237 91 243
rect 1251 237 1257 243
rect 1263 157 1269 163
rect 2447 157 2453 163
rect 97 149 103 155
rect 1263 149 1269 155
rect 1251 89 1257 95
rect 2435 89 2441 95
rect 85 81 91 87
rect 1251 81 1257 87
<< m5 >>
rect 84 2435 92 2520
rect 84 2429 85 2435
rect 91 2429 92 2435
rect 84 2287 92 2429
rect 84 2281 85 2287
rect 91 2281 92 2287
rect 84 2143 92 2281
rect 84 2137 85 2143
rect 91 2137 92 2143
rect 84 1999 92 2137
rect 84 1993 85 1999
rect 91 1993 92 1999
rect 84 1851 92 1993
rect 84 1845 85 1851
rect 91 1845 92 1851
rect 84 1711 92 1845
rect 84 1705 85 1711
rect 91 1705 92 1711
rect 84 1563 92 1705
rect 84 1557 85 1563
rect 91 1557 92 1563
rect 84 1387 92 1557
rect 84 1381 85 1387
rect 91 1381 92 1387
rect 84 1243 92 1381
rect 84 1237 85 1243
rect 91 1237 92 1243
rect 84 1103 92 1237
rect 84 1097 85 1103
rect 91 1097 92 1103
rect 84 967 92 1097
rect 84 961 85 967
rect 91 961 92 967
rect 84 823 92 961
rect 84 817 85 823
rect 91 817 92 823
rect 84 679 92 817
rect 84 673 85 679
rect 91 673 92 679
rect 84 527 92 673
rect 84 521 85 527
rect 91 521 92 527
rect 84 391 92 521
rect 84 385 85 391
rect 91 385 92 391
rect 84 243 92 385
rect 84 237 85 243
rect 91 237 92 243
rect 84 87 92 237
rect 84 81 85 87
rect 91 81 92 87
rect 84 72 92 81
rect 96 2503 104 2520
rect 96 2497 97 2503
rect 103 2497 104 2503
rect 96 2359 104 2497
rect 96 2353 97 2359
rect 103 2353 104 2359
rect 96 2219 104 2353
rect 96 2213 97 2219
rect 103 2213 104 2219
rect 96 2075 104 2213
rect 96 2069 97 2075
rect 103 2069 104 2075
rect 96 1927 104 2069
rect 96 1921 97 1927
rect 103 1921 104 1927
rect 96 1783 104 1921
rect 96 1777 97 1783
rect 103 1777 104 1783
rect 96 1639 104 1777
rect 96 1633 97 1639
rect 103 1633 104 1639
rect 96 1455 104 1633
rect 96 1449 97 1455
rect 103 1449 104 1455
rect 96 1315 104 1449
rect 96 1309 97 1315
rect 103 1309 104 1315
rect 96 1175 104 1309
rect 96 1169 97 1175
rect 103 1169 104 1175
rect 96 1035 104 1169
rect 96 1029 97 1035
rect 103 1029 104 1035
rect 96 891 104 1029
rect 96 885 97 891
rect 103 885 104 891
rect 96 751 104 885
rect 96 745 97 751
rect 103 745 104 751
rect 96 603 104 745
rect 96 597 97 603
rect 103 597 104 603
rect 96 459 104 597
rect 96 453 97 459
rect 103 453 104 459
rect 96 319 104 453
rect 96 313 97 319
rect 103 313 104 319
rect 96 155 104 313
rect 96 149 97 155
rect 103 149 104 155
rect 96 72 104 149
rect 1250 2515 1258 2520
rect 1250 2509 1251 2515
rect 1257 2509 1258 2515
rect 1250 2435 1258 2509
rect 1250 2429 1251 2435
rect 1257 2429 1258 2435
rect 1250 2379 1258 2429
rect 1250 2373 1251 2379
rect 1257 2373 1258 2379
rect 1250 2287 1258 2373
rect 1250 2281 1251 2287
rect 1257 2281 1258 2287
rect 1250 2231 1258 2281
rect 1250 2225 1251 2231
rect 1257 2225 1258 2231
rect 1250 2143 1258 2225
rect 1250 2137 1251 2143
rect 1257 2137 1258 2143
rect 1250 2091 1258 2137
rect 1250 2085 1251 2091
rect 1257 2085 1258 2091
rect 1250 1999 1258 2085
rect 1250 1993 1251 1999
rect 1257 1993 1258 1999
rect 1250 1947 1258 1993
rect 1250 1941 1251 1947
rect 1257 1941 1258 1947
rect 1250 1851 1258 1941
rect 1250 1845 1251 1851
rect 1257 1845 1258 1851
rect 1250 1807 1258 1845
rect 1250 1801 1251 1807
rect 1257 1801 1258 1807
rect 1250 1711 1258 1801
rect 1250 1705 1251 1711
rect 1257 1705 1258 1711
rect 1250 1671 1258 1705
rect 1250 1665 1251 1671
rect 1257 1665 1258 1671
rect 1250 1563 1258 1665
rect 1250 1557 1251 1563
rect 1257 1557 1258 1563
rect 1250 1531 1258 1557
rect 1250 1525 1251 1531
rect 1257 1525 1258 1531
rect 1250 1387 1258 1525
rect 1250 1381 1251 1387
rect 1257 1381 1258 1387
rect 1250 1243 1258 1381
rect 1250 1237 1251 1243
rect 1257 1237 1258 1243
rect 1250 1103 1258 1237
rect 1250 1097 1251 1103
rect 1257 1097 1258 1103
rect 1250 967 1258 1097
rect 1250 961 1251 967
rect 1257 961 1258 967
rect 1250 823 1258 961
rect 1250 817 1251 823
rect 1257 817 1258 823
rect 1250 815 1258 817
rect 1250 809 1251 815
rect 1257 809 1258 815
rect 1250 679 1258 809
rect 1250 673 1251 679
rect 1257 673 1258 679
rect 1250 535 1258 673
rect 1250 529 1251 535
rect 1257 529 1258 535
rect 1250 527 1258 529
rect 1250 521 1251 527
rect 1257 521 1258 527
rect 1250 391 1258 521
rect 1250 385 1251 391
rect 1257 385 1258 391
rect 1250 243 1258 385
rect 1250 237 1251 243
rect 1257 237 1258 243
rect 1250 95 1258 237
rect 1250 89 1251 95
rect 1257 89 1258 95
rect 1250 87 1258 89
rect 1250 81 1251 87
rect 1257 81 1258 87
rect 1250 72 1258 81
rect 1262 2503 1270 2520
rect 1262 2497 1263 2503
rect 1269 2497 1270 2503
rect 1262 2447 1270 2497
rect 1262 2441 1263 2447
rect 1269 2441 1270 2447
rect 1262 2359 1270 2441
rect 1262 2353 1263 2359
rect 1269 2353 1270 2359
rect 1262 2307 1270 2353
rect 1262 2301 1263 2307
rect 1269 2301 1270 2307
rect 1262 2219 1270 2301
rect 1262 2213 1263 2219
rect 1269 2213 1270 2219
rect 1262 2163 1270 2213
rect 1262 2157 1263 2163
rect 1269 2157 1270 2163
rect 1262 2075 1270 2157
rect 1262 2069 1263 2075
rect 1269 2069 1270 2075
rect 1262 2015 1270 2069
rect 1262 2009 1263 2015
rect 1269 2009 1270 2015
rect 1262 1927 1270 2009
rect 1262 1921 1263 1927
rect 1269 1921 1270 1927
rect 1262 1879 1270 1921
rect 1262 1873 1263 1879
rect 1269 1873 1270 1879
rect 1262 1783 1270 1873
rect 1262 1777 1263 1783
rect 1269 1777 1270 1783
rect 1262 1739 1270 1777
rect 1262 1733 1263 1739
rect 1269 1733 1270 1739
rect 1262 1639 1270 1733
rect 1262 1633 1263 1639
rect 1269 1633 1270 1639
rect 1262 1603 1270 1633
rect 1262 1597 1263 1603
rect 1269 1597 1270 1603
rect 1262 1463 1270 1597
rect 1262 1457 1263 1463
rect 1269 1457 1270 1463
rect 1262 1455 1270 1457
rect 1262 1449 1263 1455
rect 1269 1449 1270 1455
rect 1262 1315 1270 1449
rect 1262 1309 1263 1315
rect 1269 1309 1270 1315
rect 1262 1175 1270 1309
rect 1262 1169 1263 1175
rect 1269 1169 1270 1175
rect 1262 1035 1270 1169
rect 1262 1029 1263 1035
rect 1269 1029 1270 1035
rect 1262 891 1270 1029
rect 1262 885 1263 891
rect 1269 885 1270 891
rect 1262 751 1270 885
rect 1262 745 1263 751
rect 1269 745 1270 751
rect 1262 603 1270 745
rect 1262 597 1263 603
rect 1269 597 1270 603
rect 1262 459 1270 597
rect 1262 453 1263 459
rect 1269 453 1270 459
rect 1262 319 1270 453
rect 1262 313 1263 319
rect 1269 313 1270 319
rect 1262 163 1270 313
rect 1262 157 1263 163
rect 1269 157 1270 163
rect 1262 155 1270 157
rect 1262 149 1263 155
rect 1269 149 1270 155
rect 1262 72 1270 149
rect 2434 2515 2442 2520
rect 2434 2509 2435 2515
rect 2441 2509 2442 2515
rect 2434 2379 2442 2509
rect 2434 2373 2435 2379
rect 2441 2373 2442 2379
rect 2434 2231 2442 2373
rect 2434 2225 2435 2231
rect 2441 2225 2442 2231
rect 2434 2091 2442 2225
rect 2434 2085 2435 2091
rect 2441 2085 2442 2091
rect 2434 1947 2442 2085
rect 2434 1941 2435 1947
rect 2441 1941 2442 1947
rect 2434 1807 2442 1941
rect 2434 1801 2435 1807
rect 2441 1801 2442 1807
rect 2434 1671 2442 1801
rect 2434 1665 2435 1671
rect 2441 1665 2442 1671
rect 2434 1531 2442 1665
rect 2434 1525 2435 1531
rect 2441 1525 2442 1531
rect 2434 815 2442 1525
rect 2434 809 2435 815
rect 2441 809 2442 815
rect 2434 535 2442 809
rect 2434 529 2435 535
rect 2441 529 2442 535
rect 2434 95 2442 529
rect 2434 89 2435 95
rect 2441 89 2442 95
rect 2434 72 2442 89
rect 2446 2447 2454 2520
rect 2446 2441 2447 2447
rect 2453 2441 2454 2447
rect 2446 2307 2454 2441
rect 2446 2301 2447 2307
rect 2453 2301 2454 2307
rect 2446 2163 2454 2301
rect 2446 2157 2447 2163
rect 2453 2157 2454 2163
rect 2446 2015 2454 2157
rect 2446 2009 2447 2015
rect 2453 2009 2454 2015
rect 2446 1879 2454 2009
rect 2446 1873 2447 1879
rect 2453 1873 2454 1879
rect 2446 1739 2454 1873
rect 2446 1733 2447 1739
rect 2453 1733 2454 1739
rect 2446 1603 2454 1733
rect 2446 1597 2447 1603
rect 2453 1597 2454 1603
rect 2446 1463 2454 1597
rect 2446 1457 2447 1463
rect 2453 1457 2454 1463
rect 2446 163 2454 1457
rect 2446 157 2447 163
rect 2453 157 2454 163
rect 2446 72 2454 157
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__133
timestamp 1731220645
transform 1 0 2400 0 -1 2504
box 7 3 12 24
use welltap_svt  __well_tap__132
timestamp 1731220645
transform 1 0 1272 0 -1 2504
box 7 3 12 24
use welltap_svt  __well_tap__131
timestamp 1731220645
transform 1 0 2400 0 1 2384
box 7 3 12 24
use welltap_svt  __well_tap__130
timestamp 1731220645
transform 1 0 1272 0 1 2384
box 7 3 12 24
use welltap_svt  __well_tap__129
timestamp 1731220645
transform 1 0 2400 0 -1 2368
box 7 3 12 24
use welltap_svt  __well_tap__128
timestamp 1731220645
transform 1 0 1272 0 -1 2368
box 7 3 12 24
use welltap_svt  __well_tap__127
timestamp 1731220645
transform 1 0 2400 0 1 2244
box 7 3 12 24
use welltap_svt  __well_tap__126
timestamp 1731220645
transform 1 0 1272 0 1 2244
box 7 3 12 24
use welltap_svt  __well_tap__125
timestamp 1731220645
transform 1 0 2400 0 -1 2220
box 7 3 12 24
use welltap_svt  __well_tap__124
timestamp 1731220645
transform 1 0 1272 0 -1 2220
box 7 3 12 24
use welltap_svt  __well_tap__123
timestamp 1731220645
transform 1 0 2400 0 1 2100
box 7 3 12 24
use welltap_svt  __well_tap__122
timestamp 1731220645
transform 1 0 1272 0 1 2100
box 7 3 12 24
use welltap_svt  __well_tap__121
timestamp 1731220645
transform 1 0 2400 0 -1 2080
box 7 3 12 24
use welltap_svt  __well_tap__120
timestamp 1731220645
transform 1 0 1272 0 -1 2080
box 7 3 12 24
use welltap_svt  __well_tap__119
timestamp 1731220645
transform 1 0 2400 0 1 1952
box 7 3 12 24
use welltap_svt  __well_tap__118
timestamp 1731220645
transform 1 0 1272 0 1 1952
box 7 3 12 24
use welltap_svt  __well_tap__117
timestamp 1731220645
transform 1 0 2400 0 -1 1936
box 7 3 12 24
use welltap_svt  __well_tap__116
timestamp 1731220645
transform 1 0 1272 0 -1 1936
box 7 3 12 24
use welltap_svt  __well_tap__115
timestamp 1731220645
transform 1 0 2400 0 1 1816
box 7 3 12 24
use welltap_svt  __well_tap__114
timestamp 1731220645
transform 1 0 1272 0 1 1816
box 7 3 12 24
use welltap_svt  __well_tap__113
timestamp 1731220645
transform 1 0 2400 0 -1 1796
box 7 3 12 24
use welltap_svt  __well_tap__112
timestamp 1731220645
transform 1 0 1272 0 -1 1796
box 7 3 12 24
use welltap_svt  __well_tap__111
timestamp 1731220645
transform 1 0 2400 0 1 1676
box 7 3 12 24
use welltap_svt  __well_tap__110
timestamp 1731220645
transform 1 0 1272 0 1 1676
box 7 3 12 24
use welltap_svt  __well_tap__109
timestamp 1731220645
transform 1 0 2400 0 -1 1660
box 7 3 12 24
use welltap_svt  __well_tap__108
timestamp 1731220645
transform 1 0 1272 0 -1 1660
box 7 3 12 24
use welltap_svt  __well_tap__107
timestamp 1731220645
transform 1 0 2400 0 1 1540
box 7 3 12 24
use welltap_svt  __well_tap__106
timestamp 1731220645
transform 1 0 1272 0 1 1540
box 7 3 12 24
use welltap_svt  __well_tap__105
timestamp 1731220645
transform 1 0 2400 0 -1 1520
box 7 3 12 24
use welltap_svt  __well_tap__104
timestamp 1731220645
transform 1 0 1272 0 -1 1520
box 7 3 12 24
use welltap_svt  __well_tap__103
timestamp 1731220645
transform 1 0 2400 0 1 1400
box 7 3 12 24
use welltap_svt  __well_tap__102
timestamp 1731220645
transform 1 0 1272 0 1 1400
box 7 3 12 24
use welltap_svt  __well_tap__101
timestamp 1731220645
transform 1 0 2400 0 -1 1376
box 7 3 12 24
use welltap_svt  __well_tap__100
timestamp 1731220645
transform 1 0 1272 0 -1 1376
box 7 3 12 24
use welltap_svt  __well_tap__99
timestamp 1731220645
transform 1 0 2400 0 1 1256
box 7 3 12 24
use welltap_svt  __well_tap__98
timestamp 1731220645
transform 1 0 1272 0 1 1256
box 7 3 12 24
use welltap_svt  __well_tap__97
timestamp 1731220645
transform 1 0 2400 0 -1 1232
box 7 3 12 24
use welltap_svt  __well_tap__96
timestamp 1731220645
transform 1 0 1272 0 -1 1232
box 7 3 12 24
use welltap_svt  __well_tap__95
timestamp 1731220645
transform 1 0 2400 0 1 1112
box 7 3 12 24
use welltap_svt  __well_tap__94
timestamp 1731220645
transform 1 0 1272 0 1 1112
box 7 3 12 24
use welltap_svt  __well_tap__93
timestamp 1731220645
transform 1 0 2400 0 -1 1096
box 7 3 12 24
use welltap_svt  __well_tap__92
timestamp 1731220645
transform 1 0 1272 0 -1 1096
box 7 3 12 24
use welltap_svt  __well_tap__91
timestamp 1731220645
transform 1 0 2400 0 1 976
box 7 3 12 24
use welltap_svt  __well_tap__90
timestamp 1731220645
transform 1 0 1272 0 1 976
box 7 3 12 24
use welltap_svt  __well_tap__89
timestamp 1731220645
transform 1 0 2400 0 -1 952
box 7 3 12 24
use welltap_svt  __well_tap__88
timestamp 1731220645
transform 1 0 1272 0 -1 952
box 7 3 12 24
use welltap_svt  __well_tap__87
timestamp 1731220645
transform 1 0 2400 0 1 832
box 7 3 12 24
use welltap_svt  __well_tap__86
timestamp 1731220645
transform 1 0 1272 0 1 832
box 7 3 12 24
use welltap_svt  __well_tap__85
timestamp 1731220645
transform 1 0 2400 0 -1 804
box 7 3 12 24
use welltap_svt  __well_tap__84
timestamp 1731220645
transform 1 0 1272 0 -1 804
box 7 3 12 24
use welltap_svt  __well_tap__83
timestamp 1731220645
transform 1 0 2400 0 1 684
box 7 3 12 24
use welltap_svt  __well_tap__82
timestamp 1731220645
transform 1 0 1272 0 1 684
box 7 3 12 24
use welltap_svt  __well_tap__81
timestamp 1731220645
transform 1 0 2400 0 -1 664
box 7 3 12 24
use welltap_svt  __well_tap__80
timestamp 1731220645
transform 1 0 1272 0 -1 664
box 7 3 12 24
use welltap_svt  __well_tap__79
timestamp 1731220645
transform 1 0 2400 0 1 540
box 7 3 12 24
use welltap_svt  __well_tap__78
timestamp 1731220645
transform 1 0 1272 0 1 540
box 7 3 12 24
use welltap_svt  __well_tap__77
timestamp 1731220645
transform 1 0 2400 0 -1 524
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220645
transform 1 0 1272 0 -1 524
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220645
transform 1 0 2400 0 1 400
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220645
transform 1 0 1272 0 1 400
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220645
transform 1 0 2400 0 -1 380
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220645
transform 1 0 1272 0 -1 380
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220645
transform 1 0 2400 0 1 256
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220645
transform 1 0 1272 0 1 256
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220645
transform 1 0 2400 0 -1 236
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220645
transform 1 0 1272 0 -1 236
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220645
transform 1 0 2400 0 1 100
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220645
transform 1 0 1272 0 1 100
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220645
transform 1 0 1232 0 1 2440
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220645
transform 1 0 104 0 1 2440
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220645
transform 1 0 1232 0 -1 2424
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220645
transform 1 0 104 0 -1 2424
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220645
transform 1 0 1232 0 1 2296
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220645
transform 1 0 104 0 1 2296
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220645
transform 1 0 1232 0 -1 2276
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220645
transform 1 0 104 0 -1 2276
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220645
transform 1 0 1232 0 1 2156
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220645
transform 1 0 104 0 1 2156
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220645
transform 1 0 1232 0 -1 2132
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220645
transform 1 0 104 0 -1 2132
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220645
transform 1 0 1232 0 1 2012
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220645
transform 1 0 104 0 1 2012
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220645
transform 1 0 1232 0 -1 1988
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220645
transform 1 0 104 0 -1 1988
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220645
transform 1 0 1232 0 1 1864
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220645
transform 1 0 104 0 1 1864
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220645
transform 1 0 1232 0 -1 1840
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220645
transform 1 0 104 0 -1 1840
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220645
transform 1 0 1232 0 1 1720
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220645
transform 1 0 104 0 1 1720
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220645
transform 1 0 1232 0 -1 1700
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220645
transform 1 0 104 0 -1 1700
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220645
transform 1 0 1232 0 1 1576
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220645
transform 1 0 104 0 1 1576
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220645
transform 1 0 1232 0 -1 1552
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220645
transform 1 0 104 0 -1 1552
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220645
transform 1 0 1232 0 1 1392
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220645
transform 1 0 104 0 1 1392
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220645
transform 1 0 1232 0 -1 1376
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220645
transform 1 0 104 0 -1 1376
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220645
transform 1 0 1232 0 1 1252
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220645
transform 1 0 104 0 1 1252
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220645
transform 1 0 1232 0 -1 1232
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220645
transform 1 0 104 0 -1 1232
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220645
transform 1 0 1232 0 1 1112
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220645
transform 1 0 104 0 1 1112
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220645
transform 1 0 1232 0 -1 1092
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220645
transform 1 0 104 0 -1 1092
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220645
transform 1 0 1232 0 1 972
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220645
transform 1 0 104 0 1 972
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220645
transform 1 0 1232 0 -1 956
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220645
transform 1 0 104 0 -1 956
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220645
transform 1 0 1232 0 1 828
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220645
transform 1 0 104 0 1 828
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220645
transform 1 0 1232 0 -1 812
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220645
transform 1 0 104 0 -1 812
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220645
transform 1 0 1232 0 1 688
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220645
transform 1 0 104 0 1 688
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220645
transform 1 0 1232 0 -1 668
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220645
transform 1 0 104 0 -1 668
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220645
transform 1 0 1232 0 1 540
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220645
transform 1 0 104 0 1 540
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220645
transform 1 0 1232 0 -1 516
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220645
transform 1 0 104 0 -1 516
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220645
transform 1 0 1232 0 1 396
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220645
transform 1 0 104 0 1 396
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220645
transform 1 0 1232 0 -1 380
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220645
transform 1 0 104 0 -1 380
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220645
transform 1 0 1232 0 1 256
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220645
transform 1 0 104 0 1 256
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220645
transform 1 0 1232 0 -1 232
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220645
transform 1 0 104 0 -1 232
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220645
transform 1 0 1232 0 1 92
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220645
transform 1 0 104 0 1 92
box 7 3 12 24
use _0_0std_0_0cells_0_0NOR2X2  tst_5999_6
timestamp 1731220645
transform 1 0 2264 0 1 92
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5998_6
timestamp 1731220645
transform 1 0 2312 0 1 92
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5997_6
timestamp 1731220645
transform 1 0 2352 0 1 92
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5996_6
timestamp 1731220645
transform 1 0 2352 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5995_6
timestamp 1731220645
transform 1 0 2352 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5994_6
timestamp 1731220645
transform 1 0 2312 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5993_6
timestamp 1731220645
transform 1 0 2352 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5992_6
timestamp 1731220645
transform 1 0 2288 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5991_6
timestamp 1731220645
transform 1 0 2352 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5990_6
timestamp 1731220645
transform 1 0 2352 0 -1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5989_6
timestamp 1731220645
transform 1 0 2352 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5988_6
timestamp 1731220645
transform 1 0 2352 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5987_6
timestamp 1731220645
transform 1 0 2352 0 1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5986_6
timestamp 1731220645
transform 1 0 2352 0 -1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5985_6
timestamp 1731220645
transform 1 0 2296 0 -1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5984_6
timestamp 1731220645
transform 1 0 2216 0 -1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5983_6
timestamp 1731220645
transform 1 0 2304 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5982_6
timestamp 1731220645
transform 1 0 2280 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5981_6
timestamp 1731220645
transform 1 0 2280 0 -1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5980_6
timestamp 1731220645
transform 1 0 2184 0 -1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5979_6
timestamp 1731220645
transform 1 0 2096 0 -1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5978_6
timestamp 1731220645
transform 1 0 2208 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5977_6
timestamp 1731220645
transform 1 0 2128 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5976_6
timestamp 1731220645
transform 1 0 2048 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5975_6
timestamp 1731220645
transform 1 0 2032 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5974_6
timestamp 1731220645
transform 1 0 1960 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5973_6
timestamp 1731220645
transform 1 0 2104 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5972_6
timestamp 1731220645
transform 1 0 2168 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5971_6
timestamp 1731220645
transform 1 0 2232 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5970_6
timestamp 1731220645
transform 1 0 2296 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5969_6
timestamp 1731220645
transform 1 0 2248 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5968_6
timestamp 1731220645
transform 1 0 2184 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5967_6
timestamp 1731220645
transform 1 0 2128 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5966_6
timestamp 1731220645
transform 1 0 2064 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5965_6
timestamp 1731220645
transform 1 0 2064 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5964_6
timestamp 1731220645
transform 1 0 2160 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5963_6
timestamp 1731220645
transform 1 0 2264 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5962_6
timestamp 1731220645
transform 1 0 2208 0 1 92
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5961_6
timestamp 1731220645
transform 1 0 2152 0 1 92
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5960_6
timestamp 1731220645
transform 1 0 2104 0 1 92
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5959_6
timestamp 1731220645
transform 1 0 2056 0 1 92
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5958_6
timestamp 1731220645
transform 1 0 2008 0 1 92
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5957_6
timestamp 1731220645
transform 1 0 1960 0 1 92
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5956_6
timestamp 1731220645
transform 1 0 1912 0 1 92
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5955_6
timestamp 1731220645
transform 1 0 1864 0 1 92
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5954_6
timestamp 1731220645
transform 1 0 1816 0 1 92
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5953_6
timestamp 1731220645
transform 1 0 1760 0 1 92
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5952_6
timestamp 1731220645
transform 1 0 1704 0 1 92
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5951_6
timestamp 1731220645
transform 1 0 1968 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5950_6
timestamp 1731220645
transform 1 0 1880 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5949_6
timestamp 1731220645
transform 1 0 1800 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5948_6
timestamp 1731220645
transform 1 0 1728 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5947_6
timestamp 1731220645
transform 1 0 2000 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5946_6
timestamp 1731220645
transform 1 0 1928 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5945_6
timestamp 1731220645
transform 1 0 1856 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5944_6
timestamp 1731220645
transform 1 0 1792 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5943_6
timestamp 1731220645
transform 1 0 1808 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5942_6
timestamp 1731220645
transform 1 0 1728 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5941_6
timestamp 1731220645
transform 1 0 1656 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5940_6
timestamp 1731220645
transform 1 0 1584 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5939_6
timestamp 1731220645
transform 1 0 1656 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5938_6
timestamp 1731220645
transform 1 0 1888 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5937_6
timestamp 1731220645
transform 1 0 1968 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5936_6
timestamp 1731220645
transform 1 0 1888 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5935_6
timestamp 1731220645
transform 1 0 1808 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5934_6
timestamp 1731220645
transform 1 0 1728 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5933_6
timestamp 1731220645
transform 1 0 1688 0 -1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5932_6
timestamp 1731220645
transform 1 0 1792 0 -1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5931_6
timestamp 1731220645
transform 1 0 2000 0 -1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5930_6
timestamp 1731220645
transform 1 0 1896 0 -1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5929_6
timestamp 1731220645
transform 1 0 1840 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5928_6
timestamp 1731220645
transform 1 0 1784 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5927_6
timestamp 1731220645
transform 1 0 1904 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5926_6
timestamp 1731220645
transform 1 0 1968 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5925_6
timestamp 1731220645
transform 1 0 2192 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5924_6
timestamp 1731220645
transform 1 0 2112 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5923_6
timestamp 1731220645
transform 1 0 2040 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5922_6
timestamp 1731220645
transform 1 0 1968 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5921_6
timestamp 1731220645
transform 1 0 1888 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5920_6
timestamp 1731220645
transform 1 0 1808 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5919_6
timestamp 1731220645
transform 1 0 2040 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5918_6
timestamp 1731220645
transform 1 0 2104 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5917_6
timestamp 1731220645
transform 1 0 2168 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5916_6
timestamp 1731220645
transform 1 0 2232 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5915_6
timestamp 1731220645
transform 1 0 2272 0 1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5914_6
timestamp 1731220645
transform 1 0 2168 0 1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5913_6
timestamp 1731220645
transform 1 0 2072 0 1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5912_6
timestamp 1731220645
transform 1 0 1984 0 1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5911_6
timestamp 1731220645
transform 1 0 1904 0 1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5910_6
timestamp 1731220645
transform 1 0 1824 0 1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5909_6
timestamp 1731220645
transform 1 0 2136 0 -1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5908_6
timestamp 1731220645
transform 1 0 2064 0 -1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5907_6
timestamp 1731220645
transform 1 0 1992 0 -1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5906_6
timestamp 1731220645
transform 1 0 1928 0 -1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5905_6
timestamp 1731220645
transform 1 0 1864 0 -1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5904_6
timestamp 1731220645
transform 1 0 1808 0 -1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5903_6
timestamp 1731220645
transform 1 0 1752 0 -1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5902_6
timestamp 1731220645
transform 1 0 1984 0 1 824
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5901_6
timestamp 1731220645
transform 1 0 1912 0 1 824
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5900_6
timestamp 1731220645
transform 1 0 1840 0 1 824
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5899_6
timestamp 1731220645
transform 1 0 1768 0 1 824
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5898_6
timestamp 1731220645
transform 1 0 1760 0 -1 960
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5897_6
timestamp 1731220645
transform 1 0 1848 0 -1 960
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5896_6
timestamp 1731220645
transform 1 0 1936 0 -1 960
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5895_6
timestamp 1731220645
transform 1 0 2008 0 1 968
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5894_6
timestamp 1731220645
transform 1 0 1936 0 1 968
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5893_6
timestamp 1731220645
transform 1 0 1872 0 1 968
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5892_6
timestamp 1731220645
transform 1 0 1816 0 1 968
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5891_6
timestamp 1731220645
transform 1 0 1768 0 -1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5890_6
timestamp 1731220645
transform 1 0 1816 0 -1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5889_6
timestamp 1731220645
transform 1 0 1864 0 -1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5888_6
timestamp 1731220645
transform 1 0 1912 0 -1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5887_6
timestamp 1731220645
transform 1 0 1960 0 -1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5886_6
timestamp 1731220645
transform 1 0 2008 0 -1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5885_6
timestamp 1731220645
transform 1 0 2056 0 -1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5884_6
timestamp 1731220645
transform 1 0 2112 0 -1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5883_6
timestamp 1731220645
transform 1 0 2088 0 1 968
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5882_6
timestamp 1731220645
transform 1 0 2096 0 -1 960
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5881_6
timestamp 1731220645
transform 1 0 2016 0 -1 960
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5880_6
timestamp 1731220645
transform 1 0 2056 0 1 824
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5879_6
timestamp 1731220645
transform 1 0 2128 0 1 824
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5878_6
timestamp 1731220645
transform 1 0 2208 0 1 824
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5877_6
timestamp 1731220645
transform 1 0 2288 0 1 824
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5876_6
timestamp 1731220645
transform 1 0 2264 0 -1 960
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5875_6
timestamp 1731220645
transform 1 0 2176 0 -1 960
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5874_6
timestamp 1731220645
transform 1 0 2168 0 1 968
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5873_6
timestamp 1731220645
transform 1 0 2248 0 1 968
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5872_6
timestamp 1731220645
transform 1 0 2224 0 -1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5871_6
timestamp 1731220645
transform 1 0 2168 0 -1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5870_6
timestamp 1731220645
transform 1 0 2072 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5869_6
timestamp 1731220645
transform 1 0 1992 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5868_6
timestamp 1731220645
transform 1 0 1896 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5867_6
timestamp 1731220645
transform 1 0 2144 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5866_6
timestamp 1731220645
transform 1 0 2064 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5865_6
timestamp 1731220645
transform 1 0 1976 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5864_6
timestamp 1731220645
transform 1 0 1880 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5863_6
timestamp 1731220645
transform 1 0 1784 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5862_6
timestamp 1731220645
transform 1 0 2192 0 1 1248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5861_6
timestamp 1731220645
transform 1 0 2112 0 1 1248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5860_6
timestamp 1731220645
transform 1 0 2032 0 1 1248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5859_6
timestamp 1731220645
transform 1 0 1960 0 1 1248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5858_6
timestamp 1731220645
transform 1 0 1896 0 1 1248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5857_6
timestamp 1731220645
transform 1 0 1840 0 1 1248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5856_6
timestamp 1731220645
transform 1 0 1784 0 1 1248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5855_6
timestamp 1731220645
transform 1 0 1760 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5854_6
timestamp 1731220645
transform 1 0 1840 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5853_6
timestamp 1731220645
transform 1 0 1928 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5852_6
timestamp 1731220645
transform 1 0 2104 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5851_6
timestamp 1731220645
transform 1 0 2016 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5850_6
timestamp 1731220645
transform 1 0 1936 0 1 1392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5849_6
timestamp 1731220645
transform 1 0 1872 0 1 1392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5848_6
timestamp 1731220645
transform 1 0 1800 0 1 1392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5847_6
timestamp 1731220645
transform 1 0 1992 0 1 1392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5846_6
timestamp 1731220645
transform 1 0 2040 0 1 1392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5845_6
timestamp 1731220645
transform 1 0 2088 0 1 1392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5844_6
timestamp 1731220645
transform 1 0 2136 0 1 1392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5843_6
timestamp 1731220645
transform 1 0 2184 0 1 1392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5842_6
timestamp 1731220645
transform 1 0 2232 0 1 1392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5841_6
timestamp 1731220645
transform 1 0 2272 0 1 1392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5840_6
timestamp 1731220645
transform 1 0 2312 0 1 1392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5839_6
timestamp 1731220645
transform 1 0 2280 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5838_6
timestamp 1731220645
transform 1 0 2192 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5837_6
timestamp 1731220645
transform 1 0 2280 0 1 1248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5836_6
timestamp 1731220645
transform 1 0 2216 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5835_6
timestamp 1731220645
transform 1 0 2152 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5834_6
timestamp 1731220645
transform 1 0 2224 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5833_6
timestamp 1731220645
transform 1 0 2296 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5832_6
timestamp 1731220645
transform 1 0 2352 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5831_6
timestamp 1731220645
transform 1 0 2296 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5830_6
timestamp 1731220645
transform 1 0 2352 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5829_6
timestamp 1731220645
transform 1 0 2352 0 1 1248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5828_6
timestamp 1731220645
transform 1 0 2352 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5827_6
timestamp 1731220645
transform 1 0 2352 0 1 1392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5826_6
timestamp 1731220645
transform 1 0 2352 0 -1 1528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5825_6
timestamp 1731220645
transform 1 0 2208 0 -1 1528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5824_6
timestamp 1731220645
transform 1 0 2352 0 1 1532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5823_6
timestamp 1731220645
transform 1 0 2312 0 1 1532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5822_6
timestamp 1731220645
transform 1 0 2264 0 1 1532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5821_6
timestamp 1731220645
transform 1 0 2208 0 1 1532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5820_6
timestamp 1731220645
transform 1 0 2160 0 1 1532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5819_6
timestamp 1731220645
transform 1 0 2104 0 1 1532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5818_6
timestamp 1731220645
transform 1 0 2040 0 1 1532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5817_6
timestamp 1731220645
transform 1 0 1976 0 1 1532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5816_6
timestamp 1731220645
transform 1 0 1904 0 1 1532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5815_6
timestamp 1731220645
transform 1 0 2216 0 -1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5814_6
timestamp 1731220645
transform 1 0 2152 0 -1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5813_6
timestamp 1731220645
transform 1 0 2088 0 -1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5812_6
timestamp 1731220645
transform 1 0 2024 0 -1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5811_6
timestamp 1731220645
transform 1 0 1960 0 -1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5810_6
timestamp 1731220645
transform 1 0 1888 0 -1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5809_6
timestamp 1731220645
transform 1 0 1808 0 -1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5808_6
timestamp 1731220645
transform 1 0 2056 0 1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5807_6
timestamp 1731220645
transform 1 0 1992 0 1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5806_6
timestamp 1731220645
transform 1 0 1928 0 1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5805_6
timestamp 1731220645
transform 1 0 1864 0 1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5804_6
timestamp 1731220645
transform 1 0 1800 0 1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5803_6
timestamp 1731220645
transform 1 0 1728 0 1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5802_6
timestamp 1731220645
transform 1 0 1952 0 -1 1804
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5801_6
timestamp 1731220645
transform 1 0 1888 0 -1 1804
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5800_6
timestamp 1731220645
transform 1 0 1832 0 -1 1804
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5799_6
timestamp 1731220645
transform 1 0 1776 0 -1 1804
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5798_6
timestamp 1731220645
transform 1 0 1720 0 -1 1804
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5797_6
timestamp 1731220645
transform 1 0 1656 0 -1 1804
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5796_6
timestamp 1731220645
transform 1 0 1680 0 1 1808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5795_6
timestamp 1731220645
transform 1 0 1760 0 1 1808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5794_6
timestamp 1731220645
transform 1 0 1856 0 1 1808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5793_6
timestamp 1731220645
transform 1 0 2216 0 1 1808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5792_6
timestamp 1731220645
transform 1 0 2088 0 1 1808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5791_6
timestamp 1731220645
transform 1 0 1968 0 1 1808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5790_6
timestamp 1731220645
transform 1 0 1928 0 -1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5789_6
timestamp 1731220645
transform 1 0 1856 0 -1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5788_6
timestamp 1731220645
transform 1 0 1784 0 -1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5787_6
timestamp 1731220645
transform 1 0 2000 0 -1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5786_6
timestamp 1731220645
transform 1 0 2144 0 -1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5785_6
timestamp 1731220645
transform 1 0 2072 0 -1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5784_6
timestamp 1731220645
transform 1 0 1992 0 1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5783_6
timestamp 1731220645
transform 1 0 1912 0 1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5782_6
timestamp 1731220645
transform 1 0 2064 0 1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5781_6
timestamp 1731220645
transform 1 0 2128 0 1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5780_6
timestamp 1731220645
transform 1 0 2184 0 1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5779_6
timestamp 1731220645
transform 1 0 2160 0 -1 2088
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5778_6
timestamp 1731220645
transform 1 0 2088 0 -1 2088
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5777_6
timestamp 1731220645
transform 1 0 2232 0 -1 2088
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5776_6
timestamp 1731220645
transform 1 0 2304 0 -1 2088
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5775_6
timestamp 1731220645
transform 1 0 2312 0 1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5774_6
timestamp 1731220645
transform 1 0 2352 0 1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5773_6
timestamp 1731220645
transform 1 0 2352 0 -1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5772_6
timestamp 1731220645
transform 1 0 2352 0 1 1808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5771_6
timestamp 1731220645
transform 1 0 2296 0 -1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5770_6
timestamp 1731220645
transform 1 0 2216 0 -1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5769_6
timestamp 1731220645
transform 1 0 2248 0 1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5768_6
timestamp 1731220645
transform 1 0 2352 0 -1 2088
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5767_6
timestamp 1731220645
transform 1 0 2352 0 1 2092
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5766_6
timestamp 1731220645
transform 1 0 2304 0 1 2092
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5765_6
timestamp 1731220645
transform 1 0 2352 0 -1 2228
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5764_6
timestamp 1731220645
transform 1 0 2352 0 1 2236
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5763_6
timestamp 1731220645
transform 1 0 2288 0 1 2236
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5762_6
timestamp 1731220645
transform 1 0 2296 0 -1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5761_6
timestamp 1731220645
transform 1 0 2352 0 -1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5760_6
timestamp 1731220645
transform 1 0 2328 0 1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5759_6
timestamp 1731220645
transform 1 0 2216 0 -1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5758_6
timestamp 1731220645
transform 1 0 2200 0 1 2236
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5757_6
timestamp 1731220645
transform 1 0 2120 0 1 2236
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5756_6
timestamp 1731220645
transform 1 0 2176 0 -1 2228
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5755_6
timestamp 1731220645
transform 1 0 2272 0 -1 2228
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5754_6
timestamp 1731220645
transform 1 0 2232 0 1 2092
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5753_6
timestamp 1731220645
transform 1 0 2168 0 1 2092
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5752_6
timestamp 1731220645
transform 1 0 2104 0 1 2092
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5751_6
timestamp 1731220645
transform 1 0 2008 0 -1 2088
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5750_6
timestamp 1731220645
transform 1 0 1928 0 -1 2088
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5749_6
timestamp 1731220645
transform 1 0 2040 0 1 2092
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5748_6
timestamp 1731220645
transform 1 0 1968 0 1 2092
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5747_6
timestamp 1731220645
transform 1 0 1888 0 1 2092
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5746_6
timestamp 1731220645
transform 1 0 1808 0 1 2092
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5745_6
timestamp 1731220645
transform 1 0 2088 0 -1 2228
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5744_6
timestamp 1731220645
transform 1 0 2008 0 -1 2228
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5743_6
timestamp 1731220645
transform 1 0 1928 0 -1 2228
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5742_6
timestamp 1731220645
transform 1 0 1848 0 -1 2228
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5741_6
timestamp 1731220645
transform 1 0 1776 0 -1 2228
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5740_6
timestamp 1731220645
transform 1 0 2040 0 1 2236
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5739_6
timestamp 1731220645
transform 1 0 1960 0 1 2236
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5738_6
timestamp 1731220645
transform 1 0 1888 0 1 2236
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5737_6
timestamp 1731220645
transform 1 0 1816 0 1 2236
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5736_6
timestamp 1731220645
transform 1 0 1752 0 1 2236
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5735_6
timestamp 1731220645
transform 1 0 1768 0 -1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5734_6
timestamp 1731220645
transform 1 0 1848 0 -1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5733_6
timestamp 1731220645
transform 1 0 1920 0 -1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5732_6
timestamp 1731220645
transform 1 0 1992 0 -1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5731_6
timestamp 1731220645
transform 1 0 2064 0 -1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5730_6
timestamp 1731220645
transform 1 0 2136 0 -1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5729_6
timestamp 1731220645
transform 1 0 2240 0 1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5728_6
timestamp 1731220645
transform 1 0 2152 0 1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5727_6
timestamp 1731220645
transform 1 0 2072 0 1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5726_6
timestamp 1731220645
transform 1 0 1992 0 1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5725_6
timestamp 1731220645
transform 1 0 1912 0 1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5724_6
timestamp 1731220645
transform 1 0 1832 0 1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5723_6
timestamp 1731220645
transform 1 0 1968 0 -1 2512
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5722_6
timestamp 1731220645
transform 1 0 1928 0 -1 2512
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5721_6
timestamp 1731220645
transform 1 0 1888 0 -1 2512
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5720_6
timestamp 1731220645
transform 1 0 1848 0 -1 2512
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5719_6
timestamp 1731220645
transform 1 0 1808 0 -1 2512
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5718_6
timestamp 1731220645
transform 1 0 1768 0 -1 2512
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5717_6
timestamp 1731220645
transform 1 0 1728 0 -1 2512
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5716_6
timestamp 1731220645
transform 1 0 1688 0 -1 2512
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5715_6
timestamp 1731220645
transform 1 0 1648 0 -1 2512
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5714_6
timestamp 1731220645
transform 1 0 1608 0 -1 2512
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5713_6
timestamp 1731220645
transform 1 0 1568 0 -1 2512
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5712_6
timestamp 1731220645
transform 1 0 1528 0 -1 2512
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5711_6
timestamp 1731220645
transform 1 0 1752 0 1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5710_6
timestamp 1731220645
transform 1 0 1672 0 1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5709_6
timestamp 1731220645
transform 1 0 1592 0 1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5708_6
timestamp 1731220645
transform 1 0 1512 0 1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5707_6
timestamp 1731220645
transform 1 0 1448 0 1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5706_6
timestamp 1731220645
transform 1 0 1392 0 1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5705_6
timestamp 1731220645
transform 1 0 1352 0 1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5704_6
timestamp 1731220645
transform 1 0 1352 0 -1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5703_6
timestamp 1731220645
transform 1 0 1400 0 -1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5702_6
timestamp 1731220645
transform 1 0 1464 0 -1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5701_6
timestamp 1731220645
transform 1 0 1536 0 -1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5700_6
timestamp 1731220645
transform 1 0 1688 0 -1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5699_6
timestamp 1731220645
transform 1 0 1608 0 -1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5698_6
timestamp 1731220645
transform 1 0 1576 0 1 2236
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5697_6
timestamp 1731220645
transform 1 0 1536 0 1 2236
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5696_6
timestamp 1731220645
transform 1 0 1496 0 1 2236
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5695_6
timestamp 1731220645
transform 1 0 1616 0 1 2236
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5694_6
timestamp 1731220645
transform 1 0 1696 0 1 2236
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5693_6
timestamp 1731220645
transform 1 0 1656 0 1 2236
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5692_6
timestamp 1731220645
transform 1 0 1632 0 -1 2228
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5691_6
timestamp 1731220645
transform 1 0 1704 0 -1 2228
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5690_6
timestamp 1731220645
transform 1 0 1720 0 1 2092
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5689_6
timestamp 1731220645
transform 1 0 1752 0 -1 2088
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5688_6
timestamp 1731220645
transform 1 0 1840 0 -1 2088
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5687_6
timestamp 1731220645
transform 1 0 1832 0 1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5686_6
timestamp 1731220645
transform 1 0 1744 0 1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5685_6
timestamp 1731220645
transform 1 0 1656 0 1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5684_6
timestamp 1731220645
transform 1 0 1704 0 -1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5683_6
timestamp 1731220645
transform 1 0 1616 0 -1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5682_6
timestamp 1731220645
transform 1 0 1528 0 -1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5681_6
timestamp 1731220645
transform 1 0 1488 0 1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5680_6
timestamp 1731220645
transform 1 0 1416 0 1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5679_6
timestamp 1731220645
transform 1 0 1568 0 1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5678_6
timestamp 1731220645
transform 1 0 1656 0 -1 2088
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5677_6
timestamp 1731220645
transform 1 0 1560 0 -1 2088
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5676_6
timestamp 1731220645
transform 1 0 1472 0 -1 2088
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5675_6
timestamp 1731220645
transform 1 0 1392 0 -1 2088
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5674_6
timestamp 1731220645
transform 1 0 1432 0 1 2092
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5673_6
timestamp 1731220645
transform 1 0 1528 0 1 2092
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5672_6
timestamp 1731220645
transform 1 0 1624 0 1 2092
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5671_6
timestamp 1731220645
transform 1 0 1560 0 -1 2228
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5670_6
timestamp 1731220645
transform 1 0 1488 0 -1 2228
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5669_6
timestamp 1731220645
transform 1 0 1424 0 -1 2228
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5668_6
timestamp 1731220645
transform 1 0 1376 0 -1 2228
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5667_6
timestamp 1731220645
transform 1 0 1336 0 -1 2228
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5666_6
timestamp 1731220645
transform 1 0 1296 0 -1 2228
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5665_6
timestamp 1731220645
transform 1 0 1344 0 1 2092
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5664_6
timestamp 1731220645
transform 1 0 1296 0 1 2092
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5663_6
timestamp 1731220645
transform 1 0 1296 0 -1 2088
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5662_6
timestamp 1731220645
transform 1 0 1336 0 -1 2088
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5661_6
timestamp 1731220645
transform 1 0 1344 0 1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5660_6
timestamp 1731220645
transform 1 0 1296 0 1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5659_6
timestamp 1731220645
transform 1 0 1296 0 -1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5658_6
timestamp 1731220645
transform 1 0 1352 0 -1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5657_6
timestamp 1731220645
transform 1 0 1440 0 -1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5656_6
timestamp 1731220645
transform 1 0 1408 0 1 1808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5655_6
timestamp 1731220645
transform 1 0 1352 0 1 1808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5654_6
timestamp 1731220645
transform 1 0 1304 0 1 1808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5653_6
timestamp 1731220645
transform 1 0 1472 0 1 1808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5652_6
timestamp 1731220645
transform 1 0 1536 0 1 1808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5651_6
timestamp 1731220645
transform 1 0 1608 0 1 1808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5650_6
timestamp 1731220645
transform 1 0 1592 0 -1 1804
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5649_6
timestamp 1731220645
transform 1 0 1528 0 -1 1804
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5648_6
timestamp 1731220645
transform 1 0 1464 0 -1 1804
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5647_6
timestamp 1731220645
transform 1 0 1400 0 -1 1804
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5646_6
timestamp 1731220645
transform 1 0 1416 0 1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5645_6
timestamp 1731220645
transform 1 0 1496 0 1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5644_6
timestamp 1731220645
transform 1 0 1576 0 1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5643_6
timestamp 1731220645
transform 1 0 1656 0 1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5642_6
timestamp 1731220645
transform 1 0 1720 0 -1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5641_6
timestamp 1731220645
transform 1 0 1632 0 -1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5640_6
timestamp 1731220645
transform 1 0 1536 0 -1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5639_6
timestamp 1731220645
transform 1 0 1472 0 1 1532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5638_6
timestamp 1731220645
transform 1 0 1560 0 1 1532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5637_6
timestamp 1731220645
transform 1 0 1648 0 1 1532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5636_6
timestamp 1731220645
transform 1 0 1736 0 1 1532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5635_6
timestamp 1731220645
transform 1 0 1824 0 1 1532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5634_6
timestamp 1731220645
transform 1 0 2040 0 -1 1528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5633_6
timestamp 1731220645
transform 1 0 1880 0 -1 1528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5632_6
timestamp 1731220645
transform 1 0 1736 0 -1 1528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5631_6
timestamp 1731220645
transform 1 0 1608 0 -1 1528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5630_6
timestamp 1731220645
transform 1 0 1720 0 1 1392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5629_6
timestamp 1731220645
transform 1 0 1632 0 1 1392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5628_6
timestamp 1731220645
transform 1 0 1544 0 1 1392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5627_6
timestamp 1731220645
transform 1 0 1528 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5626_6
timestamp 1731220645
transform 1 0 1600 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5625_6
timestamp 1731220645
transform 1 0 1680 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5624_6
timestamp 1731220645
transform 1 0 1728 0 1 1248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5623_6
timestamp 1731220645
transform 1 0 1672 0 1 1248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5622_6
timestamp 1731220645
transform 1 0 1616 0 1 1248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5621_6
timestamp 1731220645
transform 1 0 1576 0 1 1248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5620_6
timestamp 1731220645
transform 1 0 1456 0 1 1248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5619_6
timestamp 1731220645
transform 1 0 1416 0 1 1248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5618_6
timestamp 1731220645
transform 1 0 1376 0 1 1248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5617_6
timestamp 1731220645
transform 1 0 1336 0 1 1248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5616_6
timestamp 1731220645
transform 1 0 1296 0 1 1248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5615_6
timestamp 1731220645
transform 1 0 1296 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5614_6
timestamp 1731220645
transform 1 0 1184 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5613_6
timestamp 1731220645
transform 1 0 1136 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5612_6
timestamp 1731220645
transform 1 0 1072 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5611_6
timestamp 1731220645
transform 1 0 1184 0 1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5610_6
timestamp 1731220645
transform 1 0 1144 0 1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5609_6
timestamp 1731220645
transform 1 0 1096 0 1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5608_6
timestamp 1731220645
transform 1 0 1040 0 1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5607_6
timestamp 1731220645
transform 1 0 992 0 1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5606_6
timestamp 1731220645
transform 1 0 936 0 1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5605_6
timestamp 1731220645
transform 1 0 872 0 1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5604_6
timestamp 1731220645
transform 1 0 800 0 1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5603_6
timestamp 1731220645
transform 1 0 720 0 1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5602_6
timestamp 1731220645
transform 1 0 1008 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5601_6
timestamp 1731220645
transform 1 0 944 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5600_6
timestamp 1731220645
transform 1 0 880 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5599_6
timestamp 1731220645
transform 1 0 816 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5598_6
timestamp 1731220645
transform 1 0 744 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5597_6
timestamp 1731220645
transform 1 0 672 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5596_6
timestamp 1731220645
transform 1 0 992 0 1 1244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5595_6
timestamp 1731220645
transform 1 0 928 0 1 1244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5594_6
timestamp 1731220645
transform 1 0 872 0 1 1244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5593_6
timestamp 1731220645
transform 1 0 816 0 1 1244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5592_6
timestamp 1731220645
transform 1 0 760 0 1 1244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5591_6
timestamp 1731220645
transform 1 0 696 0 1 1244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5590_6
timestamp 1731220645
transform 1 0 632 0 1 1244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5589_6
timestamp 1731220645
transform 1 0 656 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5588_6
timestamp 1731220645
transform 1 0 736 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5587_6
timestamp 1731220645
transform 1 0 808 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5586_6
timestamp 1731220645
transform 1 0 872 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5585_6
timestamp 1731220645
transform 1 0 936 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5584_6
timestamp 1731220645
transform 1 0 1000 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5583_6
timestamp 1731220645
transform 1 0 1064 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5582_6
timestamp 1731220645
transform 1 0 1184 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5581_6
timestamp 1731220645
transform 1 0 1136 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5580_6
timestamp 1731220645
transform 1 0 1064 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5579_6
timestamp 1731220645
transform 1 0 992 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5578_6
timestamp 1731220645
transform 1 0 912 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5577_6
timestamp 1731220645
transform 1 0 832 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5576_6
timestamp 1731220645
transform 1 0 736 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5575_6
timestamp 1731220645
transform 1 0 1040 0 -1 1100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5574_6
timestamp 1731220645
transform 1 0 976 0 -1 1100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5573_6
timestamp 1731220645
transform 1 0 912 0 -1 1100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5572_6
timestamp 1731220645
transform 1 0 856 0 -1 1100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5571_6
timestamp 1731220645
transform 1 0 792 0 -1 1100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5570_6
timestamp 1731220645
transform 1 0 728 0 -1 1100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5569_6
timestamp 1731220645
transform 1 0 656 0 -1 1100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5568_6
timestamp 1731220645
transform 1 0 1096 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5567_6
timestamp 1731220645
transform 1 0 992 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5566_6
timestamp 1731220645
transform 1 0 888 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5565_6
timestamp 1731220645
transform 1 0 800 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5564_6
timestamp 1731220645
transform 1 0 728 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5563_6
timestamp 1731220645
transform 1 0 664 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5562_6
timestamp 1731220645
transform 1 0 616 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5561_6
timestamp 1731220645
transform 1 0 848 0 -1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5560_6
timestamp 1731220645
transform 1 0 776 0 -1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5559_6
timestamp 1731220645
transform 1 0 704 0 -1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5558_6
timestamp 1731220645
transform 1 0 632 0 -1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5557_6
timestamp 1731220645
transform 1 0 568 0 -1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5556_6
timestamp 1731220645
transform 1 0 512 0 -1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5555_6
timestamp 1731220645
transform 1 0 456 0 -1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5554_6
timestamp 1731220645
transform 1 0 568 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5553_6
timestamp 1731220645
transform 1 0 512 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5552_6
timestamp 1731220645
transform 1 0 456 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5551_6
timestamp 1731220645
transform 1 0 392 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5550_6
timestamp 1731220645
transform 1 0 320 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5549_6
timestamp 1731220645
transform 1 0 576 0 -1 1100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5548_6
timestamp 1731220645
transform 1 0 496 0 -1 1100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5547_6
timestamp 1731220645
transform 1 0 408 0 -1 1100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5546_6
timestamp 1731220645
transform 1 0 320 0 -1 1100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5545_6
timestamp 1731220645
transform 1 0 632 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5544_6
timestamp 1731220645
transform 1 0 528 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5543_6
timestamp 1731220645
transform 1 0 424 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5542_6
timestamp 1731220645
transform 1 0 320 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5541_6
timestamp 1731220645
transform 1 0 232 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5540_6
timestamp 1731220645
transform 1 0 304 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5539_6
timestamp 1731220645
transform 1 0 392 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5538_6
timestamp 1731220645
transform 1 0 480 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5537_6
timestamp 1731220645
transform 1 0 568 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5536_6
timestamp 1731220645
transform 1 0 560 0 1 1244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5535_6
timestamp 1731220645
transform 1 0 488 0 1 1244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5534_6
timestamp 1731220645
transform 1 0 416 0 1 1244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5533_6
timestamp 1731220645
transform 1 0 344 0 1 1244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5532_6
timestamp 1731220645
transform 1 0 280 0 1 1244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5531_6
timestamp 1731220645
transform 1 0 592 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5530_6
timestamp 1731220645
transform 1 0 512 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5529_6
timestamp 1731220645
transform 1 0 432 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5528_6
timestamp 1731220645
transform 1 0 360 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5527_6
timestamp 1731220645
transform 1 0 640 0 1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5526_6
timestamp 1731220645
transform 1 0 552 0 1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5525_6
timestamp 1731220645
transform 1 0 464 0 1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5524_6
timestamp 1731220645
transform 1 0 384 0 1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5523_6
timestamp 1731220645
transform 1 0 312 0 1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5522_6
timestamp 1731220645
transform 1 0 256 0 1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5521_6
timestamp 1731220645
transform 1 0 216 0 1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5520_6
timestamp 1731220645
transform 1 0 176 0 1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5519_6
timestamp 1731220645
transform 1 0 136 0 1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5518_6
timestamp 1731220645
transform 1 0 296 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5517_6
timestamp 1731220645
transform 1 0 240 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5516_6
timestamp 1731220645
transform 1 0 200 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5515_6
timestamp 1731220645
transform 1 0 160 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5514_6
timestamp 1731220645
transform 1 0 176 0 1 1244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5513_6
timestamp 1731220645
transform 1 0 224 0 1 1244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5512_6
timestamp 1731220645
transform 1 0 224 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5511_6
timestamp 1731220645
transform 1 0 168 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5510_6
timestamp 1731220645
transform 1 0 128 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5509_6
timestamp 1731220645
transform 1 0 128 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5508_6
timestamp 1731220645
transform 1 0 168 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5507_6
timestamp 1731220645
transform 1 0 128 0 -1 1100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5506_6
timestamp 1731220645
transform 1 0 240 0 -1 1100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5505_6
timestamp 1731220645
transform 1 0 168 0 -1 1100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5504_6
timestamp 1731220645
transform 1 0 168 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5503_6
timestamp 1731220645
transform 1 0 248 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5502_6
timestamp 1731220645
transform 1 0 248 0 -1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5501_6
timestamp 1731220645
transform 1 0 208 0 -1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5500_6
timestamp 1731220645
transform 1 0 296 0 -1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5499_6
timestamp 1731220645
transform 1 0 352 0 -1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5498_6
timestamp 1731220645
transform 1 0 408 0 -1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5497_6
timestamp 1731220645
transform 1 0 632 0 1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5496_6
timestamp 1731220645
transform 1 0 536 0 1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5495_6
timestamp 1731220645
transform 1 0 440 0 1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5494_6
timestamp 1731220645
transform 1 0 352 0 1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5493_6
timestamp 1731220645
transform 1 0 280 0 1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5492_6
timestamp 1731220645
transform 1 0 224 0 1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5491_6
timestamp 1731220645
transform 1 0 184 0 1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5490_6
timestamp 1731220645
transform 1 0 496 0 -1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5489_6
timestamp 1731220645
transform 1 0 408 0 -1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5488_6
timestamp 1731220645
transform 1 0 320 0 -1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5487_6
timestamp 1731220645
transform 1 0 232 0 -1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5486_6
timestamp 1731220645
transform 1 0 168 0 -1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5485_6
timestamp 1731220645
transform 1 0 128 0 -1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5484_6
timestamp 1731220645
transform 1 0 128 0 1 680
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5483_6
timestamp 1731220645
transform 1 0 184 0 1 680
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5482_6
timestamp 1731220645
transform 1 0 192 0 -1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5481_6
timestamp 1731220645
transform 1 0 128 0 -1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5480_6
timestamp 1731220645
transform 1 0 128 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5479_6
timestamp 1731220645
transform 1 0 184 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5478_6
timestamp 1731220645
transform 1 0 264 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5477_6
timestamp 1731220645
transform 1 0 256 0 -1 524
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5476_6
timestamp 1731220645
transform 1 0 184 0 -1 524
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5475_6
timestamp 1731220645
transform 1 0 128 0 -1 524
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5474_6
timestamp 1731220645
transform 1 0 176 0 1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5473_6
timestamp 1731220645
transform 1 0 216 0 1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5472_6
timestamp 1731220645
transform 1 0 256 0 1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5471_6
timestamp 1731220645
transform 1 0 280 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5470_6
timestamp 1731220645
transform 1 0 224 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5469_6
timestamp 1731220645
transform 1 0 168 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5468_6
timestamp 1731220645
transform 1 0 128 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5467_6
timestamp 1731220645
transform 1 0 248 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5466_6
timestamp 1731220645
transform 1 0 176 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5465_6
timestamp 1731220645
transform 1 0 128 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5464_6
timestamp 1731220645
transform 1 0 128 0 -1 240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5463_6
timestamp 1731220645
transform 1 0 168 0 -1 240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5462_6
timestamp 1731220645
transform 1 0 320 0 -1 240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5461_6
timestamp 1731220645
transform 1 0 240 0 -1 240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5460_6
timestamp 1731220645
transform 1 0 208 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5459_6
timestamp 1731220645
transform 1 0 168 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5458_6
timestamp 1731220645
transform 1 0 128 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5457_6
timestamp 1731220645
transform 1 0 248 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5456_6
timestamp 1731220645
transform 1 0 288 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5455_6
timestamp 1731220645
transform 1 0 328 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5454_6
timestamp 1731220645
transform 1 0 368 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5453_6
timestamp 1731220645
transform 1 0 416 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5452_6
timestamp 1731220645
transform 1 0 464 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5451_6
timestamp 1731220645
transform 1 0 576 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5450_6
timestamp 1731220645
transform 1 0 520 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5449_6
timestamp 1731220645
transform 1 0 488 0 -1 240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5448_6
timestamp 1731220645
transform 1 0 408 0 -1 240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5447_6
timestamp 1731220645
transform 1 0 568 0 -1 240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5446_6
timestamp 1731220645
transform 1 0 544 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5445_6
timestamp 1731220645
transform 1 0 496 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5444_6
timestamp 1731220645
transform 1 0 440 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5443_6
timestamp 1731220645
transform 1 0 384 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5442_6
timestamp 1731220645
transform 1 0 320 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5441_6
timestamp 1731220645
transform 1 0 336 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5440_6
timestamp 1731220645
transform 1 0 384 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5439_6
timestamp 1731220645
transform 1 0 432 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5438_6
timestamp 1731220645
transform 1 0 488 0 1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5437_6
timestamp 1731220645
transform 1 0 424 0 1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5436_6
timestamp 1731220645
transform 1 0 360 0 1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5435_6
timestamp 1731220645
transform 1 0 304 0 1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5434_6
timestamp 1731220645
transform 1 0 328 0 -1 524
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5433_6
timestamp 1731220645
transform 1 0 408 0 -1 524
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5432_6
timestamp 1731220645
transform 1 0 488 0 -1 524
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5431_6
timestamp 1731220645
transform 1 0 568 0 -1 524
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5430_6
timestamp 1731220645
transform 1 0 528 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5429_6
timestamp 1731220645
transform 1 0 440 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5428_6
timestamp 1731220645
transform 1 0 352 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5427_6
timestamp 1731220645
transform 1 0 696 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5426_6
timestamp 1731220645
transform 1 0 616 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5425_6
timestamp 1731220645
transform 1 0 552 0 -1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5424_6
timestamp 1731220645
transform 1 0 480 0 -1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5423_6
timestamp 1731220645
transform 1 0 408 0 -1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5422_6
timestamp 1731220645
transform 1 0 344 0 -1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5421_6
timestamp 1731220645
transform 1 0 272 0 -1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5420_6
timestamp 1731220645
transform 1 0 256 0 1 680
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5419_6
timestamp 1731220645
transform 1 0 328 0 1 680
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5418_6
timestamp 1731220645
transform 1 0 392 0 1 680
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5417_6
timestamp 1731220645
transform 1 0 448 0 1 680
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5416_6
timestamp 1731220645
transform 1 0 496 0 1 680
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5415_6
timestamp 1731220645
transform 1 0 536 0 1 680
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5414_6
timestamp 1731220645
transform 1 0 576 0 1 680
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5413_6
timestamp 1731220645
transform 1 0 616 0 1 680
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5412_6
timestamp 1731220645
transform 1 0 632 0 -1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5411_6
timestamp 1731220645
transform 1 0 704 0 -1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5410_6
timestamp 1731220645
transform 1 0 776 0 -1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5409_6
timestamp 1731220645
transform 1 0 760 0 1 680
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5408_6
timestamp 1731220645
transform 1 0 712 0 1 680
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5407_6
timestamp 1731220645
transform 1 0 664 0 1 680
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5406_6
timestamp 1731220645
transform 1 0 904 0 1 680
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5405_6
timestamp 1731220645
transform 1 0 856 0 1 680
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5404_6
timestamp 1731220645
transform 1 0 808 0 1 680
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5403_6
timestamp 1731220645
transform 1 0 736 0 -1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5402_6
timestamp 1731220645
transform 1 0 664 0 -1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5401_6
timestamp 1731220645
transform 1 0 584 0 -1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5400_6
timestamp 1731220645
transform 1 0 808 0 -1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5399_6
timestamp 1731220645
transform 1 0 1008 0 -1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5398_6
timestamp 1731220645
transform 1 0 936 0 -1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5397_6
timestamp 1731220645
transform 1 0 872 0 -1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5396_6
timestamp 1731220645
transform 1 0 800 0 1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5395_6
timestamp 1731220645
transform 1 0 720 0 1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5394_6
timestamp 1731220645
transform 1 0 880 0 1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5393_6
timestamp 1731220645
transform 1 0 952 0 1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5392_6
timestamp 1731220645
transform 1 0 1152 0 1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5391_6
timestamp 1731220645
transform 1 0 1080 0 1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5390_6
timestamp 1731220645
transform 1 0 1016 0 1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5389_6
timestamp 1731220645
transform 1 0 992 0 -1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5388_6
timestamp 1731220645
transform 1 0 920 0 -1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5387_6
timestamp 1731220645
transform 1 0 1064 0 -1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5386_6
timestamp 1731220645
transform 1 0 1136 0 -1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5385_6
timestamp 1731220645
transform 1 0 1184 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5384_6
timestamp 1731220645
transform 1 0 1184 0 -1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5383_6
timestamp 1731220645
transform 1 0 1296 0 -1 960
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5382_6
timestamp 1731220645
transform 1 0 1344 0 -1 960
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5381_6
timestamp 1731220645
transform 1 0 1424 0 -1 960
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5380_6
timestamp 1731220645
transform 1 0 1504 0 -1 960
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5379_6
timestamp 1731220645
transform 1 0 1600 0 1 824
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5378_6
timestamp 1731220645
transform 1 0 1552 0 1 824
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5377_6
timestamp 1731220645
transform 1 0 1512 0 1 824
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5376_6
timestamp 1731220645
transform 1 0 1472 0 1 824
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5375_6
timestamp 1731220645
transform 1 0 1432 0 1 824
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5374_6
timestamp 1731220645
transform 1 0 1528 0 -1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5373_6
timestamp 1731220645
transform 1 0 1464 0 -1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5372_6
timestamp 1731220645
transform 1 0 1408 0 -1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5371_6
timestamp 1731220645
transform 1 0 1352 0 -1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5370_6
timestamp 1731220645
transform 1 0 1568 0 1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5369_6
timestamp 1731220645
transform 1 0 1480 0 1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5368_6
timestamp 1731220645
transform 1 0 1400 0 1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5367_6
timestamp 1731220645
transform 1 0 1336 0 1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5366_6
timestamp 1731220645
transform 1 0 1296 0 1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5365_6
timestamp 1731220645
transform 1 0 1296 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5364_6
timestamp 1731220645
transform 1 0 1184 0 -1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5363_6
timestamp 1731220645
transform 1 0 1144 0 -1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5362_6
timestamp 1731220645
transform 1 0 1088 0 -1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5361_6
timestamp 1731220645
transform 1 0 1032 0 -1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5360_6
timestamp 1731220645
transform 1 0 976 0 -1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5359_6
timestamp 1731220645
transform 1 0 912 0 -1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5358_6
timestamp 1731220645
transform 1 0 848 0 -1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5357_6
timestamp 1731220645
transform 1 0 1184 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5356_6
timestamp 1731220645
transform 1 0 1128 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5355_6
timestamp 1731220645
transform 1 0 1072 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5354_6
timestamp 1731220645
transform 1 0 1016 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5353_6
timestamp 1731220645
transform 1 0 968 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5352_6
timestamp 1731220645
transform 1 0 912 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5351_6
timestamp 1731220645
transform 1 0 848 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5350_6
timestamp 1731220645
transform 1 0 776 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5349_6
timestamp 1731220645
transform 1 0 1016 0 -1 524
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5348_6
timestamp 1731220645
transform 1 0 952 0 -1 524
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5347_6
timestamp 1731220645
transform 1 0 896 0 -1 524
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5346_6
timestamp 1731220645
transform 1 0 840 0 -1 524
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5345_6
timestamp 1731220645
transform 1 0 776 0 -1 524
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5344_6
timestamp 1731220645
transform 1 0 712 0 -1 524
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5343_6
timestamp 1731220645
transform 1 0 640 0 -1 524
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5342_6
timestamp 1731220645
transform 1 0 880 0 1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5341_6
timestamp 1731220645
transform 1 0 824 0 1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5340_6
timestamp 1731220645
transform 1 0 768 0 1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5339_6
timestamp 1731220645
transform 1 0 712 0 1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5338_6
timestamp 1731220645
transform 1 0 664 0 1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5337_6
timestamp 1731220645
transform 1 0 608 0 1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5336_6
timestamp 1731220645
transform 1 0 552 0 1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5335_6
timestamp 1731220645
transform 1 0 768 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5334_6
timestamp 1731220645
transform 1 0 720 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5333_6
timestamp 1731220645
transform 1 0 672 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5332_6
timestamp 1731220645
transform 1 0 624 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5331_6
timestamp 1731220645
transform 1 0 576 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5330_6
timestamp 1731220645
transform 1 0 528 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5329_6
timestamp 1731220645
transform 1 0 480 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5328_6
timestamp 1731220645
transform 1 0 584 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5327_6
timestamp 1731220645
transform 1 0 624 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5326_6
timestamp 1731220645
transform 1 0 672 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5325_6
timestamp 1731220645
transform 1 0 720 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5324_6
timestamp 1731220645
transform 1 0 768 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5323_6
timestamp 1731220645
transform 1 0 912 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5322_6
timestamp 1731220645
transform 1 0 864 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5321_6
timestamp 1731220645
transform 1 0 816 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5320_6
timestamp 1731220645
transform 1 0 784 0 -1 240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5319_6
timestamp 1731220645
transform 1 0 720 0 -1 240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5318_6
timestamp 1731220645
transform 1 0 648 0 -1 240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5317_6
timestamp 1731220645
transform 1 0 840 0 -1 240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5316_6
timestamp 1731220645
transform 1 0 1016 0 -1 240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5315_6
timestamp 1731220645
transform 1 0 952 0 -1 240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5314_6
timestamp 1731220645
transform 1 0 896 0 -1 240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5313_6
timestamp 1731220645
transform 1 0 720 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5312_6
timestamp 1731220645
transform 1 0 672 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5311_6
timestamp 1731220645
transform 1 0 624 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5310_6
timestamp 1731220645
transform 1 0 760 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5309_6
timestamp 1731220645
transform 1 0 800 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5308_6
timestamp 1731220645
transform 1 0 840 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5307_6
timestamp 1731220645
transform 1 0 880 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5306_6
timestamp 1731220645
transform 1 0 920 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5305_6
timestamp 1731220645
transform 1 0 968 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5304_6
timestamp 1731220645
transform 1 0 1016 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5303_6
timestamp 1731220645
transform 1 0 1064 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5302_6
timestamp 1731220645
transform 1 0 1104 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5301_6
timestamp 1731220645
transform 1 0 1144 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5300_6
timestamp 1731220645
transform 1 0 1184 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5299_6
timestamp 1731220645
transform 1 0 1296 0 1 92
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5298_6
timestamp 1731220645
transform 1 0 1336 0 1 92
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5297_6
timestamp 1731220645
transform 1 0 1376 0 1 92
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5296_6
timestamp 1731220645
transform 1 0 1416 0 1 92
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5295_6
timestamp 1731220645
transform 1 0 1456 0 1 92
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5294_6
timestamp 1731220645
transform 1 0 1640 0 1 92
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5293_6
timestamp 1731220645
transform 1 0 1576 0 1 92
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5292_6
timestamp 1731220645
transform 1 0 1512 0 1 92
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5291_6
timestamp 1731220645
transform 1 0 1440 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5290_6
timestamp 1731220645
transform 1 0 1400 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5289_6
timestamp 1731220645
transform 1 0 1360 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5288_6
timestamp 1731220645
transform 1 0 1488 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5287_6
timestamp 1731220645
transform 1 0 1544 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5286_6
timestamp 1731220645
transform 1 0 1600 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5285_6
timestamp 1731220645
transform 1 0 1664 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5284_6
timestamp 1731220645
transform 1 0 1736 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5283_6
timestamp 1731220645
transform 1 0 1688 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5282_6
timestamp 1731220645
transform 1 0 1648 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5281_6
timestamp 1731220645
transform 1 0 1608 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5280_6
timestamp 1731220645
transform 1 0 1568 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5279_6
timestamp 1731220645
transform 1 0 1528 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5278_6
timestamp 1731220645
transform 1 0 1488 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5277_6
timestamp 1731220645
transform 1 0 1584 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5276_6
timestamp 1731220645
transform 1 0 1528 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5275_6
timestamp 1731220645
transform 1 0 1480 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5274_6
timestamp 1731220645
transform 1 0 1440 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5273_6
timestamp 1731220645
transform 1 0 1520 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5272_6
timestamp 1731220645
transform 1 0 1456 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5271_6
timestamp 1731220645
transform 1 0 1392 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5270_6
timestamp 1731220645
transform 1 0 1336 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5269_6
timestamp 1731220645
transform 1 0 1296 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5268_6
timestamp 1731220645
transform 1 0 1296 0 -1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5267_6
timestamp 1731220645
transform 1 0 1184 0 -1 524
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5266_6
timestamp 1731220645
transform 1 0 1144 0 -1 524
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5265_6
timestamp 1731220645
transform 1 0 1080 0 -1 524
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5264_6
timestamp 1731220645
transform 1 0 1368 0 -1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5263_6
timestamp 1731220645
transform 1 0 1472 0 -1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5262_6
timestamp 1731220645
transform 1 0 1576 0 -1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5261_6
timestamp 1731220645
transform 1 0 1488 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5260_6
timestamp 1731220645
transform 1 0 1448 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5259_6
timestamp 1731220645
transform 1 0 1408 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5258_6
timestamp 1731220645
transform 1 0 1536 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5257_6
timestamp 1731220645
transform 1 0 1720 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5256_6
timestamp 1731220645
transform 1 0 1656 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5255_6
timestamp 1731220645
transform 1 0 1592 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5254_6
timestamp 1731220645
transform 1 0 1504 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5253_6
timestamp 1731220645
transform 1 0 1392 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5252_6
timestamp 1731220645
transform 1 0 1616 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5251_6
timestamp 1731220645
transform 1 0 1720 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5250_6
timestamp 1731220645
transform 1 0 1744 0 1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5249_6
timestamp 1731220645
transform 1 0 1656 0 1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5248_6
timestamp 1731220645
transform 1 0 1640 0 -1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5247_6
timestamp 1731220645
transform 1 0 1584 0 -1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5246_6
timestamp 1731220645
transform 1 0 1696 0 -1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5245_6
timestamp 1731220645
transform 1 0 1704 0 1 824
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5244_6
timestamp 1731220645
transform 1 0 1648 0 1 824
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5243_6
timestamp 1731220645
transform 1 0 1584 0 -1 960
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5242_6
timestamp 1731220645
transform 1 0 1672 0 -1 960
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5241_6
timestamp 1731220645
transform 1 0 1768 0 1 968
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5240_6
timestamp 1731220645
transform 1 0 1728 0 1 968
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5239_6
timestamp 1731220645
transform 1 0 1688 0 1 968
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5238_6
timestamp 1731220645
transform 1 0 1648 0 1 968
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5237_6
timestamp 1731220645
transform 1 0 1608 0 1 968
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5236_6
timestamp 1731220645
transform 1 0 1568 0 1 968
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5235_6
timestamp 1731220645
transform 1 0 1720 0 -1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5234_6
timestamp 1731220645
transform 1 0 1664 0 -1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5233_6
timestamp 1731220645
transform 1 0 1608 0 -1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5232_6
timestamp 1731220645
transform 1 0 1552 0 -1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5231_6
timestamp 1731220645
transform 1 0 1504 0 -1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5230_6
timestamp 1731220645
transform 1 0 1464 0 -1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5229_6
timestamp 1731220645
transform 1 0 1424 0 -1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5228_6
timestamp 1731220645
transform 1 0 1792 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5227_6
timestamp 1731220645
transform 1 0 1680 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5226_6
timestamp 1731220645
transform 1 0 1576 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5225_6
timestamp 1731220645
transform 1 0 1480 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5224_6
timestamp 1731220645
transform 1 0 1400 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5223_6
timestamp 1731220645
transform 1 0 1336 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5222_6
timestamp 1731220645
transform 1 0 1296 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5221_6
timestamp 1731220645
transform 1 0 1296 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5220_6
timestamp 1731220645
transform 1 0 1368 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5219_6
timestamp 1731220645
transform 1 0 1472 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5218_6
timestamp 1731220645
transform 1 0 1680 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5217_6
timestamp 1731220645
transform 1 0 1576 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5216_6
timestamp 1731220645
transform 1 0 1536 0 1 1248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5215_6
timestamp 1731220645
transform 1 0 1496 0 1 1248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5214_6
timestamp 1731220645
transform 1 0 1456 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5213_6
timestamp 1731220645
transform 1 0 1392 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5212_6
timestamp 1731220645
transform 1 0 1336 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5211_6
timestamp 1731220645
transform 1 0 1368 0 1 1392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5210_6
timestamp 1731220645
transform 1 0 1456 0 1 1392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5209_6
timestamp 1731220645
transform 1 0 1496 0 -1 1528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5208_6
timestamp 1731220645
transform 1 0 1408 0 -1 1528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5207_6
timestamp 1731220645
transform 1 0 1328 0 -1 1528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5206_6
timestamp 1731220645
transform 1 0 1320 0 1 1532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5205_6
timestamp 1731220645
transform 1 0 1392 0 1 1532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5204_6
timestamp 1731220645
transform 1 0 1440 0 -1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5203_6
timestamp 1731220645
transform 1 0 1352 0 -1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5202_6
timestamp 1731220645
transform 1 0 1296 0 -1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5201_6
timestamp 1731220645
transform 1 0 1344 0 1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5200_6
timestamp 1731220645
transform 1 0 1296 0 1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5199_6
timestamp 1731220645
transform 1 0 1184 0 1 1712
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5198_6
timestamp 1731220645
transform 1 0 1144 0 1 1712
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5197_6
timestamp 1731220645
transform 1 0 1080 0 1 1712
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5196_6
timestamp 1731220645
transform 1 0 1024 0 1 1712
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5195_6
timestamp 1731220645
transform 1 0 1184 0 -1 1848
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5194_6
timestamp 1731220645
transform 1 0 1128 0 -1 1848
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5193_6
timestamp 1731220645
transform 1 0 1056 0 -1 1848
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5192_6
timestamp 1731220645
transform 1 0 984 0 -1 1848
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5191_6
timestamp 1731220645
transform 1 0 904 0 -1 1848
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5190_6
timestamp 1731220645
transform 1 0 1112 0 1 1856
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5189_6
timestamp 1731220645
transform 1 0 1032 0 1 1856
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5188_6
timestamp 1731220645
transform 1 0 952 0 1 1856
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5187_6
timestamp 1731220645
transform 1 0 872 0 1 1856
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5186_6
timestamp 1731220645
transform 1 0 1056 0 -1 1996
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5185_6
timestamp 1731220645
transform 1 0 992 0 -1 1996
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5184_6
timestamp 1731220645
transform 1 0 928 0 -1 1996
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5183_6
timestamp 1731220645
transform 1 0 864 0 -1 1996
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5182_6
timestamp 1731220645
transform 1 0 952 0 1 2004
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5181_6
timestamp 1731220645
transform 1 0 1008 0 1 2004
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5180_6
timestamp 1731220645
transform 1 0 1064 0 1 2004
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5179_6
timestamp 1731220645
transform 1 0 1136 0 -1 2140
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5178_6
timestamp 1731220645
transform 1 0 1072 0 -1 2140
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5177_6
timestamp 1731220645
transform 1 0 1016 0 -1 2140
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5176_6
timestamp 1731220645
transform 1 0 960 0 -1 2140
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5175_6
timestamp 1731220645
transform 1 0 904 0 -1 2140
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5174_6
timestamp 1731220645
transform 1 0 848 0 -1 2140
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5173_6
timestamp 1731220645
transform 1 0 896 0 1 2004
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5172_6
timestamp 1731220645
transform 1 0 840 0 1 2004
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5171_6
timestamp 1731220645
transform 1 0 792 0 1 2004
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5170_6
timestamp 1731220645
transform 1 0 752 0 -1 1996
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5169_6
timestamp 1731220645
transform 1 0 688 0 -1 1996
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5168_6
timestamp 1731220645
transform 1 0 808 0 -1 1996
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5167_6
timestamp 1731220645
transform 1 0 792 0 1 1856
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5166_6
timestamp 1731220645
transform 1 0 712 0 1 1856
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5165_6
timestamp 1731220645
transform 1 0 632 0 1 1856
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5164_6
timestamp 1731220645
transform 1 0 624 0 -1 1848
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5163_6
timestamp 1731220645
transform 1 0 720 0 -1 1848
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5162_6
timestamp 1731220645
transform 1 0 816 0 -1 1848
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5161_6
timestamp 1731220645
transform 1 0 744 0 1 1712
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5160_6
timestamp 1731220645
transform 1 0 656 0 1 1712
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5159_6
timestamp 1731220645
transform 1 0 824 0 1 1712
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5158_6
timestamp 1731220645
transform 1 0 896 0 1 1712
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5157_6
timestamp 1731220645
transform 1 0 960 0 1 1712
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5156_6
timestamp 1731220645
transform 1 0 1152 0 -1 1708
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5155_6
timestamp 1731220645
transform 1 0 1080 0 -1 1708
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5154_6
timestamp 1731220645
transform 1 0 1008 0 -1 1708
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5153_6
timestamp 1731220645
transform 1 0 944 0 -1 1708
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5152_6
timestamp 1731220645
transform 1 0 872 0 -1 1708
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5151_6
timestamp 1731220645
transform 1 0 792 0 -1 1708
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5150_6
timestamp 1731220645
transform 1 0 704 0 -1 1708
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5149_6
timestamp 1731220645
transform 1 0 992 0 1 1568
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5148_6
timestamp 1731220645
transform 1 0 936 0 1 1568
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5147_6
timestamp 1731220645
transform 1 0 880 0 1 1568
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5146_6
timestamp 1731220645
transform 1 0 824 0 1 1568
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5145_6
timestamp 1731220645
transform 1 0 768 0 1 1568
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5144_6
timestamp 1731220645
transform 1 0 712 0 1 1568
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5143_6
timestamp 1731220645
transform 1 0 656 0 1 1568
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5142_6
timestamp 1731220645
transform 1 0 920 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5141_6
timestamp 1731220645
transform 1 0 880 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5140_6
timestamp 1731220645
transform 1 0 840 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5139_6
timestamp 1731220645
transform 1 0 800 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5138_6
timestamp 1731220645
transform 1 0 760 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5137_6
timestamp 1731220645
transform 1 0 720 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5136_6
timestamp 1731220645
transform 1 0 680 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5135_6
timestamp 1731220645
transform 1 0 640 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5134_6
timestamp 1731220645
transform 1 0 600 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5133_6
timestamp 1731220645
transform 1 0 560 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5132_6
timestamp 1731220645
transform 1 0 520 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5131_6
timestamp 1731220645
transform 1 0 480 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5130_6
timestamp 1731220645
transform 1 0 440 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5129_6
timestamp 1731220645
transform 1 0 400 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5128_6
timestamp 1731220645
transform 1 0 360 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5127_6
timestamp 1731220645
transform 1 0 320 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5126_6
timestamp 1731220645
transform 1 0 592 0 1 1568
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5125_6
timestamp 1731220645
transform 1 0 528 0 1 1568
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5124_6
timestamp 1731220645
transform 1 0 464 0 1 1568
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5123_6
timestamp 1731220645
transform 1 0 408 0 1 1568
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5122_6
timestamp 1731220645
transform 1 0 352 0 1 1568
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5121_6
timestamp 1731220645
transform 1 0 304 0 1 1568
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5120_6
timestamp 1731220645
transform 1 0 264 0 1 1568
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5119_6
timestamp 1731220645
transform 1 0 608 0 -1 1708
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5118_6
timestamp 1731220645
transform 1 0 504 0 -1 1708
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5117_6
timestamp 1731220645
transform 1 0 408 0 -1 1708
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5116_6
timestamp 1731220645
transform 1 0 312 0 -1 1708
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5115_6
timestamp 1731220645
transform 1 0 232 0 -1 1708
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5114_6
timestamp 1731220645
transform 1 0 168 0 -1 1708
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5113_6
timestamp 1731220645
transform 1 0 128 0 -1 1708
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5112_6
timestamp 1731220645
transform 1 0 560 0 1 1712
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5111_6
timestamp 1731220645
transform 1 0 464 0 1 1712
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5110_6
timestamp 1731220645
transform 1 0 368 0 1 1712
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5109_6
timestamp 1731220645
transform 1 0 280 0 1 1712
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5108_6
timestamp 1731220645
transform 1 0 208 0 1 1712
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5107_6
timestamp 1731220645
transform 1 0 168 0 1 1712
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5106_6
timestamp 1731220645
transform 1 0 128 0 1 1712
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5105_6
timestamp 1731220645
transform 1 0 128 0 -1 1848
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5104_6
timestamp 1731220645
transform 1 0 168 0 -1 1848
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5103_6
timestamp 1731220645
transform 1 0 208 0 -1 1848
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5102_6
timestamp 1731220645
transform 1 0 264 0 -1 1848
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5101_6
timestamp 1731220645
transform 1 0 528 0 -1 1848
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5100_6
timestamp 1731220645
transform 1 0 432 0 -1 1848
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_599_6
timestamp 1731220645
transform 1 0 344 0 -1 1848
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_598_6
timestamp 1731220645
transform 1 0 256 0 1 1856
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_597_6
timestamp 1731220645
transform 1 0 208 0 1 1856
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_596_6
timestamp 1731220645
transform 1 0 168 0 1 1856
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_595_6
timestamp 1731220645
transform 1 0 312 0 1 1856
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_594_6
timestamp 1731220645
transform 1 0 384 0 1 1856
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_593_6
timestamp 1731220645
transform 1 0 544 0 1 1856
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_592_6
timestamp 1731220645
transform 1 0 464 0 1 1856
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_591_6
timestamp 1731220645
transform 1 0 448 0 -1 1996
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_590_6
timestamp 1731220645
transform 1 0 400 0 -1 1996
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_589_6
timestamp 1731220645
transform 1 0 360 0 -1 1996
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_588_6
timestamp 1731220645
transform 1 0 504 0 -1 1996
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_587_6
timestamp 1731220645
transform 1 0 560 0 -1 1996
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_586_6
timestamp 1731220645
transform 1 0 624 0 -1 1996
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_585_6
timestamp 1731220645
transform 1 0 680 0 1 2004
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_584_6
timestamp 1731220645
transform 1 0 736 0 1 2004
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_583_6
timestamp 1731220645
transform 1 0 720 0 -1 2140
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_582_6
timestamp 1731220645
transform 1 0 784 0 -1 2140
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_581_6
timestamp 1731220645
transform 1 0 776 0 1 2148
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_580_6
timestamp 1731220645
transform 1 0 712 0 1 2148
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_579_6
timestamp 1731220645
transform 1 0 904 0 1 2148
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_578_6
timestamp 1731220645
transform 1 0 840 0 1 2148
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_577_6
timestamp 1731220645
transform 1 0 824 0 -1 2284
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_576_6
timestamp 1731220645
transform 1 0 904 0 -1 2284
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_575_6
timestamp 1731220645
transform 1 0 984 0 -1 2284
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_574_6
timestamp 1731220645
transform 1 0 1024 0 1 2288
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_573_6
timestamp 1731220645
transform 1 0 952 0 1 2288
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_572_6
timestamp 1731220645
transform 1 0 880 0 1 2288
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_571_6
timestamp 1731220645
transform 1 0 816 0 1 2288
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_570_6
timestamp 1731220645
transform 1 0 1040 0 -1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_569_6
timestamp 1731220645
transform 1 0 984 0 -1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_568_6
timestamp 1731220645
transform 1 0 928 0 -1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_567_6
timestamp 1731220645
transform 1 0 880 0 -1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_566_6
timestamp 1731220645
transform 1 0 832 0 -1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_565_6
timestamp 1731220645
transform 1 0 920 0 1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_564_6
timestamp 1731220645
transform 1 0 824 0 1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_563_6
timestamp 1731220645
transform 1 0 736 0 1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_562_6
timestamp 1731220645
transform 1 0 648 0 1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_561_6
timestamp 1731220645
transform 1 0 784 0 -1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_560_6
timestamp 1731220645
transform 1 0 728 0 -1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_559_6
timestamp 1731220645
transform 1 0 672 0 -1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_558_6
timestamp 1731220645
transform 1 0 608 0 -1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_557_6
timestamp 1731220645
transform 1 0 536 0 -1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_556_6
timestamp 1731220645
transform 1 0 592 0 1 2288
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_555_6
timestamp 1731220645
transform 1 0 672 0 1 2288
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_554_6
timestamp 1731220645
transform 1 0 744 0 1 2288
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_553_6
timestamp 1731220645
transform 1 0 752 0 -1 2284
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_552_6
timestamp 1731220645
transform 1 0 680 0 -1 2284
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_551_6
timestamp 1731220645
transform 1 0 608 0 -1 2284
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_550_6
timestamp 1731220645
transform 1 0 528 0 -1 2284
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_549_6
timestamp 1731220645
transform 1 0 656 0 1 2148
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_548_6
timestamp 1731220645
transform 1 0 600 0 1 2148
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_547_6
timestamp 1731220645
transform 1 0 544 0 1 2148
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_546_6
timestamp 1731220645
transform 1 0 544 0 -1 2140
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_545_6
timestamp 1731220645
transform 1 0 600 0 -1 2140
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_544_6
timestamp 1731220645
transform 1 0 656 0 -1 2140
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_543_6
timestamp 1731220645
transform 1 0 624 0 1 2004
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_542_6
timestamp 1731220645
transform 1 0 576 0 1 2004
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_541_6
timestamp 1731220645
transform 1 0 536 0 1 2004
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_540_6
timestamp 1731220645
transform 1 0 496 0 1 2004
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_539_6
timestamp 1731220645
transform 1 0 456 0 1 2004
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_538_6
timestamp 1731220645
transform 1 0 416 0 1 2004
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_537_6
timestamp 1731220645
transform 1 0 376 0 1 2004
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_536_6
timestamp 1731220645
transform 1 0 496 0 -1 2140
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_535_6
timestamp 1731220645
transform 1 0 456 0 -1 2140
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_534_6
timestamp 1731220645
transform 1 0 416 0 -1 2140
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_533_6
timestamp 1731220645
transform 1 0 376 0 -1 2140
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_532_6
timestamp 1731220645
transform 1 0 488 0 1 2148
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_531_6
timestamp 1731220645
transform 1 0 424 0 1 2148
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_530_6
timestamp 1731220645
transform 1 0 368 0 1 2148
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_529_6
timestamp 1731220645
transform 1 0 320 0 1 2148
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_528_6
timestamp 1731220645
transform 1 0 280 0 1 2148
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_527_6
timestamp 1731220645
transform 1 0 240 0 1 2148
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_526_6
timestamp 1731220645
transform 1 0 448 0 -1 2284
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_525_6
timestamp 1731220645
transform 1 0 368 0 -1 2284
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_524_6
timestamp 1731220645
transform 1 0 296 0 -1 2284
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_523_6
timestamp 1731220645
transform 1 0 224 0 -1 2284
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_522_6
timestamp 1731220645
transform 1 0 168 0 -1 2284
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_521_6
timestamp 1731220645
transform 1 0 128 0 -1 2284
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_520_6
timestamp 1731220645
transform 1 0 264 0 1 2288
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_519_6
timestamp 1731220645
transform 1 0 208 0 1 2288
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_518_6
timestamp 1731220645
transform 1 0 168 0 1 2288
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_517_6
timestamp 1731220645
transform 1 0 128 0 1 2288
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_516_6
timestamp 1731220645
transform 1 0 344 0 1 2288
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_515_6
timestamp 1731220645
transform 1 0 424 0 1 2288
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_514_6
timestamp 1731220645
transform 1 0 512 0 1 2288
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_513_6
timestamp 1731220645
transform 1 0 464 0 -1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_512_6
timestamp 1731220645
transform 1 0 384 0 -1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_511_6
timestamp 1731220645
transform 1 0 312 0 -1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_510_6
timestamp 1731220645
transform 1 0 240 0 -1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_59_6
timestamp 1731220645
transform 1 0 176 0 -1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_58_6
timestamp 1731220645
transform 1 0 128 0 -1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_57_6
timestamp 1731220645
transform 1 0 560 0 1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_56_6
timestamp 1731220645
transform 1 0 472 0 1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_55_6
timestamp 1731220645
transform 1 0 384 0 1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_54_6
timestamp 1731220645
transform 1 0 304 0 1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_53_6
timestamp 1731220645
transform 1 0 248 0 1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_52_6
timestamp 1731220645
transform 1 0 208 0 1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_51_6
timestamp 1731220645
transform 1 0 168 0 1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_50_6
timestamp 1731220645
transform 1 0 128 0 1 2432
box 4 6 36 64
<< end >>
