magic
tech sky130l
timestamp 1730767243
<< m1 >>
rect 688 1383 692 1455
rect 808 1251 812 1283
rect 912 651 916 675
rect 696 523 700 555
rect 1120 255 1124 323
<< m2c >>
rect 256 1635 260 1639
rect 344 1635 348 1639
rect 111 1621 115 1625
rect 1567 1621 1571 1625
rect 111 1603 115 1607
rect 1567 1603 1571 1607
rect 111 1569 115 1573
rect 1567 1569 1571 1573
rect 111 1551 115 1555
rect 1567 1551 1571 1555
rect 216 1535 220 1539
rect 304 1535 308 1539
rect 392 1535 396 1539
rect 384 1503 388 1507
rect 472 1499 476 1503
rect 560 1499 564 1503
rect 648 1499 652 1503
rect 111 1485 115 1489
rect 1567 1485 1571 1489
rect 111 1467 115 1471
rect 1567 1467 1571 1471
rect 688 1455 692 1459
rect 111 1413 115 1417
rect 111 1395 115 1399
rect 1567 1413 1571 1417
rect 968 1407 972 1411
rect 1567 1395 1571 1399
rect 688 1379 692 1383
rect 696 1379 700 1383
rect 784 1379 788 1383
rect 872 1379 876 1383
rect 960 1379 964 1383
rect 848 1343 852 1347
rect 968 1339 972 1343
rect 1088 1339 1092 1343
rect 1208 1339 1212 1343
rect 1328 1339 1332 1343
rect 1448 1339 1452 1343
rect 111 1325 115 1329
rect 1567 1325 1571 1329
rect 111 1307 115 1311
rect 1567 1307 1571 1311
rect 808 1283 812 1287
rect 111 1273 115 1277
rect 111 1255 115 1259
rect 1567 1273 1571 1277
rect 1080 1267 1084 1271
rect 1567 1255 1571 1259
rect 808 1247 812 1251
rect 576 1239 580 1243
rect 728 1239 732 1243
rect 896 1239 900 1243
rect 1072 1239 1076 1243
rect 1248 1239 1252 1243
rect 1432 1239 1436 1243
rect 928 1195 932 1199
rect 232 1191 236 1195
rect 448 1191 452 1195
rect 680 1191 684 1195
rect 1184 1191 1188 1195
rect 1448 1193 1452 1197
rect 111 1177 115 1181
rect 1567 1177 1571 1181
rect 111 1159 115 1163
rect 1567 1159 1571 1163
rect 111 1117 115 1121
rect 1567 1117 1571 1121
rect 111 1099 115 1103
rect 1567 1099 1571 1103
rect 168 1083 172 1087
rect 592 1083 596 1087
rect 1024 1083 1028 1087
rect 1456 1085 1460 1089
rect 272 1055 276 1059
rect 1064 1055 1068 1059
rect 1464 1055 1468 1059
rect 664 1051 668 1055
rect 111 1037 115 1041
rect 1567 1037 1571 1041
rect 111 1019 115 1023
rect 1567 1019 1571 1023
rect 111 985 115 989
rect 1567 985 1571 989
rect 111 967 115 971
rect 1567 967 1571 971
rect 448 951 452 955
rect 696 951 700 955
rect 952 951 956 955
rect 1208 951 1212 955
rect 1472 949 1476 953
rect 576 911 580 915
rect 1472 911 1476 915
rect 784 907 788 911
rect 1008 907 1012 911
rect 1240 907 1244 911
rect 111 893 115 897
rect 1567 893 1571 897
rect 111 875 115 879
rect 1567 875 1571 879
rect 111 833 115 837
rect 1567 833 1571 837
rect 968 827 972 831
rect 1128 827 1132 831
rect 111 815 115 819
rect 1567 815 1571 819
rect 808 799 812 803
rect 960 799 964 803
rect 1120 799 1124 803
rect 1288 799 1292 803
rect 1456 799 1460 803
rect 888 759 892 763
rect 1408 759 1412 763
rect 1008 755 1012 759
rect 1136 755 1140 759
rect 1272 755 1276 759
rect 111 741 115 745
rect 1567 741 1571 745
rect 111 723 115 727
rect 1567 723 1571 727
rect 111 681 115 685
rect 1567 681 1571 685
rect 912 675 916 679
rect 976 675 980 679
rect 1176 675 1180 679
rect 1384 675 1388 679
rect 111 663 115 667
rect 1567 663 1571 667
rect 768 647 772 651
rect 912 647 916 651
rect 968 647 972 651
rect 1168 647 1172 651
rect 1376 647 1380 651
rect 880 623 884 627
rect 1360 623 1364 627
rect 640 619 644 623
rect 1120 619 1124 623
rect 111 605 115 609
rect 1567 605 1571 609
rect 111 587 115 591
rect 1567 587 1571 591
rect 696 555 700 559
rect 111 545 115 549
rect 111 527 115 531
rect 1567 545 1571 549
rect 1567 527 1571 531
rect 696 519 700 523
rect 392 511 396 515
rect 624 511 628 515
rect 864 511 868 515
rect 1112 511 1116 515
rect 1360 511 1364 515
rect 768 471 772 475
rect 1376 471 1380 475
rect 184 467 188 471
rect 472 467 476 471
rect 1072 467 1076 471
rect 111 453 115 457
rect 1567 453 1571 457
rect 111 435 115 439
rect 1567 435 1571 439
rect 111 389 115 393
rect 1567 389 1571 393
rect 111 371 115 375
rect 1567 371 1571 375
rect 208 355 212 359
rect 600 355 604 359
rect 1000 355 1004 359
rect 1400 355 1404 359
rect 832 327 836 331
rect 1432 327 1436 331
rect 264 323 268 327
rect 544 323 548 327
rect 1120 323 1124 327
rect 1128 323 1132 327
rect 111 309 115 313
rect 111 291 115 295
rect 1567 309 1571 313
rect 1567 291 1571 295
rect 1120 251 1124 255
rect 111 241 115 245
rect 1567 241 1571 245
rect 704 235 708 239
rect 1208 235 1212 239
rect 111 223 115 227
rect 1567 223 1571 227
rect 456 207 460 211
rect 696 207 700 211
rect 944 207 948 211
rect 1200 207 1204 211
rect 1464 207 1468 211
rect 544 167 548 171
rect 1504 167 1508 171
rect 648 163 652 167
rect 760 163 764 167
rect 888 163 892 167
rect 1032 163 1036 167
rect 1192 163 1196 167
rect 1360 163 1364 167
rect 111 149 115 153
rect 1567 149 1571 153
rect 111 131 115 135
rect 1567 131 1571 135
<< m2 >>
rect 134 1642 140 1643
rect 134 1638 135 1642
rect 139 1638 140 1642
rect 134 1637 140 1638
rect 222 1642 228 1643
rect 222 1638 223 1642
rect 227 1638 228 1642
rect 310 1642 316 1643
rect 255 1639 261 1640
rect 255 1638 256 1639
rect 222 1637 228 1638
rect 248 1636 256 1638
rect 210 1631 216 1632
rect 210 1627 211 1631
rect 215 1630 216 1631
rect 248 1630 250 1636
rect 255 1635 256 1636
rect 260 1635 261 1639
rect 310 1638 311 1642
rect 315 1638 316 1642
rect 343 1639 349 1640
rect 343 1638 344 1639
rect 310 1637 316 1638
rect 255 1634 261 1635
rect 336 1636 344 1638
rect 215 1628 250 1630
rect 298 1631 304 1632
rect 215 1627 216 1628
rect 210 1626 216 1627
rect 298 1627 299 1631
rect 303 1630 304 1631
rect 336 1630 338 1636
rect 343 1635 344 1636
rect 348 1635 349 1639
rect 343 1634 349 1635
rect 303 1628 338 1630
rect 303 1627 304 1628
rect 298 1626 304 1627
rect 110 1625 116 1626
rect 110 1621 111 1625
rect 115 1621 116 1625
rect 110 1620 116 1621
rect 1566 1625 1572 1626
rect 1566 1621 1567 1625
rect 1571 1621 1572 1625
rect 1566 1620 1572 1621
rect 110 1607 116 1608
rect 110 1603 111 1607
rect 115 1603 116 1607
rect 110 1602 116 1603
rect 1566 1607 1572 1608
rect 1566 1603 1567 1607
rect 1571 1603 1572 1607
rect 1566 1602 1572 1603
rect 134 1596 140 1597
rect 222 1596 228 1597
rect 310 1596 316 1597
rect 134 1592 135 1596
rect 139 1592 140 1596
rect 210 1595 216 1596
rect 210 1594 211 1595
rect 205 1592 211 1594
rect 134 1591 140 1592
rect 210 1591 211 1592
rect 215 1591 216 1595
rect 222 1592 223 1596
rect 227 1592 228 1596
rect 298 1595 304 1596
rect 298 1594 299 1595
rect 293 1592 299 1594
rect 222 1591 228 1592
rect 298 1591 299 1592
rect 303 1591 304 1595
rect 310 1592 311 1596
rect 315 1592 316 1596
rect 310 1591 316 1592
rect 326 1595 332 1596
rect 326 1591 327 1595
rect 331 1594 332 1595
rect 331 1592 345 1594
rect 331 1591 332 1592
rect 210 1590 216 1591
rect 298 1590 304 1591
rect 326 1590 332 1591
rect 182 1584 188 1585
rect 270 1584 276 1585
rect 358 1584 364 1585
rect 182 1580 183 1584
rect 187 1580 188 1584
rect 258 1583 264 1584
rect 258 1582 259 1583
rect 253 1580 259 1582
rect 182 1579 188 1580
rect 258 1579 259 1580
rect 263 1579 264 1583
rect 270 1580 271 1584
rect 275 1580 276 1584
rect 346 1583 352 1584
rect 346 1582 347 1583
rect 341 1580 347 1582
rect 270 1579 276 1580
rect 346 1579 347 1580
rect 351 1579 352 1583
rect 358 1580 359 1584
rect 363 1580 364 1584
rect 358 1579 364 1580
rect 382 1583 388 1584
rect 382 1579 383 1583
rect 387 1582 388 1583
rect 387 1580 393 1582
rect 387 1579 388 1580
rect 258 1578 264 1579
rect 346 1578 352 1579
rect 382 1578 388 1579
rect 110 1573 116 1574
rect 110 1569 111 1573
rect 115 1569 116 1573
rect 110 1568 116 1569
rect 1566 1573 1572 1574
rect 1566 1569 1567 1573
rect 1571 1569 1572 1573
rect 1566 1568 1572 1569
rect 110 1555 116 1556
rect 110 1551 111 1555
rect 115 1551 116 1555
rect 110 1550 116 1551
rect 1566 1555 1572 1556
rect 1566 1551 1567 1555
rect 1571 1551 1572 1555
rect 1566 1550 1572 1551
rect 258 1547 264 1548
rect 258 1543 259 1547
rect 263 1546 264 1547
rect 346 1547 352 1548
rect 263 1544 298 1546
rect 263 1543 264 1544
rect 258 1542 264 1543
rect 215 1539 221 1540
rect 182 1538 188 1539
rect 182 1534 183 1538
rect 187 1534 188 1538
rect 215 1535 216 1539
rect 220 1538 221 1539
rect 270 1538 276 1539
rect 220 1536 266 1538
rect 220 1535 221 1536
rect 215 1534 221 1535
rect 182 1533 188 1534
rect 264 1530 266 1536
rect 270 1534 271 1538
rect 275 1534 276 1538
rect 296 1538 298 1544
rect 346 1543 347 1547
rect 351 1546 352 1547
rect 351 1544 386 1546
rect 351 1543 352 1544
rect 346 1542 352 1543
rect 303 1539 309 1540
rect 303 1538 304 1539
rect 296 1536 304 1538
rect 303 1535 304 1536
rect 308 1535 309 1539
rect 303 1534 309 1535
rect 358 1538 364 1539
rect 358 1534 359 1538
rect 363 1534 364 1538
rect 384 1538 386 1544
rect 391 1539 397 1540
rect 391 1538 392 1539
rect 384 1536 392 1538
rect 391 1535 392 1536
rect 396 1535 397 1539
rect 391 1534 397 1535
rect 270 1533 276 1534
rect 358 1533 364 1534
rect 326 1531 332 1532
rect 326 1530 327 1531
rect 264 1528 327 1530
rect 326 1527 327 1528
rect 331 1527 332 1531
rect 326 1526 332 1527
rect 382 1507 389 1508
rect 350 1506 356 1507
rect 350 1502 351 1506
rect 355 1502 356 1506
rect 382 1503 383 1507
rect 388 1503 389 1507
rect 382 1502 389 1503
rect 438 1506 444 1507
rect 438 1502 439 1506
rect 443 1502 444 1506
rect 526 1506 532 1507
rect 471 1503 477 1504
rect 471 1502 472 1503
rect 350 1501 356 1502
rect 438 1501 444 1502
rect 464 1500 472 1502
rect 426 1495 432 1496
rect 426 1491 427 1495
rect 431 1494 432 1495
rect 464 1494 466 1500
rect 471 1499 472 1500
rect 476 1499 477 1503
rect 526 1502 527 1506
rect 531 1502 532 1506
rect 614 1506 620 1507
rect 559 1503 565 1504
rect 559 1502 560 1503
rect 526 1501 532 1502
rect 471 1498 477 1499
rect 552 1500 560 1502
rect 431 1492 466 1494
rect 514 1495 520 1496
rect 431 1491 432 1492
rect 426 1490 432 1491
rect 514 1491 515 1495
rect 519 1494 520 1495
rect 552 1494 554 1500
rect 559 1499 560 1500
rect 564 1499 565 1503
rect 614 1502 615 1506
rect 619 1502 620 1506
rect 647 1503 653 1504
rect 647 1502 648 1503
rect 614 1501 620 1502
rect 559 1498 565 1499
rect 640 1500 648 1502
rect 519 1492 554 1494
rect 602 1495 608 1496
rect 519 1491 520 1492
rect 514 1490 520 1491
rect 602 1491 603 1495
rect 607 1494 608 1495
rect 640 1494 642 1500
rect 647 1499 648 1500
rect 652 1499 653 1503
rect 647 1498 653 1499
rect 607 1492 642 1494
rect 607 1491 608 1492
rect 602 1490 608 1491
rect 110 1489 116 1490
rect 110 1485 111 1489
rect 115 1485 116 1489
rect 110 1484 116 1485
rect 1566 1489 1572 1490
rect 1566 1485 1567 1489
rect 1571 1485 1572 1489
rect 1566 1484 1572 1485
rect 110 1471 116 1472
rect 110 1467 111 1471
rect 115 1467 116 1471
rect 110 1466 116 1467
rect 1566 1471 1572 1472
rect 1566 1467 1567 1471
rect 1571 1467 1572 1471
rect 1566 1466 1572 1467
rect 350 1460 356 1461
rect 438 1460 444 1461
rect 526 1460 532 1461
rect 614 1460 620 1461
rect 350 1456 351 1460
rect 355 1456 356 1460
rect 426 1459 432 1460
rect 426 1458 427 1459
rect 421 1456 427 1458
rect 350 1455 356 1456
rect 426 1455 427 1456
rect 431 1455 432 1459
rect 438 1456 439 1460
rect 443 1456 444 1460
rect 514 1459 520 1460
rect 514 1458 515 1459
rect 509 1456 515 1458
rect 438 1455 444 1456
rect 514 1455 515 1456
rect 519 1455 520 1459
rect 526 1456 527 1460
rect 531 1456 532 1460
rect 602 1459 608 1460
rect 602 1458 603 1459
rect 597 1456 603 1458
rect 526 1455 532 1456
rect 602 1455 603 1456
rect 607 1455 608 1459
rect 614 1456 615 1460
rect 619 1456 620 1460
rect 687 1459 693 1460
rect 687 1458 688 1459
rect 685 1456 688 1458
rect 614 1455 620 1456
rect 687 1455 688 1456
rect 692 1455 693 1459
rect 426 1454 432 1455
rect 514 1454 520 1455
rect 602 1454 608 1455
rect 687 1454 693 1455
rect 662 1428 668 1429
rect 750 1428 756 1429
rect 838 1428 844 1429
rect 926 1428 932 1429
rect 662 1424 663 1428
rect 667 1424 668 1428
rect 738 1427 744 1428
rect 738 1426 739 1427
rect 733 1424 739 1426
rect 662 1423 668 1424
rect 738 1423 739 1424
rect 743 1423 744 1427
rect 750 1424 751 1428
rect 755 1424 756 1428
rect 826 1427 832 1428
rect 826 1426 827 1427
rect 821 1424 827 1426
rect 750 1423 756 1424
rect 826 1423 827 1424
rect 831 1423 832 1427
rect 838 1424 839 1428
rect 843 1424 844 1428
rect 914 1427 920 1428
rect 914 1426 915 1427
rect 909 1424 915 1426
rect 838 1423 844 1424
rect 914 1423 915 1424
rect 919 1423 920 1427
rect 926 1424 927 1428
rect 931 1424 932 1428
rect 926 1423 932 1424
rect 738 1422 744 1423
rect 826 1422 832 1423
rect 914 1422 920 1423
rect 110 1417 116 1418
rect 110 1413 111 1417
rect 115 1413 116 1417
rect 110 1412 116 1413
rect 1566 1417 1572 1418
rect 1566 1413 1567 1417
rect 1571 1413 1572 1417
rect 1566 1412 1572 1413
rect 850 1411 856 1412
rect 850 1407 851 1411
rect 855 1410 856 1411
rect 967 1411 973 1412
rect 967 1410 968 1411
rect 855 1408 968 1410
rect 855 1407 856 1408
rect 850 1406 856 1407
rect 967 1407 968 1408
rect 972 1407 973 1411
rect 967 1406 973 1407
rect 110 1399 116 1400
rect 110 1395 111 1399
rect 115 1395 116 1399
rect 110 1394 116 1395
rect 1566 1399 1572 1400
rect 1566 1395 1567 1399
rect 1571 1395 1572 1399
rect 1566 1394 1572 1395
rect 738 1391 744 1392
rect 738 1387 739 1391
rect 743 1390 744 1391
rect 826 1391 832 1392
rect 743 1388 778 1390
rect 743 1387 744 1388
rect 738 1386 744 1387
rect 687 1383 693 1384
rect 662 1382 668 1383
rect 662 1378 663 1382
rect 667 1378 668 1382
rect 687 1379 688 1383
rect 692 1382 693 1383
rect 695 1383 701 1384
rect 695 1382 696 1383
rect 692 1380 696 1382
rect 692 1379 693 1380
rect 687 1378 693 1379
rect 695 1379 696 1380
rect 700 1379 701 1383
rect 695 1378 701 1379
rect 750 1382 756 1383
rect 750 1378 751 1382
rect 755 1378 756 1382
rect 776 1382 778 1388
rect 826 1387 827 1391
rect 831 1390 832 1391
rect 914 1391 920 1392
rect 831 1388 866 1390
rect 831 1387 832 1388
rect 826 1386 832 1387
rect 783 1383 789 1384
rect 783 1382 784 1383
rect 776 1380 784 1382
rect 783 1379 784 1380
rect 788 1379 789 1383
rect 783 1378 789 1379
rect 838 1382 844 1383
rect 838 1378 839 1382
rect 843 1378 844 1382
rect 864 1382 866 1388
rect 914 1387 915 1391
rect 919 1390 920 1391
rect 919 1388 954 1390
rect 919 1387 920 1388
rect 914 1386 920 1387
rect 871 1383 877 1384
rect 871 1382 872 1383
rect 864 1380 872 1382
rect 871 1379 872 1380
rect 876 1379 877 1383
rect 871 1378 877 1379
rect 926 1382 932 1383
rect 926 1378 927 1382
rect 931 1378 932 1382
rect 952 1382 954 1388
rect 959 1383 965 1384
rect 959 1382 960 1383
rect 952 1380 960 1382
rect 959 1379 960 1380
rect 964 1379 965 1383
rect 959 1378 965 1379
rect 662 1377 668 1378
rect 750 1377 756 1378
rect 838 1377 844 1378
rect 926 1377 932 1378
rect 847 1347 856 1348
rect 814 1346 820 1347
rect 814 1342 815 1346
rect 819 1342 820 1346
rect 847 1343 848 1347
rect 855 1343 856 1347
rect 847 1342 856 1343
rect 934 1346 940 1347
rect 934 1342 935 1346
rect 939 1342 940 1346
rect 1054 1346 1060 1347
rect 967 1343 973 1344
rect 967 1342 968 1343
rect 814 1341 820 1342
rect 934 1341 940 1342
rect 960 1340 968 1342
rect 906 1335 912 1336
rect 906 1331 907 1335
rect 911 1334 912 1335
rect 960 1334 962 1340
rect 967 1339 968 1340
rect 972 1339 973 1343
rect 1054 1342 1055 1346
rect 1059 1342 1060 1346
rect 1174 1346 1180 1347
rect 1087 1343 1093 1344
rect 1087 1342 1088 1343
rect 1054 1341 1060 1342
rect 967 1338 973 1339
rect 1080 1340 1088 1342
rect 911 1332 962 1334
rect 1026 1335 1032 1336
rect 911 1331 912 1332
rect 906 1330 912 1331
rect 1026 1331 1027 1335
rect 1031 1334 1032 1335
rect 1080 1334 1082 1340
rect 1087 1339 1088 1340
rect 1092 1339 1093 1343
rect 1174 1342 1175 1346
rect 1179 1342 1180 1346
rect 1294 1346 1300 1347
rect 1174 1341 1180 1342
rect 1207 1343 1213 1344
rect 1087 1338 1093 1339
rect 1207 1339 1208 1343
rect 1212 1342 1213 1343
rect 1246 1343 1252 1344
rect 1246 1342 1247 1343
rect 1212 1340 1247 1342
rect 1212 1339 1213 1340
rect 1207 1338 1213 1339
rect 1246 1339 1247 1340
rect 1251 1339 1252 1343
rect 1294 1342 1295 1346
rect 1299 1342 1300 1346
rect 1414 1346 1420 1347
rect 1327 1343 1333 1344
rect 1327 1342 1328 1343
rect 1294 1341 1300 1342
rect 1246 1338 1252 1339
rect 1320 1340 1328 1342
rect 1031 1332 1082 1334
rect 1266 1335 1272 1336
rect 1031 1331 1032 1332
rect 1026 1330 1032 1331
rect 1266 1331 1267 1335
rect 1271 1334 1272 1335
rect 1320 1334 1322 1340
rect 1327 1339 1328 1340
rect 1332 1339 1333 1343
rect 1414 1342 1415 1346
rect 1419 1342 1420 1346
rect 1447 1343 1453 1344
rect 1447 1342 1448 1343
rect 1414 1341 1420 1342
rect 1327 1338 1333 1339
rect 1440 1340 1448 1342
rect 1271 1332 1322 1334
rect 1386 1335 1392 1336
rect 1271 1331 1272 1332
rect 1266 1330 1272 1331
rect 1386 1331 1387 1335
rect 1391 1334 1392 1335
rect 1440 1334 1442 1340
rect 1447 1339 1448 1340
rect 1452 1339 1453 1343
rect 1447 1338 1453 1339
rect 1391 1332 1442 1334
rect 1391 1331 1392 1332
rect 1386 1330 1392 1331
rect 110 1329 116 1330
rect 110 1325 111 1329
rect 115 1325 116 1329
rect 110 1324 116 1325
rect 1566 1329 1572 1330
rect 1566 1325 1567 1329
rect 1571 1325 1572 1329
rect 1566 1324 1572 1325
rect 110 1311 116 1312
rect 110 1307 111 1311
rect 115 1307 116 1311
rect 110 1306 116 1307
rect 1566 1311 1572 1312
rect 1566 1307 1567 1311
rect 1571 1307 1572 1311
rect 1566 1306 1572 1307
rect 814 1300 820 1301
rect 934 1300 940 1301
rect 1054 1300 1060 1301
rect 1174 1300 1180 1301
rect 1294 1300 1300 1301
rect 1414 1300 1420 1301
rect 814 1296 815 1300
rect 819 1296 820 1300
rect 906 1299 912 1300
rect 906 1298 907 1299
rect 885 1296 907 1298
rect 814 1295 820 1296
rect 906 1295 907 1296
rect 911 1295 912 1299
rect 934 1296 935 1300
rect 939 1296 940 1300
rect 1026 1299 1032 1300
rect 1026 1298 1027 1299
rect 1005 1296 1027 1298
rect 934 1295 940 1296
rect 1026 1295 1027 1296
rect 1031 1295 1032 1299
rect 1054 1296 1055 1300
rect 1059 1296 1060 1300
rect 1054 1295 1060 1296
rect 1086 1299 1092 1300
rect 1086 1295 1087 1299
rect 1091 1295 1092 1299
rect 1174 1296 1175 1300
rect 1179 1296 1180 1300
rect 1266 1299 1272 1300
rect 1266 1298 1267 1299
rect 1245 1296 1267 1298
rect 1174 1295 1180 1296
rect 1266 1295 1267 1296
rect 1271 1295 1272 1299
rect 1294 1296 1295 1300
rect 1299 1296 1300 1300
rect 1386 1299 1392 1300
rect 1386 1298 1387 1299
rect 1365 1296 1387 1298
rect 1294 1295 1300 1296
rect 1386 1295 1387 1296
rect 1391 1295 1392 1299
rect 1414 1296 1415 1300
rect 1419 1296 1420 1300
rect 1414 1295 1420 1296
rect 1446 1299 1452 1300
rect 1446 1295 1447 1299
rect 1451 1295 1452 1299
rect 906 1294 912 1295
rect 1026 1294 1032 1295
rect 1086 1294 1092 1295
rect 1266 1294 1272 1295
rect 1386 1294 1392 1295
rect 1446 1294 1452 1295
rect 542 1288 548 1289
rect 694 1288 700 1289
rect 862 1288 868 1289
rect 1038 1288 1044 1289
rect 542 1284 543 1288
rect 547 1284 548 1288
rect 626 1287 632 1288
rect 626 1286 627 1287
rect 613 1284 627 1286
rect 542 1283 548 1284
rect 626 1283 627 1284
rect 631 1283 632 1287
rect 694 1284 695 1288
rect 699 1284 700 1288
rect 807 1287 813 1288
rect 807 1286 808 1287
rect 765 1284 808 1286
rect 694 1283 700 1284
rect 807 1283 808 1284
rect 812 1283 813 1287
rect 862 1284 863 1288
rect 867 1284 868 1288
rect 862 1283 868 1284
rect 926 1287 932 1288
rect 926 1283 927 1287
rect 931 1283 932 1287
rect 1038 1284 1039 1288
rect 1043 1284 1044 1288
rect 1038 1283 1044 1284
rect 1214 1288 1220 1289
rect 1398 1288 1404 1289
rect 1214 1284 1215 1288
rect 1219 1284 1220 1288
rect 1214 1283 1220 1284
rect 1246 1287 1252 1288
rect 1246 1283 1247 1287
rect 1251 1283 1252 1287
rect 1398 1284 1399 1288
rect 1403 1284 1404 1288
rect 1398 1283 1404 1284
rect 1438 1287 1444 1288
rect 1438 1283 1439 1287
rect 1443 1283 1444 1287
rect 626 1282 632 1283
rect 807 1282 813 1283
rect 926 1282 932 1283
rect 1246 1282 1252 1283
rect 1438 1282 1444 1283
rect 110 1277 116 1278
rect 110 1273 111 1277
rect 115 1273 116 1277
rect 110 1272 116 1273
rect 1566 1277 1572 1278
rect 1566 1273 1567 1277
rect 1571 1273 1572 1277
rect 1566 1272 1572 1273
rect 686 1271 692 1272
rect 686 1267 687 1271
rect 691 1270 692 1271
rect 1079 1271 1085 1272
rect 1079 1270 1080 1271
rect 691 1268 1080 1270
rect 691 1267 692 1268
rect 686 1266 692 1267
rect 1079 1267 1080 1268
rect 1084 1267 1085 1271
rect 1079 1266 1085 1267
rect 110 1259 116 1260
rect 110 1255 111 1259
rect 115 1255 116 1259
rect 110 1254 116 1255
rect 1566 1259 1572 1260
rect 1566 1255 1567 1259
rect 1571 1255 1572 1259
rect 1566 1254 1572 1255
rect 626 1251 632 1252
rect 626 1247 627 1251
rect 631 1250 632 1251
rect 807 1251 813 1252
rect 631 1248 722 1250
rect 631 1247 632 1248
rect 626 1246 632 1247
rect 575 1243 581 1244
rect 542 1242 548 1243
rect 542 1238 543 1242
rect 547 1238 548 1242
rect 575 1239 576 1243
rect 580 1242 581 1243
rect 686 1243 692 1244
rect 686 1242 687 1243
rect 580 1240 687 1242
rect 580 1239 581 1240
rect 575 1238 581 1239
rect 686 1239 687 1240
rect 691 1239 692 1243
rect 686 1238 692 1239
rect 694 1242 700 1243
rect 694 1238 695 1242
rect 699 1238 700 1242
rect 720 1242 722 1248
rect 807 1247 808 1251
rect 812 1250 813 1251
rect 812 1248 890 1250
rect 812 1247 813 1248
rect 807 1246 813 1247
rect 727 1243 733 1244
rect 727 1242 728 1243
rect 720 1240 728 1242
rect 727 1239 728 1240
rect 732 1239 733 1243
rect 727 1238 733 1239
rect 862 1242 868 1243
rect 862 1238 863 1242
rect 867 1238 868 1242
rect 888 1242 890 1248
rect 895 1243 901 1244
rect 1071 1243 1077 1244
rect 895 1242 896 1243
rect 888 1240 896 1242
rect 895 1239 896 1240
rect 900 1239 901 1243
rect 895 1238 901 1239
rect 1038 1242 1044 1243
rect 1038 1238 1039 1242
rect 1043 1238 1044 1242
rect 1071 1239 1072 1243
rect 1076 1242 1077 1243
rect 1086 1243 1092 1244
rect 1238 1243 1244 1244
rect 1086 1242 1087 1243
rect 1076 1240 1087 1242
rect 1076 1239 1077 1240
rect 1071 1238 1077 1239
rect 1086 1239 1087 1240
rect 1091 1239 1092 1243
rect 1086 1238 1092 1239
rect 1214 1242 1220 1243
rect 1214 1238 1215 1242
rect 1219 1238 1220 1242
rect 1238 1239 1239 1243
rect 1243 1242 1244 1243
rect 1247 1243 1253 1244
rect 1431 1243 1437 1244
rect 1247 1242 1248 1243
rect 1243 1240 1248 1242
rect 1243 1239 1244 1240
rect 1238 1238 1244 1239
rect 1247 1239 1248 1240
rect 1252 1239 1253 1243
rect 1247 1238 1253 1239
rect 1398 1242 1404 1243
rect 1398 1238 1399 1242
rect 1403 1238 1404 1242
rect 1431 1239 1432 1243
rect 1436 1242 1437 1243
rect 1446 1243 1452 1244
rect 1446 1242 1447 1243
rect 1436 1240 1447 1242
rect 1436 1239 1437 1240
rect 1431 1238 1437 1239
rect 1446 1239 1447 1240
rect 1451 1239 1452 1243
rect 1446 1238 1452 1239
rect 542 1237 548 1238
rect 694 1237 700 1238
rect 862 1237 868 1238
rect 1038 1237 1044 1238
rect 1214 1237 1220 1238
rect 1398 1237 1404 1238
rect 926 1199 933 1200
rect 1438 1199 1444 1200
rect 198 1198 204 1199
rect 198 1194 199 1198
rect 203 1194 204 1198
rect 414 1198 420 1199
rect 198 1193 204 1194
rect 231 1195 237 1196
rect 231 1191 232 1195
rect 236 1194 237 1195
rect 414 1194 415 1198
rect 419 1194 420 1198
rect 646 1198 652 1199
rect 236 1192 282 1194
rect 414 1193 420 1194
rect 447 1195 453 1196
rect 236 1191 237 1192
rect 231 1190 237 1191
rect 280 1186 282 1192
rect 447 1191 448 1195
rect 452 1194 453 1195
rect 646 1194 647 1198
rect 651 1194 652 1198
rect 894 1198 900 1199
rect 452 1192 638 1194
rect 646 1193 652 1194
rect 679 1195 685 1196
rect 452 1191 453 1192
rect 447 1190 453 1191
rect 430 1187 436 1188
rect 430 1186 431 1187
rect 280 1184 431 1186
rect 430 1183 431 1184
rect 435 1183 436 1187
rect 636 1186 638 1192
rect 679 1191 680 1195
rect 684 1194 685 1195
rect 894 1194 895 1198
rect 899 1194 900 1198
rect 926 1195 927 1199
rect 932 1195 933 1199
rect 926 1194 933 1195
rect 1150 1198 1156 1199
rect 1150 1194 1151 1198
rect 1155 1194 1156 1198
rect 1414 1198 1420 1199
rect 684 1192 806 1194
rect 894 1193 900 1194
rect 1150 1193 1156 1194
rect 1183 1195 1189 1196
rect 684 1191 685 1192
rect 679 1190 685 1191
rect 662 1187 668 1188
rect 662 1186 663 1187
rect 636 1184 663 1186
rect 430 1182 436 1183
rect 662 1183 663 1184
rect 667 1183 668 1187
rect 804 1186 806 1192
rect 1183 1191 1184 1195
rect 1188 1194 1189 1195
rect 1206 1195 1212 1196
rect 1206 1194 1207 1195
rect 1188 1192 1207 1194
rect 1188 1191 1189 1192
rect 1183 1190 1189 1191
rect 1206 1191 1207 1192
rect 1211 1191 1212 1195
rect 1414 1194 1415 1198
rect 1419 1194 1420 1198
rect 1438 1195 1439 1199
rect 1443 1198 1444 1199
rect 1443 1197 1453 1198
rect 1443 1196 1448 1197
rect 1443 1195 1444 1196
rect 1438 1194 1444 1195
rect 1414 1193 1420 1194
rect 1447 1193 1448 1196
rect 1452 1193 1453 1197
rect 1447 1192 1453 1193
rect 1206 1190 1212 1191
rect 910 1187 916 1188
rect 910 1186 911 1187
rect 804 1184 911 1186
rect 662 1182 668 1183
rect 910 1183 911 1184
rect 915 1183 916 1187
rect 910 1182 916 1183
rect 110 1181 116 1182
rect 110 1177 111 1181
rect 115 1177 116 1181
rect 110 1176 116 1177
rect 1566 1181 1572 1182
rect 1566 1177 1567 1181
rect 1571 1177 1572 1181
rect 1566 1176 1572 1177
rect 110 1163 116 1164
rect 110 1159 111 1163
rect 115 1159 116 1163
rect 110 1158 116 1159
rect 1566 1163 1572 1164
rect 1566 1159 1567 1163
rect 1571 1159 1572 1163
rect 1566 1158 1572 1159
rect 198 1152 204 1153
rect 414 1152 420 1153
rect 646 1152 652 1153
rect 894 1152 900 1153
rect 1150 1152 1156 1153
rect 1414 1152 1420 1153
rect 198 1148 199 1152
rect 203 1148 204 1152
rect 198 1147 204 1148
rect 230 1151 236 1152
rect 230 1147 231 1151
rect 235 1147 236 1151
rect 414 1148 415 1152
rect 419 1148 420 1152
rect 414 1147 420 1148
rect 430 1151 436 1152
rect 430 1147 431 1151
rect 435 1150 436 1151
rect 435 1148 449 1150
rect 646 1148 647 1152
rect 651 1148 652 1152
rect 435 1147 436 1148
rect 646 1147 652 1148
rect 662 1151 668 1152
rect 662 1147 663 1151
rect 667 1150 668 1151
rect 667 1148 681 1150
rect 894 1148 895 1152
rect 899 1148 900 1152
rect 667 1147 668 1148
rect 894 1147 900 1148
rect 910 1151 916 1152
rect 910 1147 911 1151
rect 915 1150 916 1151
rect 915 1148 929 1150
rect 1150 1148 1151 1152
rect 1155 1148 1156 1152
rect 1238 1151 1244 1152
rect 1238 1150 1239 1151
rect 1221 1148 1239 1150
rect 915 1147 916 1148
rect 1150 1147 1156 1148
rect 1238 1147 1239 1148
rect 1243 1147 1244 1151
rect 1414 1148 1415 1152
rect 1419 1148 1420 1152
rect 1414 1147 1420 1148
rect 1446 1151 1452 1152
rect 1446 1147 1447 1151
rect 1451 1147 1452 1151
rect 230 1146 236 1147
rect 430 1146 436 1147
rect 662 1146 668 1147
rect 910 1146 916 1147
rect 1238 1146 1244 1147
rect 1446 1146 1452 1147
rect 134 1132 140 1133
rect 558 1132 564 1133
rect 990 1132 996 1133
rect 1422 1132 1428 1133
rect 134 1128 135 1132
rect 139 1128 140 1132
rect 378 1131 384 1132
rect 378 1130 379 1131
rect 205 1128 379 1130
rect 134 1127 140 1128
rect 378 1127 379 1128
rect 383 1127 384 1131
rect 558 1128 559 1132
rect 563 1128 564 1132
rect 750 1131 756 1132
rect 750 1130 751 1131
rect 629 1128 751 1130
rect 558 1127 564 1128
rect 750 1127 751 1128
rect 755 1127 756 1131
rect 990 1128 991 1132
rect 995 1128 996 1132
rect 990 1127 996 1128
rect 1058 1131 1064 1132
rect 1058 1127 1059 1131
rect 1063 1127 1064 1131
rect 1422 1128 1423 1132
rect 1427 1128 1428 1132
rect 1422 1127 1428 1128
rect 1462 1131 1468 1132
rect 1462 1127 1463 1131
rect 1467 1127 1468 1131
rect 378 1126 384 1127
rect 750 1126 756 1127
rect 1058 1126 1064 1127
rect 1462 1126 1468 1127
rect 110 1121 116 1122
rect 110 1117 111 1121
rect 115 1117 116 1121
rect 110 1116 116 1117
rect 1566 1121 1572 1122
rect 1566 1117 1567 1121
rect 1571 1117 1572 1121
rect 1566 1116 1572 1117
rect 110 1103 116 1104
rect 110 1099 111 1103
rect 115 1099 116 1103
rect 110 1098 116 1099
rect 1566 1103 1572 1104
rect 1566 1099 1567 1103
rect 1571 1099 1572 1103
rect 1566 1098 1572 1099
rect 378 1095 384 1096
rect 378 1091 379 1095
rect 383 1094 384 1095
rect 750 1095 756 1096
rect 383 1092 586 1094
rect 383 1091 384 1092
rect 378 1090 384 1091
rect 167 1087 173 1088
rect 134 1086 140 1087
rect 134 1082 135 1086
rect 139 1082 140 1086
rect 167 1083 168 1087
rect 172 1086 173 1087
rect 230 1087 236 1088
rect 230 1086 231 1087
rect 172 1084 231 1086
rect 172 1083 173 1084
rect 167 1082 173 1083
rect 230 1083 231 1084
rect 235 1083 236 1087
rect 230 1082 236 1083
rect 558 1086 564 1087
rect 558 1082 559 1086
rect 563 1082 564 1086
rect 584 1086 586 1092
rect 618 1091 624 1092
rect 591 1087 597 1088
rect 591 1086 592 1087
rect 584 1084 592 1086
rect 591 1083 592 1084
rect 596 1083 597 1087
rect 618 1087 619 1091
rect 623 1090 624 1091
rect 750 1091 751 1095
rect 755 1094 756 1095
rect 755 1092 1018 1094
rect 755 1091 756 1092
rect 750 1090 756 1091
rect 623 1088 681 1090
rect 623 1087 624 1088
rect 618 1086 624 1087
rect 591 1082 597 1083
rect 134 1081 140 1082
rect 558 1081 564 1082
rect 679 1078 681 1088
rect 990 1086 996 1087
rect 990 1082 991 1086
rect 995 1082 996 1086
rect 1016 1086 1018 1092
rect 1446 1091 1452 1092
rect 1023 1087 1029 1088
rect 1446 1087 1447 1091
rect 1451 1090 1452 1091
rect 1451 1089 1461 1090
rect 1451 1088 1456 1089
rect 1451 1087 1452 1088
rect 1023 1086 1024 1087
rect 1016 1084 1024 1086
rect 1023 1083 1024 1084
rect 1028 1083 1029 1087
rect 1023 1082 1029 1083
rect 1422 1086 1428 1087
rect 1446 1086 1452 1087
rect 1422 1082 1423 1086
rect 1427 1082 1428 1086
rect 1455 1085 1456 1088
rect 1460 1085 1461 1089
rect 1455 1084 1461 1085
rect 990 1081 996 1082
rect 1422 1081 1428 1082
rect 1046 1079 1052 1080
rect 1046 1078 1047 1079
rect 679 1076 1047 1078
rect 1046 1075 1047 1076
rect 1051 1075 1052 1079
rect 1046 1074 1052 1075
rect 271 1059 277 1060
rect 238 1058 244 1059
rect 238 1054 239 1058
rect 243 1054 244 1058
rect 271 1055 272 1059
rect 276 1058 277 1059
rect 618 1059 624 1060
rect 1058 1059 1069 1060
rect 1462 1059 1469 1060
rect 618 1058 619 1059
rect 276 1056 619 1058
rect 276 1055 277 1056
rect 271 1054 277 1055
rect 618 1055 619 1056
rect 623 1055 624 1059
rect 618 1054 624 1055
rect 630 1058 636 1059
rect 630 1054 631 1058
rect 635 1054 636 1058
rect 1030 1058 1036 1059
rect 663 1055 669 1056
rect 663 1054 664 1055
rect 238 1053 244 1054
rect 630 1053 636 1054
rect 656 1052 664 1054
rect 498 1047 504 1048
rect 498 1043 499 1047
rect 503 1046 504 1047
rect 656 1046 658 1052
rect 663 1051 664 1052
rect 668 1051 669 1055
rect 1030 1054 1031 1058
rect 1035 1054 1036 1058
rect 1058 1055 1059 1059
rect 1063 1055 1064 1059
rect 1068 1055 1069 1059
rect 1058 1054 1069 1055
rect 1430 1058 1436 1059
rect 1430 1054 1431 1058
rect 1435 1054 1436 1058
rect 1462 1055 1463 1059
rect 1468 1055 1469 1059
rect 1462 1054 1469 1055
rect 1030 1053 1036 1054
rect 1430 1053 1436 1054
rect 663 1050 669 1051
rect 503 1044 658 1046
rect 503 1043 504 1044
rect 498 1042 504 1043
rect 110 1041 116 1042
rect 110 1037 111 1041
rect 115 1037 116 1041
rect 110 1036 116 1037
rect 1566 1041 1572 1042
rect 1566 1037 1567 1041
rect 1571 1037 1572 1041
rect 1566 1036 1572 1037
rect 110 1023 116 1024
rect 110 1019 111 1023
rect 115 1019 116 1023
rect 110 1018 116 1019
rect 1566 1023 1572 1024
rect 1566 1019 1567 1023
rect 1571 1019 1572 1023
rect 1566 1018 1572 1019
rect 238 1012 244 1013
rect 630 1012 636 1013
rect 1030 1012 1036 1013
rect 1430 1012 1436 1013
rect 238 1008 239 1012
rect 243 1008 244 1012
rect 498 1011 504 1012
rect 498 1010 499 1011
rect 309 1008 499 1010
rect 238 1007 244 1008
rect 498 1007 499 1008
rect 503 1007 504 1011
rect 630 1008 631 1012
rect 635 1008 636 1012
rect 630 1007 636 1008
rect 686 1011 692 1012
rect 686 1007 687 1011
rect 691 1007 692 1011
rect 1030 1008 1031 1012
rect 1035 1008 1036 1012
rect 1030 1007 1036 1008
rect 1046 1011 1052 1012
rect 1046 1007 1047 1011
rect 1051 1010 1052 1011
rect 1051 1008 1065 1010
rect 1430 1008 1431 1012
rect 1435 1008 1436 1012
rect 1051 1007 1052 1008
rect 1430 1007 1436 1008
rect 1462 1011 1468 1012
rect 1462 1007 1463 1011
rect 1467 1007 1468 1011
rect 498 1006 504 1007
rect 686 1006 692 1007
rect 1046 1006 1052 1007
rect 1462 1006 1468 1007
rect 414 1000 420 1001
rect 662 1000 668 1001
rect 918 1000 924 1001
rect 1174 1000 1180 1001
rect 1438 1000 1444 1001
rect 414 996 415 1000
rect 419 996 420 1000
rect 566 999 572 1000
rect 566 998 567 999
rect 485 996 567 998
rect 414 995 420 996
rect 566 995 567 996
rect 571 995 572 999
rect 662 996 663 1000
rect 667 996 668 1000
rect 822 999 828 1000
rect 822 998 823 999
rect 733 996 823 998
rect 662 995 668 996
rect 822 995 823 996
rect 827 995 828 999
rect 918 996 919 1000
rect 923 996 924 1000
rect 918 995 924 996
rect 950 999 956 1000
rect 950 995 951 999
rect 955 995 956 999
rect 1174 996 1175 1000
rect 1179 996 1180 1000
rect 1174 995 1180 996
rect 1206 999 1212 1000
rect 1206 995 1207 999
rect 1211 995 1212 999
rect 1438 996 1439 1000
rect 1443 996 1444 1000
rect 1438 995 1444 996
rect 1470 999 1476 1000
rect 1470 995 1471 999
rect 1475 995 1476 999
rect 566 994 572 995
rect 822 994 828 995
rect 950 994 956 995
rect 1206 994 1212 995
rect 1470 994 1476 995
rect 110 989 116 990
rect 110 985 111 989
rect 115 985 116 989
rect 110 984 116 985
rect 1566 989 1572 990
rect 1566 985 1567 989
rect 1571 985 1572 989
rect 1566 984 1572 985
rect 110 971 116 972
rect 110 967 111 971
rect 115 967 116 971
rect 110 966 116 967
rect 1566 971 1572 972
rect 1566 967 1567 971
rect 1571 967 1572 971
rect 1566 966 1572 967
rect 822 963 828 964
rect 822 959 823 963
rect 827 962 828 963
rect 827 960 946 962
rect 827 959 828 960
rect 822 958 828 959
rect 447 955 453 956
rect 686 955 692 956
rect 414 954 420 955
rect 414 950 415 954
rect 419 950 420 954
rect 447 951 448 955
rect 452 954 453 955
rect 662 954 668 955
rect 452 952 598 954
rect 452 951 453 952
rect 447 950 453 951
rect 414 949 420 950
rect 596 946 598 952
rect 662 950 663 954
rect 667 950 668 954
rect 686 951 687 955
rect 691 954 692 955
rect 695 955 701 956
rect 695 954 696 955
rect 691 952 696 954
rect 691 951 692 952
rect 686 950 692 951
rect 695 951 696 952
rect 700 951 701 955
rect 695 950 701 951
rect 918 954 924 955
rect 918 950 919 954
rect 923 950 924 954
rect 944 954 946 960
rect 951 955 957 956
rect 1207 955 1213 956
rect 951 954 952 955
rect 944 952 952 954
rect 951 951 952 952
rect 956 951 957 955
rect 951 950 957 951
rect 1174 954 1180 955
rect 1174 950 1175 954
rect 1179 950 1180 954
rect 1207 951 1208 955
rect 1212 954 1213 955
rect 1286 955 1292 956
rect 1462 955 1468 956
rect 1286 954 1287 955
rect 1212 952 1287 954
rect 1212 951 1213 952
rect 1207 950 1213 951
rect 1286 951 1287 952
rect 1291 951 1292 955
rect 1286 950 1292 951
rect 1438 954 1444 955
rect 1438 950 1439 954
rect 1443 950 1444 954
rect 1462 951 1463 955
rect 1467 954 1468 955
rect 1467 953 1477 954
rect 1467 952 1472 953
rect 1467 951 1468 952
rect 1462 950 1468 951
rect 662 949 668 950
rect 918 949 924 950
rect 1174 949 1180 950
rect 1438 949 1444 950
rect 1471 949 1472 952
rect 1476 949 1477 953
rect 1471 948 1477 949
rect 950 947 956 948
rect 950 946 951 947
rect 596 944 951 946
rect 950 943 951 944
rect 955 943 956 947
rect 950 942 956 943
rect 566 915 572 916
rect 542 914 548 915
rect 542 910 543 914
rect 547 910 548 914
rect 566 911 567 915
rect 571 914 572 915
rect 575 915 581 916
rect 1470 915 1477 916
rect 575 914 576 915
rect 571 912 576 914
rect 571 911 572 912
rect 566 910 572 911
rect 575 911 576 912
rect 580 911 581 915
rect 575 910 581 911
rect 750 914 756 915
rect 750 910 751 914
rect 755 910 756 914
rect 974 914 980 915
rect 783 911 789 912
rect 783 910 784 911
rect 542 909 548 910
rect 750 909 756 910
rect 776 908 784 910
rect 690 903 696 904
rect 690 899 691 903
rect 695 902 696 903
rect 776 902 778 908
rect 783 907 784 908
rect 788 907 789 911
rect 974 910 975 914
rect 979 910 980 914
rect 1206 914 1212 915
rect 1007 911 1013 912
rect 1007 910 1008 911
rect 974 909 980 910
rect 783 906 789 907
rect 1000 908 1008 910
rect 695 900 778 902
rect 894 903 900 904
rect 695 899 696 900
rect 690 898 696 899
rect 894 899 895 903
rect 899 902 900 903
rect 1000 902 1002 908
rect 1007 907 1008 908
rect 1012 907 1013 911
rect 1206 910 1207 914
rect 1211 910 1212 914
rect 1438 914 1444 915
rect 1239 911 1245 912
rect 1239 910 1240 911
rect 1206 909 1212 910
rect 1007 906 1013 907
rect 1232 908 1240 910
rect 899 900 1002 902
rect 1122 903 1128 904
rect 899 899 900 900
rect 894 898 900 899
rect 1122 899 1123 903
rect 1127 902 1128 903
rect 1232 902 1234 908
rect 1239 907 1240 908
rect 1244 907 1245 911
rect 1438 910 1439 914
rect 1443 910 1444 914
rect 1470 911 1471 915
rect 1476 911 1477 915
rect 1470 910 1477 911
rect 1438 909 1444 910
rect 1239 906 1245 907
rect 1127 900 1234 902
rect 1127 899 1128 900
rect 1122 898 1128 899
rect 110 897 116 898
rect 110 893 111 897
rect 115 893 116 897
rect 110 892 116 893
rect 1566 897 1572 898
rect 1566 893 1567 897
rect 1571 893 1572 897
rect 1566 892 1572 893
rect 110 879 116 880
rect 110 875 111 879
rect 115 875 116 879
rect 110 874 116 875
rect 1566 879 1572 880
rect 1566 875 1567 879
rect 1571 875 1572 879
rect 1566 874 1572 875
rect 542 868 548 869
rect 750 868 756 869
rect 974 868 980 869
rect 1206 868 1212 869
rect 1438 868 1444 869
rect 542 864 543 868
rect 547 864 548 868
rect 690 867 696 868
rect 690 866 691 867
rect 613 864 691 866
rect 542 863 548 864
rect 690 863 691 864
rect 695 863 696 867
rect 750 864 751 868
rect 755 864 756 868
rect 894 867 900 868
rect 894 866 895 867
rect 821 864 895 866
rect 750 863 756 864
rect 894 863 895 864
rect 899 863 900 867
rect 974 864 975 868
rect 979 864 980 868
rect 1122 867 1128 868
rect 1122 866 1123 867
rect 1045 864 1123 866
rect 974 863 980 864
rect 1122 863 1123 864
rect 1127 863 1128 867
rect 1206 864 1207 868
rect 1211 864 1212 868
rect 1206 863 1212 864
rect 1238 867 1244 868
rect 1238 863 1239 867
rect 1243 863 1244 867
rect 1438 864 1439 868
rect 1443 864 1444 868
rect 1438 863 1444 864
rect 1470 867 1476 868
rect 1470 863 1471 867
rect 1475 863 1476 867
rect 690 862 696 863
rect 894 862 900 863
rect 1122 862 1128 863
rect 1238 862 1244 863
rect 1470 862 1476 863
rect 774 848 780 849
rect 926 848 932 849
rect 774 844 775 848
rect 779 844 780 848
rect 878 847 884 848
rect 878 846 879 847
rect 845 844 879 846
rect 774 843 780 844
rect 878 843 879 844
rect 883 843 884 847
rect 926 844 927 848
rect 931 844 932 848
rect 926 843 932 844
rect 1086 848 1092 849
rect 1086 844 1087 848
rect 1091 844 1092 848
rect 1086 843 1092 844
rect 1254 848 1260 849
rect 1422 848 1428 849
rect 1254 844 1255 848
rect 1259 844 1260 848
rect 1254 843 1260 844
rect 1286 847 1292 848
rect 1286 843 1287 847
rect 1291 843 1292 847
rect 1422 844 1423 848
rect 1427 844 1428 848
rect 1422 843 1428 844
rect 1454 847 1460 848
rect 1454 843 1455 847
rect 1459 843 1460 847
rect 878 842 884 843
rect 1286 842 1292 843
rect 1454 842 1460 843
rect 110 837 116 838
rect 110 833 111 837
rect 115 833 116 837
rect 110 832 116 833
rect 1566 837 1572 838
rect 1566 833 1567 837
rect 1571 833 1572 837
rect 1566 832 1572 833
rect 810 831 816 832
rect 810 827 811 831
rect 815 830 816 831
rect 967 831 973 832
rect 967 830 968 831
rect 815 828 968 830
rect 815 827 816 828
rect 810 826 816 827
rect 967 827 968 828
rect 972 827 973 831
rect 967 826 973 827
rect 978 831 984 832
rect 978 827 979 831
rect 983 830 984 831
rect 1127 831 1133 832
rect 1127 830 1128 831
rect 983 828 1128 830
rect 983 827 984 828
rect 978 826 984 827
rect 1127 827 1128 828
rect 1132 827 1133 831
rect 1127 826 1133 827
rect 110 819 116 820
rect 110 815 111 819
rect 115 815 116 819
rect 110 814 116 815
rect 1566 819 1572 820
rect 1566 815 1567 819
rect 1571 815 1572 819
rect 1566 814 1572 815
rect 807 803 816 804
rect 959 803 965 804
rect 774 802 780 803
rect 774 798 775 802
rect 779 798 780 802
rect 807 799 808 803
rect 815 799 816 803
rect 807 798 816 799
rect 926 802 932 803
rect 926 798 927 802
rect 931 798 932 802
rect 959 799 960 803
rect 964 802 965 803
rect 978 803 984 804
rect 1119 803 1125 804
rect 978 802 979 803
rect 964 800 979 802
rect 964 799 965 800
rect 959 798 965 799
rect 978 799 979 800
rect 983 799 984 803
rect 978 798 984 799
rect 1086 802 1092 803
rect 1086 798 1087 802
rect 1091 798 1092 802
rect 1119 799 1120 803
rect 1124 802 1125 803
rect 1238 803 1244 804
rect 1286 803 1293 804
rect 1455 803 1461 804
rect 1238 802 1239 803
rect 1124 800 1239 802
rect 1124 799 1125 800
rect 1119 798 1125 799
rect 1238 799 1239 800
rect 1243 799 1244 803
rect 1238 798 1244 799
rect 1254 802 1260 803
rect 1254 798 1255 802
rect 1259 798 1260 802
rect 1286 799 1287 803
rect 1292 799 1293 803
rect 1286 798 1293 799
rect 1422 802 1428 803
rect 1422 798 1423 802
rect 1427 798 1428 802
rect 1455 799 1456 803
rect 1460 802 1461 803
rect 1470 803 1476 804
rect 1470 802 1471 803
rect 1460 800 1471 802
rect 1460 799 1461 800
rect 1455 798 1461 799
rect 1470 799 1471 800
rect 1475 799 1476 803
rect 1470 798 1476 799
rect 774 797 780 798
rect 926 797 932 798
rect 1086 797 1092 798
rect 1254 797 1260 798
rect 1422 797 1428 798
rect 878 763 884 764
rect 854 762 860 763
rect 854 758 855 762
rect 859 758 860 762
rect 878 759 879 763
rect 883 762 884 763
rect 887 763 893 764
rect 1407 763 1413 764
rect 887 762 888 763
rect 883 760 888 762
rect 883 759 884 760
rect 878 758 884 759
rect 887 759 888 760
rect 892 759 893 763
rect 887 758 893 759
rect 974 762 980 763
rect 974 758 975 762
rect 979 758 980 762
rect 1102 762 1108 763
rect 1007 759 1013 760
rect 1007 758 1008 759
rect 854 757 860 758
rect 974 757 980 758
rect 1000 756 1008 758
rect 946 751 952 752
rect 946 747 947 751
rect 951 750 952 751
rect 1000 750 1002 756
rect 1007 755 1008 756
rect 1012 755 1013 759
rect 1102 758 1103 762
rect 1107 758 1108 762
rect 1238 762 1244 763
rect 1135 759 1141 760
rect 1135 758 1136 759
rect 1102 757 1108 758
rect 1007 754 1013 755
rect 1128 756 1136 758
rect 951 748 1002 750
rect 1070 751 1076 752
rect 951 747 952 748
rect 946 746 952 747
rect 1070 747 1071 751
rect 1075 750 1076 751
rect 1128 750 1130 756
rect 1135 755 1136 756
rect 1140 755 1141 759
rect 1238 758 1239 762
rect 1243 758 1244 762
rect 1374 762 1380 763
rect 1238 757 1244 758
rect 1262 759 1268 760
rect 1135 754 1141 755
rect 1262 755 1263 759
rect 1267 758 1268 759
rect 1271 759 1277 760
rect 1271 758 1272 759
rect 1267 756 1272 758
rect 1267 755 1268 756
rect 1262 754 1268 755
rect 1271 755 1272 756
rect 1276 755 1277 759
rect 1374 758 1375 762
rect 1379 758 1380 762
rect 1407 759 1408 763
rect 1412 762 1413 763
rect 1454 763 1460 764
rect 1454 762 1455 763
rect 1412 760 1455 762
rect 1412 759 1413 760
rect 1407 758 1413 759
rect 1454 759 1455 760
rect 1459 759 1460 763
rect 1454 758 1460 759
rect 1374 757 1380 758
rect 1271 754 1277 755
rect 1075 748 1130 750
rect 1075 747 1076 748
rect 1070 746 1076 747
rect 110 745 116 746
rect 110 741 111 745
rect 115 741 116 745
rect 110 740 116 741
rect 1566 745 1572 746
rect 1566 741 1567 745
rect 1571 741 1572 745
rect 1566 740 1572 741
rect 110 727 116 728
rect 110 723 111 727
rect 115 723 116 727
rect 110 722 116 723
rect 1566 727 1572 728
rect 1566 723 1567 727
rect 1571 723 1572 727
rect 1566 722 1572 723
rect 854 716 860 717
rect 974 716 980 717
rect 1102 716 1108 717
rect 1238 716 1244 717
rect 1374 716 1380 717
rect 854 712 855 716
rect 859 712 860 716
rect 946 715 952 716
rect 946 714 947 715
rect 925 712 947 714
rect 854 711 860 712
rect 946 711 947 712
rect 951 711 952 715
rect 974 712 975 716
rect 979 712 980 716
rect 1070 715 1076 716
rect 1070 714 1071 715
rect 1045 712 1071 714
rect 974 711 980 712
rect 1070 711 1071 712
rect 1075 711 1076 715
rect 1102 712 1103 716
rect 1107 712 1108 716
rect 1102 711 1108 712
rect 1158 715 1164 716
rect 1158 711 1159 715
rect 1163 711 1164 715
rect 1238 712 1239 716
rect 1243 712 1244 716
rect 1238 711 1244 712
rect 1286 715 1292 716
rect 1286 711 1287 715
rect 1291 711 1292 715
rect 1374 712 1375 716
rect 1379 712 1380 716
rect 1374 711 1380 712
rect 1406 715 1412 716
rect 1406 711 1407 715
rect 1411 711 1412 715
rect 946 710 952 711
rect 1070 710 1076 711
rect 1158 710 1164 711
rect 1286 710 1292 711
rect 1406 710 1412 711
rect 734 696 740 697
rect 934 696 940 697
rect 734 692 735 696
rect 739 692 740 696
rect 870 695 876 696
rect 870 694 871 695
rect 805 692 871 694
rect 734 691 740 692
rect 870 691 871 692
rect 875 691 876 695
rect 934 692 935 696
rect 939 692 940 696
rect 934 691 940 692
rect 1134 696 1140 697
rect 1134 692 1135 696
rect 1139 692 1140 696
rect 1134 691 1140 692
rect 1342 696 1348 697
rect 1342 692 1343 696
rect 1347 692 1348 696
rect 1342 691 1348 692
rect 870 690 876 691
rect 110 685 116 686
rect 110 681 111 685
rect 115 681 116 685
rect 110 680 116 681
rect 1566 685 1572 686
rect 1566 681 1567 685
rect 1571 681 1572 685
rect 1566 680 1572 681
rect 911 679 917 680
rect 911 675 912 679
rect 916 678 917 679
rect 975 679 981 680
rect 975 678 976 679
rect 916 676 976 678
rect 916 675 917 676
rect 911 674 917 675
rect 975 675 976 676
rect 980 675 981 679
rect 975 674 981 675
rect 986 679 992 680
rect 986 675 987 679
rect 991 678 992 679
rect 1175 679 1181 680
rect 1175 678 1176 679
rect 991 676 1176 678
rect 991 675 992 676
rect 986 674 992 675
rect 1175 675 1176 676
rect 1180 675 1181 679
rect 1175 674 1181 675
rect 1374 679 1380 680
rect 1374 675 1375 679
rect 1379 678 1380 679
rect 1383 679 1389 680
rect 1383 678 1384 679
rect 1379 676 1384 678
rect 1379 675 1380 676
rect 1374 674 1380 675
rect 1383 675 1384 676
rect 1388 675 1389 679
rect 1383 674 1389 675
rect 110 667 116 668
rect 110 663 111 667
rect 115 663 116 667
rect 110 662 116 663
rect 1566 667 1572 668
rect 1566 663 1567 667
rect 1571 663 1572 667
rect 1566 662 1572 663
rect 767 651 773 652
rect 734 650 740 651
rect 734 646 735 650
rect 739 646 740 650
rect 767 647 768 651
rect 772 650 773 651
rect 911 651 917 652
rect 967 651 973 652
rect 911 650 912 651
rect 772 648 912 650
rect 772 647 773 648
rect 767 646 773 647
rect 911 647 912 648
rect 916 647 917 651
rect 911 646 917 647
rect 934 650 940 651
rect 934 646 935 650
rect 939 646 940 650
rect 967 647 968 651
rect 972 650 973 651
rect 986 651 992 652
rect 1166 651 1173 652
rect 1375 651 1381 652
rect 986 650 987 651
rect 972 648 987 650
rect 972 647 973 648
rect 967 646 973 647
rect 986 647 987 648
rect 991 647 992 651
rect 986 646 992 647
rect 1134 650 1140 651
rect 1134 646 1135 650
rect 1139 646 1140 650
rect 1166 647 1167 651
rect 1172 647 1173 651
rect 1166 646 1173 647
rect 1342 650 1348 651
rect 1342 646 1343 650
rect 1347 646 1348 650
rect 1375 647 1376 651
rect 1380 650 1381 651
rect 1406 651 1412 652
rect 1406 650 1407 651
rect 1380 648 1407 650
rect 1380 647 1381 648
rect 1375 646 1381 647
rect 1406 647 1407 648
rect 1411 647 1412 651
rect 1406 646 1412 647
rect 734 645 740 646
rect 934 645 940 646
rect 1134 645 1140 646
rect 1342 645 1348 646
rect 870 627 876 628
rect 606 626 612 627
rect 606 622 607 626
rect 611 622 612 626
rect 846 626 852 627
rect 606 621 612 622
rect 639 623 645 624
rect 639 619 640 623
rect 644 622 645 623
rect 846 622 847 626
rect 851 622 852 626
rect 870 623 871 627
rect 875 626 876 627
rect 879 627 885 628
rect 1359 627 1365 628
rect 879 626 880 627
rect 875 624 880 626
rect 875 623 876 624
rect 870 622 876 623
rect 879 623 880 624
rect 884 623 885 627
rect 879 622 885 623
rect 1086 626 1092 627
rect 1086 622 1087 626
rect 1091 622 1092 626
rect 1326 626 1332 627
rect 644 620 782 622
rect 846 621 852 622
rect 1086 621 1092 622
rect 1118 623 1125 624
rect 644 619 645 620
rect 639 618 645 619
rect 780 614 782 620
rect 1118 619 1119 623
rect 1124 619 1125 623
rect 1326 622 1327 626
rect 1331 622 1332 626
rect 1359 623 1360 627
rect 1364 626 1365 627
rect 1374 627 1380 628
rect 1374 626 1375 627
rect 1364 624 1375 626
rect 1364 623 1365 624
rect 1359 622 1365 623
rect 1374 623 1375 624
rect 1379 623 1380 627
rect 1374 622 1380 623
rect 1326 621 1332 622
rect 1118 618 1125 619
rect 862 615 868 616
rect 862 614 863 615
rect 780 612 863 614
rect 862 611 863 612
rect 867 611 868 615
rect 862 610 868 611
rect 110 609 116 610
rect 110 605 111 609
rect 115 605 116 609
rect 110 604 116 605
rect 1566 609 1572 610
rect 1566 605 1567 609
rect 1571 605 1572 609
rect 1566 604 1572 605
rect 110 591 116 592
rect 110 587 111 591
rect 115 587 116 591
rect 110 586 116 587
rect 1566 591 1572 592
rect 1566 587 1567 591
rect 1571 587 1572 591
rect 1566 586 1572 587
rect 606 580 612 581
rect 606 576 607 580
rect 611 576 612 580
rect 846 580 852 581
rect 1086 580 1092 581
rect 1326 580 1332 581
rect 606 575 612 576
rect 390 571 396 572
rect 390 567 391 571
rect 395 570 396 571
rect 640 570 642 577
rect 846 576 847 580
rect 851 576 852 580
rect 846 575 852 576
rect 862 579 868 580
rect 862 575 863 579
rect 867 578 868 579
rect 867 576 881 578
rect 1086 576 1087 580
rect 1091 576 1092 580
rect 1262 579 1268 580
rect 1262 578 1263 579
rect 1157 576 1263 578
rect 867 575 868 576
rect 1086 575 1092 576
rect 1262 575 1263 576
rect 1267 575 1268 579
rect 1326 576 1327 580
rect 1331 576 1332 580
rect 1326 575 1332 576
rect 1358 579 1364 580
rect 1358 575 1359 579
rect 1363 575 1364 579
rect 862 574 868 575
rect 1262 574 1268 575
rect 1358 574 1364 575
rect 395 568 642 570
rect 395 567 396 568
rect 390 566 396 567
rect 358 560 364 561
rect 590 560 596 561
rect 830 560 836 561
rect 1078 560 1084 561
rect 1326 560 1332 561
rect 358 556 359 560
rect 363 556 364 560
rect 506 559 512 560
rect 506 558 507 559
rect 429 556 507 558
rect 358 555 364 556
rect 506 555 507 556
rect 511 555 512 559
rect 590 556 591 560
rect 595 556 596 560
rect 695 559 701 560
rect 695 558 696 559
rect 661 556 696 558
rect 590 555 596 556
rect 695 555 696 556
rect 700 555 701 559
rect 830 556 831 560
rect 835 556 836 560
rect 830 555 836 556
rect 862 559 868 560
rect 862 555 863 559
rect 867 555 868 559
rect 1078 556 1079 560
rect 1083 556 1084 560
rect 1078 555 1084 556
rect 1118 559 1124 560
rect 1118 555 1119 559
rect 1123 555 1124 559
rect 1326 556 1327 560
rect 1331 556 1332 560
rect 1326 555 1332 556
rect 1374 559 1380 560
rect 1374 555 1375 559
rect 1379 555 1380 559
rect 506 554 512 555
rect 695 554 701 555
rect 862 554 868 555
rect 1118 554 1124 555
rect 1374 554 1380 555
rect 110 549 116 550
rect 110 545 111 549
rect 115 545 116 549
rect 110 544 116 545
rect 1566 549 1572 550
rect 1566 545 1567 549
rect 1571 545 1572 549
rect 1566 544 1572 545
rect 110 531 116 532
rect 110 527 111 531
rect 115 527 116 531
rect 110 526 116 527
rect 1566 531 1572 532
rect 1566 527 1567 531
rect 1571 527 1572 531
rect 1566 526 1572 527
rect 506 523 512 524
rect 506 519 507 523
rect 511 522 512 523
rect 695 523 701 524
rect 511 520 618 522
rect 511 519 512 520
rect 506 518 512 519
rect 390 515 397 516
rect 358 514 364 515
rect 358 510 359 514
rect 363 510 364 514
rect 390 511 391 515
rect 396 511 397 515
rect 390 510 397 511
rect 590 514 596 515
rect 590 510 591 514
rect 595 510 596 514
rect 616 514 618 520
rect 695 519 696 523
rect 700 522 701 523
rect 700 520 858 522
rect 700 519 701 520
rect 695 518 701 519
rect 623 515 629 516
rect 623 514 624 515
rect 616 512 624 514
rect 623 511 624 512
rect 628 511 629 515
rect 623 510 629 511
rect 830 514 836 515
rect 830 510 831 514
rect 835 510 836 514
rect 856 514 858 520
rect 863 515 869 516
rect 1106 515 1117 516
rect 1358 515 1365 516
rect 863 514 864 515
rect 856 512 864 514
rect 863 511 864 512
rect 868 511 869 515
rect 863 510 869 511
rect 1078 514 1084 515
rect 1078 510 1079 514
rect 1083 510 1084 514
rect 1106 511 1107 515
rect 1111 511 1112 515
rect 1116 511 1117 515
rect 1106 510 1117 511
rect 1326 514 1332 515
rect 1326 510 1327 514
rect 1331 510 1332 514
rect 1358 511 1359 515
rect 1364 511 1365 515
rect 1358 510 1365 511
rect 358 509 364 510
rect 590 509 596 510
rect 830 509 836 510
rect 1078 509 1084 510
rect 1326 509 1332 510
rect 767 475 773 476
rect 150 474 156 475
rect 150 470 151 474
rect 155 470 156 474
rect 438 474 444 475
rect 150 469 156 470
rect 183 471 189 472
rect 183 467 184 471
rect 188 470 189 471
rect 438 470 439 474
rect 443 470 444 474
rect 734 474 740 475
rect 188 468 330 470
rect 438 469 444 470
rect 471 471 477 472
rect 188 467 189 468
rect 183 466 189 467
rect 328 462 330 468
rect 471 467 472 471
rect 476 470 477 471
rect 734 470 735 474
rect 739 470 740 474
rect 767 471 768 475
rect 772 474 773 475
rect 862 475 868 476
rect 1374 475 1381 476
rect 862 474 863 475
rect 772 472 863 474
rect 772 471 773 472
rect 767 470 773 471
rect 862 471 863 472
rect 867 471 868 475
rect 862 470 868 471
rect 1038 474 1044 475
rect 1038 470 1039 474
rect 1043 470 1044 474
rect 1342 474 1348 475
rect 476 468 681 470
rect 734 469 740 470
rect 1038 469 1044 470
rect 1070 471 1077 472
rect 476 467 477 468
rect 471 466 477 467
rect 454 463 460 464
rect 454 462 455 463
rect 328 460 455 462
rect 454 459 455 460
rect 459 459 460 463
rect 679 462 681 468
rect 1070 467 1071 471
rect 1076 467 1077 471
rect 1342 470 1343 474
rect 1347 470 1348 474
rect 1374 471 1375 475
rect 1380 471 1381 475
rect 1374 470 1381 471
rect 1342 469 1348 470
rect 1070 466 1077 467
rect 750 463 756 464
rect 750 462 751 463
rect 679 460 751 462
rect 454 458 460 459
rect 750 459 751 460
rect 755 459 756 463
rect 750 458 756 459
rect 110 457 116 458
rect 110 453 111 457
rect 115 453 116 457
rect 110 452 116 453
rect 1566 457 1572 458
rect 1566 453 1567 457
rect 1571 453 1572 457
rect 1566 452 1572 453
rect 110 439 116 440
rect 110 435 111 439
rect 115 435 116 439
rect 110 434 116 435
rect 1566 439 1572 440
rect 1566 435 1567 439
rect 1571 435 1572 439
rect 1566 434 1572 435
rect 1106 431 1112 432
rect 150 428 156 429
rect 438 428 444 429
rect 734 428 740 429
rect 1038 428 1044 429
rect 150 424 151 428
rect 155 424 156 428
rect 150 423 156 424
rect 206 427 212 428
rect 206 423 207 427
rect 211 423 212 427
rect 438 424 439 428
rect 443 424 444 428
rect 438 423 444 424
rect 454 427 460 428
rect 454 423 455 427
rect 459 426 460 427
rect 459 424 473 426
rect 734 424 735 428
rect 739 424 740 428
rect 459 423 460 424
rect 734 423 740 424
rect 750 427 756 428
rect 750 423 751 427
rect 755 426 756 427
rect 755 424 769 426
rect 1038 424 1039 428
rect 1043 424 1044 428
rect 1106 427 1107 431
rect 1111 427 1112 431
rect 1106 426 1112 427
rect 1342 428 1348 429
rect 755 423 756 424
rect 1038 423 1044 424
rect 1342 424 1343 428
rect 1347 424 1348 428
rect 1342 423 1348 424
rect 1398 427 1404 428
rect 1398 423 1399 427
rect 1403 423 1404 427
rect 206 422 212 423
rect 454 422 460 423
rect 750 422 756 423
rect 1398 422 1404 423
rect 174 404 180 405
rect 566 404 572 405
rect 966 404 972 405
rect 1366 404 1372 405
rect 174 400 175 404
rect 179 400 180 404
rect 498 403 504 404
rect 498 402 499 403
rect 245 400 499 402
rect 174 399 180 400
rect 498 399 499 400
rect 503 399 504 403
rect 566 400 567 404
rect 571 400 572 404
rect 830 403 836 404
rect 830 402 831 403
rect 637 400 831 402
rect 566 399 572 400
rect 830 399 831 400
rect 835 399 836 403
rect 966 400 967 404
rect 971 400 972 404
rect 1070 403 1076 404
rect 1070 402 1071 403
rect 1037 400 1071 402
rect 966 399 972 400
rect 1070 399 1071 400
rect 1075 399 1076 403
rect 1366 400 1367 404
rect 1371 400 1372 404
rect 1366 399 1372 400
rect 1430 403 1436 404
rect 1430 399 1431 403
rect 1435 399 1436 403
rect 498 398 504 399
rect 830 398 836 399
rect 1070 398 1076 399
rect 1430 398 1436 399
rect 110 393 116 394
rect 110 389 111 393
rect 115 389 116 393
rect 110 388 116 389
rect 1566 393 1572 394
rect 1566 389 1567 393
rect 1571 389 1572 393
rect 1566 388 1572 389
rect 110 375 116 376
rect 110 371 111 375
rect 115 371 116 375
rect 110 370 116 371
rect 1566 375 1572 376
rect 1566 371 1567 375
rect 1571 371 1572 375
rect 1566 370 1572 371
rect 498 367 504 368
rect 498 363 499 367
rect 503 366 504 367
rect 503 364 594 366
rect 503 363 504 364
rect 498 362 504 363
rect 206 359 213 360
rect 174 358 180 359
rect 174 354 175 358
rect 179 354 180 358
rect 206 355 207 359
rect 212 355 213 359
rect 206 354 213 355
rect 566 358 572 359
rect 566 354 567 358
rect 571 354 572 358
rect 592 358 594 364
rect 599 359 605 360
rect 999 359 1005 360
rect 599 358 600 359
rect 592 356 600 358
rect 599 355 600 356
rect 604 355 605 359
rect 599 354 605 355
rect 966 358 972 359
rect 966 354 967 358
rect 971 354 972 358
rect 999 355 1000 359
rect 1004 358 1005 359
rect 1126 359 1132 360
rect 1398 359 1405 360
rect 1126 358 1127 359
rect 1004 356 1127 358
rect 1004 355 1005 356
rect 999 354 1005 355
rect 1126 355 1127 356
rect 1131 355 1132 359
rect 1126 354 1132 355
rect 1366 358 1372 359
rect 1366 354 1367 358
rect 1371 354 1372 358
rect 1398 355 1399 359
rect 1404 355 1405 359
rect 1398 354 1405 355
rect 174 353 180 354
rect 566 353 572 354
rect 966 353 972 354
rect 1366 353 1372 354
rect 830 331 837 332
rect 1430 331 1437 332
rect 230 330 236 331
rect 230 326 231 330
rect 235 326 236 330
rect 510 330 516 331
rect 230 325 236 326
rect 263 327 269 328
rect 263 323 264 327
rect 268 326 269 327
rect 510 326 511 330
rect 515 326 516 330
rect 798 330 804 331
rect 268 324 406 326
rect 510 325 516 326
rect 543 327 549 328
rect 268 323 269 324
rect 263 322 269 323
rect 404 318 406 324
rect 543 323 544 327
rect 548 326 549 327
rect 798 326 799 330
rect 803 326 804 330
rect 830 327 831 331
rect 836 327 837 331
rect 830 326 837 327
rect 1094 330 1100 331
rect 1094 326 1095 330
rect 1099 326 1100 330
rect 1398 330 1404 331
rect 548 324 681 326
rect 798 325 804 326
rect 1094 325 1100 326
rect 1119 327 1125 328
rect 548 323 549 324
rect 543 322 549 323
rect 526 319 532 320
rect 526 318 527 319
rect 404 316 527 318
rect 526 315 527 316
rect 531 315 532 319
rect 679 318 681 324
rect 1119 323 1120 327
rect 1124 326 1125 327
rect 1127 327 1133 328
rect 1127 326 1128 327
rect 1124 324 1128 326
rect 1124 323 1125 324
rect 1119 322 1125 323
rect 1127 323 1128 324
rect 1132 323 1133 327
rect 1398 326 1399 330
rect 1403 326 1404 330
rect 1430 327 1431 331
rect 1436 327 1437 331
rect 1430 326 1437 327
rect 1398 325 1404 326
rect 1127 322 1133 323
rect 814 319 820 320
rect 814 318 815 319
rect 679 316 815 318
rect 526 314 532 315
rect 814 315 815 316
rect 819 315 820 319
rect 814 314 820 315
rect 110 313 116 314
rect 110 309 111 313
rect 115 309 116 313
rect 110 308 116 309
rect 1566 313 1572 314
rect 1566 309 1567 313
rect 1571 309 1572 313
rect 1566 308 1572 309
rect 110 295 116 296
rect 110 291 111 295
rect 115 291 116 295
rect 110 290 116 291
rect 1566 295 1572 296
rect 1566 291 1567 295
rect 1571 291 1572 295
rect 1566 290 1572 291
rect 230 284 236 285
rect 510 284 516 285
rect 798 284 804 285
rect 1094 284 1100 285
rect 1398 284 1404 285
rect 230 280 231 284
rect 235 280 236 284
rect 446 283 452 284
rect 446 282 447 283
rect 301 280 447 282
rect 230 279 236 280
rect 446 279 447 280
rect 451 279 452 283
rect 510 280 511 284
rect 515 280 516 284
rect 510 279 516 280
rect 526 283 532 284
rect 526 279 527 283
rect 531 282 532 283
rect 531 280 545 282
rect 798 280 799 284
rect 803 280 804 284
rect 531 279 532 280
rect 798 279 804 280
rect 814 283 820 284
rect 814 279 815 283
rect 819 282 820 283
rect 819 280 833 282
rect 1094 280 1095 284
rect 1099 280 1100 284
rect 819 279 820 280
rect 1094 279 1100 280
rect 1126 283 1132 284
rect 1126 279 1127 283
rect 1131 279 1132 283
rect 1398 280 1399 284
rect 1403 280 1404 284
rect 1398 279 1404 280
rect 1454 283 1460 284
rect 1454 279 1455 283
rect 1459 279 1460 283
rect 446 278 452 279
rect 526 278 532 279
rect 814 278 820 279
rect 1126 278 1132 279
rect 1454 278 1460 279
rect 422 256 428 257
rect 662 256 668 257
rect 422 252 423 256
rect 427 252 428 256
rect 566 255 572 256
rect 566 254 567 255
rect 493 252 567 254
rect 422 251 428 252
rect 566 251 567 252
rect 571 251 572 255
rect 662 252 663 256
rect 667 252 668 256
rect 662 251 668 252
rect 910 256 916 257
rect 1166 256 1172 257
rect 910 252 911 256
rect 915 252 916 256
rect 1119 255 1125 256
rect 1119 254 1120 255
rect 981 252 1120 254
rect 910 251 916 252
rect 1119 251 1120 252
rect 1124 251 1125 255
rect 1166 252 1167 256
rect 1171 252 1172 256
rect 1166 251 1172 252
rect 1430 256 1436 257
rect 1430 252 1431 256
rect 1435 252 1436 256
rect 1430 251 1436 252
rect 1498 255 1504 256
rect 1498 251 1499 255
rect 1503 251 1504 255
rect 566 250 572 251
rect 1119 250 1125 251
rect 1498 250 1504 251
rect 110 245 116 246
rect 110 241 111 245
rect 115 241 116 245
rect 110 240 116 241
rect 1566 245 1572 246
rect 1566 241 1567 245
rect 1571 241 1572 245
rect 1566 240 1572 241
rect 574 239 580 240
rect 574 235 575 239
rect 579 238 580 239
rect 703 239 709 240
rect 703 238 704 239
rect 579 236 704 238
rect 579 235 580 236
rect 574 234 580 235
rect 703 235 704 236
rect 708 235 709 239
rect 703 234 709 235
rect 946 239 952 240
rect 946 235 947 239
rect 951 238 952 239
rect 1207 239 1213 240
rect 1207 238 1208 239
rect 951 236 1208 238
rect 951 235 952 236
rect 946 234 952 235
rect 1207 235 1208 236
rect 1212 235 1213 239
rect 1207 234 1213 235
rect 110 227 116 228
rect 110 223 111 227
rect 115 223 116 227
rect 110 222 116 223
rect 1566 227 1572 228
rect 1566 223 1567 227
rect 1571 223 1572 227
rect 1566 222 1572 223
rect 566 219 572 220
rect 566 215 567 219
rect 571 218 572 219
rect 571 216 690 218
rect 571 215 572 216
rect 566 214 572 215
rect 446 211 452 212
rect 422 210 428 211
rect 422 206 423 210
rect 427 206 428 210
rect 446 207 447 211
rect 451 210 452 211
rect 455 211 461 212
rect 455 210 456 211
rect 451 208 456 210
rect 451 207 452 208
rect 446 206 452 207
rect 455 207 456 208
rect 460 207 461 211
rect 455 206 461 207
rect 662 210 668 211
rect 662 206 663 210
rect 667 206 668 210
rect 688 210 690 216
rect 695 211 701 212
rect 943 211 952 212
rect 1198 211 1205 212
rect 1454 211 1460 212
rect 695 210 696 211
rect 688 208 696 210
rect 695 207 696 208
rect 700 207 701 211
rect 695 206 701 207
rect 910 210 916 211
rect 910 206 911 210
rect 915 206 916 210
rect 943 207 944 211
rect 951 207 952 211
rect 943 206 952 207
rect 1166 210 1172 211
rect 1166 206 1167 210
rect 1171 206 1172 210
rect 1198 207 1199 211
rect 1204 207 1205 211
rect 1198 206 1205 207
rect 1430 210 1436 211
rect 1430 206 1431 210
rect 1435 206 1436 210
rect 1454 207 1455 211
rect 1459 210 1460 211
rect 1463 211 1469 212
rect 1463 210 1464 211
rect 1459 208 1464 210
rect 1459 207 1460 208
rect 1454 206 1460 207
rect 1463 207 1464 208
rect 1468 207 1469 211
rect 1463 206 1469 207
rect 422 205 428 206
rect 662 205 668 206
rect 910 205 916 206
rect 1166 205 1172 206
rect 1430 205 1436 206
rect 543 171 549 172
rect 510 170 516 171
rect 510 166 511 170
rect 515 166 516 170
rect 543 167 544 171
rect 548 170 549 171
rect 574 171 580 172
rect 1498 171 1509 172
rect 574 170 575 171
rect 548 168 575 170
rect 548 167 549 168
rect 543 166 549 167
rect 574 167 575 168
rect 579 167 580 171
rect 574 166 580 167
rect 614 170 620 171
rect 614 166 615 170
rect 619 166 620 170
rect 726 170 732 171
rect 647 167 653 168
rect 647 166 648 167
rect 510 165 516 166
rect 614 165 620 166
rect 640 164 648 166
rect 594 159 600 160
rect 594 155 595 159
rect 599 158 600 159
rect 640 158 642 164
rect 647 163 648 164
rect 652 163 653 167
rect 726 166 727 170
rect 731 166 732 170
rect 854 170 860 171
rect 759 167 765 168
rect 759 166 760 167
rect 726 165 732 166
rect 647 162 653 163
rect 752 164 760 166
rect 599 156 642 158
rect 718 159 724 160
rect 599 155 600 156
rect 594 154 600 155
rect 718 155 719 159
rect 723 158 724 159
rect 752 158 754 164
rect 759 163 760 164
rect 764 163 765 167
rect 854 166 855 170
rect 859 166 860 170
rect 998 170 1004 171
rect 887 167 893 168
rect 887 166 888 167
rect 854 165 860 166
rect 759 162 765 163
rect 880 164 888 166
rect 723 156 754 158
rect 822 159 828 160
rect 723 155 724 156
rect 718 154 724 155
rect 822 155 823 159
rect 827 158 828 159
rect 880 158 882 164
rect 887 163 888 164
rect 892 163 893 167
rect 998 166 999 170
rect 1003 166 1004 170
rect 1158 170 1164 171
rect 1031 167 1037 168
rect 1031 166 1032 167
rect 998 165 1004 166
rect 887 162 893 163
rect 1024 164 1032 166
rect 827 156 882 158
rect 958 159 964 160
rect 827 155 828 156
rect 822 154 828 155
rect 958 155 959 159
rect 963 158 964 159
rect 1024 158 1026 164
rect 1031 163 1032 164
rect 1036 163 1037 167
rect 1158 166 1159 170
rect 1163 166 1164 170
rect 1326 170 1332 171
rect 1191 167 1197 168
rect 1191 166 1192 167
rect 1158 165 1164 166
rect 1031 162 1037 163
rect 1184 164 1192 166
rect 963 156 1026 158
rect 1110 159 1116 160
rect 963 155 964 156
rect 958 154 964 155
rect 1110 155 1111 159
rect 1115 158 1116 159
rect 1184 158 1186 164
rect 1191 163 1192 164
rect 1196 163 1197 167
rect 1326 166 1327 170
rect 1331 166 1332 170
rect 1470 170 1476 171
rect 1326 165 1332 166
rect 1359 167 1365 168
rect 1191 162 1197 163
rect 1359 163 1360 167
rect 1364 166 1365 167
rect 1470 166 1471 170
rect 1475 166 1476 170
rect 1498 167 1499 171
rect 1503 167 1504 171
rect 1508 167 1509 171
rect 1498 166 1509 167
rect 1364 164 1434 166
rect 1470 165 1476 166
rect 1364 163 1365 164
rect 1359 162 1365 163
rect 1115 156 1186 158
rect 1432 158 1434 164
rect 1486 159 1492 160
rect 1486 158 1487 159
rect 1432 156 1487 158
rect 1115 155 1116 156
rect 1110 154 1116 155
rect 1486 155 1487 156
rect 1491 155 1492 159
rect 1486 154 1492 155
rect 110 153 116 154
rect 110 149 111 153
rect 115 149 116 153
rect 110 148 116 149
rect 1566 153 1572 154
rect 1566 149 1567 153
rect 1571 149 1572 153
rect 1566 148 1572 149
rect 110 135 116 136
rect 110 131 111 135
rect 115 131 116 135
rect 110 130 116 131
rect 1566 135 1572 136
rect 1566 131 1567 135
rect 1571 131 1572 135
rect 1566 130 1572 131
rect 510 124 516 125
rect 614 124 620 125
rect 726 124 732 125
rect 854 124 860 125
rect 998 124 1004 125
rect 1158 124 1164 125
rect 1326 124 1332 125
rect 510 120 511 124
rect 515 120 516 124
rect 594 123 600 124
rect 594 122 595 123
rect 581 120 595 122
rect 510 119 516 120
rect 594 119 595 120
rect 599 119 600 123
rect 614 120 615 124
rect 619 120 620 124
rect 718 123 724 124
rect 718 122 719 123
rect 685 120 719 122
rect 614 119 620 120
rect 718 119 719 120
rect 723 119 724 123
rect 726 120 727 124
rect 731 120 732 124
rect 822 123 828 124
rect 822 122 823 123
rect 797 120 823 122
rect 726 119 732 120
rect 822 119 823 120
rect 827 119 828 123
rect 854 120 855 124
rect 859 120 860 124
rect 958 123 964 124
rect 958 122 959 123
rect 925 120 959 122
rect 854 119 860 120
rect 958 119 959 120
rect 963 119 964 123
rect 998 120 999 124
rect 1003 120 1004 124
rect 1110 123 1116 124
rect 1110 122 1111 123
rect 1069 120 1111 122
rect 998 119 1004 120
rect 1110 119 1111 120
rect 1115 119 1116 123
rect 1158 120 1159 124
rect 1163 120 1164 124
rect 1158 119 1164 120
rect 1198 123 1204 124
rect 1198 119 1199 123
rect 1203 119 1204 123
rect 1326 120 1327 124
rect 1331 120 1332 124
rect 1326 119 1332 120
rect 1470 124 1476 125
rect 1470 120 1471 124
rect 1475 120 1476 124
rect 1470 119 1476 120
rect 1486 123 1492 124
rect 1486 119 1487 123
rect 1491 122 1492 123
rect 1491 120 1505 122
rect 1491 119 1492 120
rect 594 118 600 119
rect 718 118 724 119
rect 822 118 828 119
rect 958 118 964 119
rect 1110 118 1116 119
rect 1198 118 1204 119
rect 1486 118 1492 119
<< m3c >>
rect 135 1638 139 1642
rect 223 1638 227 1642
rect 211 1627 215 1631
rect 311 1638 315 1642
rect 299 1627 303 1631
rect 111 1621 115 1625
rect 1567 1621 1571 1625
rect 111 1603 115 1607
rect 1567 1603 1571 1607
rect 135 1592 139 1596
rect 211 1591 215 1595
rect 223 1592 227 1596
rect 299 1591 303 1595
rect 311 1592 315 1596
rect 327 1591 331 1595
rect 183 1580 187 1584
rect 259 1579 263 1583
rect 271 1580 275 1584
rect 347 1579 351 1583
rect 359 1580 363 1584
rect 383 1579 387 1583
rect 111 1569 115 1573
rect 1567 1569 1571 1573
rect 111 1551 115 1555
rect 1567 1551 1571 1555
rect 259 1543 263 1547
rect 183 1534 187 1538
rect 271 1534 275 1538
rect 347 1543 351 1547
rect 359 1534 363 1538
rect 327 1527 331 1531
rect 351 1502 355 1506
rect 383 1503 384 1507
rect 384 1503 387 1507
rect 439 1502 443 1506
rect 427 1491 431 1495
rect 527 1502 531 1506
rect 515 1491 519 1495
rect 615 1502 619 1506
rect 603 1491 607 1495
rect 111 1485 115 1489
rect 1567 1485 1571 1489
rect 111 1467 115 1471
rect 1567 1467 1571 1471
rect 351 1456 355 1460
rect 427 1455 431 1459
rect 439 1456 443 1460
rect 515 1455 519 1459
rect 527 1456 531 1460
rect 603 1455 607 1459
rect 615 1456 619 1460
rect 663 1424 667 1428
rect 739 1423 743 1427
rect 751 1424 755 1428
rect 827 1423 831 1427
rect 839 1424 843 1428
rect 915 1423 919 1427
rect 927 1424 931 1428
rect 111 1413 115 1417
rect 1567 1413 1571 1417
rect 851 1407 855 1411
rect 111 1395 115 1399
rect 1567 1395 1571 1399
rect 739 1387 743 1391
rect 663 1378 667 1382
rect 751 1378 755 1382
rect 827 1387 831 1391
rect 839 1378 843 1382
rect 915 1387 919 1391
rect 927 1378 931 1382
rect 815 1342 819 1346
rect 851 1343 852 1347
rect 852 1343 855 1347
rect 935 1342 939 1346
rect 907 1331 911 1335
rect 1055 1342 1059 1346
rect 1027 1331 1031 1335
rect 1175 1342 1179 1346
rect 1247 1339 1251 1343
rect 1295 1342 1299 1346
rect 1267 1331 1271 1335
rect 1415 1342 1419 1346
rect 1387 1331 1391 1335
rect 111 1325 115 1329
rect 1567 1325 1571 1329
rect 111 1307 115 1311
rect 1567 1307 1571 1311
rect 815 1296 819 1300
rect 907 1295 911 1299
rect 935 1296 939 1300
rect 1027 1295 1031 1299
rect 1055 1296 1059 1300
rect 1087 1295 1091 1299
rect 1175 1296 1179 1300
rect 1267 1295 1271 1299
rect 1295 1296 1299 1300
rect 1387 1295 1391 1299
rect 1415 1296 1419 1300
rect 1447 1295 1451 1299
rect 543 1284 547 1288
rect 627 1283 631 1287
rect 695 1284 699 1288
rect 863 1284 867 1288
rect 927 1283 931 1287
rect 1039 1284 1043 1288
rect 1215 1284 1219 1288
rect 1247 1283 1251 1287
rect 1399 1284 1403 1288
rect 1439 1283 1443 1287
rect 111 1273 115 1277
rect 1567 1273 1571 1277
rect 687 1267 691 1271
rect 111 1255 115 1259
rect 1567 1255 1571 1259
rect 627 1247 631 1251
rect 543 1238 547 1242
rect 687 1239 691 1243
rect 695 1238 699 1242
rect 863 1238 867 1242
rect 1039 1238 1043 1242
rect 1087 1239 1091 1243
rect 1215 1238 1219 1242
rect 1239 1239 1243 1243
rect 1399 1238 1403 1242
rect 1447 1239 1451 1243
rect 199 1194 203 1198
rect 415 1194 419 1198
rect 647 1194 651 1198
rect 431 1183 435 1187
rect 895 1194 899 1198
rect 927 1195 928 1199
rect 928 1195 931 1199
rect 1151 1194 1155 1198
rect 663 1183 667 1187
rect 1207 1191 1211 1195
rect 1415 1194 1419 1198
rect 1439 1195 1443 1199
rect 911 1183 915 1187
rect 111 1177 115 1181
rect 1567 1177 1571 1181
rect 111 1159 115 1163
rect 1567 1159 1571 1163
rect 199 1148 203 1152
rect 231 1147 235 1151
rect 415 1148 419 1152
rect 431 1147 435 1151
rect 647 1148 651 1152
rect 663 1147 667 1151
rect 895 1148 899 1152
rect 911 1147 915 1151
rect 1151 1148 1155 1152
rect 1239 1147 1243 1151
rect 1415 1148 1419 1152
rect 1447 1147 1451 1151
rect 135 1128 139 1132
rect 379 1127 383 1131
rect 559 1128 563 1132
rect 751 1127 755 1131
rect 991 1128 995 1132
rect 1059 1127 1063 1131
rect 1423 1128 1427 1132
rect 1463 1127 1467 1131
rect 111 1117 115 1121
rect 1567 1117 1571 1121
rect 111 1099 115 1103
rect 1567 1099 1571 1103
rect 379 1091 383 1095
rect 135 1082 139 1086
rect 231 1083 235 1087
rect 559 1082 563 1086
rect 619 1087 623 1091
rect 751 1091 755 1095
rect 991 1082 995 1086
rect 1447 1087 1451 1091
rect 1423 1082 1427 1086
rect 1047 1075 1051 1079
rect 239 1054 243 1058
rect 619 1055 623 1059
rect 631 1054 635 1058
rect 499 1043 503 1047
rect 1031 1054 1035 1058
rect 1059 1055 1063 1059
rect 1431 1054 1435 1058
rect 1463 1055 1464 1059
rect 1464 1055 1467 1059
rect 111 1037 115 1041
rect 1567 1037 1571 1041
rect 111 1019 115 1023
rect 1567 1019 1571 1023
rect 239 1008 243 1012
rect 499 1007 503 1011
rect 631 1008 635 1012
rect 687 1007 691 1011
rect 1031 1008 1035 1012
rect 1047 1007 1051 1011
rect 1431 1008 1435 1012
rect 1463 1007 1467 1011
rect 415 996 419 1000
rect 567 995 571 999
rect 663 996 667 1000
rect 823 995 827 999
rect 919 996 923 1000
rect 951 995 955 999
rect 1175 996 1179 1000
rect 1207 995 1211 999
rect 1439 996 1443 1000
rect 1471 995 1475 999
rect 111 985 115 989
rect 1567 985 1571 989
rect 111 967 115 971
rect 1567 967 1571 971
rect 823 959 827 963
rect 415 950 419 954
rect 663 950 667 954
rect 687 951 691 955
rect 919 950 923 954
rect 1175 950 1179 954
rect 1287 951 1291 955
rect 1439 950 1443 954
rect 1463 951 1467 955
rect 951 943 955 947
rect 543 910 547 914
rect 567 911 571 915
rect 751 910 755 914
rect 691 899 695 903
rect 975 910 979 914
rect 895 899 899 903
rect 1207 910 1211 914
rect 1123 899 1127 903
rect 1439 910 1443 914
rect 1471 911 1472 915
rect 1472 911 1475 915
rect 111 893 115 897
rect 1567 893 1571 897
rect 111 875 115 879
rect 1567 875 1571 879
rect 543 864 547 868
rect 691 863 695 867
rect 751 864 755 868
rect 895 863 899 867
rect 975 864 979 868
rect 1123 863 1127 867
rect 1207 864 1211 868
rect 1239 863 1243 867
rect 1439 864 1443 868
rect 1471 863 1475 867
rect 775 844 779 848
rect 879 843 883 847
rect 927 844 931 848
rect 1087 844 1091 848
rect 1255 844 1259 848
rect 1287 843 1291 847
rect 1423 844 1427 848
rect 1455 843 1459 847
rect 111 833 115 837
rect 1567 833 1571 837
rect 811 827 815 831
rect 979 827 983 831
rect 111 815 115 819
rect 1567 815 1571 819
rect 775 798 779 802
rect 811 799 812 803
rect 812 799 815 803
rect 927 798 931 802
rect 979 799 983 803
rect 1087 798 1091 802
rect 1239 799 1243 803
rect 1255 798 1259 802
rect 1287 799 1288 803
rect 1288 799 1291 803
rect 1423 798 1427 802
rect 1471 799 1475 803
rect 855 758 859 762
rect 879 759 883 763
rect 975 758 979 762
rect 947 747 951 751
rect 1103 758 1107 762
rect 1071 747 1075 751
rect 1239 758 1243 762
rect 1263 755 1267 759
rect 1375 758 1379 762
rect 1455 759 1459 763
rect 111 741 115 745
rect 1567 741 1571 745
rect 111 723 115 727
rect 1567 723 1571 727
rect 855 712 859 716
rect 947 711 951 715
rect 975 712 979 716
rect 1071 711 1075 715
rect 1103 712 1107 716
rect 1159 711 1163 715
rect 1239 712 1243 716
rect 1287 711 1291 715
rect 1375 712 1379 716
rect 1407 711 1411 715
rect 735 692 739 696
rect 871 691 875 695
rect 935 692 939 696
rect 1135 692 1139 696
rect 1343 692 1347 696
rect 111 681 115 685
rect 1567 681 1571 685
rect 987 675 991 679
rect 1375 675 1379 679
rect 111 663 115 667
rect 1567 663 1571 667
rect 735 646 739 650
rect 935 646 939 650
rect 987 647 991 651
rect 1135 646 1139 650
rect 1167 647 1168 651
rect 1168 647 1171 651
rect 1343 646 1347 650
rect 1407 647 1411 651
rect 607 622 611 626
rect 847 622 851 626
rect 871 623 875 627
rect 1087 622 1091 626
rect 1119 619 1120 623
rect 1120 619 1123 623
rect 1327 622 1331 626
rect 1375 623 1379 627
rect 863 611 867 615
rect 111 605 115 609
rect 1567 605 1571 609
rect 111 587 115 591
rect 1567 587 1571 591
rect 607 576 611 580
rect 391 567 395 571
rect 847 576 851 580
rect 863 575 867 579
rect 1087 576 1091 580
rect 1263 575 1267 579
rect 1327 576 1331 580
rect 1359 575 1363 579
rect 359 556 363 560
rect 507 555 511 559
rect 591 556 595 560
rect 831 556 835 560
rect 863 555 867 559
rect 1079 556 1083 560
rect 1119 555 1123 559
rect 1327 556 1331 560
rect 1375 555 1379 559
rect 111 545 115 549
rect 1567 545 1571 549
rect 111 527 115 531
rect 1567 527 1571 531
rect 507 519 511 523
rect 359 510 363 514
rect 391 511 392 515
rect 392 511 395 515
rect 591 510 595 514
rect 831 510 835 514
rect 1079 510 1083 514
rect 1107 511 1111 515
rect 1327 510 1331 514
rect 1359 511 1360 515
rect 1360 511 1363 515
rect 151 470 155 474
rect 439 470 443 474
rect 735 470 739 474
rect 863 471 867 475
rect 1039 470 1043 474
rect 455 459 459 463
rect 1071 467 1072 471
rect 1072 467 1075 471
rect 1343 470 1347 474
rect 1375 471 1376 475
rect 1376 471 1379 475
rect 751 459 755 463
rect 111 453 115 457
rect 1567 453 1571 457
rect 111 435 115 439
rect 1567 435 1571 439
rect 151 424 155 428
rect 207 423 211 427
rect 439 424 443 428
rect 455 423 459 427
rect 735 424 739 428
rect 751 423 755 427
rect 1039 424 1043 428
rect 1107 427 1111 431
rect 1343 424 1347 428
rect 1399 423 1403 427
rect 175 400 179 404
rect 499 399 503 403
rect 567 400 571 404
rect 831 399 835 403
rect 967 400 971 404
rect 1071 399 1075 403
rect 1367 400 1371 404
rect 1431 399 1435 403
rect 111 389 115 393
rect 1567 389 1571 393
rect 111 371 115 375
rect 1567 371 1571 375
rect 499 363 503 367
rect 175 354 179 358
rect 207 355 208 359
rect 208 355 211 359
rect 567 354 571 358
rect 967 354 971 358
rect 1127 355 1131 359
rect 1367 354 1371 358
rect 1399 355 1400 359
rect 1400 355 1403 359
rect 231 326 235 330
rect 511 326 515 330
rect 799 326 803 330
rect 831 327 832 331
rect 832 327 835 331
rect 1095 326 1099 330
rect 527 315 531 319
rect 1399 326 1403 330
rect 1431 327 1432 331
rect 1432 327 1435 331
rect 815 315 819 319
rect 111 309 115 313
rect 1567 309 1571 313
rect 111 291 115 295
rect 1567 291 1571 295
rect 231 280 235 284
rect 447 279 451 283
rect 511 280 515 284
rect 527 279 531 283
rect 799 280 803 284
rect 815 279 819 283
rect 1095 280 1099 284
rect 1127 279 1131 283
rect 1399 280 1403 284
rect 1455 279 1459 283
rect 423 252 427 256
rect 567 251 571 255
rect 663 252 667 256
rect 911 252 915 256
rect 1167 252 1171 256
rect 1431 252 1435 256
rect 1499 251 1503 255
rect 111 241 115 245
rect 1567 241 1571 245
rect 575 235 579 239
rect 947 235 951 239
rect 111 223 115 227
rect 1567 223 1571 227
rect 567 215 571 219
rect 423 206 427 210
rect 447 207 451 211
rect 663 206 667 210
rect 911 206 915 210
rect 947 207 948 211
rect 948 207 951 211
rect 1167 206 1171 210
rect 1199 207 1200 211
rect 1200 207 1203 211
rect 1431 206 1435 210
rect 1455 207 1459 211
rect 511 166 515 170
rect 575 167 579 171
rect 615 166 619 170
rect 595 155 599 159
rect 727 166 731 170
rect 719 155 723 159
rect 855 166 859 170
rect 823 155 827 159
rect 999 166 1003 170
rect 959 155 963 159
rect 1159 166 1163 170
rect 1111 155 1115 159
rect 1327 166 1331 170
rect 1471 166 1475 170
rect 1499 167 1503 171
rect 1487 155 1491 159
rect 111 149 115 153
rect 1567 149 1571 153
rect 111 131 115 135
rect 1567 131 1571 135
rect 511 120 515 124
rect 595 119 599 123
rect 615 120 619 124
rect 719 119 723 123
rect 727 120 731 124
rect 823 119 827 123
rect 855 120 859 124
rect 959 119 963 123
rect 999 120 1003 124
rect 1111 119 1115 123
rect 1159 120 1163 124
rect 1199 119 1203 123
rect 1327 120 1331 124
rect 1471 120 1475 124
rect 1487 119 1491 123
<< m3 >>
rect 111 1654 115 1655
rect 111 1649 115 1650
rect 135 1654 139 1655
rect 135 1649 139 1650
rect 223 1654 227 1655
rect 223 1649 227 1650
rect 311 1654 315 1655
rect 311 1649 315 1650
rect 1567 1654 1571 1655
rect 1567 1649 1571 1650
rect 112 1626 114 1649
rect 136 1643 138 1649
rect 224 1643 226 1649
rect 312 1643 314 1649
rect 134 1642 140 1643
rect 134 1638 135 1642
rect 139 1638 140 1642
rect 134 1637 140 1638
rect 222 1642 228 1643
rect 222 1638 223 1642
rect 227 1638 228 1642
rect 222 1637 228 1638
rect 310 1642 316 1643
rect 310 1638 311 1642
rect 315 1638 316 1642
rect 310 1637 316 1638
rect 210 1631 216 1632
rect 210 1627 211 1631
rect 215 1627 216 1631
rect 210 1626 216 1627
rect 298 1631 304 1632
rect 298 1627 299 1631
rect 303 1627 304 1631
rect 298 1626 304 1627
rect 1568 1626 1570 1649
rect 110 1625 116 1626
rect 110 1621 111 1625
rect 115 1621 116 1625
rect 110 1620 116 1621
rect 110 1607 116 1608
rect 110 1603 111 1607
rect 115 1603 116 1607
rect 110 1602 116 1603
rect 112 1591 114 1602
rect 134 1596 140 1597
rect 212 1596 214 1626
rect 222 1596 228 1597
rect 300 1596 302 1626
rect 1566 1625 1572 1626
rect 1566 1621 1567 1625
rect 1571 1621 1572 1625
rect 1566 1620 1572 1621
rect 1566 1607 1572 1608
rect 1566 1603 1567 1607
rect 1571 1603 1572 1607
rect 1566 1602 1572 1603
rect 310 1596 316 1597
rect 134 1592 135 1596
rect 139 1592 140 1596
rect 134 1591 140 1592
rect 210 1595 216 1596
rect 210 1591 211 1595
rect 215 1591 216 1595
rect 222 1592 223 1596
rect 227 1592 228 1596
rect 222 1591 228 1592
rect 298 1595 304 1596
rect 298 1591 299 1595
rect 303 1591 304 1595
rect 310 1592 311 1596
rect 315 1592 316 1596
rect 310 1591 316 1592
rect 326 1595 332 1596
rect 326 1591 327 1595
rect 331 1591 332 1595
rect 1568 1591 1570 1602
rect 111 1590 115 1591
rect 111 1585 115 1586
rect 135 1590 139 1591
rect 135 1585 139 1586
rect 183 1590 187 1591
rect 210 1590 216 1591
rect 223 1590 227 1591
rect 183 1585 187 1586
rect 223 1585 227 1586
rect 271 1590 275 1591
rect 298 1590 304 1591
rect 311 1590 315 1591
rect 326 1590 332 1591
rect 359 1590 363 1591
rect 271 1585 275 1586
rect 311 1585 315 1586
rect 112 1574 114 1585
rect 182 1584 188 1585
rect 270 1584 276 1585
rect 182 1580 183 1584
rect 187 1580 188 1584
rect 182 1579 188 1580
rect 258 1583 264 1584
rect 258 1579 259 1583
rect 263 1579 264 1583
rect 270 1580 271 1584
rect 275 1580 276 1584
rect 270 1579 276 1580
rect 258 1578 264 1579
rect 110 1573 116 1574
rect 110 1569 111 1573
rect 115 1569 116 1573
rect 110 1568 116 1569
rect 110 1555 116 1556
rect 110 1551 111 1555
rect 115 1551 116 1555
rect 110 1550 116 1551
rect 112 1519 114 1550
rect 260 1548 262 1578
rect 258 1547 264 1548
rect 258 1543 259 1547
rect 263 1543 264 1547
rect 258 1542 264 1543
rect 182 1538 188 1539
rect 182 1534 183 1538
rect 187 1534 188 1538
rect 182 1533 188 1534
rect 270 1538 276 1539
rect 270 1534 271 1538
rect 275 1534 276 1538
rect 270 1533 276 1534
rect 184 1519 186 1533
rect 272 1519 274 1533
rect 328 1532 330 1590
rect 359 1585 363 1586
rect 1567 1590 1571 1591
rect 1567 1585 1571 1586
rect 358 1584 364 1585
rect 346 1583 352 1584
rect 346 1579 347 1583
rect 351 1579 352 1583
rect 358 1580 359 1584
rect 363 1580 364 1584
rect 358 1579 364 1580
rect 382 1583 388 1584
rect 382 1579 383 1583
rect 387 1579 388 1583
rect 346 1578 352 1579
rect 382 1578 388 1579
rect 348 1548 350 1578
rect 346 1547 352 1548
rect 346 1543 347 1547
rect 351 1543 352 1547
rect 346 1542 352 1543
rect 358 1538 364 1539
rect 358 1534 359 1538
rect 363 1534 364 1538
rect 358 1533 364 1534
rect 326 1531 332 1532
rect 326 1527 327 1531
rect 331 1527 332 1531
rect 326 1526 332 1527
rect 360 1519 362 1533
rect 111 1518 115 1519
rect 111 1513 115 1514
rect 183 1518 187 1519
rect 183 1513 187 1514
rect 271 1518 275 1519
rect 271 1513 275 1514
rect 351 1518 355 1519
rect 351 1513 355 1514
rect 359 1518 363 1519
rect 359 1513 363 1514
rect 112 1490 114 1513
rect 352 1507 354 1513
rect 384 1508 386 1578
rect 1568 1574 1570 1585
rect 1566 1573 1572 1574
rect 1566 1569 1567 1573
rect 1571 1569 1572 1573
rect 1566 1568 1572 1569
rect 1566 1555 1572 1556
rect 1566 1551 1567 1555
rect 1571 1551 1572 1555
rect 1566 1550 1572 1551
rect 1568 1519 1570 1550
rect 439 1518 443 1519
rect 439 1513 443 1514
rect 527 1518 531 1519
rect 527 1513 531 1514
rect 615 1518 619 1519
rect 615 1513 619 1514
rect 1567 1518 1571 1519
rect 1567 1513 1571 1514
rect 382 1507 388 1508
rect 440 1507 442 1513
rect 528 1507 530 1513
rect 616 1507 618 1513
rect 350 1506 356 1507
rect 350 1502 351 1506
rect 355 1502 356 1506
rect 382 1503 383 1507
rect 387 1503 388 1507
rect 382 1502 388 1503
rect 438 1506 444 1507
rect 438 1502 439 1506
rect 443 1502 444 1506
rect 350 1501 356 1502
rect 438 1501 444 1502
rect 526 1506 532 1507
rect 526 1502 527 1506
rect 531 1502 532 1506
rect 526 1501 532 1502
rect 614 1506 620 1507
rect 614 1502 615 1506
rect 619 1502 620 1506
rect 614 1501 620 1502
rect 426 1495 432 1496
rect 426 1491 427 1495
rect 431 1491 432 1495
rect 426 1490 432 1491
rect 514 1495 520 1496
rect 514 1491 515 1495
rect 519 1491 520 1495
rect 514 1490 520 1491
rect 602 1495 608 1496
rect 602 1491 603 1495
rect 607 1491 608 1495
rect 602 1490 608 1491
rect 1568 1490 1570 1513
rect 110 1489 116 1490
rect 110 1485 111 1489
rect 115 1485 116 1489
rect 110 1484 116 1485
rect 110 1471 116 1472
rect 110 1467 111 1471
rect 115 1467 116 1471
rect 110 1466 116 1467
rect 112 1435 114 1466
rect 350 1460 356 1461
rect 428 1460 430 1490
rect 438 1460 444 1461
rect 516 1460 518 1490
rect 526 1460 532 1461
rect 604 1460 606 1490
rect 1566 1489 1572 1490
rect 1566 1485 1567 1489
rect 1571 1485 1572 1489
rect 1566 1484 1572 1485
rect 1566 1471 1572 1472
rect 1566 1467 1567 1471
rect 1571 1467 1572 1471
rect 1566 1466 1572 1467
rect 614 1460 620 1461
rect 350 1456 351 1460
rect 355 1456 356 1460
rect 350 1455 356 1456
rect 426 1459 432 1460
rect 426 1455 427 1459
rect 431 1455 432 1459
rect 438 1456 439 1460
rect 443 1456 444 1460
rect 438 1455 444 1456
rect 514 1459 520 1460
rect 514 1455 515 1459
rect 519 1455 520 1459
rect 526 1456 527 1460
rect 531 1456 532 1460
rect 526 1455 532 1456
rect 602 1459 608 1460
rect 602 1455 603 1459
rect 607 1455 608 1459
rect 614 1456 615 1460
rect 619 1456 620 1460
rect 614 1455 620 1456
rect 352 1435 354 1455
rect 426 1454 432 1455
rect 440 1435 442 1455
rect 514 1454 520 1455
rect 528 1435 530 1455
rect 602 1454 608 1455
rect 616 1435 618 1455
rect 1568 1435 1570 1466
rect 111 1434 115 1435
rect 111 1429 115 1430
rect 351 1434 355 1435
rect 351 1429 355 1430
rect 439 1434 443 1435
rect 439 1429 443 1430
rect 527 1434 531 1435
rect 527 1429 531 1430
rect 615 1434 619 1435
rect 615 1429 619 1430
rect 663 1434 667 1435
rect 663 1429 667 1430
rect 751 1434 755 1435
rect 751 1429 755 1430
rect 839 1434 843 1435
rect 839 1429 843 1430
rect 927 1434 931 1435
rect 927 1429 931 1430
rect 1567 1434 1571 1435
rect 1567 1429 1571 1430
rect 112 1418 114 1429
rect 662 1428 668 1429
rect 750 1428 756 1429
rect 838 1428 844 1429
rect 926 1428 932 1429
rect 662 1424 663 1428
rect 667 1424 668 1428
rect 662 1423 668 1424
rect 738 1427 744 1428
rect 738 1423 739 1427
rect 743 1423 744 1427
rect 750 1424 751 1428
rect 755 1424 756 1428
rect 750 1423 756 1424
rect 826 1427 832 1428
rect 826 1423 827 1427
rect 831 1423 832 1427
rect 838 1424 839 1428
rect 843 1424 844 1428
rect 838 1423 844 1424
rect 914 1427 920 1428
rect 914 1423 915 1427
rect 919 1423 920 1427
rect 926 1424 927 1428
rect 931 1424 932 1428
rect 926 1423 932 1424
rect 738 1422 744 1423
rect 826 1422 832 1423
rect 914 1422 920 1423
rect 110 1417 116 1418
rect 110 1413 111 1417
rect 115 1413 116 1417
rect 110 1412 116 1413
rect 110 1399 116 1400
rect 110 1395 111 1399
rect 115 1395 116 1399
rect 110 1394 116 1395
rect 112 1359 114 1394
rect 740 1392 742 1422
rect 828 1392 830 1422
rect 850 1411 856 1412
rect 850 1407 851 1411
rect 855 1407 856 1411
rect 850 1406 856 1407
rect 738 1391 744 1392
rect 738 1387 739 1391
rect 743 1387 744 1391
rect 738 1386 744 1387
rect 826 1391 832 1392
rect 826 1387 827 1391
rect 831 1387 832 1391
rect 826 1386 832 1387
rect 662 1382 668 1383
rect 662 1378 663 1382
rect 667 1378 668 1382
rect 662 1377 668 1378
rect 750 1382 756 1383
rect 750 1378 751 1382
rect 755 1378 756 1382
rect 750 1377 756 1378
rect 838 1382 844 1383
rect 838 1378 839 1382
rect 843 1378 844 1382
rect 838 1377 844 1378
rect 664 1359 666 1377
rect 752 1359 754 1377
rect 840 1359 842 1377
rect 111 1358 115 1359
rect 111 1353 115 1354
rect 663 1358 667 1359
rect 663 1353 667 1354
rect 751 1358 755 1359
rect 751 1353 755 1354
rect 815 1358 819 1359
rect 815 1353 819 1354
rect 839 1358 843 1359
rect 839 1353 843 1354
rect 112 1330 114 1353
rect 816 1347 818 1353
rect 852 1348 854 1406
rect 916 1392 918 1422
rect 1568 1418 1570 1429
rect 1566 1417 1572 1418
rect 1566 1413 1567 1417
rect 1571 1413 1572 1417
rect 1566 1412 1572 1413
rect 1566 1399 1572 1400
rect 1566 1395 1567 1399
rect 1571 1395 1572 1399
rect 1566 1394 1572 1395
rect 914 1391 920 1392
rect 914 1387 915 1391
rect 919 1387 920 1391
rect 914 1386 920 1387
rect 926 1382 932 1383
rect 926 1378 927 1382
rect 931 1378 932 1382
rect 926 1377 932 1378
rect 928 1359 930 1377
rect 1568 1359 1570 1394
rect 927 1358 931 1359
rect 927 1353 931 1354
rect 935 1358 939 1359
rect 935 1353 939 1354
rect 1055 1358 1059 1359
rect 1055 1353 1059 1354
rect 1175 1358 1179 1359
rect 1175 1353 1179 1354
rect 1295 1358 1299 1359
rect 1295 1353 1299 1354
rect 1415 1358 1419 1359
rect 1415 1353 1419 1354
rect 1567 1358 1571 1359
rect 1567 1353 1571 1354
rect 850 1347 856 1348
rect 936 1347 938 1353
rect 1056 1347 1058 1353
rect 1176 1347 1178 1353
rect 1296 1347 1298 1353
rect 1416 1347 1418 1353
rect 814 1346 820 1347
rect 814 1342 815 1346
rect 819 1342 820 1346
rect 850 1343 851 1347
rect 855 1343 856 1347
rect 850 1342 856 1343
rect 934 1346 940 1347
rect 934 1342 935 1346
rect 939 1342 940 1346
rect 814 1341 820 1342
rect 934 1341 940 1342
rect 1054 1346 1060 1347
rect 1054 1342 1055 1346
rect 1059 1342 1060 1346
rect 1054 1341 1060 1342
rect 1174 1346 1180 1347
rect 1174 1342 1175 1346
rect 1179 1342 1180 1346
rect 1294 1346 1300 1347
rect 1174 1341 1180 1342
rect 1246 1343 1252 1344
rect 1246 1339 1247 1343
rect 1251 1339 1252 1343
rect 1294 1342 1295 1346
rect 1299 1342 1300 1346
rect 1294 1341 1300 1342
rect 1414 1346 1420 1347
rect 1414 1342 1415 1346
rect 1419 1342 1420 1346
rect 1414 1341 1420 1342
rect 1246 1338 1252 1339
rect 906 1335 912 1336
rect 906 1331 907 1335
rect 911 1331 912 1335
rect 906 1330 912 1331
rect 1026 1335 1032 1336
rect 1026 1331 1027 1335
rect 1031 1331 1032 1335
rect 1026 1330 1032 1331
rect 110 1329 116 1330
rect 110 1325 111 1329
rect 115 1325 116 1329
rect 110 1324 116 1325
rect 110 1311 116 1312
rect 110 1307 111 1311
rect 115 1307 116 1311
rect 110 1306 116 1307
rect 112 1295 114 1306
rect 814 1300 820 1301
rect 908 1300 910 1330
rect 934 1300 940 1301
rect 1028 1300 1030 1330
rect 1054 1300 1060 1301
rect 1174 1300 1180 1301
rect 814 1296 815 1300
rect 819 1296 820 1300
rect 814 1295 820 1296
rect 906 1299 912 1300
rect 906 1295 907 1299
rect 911 1295 912 1299
rect 934 1296 935 1300
rect 939 1296 940 1300
rect 934 1295 940 1296
rect 1026 1299 1032 1300
rect 1026 1295 1027 1299
rect 1031 1295 1032 1299
rect 1054 1296 1055 1300
rect 1059 1296 1060 1300
rect 1054 1295 1060 1296
rect 1086 1299 1092 1300
rect 1086 1295 1087 1299
rect 1091 1295 1092 1299
rect 1174 1296 1175 1300
rect 1179 1296 1180 1300
rect 1174 1295 1180 1296
rect 111 1294 115 1295
rect 111 1289 115 1290
rect 543 1294 547 1295
rect 543 1289 547 1290
rect 695 1294 699 1295
rect 695 1289 699 1290
rect 815 1294 819 1295
rect 815 1289 819 1290
rect 863 1294 867 1295
rect 906 1294 912 1295
rect 935 1294 939 1295
rect 1026 1294 1032 1295
rect 1039 1294 1043 1295
rect 863 1289 867 1290
rect 935 1289 939 1290
rect 1039 1289 1043 1290
rect 1055 1294 1059 1295
rect 1086 1294 1092 1295
rect 1175 1294 1179 1295
rect 1055 1289 1059 1290
rect 112 1278 114 1289
rect 542 1288 548 1289
rect 694 1288 700 1289
rect 542 1284 543 1288
rect 547 1284 548 1288
rect 542 1283 548 1284
rect 626 1287 632 1288
rect 626 1283 627 1287
rect 631 1283 632 1287
rect 694 1284 695 1288
rect 699 1284 700 1288
rect 694 1283 700 1284
rect 862 1288 868 1289
rect 1038 1288 1044 1289
rect 862 1284 863 1288
rect 867 1284 868 1288
rect 862 1283 868 1284
rect 926 1287 932 1288
rect 926 1283 927 1287
rect 931 1283 932 1287
rect 1038 1284 1039 1288
rect 1043 1284 1044 1288
rect 1038 1283 1044 1284
rect 626 1282 632 1283
rect 926 1282 932 1283
rect 110 1277 116 1278
rect 110 1273 111 1277
rect 115 1273 116 1277
rect 110 1272 116 1273
rect 110 1259 116 1260
rect 110 1255 111 1259
rect 115 1255 116 1259
rect 110 1254 116 1255
rect 112 1211 114 1254
rect 628 1252 630 1282
rect 686 1271 692 1272
rect 686 1267 687 1271
rect 691 1267 692 1271
rect 686 1266 692 1267
rect 626 1251 632 1252
rect 626 1247 627 1251
rect 631 1247 632 1251
rect 626 1246 632 1247
rect 688 1244 690 1266
rect 686 1243 692 1244
rect 542 1242 548 1243
rect 542 1238 543 1242
rect 547 1238 548 1242
rect 686 1239 687 1243
rect 691 1239 692 1243
rect 686 1238 692 1239
rect 694 1242 700 1243
rect 694 1238 695 1242
rect 699 1238 700 1242
rect 542 1237 548 1238
rect 694 1237 700 1238
rect 862 1242 868 1243
rect 862 1238 863 1242
rect 867 1238 868 1242
rect 862 1237 868 1238
rect 544 1211 546 1237
rect 696 1211 698 1237
rect 864 1211 866 1237
rect 111 1210 115 1211
rect 111 1205 115 1206
rect 199 1210 203 1211
rect 199 1205 203 1206
rect 415 1210 419 1211
rect 415 1205 419 1206
rect 543 1210 547 1211
rect 543 1205 547 1206
rect 647 1210 651 1211
rect 647 1205 651 1206
rect 695 1210 699 1211
rect 695 1205 699 1206
rect 863 1210 867 1211
rect 863 1205 867 1206
rect 895 1210 899 1211
rect 895 1205 899 1206
rect 112 1182 114 1205
rect 200 1199 202 1205
rect 416 1199 418 1205
rect 648 1199 650 1205
rect 896 1199 898 1205
rect 928 1200 930 1282
rect 1088 1244 1090 1294
rect 1175 1289 1179 1290
rect 1215 1294 1219 1295
rect 1215 1289 1219 1290
rect 1214 1288 1220 1289
rect 1248 1288 1250 1338
rect 1266 1335 1272 1336
rect 1266 1331 1267 1335
rect 1271 1331 1272 1335
rect 1266 1330 1272 1331
rect 1386 1335 1392 1336
rect 1386 1331 1387 1335
rect 1391 1331 1392 1335
rect 1386 1330 1392 1331
rect 1568 1330 1570 1353
rect 1268 1300 1270 1330
rect 1294 1300 1300 1301
rect 1388 1300 1390 1330
rect 1566 1329 1572 1330
rect 1566 1325 1567 1329
rect 1571 1325 1572 1329
rect 1566 1324 1572 1325
rect 1566 1311 1572 1312
rect 1566 1307 1567 1311
rect 1571 1307 1572 1311
rect 1566 1306 1572 1307
rect 1414 1300 1420 1301
rect 1266 1299 1272 1300
rect 1266 1295 1267 1299
rect 1271 1295 1272 1299
rect 1294 1296 1295 1300
rect 1299 1296 1300 1300
rect 1294 1295 1300 1296
rect 1386 1299 1392 1300
rect 1386 1295 1387 1299
rect 1391 1295 1392 1299
rect 1414 1296 1415 1300
rect 1419 1296 1420 1300
rect 1414 1295 1420 1296
rect 1446 1299 1452 1300
rect 1446 1295 1447 1299
rect 1451 1295 1452 1299
rect 1568 1295 1570 1306
rect 1266 1294 1272 1295
rect 1295 1294 1299 1295
rect 1386 1294 1392 1295
rect 1399 1294 1403 1295
rect 1295 1289 1299 1290
rect 1399 1289 1403 1290
rect 1415 1294 1419 1295
rect 1446 1294 1452 1295
rect 1567 1294 1571 1295
rect 1415 1289 1419 1290
rect 1398 1288 1404 1289
rect 1214 1284 1215 1288
rect 1219 1284 1220 1288
rect 1214 1283 1220 1284
rect 1246 1287 1252 1288
rect 1246 1283 1247 1287
rect 1251 1283 1252 1287
rect 1398 1284 1399 1288
rect 1403 1284 1404 1288
rect 1398 1283 1404 1284
rect 1438 1287 1444 1288
rect 1438 1283 1439 1287
rect 1443 1283 1444 1287
rect 1246 1282 1252 1283
rect 1438 1282 1444 1283
rect 1086 1243 1092 1244
rect 1238 1243 1244 1244
rect 1038 1242 1044 1243
rect 1038 1238 1039 1242
rect 1043 1238 1044 1242
rect 1086 1239 1087 1243
rect 1091 1239 1092 1243
rect 1086 1238 1092 1239
rect 1214 1242 1220 1243
rect 1214 1238 1215 1242
rect 1219 1238 1220 1242
rect 1238 1239 1239 1243
rect 1243 1239 1244 1243
rect 1238 1238 1244 1239
rect 1398 1242 1404 1243
rect 1398 1238 1399 1242
rect 1403 1238 1404 1242
rect 1038 1237 1044 1238
rect 1214 1237 1220 1238
rect 1040 1211 1042 1237
rect 1216 1211 1218 1237
rect 1039 1210 1043 1211
rect 1039 1205 1043 1206
rect 1151 1210 1155 1211
rect 1151 1205 1155 1206
rect 1215 1210 1219 1211
rect 1215 1205 1219 1206
rect 926 1199 932 1200
rect 1152 1199 1154 1205
rect 198 1198 204 1199
rect 198 1194 199 1198
rect 203 1194 204 1198
rect 198 1193 204 1194
rect 414 1198 420 1199
rect 414 1194 415 1198
rect 419 1194 420 1198
rect 414 1193 420 1194
rect 646 1198 652 1199
rect 646 1194 647 1198
rect 651 1194 652 1198
rect 646 1193 652 1194
rect 894 1198 900 1199
rect 894 1194 895 1198
rect 899 1194 900 1198
rect 926 1195 927 1199
rect 931 1195 932 1199
rect 926 1194 932 1195
rect 1150 1198 1156 1199
rect 1150 1194 1151 1198
rect 1155 1194 1156 1198
rect 894 1193 900 1194
rect 1150 1193 1156 1194
rect 1206 1195 1212 1196
rect 1206 1191 1207 1195
rect 1211 1191 1212 1195
rect 1206 1190 1212 1191
rect 430 1187 436 1188
rect 430 1183 431 1187
rect 435 1183 436 1187
rect 430 1182 436 1183
rect 662 1187 668 1188
rect 662 1183 663 1187
rect 667 1183 668 1187
rect 662 1182 668 1183
rect 910 1187 916 1188
rect 910 1183 911 1187
rect 915 1183 916 1187
rect 910 1182 916 1183
rect 110 1181 116 1182
rect 110 1177 111 1181
rect 115 1177 116 1181
rect 110 1176 116 1177
rect 110 1163 116 1164
rect 110 1159 111 1163
rect 115 1159 116 1163
rect 110 1158 116 1159
rect 112 1139 114 1158
rect 198 1152 204 1153
rect 414 1152 420 1153
rect 432 1152 434 1182
rect 646 1152 652 1153
rect 664 1152 666 1182
rect 894 1152 900 1153
rect 912 1152 914 1182
rect 1150 1152 1156 1153
rect 198 1148 199 1152
rect 203 1148 204 1152
rect 198 1147 204 1148
rect 230 1151 236 1152
rect 230 1147 231 1151
rect 235 1147 236 1151
rect 414 1148 415 1152
rect 419 1148 420 1152
rect 414 1147 420 1148
rect 430 1151 436 1152
rect 430 1147 431 1151
rect 435 1147 436 1151
rect 646 1148 647 1152
rect 651 1148 652 1152
rect 646 1147 652 1148
rect 662 1151 668 1152
rect 662 1147 663 1151
rect 667 1147 668 1151
rect 894 1148 895 1152
rect 899 1148 900 1152
rect 894 1147 900 1148
rect 910 1151 916 1152
rect 910 1147 911 1151
rect 915 1147 916 1151
rect 1150 1148 1151 1152
rect 1155 1148 1156 1152
rect 1150 1147 1156 1148
rect 200 1139 202 1147
rect 230 1146 236 1147
rect 111 1138 115 1139
rect 111 1133 115 1134
rect 135 1138 139 1139
rect 135 1133 139 1134
rect 199 1138 203 1139
rect 199 1133 203 1134
rect 112 1122 114 1133
rect 134 1132 140 1133
rect 134 1128 135 1132
rect 139 1128 140 1132
rect 134 1127 140 1128
rect 110 1121 116 1122
rect 110 1117 111 1121
rect 115 1117 116 1121
rect 110 1116 116 1117
rect 110 1103 116 1104
rect 110 1099 111 1103
rect 115 1099 116 1103
rect 110 1098 116 1099
rect 112 1071 114 1098
rect 232 1088 234 1146
rect 416 1139 418 1147
rect 430 1146 436 1147
rect 648 1139 650 1147
rect 662 1146 668 1147
rect 896 1139 898 1147
rect 910 1146 916 1147
rect 1152 1139 1154 1147
rect 415 1138 419 1139
rect 415 1133 419 1134
rect 559 1138 563 1139
rect 559 1133 563 1134
rect 647 1138 651 1139
rect 647 1133 651 1134
rect 895 1138 899 1139
rect 895 1133 899 1134
rect 991 1138 995 1139
rect 991 1133 995 1134
rect 1151 1138 1155 1139
rect 1151 1133 1155 1134
rect 558 1132 564 1133
rect 990 1132 996 1133
rect 378 1131 384 1132
rect 378 1127 379 1131
rect 383 1127 384 1131
rect 558 1128 559 1132
rect 563 1128 564 1132
rect 558 1127 564 1128
rect 750 1131 756 1132
rect 750 1127 751 1131
rect 755 1127 756 1131
rect 990 1128 991 1132
rect 995 1128 996 1132
rect 990 1127 996 1128
rect 1058 1131 1064 1132
rect 1058 1127 1059 1131
rect 1063 1127 1064 1131
rect 378 1126 384 1127
rect 750 1126 756 1127
rect 1058 1126 1064 1127
rect 380 1096 382 1126
rect 752 1096 754 1126
rect 378 1095 384 1096
rect 378 1091 379 1095
rect 383 1091 384 1095
rect 750 1095 756 1096
rect 378 1090 384 1091
rect 618 1091 624 1092
rect 230 1087 236 1088
rect 618 1087 619 1091
rect 623 1087 624 1091
rect 750 1091 751 1095
rect 755 1091 756 1095
rect 750 1090 756 1091
rect 134 1086 140 1087
rect 134 1082 135 1086
rect 139 1082 140 1086
rect 230 1083 231 1087
rect 235 1083 236 1087
rect 230 1082 236 1083
rect 558 1086 564 1087
rect 618 1086 624 1087
rect 990 1086 996 1087
rect 558 1082 559 1086
rect 563 1082 564 1086
rect 134 1081 140 1082
rect 558 1081 564 1082
rect 136 1071 138 1081
rect 560 1071 562 1081
rect 111 1070 115 1071
rect 111 1065 115 1066
rect 135 1070 139 1071
rect 135 1065 139 1066
rect 239 1070 243 1071
rect 239 1065 243 1066
rect 559 1070 563 1071
rect 559 1065 563 1066
rect 112 1042 114 1065
rect 240 1059 242 1065
rect 620 1060 622 1086
rect 990 1082 991 1086
rect 995 1082 996 1086
rect 990 1081 996 1082
rect 992 1071 994 1081
rect 1046 1079 1052 1080
rect 1046 1075 1047 1079
rect 1051 1075 1052 1079
rect 1046 1074 1052 1075
rect 631 1070 635 1071
rect 631 1065 635 1066
rect 991 1070 995 1071
rect 991 1065 995 1066
rect 1031 1070 1035 1071
rect 1031 1065 1035 1066
rect 618 1059 624 1060
rect 632 1059 634 1065
rect 1032 1059 1034 1065
rect 238 1058 244 1059
rect 238 1054 239 1058
rect 243 1054 244 1058
rect 618 1055 619 1059
rect 623 1055 624 1059
rect 618 1054 624 1055
rect 630 1058 636 1059
rect 630 1054 631 1058
rect 635 1054 636 1058
rect 238 1053 244 1054
rect 630 1053 636 1054
rect 1030 1058 1036 1059
rect 1030 1054 1031 1058
rect 1035 1054 1036 1058
rect 1030 1053 1036 1054
rect 498 1047 504 1048
rect 498 1043 499 1047
rect 503 1043 504 1047
rect 498 1042 504 1043
rect 110 1041 116 1042
rect 110 1037 111 1041
rect 115 1037 116 1041
rect 110 1036 116 1037
rect 110 1023 116 1024
rect 110 1019 111 1023
rect 115 1019 116 1023
rect 110 1018 116 1019
rect 112 1007 114 1018
rect 238 1012 244 1013
rect 500 1012 502 1042
rect 630 1012 636 1013
rect 1030 1012 1036 1013
rect 1048 1012 1050 1074
rect 1060 1060 1062 1126
rect 1058 1059 1064 1060
rect 1058 1055 1059 1059
rect 1063 1055 1064 1059
rect 1058 1054 1064 1055
rect 238 1008 239 1012
rect 243 1008 244 1012
rect 238 1007 244 1008
rect 498 1011 504 1012
rect 498 1007 499 1011
rect 503 1007 504 1011
rect 630 1008 631 1012
rect 635 1008 636 1012
rect 630 1007 636 1008
rect 686 1011 692 1012
rect 686 1007 687 1011
rect 691 1007 692 1011
rect 1030 1008 1031 1012
rect 1035 1008 1036 1012
rect 1030 1007 1036 1008
rect 1046 1011 1052 1012
rect 1046 1007 1047 1011
rect 1051 1007 1052 1011
rect 111 1006 115 1007
rect 111 1001 115 1002
rect 239 1006 243 1007
rect 239 1001 243 1002
rect 415 1006 419 1007
rect 498 1006 504 1007
rect 631 1006 635 1007
rect 415 1001 419 1002
rect 631 1001 635 1002
rect 663 1006 667 1007
rect 686 1006 692 1007
rect 919 1006 923 1007
rect 663 1001 667 1002
rect 112 990 114 1001
rect 414 1000 420 1001
rect 662 1000 668 1001
rect 414 996 415 1000
rect 419 996 420 1000
rect 414 995 420 996
rect 566 999 572 1000
rect 566 995 567 999
rect 571 995 572 999
rect 662 996 663 1000
rect 667 996 668 1000
rect 662 995 668 996
rect 566 994 572 995
rect 110 989 116 990
rect 110 985 111 989
rect 115 985 116 989
rect 110 984 116 985
rect 110 971 116 972
rect 110 967 111 971
rect 115 967 116 971
rect 110 966 116 967
rect 112 927 114 966
rect 414 954 420 955
rect 414 950 415 954
rect 419 950 420 954
rect 414 949 420 950
rect 416 927 418 949
rect 111 926 115 927
rect 111 921 115 922
rect 415 926 419 927
rect 415 921 419 922
rect 543 926 547 927
rect 543 921 547 922
rect 112 898 114 921
rect 544 915 546 921
rect 568 916 570 994
rect 688 956 690 1006
rect 919 1001 923 1002
rect 1031 1006 1035 1007
rect 1046 1006 1052 1007
rect 1175 1006 1179 1007
rect 1031 1001 1035 1002
rect 1175 1001 1179 1002
rect 918 1000 924 1001
rect 1174 1000 1180 1001
rect 1208 1000 1210 1190
rect 1240 1152 1242 1238
rect 1398 1237 1404 1238
rect 1400 1211 1402 1237
rect 1399 1210 1403 1211
rect 1399 1205 1403 1206
rect 1415 1210 1419 1211
rect 1415 1205 1419 1206
rect 1416 1199 1418 1205
rect 1440 1200 1442 1282
rect 1448 1244 1450 1294
rect 1567 1289 1571 1290
rect 1568 1278 1570 1289
rect 1566 1277 1572 1278
rect 1566 1273 1567 1277
rect 1571 1273 1572 1277
rect 1566 1272 1572 1273
rect 1566 1259 1572 1260
rect 1566 1255 1567 1259
rect 1571 1255 1572 1259
rect 1566 1254 1572 1255
rect 1446 1243 1452 1244
rect 1446 1239 1447 1243
rect 1451 1239 1452 1243
rect 1446 1238 1452 1239
rect 1568 1211 1570 1254
rect 1567 1210 1571 1211
rect 1567 1205 1571 1206
rect 1438 1199 1444 1200
rect 1414 1198 1420 1199
rect 1414 1194 1415 1198
rect 1419 1194 1420 1198
rect 1438 1195 1439 1199
rect 1443 1195 1444 1199
rect 1438 1194 1444 1195
rect 1414 1193 1420 1194
rect 1568 1182 1570 1205
rect 1566 1181 1572 1182
rect 1566 1177 1567 1181
rect 1571 1177 1572 1181
rect 1566 1176 1572 1177
rect 1566 1163 1572 1164
rect 1566 1159 1567 1163
rect 1571 1159 1572 1163
rect 1566 1158 1572 1159
rect 1414 1152 1420 1153
rect 1238 1151 1244 1152
rect 1238 1147 1239 1151
rect 1243 1147 1244 1151
rect 1414 1148 1415 1152
rect 1419 1148 1420 1152
rect 1414 1147 1420 1148
rect 1446 1151 1452 1152
rect 1446 1147 1447 1151
rect 1451 1147 1452 1151
rect 1238 1146 1244 1147
rect 1416 1139 1418 1147
rect 1446 1146 1452 1147
rect 1415 1138 1419 1139
rect 1415 1133 1419 1134
rect 1423 1138 1427 1139
rect 1423 1133 1427 1134
rect 1422 1132 1428 1133
rect 1422 1128 1423 1132
rect 1427 1128 1428 1132
rect 1422 1127 1428 1128
rect 1448 1092 1450 1146
rect 1568 1139 1570 1158
rect 1567 1138 1571 1139
rect 1567 1133 1571 1134
rect 1462 1131 1468 1132
rect 1462 1127 1463 1131
rect 1467 1127 1468 1131
rect 1462 1126 1468 1127
rect 1446 1091 1452 1092
rect 1446 1087 1447 1091
rect 1451 1087 1452 1091
rect 1422 1086 1428 1087
rect 1446 1086 1452 1087
rect 1422 1082 1423 1086
rect 1427 1082 1428 1086
rect 1422 1081 1428 1082
rect 1424 1071 1426 1081
rect 1423 1070 1427 1071
rect 1423 1065 1427 1066
rect 1431 1070 1435 1071
rect 1431 1065 1435 1066
rect 1432 1059 1434 1065
rect 1464 1060 1466 1126
rect 1568 1122 1570 1133
rect 1566 1121 1572 1122
rect 1566 1117 1567 1121
rect 1571 1117 1572 1121
rect 1566 1116 1572 1117
rect 1566 1103 1572 1104
rect 1566 1099 1567 1103
rect 1571 1099 1572 1103
rect 1566 1098 1572 1099
rect 1568 1071 1570 1098
rect 1567 1070 1571 1071
rect 1567 1065 1571 1066
rect 1462 1059 1468 1060
rect 1430 1058 1436 1059
rect 1430 1054 1431 1058
rect 1435 1054 1436 1058
rect 1462 1055 1463 1059
rect 1467 1055 1468 1059
rect 1462 1054 1468 1055
rect 1430 1053 1436 1054
rect 1568 1042 1570 1065
rect 1566 1041 1572 1042
rect 1566 1037 1567 1041
rect 1571 1037 1572 1041
rect 1566 1036 1572 1037
rect 1566 1023 1572 1024
rect 1566 1019 1567 1023
rect 1571 1019 1572 1023
rect 1566 1018 1572 1019
rect 1430 1012 1436 1013
rect 1430 1008 1431 1012
rect 1435 1008 1436 1012
rect 1430 1007 1436 1008
rect 1462 1011 1468 1012
rect 1462 1007 1463 1011
rect 1467 1007 1468 1011
rect 1568 1007 1570 1018
rect 1431 1006 1435 1007
rect 1431 1001 1435 1002
rect 1439 1006 1443 1007
rect 1462 1006 1468 1007
rect 1567 1006 1571 1007
rect 1439 1001 1443 1002
rect 1438 1000 1444 1001
rect 822 999 828 1000
rect 822 995 823 999
rect 827 995 828 999
rect 918 996 919 1000
rect 923 996 924 1000
rect 918 995 924 996
rect 950 999 956 1000
rect 950 995 951 999
rect 955 995 956 999
rect 1174 996 1175 1000
rect 1179 996 1180 1000
rect 1174 995 1180 996
rect 1206 999 1212 1000
rect 1206 995 1207 999
rect 1211 995 1212 999
rect 1438 996 1439 1000
rect 1443 996 1444 1000
rect 1438 995 1444 996
rect 822 994 828 995
rect 950 994 956 995
rect 1206 994 1212 995
rect 824 964 826 994
rect 822 963 828 964
rect 822 959 823 963
rect 827 959 828 963
rect 822 958 828 959
rect 686 955 692 956
rect 662 954 668 955
rect 662 950 663 954
rect 667 950 668 954
rect 686 951 687 955
rect 691 951 692 955
rect 686 950 692 951
rect 918 954 924 955
rect 918 950 919 954
rect 923 950 924 954
rect 662 949 668 950
rect 918 949 924 950
rect 664 927 666 949
rect 920 927 922 949
rect 952 948 954 994
rect 1464 956 1466 1006
rect 1567 1001 1571 1002
rect 1470 999 1476 1000
rect 1470 995 1471 999
rect 1475 995 1476 999
rect 1470 994 1476 995
rect 1286 955 1292 956
rect 1462 955 1468 956
rect 1174 954 1180 955
rect 1174 950 1175 954
rect 1179 950 1180 954
rect 1286 951 1287 955
rect 1291 951 1292 955
rect 1286 950 1292 951
rect 1438 954 1444 955
rect 1438 950 1439 954
rect 1443 950 1444 954
rect 1462 951 1463 955
rect 1467 951 1468 955
rect 1462 950 1468 951
rect 1174 949 1180 950
rect 950 947 956 948
rect 950 943 951 947
rect 955 943 956 947
rect 950 942 956 943
rect 1176 927 1178 949
rect 663 926 667 927
rect 663 921 667 922
rect 751 926 755 927
rect 751 921 755 922
rect 919 926 923 927
rect 919 921 923 922
rect 975 926 979 927
rect 975 921 979 922
rect 1175 926 1179 927
rect 1175 921 1179 922
rect 1207 926 1211 927
rect 1207 921 1211 922
rect 566 915 572 916
rect 752 915 754 921
rect 976 915 978 921
rect 1208 915 1210 921
rect 542 914 548 915
rect 542 910 543 914
rect 547 910 548 914
rect 566 911 567 915
rect 571 911 572 915
rect 566 910 572 911
rect 750 914 756 915
rect 750 910 751 914
rect 755 910 756 914
rect 542 909 548 910
rect 750 909 756 910
rect 974 914 980 915
rect 974 910 975 914
rect 979 910 980 914
rect 974 909 980 910
rect 1206 914 1212 915
rect 1206 910 1207 914
rect 1211 910 1212 914
rect 1206 909 1212 910
rect 690 903 696 904
rect 690 899 691 903
rect 695 899 696 903
rect 690 898 696 899
rect 894 903 900 904
rect 894 899 895 903
rect 899 899 900 903
rect 894 898 900 899
rect 1122 903 1128 904
rect 1122 899 1123 903
rect 1127 899 1128 903
rect 1122 898 1128 899
rect 110 897 116 898
rect 110 893 111 897
rect 115 893 116 897
rect 110 892 116 893
rect 110 879 116 880
rect 110 875 111 879
rect 115 875 116 879
rect 110 874 116 875
rect 112 855 114 874
rect 542 868 548 869
rect 692 868 694 898
rect 750 868 756 869
rect 896 868 898 898
rect 974 868 980 869
rect 1124 868 1126 898
rect 1206 868 1212 869
rect 542 864 543 868
rect 547 864 548 868
rect 542 863 548 864
rect 690 867 696 868
rect 690 863 691 867
rect 695 863 696 867
rect 750 864 751 868
rect 755 864 756 868
rect 750 863 756 864
rect 894 867 900 868
rect 894 863 895 867
rect 899 863 900 867
rect 974 864 975 868
rect 979 864 980 868
rect 974 863 980 864
rect 1122 867 1128 868
rect 1122 863 1123 867
rect 1127 863 1128 867
rect 1206 864 1207 868
rect 1211 864 1212 868
rect 1206 863 1212 864
rect 1238 867 1244 868
rect 1238 863 1239 867
rect 1243 863 1244 867
rect 544 855 546 863
rect 690 862 696 863
rect 752 855 754 863
rect 894 862 900 863
rect 976 855 978 863
rect 1122 862 1128 863
rect 1208 855 1210 863
rect 1238 862 1244 863
rect 111 854 115 855
rect 111 849 115 850
rect 543 854 547 855
rect 543 849 547 850
rect 751 854 755 855
rect 751 849 755 850
rect 775 854 779 855
rect 775 849 779 850
rect 927 854 931 855
rect 927 849 931 850
rect 975 854 979 855
rect 975 849 979 850
rect 1087 854 1091 855
rect 1087 849 1091 850
rect 1207 854 1211 855
rect 1207 849 1211 850
rect 112 838 114 849
rect 774 848 780 849
rect 926 848 932 849
rect 774 844 775 848
rect 779 844 780 848
rect 774 843 780 844
rect 878 847 884 848
rect 878 843 879 847
rect 883 843 884 847
rect 926 844 927 848
rect 931 844 932 848
rect 926 843 932 844
rect 1086 848 1092 849
rect 1086 844 1087 848
rect 1091 844 1092 848
rect 1086 843 1092 844
rect 878 842 884 843
rect 110 837 116 838
rect 110 833 111 837
rect 115 833 116 837
rect 110 832 116 833
rect 810 831 816 832
rect 810 827 811 831
rect 815 827 816 831
rect 810 826 816 827
rect 110 819 116 820
rect 110 815 111 819
rect 115 815 116 819
rect 110 814 116 815
rect 112 775 114 814
rect 812 804 814 826
rect 810 803 816 804
rect 774 802 780 803
rect 774 798 775 802
rect 779 798 780 802
rect 810 799 811 803
rect 815 799 816 803
rect 810 798 816 799
rect 774 797 780 798
rect 776 775 778 797
rect 111 774 115 775
rect 111 769 115 770
rect 775 774 779 775
rect 775 769 779 770
rect 855 774 859 775
rect 855 769 859 770
rect 112 746 114 769
rect 856 763 858 769
rect 880 764 882 842
rect 978 831 984 832
rect 978 827 979 831
rect 983 827 984 831
rect 978 826 984 827
rect 980 804 982 826
rect 1240 804 1242 862
rect 1255 854 1259 855
rect 1255 849 1259 850
rect 1254 848 1260 849
rect 1288 848 1290 950
rect 1438 949 1444 950
rect 1440 927 1442 949
rect 1439 926 1443 927
rect 1439 921 1443 922
rect 1440 915 1442 921
rect 1472 916 1474 994
rect 1568 990 1570 1001
rect 1566 989 1572 990
rect 1566 985 1567 989
rect 1571 985 1572 989
rect 1566 984 1572 985
rect 1566 971 1572 972
rect 1566 967 1567 971
rect 1571 967 1572 971
rect 1566 966 1572 967
rect 1568 927 1570 966
rect 1567 926 1571 927
rect 1567 921 1571 922
rect 1470 915 1476 916
rect 1438 914 1444 915
rect 1438 910 1439 914
rect 1443 910 1444 914
rect 1470 911 1471 915
rect 1475 911 1476 915
rect 1470 910 1476 911
rect 1438 909 1444 910
rect 1568 898 1570 921
rect 1566 897 1572 898
rect 1566 893 1567 897
rect 1571 893 1572 897
rect 1566 892 1572 893
rect 1566 879 1572 880
rect 1566 875 1567 879
rect 1571 875 1572 879
rect 1566 874 1572 875
rect 1438 868 1444 869
rect 1438 864 1439 868
rect 1443 864 1444 868
rect 1438 863 1444 864
rect 1470 867 1476 868
rect 1470 863 1471 867
rect 1475 863 1476 867
rect 1440 855 1442 863
rect 1470 862 1476 863
rect 1423 854 1427 855
rect 1423 849 1427 850
rect 1439 854 1443 855
rect 1439 849 1443 850
rect 1422 848 1428 849
rect 1254 844 1255 848
rect 1259 844 1260 848
rect 1254 843 1260 844
rect 1286 847 1292 848
rect 1286 843 1287 847
rect 1291 843 1292 847
rect 1422 844 1423 848
rect 1427 844 1428 848
rect 1422 843 1428 844
rect 1454 847 1460 848
rect 1454 843 1455 847
rect 1459 843 1460 847
rect 1286 842 1292 843
rect 1454 842 1460 843
rect 978 803 984 804
rect 1238 803 1244 804
rect 1286 803 1292 804
rect 926 802 932 803
rect 926 798 927 802
rect 931 798 932 802
rect 978 799 979 803
rect 983 799 984 803
rect 978 798 984 799
rect 1086 802 1092 803
rect 1086 798 1087 802
rect 1091 798 1092 802
rect 1238 799 1239 803
rect 1243 799 1244 803
rect 1238 798 1244 799
rect 1254 802 1260 803
rect 1254 798 1255 802
rect 1259 798 1260 802
rect 1286 799 1287 803
rect 1291 799 1292 803
rect 1286 798 1292 799
rect 1422 802 1428 803
rect 1422 798 1423 802
rect 1427 798 1428 802
rect 926 797 932 798
rect 1086 797 1092 798
rect 1254 797 1260 798
rect 928 775 930 797
rect 1088 775 1090 797
rect 1256 775 1258 797
rect 927 774 931 775
rect 927 769 931 770
rect 975 774 979 775
rect 975 769 979 770
rect 1087 774 1091 775
rect 1087 769 1091 770
rect 1103 774 1107 775
rect 1103 769 1107 770
rect 1239 774 1243 775
rect 1239 769 1243 770
rect 1255 774 1259 775
rect 1255 769 1259 770
rect 878 763 884 764
rect 976 763 978 769
rect 1104 763 1106 769
rect 1240 763 1242 769
rect 854 762 860 763
rect 854 758 855 762
rect 859 758 860 762
rect 878 759 879 763
rect 883 759 884 763
rect 878 758 884 759
rect 974 762 980 763
rect 974 758 975 762
rect 979 758 980 762
rect 854 757 860 758
rect 974 757 980 758
rect 1102 762 1108 763
rect 1102 758 1103 762
rect 1107 758 1108 762
rect 1102 757 1108 758
rect 1238 762 1244 763
rect 1238 758 1239 762
rect 1243 758 1244 762
rect 1238 757 1244 758
rect 1262 759 1268 760
rect 1262 755 1263 759
rect 1267 755 1268 759
rect 1262 754 1268 755
rect 946 751 952 752
rect 946 747 947 751
rect 951 747 952 751
rect 946 746 952 747
rect 1070 751 1076 752
rect 1070 747 1071 751
rect 1075 747 1076 751
rect 1070 746 1076 747
rect 110 745 116 746
rect 110 741 111 745
rect 115 741 116 745
rect 110 740 116 741
rect 110 727 116 728
rect 110 723 111 727
rect 115 723 116 727
rect 110 722 116 723
rect 112 703 114 722
rect 854 716 860 717
rect 948 716 950 746
rect 974 716 980 717
rect 1072 716 1074 746
rect 1102 716 1108 717
rect 1238 716 1244 717
rect 854 712 855 716
rect 859 712 860 716
rect 854 711 860 712
rect 946 715 952 716
rect 946 711 947 715
rect 951 711 952 715
rect 974 712 975 716
rect 979 712 980 716
rect 974 711 980 712
rect 1070 715 1076 716
rect 1070 711 1071 715
rect 1075 711 1076 715
rect 1102 712 1103 716
rect 1107 712 1108 716
rect 1102 711 1108 712
rect 1158 715 1164 716
rect 1158 711 1159 715
rect 1163 711 1164 715
rect 1238 712 1239 716
rect 1243 712 1244 716
rect 1238 711 1244 712
rect 856 703 858 711
rect 946 710 952 711
rect 976 703 978 711
rect 1070 710 1076 711
rect 1104 703 1106 711
rect 1158 710 1164 711
rect 111 702 115 703
rect 111 697 115 698
rect 735 702 739 703
rect 735 697 739 698
rect 855 702 859 703
rect 855 697 859 698
rect 935 702 939 703
rect 935 697 939 698
rect 975 702 979 703
rect 975 697 979 698
rect 1103 702 1107 703
rect 1103 697 1107 698
rect 1135 702 1139 703
rect 1135 697 1139 698
rect 112 686 114 697
rect 734 696 740 697
rect 934 696 940 697
rect 734 692 735 696
rect 739 692 740 696
rect 734 691 740 692
rect 870 695 876 696
rect 870 691 871 695
rect 875 691 876 695
rect 934 692 935 696
rect 939 692 940 696
rect 934 691 940 692
rect 1134 696 1140 697
rect 1134 692 1135 696
rect 1139 692 1140 696
rect 1134 691 1140 692
rect 870 690 876 691
rect 110 685 116 686
rect 110 681 111 685
rect 115 681 116 685
rect 110 680 116 681
rect 110 667 116 668
rect 110 663 111 667
rect 115 663 116 667
rect 110 662 116 663
rect 112 639 114 662
rect 734 650 740 651
rect 734 646 735 650
rect 739 646 740 650
rect 734 645 740 646
rect 736 639 738 645
rect 111 638 115 639
rect 111 633 115 634
rect 607 638 611 639
rect 607 633 611 634
rect 735 638 739 639
rect 735 633 739 634
rect 847 638 851 639
rect 847 633 851 634
rect 112 610 114 633
rect 608 627 610 633
rect 848 627 850 633
rect 872 628 874 690
rect 986 679 992 680
rect 986 675 987 679
rect 991 675 992 679
rect 986 674 992 675
rect 988 652 990 674
rect 1160 673 1162 710
rect 1240 703 1242 711
rect 1239 702 1243 703
rect 1239 697 1243 698
rect 1160 671 1170 673
rect 1168 652 1170 671
rect 986 651 992 652
rect 1166 651 1172 652
rect 934 650 940 651
rect 934 646 935 650
rect 939 646 940 650
rect 986 647 987 651
rect 991 647 992 651
rect 986 646 992 647
rect 1134 650 1140 651
rect 1134 646 1135 650
rect 1139 646 1140 650
rect 1166 647 1167 651
rect 1171 647 1172 651
rect 1166 646 1172 647
rect 934 645 940 646
rect 1134 645 1140 646
rect 936 639 938 645
rect 1136 639 1138 645
rect 935 638 939 639
rect 935 633 939 634
rect 1087 638 1091 639
rect 1087 633 1091 634
rect 1135 638 1139 639
rect 1135 633 1139 634
rect 870 627 876 628
rect 1088 627 1090 633
rect 606 626 612 627
rect 606 622 607 626
rect 611 622 612 626
rect 606 621 612 622
rect 846 626 852 627
rect 846 622 847 626
rect 851 622 852 626
rect 870 623 871 627
rect 875 623 876 627
rect 870 622 876 623
rect 1086 626 1092 627
rect 1086 622 1087 626
rect 1091 622 1092 626
rect 846 621 852 622
rect 1086 621 1092 622
rect 1118 623 1124 624
rect 1118 619 1119 623
rect 1123 619 1124 623
rect 1118 618 1124 619
rect 862 615 868 616
rect 862 611 863 615
rect 867 611 868 615
rect 862 610 868 611
rect 110 609 116 610
rect 110 605 111 609
rect 115 605 116 609
rect 110 604 116 605
rect 110 591 116 592
rect 110 587 111 591
rect 115 587 116 591
rect 110 586 116 587
rect 112 567 114 586
rect 606 580 612 581
rect 606 576 607 580
rect 611 576 612 580
rect 606 575 612 576
rect 846 580 852 581
rect 864 580 866 610
rect 1086 580 1092 581
rect 846 576 847 580
rect 851 576 852 580
rect 846 575 852 576
rect 862 579 868 580
rect 862 575 863 579
rect 867 575 868 579
rect 1086 576 1087 580
rect 1091 576 1092 580
rect 1086 575 1092 576
rect 390 571 396 572
rect 390 567 391 571
rect 395 567 396 571
rect 608 567 610 575
rect 848 567 850 575
rect 862 574 868 575
rect 1088 567 1090 575
rect 111 566 115 567
rect 111 561 115 562
rect 359 566 363 567
rect 390 566 396 567
rect 591 566 595 567
rect 359 561 363 562
rect 112 550 114 561
rect 358 560 364 561
rect 358 556 359 560
rect 363 556 364 560
rect 358 555 364 556
rect 110 549 116 550
rect 110 545 111 549
rect 115 545 116 549
rect 110 544 116 545
rect 110 531 116 532
rect 110 527 111 531
rect 115 527 116 531
rect 110 526 116 527
rect 112 487 114 526
rect 392 516 394 566
rect 591 561 595 562
rect 607 566 611 567
rect 607 561 611 562
rect 831 566 835 567
rect 831 561 835 562
rect 847 566 851 567
rect 847 561 851 562
rect 1079 566 1083 567
rect 1079 561 1083 562
rect 1087 566 1091 567
rect 1087 561 1091 562
rect 590 560 596 561
rect 506 559 512 560
rect 506 555 507 559
rect 511 555 512 559
rect 590 556 591 560
rect 595 556 596 560
rect 590 555 596 556
rect 830 560 836 561
rect 1078 560 1084 561
rect 1120 560 1122 618
rect 1264 580 1266 754
rect 1288 716 1290 798
rect 1422 797 1428 798
rect 1424 775 1426 797
rect 1375 774 1379 775
rect 1375 769 1379 770
rect 1423 774 1427 775
rect 1423 769 1427 770
rect 1376 763 1378 769
rect 1456 764 1458 842
rect 1472 804 1474 862
rect 1568 855 1570 874
rect 1567 854 1571 855
rect 1567 849 1571 850
rect 1568 838 1570 849
rect 1566 837 1572 838
rect 1566 833 1567 837
rect 1571 833 1572 837
rect 1566 832 1572 833
rect 1566 819 1572 820
rect 1566 815 1567 819
rect 1571 815 1572 819
rect 1566 814 1572 815
rect 1470 803 1476 804
rect 1470 799 1471 803
rect 1475 799 1476 803
rect 1470 798 1476 799
rect 1568 775 1570 814
rect 1567 774 1571 775
rect 1567 769 1571 770
rect 1454 763 1460 764
rect 1374 762 1380 763
rect 1374 758 1375 762
rect 1379 758 1380 762
rect 1454 759 1455 763
rect 1459 759 1460 763
rect 1454 758 1460 759
rect 1374 757 1380 758
rect 1568 746 1570 769
rect 1566 745 1572 746
rect 1566 741 1567 745
rect 1571 741 1572 745
rect 1566 740 1572 741
rect 1566 727 1572 728
rect 1566 723 1567 727
rect 1571 723 1572 727
rect 1566 722 1572 723
rect 1374 716 1380 717
rect 1286 715 1292 716
rect 1286 711 1287 715
rect 1291 711 1292 715
rect 1374 712 1375 716
rect 1379 712 1380 716
rect 1374 711 1380 712
rect 1406 715 1412 716
rect 1406 711 1407 715
rect 1411 711 1412 715
rect 1286 710 1292 711
rect 1376 703 1378 711
rect 1406 710 1412 711
rect 1343 702 1347 703
rect 1343 697 1347 698
rect 1375 702 1379 703
rect 1375 697 1379 698
rect 1342 696 1348 697
rect 1342 692 1343 696
rect 1347 692 1348 696
rect 1342 691 1348 692
rect 1374 679 1380 680
rect 1374 675 1375 679
rect 1379 675 1380 679
rect 1374 674 1380 675
rect 1342 650 1348 651
rect 1342 646 1343 650
rect 1347 646 1348 650
rect 1342 645 1348 646
rect 1344 639 1346 645
rect 1327 638 1331 639
rect 1327 633 1331 634
rect 1343 638 1347 639
rect 1343 633 1347 634
rect 1328 627 1330 633
rect 1376 628 1378 674
rect 1408 652 1410 710
rect 1568 703 1570 722
rect 1567 702 1571 703
rect 1567 697 1571 698
rect 1568 686 1570 697
rect 1566 685 1572 686
rect 1566 681 1567 685
rect 1571 681 1572 685
rect 1566 680 1572 681
rect 1566 667 1572 668
rect 1566 663 1567 667
rect 1571 663 1572 667
rect 1566 662 1572 663
rect 1406 651 1412 652
rect 1406 647 1407 651
rect 1411 647 1412 651
rect 1406 646 1412 647
rect 1568 639 1570 662
rect 1567 638 1571 639
rect 1567 633 1571 634
rect 1374 627 1380 628
rect 1326 626 1332 627
rect 1326 622 1327 626
rect 1331 622 1332 626
rect 1374 623 1375 627
rect 1379 623 1380 627
rect 1374 622 1380 623
rect 1326 621 1332 622
rect 1568 610 1570 633
rect 1566 609 1572 610
rect 1566 605 1567 609
rect 1571 605 1572 609
rect 1566 604 1572 605
rect 1566 591 1572 592
rect 1566 587 1567 591
rect 1571 587 1572 591
rect 1566 586 1572 587
rect 1326 580 1332 581
rect 1262 579 1268 580
rect 1262 575 1263 579
rect 1267 575 1268 579
rect 1326 576 1327 580
rect 1331 576 1332 580
rect 1326 575 1332 576
rect 1358 579 1364 580
rect 1358 575 1359 579
rect 1363 575 1364 579
rect 1262 574 1268 575
rect 1328 567 1330 575
rect 1358 574 1364 575
rect 1327 566 1331 567
rect 1327 561 1331 562
rect 1326 560 1332 561
rect 830 556 831 560
rect 835 556 836 560
rect 830 555 836 556
rect 862 559 868 560
rect 862 555 863 559
rect 867 555 868 559
rect 1078 556 1079 560
rect 1083 556 1084 560
rect 1078 555 1084 556
rect 1118 559 1124 560
rect 1118 555 1119 559
rect 1123 555 1124 559
rect 1326 556 1327 560
rect 1331 556 1332 560
rect 1326 555 1332 556
rect 506 554 512 555
rect 862 554 868 555
rect 1118 554 1124 555
rect 508 524 510 554
rect 506 523 512 524
rect 506 519 507 523
rect 511 519 512 523
rect 506 518 512 519
rect 390 515 396 516
rect 358 514 364 515
rect 358 510 359 514
rect 363 510 364 514
rect 390 511 391 515
rect 395 511 396 515
rect 390 510 396 511
rect 590 514 596 515
rect 590 510 591 514
rect 595 510 596 514
rect 358 509 364 510
rect 590 509 596 510
rect 830 514 836 515
rect 830 510 831 514
rect 835 510 836 514
rect 830 509 836 510
rect 360 487 362 509
rect 592 487 594 509
rect 832 487 834 509
rect 111 486 115 487
rect 111 481 115 482
rect 151 486 155 487
rect 151 481 155 482
rect 359 486 363 487
rect 359 481 363 482
rect 439 486 443 487
rect 439 481 443 482
rect 591 486 595 487
rect 591 481 595 482
rect 735 486 739 487
rect 735 481 739 482
rect 831 486 835 487
rect 831 481 835 482
rect 112 458 114 481
rect 152 475 154 481
rect 440 475 442 481
rect 736 475 738 481
rect 864 476 866 554
rect 1360 516 1362 574
rect 1568 567 1570 586
rect 1567 566 1571 567
rect 1567 561 1571 562
rect 1374 559 1380 560
rect 1374 555 1375 559
rect 1379 555 1380 559
rect 1374 554 1380 555
rect 1106 515 1112 516
rect 1358 515 1364 516
rect 1078 514 1084 515
rect 1078 510 1079 514
rect 1083 510 1084 514
rect 1106 511 1107 515
rect 1111 511 1112 515
rect 1106 510 1112 511
rect 1326 514 1332 515
rect 1326 510 1327 514
rect 1331 510 1332 514
rect 1358 511 1359 515
rect 1363 511 1364 515
rect 1358 510 1364 511
rect 1078 509 1084 510
rect 1080 487 1082 509
rect 1039 486 1043 487
rect 1039 481 1043 482
rect 1079 486 1083 487
rect 1079 481 1083 482
rect 862 475 868 476
rect 1040 475 1042 481
rect 150 474 156 475
rect 150 470 151 474
rect 155 470 156 474
rect 150 469 156 470
rect 438 474 444 475
rect 438 470 439 474
rect 443 470 444 474
rect 438 469 444 470
rect 734 474 740 475
rect 734 470 735 474
rect 739 470 740 474
rect 862 471 863 475
rect 867 471 868 475
rect 862 470 868 471
rect 1038 474 1044 475
rect 1038 470 1039 474
rect 1043 470 1044 474
rect 734 469 740 470
rect 1038 469 1044 470
rect 1070 471 1076 472
rect 1070 467 1071 471
rect 1075 467 1076 471
rect 1070 466 1076 467
rect 454 463 460 464
rect 454 459 455 463
rect 459 459 460 463
rect 454 458 460 459
rect 750 463 756 464
rect 750 459 751 463
rect 755 459 756 463
rect 750 458 756 459
rect 110 457 116 458
rect 110 453 111 457
rect 115 453 116 457
rect 110 452 116 453
rect 110 439 116 440
rect 110 435 111 439
rect 115 435 116 439
rect 110 434 116 435
rect 112 411 114 434
rect 150 428 156 429
rect 438 428 444 429
rect 456 428 458 458
rect 734 428 740 429
rect 752 428 754 458
rect 1038 428 1044 429
rect 150 424 151 428
rect 155 424 156 428
rect 150 423 156 424
rect 206 427 212 428
rect 206 423 207 427
rect 211 423 212 427
rect 438 424 439 428
rect 443 424 444 428
rect 438 423 444 424
rect 454 427 460 428
rect 454 423 455 427
rect 459 423 460 427
rect 734 424 735 428
rect 739 424 740 428
rect 734 423 740 424
rect 750 427 756 428
rect 750 423 751 427
rect 755 423 756 427
rect 1038 424 1039 428
rect 1043 424 1044 428
rect 1038 423 1044 424
rect 152 411 154 423
rect 206 422 212 423
rect 111 410 115 411
rect 111 405 115 406
rect 151 410 155 411
rect 151 405 155 406
rect 175 410 179 411
rect 175 405 179 406
rect 112 394 114 405
rect 174 404 180 405
rect 174 400 175 404
rect 179 400 180 404
rect 174 399 180 400
rect 110 393 116 394
rect 110 389 111 393
rect 115 389 116 393
rect 110 388 116 389
rect 110 375 116 376
rect 110 371 111 375
rect 115 371 116 375
rect 110 370 116 371
rect 112 343 114 370
rect 208 360 210 422
rect 440 411 442 423
rect 454 422 460 423
rect 736 411 738 423
rect 750 422 756 423
rect 1040 411 1042 423
rect 439 410 443 411
rect 439 405 443 406
rect 567 410 571 411
rect 567 405 571 406
rect 735 410 739 411
rect 735 405 739 406
rect 967 410 971 411
rect 967 405 971 406
rect 1039 410 1043 411
rect 1039 405 1043 406
rect 566 404 572 405
rect 966 404 972 405
rect 1072 404 1074 466
rect 1108 432 1110 510
rect 1326 509 1332 510
rect 1328 487 1330 509
rect 1327 486 1331 487
rect 1327 481 1331 482
rect 1343 486 1347 487
rect 1343 481 1347 482
rect 1344 475 1346 481
rect 1376 476 1378 554
rect 1568 550 1570 561
rect 1566 549 1572 550
rect 1566 545 1567 549
rect 1571 545 1572 549
rect 1566 544 1572 545
rect 1566 531 1572 532
rect 1566 527 1567 531
rect 1571 527 1572 531
rect 1566 526 1572 527
rect 1568 487 1570 526
rect 1567 486 1571 487
rect 1567 481 1571 482
rect 1374 475 1380 476
rect 1342 474 1348 475
rect 1342 470 1343 474
rect 1347 470 1348 474
rect 1374 471 1375 475
rect 1379 471 1380 475
rect 1374 470 1380 471
rect 1342 469 1348 470
rect 1568 458 1570 481
rect 1566 457 1572 458
rect 1566 453 1567 457
rect 1571 453 1572 457
rect 1566 452 1572 453
rect 1566 439 1572 440
rect 1566 435 1567 439
rect 1571 435 1572 439
rect 1566 434 1572 435
rect 1106 431 1112 432
rect 1106 427 1107 431
rect 1111 427 1112 431
rect 1106 426 1112 427
rect 1342 428 1348 429
rect 1342 424 1343 428
rect 1347 424 1348 428
rect 1342 423 1348 424
rect 1398 427 1404 428
rect 1398 423 1399 427
rect 1403 423 1404 427
rect 1344 411 1346 423
rect 1398 422 1404 423
rect 1343 410 1347 411
rect 1343 405 1347 406
rect 1367 410 1371 411
rect 1367 405 1371 406
rect 1366 404 1372 405
rect 498 403 504 404
rect 498 399 499 403
rect 503 399 504 403
rect 566 400 567 404
rect 571 400 572 404
rect 566 399 572 400
rect 830 403 836 404
rect 830 399 831 403
rect 835 399 836 403
rect 966 400 967 404
rect 971 400 972 404
rect 966 399 972 400
rect 1070 403 1076 404
rect 1070 399 1071 403
rect 1075 399 1076 403
rect 1366 400 1367 404
rect 1371 400 1372 404
rect 1366 399 1372 400
rect 498 398 504 399
rect 830 398 836 399
rect 1070 398 1076 399
rect 500 368 502 398
rect 498 367 504 368
rect 498 363 499 367
rect 503 363 504 367
rect 498 362 504 363
rect 206 359 212 360
rect 174 358 180 359
rect 174 354 175 358
rect 179 354 180 358
rect 206 355 207 359
rect 211 355 212 359
rect 206 354 212 355
rect 566 358 572 359
rect 566 354 567 358
rect 571 354 572 358
rect 174 353 180 354
rect 566 353 572 354
rect 176 343 178 353
rect 568 343 570 353
rect 111 342 115 343
rect 111 337 115 338
rect 175 342 179 343
rect 175 337 179 338
rect 231 342 235 343
rect 231 337 235 338
rect 511 342 515 343
rect 511 337 515 338
rect 567 342 571 343
rect 567 337 571 338
rect 799 342 803 343
rect 799 337 803 338
rect 112 314 114 337
rect 232 331 234 337
rect 512 331 514 337
rect 800 331 802 337
rect 832 332 834 398
rect 1400 360 1402 422
rect 1568 411 1570 434
rect 1567 410 1571 411
rect 1567 405 1571 406
rect 1430 403 1436 404
rect 1430 399 1431 403
rect 1435 399 1436 403
rect 1430 398 1436 399
rect 1126 359 1132 360
rect 1398 359 1404 360
rect 966 358 972 359
rect 966 354 967 358
rect 971 354 972 358
rect 1126 355 1127 359
rect 1131 355 1132 359
rect 1126 354 1132 355
rect 1366 358 1372 359
rect 1366 354 1367 358
rect 1371 354 1372 358
rect 1398 355 1399 359
rect 1403 355 1404 359
rect 1398 354 1404 355
rect 966 353 972 354
rect 968 343 970 353
rect 967 342 971 343
rect 967 337 971 338
rect 1095 342 1099 343
rect 1095 337 1099 338
rect 830 331 836 332
rect 1096 331 1098 337
rect 230 330 236 331
rect 230 326 231 330
rect 235 326 236 330
rect 230 325 236 326
rect 510 330 516 331
rect 510 326 511 330
rect 515 326 516 330
rect 510 325 516 326
rect 798 330 804 331
rect 798 326 799 330
rect 803 326 804 330
rect 830 327 831 331
rect 835 327 836 331
rect 830 326 836 327
rect 1094 330 1100 331
rect 1094 326 1095 330
rect 1099 326 1100 330
rect 798 325 804 326
rect 1094 325 1100 326
rect 526 319 532 320
rect 526 315 527 319
rect 531 315 532 319
rect 526 314 532 315
rect 814 319 820 320
rect 814 315 815 319
rect 819 315 820 319
rect 814 314 820 315
rect 110 313 116 314
rect 110 309 111 313
rect 115 309 116 313
rect 110 308 116 309
rect 110 295 116 296
rect 110 291 111 295
rect 115 291 116 295
rect 110 290 116 291
rect 112 263 114 290
rect 230 284 236 285
rect 510 284 516 285
rect 528 284 530 314
rect 798 284 804 285
rect 816 284 818 314
rect 1094 284 1100 285
rect 1128 284 1130 354
rect 1366 353 1372 354
rect 1368 343 1370 353
rect 1367 342 1371 343
rect 1367 337 1371 338
rect 1399 342 1403 343
rect 1399 337 1403 338
rect 1400 331 1402 337
rect 1432 332 1434 398
rect 1568 394 1570 405
rect 1566 393 1572 394
rect 1566 389 1567 393
rect 1571 389 1572 393
rect 1566 388 1572 389
rect 1566 375 1572 376
rect 1566 371 1567 375
rect 1571 371 1572 375
rect 1566 370 1572 371
rect 1568 343 1570 370
rect 1567 342 1571 343
rect 1567 337 1571 338
rect 1430 331 1436 332
rect 1398 330 1404 331
rect 1398 326 1399 330
rect 1403 326 1404 330
rect 1430 327 1431 331
rect 1435 327 1436 331
rect 1430 326 1436 327
rect 1398 325 1404 326
rect 1568 314 1570 337
rect 1566 313 1572 314
rect 1566 309 1567 313
rect 1571 309 1572 313
rect 1566 308 1572 309
rect 1566 295 1572 296
rect 1566 291 1567 295
rect 1571 291 1572 295
rect 1566 290 1572 291
rect 1398 284 1404 285
rect 230 280 231 284
rect 235 280 236 284
rect 230 279 236 280
rect 446 283 452 284
rect 446 279 447 283
rect 451 279 452 283
rect 510 280 511 284
rect 515 280 516 284
rect 510 279 516 280
rect 526 283 532 284
rect 526 279 527 283
rect 531 279 532 283
rect 798 280 799 284
rect 803 280 804 284
rect 798 279 804 280
rect 814 283 820 284
rect 814 279 815 283
rect 819 279 820 283
rect 1094 280 1095 284
rect 1099 280 1100 284
rect 1094 279 1100 280
rect 1126 283 1132 284
rect 1126 279 1127 283
rect 1131 279 1132 283
rect 1398 280 1399 284
rect 1403 280 1404 284
rect 1398 279 1404 280
rect 1454 283 1460 284
rect 1454 279 1455 283
rect 1459 279 1460 283
rect 232 263 234 279
rect 446 278 452 279
rect 111 262 115 263
rect 111 257 115 258
rect 231 262 235 263
rect 231 257 235 258
rect 423 262 427 263
rect 423 257 427 258
rect 112 246 114 257
rect 422 256 428 257
rect 422 252 423 256
rect 427 252 428 256
rect 422 251 428 252
rect 110 245 116 246
rect 110 241 111 245
rect 115 241 116 245
rect 110 240 116 241
rect 110 227 116 228
rect 110 223 111 227
rect 115 223 116 227
rect 110 222 116 223
rect 112 183 114 222
rect 448 212 450 278
rect 512 263 514 279
rect 526 278 532 279
rect 800 263 802 279
rect 814 278 820 279
rect 1096 263 1098 279
rect 1126 278 1132 279
rect 1400 263 1402 279
rect 1454 278 1460 279
rect 511 262 515 263
rect 511 257 515 258
rect 663 262 667 263
rect 663 257 667 258
rect 799 262 803 263
rect 799 257 803 258
rect 911 262 915 263
rect 911 257 915 258
rect 1095 262 1099 263
rect 1095 257 1099 258
rect 1167 262 1171 263
rect 1167 257 1171 258
rect 1399 262 1403 263
rect 1399 257 1403 258
rect 1431 262 1435 263
rect 1431 257 1435 258
rect 662 256 668 257
rect 566 255 572 256
rect 566 251 567 255
rect 571 251 572 255
rect 662 252 663 256
rect 667 252 668 256
rect 662 251 668 252
rect 910 256 916 257
rect 910 252 911 256
rect 915 252 916 256
rect 910 251 916 252
rect 1166 256 1172 257
rect 1166 252 1167 256
rect 1171 252 1172 256
rect 1166 251 1172 252
rect 1430 256 1436 257
rect 1430 252 1431 256
rect 1435 252 1436 256
rect 1430 251 1436 252
rect 566 250 572 251
rect 568 220 570 250
rect 574 239 580 240
rect 574 235 575 239
rect 579 235 580 239
rect 574 234 580 235
rect 946 239 952 240
rect 946 235 947 239
rect 951 235 952 239
rect 946 234 952 235
rect 566 219 572 220
rect 566 215 567 219
rect 571 215 572 219
rect 566 214 572 215
rect 446 211 452 212
rect 422 210 428 211
rect 422 206 423 210
rect 427 206 428 210
rect 446 207 447 211
rect 451 207 452 211
rect 446 206 452 207
rect 422 205 428 206
rect 424 183 426 205
rect 111 182 115 183
rect 111 177 115 178
rect 423 182 427 183
rect 423 177 427 178
rect 511 182 515 183
rect 511 177 515 178
rect 112 154 114 177
rect 512 171 514 177
rect 576 172 578 234
rect 948 212 950 234
rect 1456 212 1458 278
rect 1568 263 1570 290
rect 1567 262 1571 263
rect 1567 257 1571 258
rect 1498 255 1504 256
rect 1498 251 1499 255
rect 1503 251 1504 255
rect 1498 250 1504 251
rect 946 211 952 212
rect 1198 211 1204 212
rect 1454 211 1460 212
rect 662 210 668 211
rect 662 206 663 210
rect 667 206 668 210
rect 662 205 668 206
rect 910 210 916 211
rect 910 206 911 210
rect 915 206 916 210
rect 946 207 947 211
rect 951 207 952 211
rect 946 206 952 207
rect 1166 210 1172 211
rect 1166 206 1167 210
rect 1171 206 1172 210
rect 1198 207 1199 211
rect 1203 207 1204 211
rect 1198 206 1204 207
rect 1430 210 1436 211
rect 1430 206 1431 210
rect 1435 206 1436 210
rect 1454 207 1455 211
rect 1459 207 1460 211
rect 1454 206 1460 207
rect 910 205 916 206
rect 1166 205 1172 206
rect 664 183 666 205
rect 912 183 914 205
rect 1168 183 1170 205
rect 615 182 619 183
rect 615 177 619 178
rect 663 182 667 183
rect 663 177 667 178
rect 727 182 731 183
rect 727 177 731 178
rect 855 182 859 183
rect 855 177 859 178
rect 911 182 915 183
rect 911 177 915 178
rect 999 182 1003 183
rect 999 177 1003 178
rect 1159 182 1163 183
rect 1159 177 1163 178
rect 1167 182 1171 183
rect 1167 177 1171 178
rect 574 171 580 172
rect 616 171 618 177
rect 728 171 730 177
rect 856 171 858 177
rect 1000 171 1002 177
rect 1160 171 1162 177
rect 510 170 516 171
rect 510 166 511 170
rect 515 166 516 170
rect 574 167 575 171
rect 579 167 580 171
rect 574 166 580 167
rect 614 170 620 171
rect 614 166 615 170
rect 619 166 620 170
rect 510 165 516 166
rect 614 165 620 166
rect 726 170 732 171
rect 726 166 727 170
rect 731 166 732 170
rect 726 165 732 166
rect 854 170 860 171
rect 854 166 855 170
rect 859 166 860 170
rect 854 165 860 166
rect 998 170 1004 171
rect 998 166 999 170
rect 1003 166 1004 170
rect 998 165 1004 166
rect 1158 170 1164 171
rect 1158 166 1159 170
rect 1163 166 1164 170
rect 1158 165 1164 166
rect 594 159 600 160
rect 594 155 595 159
rect 599 155 600 159
rect 594 154 600 155
rect 718 159 724 160
rect 718 155 719 159
rect 723 155 724 159
rect 718 154 724 155
rect 822 159 828 160
rect 822 155 823 159
rect 827 155 828 159
rect 822 154 828 155
rect 958 159 964 160
rect 958 155 959 159
rect 963 155 964 159
rect 958 154 964 155
rect 1110 159 1116 160
rect 1110 155 1111 159
rect 1115 155 1116 159
rect 1110 154 1116 155
rect 110 153 116 154
rect 110 149 111 153
rect 115 149 116 153
rect 110 148 116 149
rect 110 135 116 136
rect 110 131 111 135
rect 115 131 116 135
rect 110 130 116 131
rect 112 119 114 130
rect 510 124 516 125
rect 596 124 598 154
rect 614 124 620 125
rect 720 124 722 154
rect 726 124 732 125
rect 824 124 826 154
rect 854 124 860 125
rect 960 124 962 154
rect 998 124 1004 125
rect 1112 124 1114 154
rect 1158 124 1164 125
rect 1200 124 1202 206
rect 1430 205 1436 206
rect 1432 183 1434 205
rect 1327 182 1331 183
rect 1327 177 1331 178
rect 1431 182 1435 183
rect 1431 177 1435 178
rect 1471 182 1475 183
rect 1471 177 1475 178
rect 1328 171 1330 177
rect 1472 171 1474 177
rect 1500 172 1502 250
rect 1568 246 1570 257
rect 1566 245 1572 246
rect 1566 241 1567 245
rect 1571 241 1572 245
rect 1566 240 1572 241
rect 1566 227 1572 228
rect 1566 223 1567 227
rect 1571 223 1572 227
rect 1566 222 1572 223
rect 1568 183 1570 222
rect 1567 182 1571 183
rect 1567 177 1571 178
rect 1498 171 1504 172
rect 1326 170 1332 171
rect 1326 166 1327 170
rect 1331 166 1332 170
rect 1326 165 1332 166
rect 1470 170 1476 171
rect 1470 166 1471 170
rect 1475 166 1476 170
rect 1498 167 1499 171
rect 1503 167 1504 171
rect 1498 166 1504 167
rect 1470 165 1476 166
rect 1486 159 1492 160
rect 1486 155 1487 159
rect 1491 155 1492 159
rect 1486 154 1492 155
rect 1568 154 1570 177
rect 1326 124 1332 125
rect 510 120 511 124
rect 515 120 516 124
rect 510 119 516 120
rect 594 123 600 124
rect 594 119 595 123
rect 599 119 600 123
rect 614 120 615 124
rect 619 120 620 124
rect 614 119 620 120
rect 718 123 724 124
rect 718 119 719 123
rect 723 119 724 123
rect 726 120 727 124
rect 731 120 732 124
rect 726 119 732 120
rect 822 123 828 124
rect 822 119 823 123
rect 827 119 828 123
rect 854 120 855 124
rect 859 120 860 124
rect 854 119 860 120
rect 958 123 964 124
rect 958 119 959 123
rect 963 119 964 123
rect 998 120 999 124
rect 1003 120 1004 124
rect 998 119 1004 120
rect 1110 123 1116 124
rect 1110 119 1111 123
rect 1115 119 1116 123
rect 1158 120 1159 124
rect 1163 120 1164 124
rect 1158 119 1164 120
rect 1198 123 1204 124
rect 1198 119 1199 123
rect 1203 119 1204 123
rect 1326 120 1327 124
rect 1331 120 1332 124
rect 1326 119 1332 120
rect 1470 124 1476 125
rect 1488 124 1490 154
rect 1566 153 1572 154
rect 1566 149 1567 153
rect 1571 149 1572 153
rect 1566 148 1572 149
rect 1566 135 1572 136
rect 1566 131 1567 135
rect 1571 131 1572 135
rect 1566 130 1572 131
rect 1470 120 1471 124
rect 1475 120 1476 124
rect 1470 119 1476 120
rect 1486 123 1492 124
rect 1486 119 1487 123
rect 1491 119 1492 123
rect 1568 119 1570 130
rect 111 118 115 119
rect 111 113 115 114
rect 511 118 515 119
rect 594 118 600 119
rect 615 118 619 119
rect 718 118 724 119
rect 727 118 731 119
rect 822 118 828 119
rect 855 118 859 119
rect 958 118 964 119
rect 999 118 1003 119
rect 1110 118 1116 119
rect 1159 118 1163 119
rect 1198 118 1204 119
rect 1327 118 1331 119
rect 511 113 515 114
rect 615 113 619 114
rect 727 113 731 114
rect 855 113 859 114
rect 999 113 1003 114
rect 1159 113 1163 114
rect 1327 113 1331 114
rect 1471 118 1475 119
rect 1486 118 1492 119
rect 1567 118 1571 119
rect 1471 113 1475 114
rect 1567 113 1571 114
<< m4c >>
rect 111 1650 115 1654
rect 135 1650 139 1654
rect 223 1650 227 1654
rect 311 1650 315 1654
rect 1567 1650 1571 1654
rect 111 1586 115 1590
rect 135 1586 139 1590
rect 183 1586 187 1590
rect 223 1586 227 1590
rect 271 1586 275 1590
rect 311 1586 315 1590
rect 359 1586 363 1590
rect 1567 1586 1571 1590
rect 111 1514 115 1518
rect 183 1514 187 1518
rect 271 1514 275 1518
rect 351 1514 355 1518
rect 359 1514 363 1518
rect 439 1514 443 1518
rect 527 1514 531 1518
rect 615 1514 619 1518
rect 1567 1514 1571 1518
rect 111 1430 115 1434
rect 351 1430 355 1434
rect 439 1430 443 1434
rect 527 1430 531 1434
rect 615 1430 619 1434
rect 663 1430 667 1434
rect 751 1430 755 1434
rect 839 1430 843 1434
rect 927 1430 931 1434
rect 1567 1430 1571 1434
rect 111 1354 115 1358
rect 663 1354 667 1358
rect 751 1354 755 1358
rect 815 1354 819 1358
rect 839 1354 843 1358
rect 927 1354 931 1358
rect 935 1354 939 1358
rect 1055 1354 1059 1358
rect 1175 1354 1179 1358
rect 1295 1354 1299 1358
rect 1415 1354 1419 1358
rect 1567 1354 1571 1358
rect 111 1290 115 1294
rect 543 1290 547 1294
rect 695 1290 699 1294
rect 815 1290 819 1294
rect 863 1290 867 1294
rect 935 1290 939 1294
rect 1039 1290 1043 1294
rect 1055 1290 1059 1294
rect 111 1206 115 1210
rect 199 1206 203 1210
rect 415 1206 419 1210
rect 543 1206 547 1210
rect 647 1206 651 1210
rect 695 1206 699 1210
rect 863 1206 867 1210
rect 895 1206 899 1210
rect 1175 1290 1179 1294
rect 1215 1290 1219 1294
rect 1295 1290 1299 1294
rect 1399 1290 1403 1294
rect 1415 1290 1419 1294
rect 1039 1206 1043 1210
rect 1151 1206 1155 1210
rect 1215 1206 1219 1210
rect 111 1134 115 1138
rect 135 1134 139 1138
rect 199 1134 203 1138
rect 415 1134 419 1138
rect 559 1134 563 1138
rect 647 1134 651 1138
rect 895 1134 899 1138
rect 991 1134 995 1138
rect 1151 1134 1155 1138
rect 111 1066 115 1070
rect 135 1066 139 1070
rect 239 1066 243 1070
rect 559 1066 563 1070
rect 631 1066 635 1070
rect 991 1066 995 1070
rect 1031 1066 1035 1070
rect 111 1002 115 1006
rect 239 1002 243 1006
rect 415 1002 419 1006
rect 631 1002 635 1006
rect 663 1002 667 1006
rect 111 922 115 926
rect 415 922 419 926
rect 543 922 547 926
rect 919 1002 923 1006
rect 1031 1002 1035 1006
rect 1175 1002 1179 1006
rect 1399 1206 1403 1210
rect 1415 1206 1419 1210
rect 1567 1290 1571 1294
rect 1567 1206 1571 1210
rect 1415 1134 1419 1138
rect 1423 1134 1427 1138
rect 1567 1134 1571 1138
rect 1423 1066 1427 1070
rect 1431 1066 1435 1070
rect 1567 1066 1571 1070
rect 1431 1002 1435 1006
rect 1439 1002 1443 1006
rect 1567 1002 1571 1006
rect 663 922 667 926
rect 751 922 755 926
rect 919 922 923 926
rect 975 922 979 926
rect 1175 922 1179 926
rect 1207 922 1211 926
rect 111 850 115 854
rect 543 850 547 854
rect 751 850 755 854
rect 775 850 779 854
rect 927 850 931 854
rect 975 850 979 854
rect 1087 850 1091 854
rect 1207 850 1211 854
rect 111 770 115 774
rect 775 770 779 774
rect 855 770 859 774
rect 1255 850 1259 854
rect 1439 922 1443 926
rect 1567 922 1571 926
rect 1423 850 1427 854
rect 1439 850 1443 854
rect 927 770 931 774
rect 975 770 979 774
rect 1087 770 1091 774
rect 1103 770 1107 774
rect 1239 770 1243 774
rect 1255 770 1259 774
rect 111 698 115 702
rect 735 698 739 702
rect 855 698 859 702
rect 935 698 939 702
rect 975 698 979 702
rect 1103 698 1107 702
rect 1135 698 1139 702
rect 111 634 115 638
rect 607 634 611 638
rect 735 634 739 638
rect 847 634 851 638
rect 1239 698 1243 702
rect 935 634 939 638
rect 1087 634 1091 638
rect 1135 634 1139 638
rect 111 562 115 566
rect 359 562 363 566
rect 591 562 595 566
rect 607 562 611 566
rect 831 562 835 566
rect 847 562 851 566
rect 1079 562 1083 566
rect 1087 562 1091 566
rect 1375 770 1379 774
rect 1423 770 1427 774
rect 1567 850 1571 854
rect 1567 770 1571 774
rect 1343 698 1347 702
rect 1375 698 1379 702
rect 1327 634 1331 638
rect 1343 634 1347 638
rect 1567 698 1571 702
rect 1567 634 1571 638
rect 1327 562 1331 566
rect 111 482 115 486
rect 151 482 155 486
rect 359 482 363 486
rect 439 482 443 486
rect 591 482 595 486
rect 735 482 739 486
rect 831 482 835 486
rect 1567 562 1571 566
rect 1039 482 1043 486
rect 1079 482 1083 486
rect 111 406 115 410
rect 151 406 155 410
rect 175 406 179 410
rect 439 406 443 410
rect 567 406 571 410
rect 735 406 739 410
rect 967 406 971 410
rect 1039 406 1043 410
rect 1327 482 1331 486
rect 1343 482 1347 486
rect 1567 482 1571 486
rect 1343 406 1347 410
rect 1367 406 1371 410
rect 111 338 115 342
rect 175 338 179 342
rect 231 338 235 342
rect 511 338 515 342
rect 567 338 571 342
rect 799 338 803 342
rect 1567 406 1571 410
rect 967 338 971 342
rect 1095 338 1099 342
rect 1367 338 1371 342
rect 1399 338 1403 342
rect 1567 338 1571 342
rect 111 258 115 262
rect 231 258 235 262
rect 423 258 427 262
rect 511 258 515 262
rect 663 258 667 262
rect 799 258 803 262
rect 911 258 915 262
rect 1095 258 1099 262
rect 1167 258 1171 262
rect 1399 258 1403 262
rect 1431 258 1435 262
rect 111 178 115 182
rect 423 178 427 182
rect 511 178 515 182
rect 1567 258 1571 262
rect 615 178 619 182
rect 663 178 667 182
rect 727 178 731 182
rect 855 178 859 182
rect 911 178 915 182
rect 999 178 1003 182
rect 1159 178 1163 182
rect 1167 178 1171 182
rect 1327 178 1331 182
rect 1431 178 1435 182
rect 1471 178 1475 182
rect 1567 178 1571 182
rect 111 114 115 118
rect 511 114 515 118
rect 615 114 619 118
rect 727 114 731 118
rect 855 114 859 118
rect 999 114 1003 118
rect 1159 114 1163 118
rect 1327 114 1331 118
rect 1471 114 1475 118
rect 1567 114 1571 118
<< m4 >>
rect 96 1649 97 1655
rect 103 1654 1603 1655
rect 103 1650 111 1654
rect 115 1650 135 1654
rect 139 1650 223 1654
rect 227 1650 311 1654
rect 315 1650 1567 1654
rect 1571 1650 1603 1654
rect 103 1649 1603 1650
rect 1609 1649 1610 1655
rect 84 1585 85 1591
rect 91 1590 1591 1591
rect 91 1586 111 1590
rect 115 1586 135 1590
rect 139 1586 183 1590
rect 187 1586 223 1590
rect 227 1586 271 1590
rect 275 1586 311 1590
rect 315 1586 359 1590
rect 363 1586 1567 1590
rect 1571 1586 1591 1590
rect 91 1585 1591 1586
rect 1597 1585 1598 1591
rect 96 1513 97 1519
rect 103 1518 1603 1519
rect 103 1514 111 1518
rect 115 1514 183 1518
rect 187 1514 271 1518
rect 275 1514 351 1518
rect 355 1514 359 1518
rect 363 1514 439 1518
rect 443 1514 527 1518
rect 531 1514 615 1518
rect 619 1514 1567 1518
rect 1571 1514 1603 1518
rect 103 1513 1603 1514
rect 1609 1513 1610 1519
rect 84 1429 85 1435
rect 91 1434 1591 1435
rect 91 1430 111 1434
rect 115 1430 351 1434
rect 355 1430 439 1434
rect 443 1430 527 1434
rect 531 1430 615 1434
rect 619 1430 663 1434
rect 667 1430 751 1434
rect 755 1430 839 1434
rect 843 1430 927 1434
rect 931 1430 1567 1434
rect 1571 1430 1591 1434
rect 91 1429 1591 1430
rect 1597 1429 1598 1435
rect 96 1353 97 1359
rect 103 1358 1603 1359
rect 103 1354 111 1358
rect 115 1354 663 1358
rect 667 1354 751 1358
rect 755 1354 815 1358
rect 819 1354 839 1358
rect 843 1354 927 1358
rect 931 1354 935 1358
rect 939 1354 1055 1358
rect 1059 1354 1175 1358
rect 1179 1354 1295 1358
rect 1299 1354 1415 1358
rect 1419 1354 1567 1358
rect 1571 1354 1603 1358
rect 103 1353 1603 1354
rect 1609 1353 1610 1359
rect 84 1289 85 1295
rect 91 1294 1591 1295
rect 91 1290 111 1294
rect 115 1290 543 1294
rect 547 1290 695 1294
rect 699 1290 815 1294
rect 819 1290 863 1294
rect 867 1290 935 1294
rect 939 1290 1039 1294
rect 1043 1290 1055 1294
rect 1059 1290 1175 1294
rect 1179 1290 1215 1294
rect 1219 1290 1295 1294
rect 1299 1290 1399 1294
rect 1403 1290 1415 1294
rect 1419 1290 1567 1294
rect 1571 1290 1591 1294
rect 91 1289 1591 1290
rect 1597 1289 1598 1295
rect 96 1205 97 1211
rect 103 1210 1603 1211
rect 103 1206 111 1210
rect 115 1206 199 1210
rect 203 1206 415 1210
rect 419 1206 543 1210
rect 547 1206 647 1210
rect 651 1206 695 1210
rect 699 1206 863 1210
rect 867 1206 895 1210
rect 899 1206 1039 1210
rect 1043 1206 1151 1210
rect 1155 1206 1215 1210
rect 1219 1206 1399 1210
rect 1403 1206 1415 1210
rect 1419 1206 1567 1210
rect 1571 1206 1603 1210
rect 103 1205 1603 1206
rect 1609 1205 1610 1211
rect 84 1133 85 1139
rect 91 1138 1591 1139
rect 91 1134 111 1138
rect 115 1134 135 1138
rect 139 1134 199 1138
rect 203 1134 415 1138
rect 419 1134 559 1138
rect 563 1134 647 1138
rect 651 1134 895 1138
rect 899 1134 991 1138
rect 995 1134 1151 1138
rect 1155 1134 1415 1138
rect 1419 1134 1423 1138
rect 1427 1134 1567 1138
rect 1571 1134 1591 1138
rect 91 1133 1591 1134
rect 1597 1133 1598 1139
rect 96 1065 97 1071
rect 103 1070 1603 1071
rect 103 1066 111 1070
rect 115 1066 135 1070
rect 139 1066 239 1070
rect 243 1066 559 1070
rect 563 1066 631 1070
rect 635 1066 991 1070
rect 995 1066 1031 1070
rect 1035 1066 1423 1070
rect 1427 1066 1431 1070
rect 1435 1066 1567 1070
rect 1571 1066 1603 1070
rect 103 1065 1603 1066
rect 1609 1065 1610 1071
rect 84 1001 85 1007
rect 91 1006 1591 1007
rect 91 1002 111 1006
rect 115 1002 239 1006
rect 243 1002 415 1006
rect 419 1002 631 1006
rect 635 1002 663 1006
rect 667 1002 919 1006
rect 923 1002 1031 1006
rect 1035 1002 1175 1006
rect 1179 1002 1431 1006
rect 1435 1002 1439 1006
rect 1443 1002 1567 1006
rect 1571 1002 1591 1006
rect 91 1001 1591 1002
rect 1597 1001 1598 1007
rect 96 921 97 927
rect 103 926 1603 927
rect 103 922 111 926
rect 115 922 415 926
rect 419 922 543 926
rect 547 922 663 926
rect 667 922 751 926
rect 755 922 919 926
rect 923 922 975 926
rect 979 922 1175 926
rect 1179 922 1207 926
rect 1211 922 1439 926
rect 1443 922 1567 926
rect 1571 922 1603 926
rect 103 921 1603 922
rect 1609 921 1610 927
rect 84 849 85 855
rect 91 854 1591 855
rect 91 850 111 854
rect 115 850 543 854
rect 547 850 751 854
rect 755 850 775 854
rect 779 850 927 854
rect 931 850 975 854
rect 979 850 1087 854
rect 1091 850 1207 854
rect 1211 850 1255 854
rect 1259 850 1423 854
rect 1427 850 1439 854
rect 1443 850 1567 854
rect 1571 850 1591 854
rect 91 849 1591 850
rect 1597 849 1598 855
rect 96 769 97 775
rect 103 774 1603 775
rect 103 770 111 774
rect 115 770 775 774
rect 779 770 855 774
rect 859 770 927 774
rect 931 770 975 774
rect 979 770 1087 774
rect 1091 770 1103 774
rect 1107 770 1239 774
rect 1243 770 1255 774
rect 1259 770 1375 774
rect 1379 770 1423 774
rect 1427 770 1567 774
rect 1571 770 1603 774
rect 103 769 1603 770
rect 1609 769 1610 775
rect 84 697 85 703
rect 91 702 1591 703
rect 91 698 111 702
rect 115 698 735 702
rect 739 698 855 702
rect 859 698 935 702
rect 939 698 975 702
rect 979 698 1103 702
rect 1107 698 1135 702
rect 1139 698 1239 702
rect 1243 698 1343 702
rect 1347 698 1375 702
rect 1379 698 1567 702
rect 1571 698 1591 702
rect 91 697 1591 698
rect 1597 697 1598 703
rect 96 633 97 639
rect 103 638 1603 639
rect 103 634 111 638
rect 115 634 607 638
rect 611 634 735 638
rect 739 634 847 638
rect 851 634 935 638
rect 939 634 1087 638
rect 1091 634 1135 638
rect 1139 634 1327 638
rect 1331 634 1343 638
rect 1347 634 1567 638
rect 1571 634 1603 638
rect 103 633 1603 634
rect 1609 633 1610 639
rect 84 561 85 567
rect 91 566 1591 567
rect 91 562 111 566
rect 115 562 359 566
rect 363 562 591 566
rect 595 562 607 566
rect 611 562 831 566
rect 835 562 847 566
rect 851 562 1079 566
rect 1083 562 1087 566
rect 1091 562 1327 566
rect 1331 562 1567 566
rect 1571 562 1591 566
rect 91 561 1591 562
rect 1597 561 1598 567
rect 96 481 97 487
rect 103 486 1603 487
rect 103 482 111 486
rect 115 482 151 486
rect 155 482 359 486
rect 363 482 439 486
rect 443 482 591 486
rect 595 482 735 486
rect 739 482 831 486
rect 835 482 1039 486
rect 1043 482 1079 486
rect 1083 482 1327 486
rect 1331 482 1343 486
rect 1347 482 1567 486
rect 1571 482 1603 486
rect 103 481 1603 482
rect 1609 481 1610 487
rect 84 405 85 411
rect 91 410 1591 411
rect 91 406 111 410
rect 115 406 151 410
rect 155 406 175 410
rect 179 406 439 410
rect 443 406 567 410
rect 571 406 735 410
rect 739 406 967 410
rect 971 406 1039 410
rect 1043 406 1343 410
rect 1347 406 1367 410
rect 1371 406 1567 410
rect 1571 406 1591 410
rect 91 405 1591 406
rect 1597 405 1598 411
rect 96 337 97 343
rect 103 342 1603 343
rect 103 338 111 342
rect 115 338 175 342
rect 179 338 231 342
rect 235 338 511 342
rect 515 338 567 342
rect 571 338 799 342
rect 803 338 967 342
rect 971 338 1095 342
rect 1099 338 1367 342
rect 1371 338 1399 342
rect 1403 338 1567 342
rect 1571 338 1603 342
rect 103 337 1603 338
rect 1609 337 1610 343
rect 84 257 85 263
rect 91 262 1591 263
rect 91 258 111 262
rect 115 258 231 262
rect 235 258 423 262
rect 427 258 511 262
rect 515 258 663 262
rect 667 258 799 262
rect 803 258 911 262
rect 915 258 1095 262
rect 1099 258 1167 262
rect 1171 258 1399 262
rect 1403 258 1431 262
rect 1435 258 1567 262
rect 1571 258 1591 262
rect 91 257 1591 258
rect 1597 257 1598 263
rect 96 177 97 183
rect 103 182 1603 183
rect 103 178 111 182
rect 115 178 423 182
rect 427 178 511 182
rect 515 178 615 182
rect 619 178 663 182
rect 667 178 727 182
rect 731 178 855 182
rect 859 178 911 182
rect 915 178 999 182
rect 1003 178 1159 182
rect 1163 178 1167 182
rect 1171 178 1327 182
rect 1331 178 1431 182
rect 1435 178 1471 182
rect 1475 178 1567 182
rect 1571 178 1603 182
rect 103 177 1603 178
rect 1609 177 1610 183
rect 84 113 85 119
rect 91 118 1591 119
rect 91 114 111 118
rect 115 114 511 118
rect 515 114 615 118
rect 619 114 727 118
rect 731 114 855 118
rect 859 114 999 118
rect 1003 114 1159 118
rect 1163 114 1327 118
rect 1331 114 1471 118
rect 1475 114 1567 118
rect 1571 114 1591 118
rect 91 113 1591 114
rect 1597 113 1598 119
<< m5c >>
rect 97 1649 103 1655
rect 1603 1649 1609 1655
rect 85 1585 91 1591
rect 1591 1585 1597 1591
rect 97 1513 103 1519
rect 1603 1513 1609 1519
rect 85 1429 91 1435
rect 1591 1429 1597 1435
rect 97 1353 103 1359
rect 1603 1353 1609 1359
rect 85 1289 91 1295
rect 1591 1289 1597 1295
rect 97 1205 103 1211
rect 1603 1205 1609 1211
rect 85 1133 91 1139
rect 1591 1133 1597 1139
rect 97 1065 103 1071
rect 1603 1065 1609 1071
rect 85 1001 91 1007
rect 1591 1001 1597 1007
rect 97 921 103 927
rect 1603 921 1609 927
rect 85 849 91 855
rect 1591 849 1597 855
rect 97 769 103 775
rect 1603 769 1609 775
rect 85 697 91 703
rect 1591 697 1597 703
rect 97 633 103 639
rect 1603 633 1609 639
rect 85 561 91 567
rect 1591 561 1597 567
rect 97 481 103 487
rect 1603 481 1609 487
rect 85 405 91 411
rect 1591 405 1597 411
rect 97 337 103 343
rect 1603 337 1609 343
rect 85 257 91 263
rect 1591 257 1597 263
rect 97 177 103 183
rect 1603 177 1609 183
rect 85 113 91 119
rect 1591 113 1597 119
<< m5 >>
rect 84 1591 92 1656
rect 84 1585 85 1591
rect 91 1585 92 1591
rect 84 1435 92 1585
rect 84 1429 85 1435
rect 91 1429 92 1435
rect 84 1295 92 1429
rect 84 1289 85 1295
rect 91 1289 92 1295
rect 84 1139 92 1289
rect 84 1133 85 1139
rect 91 1133 92 1139
rect 84 1007 92 1133
rect 84 1001 85 1007
rect 91 1001 92 1007
rect 84 855 92 1001
rect 84 849 85 855
rect 91 849 92 855
rect 84 703 92 849
rect 84 697 85 703
rect 91 697 92 703
rect 84 567 92 697
rect 84 561 85 567
rect 91 561 92 567
rect 84 411 92 561
rect 84 405 85 411
rect 91 405 92 411
rect 84 263 92 405
rect 84 257 85 263
rect 91 257 92 263
rect 84 119 92 257
rect 84 113 85 119
rect 91 113 92 119
rect 84 72 92 113
rect 96 1655 104 1656
rect 96 1649 97 1655
rect 103 1649 104 1655
rect 96 1519 104 1649
rect 96 1513 97 1519
rect 103 1513 104 1519
rect 96 1359 104 1513
rect 96 1353 97 1359
rect 103 1353 104 1359
rect 96 1211 104 1353
rect 96 1205 97 1211
rect 103 1205 104 1211
rect 96 1071 104 1205
rect 96 1065 97 1071
rect 103 1065 104 1071
rect 96 927 104 1065
rect 96 921 97 927
rect 103 921 104 927
rect 96 775 104 921
rect 96 769 97 775
rect 103 769 104 775
rect 96 639 104 769
rect 96 633 97 639
rect 103 633 104 639
rect 96 487 104 633
rect 96 481 97 487
rect 103 481 104 487
rect 96 343 104 481
rect 96 337 97 343
rect 103 337 104 343
rect 96 183 104 337
rect 96 177 97 183
rect 103 177 104 183
rect 96 72 104 177
rect 1590 1591 1598 1656
rect 1590 1585 1591 1591
rect 1597 1585 1598 1591
rect 1590 1435 1598 1585
rect 1590 1429 1591 1435
rect 1597 1429 1598 1435
rect 1590 1295 1598 1429
rect 1590 1289 1591 1295
rect 1597 1289 1598 1295
rect 1590 1139 1598 1289
rect 1590 1133 1591 1139
rect 1597 1133 1598 1139
rect 1590 1007 1598 1133
rect 1590 1001 1591 1007
rect 1597 1001 1598 1007
rect 1590 855 1598 1001
rect 1590 849 1591 855
rect 1597 849 1598 855
rect 1590 703 1598 849
rect 1590 697 1591 703
rect 1597 697 1598 703
rect 1590 567 1598 697
rect 1590 561 1591 567
rect 1597 561 1598 567
rect 1590 411 1598 561
rect 1590 405 1591 411
rect 1597 405 1598 411
rect 1590 263 1598 405
rect 1590 257 1591 263
rect 1597 257 1598 263
rect 1590 119 1598 257
rect 1590 113 1591 119
rect 1597 113 1598 119
rect 1590 72 1598 113
rect 1602 1655 1610 1656
rect 1602 1649 1603 1655
rect 1609 1649 1610 1655
rect 1602 1519 1610 1649
rect 1602 1513 1603 1519
rect 1609 1513 1610 1519
rect 1602 1359 1610 1513
rect 1602 1353 1603 1359
rect 1609 1353 1610 1359
rect 1602 1211 1610 1353
rect 1602 1205 1603 1211
rect 1609 1205 1610 1211
rect 1602 1071 1610 1205
rect 1602 1065 1603 1071
rect 1609 1065 1610 1071
rect 1602 927 1610 1065
rect 1602 921 1603 927
rect 1609 921 1610 927
rect 1602 775 1610 921
rect 1602 769 1603 775
rect 1609 769 1610 775
rect 1602 639 1610 769
rect 1602 633 1603 639
rect 1609 633 1610 639
rect 1602 487 1610 633
rect 1602 481 1603 487
rect 1609 481 1610 487
rect 1602 343 1610 481
rect 1602 337 1603 343
rect 1609 337 1610 343
rect 1602 183 1610 337
rect 1602 177 1603 183
rect 1609 177 1610 183
rect 1602 72 1610 177
use welltap_svt  __well_tap__0
timestamp 1730767243
transform 1 0 104 0 1 128
box 8 4 12 24
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__0
timestamp 1730767243
transform 1 0 104 0 1 128
box 8 4 12 24
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use _0_0cell_0_0gcelem3x0  celem_562_6_acx0
timestamp 1730767243
transform 1 0 504 0 1 116
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_562_6_acx0
timestamp 1730767243
transform 1 0 504 0 1 116
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_563_6_acx0
timestamp 1730767243
transform 1 0 608 0 1 116
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_563_6_acx0
timestamp 1730767243
transform 1 0 608 0 1 116
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_564_6_acx0
timestamp 1730767243
transform 1 0 720 0 1 116
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_564_6_acx0
timestamp 1730767243
transform 1 0 720 0 1 116
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_565_6_acx0
timestamp 1730767243
transform 1 0 848 0 1 116
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_565_6_acx0
timestamp 1730767243
transform 1 0 848 0 1 116
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_566_6_acx0
timestamp 1730767243
transform 1 0 992 0 1 116
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_566_6_acx0
timestamp 1730767243
transform 1 0 992 0 1 116
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_567_6_acx0
timestamp 1730767243
transform 1 0 1152 0 1 116
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_567_6_acx0
timestamp 1730767243
transform 1 0 1152 0 1 116
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_599_6_acx0
timestamp 1730767243
transform 1 0 1320 0 1 116
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_599_6_acx0
timestamp 1730767243
transform 1 0 1320 0 1 116
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_598_6_acx0
timestamp 1730767243
transform 1 0 1464 0 1 116
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_598_6_acx0
timestamp 1730767243
transform 1 0 1464 0 1 116
box 8 4 79 60
use welltap_svt  __well_tap__1
timestamp 1730767243
transform 1 0 1560 0 1 128
box 8 4 12 24
use welltap_svt  __well_tap__1
timestamp 1730767243
transform 1 0 1560 0 1 128
box 8 4 12 24
use welltap_svt  __well_tap__2
timestamp 1730767243
transform 1 0 104 0 -1 248
box 8 4 12 24
use welltap_svt  __well_tap__2
timestamp 1730767243
transform 1 0 104 0 -1 248
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_560_6_acx0
timestamp 1730767243
transform 1 0 416 0 -1 260
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_560_6_acx0
timestamp 1730767243
transform 1 0 416 0 -1 260
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_561_6_acx0
timestamp 1730767243
transform 1 0 656 0 -1 260
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_561_6_acx0
timestamp 1730767243
transform 1 0 656 0 -1 260
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_569_6_acx0
timestamp 1730767243
transform 1 0 904 0 -1 260
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_569_6_acx0
timestamp 1730767243
transform 1 0 904 0 -1 260
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_568_6_acx0
timestamp 1730767243
transform 1 0 1160 0 -1 260
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_568_6_acx0
timestamp 1730767243
transform 1 0 1160 0 -1 260
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_597_6_acx0
timestamp 1730767243
transform 1 0 1424 0 -1 260
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_597_6_acx0
timestamp 1730767243
transform 1 0 1424 0 -1 260
box 8 4 79 60
use welltap_svt  __well_tap__3
timestamp 1730767243
transform 1 0 1560 0 -1 248
box 8 4 12 24
use welltap_svt  __well_tap__3
timestamp 1730767243
transform 1 0 1560 0 -1 248
box 8 4 12 24
use welltap_svt  __well_tap__4
timestamp 1730767243
transform 1 0 104 0 1 288
box 8 4 12 24
use welltap_svt  __well_tap__4
timestamp 1730767243
transform 1 0 104 0 1 288
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_559_6_acx0
timestamp 1730767243
transform 1 0 224 0 1 276
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_559_6_acx0
timestamp 1730767243
transform 1 0 224 0 1 276
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_558_6_acx0
timestamp 1730767243
transform 1 0 504 0 1 276
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_558_6_acx0
timestamp 1730767243
transform 1 0 504 0 1 276
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_557_6_acx0
timestamp 1730767243
transform 1 0 792 0 1 276
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_557_6_acx0
timestamp 1730767243
transform 1 0 792 0 1 276
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_570_6_acx0
timestamp 1730767243
transform 1 0 1088 0 1 276
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_570_6_acx0
timestamp 1730767243
transform 1 0 1088 0 1 276
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_596_6_acx0
timestamp 1730767243
transform 1 0 1392 0 1 276
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_596_6_acx0
timestamp 1730767243
transform 1 0 1392 0 1 276
box 8 4 79 60
use welltap_svt  __well_tap__5
timestamp 1730767243
transform 1 0 1560 0 1 288
box 8 4 12 24
use welltap_svt  __well_tap__5
timestamp 1730767243
transform 1 0 1560 0 1 288
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_554_6_acx0
timestamp 1730767243
transform 1 0 144 0 1 420
box 8 4 79 60
use welltap_svt  __well_tap__6
timestamp 1730767243
transform 1 0 104 0 -1 396
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_554_6_acx0
timestamp 1730767243
transform 1 0 144 0 1 420
box 8 4 79 60
use welltap_svt  __well_tap__6
timestamp 1730767243
transform 1 0 104 0 -1 396
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_555_6_acx0
timestamp 1730767243
transform 1 0 168 0 -1 408
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_555_6_acx0
timestamp 1730767243
transform 1 0 168 0 -1 408
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_553_6_acx0
timestamp 1730767243
transform 1 0 432 0 1 420
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_553_6_acx0
timestamp 1730767243
transform 1 0 432 0 1 420
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_556_6_acx0
timestamp 1730767243
transform 1 0 560 0 -1 408
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_556_6_acx0
timestamp 1730767243
transform 1 0 560 0 -1 408
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_552_6_acx0
timestamp 1730767243
transform 1 0 728 0 1 420
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_552_6_acx0
timestamp 1730767243
transform 1 0 728 0 1 420
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_571_6_acx0
timestamp 1730767243
transform 1 0 960 0 -1 408
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_571_6_acx0
timestamp 1730767243
transform 1 0 960 0 -1 408
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_572_6_acx0
timestamp 1730767243
transform 1 0 1032 0 1 420
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_572_6_acx0
timestamp 1730767243
transform 1 0 1032 0 1 420
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_594_6_acx0
timestamp 1730767243
transform 1 0 1336 0 1 420
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_595_6_acx0
timestamp 1730767243
transform 1 0 1360 0 -1 408
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_594_6_acx0
timestamp 1730767243
transform 1 0 1336 0 1 420
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_595_6_acx0
timestamp 1730767243
transform 1 0 1360 0 -1 408
box 8 4 79 60
use welltap_svt  __well_tap__7
timestamp 1730767243
transform 1 0 1560 0 -1 396
box 8 4 12 24
use welltap_svt  __well_tap__7
timestamp 1730767243
transform 1 0 1560 0 -1 396
box 8 4 12 24
use welltap_svt  __well_tap__8
timestamp 1730767243
transform 1 0 104 0 1 432
box 8 4 12 24
use welltap_svt  __well_tap__8
timestamp 1730767243
transform 1 0 104 0 1 432
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_549_6_acx0
timestamp 1730767243
transform 1 0 352 0 -1 564
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_549_6_acx0
timestamp 1730767243
transform 1 0 352 0 -1 564
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_550_6_acx0
timestamp 1730767243
transform 1 0 584 0 -1 564
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_550_6_acx0
timestamp 1730767243
transform 1 0 584 0 -1 564
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_551_6_acx0
timestamp 1730767243
transform 1 0 824 0 -1 564
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_551_6_acx0
timestamp 1730767243
transform 1 0 824 0 -1 564
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_573_6_acx0
timestamp 1730767243
transform 1 0 1072 0 -1 564
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_573_6_acx0
timestamp 1730767243
transform 1 0 1072 0 -1 564
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_593_6_acx0
timestamp 1730767243
transform 1 0 1320 0 -1 564
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_593_6_acx0
timestamp 1730767243
transform 1 0 1320 0 -1 564
box 8 4 79 60
use welltap_svt  __well_tap__9
timestamp 1730767243
transform 1 0 1560 0 1 432
box 8 4 12 24
use welltap_svt  __well_tap__9
timestamp 1730767243
transform 1 0 1560 0 1 432
box 8 4 12 24
use welltap_svt  __well_tap__10
timestamp 1730767243
transform 1 0 104 0 -1 552
box 8 4 12 24
use welltap_svt  __well_tap__12
timestamp 1730767243
transform 1 0 104 0 1 584
box 8 4 12 24
use welltap_svt  __well_tap__10
timestamp 1730767243
transform 1 0 104 0 -1 552
box 8 4 12 24
use welltap_svt  __well_tap__12
timestamp 1730767243
transform 1 0 104 0 1 584
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_548_6_acx0
timestamp 1730767243
transform 1 0 600 0 1 572
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_548_6_acx0
timestamp 1730767243
transform 1 0 600 0 1 572
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_547_6_acx0
timestamp 1730767243
transform 1 0 840 0 1 572
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_547_6_acx0
timestamp 1730767243
transform 1 0 840 0 1 572
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_574_6_acx0
timestamp 1730767243
transform 1 0 1080 0 1 572
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_574_6_acx0
timestamp 1730767243
transform 1 0 1080 0 1 572
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_592_6_acx0
timestamp 1730767243
transform 1 0 1320 0 1 572
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_592_6_acx0
timestamp 1730767243
transform 1 0 1320 0 1 572
box 8 4 79 60
use welltap_svt  __well_tap__11
timestamp 1730767243
transform 1 0 1560 0 -1 552
box 8 4 12 24
use welltap_svt  __well_tap__13
timestamp 1730767243
transform 1 0 1560 0 1 584
box 8 4 12 24
use welltap_svt  __well_tap__11
timestamp 1730767243
transform 1 0 1560 0 -1 552
box 8 4 12 24
use welltap_svt  __well_tap__13
timestamp 1730767243
transform 1 0 1560 0 1 584
box 8 4 12 24
use welltap_svt  __well_tap__14
timestamp 1730767243
transform 1 0 104 0 -1 688
box 8 4 12 24
use welltap_svt  __well_tap__14
timestamp 1730767243
transform 1 0 104 0 -1 688
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_546_6_acx0
timestamp 1730767243
transform 1 0 728 0 -1 700
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_546_6_acx0
timestamp 1730767243
transform 1 0 728 0 -1 700
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_545_6_acx0
timestamp 1730767243
transform 1 0 928 0 -1 700
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_545_6_acx0
timestamp 1730767243
transform 1 0 928 0 -1 700
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_544_6_acx0
timestamp 1730767243
transform 1 0 1128 0 -1 700
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_544_6_acx0
timestamp 1730767243
transform 1 0 1128 0 -1 700
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_591_6_acx0
timestamp 1730767243
transform 1 0 1336 0 -1 700
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_591_6_acx0
timestamp 1730767243
transform 1 0 1336 0 -1 700
box 8 4 79 60
use welltap_svt  __well_tap__15
timestamp 1730767243
transform 1 0 1560 0 -1 688
box 8 4 12 24
use welltap_svt  __well_tap__15
timestamp 1730767243
transform 1 0 1560 0 -1 688
box 8 4 12 24
use welltap_svt  __well_tap__16
timestamp 1730767243
transform 1 0 104 0 1 720
box 8 4 12 24
use welltap_svt  __well_tap__16
timestamp 1730767243
transform 1 0 104 0 1 720
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_541_6_acx0
timestamp 1730767243
transform 1 0 848 0 1 708
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_541_6_acx0
timestamp 1730767243
transform 1 0 848 0 1 708
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_542_6_acx0
timestamp 1730767243
transform 1 0 968 0 1 708
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_542_6_acx0
timestamp 1730767243
transform 1 0 968 0 1 708
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_543_6_acx0
timestamp 1730767243
transform 1 0 1096 0 1 708
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_543_6_acx0
timestamp 1730767243
transform 1 0 1096 0 1 708
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_575_6_acx0
timestamp 1730767243
transform 1 0 1232 0 1 708
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_575_6_acx0
timestamp 1730767243
transform 1 0 1232 0 1 708
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_590_6_acx0
timestamp 1730767243
transform 1 0 1368 0 1 708
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_590_6_acx0
timestamp 1730767243
transform 1 0 1368 0 1 708
box 8 4 79 60
use welltap_svt  __well_tap__17
timestamp 1730767243
transform 1 0 1560 0 1 720
box 8 4 12 24
use welltap_svt  __well_tap__17
timestamp 1730767243
transform 1 0 1560 0 1 720
box 8 4 12 24
use welltap_svt  __well_tap__18
timestamp 1730767243
transform 1 0 104 0 -1 840
box 8 4 12 24
use welltap_svt  __well_tap__20
timestamp 1730767243
transform 1 0 104 0 1 872
box 8 4 12 24
use welltap_svt  __well_tap__18
timestamp 1730767243
transform 1 0 104 0 -1 840
box 8 4 12 24
use welltap_svt  __well_tap__20
timestamp 1730767243
transform 1 0 104 0 1 872
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_534_6_acx0
timestamp 1730767243
transform 1 0 536 0 1 860
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_534_6_acx0
timestamp 1730767243
transform 1 0 536 0 1 860
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_535_6_acx0
timestamp 1730767243
transform 1 0 744 0 1 860
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_540_6_acx0
timestamp 1730767243
transform 1 0 768 0 -1 852
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_535_6_acx0
timestamp 1730767243
transform 1 0 744 0 1 860
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_540_6_acx0
timestamp 1730767243
transform 1 0 768 0 -1 852
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_536_6_acx0
timestamp 1730767243
transform 1 0 968 0 1 860
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_539_6_acx0
timestamp 1730767243
transform 1 0 920 0 -1 852
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_536_6_acx0
timestamp 1730767243
transform 1 0 968 0 1 860
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_539_6_acx0
timestamp 1730767243
transform 1 0 920 0 -1 852
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_538_6_acx0
timestamp 1730767243
transform 1 0 1080 0 -1 852
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_538_6_acx0
timestamp 1730767243
transform 1 0 1080 0 -1 852
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_537_6_acx0
timestamp 1730767243
transform 1 0 1200 0 1 860
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_537_6_acx0
timestamp 1730767243
transform 1 0 1200 0 1 860
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_576_6_acx0
timestamp 1730767243
transform 1 0 1248 0 -1 852
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_576_6_acx0
timestamp 1730767243
transform 1 0 1248 0 -1 852
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_589_6_acx0
timestamp 1730767243
transform 1 0 1416 0 -1 852
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_589_6_acx0
timestamp 1730767243
transform 1 0 1416 0 -1 852
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_588_6_acx0
timestamp 1730767243
transform 1 0 1432 0 1 860
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_588_6_acx0
timestamp 1730767243
transform 1 0 1432 0 1 860
box 8 4 79 60
use welltap_svt  __well_tap__19
timestamp 1730767243
transform 1 0 1560 0 -1 840
box 8 4 12 24
use welltap_svt  __well_tap__21
timestamp 1730767243
transform 1 0 1560 0 1 872
box 8 4 12 24
use welltap_svt  __well_tap__19
timestamp 1730767243
transform 1 0 1560 0 -1 840
box 8 4 12 24
use welltap_svt  __well_tap__21
timestamp 1730767243
transform 1 0 1560 0 1 872
box 8 4 12 24
use welltap_svt  __well_tap__22
timestamp 1730767243
transform 1 0 104 0 -1 992
box 8 4 12 24
use welltap_svt  __well_tap__22
timestamp 1730767243
transform 1 0 104 0 -1 992
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_533_6_acx0
timestamp 1730767243
transform 1 0 408 0 -1 1004
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_533_6_acx0
timestamp 1730767243
transform 1 0 408 0 -1 1004
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_531_6_acx0
timestamp 1730767243
transform 1 0 656 0 -1 1004
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_531_6_acx0
timestamp 1730767243
transform 1 0 656 0 -1 1004
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_532_6_acx0
timestamp 1730767243
transform 1 0 912 0 -1 1004
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_532_6_acx0
timestamp 1730767243
transform 1 0 912 0 -1 1004
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_577_6_acx0
timestamp 1730767243
transform 1 0 1168 0 -1 1004
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_577_6_acx0
timestamp 1730767243
transform 1 0 1168 0 -1 1004
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_587_6_acx0
timestamp 1730767243
transform 1 0 1432 0 -1 1004
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_587_6_acx0
timestamp 1730767243
transform 1 0 1432 0 -1 1004
box 8 4 79 60
use welltap_svt  __well_tap__23
timestamp 1730767243
transform 1 0 1560 0 -1 992
box 8 4 12 24
use welltap_svt  __well_tap__23
timestamp 1730767243
transform 1 0 1560 0 -1 992
box 8 4 12 24
use welltap_svt  __well_tap__24
timestamp 1730767243
transform 1 0 104 0 1 1016
box 8 4 12 24
use welltap_svt  __well_tap__24
timestamp 1730767243
transform 1 0 104 0 1 1016
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_529_6_acx0
timestamp 1730767243
transform 1 0 232 0 1 1004
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_529_6_acx0
timestamp 1730767243
transform 1 0 232 0 1 1004
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_530_6_acx0
timestamp 1730767243
transform 1 0 624 0 1 1004
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_530_6_acx0
timestamp 1730767243
transform 1 0 624 0 1 1004
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_528_6_acx0
timestamp 1730767243
transform 1 0 1024 0 1 1004
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_528_6_acx0
timestamp 1730767243
transform 1 0 1024 0 1 1004
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_586_6_acx0
timestamp 1730767243
transform 1 0 1424 0 1 1004
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_586_6_acx0
timestamp 1730767243
transform 1 0 1424 0 1 1004
box 8 4 79 60
use welltap_svt  __well_tap__25
timestamp 1730767243
transform 1 0 1560 0 1 1016
box 8 4 12 24
use welltap_svt  __well_tap__25
timestamp 1730767243
transform 1 0 1560 0 1 1016
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_525_6_acx0
timestamp 1730767243
transform 1 0 128 0 -1 1136
box 8 4 79 60
use welltap_svt  __well_tap__26
timestamp 1730767243
transform 1 0 104 0 -1 1124
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_525_6_acx0
timestamp 1730767243
transform 1 0 128 0 -1 1136
box 8 4 79 60
use welltap_svt  __well_tap__26
timestamp 1730767243
transform 1 0 104 0 -1 1124
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_524_6_acx0
timestamp 1730767243
transform 1 0 192 0 1 1144
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_524_6_acx0
timestamp 1730767243
transform 1 0 192 0 1 1144
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_523_6_acx0
timestamp 1730767243
transform 1 0 408 0 1 1144
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_523_6_acx0
timestamp 1730767243
transform 1 0 408 0 1 1144
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_526_6_acx0
timestamp 1730767243
transform 1 0 552 0 -1 1136
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_526_6_acx0
timestamp 1730767243
transform 1 0 552 0 -1 1136
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_522_6_acx0
timestamp 1730767243
transform 1 0 640 0 1 1144
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_522_6_acx0
timestamp 1730767243
transform 1 0 640 0 1 1144
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_521_6_acx0
timestamp 1730767243
transform 1 0 888 0 1 1144
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_521_6_acx0
timestamp 1730767243
transform 1 0 888 0 1 1144
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_527_6_acx0
timestamp 1730767243
transform 1 0 984 0 -1 1136
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_527_6_acx0
timestamp 1730767243
transform 1 0 984 0 -1 1136
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_578_6_acx0
timestamp 1730767243
transform 1 0 1144 0 1 1144
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_578_6_acx0
timestamp 1730767243
transform 1 0 1144 0 1 1144
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_584_6_acx0
timestamp 1730767243
transform 1 0 1408 0 1 1144
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_585_6_acx0
timestamp 1730767243
transform 1 0 1416 0 -1 1136
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_584_6_acx0
timestamp 1730767243
transform 1 0 1408 0 1 1144
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_585_6_acx0
timestamp 1730767243
transform 1 0 1416 0 -1 1136
box 8 4 79 60
use welltap_svt  __well_tap__27
timestamp 1730767243
transform 1 0 1560 0 -1 1124
box 8 4 12 24
use welltap_svt  __well_tap__27
timestamp 1730767243
transform 1 0 1560 0 -1 1124
box 8 4 12 24
use welltap_svt  __well_tap__28
timestamp 1730767243
transform 1 0 104 0 1 1156
box 8 4 12 24
use welltap_svt  __well_tap__28
timestamp 1730767243
transform 1 0 104 0 1 1156
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_518_6_acx0
timestamp 1730767243
transform 1 0 536 0 -1 1292
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_518_6_acx0
timestamp 1730767243
transform 1 0 536 0 -1 1292
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_519_6_acx0
timestamp 1730767243
transform 1 0 688 0 -1 1292
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_519_6_acx0
timestamp 1730767243
transform 1 0 688 0 -1 1292
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_520_6_acx0
timestamp 1730767243
transform 1 0 856 0 -1 1292
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_520_6_acx0
timestamp 1730767243
transform 1 0 856 0 -1 1292
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_517_6_acx0
timestamp 1730767243
transform 1 0 1032 0 -1 1292
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_517_6_acx0
timestamp 1730767243
transform 1 0 1032 0 -1 1292
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_579_6_acx0
timestamp 1730767243
transform 1 0 1208 0 -1 1292
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_579_6_acx0
timestamp 1730767243
transform 1 0 1208 0 -1 1292
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_583_6_acx0
timestamp 1730767243
transform 1 0 1392 0 -1 1292
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_583_6_acx0
timestamp 1730767243
transform 1 0 1392 0 -1 1292
box 8 4 79 60
use welltap_svt  __well_tap__29
timestamp 1730767243
transform 1 0 1560 0 1 1156
box 8 4 12 24
use welltap_svt  __well_tap__29
timestamp 1730767243
transform 1 0 1560 0 1 1156
box 8 4 12 24
use welltap_svt  __well_tap__30
timestamp 1730767243
transform 1 0 104 0 -1 1280
box 8 4 12 24
use welltap_svt  __well_tap__32
timestamp 1730767243
transform 1 0 104 0 1 1304
box 8 4 12 24
use welltap_svt  __well_tap__30
timestamp 1730767243
transform 1 0 104 0 -1 1280
box 8 4 12 24
use welltap_svt  __well_tap__32
timestamp 1730767243
transform 1 0 104 0 1 1304
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_514_6_acx0
timestamp 1730767243
transform 1 0 808 0 1 1292
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_514_6_acx0
timestamp 1730767243
transform 1 0 808 0 1 1292
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_515_6_acx0
timestamp 1730767243
transform 1 0 928 0 1 1292
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_515_6_acx0
timestamp 1730767243
transform 1 0 928 0 1 1292
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_516_6_acx0
timestamp 1730767243
transform 1 0 1048 0 1 1292
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_516_6_acx0
timestamp 1730767243
transform 1 0 1048 0 1 1292
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_580_6_acx0
timestamp 1730767243
transform 1 0 1168 0 1 1292
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_580_6_acx0
timestamp 1730767243
transform 1 0 1168 0 1 1292
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_581_6_acx0
timestamp 1730767243
transform 1 0 1288 0 1 1292
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_581_6_acx0
timestamp 1730767243
transform 1 0 1288 0 1 1292
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_582_6_acx0
timestamp 1730767243
transform 1 0 1408 0 1 1292
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_582_6_acx0
timestamp 1730767243
transform 1 0 1408 0 1 1292
box 8 4 79 60
use welltap_svt  __well_tap__31
timestamp 1730767243
transform 1 0 1560 0 -1 1280
box 8 4 12 24
use welltap_svt  __well_tap__33
timestamp 1730767243
transform 1 0 1560 0 1 1304
box 8 4 12 24
use welltap_svt  __well_tap__31
timestamp 1730767243
transform 1 0 1560 0 -1 1280
box 8 4 12 24
use welltap_svt  __well_tap__33
timestamp 1730767243
transform 1 0 1560 0 1 1304
box 8 4 12 24
use welltap_svt  __well_tap__34
timestamp 1730767243
transform 1 0 104 0 -1 1420
box 8 4 12 24
use welltap_svt  __well_tap__34
timestamp 1730767243
transform 1 0 104 0 -1 1420
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_510_6_acx0
timestamp 1730767243
transform 1 0 656 0 -1 1432
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_510_6_acx0
timestamp 1730767243
transform 1 0 656 0 -1 1432
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_511_6_acx0
timestamp 1730767243
transform 1 0 744 0 -1 1432
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_511_6_acx0
timestamp 1730767243
transform 1 0 744 0 -1 1432
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_512_6_acx0
timestamp 1730767243
transform 1 0 832 0 -1 1432
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_512_6_acx0
timestamp 1730767243
transform 1 0 832 0 -1 1432
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_513_6_acx0
timestamp 1730767243
transform 1 0 920 0 -1 1432
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_513_6_acx0
timestamp 1730767243
transform 1 0 920 0 -1 1432
box 8 4 79 60
use welltap_svt  __well_tap__35
timestamp 1730767243
transform 1 0 1560 0 -1 1420
box 8 4 12 24
use welltap_svt  __well_tap__35
timestamp 1730767243
transform 1 0 1560 0 -1 1420
box 8 4 12 24
use welltap_svt  __well_tap__36
timestamp 1730767243
transform 1 0 104 0 1 1464
box 8 4 12 24
use welltap_svt  __well_tap__36
timestamp 1730767243
transform 1 0 104 0 1 1464
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_56_6_acx0
timestamp 1730767243
transform 1 0 344 0 1 1452
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_56_6_acx0
timestamp 1730767243
transform 1 0 344 0 1 1452
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_57_6_acx0
timestamp 1730767243
transform 1 0 432 0 1 1452
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_58_6_acx0
timestamp 1730767243
transform 1 0 520 0 1 1452
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_57_6_acx0
timestamp 1730767243
transform 1 0 432 0 1 1452
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_58_6_acx0
timestamp 1730767243
transform 1 0 520 0 1 1452
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_59_6_acx0
timestamp 1730767243
transform 1 0 608 0 1 1452
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_59_6_acx0
timestamp 1730767243
transform 1 0 608 0 1 1452
box 8 4 79 60
use welltap_svt  __well_tap__37
timestamp 1730767243
transform 1 0 1560 0 1 1464
box 8 4 12 24
use welltap_svt  __well_tap__37
timestamp 1730767243
transform 1 0 1560 0 1 1464
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_50_6_acx0
timestamp 1730767243
transform 1 0 128 0 1 1588
box 8 4 79 60
use welltap_svt  __well_tap__38
timestamp 1730767243
transform 1 0 104 0 -1 1576
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_50_6_acx0
timestamp 1730767243
transform 1 0 128 0 1 1588
box 8 4 79 60
use welltap_svt  __well_tap__38
timestamp 1730767243
transform 1 0 104 0 -1 1576
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_51_6_acx0
timestamp 1730767243
transform 1 0 216 0 1 1588
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_53_6_acx0
timestamp 1730767243
transform 1 0 176 0 -1 1588
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_51_6_acx0
timestamp 1730767243
transform 1 0 216 0 1 1588
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_53_6_acx0
timestamp 1730767243
transform 1 0 176 0 -1 1588
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_52_6_acx0
timestamp 1730767243
transform 1 0 304 0 1 1588
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_54_6_acx0
timestamp 1730767243
transform 1 0 264 0 -1 1588
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_52_6_acx0
timestamp 1730767243
transform 1 0 304 0 1 1588
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_54_6_acx0
timestamp 1730767243
transform 1 0 264 0 -1 1588
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_55_6_acx0
timestamp 1730767243
transform 1 0 352 0 -1 1588
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_55_6_acx0
timestamp 1730767243
transform 1 0 352 0 -1 1588
box 8 4 79 60
use welltap_svt  __well_tap__39
timestamp 1730767243
transform 1 0 1560 0 -1 1576
box 8 4 12 24
use welltap_svt  __well_tap__39
timestamp 1730767243
transform 1 0 1560 0 -1 1576
box 8 4 12 24
use welltap_svt  __well_tap__40
timestamp 1730767243
transform 1 0 104 0 1 1600
box 8 4 12 24
use welltap_svt  __well_tap__40
timestamp 1730767243
transform 1 0 104 0 1 1600
box 8 4 12 24
use welltap_svt  __well_tap__41
timestamp 1730767243
transform 1 0 1560 0 1 1600
box 8 4 12 24
use welltap_svt  __well_tap__41
timestamp 1730767243
transform 1 0 1560 0 1 1600
box 8 4 12 24
<< end >>
