magic
tech sky130l
timestamp 1731001260
<< m1 >>
rect 12 59 13 62
rect 9 54 13 59
rect 8 48 13 54
rect 36 59 37 62
rect 33 53 37 59
rect 47 59 48 62
rect 44 53 48 59
rect 16 50 20 52
rect 19 48 20 50
rect 24 49 37 53
rect 40 50 48 53
rect 55 56 56 59
rect 55 51 59 56
rect 51 50 59 51
rect 8 40 13 43
rect 16 34 19 47
rect 24 42 28 49
rect 40 48 44 50
rect 54 47 59 50
rect 51 45 54 47
rect 49 42 54 45
rect 60 40 65 43
rect 56 36 60 37
rect 23 25 26 36
rect 33 33 34 36
rect 37 33 38 36
rect 59 33 60 36
rect 67 33 68 36
rect 71 33 72 36
rect 8 15 12 20
rect 22 19 23 22
rect 26 19 27 22
rect 34 19 37 30
rect 56 23 60 33
rect 75 26 80 29
rect 8 12 9 15
rect 8 6 12 12
rect 41 15 44 23
rect 56 22 64 23
rect 41 11 44 12
rect 50 11 53 20
rect 56 19 61 22
rect 56 18 64 19
rect 56 12 60 18
rect 68 11 71 20
rect 8 3 9 6
<< m2c >>
rect 9 59 12 62
rect 33 59 36 62
rect 44 59 47 62
rect 16 47 19 50
rect 56 56 59 59
rect 51 47 54 50
rect 34 33 37 36
rect 56 33 59 36
rect 68 33 71 36
rect 23 19 26 22
rect 9 12 12 15
rect 41 12 44 15
rect 61 19 64 22
rect 9 3 12 6
<< m2 >>
rect 8 62 13 63
rect 8 59 9 62
rect 12 59 13 62
rect 8 58 13 59
rect 32 62 37 63
rect 32 59 33 62
rect 36 59 37 62
rect 32 58 37 59
rect 43 62 48 63
rect 43 59 44 62
rect 47 59 48 62
rect 43 58 48 59
rect 55 59 60 60
rect 55 56 56 59
rect 59 56 60 59
rect 55 55 60 56
rect 15 50 55 51
rect 15 47 16 50
rect 19 47 51 50
rect 54 47 55 50
rect 15 46 55 47
rect 8 39 65 44
rect 33 36 72 37
rect 33 33 34 36
rect 37 33 56 36
rect 59 33 68 36
rect 71 33 72 36
rect 33 32 72 33
rect 22 25 80 30
rect 22 22 65 23
rect 22 19 23 22
rect 26 19 61 22
rect 64 19 65 22
rect 22 18 65 19
rect 8 15 46 16
rect 8 12 9 15
rect 12 12 41 15
rect 44 12 46 15
rect 8 11 46 12
rect 49 11 72 16
rect 8 6 13 7
rect 8 3 9 6
rect 12 3 13 6
rect 8 2 13 3
<< labels >>
rlabel m2 s 12 59 13 62 6 A
port 1 nsew signal input
rlabel m2 s 9 59 12 62 6 A
port 1 nsew signal input
rlabel m2 s 8 58 13 59 6 A
port 1 nsew signal input
rlabel m2 s 8 59 9 62 6 A
port 1 nsew signal input
rlabel m2 s 8 62 13 63 6 A
port 1 nsew signal input
rlabel m2c s 9 59 12 62 6 A
port 1 nsew signal input
rlabel m1 s 12 59 13 62 6 A
port 1 nsew signal input
rlabel m1 s 10 50 13 53 6 A
port 1 nsew signal input
rlabel m1 s 9 54 13 59 6 A
port 1 nsew signal input
rlabel m1 s 9 59 12 62 6 A
port 1 nsew signal input
rlabel m1 s 8 48 13 50 6 A
port 1 nsew signal input
rlabel m1 s 8 50 10 53 6 A
port 1 nsew signal input
rlabel m1 s 8 53 13 54 6 A
port 1 nsew signal input
rlabel m2 s 47 59 48 62 6 B
port 2 nsew signal input
rlabel m2 s 44 59 47 62 6 B
port 2 nsew signal input
rlabel m2 s 43 58 48 59 6 B
port 2 nsew signal input
rlabel m2 s 43 59 44 62 6 B
port 2 nsew signal input
rlabel m2 s 43 62 48 63 6 B
port 2 nsew signal input
rlabel m2c s 44 59 47 62 6 B
port 2 nsew signal input
rlabel m1 s 47 59 48 62 6 B
port 2 nsew signal input
rlabel m1 s 47 50 48 53 6 B
port 2 nsew signal input
rlabel m1 s 44 53 48 59 6 B
port 2 nsew signal input
rlabel m1 s 44 59 47 62 6 B
port 2 nsew signal input
rlabel m1 s 44 50 47 53 6 B
port 2 nsew signal input
rlabel m1 s 40 48 44 53 6 B
port 2 nsew signal input
rlabel m2 s 36 59 37 62 6 S
port 3 nsew signal input
rlabel m2 s 33 59 36 62 6 S
port 3 nsew signal input
rlabel m2 s 32 58 37 59 6 S
port 3 nsew signal input
rlabel m2 s 32 59 33 62 6 S
port 3 nsew signal input
rlabel m2 s 32 62 37 63 6 S
port 3 nsew signal input
rlabel m2c s 33 59 36 62 6 S
port 3 nsew signal input
rlabel m1 s 36 59 37 62 6 S
port 3 nsew signal input
rlabel m1 s 33 53 37 59 6 S
port 3 nsew signal input
rlabel m1 s 33 59 36 62 6 S
port 3 nsew signal input
rlabel m1 s 36 50 37 53 6 S
port 3 nsew signal input
rlabel m1 s 27 43 28 46 6 S
port 3 nsew signal input
rlabel m1 s 33 50 36 53 6 S
port 3 nsew signal input
rlabel m1 s 24 42 28 43 6 S
port 3 nsew signal input
rlabel m1 s 24 43 27 46 6 S
port 3 nsew signal input
rlabel m1 s 24 46 28 49 6 S
port 3 nsew signal input
rlabel m1 s 24 49 37 50 6 S
port 3 nsew signal input
rlabel m1 s 24 50 33 53 6 S
port 3 nsew signal input
rlabel m2 s 71 33 72 36 6 Y
port 4 nsew signal output
rlabel m2 s 68 33 71 36 6 Y
port 4 nsew signal output
rlabel m2 s 59 33 68 36 6 Y
port 4 nsew signal output
rlabel m2 s 56 33 59 36 6 Y
port 4 nsew signal output
rlabel m2 s 37 33 56 36 6 Y
port 4 nsew signal output
rlabel m2 s 34 33 37 36 6 Y
port 4 nsew signal output
rlabel m2 s 64 19 65 22 6 Y
port 4 nsew signal output
rlabel m2 s 33 32 72 33 6 Y
port 4 nsew signal output
rlabel m2 s 33 33 34 36 6 Y
port 4 nsew signal output
rlabel m2 s 33 36 72 37 6 Y
port 4 nsew signal output
rlabel m2 s 61 19 64 22 6 Y
port 4 nsew signal output
rlabel m2 s 26 19 61 22 6 Y
port 4 nsew signal output
rlabel m2 s 23 19 26 22 6 Y
port 4 nsew signal output
rlabel m2 s 22 18 65 19 6 Y
port 4 nsew signal output
rlabel m2 s 22 19 23 22 6 Y
port 4 nsew signal output
rlabel m2 s 22 22 65 23 6 Y
port 4 nsew signal output
rlabel m2c s 68 33 71 36 6 Y
port 4 nsew signal output
rlabel m2c s 61 19 64 22 6 Y
port 4 nsew signal output
rlabel m2c s 56 33 59 36 6 Y
port 4 nsew signal output
rlabel m2c s 34 33 37 36 6 Y
port 4 nsew signal output
rlabel m2c s 23 19 26 22 6 Y
port 4 nsew signal output
rlabel m1 s 71 33 72 36 6 Y
port 4 nsew signal output
rlabel m1 s 68 33 71 36 6 Y
port 4 nsew signal output
rlabel m1 s 67 33 68 36 6 Y
port 4 nsew signal output
rlabel m1 s 61 19 64 22 6 Y
port 4 nsew signal output
rlabel m1 s 59 33 60 36 6 Y
port 4 nsew signal output
rlabel m1 s 56 12 60 18 6 Y
port 4 nsew signal output
rlabel m1 s 56 18 64 19 6 Y
port 4 nsew signal output
rlabel m1 s 56 19 61 22 6 Y
port 4 nsew signal output
rlabel m1 s 56 22 64 23 6 Y
port 4 nsew signal output
rlabel m1 s 56 23 60 33 6 Y
port 4 nsew signal output
rlabel m1 s 56 33 59 36 6 Y
port 4 nsew signal output
rlabel m1 s 56 36 60 37 6 Y
port 4 nsew signal output
rlabel m1 s 37 33 38 36 6 Y
port 4 nsew signal output
rlabel m1 s 34 33 37 36 6 Y
port 4 nsew signal output
rlabel m1 s 33 33 34 36 6 Y
port 4 nsew signal output
rlabel m1 s 26 19 27 22 6 Y
port 4 nsew signal output
rlabel m1 s 23 19 26 22 6 Y
port 4 nsew signal output
rlabel m1 s 22 19 23 22 6 Y
port 4 nsew signal output
rlabel m2 s 59 56 60 59 6 Vdd
port 5 nsew power input
rlabel m2 s 56 56 59 59 6 Vdd
port 5 nsew power input
rlabel m2 s 55 55 60 56 6 Vdd
port 5 nsew power input
rlabel m2 s 55 56 56 59 6 Vdd
port 5 nsew power input
rlabel m2 s 55 59 60 60 6 Vdd
port 5 nsew power input
rlabel m2 s 54 47 55 50 6 Vdd
port 5 nsew power input
rlabel m2 s 51 47 54 50 6 Vdd
port 5 nsew power input
rlabel m2 s 19 47 51 50 6 Vdd
port 5 nsew power input
rlabel m2 s 16 47 19 50 6 Vdd
port 5 nsew power input
rlabel m2 s 15 46 55 47 6 Vdd
port 5 nsew power input
rlabel m2 s 15 47 16 50 6 Vdd
port 5 nsew power input
rlabel m2 s 15 50 55 51 6 Vdd
port 5 nsew power input
rlabel m2c s 56 56 59 59 6 Vdd
port 5 nsew power input
rlabel m2c s 51 47 54 50 6 Vdd
port 5 nsew power input
rlabel m2c s 16 47 19 50 6 Vdd
port 5 nsew power input
rlabel m1 s 56 56 59 59 6 Vdd
port 5 nsew power input
rlabel m1 s 55 51 59 56 6 Vdd
port 5 nsew power input
rlabel m1 s 55 56 56 59 6 Vdd
port 5 nsew power input
rlabel m1 s 54 47 59 50 6 Vdd
port 5 nsew power input
rlabel m1 s 53 42 54 45 6 Vdd
port 5 nsew power input
rlabel m1 s 51 45 54 47 6 Vdd
port 5 nsew power input
rlabel m1 s 51 47 54 50 6 Vdd
port 5 nsew power input
rlabel m1 s 51 50 59 51 6 Vdd
port 5 nsew power input
rlabel m1 s 50 42 53 45 6 Vdd
port 5 nsew power input
rlabel m1 s 49 42 50 45 6 Vdd
port 5 nsew power input
rlabel m1 s 19 48 20 50 6 Vdd
port 5 nsew power input
rlabel m1 s 16 47 19 50 6 Vdd
port 5 nsew power input
rlabel m1 s 16 50 20 52 6 Vdd
port 5 nsew power input
rlabel m1 s 16 34 19 35 6 Vdd
port 5 nsew power input
rlabel m1 s 16 35 19 38 6 Vdd
port 5 nsew power input
rlabel m1 s 16 38 19 47 6 Vdd
port 5 nsew power input
rlabel m2 s 44 12 46 15 6 GND
port 6 nsew ground input
rlabel m2 s 41 12 44 15 6 GND
port 6 nsew ground input
rlabel m2 s 12 3 13 6 6 GND
port 6 nsew ground input
rlabel m2 s 12 12 41 15 6 GND
port 6 nsew ground input
rlabel m2 s 9 3 12 6 6 GND
port 6 nsew ground input
rlabel m2 s 9 12 12 15 6 GND
port 6 nsew ground input
rlabel m2 s 8 2 13 3 6 GND
port 6 nsew ground input
rlabel m2 s 8 3 9 6 6 GND
port 6 nsew ground input
rlabel m2 s 8 6 13 7 6 GND
port 6 nsew ground input
rlabel m2 s 8 11 46 12 6 GND
port 6 nsew ground input
rlabel m2 s 8 12 9 15 6 GND
port 6 nsew ground input
rlabel m2 s 8 15 46 16 6 GND
port 6 nsew ground input
rlabel m2c s 41 12 44 15 6 GND
port 6 nsew ground input
rlabel m2c s 9 3 12 6 6 GND
port 6 nsew ground input
rlabel m2c s 9 12 12 15 6 GND
port 6 nsew ground input
rlabel m1 s 41 11 44 12 6 GND
port 6 nsew ground input
rlabel m1 s 41 12 44 15 6 GND
port 6 nsew ground input
rlabel m1 s 41 15 44 19 6 GND
port 6 nsew ground input
rlabel m1 s 41 19 44 22 6 GND
port 6 nsew ground input
rlabel m1 s 41 22 44 23 6 GND
port 6 nsew ground input
rlabel m1 s 9 3 12 6 6 GND
port 6 nsew ground input
rlabel m1 s 9 12 12 15 6 GND
port 6 nsew ground input
rlabel m1 s 9 16 12 19 6 GND
port 6 nsew ground input
rlabel m1 s 8 3 9 6 6 GND
port 6 nsew ground input
rlabel m1 s 8 6 12 12 6 GND
port 6 nsew ground input
rlabel m1 s 8 12 9 15 6 GND
port 6 nsew ground input
rlabel m1 s 8 15 12 16 6 GND
port 6 nsew ground input
rlabel m1 s 8 16 9 19 6 GND
port 6 nsew ground input
rlabel m1 s 8 19 12 20 6 GND
port 6 nsew ground input
<< properties >>
string LEFsite CoreSite
string LEFclass CORE
string FIXED_BBOX 0 0 88 64
string LEFsymmetry X Y
string LEFview TRUE
<< end >>
