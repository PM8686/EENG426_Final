magic
tech sky130l
timestamp 1731220619
<< m2 >>
rect 1342 2196 1348 2197
rect 1342 2192 1343 2196
rect 1347 2192 1348 2196
rect 1342 2191 1348 2192
rect 1382 2196 1388 2197
rect 1382 2192 1383 2196
rect 1387 2192 1388 2196
rect 1382 2191 1388 2192
rect 1422 2196 1428 2197
rect 1422 2192 1423 2196
rect 1427 2192 1428 2196
rect 1422 2191 1428 2192
rect 1462 2196 1468 2197
rect 1462 2192 1463 2196
rect 1467 2192 1468 2196
rect 1462 2191 1468 2192
rect 1502 2196 1508 2197
rect 1502 2192 1503 2196
rect 1507 2192 1508 2196
rect 1502 2191 1508 2192
rect 1542 2196 1548 2197
rect 1542 2192 1543 2196
rect 1547 2192 1548 2196
rect 1542 2191 1548 2192
rect 1582 2196 1588 2197
rect 1582 2192 1583 2196
rect 1587 2192 1588 2196
rect 1582 2191 1588 2192
rect 1622 2196 1628 2197
rect 1622 2192 1623 2196
rect 1627 2192 1628 2196
rect 1622 2191 1628 2192
rect 1662 2196 1668 2197
rect 1662 2192 1663 2196
rect 1667 2192 1668 2196
rect 1662 2191 1668 2192
rect 1702 2196 1708 2197
rect 1702 2192 1703 2196
rect 1707 2192 1708 2196
rect 1702 2191 1708 2192
rect 1742 2196 1748 2197
rect 1742 2192 1743 2196
rect 1747 2192 1748 2196
rect 1742 2191 1748 2192
rect 1782 2196 1788 2197
rect 1782 2192 1783 2196
rect 1787 2192 1788 2196
rect 1782 2191 1788 2192
rect 1822 2196 1828 2197
rect 1822 2192 1823 2196
rect 1827 2192 1828 2196
rect 1822 2191 1828 2192
rect 1134 2188 1140 2189
rect 1134 2184 1135 2188
rect 1139 2184 1140 2188
rect 1134 2183 1140 2184
rect 2118 2188 2124 2189
rect 2118 2184 2119 2188
rect 2123 2184 2124 2188
rect 2118 2183 2124 2184
rect 1134 2171 1140 2172
rect 1134 2167 1135 2171
rect 1139 2167 1140 2171
rect 2118 2171 2124 2172
rect 1134 2166 1140 2167
rect 1342 2168 1348 2169
rect 1342 2164 1343 2168
rect 1347 2164 1348 2168
rect 1342 2163 1348 2164
rect 1382 2168 1388 2169
rect 1382 2164 1383 2168
rect 1387 2164 1388 2168
rect 1382 2163 1388 2164
rect 1422 2168 1428 2169
rect 1422 2164 1423 2168
rect 1427 2164 1428 2168
rect 1422 2163 1428 2164
rect 1462 2168 1468 2169
rect 1462 2164 1463 2168
rect 1467 2164 1468 2168
rect 1462 2163 1468 2164
rect 1502 2168 1508 2169
rect 1502 2164 1503 2168
rect 1507 2164 1508 2168
rect 1502 2163 1508 2164
rect 1542 2168 1548 2169
rect 1542 2164 1543 2168
rect 1547 2164 1548 2168
rect 1542 2163 1548 2164
rect 1582 2168 1588 2169
rect 1582 2164 1583 2168
rect 1587 2164 1588 2168
rect 1582 2163 1588 2164
rect 1622 2168 1628 2169
rect 1622 2164 1623 2168
rect 1627 2164 1628 2168
rect 1622 2163 1628 2164
rect 1662 2168 1668 2169
rect 1662 2164 1663 2168
rect 1667 2164 1668 2168
rect 1662 2163 1668 2164
rect 1702 2168 1708 2169
rect 1702 2164 1703 2168
rect 1707 2164 1708 2168
rect 1702 2163 1708 2164
rect 1742 2168 1748 2169
rect 1742 2164 1743 2168
rect 1747 2164 1748 2168
rect 1742 2163 1748 2164
rect 1782 2168 1788 2169
rect 1782 2164 1783 2168
rect 1787 2164 1788 2168
rect 1782 2163 1788 2164
rect 1822 2168 1828 2169
rect 1822 2164 1823 2168
rect 1827 2164 1828 2168
rect 2118 2167 2119 2171
rect 2123 2167 2124 2171
rect 2118 2166 2124 2167
rect 1822 2163 1828 2164
rect 1286 2156 1292 2157
rect 1134 2153 1140 2154
rect 1134 2149 1135 2153
rect 1139 2149 1140 2153
rect 1286 2152 1287 2156
rect 1291 2152 1292 2156
rect 1286 2151 1292 2152
rect 1326 2156 1332 2157
rect 1326 2152 1327 2156
rect 1331 2152 1332 2156
rect 1326 2151 1332 2152
rect 1366 2156 1372 2157
rect 1366 2152 1367 2156
rect 1371 2152 1372 2156
rect 1366 2151 1372 2152
rect 1414 2156 1420 2157
rect 1414 2152 1415 2156
rect 1419 2152 1420 2156
rect 1414 2151 1420 2152
rect 1462 2156 1468 2157
rect 1462 2152 1463 2156
rect 1467 2152 1468 2156
rect 1462 2151 1468 2152
rect 1518 2156 1524 2157
rect 1518 2152 1519 2156
rect 1523 2152 1524 2156
rect 1518 2151 1524 2152
rect 1574 2156 1580 2157
rect 1574 2152 1575 2156
rect 1579 2152 1580 2156
rect 1574 2151 1580 2152
rect 1622 2156 1628 2157
rect 1622 2152 1623 2156
rect 1627 2152 1628 2156
rect 1622 2151 1628 2152
rect 1670 2156 1676 2157
rect 1670 2152 1671 2156
rect 1675 2152 1676 2156
rect 1670 2151 1676 2152
rect 1718 2156 1724 2157
rect 1718 2152 1719 2156
rect 1723 2152 1724 2156
rect 1718 2151 1724 2152
rect 1774 2156 1780 2157
rect 1774 2152 1775 2156
rect 1779 2152 1780 2156
rect 1774 2151 1780 2152
rect 1830 2156 1836 2157
rect 1830 2152 1831 2156
rect 1835 2152 1836 2156
rect 1830 2151 1836 2152
rect 1886 2156 1892 2157
rect 1886 2152 1887 2156
rect 1891 2152 1892 2156
rect 1886 2151 1892 2152
rect 2118 2153 2124 2154
rect 1134 2148 1140 2149
rect 2118 2149 2119 2153
rect 2123 2149 2124 2153
rect 2118 2148 2124 2149
rect 1134 2136 1140 2137
rect 1134 2132 1135 2136
rect 1139 2132 1140 2136
rect 1134 2131 1140 2132
rect 2118 2136 2124 2137
rect 2118 2132 2119 2136
rect 2123 2132 2124 2136
rect 2118 2131 2124 2132
rect 1286 2128 1292 2129
rect 1286 2124 1287 2128
rect 1291 2124 1292 2128
rect 1286 2123 1292 2124
rect 1326 2128 1332 2129
rect 1326 2124 1327 2128
rect 1331 2124 1332 2128
rect 1326 2123 1332 2124
rect 1366 2128 1372 2129
rect 1366 2124 1367 2128
rect 1371 2124 1372 2128
rect 1366 2123 1372 2124
rect 1414 2128 1420 2129
rect 1414 2124 1415 2128
rect 1419 2124 1420 2128
rect 1414 2123 1420 2124
rect 1462 2128 1468 2129
rect 1462 2124 1463 2128
rect 1467 2124 1468 2128
rect 1462 2123 1468 2124
rect 1518 2128 1524 2129
rect 1518 2124 1519 2128
rect 1523 2124 1524 2128
rect 1518 2123 1524 2124
rect 1574 2128 1580 2129
rect 1574 2124 1575 2128
rect 1579 2124 1580 2128
rect 1574 2123 1580 2124
rect 1622 2128 1628 2129
rect 1622 2124 1623 2128
rect 1627 2124 1628 2128
rect 1622 2123 1628 2124
rect 1670 2128 1676 2129
rect 1670 2124 1671 2128
rect 1675 2124 1676 2128
rect 1670 2123 1676 2124
rect 1718 2128 1724 2129
rect 1718 2124 1719 2128
rect 1723 2124 1724 2128
rect 1718 2123 1724 2124
rect 1774 2128 1780 2129
rect 1774 2124 1775 2128
rect 1779 2124 1780 2128
rect 1774 2123 1780 2124
rect 1830 2128 1836 2129
rect 1830 2124 1831 2128
rect 1835 2124 1836 2128
rect 1830 2123 1836 2124
rect 1886 2128 1892 2129
rect 1886 2124 1887 2128
rect 1891 2124 1892 2128
rect 1886 2123 1892 2124
rect 1222 2088 1228 2089
rect 1222 2084 1223 2088
rect 1227 2084 1228 2088
rect 1222 2083 1228 2084
rect 1278 2088 1284 2089
rect 1278 2084 1279 2088
rect 1283 2084 1284 2088
rect 1278 2083 1284 2084
rect 1342 2088 1348 2089
rect 1342 2084 1343 2088
rect 1347 2084 1348 2088
rect 1342 2083 1348 2084
rect 1422 2088 1428 2089
rect 1422 2084 1423 2088
rect 1427 2084 1428 2088
rect 1422 2083 1428 2084
rect 1502 2088 1508 2089
rect 1502 2084 1503 2088
rect 1507 2084 1508 2088
rect 1502 2083 1508 2084
rect 1582 2088 1588 2089
rect 1582 2084 1583 2088
rect 1587 2084 1588 2088
rect 1582 2083 1588 2084
rect 1662 2088 1668 2089
rect 1662 2084 1663 2088
rect 1667 2084 1668 2088
rect 1662 2083 1668 2084
rect 1742 2088 1748 2089
rect 1742 2084 1743 2088
rect 1747 2084 1748 2088
rect 1742 2083 1748 2084
rect 1830 2088 1836 2089
rect 1830 2084 1831 2088
rect 1835 2084 1836 2088
rect 1830 2083 1836 2084
rect 1918 2088 1924 2089
rect 1918 2084 1919 2088
rect 1923 2084 1924 2088
rect 1918 2083 1924 2084
rect 2006 2088 2012 2089
rect 2006 2084 2007 2088
rect 2011 2084 2012 2088
rect 2006 2083 2012 2084
rect 2070 2088 2076 2089
rect 2070 2084 2071 2088
rect 2075 2084 2076 2088
rect 2070 2083 2076 2084
rect 1134 2080 1140 2081
rect 1134 2076 1135 2080
rect 1139 2076 1140 2080
rect 1134 2075 1140 2076
rect 2118 2080 2124 2081
rect 2118 2076 2119 2080
rect 2123 2076 2124 2080
rect 2118 2075 2124 2076
rect 1134 2063 1140 2064
rect 1134 2059 1135 2063
rect 1139 2059 1140 2063
rect 2118 2063 2124 2064
rect 1134 2058 1140 2059
rect 1222 2060 1228 2061
rect 1222 2056 1223 2060
rect 1227 2056 1228 2060
rect 1222 2055 1228 2056
rect 1278 2060 1284 2061
rect 1278 2056 1279 2060
rect 1283 2056 1284 2060
rect 1278 2055 1284 2056
rect 1342 2060 1348 2061
rect 1342 2056 1343 2060
rect 1347 2056 1348 2060
rect 1342 2055 1348 2056
rect 1422 2060 1428 2061
rect 1422 2056 1423 2060
rect 1427 2056 1428 2060
rect 1422 2055 1428 2056
rect 1502 2060 1508 2061
rect 1502 2056 1503 2060
rect 1507 2056 1508 2060
rect 1502 2055 1508 2056
rect 1582 2060 1588 2061
rect 1582 2056 1583 2060
rect 1587 2056 1588 2060
rect 1582 2055 1588 2056
rect 1662 2060 1668 2061
rect 1662 2056 1663 2060
rect 1667 2056 1668 2060
rect 1662 2055 1668 2056
rect 1742 2060 1748 2061
rect 1742 2056 1743 2060
rect 1747 2056 1748 2060
rect 1742 2055 1748 2056
rect 1830 2060 1836 2061
rect 1830 2056 1831 2060
rect 1835 2056 1836 2060
rect 1830 2055 1836 2056
rect 1918 2060 1924 2061
rect 1918 2056 1919 2060
rect 1923 2056 1924 2060
rect 1918 2055 1924 2056
rect 2006 2060 2012 2061
rect 2006 2056 2007 2060
rect 2011 2056 2012 2060
rect 2006 2055 2012 2056
rect 2070 2060 2076 2061
rect 2070 2056 2071 2060
rect 2075 2056 2076 2060
rect 2118 2059 2119 2063
rect 2123 2059 2124 2063
rect 2118 2058 2124 2059
rect 2070 2055 2076 2056
rect 1182 2048 1188 2049
rect 1134 2045 1140 2046
rect 1134 2041 1135 2045
rect 1139 2041 1140 2045
rect 1182 2044 1183 2048
rect 1187 2044 1188 2048
rect 1182 2043 1188 2044
rect 1238 2048 1244 2049
rect 1238 2044 1239 2048
rect 1243 2044 1244 2048
rect 1238 2043 1244 2044
rect 1310 2048 1316 2049
rect 1310 2044 1311 2048
rect 1315 2044 1316 2048
rect 1310 2043 1316 2044
rect 1398 2048 1404 2049
rect 1398 2044 1399 2048
rect 1403 2044 1404 2048
rect 1398 2043 1404 2044
rect 1486 2048 1492 2049
rect 1486 2044 1487 2048
rect 1491 2044 1492 2048
rect 1486 2043 1492 2044
rect 1582 2048 1588 2049
rect 1582 2044 1583 2048
rect 1587 2044 1588 2048
rect 1582 2043 1588 2044
rect 1670 2048 1676 2049
rect 1670 2044 1671 2048
rect 1675 2044 1676 2048
rect 1670 2043 1676 2044
rect 1758 2048 1764 2049
rect 1758 2044 1759 2048
rect 1763 2044 1764 2048
rect 1758 2043 1764 2044
rect 1838 2048 1844 2049
rect 1838 2044 1839 2048
rect 1843 2044 1844 2048
rect 1838 2043 1844 2044
rect 1918 2048 1924 2049
rect 1918 2044 1919 2048
rect 1923 2044 1924 2048
rect 1918 2043 1924 2044
rect 2006 2048 2012 2049
rect 2006 2044 2007 2048
rect 2011 2044 2012 2048
rect 2006 2043 2012 2044
rect 2070 2048 2076 2049
rect 2070 2044 2071 2048
rect 2075 2044 2076 2048
rect 2070 2043 2076 2044
rect 2118 2045 2124 2046
rect 1134 2040 1140 2041
rect 2118 2041 2119 2045
rect 2123 2041 2124 2045
rect 2118 2040 2124 2041
rect 1134 2028 1140 2029
rect 1134 2024 1135 2028
rect 1139 2024 1140 2028
rect 1134 2023 1140 2024
rect 2118 2028 2124 2029
rect 2118 2024 2119 2028
rect 2123 2024 2124 2028
rect 2118 2023 2124 2024
rect 1182 2020 1188 2021
rect 190 2016 196 2017
rect 190 2012 191 2016
rect 195 2012 196 2016
rect 190 2011 196 2012
rect 230 2016 236 2017
rect 230 2012 231 2016
rect 235 2012 236 2016
rect 230 2011 236 2012
rect 286 2016 292 2017
rect 286 2012 287 2016
rect 291 2012 292 2016
rect 286 2011 292 2012
rect 350 2016 356 2017
rect 350 2012 351 2016
rect 355 2012 356 2016
rect 350 2011 356 2012
rect 422 2016 428 2017
rect 422 2012 423 2016
rect 427 2012 428 2016
rect 422 2011 428 2012
rect 494 2016 500 2017
rect 494 2012 495 2016
rect 499 2012 500 2016
rect 494 2011 500 2012
rect 574 2016 580 2017
rect 574 2012 575 2016
rect 579 2012 580 2016
rect 574 2011 580 2012
rect 646 2016 652 2017
rect 646 2012 647 2016
rect 651 2012 652 2016
rect 646 2011 652 2012
rect 718 2016 724 2017
rect 718 2012 719 2016
rect 723 2012 724 2016
rect 718 2011 724 2012
rect 782 2016 788 2017
rect 782 2012 783 2016
rect 787 2012 788 2016
rect 782 2011 788 2012
rect 838 2016 844 2017
rect 838 2012 839 2016
rect 843 2012 844 2016
rect 838 2011 844 2012
rect 894 2016 900 2017
rect 894 2012 895 2016
rect 899 2012 900 2016
rect 894 2011 900 2012
rect 950 2016 956 2017
rect 950 2012 951 2016
rect 955 2012 956 2016
rect 950 2011 956 2012
rect 1006 2016 1012 2017
rect 1006 2012 1007 2016
rect 1011 2012 1012 2016
rect 1006 2011 1012 2012
rect 1046 2016 1052 2017
rect 1046 2012 1047 2016
rect 1051 2012 1052 2016
rect 1182 2016 1183 2020
rect 1187 2016 1188 2020
rect 1182 2015 1188 2016
rect 1238 2020 1244 2021
rect 1238 2016 1239 2020
rect 1243 2016 1244 2020
rect 1238 2015 1244 2016
rect 1310 2020 1316 2021
rect 1310 2016 1311 2020
rect 1315 2016 1316 2020
rect 1310 2015 1316 2016
rect 1398 2020 1404 2021
rect 1398 2016 1399 2020
rect 1403 2016 1404 2020
rect 1398 2015 1404 2016
rect 1486 2020 1492 2021
rect 1486 2016 1487 2020
rect 1491 2016 1492 2020
rect 1486 2015 1492 2016
rect 1582 2020 1588 2021
rect 1582 2016 1583 2020
rect 1587 2016 1588 2020
rect 1582 2015 1588 2016
rect 1670 2020 1676 2021
rect 1670 2016 1671 2020
rect 1675 2016 1676 2020
rect 1670 2015 1676 2016
rect 1758 2020 1764 2021
rect 1758 2016 1759 2020
rect 1763 2016 1764 2020
rect 1758 2015 1764 2016
rect 1838 2020 1844 2021
rect 1838 2016 1839 2020
rect 1843 2016 1844 2020
rect 1838 2015 1844 2016
rect 1918 2020 1924 2021
rect 1918 2016 1919 2020
rect 1923 2016 1924 2020
rect 1918 2015 1924 2016
rect 2006 2020 2012 2021
rect 2006 2016 2007 2020
rect 2011 2016 2012 2020
rect 2006 2015 2012 2016
rect 2070 2020 2076 2021
rect 2070 2016 2071 2020
rect 2075 2016 2076 2020
rect 2070 2015 2076 2016
rect 1046 2011 1052 2012
rect 110 2008 116 2009
rect 110 2004 111 2008
rect 115 2004 116 2008
rect 110 2003 116 2004
rect 1094 2008 1100 2009
rect 1094 2004 1095 2008
rect 1099 2004 1100 2008
rect 1094 2003 1100 2004
rect 110 1991 116 1992
rect 110 1987 111 1991
rect 115 1987 116 1991
rect 1094 1991 1100 1992
rect 110 1986 116 1987
rect 190 1988 196 1989
rect 190 1984 191 1988
rect 195 1984 196 1988
rect 190 1983 196 1984
rect 230 1988 236 1989
rect 230 1984 231 1988
rect 235 1984 236 1988
rect 230 1983 236 1984
rect 286 1988 292 1989
rect 286 1984 287 1988
rect 291 1984 292 1988
rect 286 1983 292 1984
rect 350 1988 356 1989
rect 350 1984 351 1988
rect 355 1984 356 1988
rect 350 1983 356 1984
rect 422 1988 428 1989
rect 422 1984 423 1988
rect 427 1984 428 1988
rect 422 1983 428 1984
rect 494 1988 500 1989
rect 494 1984 495 1988
rect 499 1984 500 1988
rect 494 1983 500 1984
rect 574 1988 580 1989
rect 574 1984 575 1988
rect 579 1984 580 1988
rect 574 1983 580 1984
rect 646 1988 652 1989
rect 646 1984 647 1988
rect 651 1984 652 1988
rect 646 1983 652 1984
rect 718 1988 724 1989
rect 718 1984 719 1988
rect 723 1984 724 1988
rect 718 1983 724 1984
rect 782 1988 788 1989
rect 782 1984 783 1988
rect 787 1984 788 1988
rect 782 1983 788 1984
rect 838 1988 844 1989
rect 838 1984 839 1988
rect 843 1984 844 1988
rect 838 1983 844 1984
rect 894 1988 900 1989
rect 894 1984 895 1988
rect 899 1984 900 1988
rect 894 1983 900 1984
rect 950 1988 956 1989
rect 950 1984 951 1988
rect 955 1984 956 1988
rect 950 1983 956 1984
rect 1006 1988 1012 1989
rect 1006 1984 1007 1988
rect 1011 1984 1012 1988
rect 1006 1983 1012 1984
rect 1046 1988 1052 1989
rect 1046 1984 1047 1988
rect 1051 1984 1052 1988
rect 1094 1987 1095 1991
rect 1099 1987 1100 1991
rect 1094 1986 1100 1987
rect 1046 1983 1052 1984
rect 1302 1984 1308 1985
rect 1302 1980 1303 1984
rect 1307 1980 1308 1984
rect 1302 1979 1308 1980
rect 1382 1984 1388 1985
rect 1382 1980 1383 1984
rect 1387 1980 1388 1984
rect 1382 1979 1388 1980
rect 1462 1984 1468 1985
rect 1462 1980 1463 1984
rect 1467 1980 1468 1984
rect 1462 1979 1468 1980
rect 1542 1984 1548 1985
rect 1542 1980 1543 1984
rect 1547 1980 1548 1984
rect 1542 1979 1548 1980
rect 1614 1984 1620 1985
rect 1614 1980 1615 1984
rect 1619 1980 1620 1984
rect 1614 1979 1620 1980
rect 1686 1984 1692 1985
rect 1686 1980 1687 1984
rect 1691 1980 1692 1984
rect 1686 1979 1692 1980
rect 1750 1984 1756 1985
rect 1750 1980 1751 1984
rect 1755 1980 1756 1984
rect 1750 1979 1756 1980
rect 1814 1984 1820 1985
rect 1814 1980 1815 1984
rect 1819 1980 1820 1984
rect 1814 1979 1820 1980
rect 1878 1984 1884 1985
rect 1878 1980 1879 1984
rect 1883 1980 1884 1984
rect 1878 1979 1884 1980
rect 1950 1984 1956 1985
rect 1950 1980 1951 1984
rect 1955 1980 1956 1984
rect 1950 1979 1956 1980
rect 2022 1984 2028 1985
rect 2022 1980 2023 1984
rect 2027 1980 2028 1984
rect 2022 1979 2028 1980
rect 2070 1984 2076 1985
rect 2070 1980 2071 1984
rect 2075 1980 2076 1984
rect 2070 1979 2076 1980
rect 190 1976 196 1977
rect 110 1973 116 1974
rect 110 1969 111 1973
rect 115 1969 116 1973
rect 190 1972 191 1976
rect 195 1972 196 1976
rect 190 1971 196 1972
rect 246 1976 252 1977
rect 246 1972 247 1976
rect 251 1972 252 1976
rect 246 1971 252 1972
rect 310 1976 316 1977
rect 310 1972 311 1976
rect 315 1972 316 1976
rect 310 1971 316 1972
rect 374 1976 380 1977
rect 374 1972 375 1976
rect 379 1972 380 1976
rect 374 1971 380 1972
rect 446 1976 452 1977
rect 446 1972 447 1976
rect 451 1972 452 1976
rect 446 1971 452 1972
rect 518 1976 524 1977
rect 518 1972 519 1976
rect 523 1972 524 1976
rect 518 1971 524 1972
rect 590 1976 596 1977
rect 590 1972 591 1976
rect 595 1972 596 1976
rect 590 1971 596 1972
rect 654 1976 660 1977
rect 654 1972 655 1976
rect 659 1972 660 1976
rect 654 1971 660 1972
rect 718 1976 724 1977
rect 718 1972 719 1976
rect 723 1972 724 1976
rect 718 1971 724 1972
rect 774 1976 780 1977
rect 774 1972 775 1976
rect 779 1972 780 1976
rect 774 1971 780 1972
rect 822 1976 828 1977
rect 822 1972 823 1976
rect 827 1972 828 1976
rect 822 1971 828 1972
rect 870 1976 876 1977
rect 870 1972 871 1976
rect 875 1972 876 1976
rect 870 1971 876 1972
rect 918 1976 924 1977
rect 918 1972 919 1976
rect 923 1972 924 1976
rect 918 1971 924 1972
rect 966 1976 972 1977
rect 966 1972 967 1976
rect 971 1972 972 1976
rect 966 1971 972 1972
rect 1006 1976 1012 1977
rect 1006 1972 1007 1976
rect 1011 1972 1012 1976
rect 1006 1971 1012 1972
rect 1046 1976 1052 1977
rect 1046 1972 1047 1976
rect 1051 1972 1052 1976
rect 1134 1976 1140 1977
rect 1046 1971 1052 1972
rect 1094 1973 1100 1974
rect 110 1968 116 1969
rect 1094 1969 1095 1973
rect 1099 1969 1100 1973
rect 1134 1972 1135 1976
rect 1139 1972 1140 1976
rect 1134 1971 1140 1972
rect 2118 1976 2124 1977
rect 2118 1972 2119 1976
rect 2123 1972 2124 1976
rect 2118 1971 2124 1972
rect 1094 1968 1100 1969
rect 1134 1959 1140 1960
rect 110 1956 116 1957
rect 110 1952 111 1956
rect 115 1952 116 1956
rect 110 1951 116 1952
rect 1094 1956 1100 1957
rect 1094 1952 1095 1956
rect 1099 1952 1100 1956
rect 1134 1955 1135 1959
rect 1139 1955 1140 1959
rect 2118 1959 2124 1960
rect 1134 1954 1140 1955
rect 1302 1956 1308 1957
rect 1094 1951 1100 1952
rect 1302 1952 1303 1956
rect 1307 1952 1308 1956
rect 1302 1951 1308 1952
rect 1382 1956 1388 1957
rect 1382 1952 1383 1956
rect 1387 1952 1388 1956
rect 1382 1951 1388 1952
rect 1462 1956 1468 1957
rect 1462 1952 1463 1956
rect 1467 1952 1468 1956
rect 1462 1951 1468 1952
rect 1542 1956 1548 1957
rect 1542 1952 1543 1956
rect 1547 1952 1548 1956
rect 1542 1951 1548 1952
rect 1614 1956 1620 1957
rect 1614 1952 1615 1956
rect 1619 1952 1620 1956
rect 1614 1951 1620 1952
rect 1686 1956 1692 1957
rect 1686 1952 1687 1956
rect 1691 1952 1692 1956
rect 1686 1951 1692 1952
rect 1750 1956 1756 1957
rect 1750 1952 1751 1956
rect 1755 1952 1756 1956
rect 1750 1951 1756 1952
rect 1814 1956 1820 1957
rect 1814 1952 1815 1956
rect 1819 1952 1820 1956
rect 1814 1951 1820 1952
rect 1878 1956 1884 1957
rect 1878 1952 1879 1956
rect 1883 1952 1884 1956
rect 1878 1951 1884 1952
rect 1950 1956 1956 1957
rect 1950 1952 1951 1956
rect 1955 1952 1956 1956
rect 1950 1951 1956 1952
rect 2022 1956 2028 1957
rect 2022 1952 2023 1956
rect 2027 1952 2028 1956
rect 2022 1951 2028 1952
rect 2070 1956 2076 1957
rect 2070 1952 2071 1956
rect 2075 1952 2076 1956
rect 2118 1955 2119 1959
rect 2123 1955 2124 1959
rect 2118 1954 2124 1955
rect 2070 1951 2076 1952
rect 190 1948 196 1949
rect 190 1944 191 1948
rect 195 1944 196 1948
rect 190 1943 196 1944
rect 246 1948 252 1949
rect 246 1944 247 1948
rect 251 1944 252 1948
rect 246 1943 252 1944
rect 310 1948 316 1949
rect 310 1944 311 1948
rect 315 1944 316 1948
rect 310 1943 316 1944
rect 374 1948 380 1949
rect 374 1944 375 1948
rect 379 1944 380 1948
rect 374 1943 380 1944
rect 446 1948 452 1949
rect 446 1944 447 1948
rect 451 1944 452 1948
rect 446 1943 452 1944
rect 518 1948 524 1949
rect 518 1944 519 1948
rect 523 1944 524 1948
rect 518 1943 524 1944
rect 590 1948 596 1949
rect 590 1944 591 1948
rect 595 1944 596 1948
rect 590 1943 596 1944
rect 654 1948 660 1949
rect 654 1944 655 1948
rect 659 1944 660 1948
rect 654 1943 660 1944
rect 718 1948 724 1949
rect 718 1944 719 1948
rect 723 1944 724 1948
rect 718 1943 724 1944
rect 774 1948 780 1949
rect 774 1944 775 1948
rect 779 1944 780 1948
rect 774 1943 780 1944
rect 822 1948 828 1949
rect 822 1944 823 1948
rect 827 1944 828 1948
rect 822 1943 828 1944
rect 870 1948 876 1949
rect 870 1944 871 1948
rect 875 1944 876 1948
rect 870 1943 876 1944
rect 918 1948 924 1949
rect 918 1944 919 1948
rect 923 1944 924 1948
rect 918 1943 924 1944
rect 966 1948 972 1949
rect 966 1944 967 1948
rect 971 1944 972 1948
rect 966 1943 972 1944
rect 1006 1948 1012 1949
rect 1006 1944 1007 1948
rect 1011 1944 1012 1948
rect 1006 1943 1012 1944
rect 1046 1948 1052 1949
rect 1046 1944 1047 1948
rect 1051 1944 1052 1948
rect 1046 1943 1052 1944
rect 1158 1940 1164 1941
rect 1134 1937 1140 1938
rect 1134 1933 1135 1937
rect 1139 1933 1140 1937
rect 1158 1936 1159 1940
rect 1163 1936 1164 1940
rect 1158 1935 1164 1936
rect 1222 1940 1228 1941
rect 1222 1936 1223 1940
rect 1227 1936 1228 1940
rect 1222 1935 1228 1936
rect 1302 1940 1308 1941
rect 1302 1936 1303 1940
rect 1307 1936 1308 1940
rect 1302 1935 1308 1936
rect 1382 1940 1388 1941
rect 1382 1936 1383 1940
rect 1387 1936 1388 1940
rect 1382 1935 1388 1936
rect 1462 1940 1468 1941
rect 1462 1936 1463 1940
rect 1467 1936 1468 1940
rect 1462 1935 1468 1936
rect 1534 1940 1540 1941
rect 1534 1936 1535 1940
rect 1539 1936 1540 1940
rect 1534 1935 1540 1936
rect 1614 1940 1620 1941
rect 1614 1936 1615 1940
rect 1619 1936 1620 1940
rect 1614 1935 1620 1936
rect 1694 1940 1700 1941
rect 1694 1936 1695 1940
rect 1699 1936 1700 1940
rect 1694 1935 1700 1936
rect 1782 1940 1788 1941
rect 1782 1936 1783 1940
rect 1787 1936 1788 1940
rect 1782 1935 1788 1936
rect 1878 1940 1884 1941
rect 1878 1936 1879 1940
rect 1883 1936 1884 1940
rect 1878 1935 1884 1936
rect 1982 1940 1988 1941
rect 1982 1936 1983 1940
rect 1987 1936 1988 1940
rect 1982 1935 1988 1936
rect 2070 1940 2076 1941
rect 2070 1936 2071 1940
rect 2075 1936 2076 1940
rect 2070 1935 2076 1936
rect 2118 1937 2124 1938
rect 1134 1932 1140 1933
rect 2118 1933 2119 1937
rect 2123 1933 2124 1937
rect 2118 1932 2124 1933
rect 1134 1920 1140 1921
rect 1134 1916 1135 1920
rect 1139 1916 1140 1920
rect 1134 1915 1140 1916
rect 2118 1920 2124 1921
rect 2118 1916 2119 1920
rect 2123 1916 2124 1920
rect 2118 1915 2124 1916
rect 134 1912 140 1913
rect 134 1908 135 1912
rect 139 1908 140 1912
rect 134 1907 140 1908
rect 174 1912 180 1913
rect 174 1908 175 1912
rect 179 1908 180 1912
rect 174 1907 180 1908
rect 230 1912 236 1913
rect 230 1908 231 1912
rect 235 1908 236 1912
rect 230 1907 236 1908
rect 294 1912 300 1913
rect 294 1908 295 1912
rect 299 1908 300 1912
rect 294 1907 300 1908
rect 366 1912 372 1913
rect 366 1908 367 1912
rect 371 1908 372 1912
rect 366 1907 372 1908
rect 430 1912 436 1913
rect 430 1908 431 1912
rect 435 1908 436 1912
rect 430 1907 436 1908
rect 494 1912 500 1913
rect 494 1908 495 1912
rect 499 1908 500 1912
rect 494 1907 500 1908
rect 558 1912 564 1913
rect 558 1908 559 1912
rect 563 1908 564 1912
rect 558 1907 564 1908
rect 614 1912 620 1913
rect 614 1908 615 1912
rect 619 1908 620 1912
rect 614 1907 620 1908
rect 670 1912 676 1913
rect 670 1908 671 1912
rect 675 1908 676 1912
rect 670 1907 676 1908
rect 726 1912 732 1913
rect 726 1908 727 1912
rect 731 1908 732 1912
rect 726 1907 732 1908
rect 782 1912 788 1913
rect 782 1908 783 1912
rect 787 1908 788 1912
rect 782 1907 788 1908
rect 846 1912 852 1913
rect 846 1908 847 1912
rect 851 1908 852 1912
rect 846 1907 852 1908
rect 1158 1912 1164 1913
rect 1158 1908 1159 1912
rect 1163 1908 1164 1912
rect 1158 1907 1164 1908
rect 1222 1912 1228 1913
rect 1222 1908 1223 1912
rect 1227 1908 1228 1912
rect 1222 1907 1228 1908
rect 1302 1912 1308 1913
rect 1302 1908 1303 1912
rect 1307 1908 1308 1912
rect 1302 1907 1308 1908
rect 1382 1912 1388 1913
rect 1382 1908 1383 1912
rect 1387 1908 1388 1912
rect 1382 1907 1388 1908
rect 1462 1912 1468 1913
rect 1462 1908 1463 1912
rect 1467 1908 1468 1912
rect 1462 1907 1468 1908
rect 1534 1912 1540 1913
rect 1534 1908 1535 1912
rect 1539 1908 1540 1912
rect 1534 1907 1540 1908
rect 1614 1912 1620 1913
rect 1614 1908 1615 1912
rect 1619 1908 1620 1912
rect 1614 1907 1620 1908
rect 1694 1912 1700 1913
rect 1694 1908 1695 1912
rect 1699 1908 1700 1912
rect 1694 1907 1700 1908
rect 1782 1912 1788 1913
rect 1782 1908 1783 1912
rect 1787 1908 1788 1912
rect 1782 1907 1788 1908
rect 1878 1912 1884 1913
rect 1878 1908 1879 1912
rect 1883 1908 1884 1912
rect 1878 1907 1884 1908
rect 1982 1912 1988 1913
rect 1982 1908 1983 1912
rect 1987 1908 1988 1912
rect 1982 1907 1988 1908
rect 2070 1912 2076 1913
rect 2070 1908 2071 1912
rect 2075 1908 2076 1912
rect 2070 1907 2076 1908
rect 110 1904 116 1905
rect 110 1900 111 1904
rect 115 1900 116 1904
rect 110 1899 116 1900
rect 1094 1904 1100 1905
rect 1094 1900 1095 1904
rect 1099 1900 1100 1904
rect 1094 1899 1100 1900
rect 110 1887 116 1888
rect 110 1883 111 1887
rect 115 1883 116 1887
rect 1094 1887 1100 1888
rect 110 1882 116 1883
rect 134 1884 140 1885
rect 134 1880 135 1884
rect 139 1880 140 1884
rect 134 1879 140 1880
rect 174 1884 180 1885
rect 174 1880 175 1884
rect 179 1880 180 1884
rect 174 1879 180 1880
rect 230 1884 236 1885
rect 230 1880 231 1884
rect 235 1880 236 1884
rect 230 1879 236 1880
rect 294 1884 300 1885
rect 294 1880 295 1884
rect 299 1880 300 1884
rect 294 1879 300 1880
rect 366 1884 372 1885
rect 366 1880 367 1884
rect 371 1880 372 1884
rect 366 1879 372 1880
rect 430 1884 436 1885
rect 430 1880 431 1884
rect 435 1880 436 1884
rect 430 1879 436 1880
rect 494 1884 500 1885
rect 494 1880 495 1884
rect 499 1880 500 1884
rect 494 1879 500 1880
rect 558 1884 564 1885
rect 558 1880 559 1884
rect 563 1880 564 1884
rect 558 1879 564 1880
rect 614 1884 620 1885
rect 614 1880 615 1884
rect 619 1880 620 1884
rect 614 1879 620 1880
rect 670 1884 676 1885
rect 670 1880 671 1884
rect 675 1880 676 1884
rect 670 1879 676 1880
rect 726 1884 732 1885
rect 726 1880 727 1884
rect 731 1880 732 1884
rect 726 1879 732 1880
rect 782 1884 788 1885
rect 782 1880 783 1884
rect 787 1880 788 1884
rect 782 1879 788 1880
rect 846 1884 852 1885
rect 846 1880 847 1884
rect 851 1880 852 1884
rect 1094 1883 1095 1887
rect 1099 1883 1100 1887
rect 1094 1882 1100 1883
rect 846 1879 852 1880
rect 1158 1872 1164 1873
rect 134 1868 140 1869
rect 110 1865 116 1866
rect 110 1861 111 1865
rect 115 1861 116 1865
rect 134 1864 135 1868
rect 139 1864 140 1868
rect 134 1863 140 1864
rect 198 1868 204 1869
rect 198 1864 199 1868
rect 203 1864 204 1868
rect 198 1863 204 1864
rect 270 1868 276 1869
rect 270 1864 271 1868
rect 275 1864 276 1868
rect 270 1863 276 1864
rect 334 1868 340 1869
rect 334 1864 335 1868
rect 339 1864 340 1868
rect 334 1863 340 1864
rect 398 1868 404 1869
rect 398 1864 399 1868
rect 403 1864 404 1868
rect 398 1863 404 1864
rect 454 1868 460 1869
rect 454 1864 455 1868
rect 459 1864 460 1868
rect 454 1863 460 1864
rect 502 1868 508 1869
rect 502 1864 503 1868
rect 507 1864 508 1868
rect 502 1863 508 1864
rect 550 1868 556 1869
rect 550 1864 551 1868
rect 555 1864 556 1868
rect 550 1863 556 1864
rect 598 1868 604 1869
rect 598 1864 599 1868
rect 603 1864 604 1868
rect 598 1863 604 1864
rect 646 1868 652 1869
rect 646 1864 647 1868
rect 651 1864 652 1868
rect 646 1863 652 1864
rect 694 1868 700 1869
rect 694 1864 695 1868
rect 699 1864 700 1868
rect 694 1863 700 1864
rect 750 1868 756 1869
rect 750 1864 751 1868
rect 755 1864 756 1868
rect 1158 1868 1159 1872
rect 1163 1868 1164 1872
rect 1158 1867 1164 1868
rect 1198 1872 1204 1873
rect 1198 1868 1199 1872
rect 1203 1868 1204 1872
rect 1198 1867 1204 1868
rect 1262 1872 1268 1873
rect 1262 1868 1263 1872
rect 1267 1868 1268 1872
rect 1262 1867 1268 1868
rect 1326 1872 1332 1873
rect 1326 1868 1327 1872
rect 1331 1868 1332 1872
rect 1326 1867 1332 1868
rect 1390 1872 1396 1873
rect 1390 1868 1391 1872
rect 1395 1868 1396 1872
rect 1390 1867 1396 1868
rect 1446 1872 1452 1873
rect 1446 1868 1447 1872
rect 1451 1868 1452 1872
rect 1446 1867 1452 1868
rect 1502 1872 1508 1873
rect 1502 1868 1503 1872
rect 1507 1868 1508 1872
rect 1502 1867 1508 1868
rect 1558 1872 1564 1873
rect 1558 1868 1559 1872
rect 1563 1868 1564 1872
rect 1558 1867 1564 1868
rect 1630 1872 1636 1873
rect 1630 1868 1631 1872
rect 1635 1868 1636 1872
rect 1630 1867 1636 1868
rect 1710 1872 1716 1873
rect 1710 1868 1711 1872
rect 1715 1868 1716 1872
rect 1710 1867 1716 1868
rect 1798 1872 1804 1873
rect 1798 1868 1799 1872
rect 1803 1868 1804 1872
rect 1798 1867 1804 1868
rect 1894 1872 1900 1873
rect 1894 1868 1895 1872
rect 1899 1868 1900 1872
rect 1894 1867 1900 1868
rect 1990 1872 1996 1873
rect 1990 1868 1991 1872
rect 1995 1868 1996 1872
rect 1990 1867 1996 1868
rect 2070 1872 2076 1873
rect 2070 1868 2071 1872
rect 2075 1868 2076 1872
rect 2070 1867 2076 1868
rect 750 1863 756 1864
rect 1094 1865 1100 1866
rect 110 1860 116 1861
rect 1094 1861 1095 1865
rect 1099 1861 1100 1865
rect 1094 1860 1100 1861
rect 1134 1864 1140 1865
rect 1134 1860 1135 1864
rect 1139 1860 1140 1864
rect 1134 1859 1140 1860
rect 2118 1864 2124 1865
rect 2118 1860 2119 1864
rect 2123 1860 2124 1864
rect 2118 1859 2124 1860
rect 110 1848 116 1849
rect 110 1844 111 1848
rect 115 1844 116 1848
rect 110 1843 116 1844
rect 1094 1848 1100 1849
rect 1094 1844 1095 1848
rect 1099 1844 1100 1848
rect 1094 1843 1100 1844
rect 1134 1847 1140 1848
rect 1134 1843 1135 1847
rect 1139 1843 1140 1847
rect 2118 1847 2124 1848
rect 1134 1842 1140 1843
rect 1158 1844 1164 1845
rect 134 1840 140 1841
rect 134 1836 135 1840
rect 139 1836 140 1840
rect 134 1835 140 1836
rect 198 1840 204 1841
rect 198 1836 199 1840
rect 203 1836 204 1840
rect 198 1835 204 1836
rect 270 1840 276 1841
rect 270 1836 271 1840
rect 275 1836 276 1840
rect 270 1835 276 1836
rect 334 1840 340 1841
rect 334 1836 335 1840
rect 339 1836 340 1840
rect 334 1835 340 1836
rect 398 1840 404 1841
rect 398 1836 399 1840
rect 403 1836 404 1840
rect 398 1835 404 1836
rect 454 1840 460 1841
rect 454 1836 455 1840
rect 459 1836 460 1840
rect 454 1835 460 1836
rect 502 1840 508 1841
rect 502 1836 503 1840
rect 507 1836 508 1840
rect 502 1835 508 1836
rect 550 1840 556 1841
rect 550 1836 551 1840
rect 555 1836 556 1840
rect 550 1835 556 1836
rect 598 1840 604 1841
rect 598 1836 599 1840
rect 603 1836 604 1840
rect 598 1835 604 1836
rect 646 1840 652 1841
rect 646 1836 647 1840
rect 651 1836 652 1840
rect 646 1835 652 1836
rect 694 1840 700 1841
rect 694 1836 695 1840
rect 699 1836 700 1840
rect 694 1835 700 1836
rect 750 1840 756 1841
rect 750 1836 751 1840
rect 755 1836 756 1840
rect 1158 1840 1159 1844
rect 1163 1840 1164 1844
rect 1158 1839 1164 1840
rect 1198 1844 1204 1845
rect 1198 1840 1199 1844
rect 1203 1840 1204 1844
rect 1198 1839 1204 1840
rect 1262 1844 1268 1845
rect 1262 1840 1263 1844
rect 1267 1840 1268 1844
rect 1262 1839 1268 1840
rect 1326 1844 1332 1845
rect 1326 1840 1327 1844
rect 1331 1840 1332 1844
rect 1326 1839 1332 1840
rect 1390 1844 1396 1845
rect 1390 1840 1391 1844
rect 1395 1840 1396 1844
rect 1390 1839 1396 1840
rect 1446 1844 1452 1845
rect 1446 1840 1447 1844
rect 1451 1840 1452 1844
rect 1446 1839 1452 1840
rect 1502 1844 1508 1845
rect 1502 1840 1503 1844
rect 1507 1840 1508 1844
rect 1502 1839 1508 1840
rect 1558 1844 1564 1845
rect 1558 1840 1559 1844
rect 1563 1840 1564 1844
rect 1558 1839 1564 1840
rect 1630 1844 1636 1845
rect 1630 1840 1631 1844
rect 1635 1840 1636 1844
rect 1630 1839 1636 1840
rect 1710 1844 1716 1845
rect 1710 1840 1711 1844
rect 1715 1840 1716 1844
rect 1710 1839 1716 1840
rect 1798 1844 1804 1845
rect 1798 1840 1799 1844
rect 1803 1840 1804 1844
rect 1798 1839 1804 1840
rect 1894 1844 1900 1845
rect 1894 1840 1895 1844
rect 1899 1840 1900 1844
rect 1894 1839 1900 1840
rect 1990 1844 1996 1845
rect 1990 1840 1991 1844
rect 1995 1840 1996 1844
rect 1990 1839 1996 1840
rect 2070 1844 2076 1845
rect 2070 1840 2071 1844
rect 2075 1840 2076 1844
rect 2118 1843 2119 1847
rect 2123 1843 2124 1847
rect 2118 1842 2124 1843
rect 2070 1839 2076 1840
rect 750 1835 756 1836
rect 1158 1832 1164 1833
rect 1134 1829 1140 1830
rect 1134 1825 1135 1829
rect 1139 1825 1140 1829
rect 1158 1828 1159 1832
rect 1163 1828 1164 1832
rect 1158 1827 1164 1828
rect 1230 1832 1236 1833
rect 1230 1828 1231 1832
rect 1235 1828 1236 1832
rect 1230 1827 1236 1828
rect 1302 1832 1308 1833
rect 1302 1828 1303 1832
rect 1307 1828 1308 1832
rect 1302 1827 1308 1828
rect 1382 1832 1388 1833
rect 1382 1828 1383 1832
rect 1387 1828 1388 1832
rect 1382 1827 1388 1828
rect 1462 1832 1468 1833
rect 1462 1828 1463 1832
rect 1467 1828 1468 1832
rect 1462 1827 1468 1828
rect 1550 1832 1556 1833
rect 1550 1828 1551 1832
rect 1555 1828 1556 1832
rect 1550 1827 1556 1828
rect 1646 1832 1652 1833
rect 1646 1828 1647 1832
rect 1651 1828 1652 1832
rect 1646 1827 1652 1828
rect 1750 1832 1756 1833
rect 1750 1828 1751 1832
rect 1755 1828 1756 1832
rect 1750 1827 1756 1828
rect 1854 1832 1860 1833
rect 1854 1828 1855 1832
rect 1859 1828 1860 1832
rect 1854 1827 1860 1828
rect 1966 1832 1972 1833
rect 1966 1828 1967 1832
rect 1971 1828 1972 1832
rect 1966 1827 1972 1828
rect 2070 1832 2076 1833
rect 2070 1828 2071 1832
rect 2075 1828 2076 1832
rect 2070 1827 2076 1828
rect 2118 1829 2124 1830
rect 1134 1824 1140 1825
rect 2118 1825 2119 1829
rect 2123 1825 2124 1829
rect 2118 1824 2124 1825
rect 1134 1812 1140 1813
rect 1134 1808 1135 1812
rect 1139 1808 1140 1812
rect 1134 1807 1140 1808
rect 2118 1812 2124 1813
rect 2118 1808 2119 1812
rect 2123 1808 2124 1812
rect 2118 1807 2124 1808
rect 1158 1804 1164 1805
rect 1158 1800 1159 1804
rect 1163 1800 1164 1804
rect 1158 1799 1164 1800
rect 1230 1804 1236 1805
rect 1230 1800 1231 1804
rect 1235 1800 1236 1804
rect 1230 1799 1236 1800
rect 1302 1804 1308 1805
rect 1302 1800 1303 1804
rect 1307 1800 1308 1804
rect 1302 1799 1308 1800
rect 1382 1804 1388 1805
rect 1382 1800 1383 1804
rect 1387 1800 1388 1804
rect 1382 1799 1388 1800
rect 1462 1804 1468 1805
rect 1462 1800 1463 1804
rect 1467 1800 1468 1804
rect 1462 1799 1468 1800
rect 1550 1804 1556 1805
rect 1550 1800 1551 1804
rect 1555 1800 1556 1804
rect 1550 1799 1556 1800
rect 1646 1804 1652 1805
rect 1646 1800 1647 1804
rect 1651 1800 1652 1804
rect 1646 1799 1652 1800
rect 1750 1804 1756 1805
rect 1750 1800 1751 1804
rect 1755 1800 1756 1804
rect 1750 1799 1756 1800
rect 1854 1804 1860 1805
rect 1854 1800 1855 1804
rect 1859 1800 1860 1804
rect 1854 1799 1860 1800
rect 1966 1804 1972 1805
rect 1966 1800 1967 1804
rect 1971 1800 1972 1804
rect 1966 1799 1972 1800
rect 2070 1804 2076 1805
rect 2070 1800 2071 1804
rect 2075 1800 2076 1804
rect 2070 1799 2076 1800
rect 150 1796 156 1797
rect 150 1792 151 1796
rect 155 1792 156 1796
rect 150 1791 156 1792
rect 214 1796 220 1797
rect 214 1792 215 1796
rect 219 1792 220 1796
rect 214 1791 220 1792
rect 270 1796 276 1797
rect 270 1792 271 1796
rect 275 1792 276 1796
rect 270 1791 276 1792
rect 326 1796 332 1797
rect 326 1792 327 1796
rect 331 1792 332 1796
rect 326 1791 332 1792
rect 382 1796 388 1797
rect 382 1792 383 1796
rect 387 1792 388 1796
rect 382 1791 388 1792
rect 430 1796 436 1797
rect 430 1792 431 1796
rect 435 1792 436 1796
rect 430 1791 436 1792
rect 478 1796 484 1797
rect 478 1792 479 1796
rect 483 1792 484 1796
rect 478 1791 484 1792
rect 526 1796 532 1797
rect 526 1792 527 1796
rect 531 1792 532 1796
rect 526 1791 532 1792
rect 574 1796 580 1797
rect 574 1792 575 1796
rect 579 1792 580 1796
rect 574 1791 580 1792
rect 622 1796 628 1797
rect 622 1792 623 1796
rect 627 1792 628 1796
rect 622 1791 628 1792
rect 670 1796 676 1797
rect 670 1792 671 1796
rect 675 1792 676 1796
rect 670 1791 676 1792
rect 726 1796 732 1797
rect 726 1792 727 1796
rect 731 1792 732 1796
rect 726 1791 732 1792
rect 110 1788 116 1789
rect 110 1784 111 1788
rect 115 1784 116 1788
rect 110 1783 116 1784
rect 1094 1788 1100 1789
rect 1094 1784 1095 1788
rect 1099 1784 1100 1788
rect 1094 1783 1100 1784
rect 110 1771 116 1772
rect 110 1767 111 1771
rect 115 1767 116 1771
rect 1094 1771 1100 1772
rect 110 1766 116 1767
rect 150 1768 156 1769
rect 150 1764 151 1768
rect 155 1764 156 1768
rect 150 1763 156 1764
rect 214 1768 220 1769
rect 214 1764 215 1768
rect 219 1764 220 1768
rect 214 1763 220 1764
rect 270 1768 276 1769
rect 270 1764 271 1768
rect 275 1764 276 1768
rect 270 1763 276 1764
rect 326 1768 332 1769
rect 326 1764 327 1768
rect 331 1764 332 1768
rect 326 1763 332 1764
rect 382 1768 388 1769
rect 382 1764 383 1768
rect 387 1764 388 1768
rect 382 1763 388 1764
rect 430 1768 436 1769
rect 430 1764 431 1768
rect 435 1764 436 1768
rect 430 1763 436 1764
rect 478 1768 484 1769
rect 478 1764 479 1768
rect 483 1764 484 1768
rect 478 1763 484 1764
rect 526 1768 532 1769
rect 526 1764 527 1768
rect 531 1764 532 1768
rect 526 1763 532 1764
rect 574 1768 580 1769
rect 574 1764 575 1768
rect 579 1764 580 1768
rect 574 1763 580 1764
rect 622 1768 628 1769
rect 622 1764 623 1768
rect 627 1764 628 1768
rect 622 1763 628 1764
rect 670 1768 676 1769
rect 670 1764 671 1768
rect 675 1764 676 1768
rect 670 1763 676 1764
rect 726 1768 732 1769
rect 726 1764 727 1768
rect 731 1764 732 1768
rect 1094 1767 1095 1771
rect 1099 1767 1100 1771
rect 1094 1766 1100 1767
rect 1190 1768 1196 1769
rect 726 1763 732 1764
rect 1190 1764 1191 1768
rect 1195 1764 1196 1768
rect 1190 1763 1196 1764
rect 1254 1768 1260 1769
rect 1254 1764 1255 1768
rect 1259 1764 1260 1768
rect 1254 1763 1260 1764
rect 1318 1768 1324 1769
rect 1318 1764 1319 1768
rect 1323 1764 1324 1768
rect 1318 1763 1324 1764
rect 1382 1768 1388 1769
rect 1382 1764 1383 1768
rect 1387 1764 1388 1768
rect 1382 1763 1388 1764
rect 1454 1768 1460 1769
rect 1454 1764 1455 1768
rect 1459 1764 1460 1768
rect 1454 1763 1460 1764
rect 1526 1768 1532 1769
rect 1526 1764 1527 1768
rect 1531 1764 1532 1768
rect 1526 1763 1532 1764
rect 1606 1768 1612 1769
rect 1606 1764 1607 1768
rect 1611 1764 1612 1768
rect 1606 1763 1612 1764
rect 1686 1768 1692 1769
rect 1686 1764 1687 1768
rect 1691 1764 1692 1768
rect 1686 1763 1692 1764
rect 1766 1768 1772 1769
rect 1766 1764 1767 1768
rect 1771 1764 1772 1768
rect 1766 1763 1772 1764
rect 1846 1768 1852 1769
rect 1846 1764 1847 1768
rect 1851 1764 1852 1768
rect 1846 1763 1852 1764
rect 1926 1768 1932 1769
rect 1926 1764 1927 1768
rect 1931 1764 1932 1768
rect 1926 1763 1932 1764
rect 2006 1768 2012 1769
rect 2006 1764 2007 1768
rect 2011 1764 2012 1768
rect 2006 1763 2012 1764
rect 2070 1768 2076 1769
rect 2070 1764 2071 1768
rect 2075 1764 2076 1768
rect 2070 1763 2076 1764
rect 1134 1760 1140 1761
rect 230 1756 236 1757
rect 110 1753 116 1754
rect 110 1749 111 1753
rect 115 1749 116 1753
rect 230 1752 231 1756
rect 235 1752 236 1756
rect 230 1751 236 1752
rect 294 1756 300 1757
rect 294 1752 295 1756
rect 299 1752 300 1756
rect 294 1751 300 1752
rect 350 1756 356 1757
rect 350 1752 351 1756
rect 355 1752 356 1756
rect 350 1751 356 1752
rect 414 1756 420 1757
rect 414 1752 415 1756
rect 419 1752 420 1756
rect 414 1751 420 1752
rect 478 1756 484 1757
rect 478 1752 479 1756
rect 483 1752 484 1756
rect 478 1751 484 1752
rect 542 1756 548 1757
rect 542 1752 543 1756
rect 547 1752 548 1756
rect 542 1751 548 1752
rect 614 1756 620 1757
rect 614 1752 615 1756
rect 619 1752 620 1756
rect 614 1751 620 1752
rect 686 1756 692 1757
rect 686 1752 687 1756
rect 691 1752 692 1756
rect 686 1751 692 1752
rect 758 1756 764 1757
rect 758 1752 759 1756
rect 763 1752 764 1756
rect 758 1751 764 1752
rect 830 1756 836 1757
rect 830 1752 831 1756
rect 835 1752 836 1756
rect 830 1751 836 1752
rect 910 1756 916 1757
rect 910 1752 911 1756
rect 915 1752 916 1756
rect 910 1751 916 1752
rect 990 1756 996 1757
rect 990 1752 991 1756
rect 995 1752 996 1756
rect 1134 1756 1135 1760
rect 1139 1756 1140 1760
rect 1134 1755 1140 1756
rect 2118 1760 2124 1761
rect 2118 1756 2119 1760
rect 2123 1756 2124 1760
rect 2118 1755 2124 1756
rect 990 1751 996 1752
rect 1094 1753 1100 1754
rect 110 1748 116 1749
rect 1094 1749 1095 1753
rect 1099 1749 1100 1753
rect 1094 1748 1100 1749
rect 1134 1743 1140 1744
rect 1134 1739 1135 1743
rect 1139 1739 1140 1743
rect 2118 1743 2124 1744
rect 1134 1738 1140 1739
rect 1190 1740 1196 1741
rect 110 1736 116 1737
rect 110 1732 111 1736
rect 115 1732 116 1736
rect 110 1731 116 1732
rect 1094 1736 1100 1737
rect 1094 1732 1095 1736
rect 1099 1732 1100 1736
rect 1190 1736 1191 1740
rect 1195 1736 1196 1740
rect 1190 1735 1196 1736
rect 1254 1740 1260 1741
rect 1254 1736 1255 1740
rect 1259 1736 1260 1740
rect 1254 1735 1260 1736
rect 1318 1740 1324 1741
rect 1318 1736 1319 1740
rect 1323 1736 1324 1740
rect 1318 1735 1324 1736
rect 1382 1740 1388 1741
rect 1382 1736 1383 1740
rect 1387 1736 1388 1740
rect 1382 1735 1388 1736
rect 1454 1740 1460 1741
rect 1454 1736 1455 1740
rect 1459 1736 1460 1740
rect 1454 1735 1460 1736
rect 1526 1740 1532 1741
rect 1526 1736 1527 1740
rect 1531 1736 1532 1740
rect 1526 1735 1532 1736
rect 1606 1740 1612 1741
rect 1606 1736 1607 1740
rect 1611 1736 1612 1740
rect 1606 1735 1612 1736
rect 1686 1740 1692 1741
rect 1686 1736 1687 1740
rect 1691 1736 1692 1740
rect 1686 1735 1692 1736
rect 1766 1740 1772 1741
rect 1766 1736 1767 1740
rect 1771 1736 1772 1740
rect 1766 1735 1772 1736
rect 1846 1740 1852 1741
rect 1846 1736 1847 1740
rect 1851 1736 1852 1740
rect 1846 1735 1852 1736
rect 1926 1740 1932 1741
rect 1926 1736 1927 1740
rect 1931 1736 1932 1740
rect 1926 1735 1932 1736
rect 2006 1740 2012 1741
rect 2006 1736 2007 1740
rect 2011 1736 2012 1740
rect 2006 1735 2012 1736
rect 2070 1740 2076 1741
rect 2070 1736 2071 1740
rect 2075 1736 2076 1740
rect 2118 1739 2119 1743
rect 2123 1739 2124 1743
rect 2118 1738 2124 1739
rect 2070 1735 2076 1736
rect 1094 1731 1100 1732
rect 230 1728 236 1729
rect 230 1724 231 1728
rect 235 1724 236 1728
rect 230 1723 236 1724
rect 294 1728 300 1729
rect 294 1724 295 1728
rect 299 1724 300 1728
rect 294 1723 300 1724
rect 350 1728 356 1729
rect 350 1724 351 1728
rect 355 1724 356 1728
rect 350 1723 356 1724
rect 414 1728 420 1729
rect 414 1724 415 1728
rect 419 1724 420 1728
rect 414 1723 420 1724
rect 478 1728 484 1729
rect 478 1724 479 1728
rect 483 1724 484 1728
rect 478 1723 484 1724
rect 542 1728 548 1729
rect 542 1724 543 1728
rect 547 1724 548 1728
rect 542 1723 548 1724
rect 614 1728 620 1729
rect 614 1724 615 1728
rect 619 1724 620 1728
rect 614 1723 620 1724
rect 686 1728 692 1729
rect 686 1724 687 1728
rect 691 1724 692 1728
rect 686 1723 692 1724
rect 758 1728 764 1729
rect 758 1724 759 1728
rect 763 1724 764 1728
rect 758 1723 764 1724
rect 830 1728 836 1729
rect 830 1724 831 1728
rect 835 1724 836 1728
rect 830 1723 836 1724
rect 910 1728 916 1729
rect 910 1724 911 1728
rect 915 1724 916 1728
rect 910 1723 916 1724
rect 990 1728 996 1729
rect 990 1724 991 1728
rect 995 1724 996 1728
rect 1246 1728 1252 1729
rect 990 1723 996 1724
rect 1134 1725 1140 1726
rect 1134 1721 1135 1725
rect 1139 1721 1140 1725
rect 1246 1724 1247 1728
rect 1251 1724 1252 1728
rect 1246 1723 1252 1724
rect 1294 1728 1300 1729
rect 1294 1724 1295 1728
rect 1299 1724 1300 1728
rect 1294 1723 1300 1724
rect 1342 1728 1348 1729
rect 1342 1724 1343 1728
rect 1347 1724 1348 1728
rect 1342 1723 1348 1724
rect 1398 1728 1404 1729
rect 1398 1724 1399 1728
rect 1403 1724 1404 1728
rect 1398 1723 1404 1724
rect 1462 1728 1468 1729
rect 1462 1724 1463 1728
rect 1467 1724 1468 1728
rect 1462 1723 1468 1724
rect 1526 1728 1532 1729
rect 1526 1724 1527 1728
rect 1531 1724 1532 1728
rect 1526 1723 1532 1724
rect 1598 1728 1604 1729
rect 1598 1724 1599 1728
rect 1603 1724 1604 1728
rect 1598 1723 1604 1724
rect 1670 1728 1676 1729
rect 1670 1724 1671 1728
rect 1675 1724 1676 1728
rect 1670 1723 1676 1724
rect 1742 1728 1748 1729
rect 1742 1724 1743 1728
rect 1747 1724 1748 1728
rect 1742 1723 1748 1724
rect 1806 1728 1812 1729
rect 1806 1724 1807 1728
rect 1811 1724 1812 1728
rect 1806 1723 1812 1724
rect 1878 1728 1884 1729
rect 1878 1724 1879 1728
rect 1883 1724 1884 1728
rect 1878 1723 1884 1724
rect 1950 1728 1956 1729
rect 1950 1724 1951 1728
rect 1955 1724 1956 1728
rect 1950 1723 1956 1724
rect 2022 1728 2028 1729
rect 2022 1724 2023 1728
rect 2027 1724 2028 1728
rect 2022 1723 2028 1724
rect 2070 1728 2076 1729
rect 2070 1724 2071 1728
rect 2075 1724 2076 1728
rect 2070 1723 2076 1724
rect 2118 1725 2124 1726
rect 1134 1720 1140 1721
rect 2118 1721 2119 1725
rect 2123 1721 2124 1725
rect 2118 1720 2124 1721
rect 1134 1708 1140 1709
rect 1134 1704 1135 1708
rect 1139 1704 1140 1708
rect 1134 1703 1140 1704
rect 2118 1708 2124 1709
rect 2118 1704 2119 1708
rect 2123 1704 2124 1708
rect 2118 1703 2124 1704
rect 1246 1700 1252 1701
rect 1246 1696 1247 1700
rect 1251 1696 1252 1700
rect 1246 1695 1252 1696
rect 1294 1700 1300 1701
rect 1294 1696 1295 1700
rect 1299 1696 1300 1700
rect 1294 1695 1300 1696
rect 1342 1700 1348 1701
rect 1342 1696 1343 1700
rect 1347 1696 1348 1700
rect 1342 1695 1348 1696
rect 1398 1700 1404 1701
rect 1398 1696 1399 1700
rect 1403 1696 1404 1700
rect 1398 1695 1404 1696
rect 1462 1700 1468 1701
rect 1462 1696 1463 1700
rect 1467 1696 1468 1700
rect 1462 1695 1468 1696
rect 1526 1700 1532 1701
rect 1526 1696 1527 1700
rect 1531 1696 1532 1700
rect 1526 1695 1532 1696
rect 1598 1700 1604 1701
rect 1598 1696 1599 1700
rect 1603 1696 1604 1700
rect 1598 1695 1604 1696
rect 1670 1700 1676 1701
rect 1670 1696 1671 1700
rect 1675 1696 1676 1700
rect 1670 1695 1676 1696
rect 1742 1700 1748 1701
rect 1742 1696 1743 1700
rect 1747 1696 1748 1700
rect 1742 1695 1748 1696
rect 1806 1700 1812 1701
rect 1806 1696 1807 1700
rect 1811 1696 1812 1700
rect 1806 1695 1812 1696
rect 1878 1700 1884 1701
rect 1878 1696 1879 1700
rect 1883 1696 1884 1700
rect 1878 1695 1884 1696
rect 1950 1700 1956 1701
rect 1950 1696 1951 1700
rect 1955 1696 1956 1700
rect 1950 1695 1956 1696
rect 2022 1700 2028 1701
rect 2022 1696 2023 1700
rect 2027 1696 2028 1700
rect 2022 1695 2028 1696
rect 2070 1700 2076 1701
rect 2070 1696 2071 1700
rect 2075 1696 2076 1700
rect 2070 1695 2076 1696
rect 134 1688 140 1689
rect 134 1684 135 1688
rect 139 1684 140 1688
rect 134 1683 140 1684
rect 198 1688 204 1689
rect 198 1684 199 1688
rect 203 1684 204 1688
rect 198 1683 204 1684
rect 278 1688 284 1689
rect 278 1684 279 1688
rect 283 1684 284 1688
rect 278 1683 284 1684
rect 366 1688 372 1689
rect 366 1684 367 1688
rect 371 1684 372 1688
rect 366 1683 372 1684
rect 462 1688 468 1689
rect 462 1684 463 1688
rect 467 1684 468 1688
rect 462 1683 468 1684
rect 550 1688 556 1689
rect 550 1684 551 1688
rect 555 1684 556 1688
rect 550 1683 556 1684
rect 638 1688 644 1689
rect 638 1684 639 1688
rect 643 1684 644 1688
rect 638 1683 644 1684
rect 718 1688 724 1689
rect 718 1684 719 1688
rect 723 1684 724 1688
rect 718 1683 724 1684
rect 790 1688 796 1689
rect 790 1684 791 1688
rect 795 1684 796 1688
rect 790 1683 796 1684
rect 854 1688 860 1689
rect 854 1684 855 1688
rect 859 1684 860 1688
rect 854 1683 860 1684
rect 918 1688 924 1689
rect 918 1684 919 1688
rect 923 1684 924 1688
rect 918 1683 924 1684
rect 982 1688 988 1689
rect 982 1684 983 1688
rect 987 1684 988 1688
rect 982 1683 988 1684
rect 1046 1688 1052 1689
rect 1046 1684 1047 1688
rect 1051 1684 1052 1688
rect 1046 1683 1052 1684
rect 110 1680 116 1681
rect 110 1676 111 1680
rect 115 1676 116 1680
rect 110 1675 116 1676
rect 1094 1680 1100 1681
rect 1094 1676 1095 1680
rect 1099 1676 1100 1680
rect 1094 1675 1100 1676
rect 110 1663 116 1664
rect 110 1659 111 1663
rect 115 1659 116 1663
rect 1094 1663 1100 1664
rect 110 1658 116 1659
rect 134 1660 140 1661
rect 134 1656 135 1660
rect 139 1656 140 1660
rect 134 1655 140 1656
rect 198 1660 204 1661
rect 198 1656 199 1660
rect 203 1656 204 1660
rect 198 1655 204 1656
rect 278 1660 284 1661
rect 278 1656 279 1660
rect 283 1656 284 1660
rect 278 1655 284 1656
rect 366 1660 372 1661
rect 366 1656 367 1660
rect 371 1656 372 1660
rect 366 1655 372 1656
rect 462 1660 468 1661
rect 462 1656 463 1660
rect 467 1656 468 1660
rect 462 1655 468 1656
rect 550 1660 556 1661
rect 550 1656 551 1660
rect 555 1656 556 1660
rect 550 1655 556 1656
rect 638 1660 644 1661
rect 638 1656 639 1660
rect 643 1656 644 1660
rect 638 1655 644 1656
rect 718 1660 724 1661
rect 718 1656 719 1660
rect 723 1656 724 1660
rect 718 1655 724 1656
rect 790 1660 796 1661
rect 790 1656 791 1660
rect 795 1656 796 1660
rect 790 1655 796 1656
rect 854 1660 860 1661
rect 854 1656 855 1660
rect 859 1656 860 1660
rect 854 1655 860 1656
rect 918 1660 924 1661
rect 918 1656 919 1660
rect 923 1656 924 1660
rect 918 1655 924 1656
rect 982 1660 988 1661
rect 982 1656 983 1660
rect 987 1656 988 1660
rect 982 1655 988 1656
rect 1046 1660 1052 1661
rect 1046 1656 1047 1660
rect 1051 1656 1052 1660
rect 1094 1659 1095 1663
rect 1099 1659 1100 1663
rect 1094 1658 1100 1659
rect 1262 1660 1268 1661
rect 1046 1655 1052 1656
rect 1262 1656 1263 1660
rect 1267 1656 1268 1660
rect 1262 1655 1268 1656
rect 1302 1660 1308 1661
rect 1302 1656 1303 1660
rect 1307 1656 1308 1660
rect 1302 1655 1308 1656
rect 1342 1660 1348 1661
rect 1342 1656 1343 1660
rect 1347 1656 1348 1660
rect 1342 1655 1348 1656
rect 1390 1660 1396 1661
rect 1390 1656 1391 1660
rect 1395 1656 1396 1660
rect 1390 1655 1396 1656
rect 1446 1660 1452 1661
rect 1446 1656 1447 1660
rect 1451 1656 1452 1660
rect 1446 1655 1452 1656
rect 1502 1660 1508 1661
rect 1502 1656 1503 1660
rect 1507 1656 1508 1660
rect 1502 1655 1508 1656
rect 1566 1660 1572 1661
rect 1566 1656 1567 1660
rect 1571 1656 1572 1660
rect 1566 1655 1572 1656
rect 1630 1660 1636 1661
rect 1630 1656 1631 1660
rect 1635 1656 1636 1660
rect 1630 1655 1636 1656
rect 1694 1660 1700 1661
rect 1694 1656 1695 1660
rect 1699 1656 1700 1660
rect 1694 1655 1700 1656
rect 1758 1660 1764 1661
rect 1758 1656 1759 1660
rect 1763 1656 1764 1660
rect 1758 1655 1764 1656
rect 1830 1660 1836 1661
rect 1830 1656 1831 1660
rect 1835 1656 1836 1660
rect 1830 1655 1836 1656
rect 1910 1660 1916 1661
rect 1910 1656 1911 1660
rect 1915 1656 1916 1660
rect 1910 1655 1916 1656
rect 1998 1660 2004 1661
rect 1998 1656 1999 1660
rect 2003 1656 2004 1660
rect 1998 1655 2004 1656
rect 2070 1660 2076 1661
rect 2070 1656 2071 1660
rect 2075 1656 2076 1660
rect 2070 1655 2076 1656
rect 1134 1652 1140 1653
rect 1134 1648 1135 1652
rect 1139 1648 1140 1652
rect 1134 1647 1140 1648
rect 2118 1652 2124 1653
rect 2118 1648 2119 1652
rect 2123 1648 2124 1652
rect 2118 1647 2124 1648
rect 134 1644 140 1645
rect 110 1641 116 1642
rect 110 1637 111 1641
rect 115 1637 116 1641
rect 134 1640 135 1644
rect 139 1640 140 1644
rect 134 1639 140 1640
rect 182 1644 188 1645
rect 182 1640 183 1644
rect 187 1640 188 1644
rect 182 1639 188 1640
rect 262 1644 268 1645
rect 262 1640 263 1644
rect 267 1640 268 1644
rect 262 1639 268 1640
rect 342 1644 348 1645
rect 342 1640 343 1644
rect 347 1640 348 1644
rect 342 1639 348 1640
rect 422 1644 428 1645
rect 422 1640 423 1644
rect 427 1640 428 1644
rect 422 1639 428 1640
rect 502 1644 508 1645
rect 502 1640 503 1644
rect 507 1640 508 1644
rect 502 1639 508 1640
rect 582 1644 588 1645
rect 582 1640 583 1644
rect 587 1640 588 1644
rect 582 1639 588 1640
rect 654 1644 660 1645
rect 654 1640 655 1644
rect 659 1640 660 1644
rect 654 1639 660 1640
rect 726 1644 732 1645
rect 726 1640 727 1644
rect 731 1640 732 1644
rect 726 1639 732 1640
rect 790 1644 796 1645
rect 790 1640 791 1644
rect 795 1640 796 1644
rect 790 1639 796 1640
rect 846 1644 852 1645
rect 846 1640 847 1644
rect 851 1640 852 1644
rect 846 1639 852 1640
rect 902 1644 908 1645
rect 902 1640 903 1644
rect 907 1640 908 1644
rect 902 1639 908 1640
rect 958 1644 964 1645
rect 958 1640 959 1644
rect 963 1640 964 1644
rect 958 1639 964 1640
rect 1006 1644 1012 1645
rect 1006 1640 1007 1644
rect 1011 1640 1012 1644
rect 1006 1639 1012 1640
rect 1046 1644 1052 1645
rect 1046 1640 1047 1644
rect 1051 1640 1052 1644
rect 1046 1639 1052 1640
rect 1094 1641 1100 1642
rect 110 1636 116 1637
rect 1094 1637 1095 1641
rect 1099 1637 1100 1641
rect 1094 1636 1100 1637
rect 1134 1635 1140 1636
rect 1134 1631 1135 1635
rect 1139 1631 1140 1635
rect 2118 1635 2124 1636
rect 1134 1630 1140 1631
rect 1262 1632 1268 1633
rect 1262 1628 1263 1632
rect 1267 1628 1268 1632
rect 1262 1627 1268 1628
rect 1302 1632 1308 1633
rect 1302 1628 1303 1632
rect 1307 1628 1308 1632
rect 1302 1627 1308 1628
rect 1342 1632 1348 1633
rect 1342 1628 1343 1632
rect 1347 1628 1348 1632
rect 1342 1627 1348 1628
rect 1390 1632 1396 1633
rect 1390 1628 1391 1632
rect 1395 1628 1396 1632
rect 1390 1627 1396 1628
rect 1446 1632 1452 1633
rect 1446 1628 1447 1632
rect 1451 1628 1452 1632
rect 1446 1627 1452 1628
rect 1502 1632 1508 1633
rect 1502 1628 1503 1632
rect 1507 1628 1508 1632
rect 1502 1627 1508 1628
rect 1566 1632 1572 1633
rect 1566 1628 1567 1632
rect 1571 1628 1572 1632
rect 1566 1627 1572 1628
rect 1630 1632 1636 1633
rect 1630 1628 1631 1632
rect 1635 1628 1636 1632
rect 1630 1627 1636 1628
rect 1694 1632 1700 1633
rect 1694 1628 1695 1632
rect 1699 1628 1700 1632
rect 1694 1627 1700 1628
rect 1758 1632 1764 1633
rect 1758 1628 1759 1632
rect 1763 1628 1764 1632
rect 1758 1627 1764 1628
rect 1830 1632 1836 1633
rect 1830 1628 1831 1632
rect 1835 1628 1836 1632
rect 1830 1627 1836 1628
rect 1910 1632 1916 1633
rect 1910 1628 1911 1632
rect 1915 1628 1916 1632
rect 1910 1627 1916 1628
rect 1998 1632 2004 1633
rect 1998 1628 1999 1632
rect 2003 1628 2004 1632
rect 1998 1627 2004 1628
rect 2070 1632 2076 1633
rect 2070 1628 2071 1632
rect 2075 1628 2076 1632
rect 2118 1631 2119 1635
rect 2123 1631 2124 1635
rect 2118 1630 2124 1631
rect 2070 1627 2076 1628
rect 110 1624 116 1625
rect 110 1620 111 1624
rect 115 1620 116 1624
rect 110 1619 116 1620
rect 1094 1624 1100 1625
rect 1094 1620 1095 1624
rect 1099 1620 1100 1624
rect 1094 1619 1100 1620
rect 134 1616 140 1617
rect 134 1612 135 1616
rect 139 1612 140 1616
rect 134 1611 140 1612
rect 182 1616 188 1617
rect 182 1612 183 1616
rect 187 1612 188 1616
rect 182 1611 188 1612
rect 262 1616 268 1617
rect 262 1612 263 1616
rect 267 1612 268 1616
rect 262 1611 268 1612
rect 342 1616 348 1617
rect 342 1612 343 1616
rect 347 1612 348 1616
rect 342 1611 348 1612
rect 422 1616 428 1617
rect 422 1612 423 1616
rect 427 1612 428 1616
rect 422 1611 428 1612
rect 502 1616 508 1617
rect 502 1612 503 1616
rect 507 1612 508 1616
rect 502 1611 508 1612
rect 582 1616 588 1617
rect 582 1612 583 1616
rect 587 1612 588 1616
rect 582 1611 588 1612
rect 654 1616 660 1617
rect 654 1612 655 1616
rect 659 1612 660 1616
rect 654 1611 660 1612
rect 726 1616 732 1617
rect 726 1612 727 1616
rect 731 1612 732 1616
rect 726 1611 732 1612
rect 790 1616 796 1617
rect 790 1612 791 1616
rect 795 1612 796 1616
rect 790 1611 796 1612
rect 846 1616 852 1617
rect 846 1612 847 1616
rect 851 1612 852 1616
rect 846 1611 852 1612
rect 902 1616 908 1617
rect 902 1612 903 1616
rect 907 1612 908 1616
rect 902 1611 908 1612
rect 958 1616 964 1617
rect 958 1612 959 1616
rect 963 1612 964 1616
rect 958 1611 964 1612
rect 1006 1616 1012 1617
rect 1006 1612 1007 1616
rect 1011 1612 1012 1616
rect 1006 1611 1012 1612
rect 1046 1616 1052 1617
rect 1046 1612 1047 1616
rect 1051 1612 1052 1616
rect 1046 1611 1052 1612
rect 1158 1608 1164 1609
rect 1134 1605 1140 1606
rect 1134 1601 1135 1605
rect 1139 1601 1140 1605
rect 1158 1604 1159 1608
rect 1163 1604 1164 1608
rect 1158 1603 1164 1604
rect 1214 1608 1220 1609
rect 1214 1604 1215 1608
rect 1219 1604 1220 1608
rect 1214 1603 1220 1604
rect 1302 1608 1308 1609
rect 1302 1604 1303 1608
rect 1307 1604 1308 1608
rect 1302 1603 1308 1604
rect 1382 1608 1388 1609
rect 1382 1604 1383 1608
rect 1387 1604 1388 1608
rect 1382 1603 1388 1604
rect 1462 1608 1468 1609
rect 1462 1604 1463 1608
rect 1467 1604 1468 1608
rect 1462 1603 1468 1604
rect 1542 1608 1548 1609
rect 1542 1604 1543 1608
rect 1547 1604 1548 1608
rect 1542 1603 1548 1604
rect 1622 1608 1628 1609
rect 1622 1604 1623 1608
rect 1627 1604 1628 1608
rect 1622 1603 1628 1604
rect 1710 1608 1716 1609
rect 1710 1604 1711 1608
rect 1715 1604 1716 1608
rect 1710 1603 1716 1604
rect 1798 1608 1804 1609
rect 1798 1604 1799 1608
rect 1803 1604 1804 1608
rect 1798 1603 1804 1604
rect 1886 1608 1892 1609
rect 1886 1604 1887 1608
rect 1891 1604 1892 1608
rect 1886 1603 1892 1604
rect 1982 1608 1988 1609
rect 1982 1604 1983 1608
rect 1987 1604 1988 1608
rect 1982 1603 1988 1604
rect 2070 1608 2076 1609
rect 2070 1604 2071 1608
rect 2075 1604 2076 1608
rect 2070 1603 2076 1604
rect 2118 1605 2124 1606
rect 1134 1600 1140 1601
rect 2118 1601 2119 1605
rect 2123 1601 2124 1605
rect 2118 1600 2124 1601
rect 1134 1588 1140 1589
rect 1134 1584 1135 1588
rect 1139 1584 1140 1588
rect 1134 1583 1140 1584
rect 2118 1588 2124 1589
rect 2118 1584 2119 1588
rect 2123 1584 2124 1588
rect 2118 1583 2124 1584
rect 134 1580 140 1581
rect 134 1576 135 1580
rect 139 1576 140 1580
rect 134 1575 140 1576
rect 174 1580 180 1581
rect 174 1576 175 1580
rect 179 1576 180 1580
rect 174 1575 180 1576
rect 230 1580 236 1581
rect 230 1576 231 1580
rect 235 1576 236 1580
rect 230 1575 236 1576
rect 302 1580 308 1581
rect 302 1576 303 1580
rect 307 1576 308 1580
rect 302 1575 308 1576
rect 374 1580 380 1581
rect 374 1576 375 1580
rect 379 1576 380 1580
rect 374 1575 380 1576
rect 454 1580 460 1581
rect 454 1576 455 1580
rect 459 1576 460 1580
rect 454 1575 460 1576
rect 526 1580 532 1581
rect 526 1576 527 1580
rect 531 1576 532 1580
rect 526 1575 532 1576
rect 598 1580 604 1581
rect 598 1576 599 1580
rect 603 1576 604 1580
rect 598 1575 604 1576
rect 670 1580 676 1581
rect 670 1576 671 1580
rect 675 1576 676 1580
rect 670 1575 676 1576
rect 742 1580 748 1581
rect 742 1576 743 1580
rect 747 1576 748 1580
rect 742 1575 748 1576
rect 814 1580 820 1581
rect 814 1576 815 1580
rect 819 1576 820 1580
rect 814 1575 820 1576
rect 886 1580 892 1581
rect 886 1576 887 1580
rect 891 1576 892 1580
rect 886 1575 892 1576
rect 1158 1580 1164 1581
rect 1158 1576 1159 1580
rect 1163 1576 1164 1580
rect 1158 1575 1164 1576
rect 1214 1580 1220 1581
rect 1214 1576 1215 1580
rect 1219 1576 1220 1580
rect 1214 1575 1220 1576
rect 1302 1580 1308 1581
rect 1302 1576 1303 1580
rect 1307 1576 1308 1580
rect 1302 1575 1308 1576
rect 1382 1580 1388 1581
rect 1382 1576 1383 1580
rect 1387 1576 1388 1580
rect 1382 1575 1388 1576
rect 1462 1580 1468 1581
rect 1462 1576 1463 1580
rect 1467 1576 1468 1580
rect 1462 1575 1468 1576
rect 1542 1580 1548 1581
rect 1542 1576 1543 1580
rect 1547 1576 1548 1580
rect 1542 1575 1548 1576
rect 1622 1580 1628 1581
rect 1622 1576 1623 1580
rect 1627 1576 1628 1580
rect 1622 1575 1628 1576
rect 1710 1580 1716 1581
rect 1710 1576 1711 1580
rect 1715 1576 1716 1580
rect 1710 1575 1716 1576
rect 1798 1580 1804 1581
rect 1798 1576 1799 1580
rect 1803 1576 1804 1580
rect 1798 1575 1804 1576
rect 1886 1580 1892 1581
rect 1886 1576 1887 1580
rect 1891 1576 1892 1580
rect 1886 1575 1892 1576
rect 1982 1580 1988 1581
rect 1982 1576 1983 1580
rect 1987 1576 1988 1580
rect 1982 1575 1988 1576
rect 2070 1580 2076 1581
rect 2070 1576 2071 1580
rect 2075 1576 2076 1580
rect 2070 1575 2076 1576
rect 110 1572 116 1573
rect 110 1568 111 1572
rect 115 1568 116 1572
rect 110 1567 116 1568
rect 1094 1572 1100 1573
rect 1094 1568 1095 1572
rect 1099 1568 1100 1572
rect 1094 1567 1100 1568
rect 110 1555 116 1556
rect 110 1551 111 1555
rect 115 1551 116 1555
rect 1094 1555 1100 1556
rect 110 1550 116 1551
rect 134 1552 140 1553
rect 134 1548 135 1552
rect 139 1548 140 1552
rect 134 1547 140 1548
rect 174 1552 180 1553
rect 174 1548 175 1552
rect 179 1548 180 1552
rect 174 1547 180 1548
rect 230 1552 236 1553
rect 230 1548 231 1552
rect 235 1548 236 1552
rect 230 1547 236 1548
rect 302 1552 308 1553
rect 302 1548 303 1552
rect 307 1548 308 1552
rect 302 1547 308 1548
rect 374 1552 380 1553
rect 374 1548 375 1552
rect 379 1548 380 1552
rect 374 1547 380 1548
rect 454 1552 460 1553
rect 454 1548 455 1552
rect 459 1548 460 1552
rect 454 1547 460 1548
rect 526 1552 532 1553
rect 526 1548 527 1552
rect 531 1548 532 1552
rect 526 1547 532 1548
rect 598 1552 604 1553
rect 598 1548 599 1552
rect 603 1548 604 1552
rect 598 1547 604 1548
rect 670 1552 676 1553
rect 670 1548 671 1552
rect 675 1548 676 1552
rect 670 1547 676 1548
rect 742 1552 748 1553
rect 742 1548 743 1552
rect 747 1548 748 1552
rect 742 1547 748 1548
rect 814 1552 820 1553
rect 814 1548 815 1552
rect 819 1548 820 1552
rect 814 1547 820 1548
rect 886 1552 892 1553
rect 886 1548 887 1552
rect 891 1548 892 1552
rect 1094 1551 1095 1555
rect 1099 1551 1100 1555
rect 1094 1550 1100 1551
rect 886 1547 892 1548
rect 1158 1544 1164 1545
rect 134 1540 140 1541
rect 110 1537 116 1538
rect 110 1533 111 1537
rect 115 1533 116 1537
rect 134 1536 135 1540
rect 139 1536 140 1540
rect 134 1535 140 1536
rect 174 1540 180 1541
rect 174 1536 175 1540
rect 179 1536 180 1540
rect 174 1535 180 1536
rect 230 1540 236 1541
rect 230 1536 231 1540
rect 235 1536 236 1540
rect 230 1535 236 1536
rect 310 1540 316 1541
rect 310 1536 311 1540
rect 315 1536 316 1540
rect 310 1535 316 1536
rect 390 1540 396 1541
rect 390 1536 391 1540
rect 395 1536 396 1540
rect 390 1535 396 1536
rect 478 1540 484 1541
rect 478 1536 479 1540
rect 483 1536 484 1540
rect 478 1535 484 1536
rect 566 1540 572 1541
rect 566 1536 567 1540
rect 571 1536 572 1540
rect 566 1535 572 1536
rect 654 1540 660 1541
rect 654 1536 655 1540
rect 659 1536 660 1540
rect 654 1535 660 1536
rect 742 1540 748 1541
rect 742 1536 743 1540
rect 747 1536 748 1540
rect 742 1535 748 1536
rect 822 1540 828 1541
rect 822 1536 823 1540
rect 827 1536 828 1540
rect 822 1535 828 1536
rect 910 1540 916 1541
rect 910 1536 911 1540
rect 915 1536 916 1540
rect 910 1535 916 1536
rect 998 1540 1004 1541
rect 998 1536 999 1540
rect 1003 1536 1004 1540
rect 1158 1540 1159 1544
rect 1163 1540 1164 1544
rect 1158 1539 1164 1540
rect 1198 1544 1204 1545
rect 1198 1540 1199 1544
rect 1203 1540 1204 1544
rect 1198 1539 1204 1540
rect 1246 1544 1252 1545
rect 1246 1540 1247 1544
rect 1251 1540 1252 1544
rect 1246 1539 1252 1540
rect 1318 1544 1324 1545
rect 1318 1540 1319 1544
rect 1323 1540 1324 1544
rect 1318 1539 1324 1540
rect 1398 1544 1404 1545
rect 1398 1540 1399 1544
rect 1403 1540 1404 1544
rect 1398 1539 1404 1540
rect 1478 1544 1484 1545
rect 1478 1540 1479 1544
rect 1483 1540 1484 1544
rect 1478 1539 1484 1540
rect 1558 1544 1564 1545
rect 1558 1540 1559 1544
rect 1563 1540 1564 1544
rect 1558 1539 1564 1540
rect 1646 1544 1652 1545
rect 1646 1540 1647 1544
rect 1651 1540 1652 1544
rect 1646 1539 1652 1540
rect 1734 1544 1740 1545
rect 1734 1540 1735 1544
rect 1739 1540 1740 1544
rect 1734 1539 1740 1540
rect 1822 1544 1828 1545
rect 1822 1540 1823 1544
rect 1827 1540 1828 1544
rect 1822 1539 1828 1540
rect 1910 1544 1916 1545
rect 1910 1540 1911 1544
rect 1915 1540 1916 1544
rect 1910 1539 1916 1540
rect 1998 1544 2004 1545
rect 1998 1540 1999 1544
rect 2003 1540 2004 1544
rect 1998 1539 2004 1540
rect 2070 1544 2076 1545
rect 2070 1540 2071 1544
rect 2075 1540 2076 1544
rect 2070 1539 2076 1540
rect 998 1535 1004 1536
rect 1094 1537 1100 1538
rect 110 1532 116 1533
rect 1094 1533 1095 1537
rect 1099 1533 1100 1537
rect 1094 1532 1100 1533
rect 1134 1536 1140 1537
rect 1134 1532 1135 1536
rect 1139 1532 1140 1536
rect 1134 1531 1140 1532
rect 2118 1536 2124 1537
rect 2118 1532 2119 1536
rect 2123 1532 2124 1536
rect 2118 1531 2124 1532
rect 110 1520 116 1521
rect 110 1516 111 1520
rect 115 1516 116 1520
rect 110 1515 116 1516
rect 1094 1520 1100 1521
rect 1094 1516 1095 1520
rect 1099 1516 1100 1520
rect 1094 1515 1100 1516
rect 1134 1519 1140 1520
rect 1134 1515 1135 1519
rect 1139 1515 1140 1519
rect 2118 1519 2124 1520
rect 1134 1514 1140 1515
rect 1158 1516 1164 1517
rect 134 1512 140 1513
rect 134 1508 135 1512
rect 139 1508 140 1512
rect 134 1507 140 1508
rect 174 1512 180 1513
rect 174 1508 175 1512
rect 179 1508 180 1512
rect 174 1507 180 1508
rect 230 1512 236 1513
rect 230 1508 231 1512
rect 235 1508 236 1512
rect 230 1507 236 1508
rect 310 1512 316 1513
rect 310 1508 311 1512
rect 315 1508 316 1512
rect 310 1507 316 1508
rect 390 1512 396 1513
rect 390 1508 391 1512
rect 395 1508 396 1512
rect 390 1507 396 1508
rect 478 1512 484 1513
rect 478 1508 479 1512
rect 483 1508 484 1512
rect 478 1507 484 1508
rect 566 1512 572 1513
rect 566 1508 567 1512
rect 571 1508 572 1512
rect 566 1507 572 1508
rect 654 1512 660 1513
rect 654 1508 655 1512
rect 659 1508 660 1512
rect 654 1507 660 1508
rect 742 1512 748 1513
rect 742 1508 743 1512
rect 747 1508 748 1512
rect 742 1507 748 1508
rect 822 1512 828 1513
rect 822 1508 823 1512
rect 827 1508 828 1512
rect 822 1507 828 1508
rect 910 1512 916 1513
rect 910 1508 911 1512
rect 915 1508 916 1512
rect 910 1507 916 1508
rect 998 1512 1004 1513
rect 998 1508 999 1512
rect 1003 1508 1004 1512
rect 1158 1512 1159 1516
rect 1163 1512 1164 1516
rect 1158 1511 1164 1512
rect 1198 1516 1204 1517
rect 1198 1512 1199 1516
rect 1203 1512 1204 1516
rect 1198 1511 1204 1512
rect 1246 1516 1252 1517
rect 1246 1512 1247 1516
rect 1251 1512 1252 1516
rect 1246 1511 1252 1512
rect 1318 1516 1324 1517
rect 1318 1512 1319 1516
rect 1323 1512 1324 1516
rect 1318 1511 1324 1512
rect 1398 1516 1404 1517
rect 1398 1512 1399 1516
rect 1403 1512 1404 1516
rect 1398 1511 1404 1512
rect 1478 1516 1484 1517
rect 1478 1512 1479 1516
rect 1483 1512 1484 1516
rect 1478 1511 1484 1512
rect 1558 1516 1564 1517
rect 1558 1512 1559 1516
rect 1563 1512 1564 1516
rect 1558 1511 1564 1512
rect 1646 1516 1652 1517
rect 1646 1512 1647 1516
rect 1651 1512 1652 1516
rect 1646 1511 1652 1512
rect 1734 1516 1740 1517
rect 1734 1512 1735 1516
rect 1739 1512 1740 1516
rect 1734 1511 1740 1512
rect 1822 1516 1828 1517
rect 1822 1512 1823 1516
rect 1827 1512 1828 1516
rect 1822 1511 1828 1512
rect 1910 1516 1916 1517
rect 1910 1512 1911 1516
rect 1915 1512 1916 1516
rect 1910 1511 1916 1512
rect 1998 1516 2004 1517
rect 1998 1512 1999 1516
rect 2003 1512 2004 1516
rect 1998 1511 2004 1512
rect 2070 1516 2076 1517
rect 2070 1512 2071 1516
rect 2075 1512 2076 1516
rect 2118 1515 2119 1519
rect 2123 1515 2124 1519
rect 2118 1514 2124 1515
rect 2070 1511 2076 1512
rect 998 1507 1004 1508
rect 1158 1504 1164 1505
rect 1134 1501 1140 1502
rect 1134 1497 1135 1501
rect 1139 1497 1140 1501
rect 1158 1500 1159 1504
rect 1163 1500 1164 1504
rect 1158 1499 1164 1500
rect 1198 1504 1204 1505
rect 1198 1500 1199 1504
rect 1203 1500 1204 1504
rect 1198 1499 1204 1500
rect 1238 1504 1244 1505
rect 1238 1500 1239 1504
rect 1243 1500 1244 1504
rect 1238 1499 1244 1500
rect 1302 1504 1308 1505
rect 1302 1500 1303 1504
rect 1307 1500 1308 1504
rect 1302 1499 1308 1500
rect 1374 1504 1380 1505
rect 1374 1500 1375 1504
rect 1379 1500 1380 1504
rect 1374 1499 1380 1500
rect 1454 1504 1460 1505
rect 1454 1500 1455 1504
rect 1459 1500 1460 1504
rect 1454 1499 1460 1500
rect 1542 1504 1548 1505
rect 1542 1500 1543 1504
rect 1547 1500 1548 1504
rect 1542 1499 1548 1500
rect 1622 1504 1628 1505
rect 1622 1500 1623 1504
rect 1627 1500 1628 1504
rect 1622 1499 1628 1500
rect 1702 1504 1708 1505
rect 1702 1500 1703 1504
rect 1707 1500 1708 1504
rect 1702 1499 1708 1500
rect 1774 1504 1780 1505
rect 1774 1500 1775 1504
rect 1779 1500 1780 1504
rect 1774 1499 1780 1500
rect 1846 1504 1852 1505
rect 1846 1500 1847 1504
rect 1851 1500 1852 1504
rect 1846 1499 1852 1500
rect 1918 1504 1924 1505
rect 1918 1500 1919 1504
rect 1923 1500 1924 1504
rect 1918 1499 1924 1500
rect 1990 1504 1996 1505
rect 1990 1500 1991 1504
rect 1995 1500 1996 1504
rect 1990 1499 1996 1500
rect 2062 1504 2068 1505
rect 2062 1500 2063 1504
rect 2067 1500 2068 1504
rect 2062 1499 2068 1500
rect 2118 1501 2124 1502
rect 1134 1496 1140 1497
rect 2118 1497 2119 1501
rect 2123 1497 2124 1501
rect 2118 1496 2124 1497
rect 1134 1484 1140 1485
rect 1134 1480 1135 1484
rect 1139 1480 1140 1484
rect 1134 1479 1140 1480
rect 2118 1484 2124 1485
rect 2118 1480 2119 1484
rect 2123 1480 2124 1484
rect 2118 1479 2124 1480
rect 134 1476 140 1477
rect 134 1472 135 1476
rect 139 1472 140 1476
rect 134 1471 140 1472
rect 198 1476 204 1477
rect 198 1472 199 1476
rect 203 1472 204 1476
rect 198 1471 204 1472
rect 278 1476 284 1477
rect 278 1472 279 1476
rect 283 1472 284 1476
rect 278 1471 284 1472
rect 358 1476 364 1477
rect 358 1472 359 1476
rect 363 1472 364 1476
rect 358 1471 364 1472
rect 438 1476 444 1477
rect 438 1472 439 1476
rect 443 1472 444 1476
rect 438 1471 444 1472
rect 518 1476 524 1477
rect 518 1472 519 1476
rect 523 1472 524 1476
rect 518 1471 524 1472
rect 598 1476 604 1477
rect 598 1472 599 1476
rect 603 1472 604 1476
rect 598 1471 604 1472
rect 678 1476 684 1477
rect 678 1472 679 1476
rect 683 1472 684 1476
rect 678 1471 684 1472
rect 766 1476 772 1477
rect 766 1472 767 1476
rect 771 1472 772 1476
rect 766 1471 772 1472
rect 854 1476 860 1477
rect 854 1472 855 1476
rect 859 1472 860 1476
rect 854 1471 860 1472
rect 942 1476 948 1477
rect 942 1472 943 1476
rect 947 1472 948 1476
rect 942 1471 948 1472
rect 1030 1476 1036 1477
rect 1030 1472 1031 1476
rect 1035 1472 1036 1476
rect 1030 1471 1036 1472
rect 1158 1476 1164 1477
rect 1158 1472 1159 1476
rect 1163 1472 1164 1476
rect 1158 1471 1164 1472
rect 1198 1476 1204 1477
rect 1198 1472 1199 1476
rect 1203 1472 1204 1476
rect 1198 1471 1204 1472
rect 1238 1476 1244 1477
rect 1238 1472 1239 1476
rect 1243 1472 1244 1476
rect 1238 1471 1244 1472
rect 1302 1476 1308 1477
rect 1302 1472 1303 1476
rect 1307 1472 1308 1476
rect 1302 1471 1308 1472
rect 1374 1476 1380 1477
rect 1374 1472 1375 1476
rect 1379 1472 1380 1476
rect 1374 1471 1380 1472
rect 1454 1476 1460 1477
rect 1454 1472 1455 1476
rect 1459 1472 1460 1476
rect 1454 1471 1460 1472
rect 1542 1476 1548 1477
rect 1542 1472 1543 1476
rect 1547 1472 1548 1476
rect 1542 1471 1548 1472
rect 1622 1476 1628 1477
rect 1622 1472 1623 1476
rect 1627 1472 1628 1476
rect 1622 1471 1628 1472
rect 1702 1476 1708 1477
rect 1702 1472 1703 1476
rect 1707 1472 1708 1476
rect 1702 1471 1708 1472
rect 1774 1476 1780 1477
rect 1774 1472 1775 1476
rect 1779 1472 1780 1476
rect 1774 1471 1780 1472
rect 1846 1476 1852 1477
rect 1846 1472 1847 1476
rect 1851 1472 1852 1476
rect 1846 1471 1852 1472
rect 1918 1476 1924 1477
rect 1918 1472 1919 1476
rect 1923 1472 1924 1476
rect 1918 1471 1924 1472
rect 1990 1476 1996 1477
rect 1990 1472 1991 1476
rect 1995 1472 1996 1476
rect 1990 1471 1996 1472
rect 2062 1476 2068 1477
rect 2062 1472 2063 1476
rect 2067 1472 2068 1476
rect 2062 1471 2068 1472
rect 110 1468 116 1469
rect 110 1464 111 1468
rect 115 1464 116 1468
rect 110 1463 116 1464
rect 1094 1468 1100 1469
rect 1094 1464 1095 1468
rect 1099 1464 1100 1468
rect 1094 1463 1100 1464
rect 110 1451 116 1452
rect 110 1447 111 1451
rect 115 1447 116 1451
rect 1094 1451 1100 1452
rect 110 1446 116 1447
rect 134 1448 140 1449
rect 134 1444 135 1448
rect 139 1444 140 1448
rect 134 1443 140 1444
rect 198 1448 204 1449
rect 198 1444 199 1448
rect 203 1444 204 1448
rect 198 1443 204 1444
rect 278 1448 284 1449
rect 278 1444 279 1448
rect 283 1444 284 1448
rect 278 1443 284 1444
rect 358 1448 364 1449
rect 358 1444 359 1448
rect 363 1444 364 1448
rect 358 1443 364 1444
rect 438 1448 444 1449
rect 438 1444 439 1448
rect 443 1444 444 1448
rect 438 1443 444 1444
rect 518 1448 524 1449
rect 518 1444 519 1448
rect 523 1444 524 1448
rect 518 1443 524 1444
rect 598 1448 604 1449
rect 598 1444 599 1448
rect 603 1444 604 1448
rect 598 1443 604 1444
rect 678 1448 684 1449
rect 678 1444 679 1448
rect 683 1444 684 1448
rect 678 1443 684 1444
rect 766 1448 772 1449
rect 766 1444 767 1448
rect 771 1444 772 1448
rect 766 1443 772 1444
rect 854 1448 860 1449
rect 854 1444 855 1448
rect 859 1444 860 1448
rect 854 1443 860 1444
rect 942 1448 948 1449
rect 942 1444 943 1448
rect 947 1444 948 1448
rect 942 1443 948 1444
rect 1030 1448 1036 1449
rect 1030 1444 1031 1448
rect 1035 1444 1036 1448
rect 1094 1447 1095 1451
rect 1099 1447 1100 1451
rect 1094 1446 1100 1447
rect 1030 1443 1036 1444
rect 134 1436 140 1437
rect 110 1433 116 1434
rect 110 1429 111 1433
rect 115 1429 116 1433
rect 134 1432 135 1436
rect 139 1432 140 1436
rect 134 1431 140 1432
rect 190 1436 196 1437
rect 190 1432 191 1436
rect 195 1432 196 1436
rect 190 1431 196 1432
rect 262 1436 268 1437
rect 262 1432 263 1436
rect 267 1432 268 1436
rect 262 1431 268 1432
rect 334 1436 340 1437
rect 334 1432 335 1436
rect 339 1432 340 1436
rect 334 1431 340 1432
rect 406 1436 412 1437
rect 406 1432 407 1436
rect 411 1432 412 1436
rect 406 1431 412 1432
rect 478 1436 484 1437
rect 478 1432 479 1436
rect 483 1432 484 1436
rect 478 1431 484 1432
rect 550 1436 556 1437
rect 550 1432 551 1436
rect 555 1432 556 1436
rect 550 1431 556 1432
rect 630 1436 636 1437
rect 630 1432 631 1436
rect 635 1432 636 1436
rect 630 1431 636 1432
rect 710 1436 716 1437
rect 710 1432 711 1436
rect 715 1432 716 1436
rect 710 1431 716 1432
rect 798 1436 804 1437
rect 798 1432 799 1436
rect 803 1432 804 1436
rect 798 1431 804 1432
rect 886 1436 892 1437
rect 886 1432 887 1436
rect 891 1432 892 1436
rect 886 1431 892 1432
rect 974 1436 980 1437
rect 974 1432 975 1436
rect 979 1432 980 1436
rect 974 1431 980 1432
rect 1046 1436 1052 1437
rect 1046 1432 1047 1436
rect 1051 1432 1052 1436
rect 1278 1436 1284 1437
rect 1046 1431 1052 1432
rect 1094 1433 1100 1434
rect 110 1428 116 1429
rect 1094 1429 1095 1433
rect 1099 1429 1100 1433
rect 1278 1432 1279 1436
rect 1283 1432 1284 1436
rect 1278 1431 1284 1432
rect 1326 1436 1332 1437
rect 1326 1432 1327 1436
rect 1331 1432 1332 1436
rect 1326 1431 1332 1432
rect 1382 1436 1388 1437
rect 1382 1432 1383 1436
rect 1387 1432 1388 1436
rect 1382 1431 1388 1432
rect 1438 1436 1444 1437
rect 1438 1432 1439 1436
rect 1443 1432 1444 1436
rect 1438 1431 1444 1432
rect 1494 1436 1500 1437
rect 1494 1432 1495 1436
rect 1499 1432 1500 1436
rect 1494 1431 1500 1432
rect 1550 1436 1556 1437
rect 1550 1432 1551 1436
rect 1555 1432 1556 1436
rect 1550 1431 1556 1432
rect 1606 1436 1612 1437
rect 1606 1432 1607 1436
rect 1611 1432 1612 1436
rect 1606 1431 1612 1432
rect 1670 1436 1676 1437
rect 1670 1432 1671 1436
rect 1675 1432 1676 1436
rect 1670 1431 1676 1432
rect 1734 1436 1740 1437
rect 1734 1432 1735 1436
rect 1739 1432 1740 1436
rect 1734 1431 1740 1432
rect 1806 1436 1812 1437
rect 1806 1432 1807 1436
rect 1811 1432 1812 1436
rect 1806 1431 1812 1432
rect 1886 1436 1892 1437
rect 1886 1432 1887 1436
rect 1891 1432 1892 1436
rect 1886 1431 1892 1432
rect 1974 1436 1980 1437
rect 1974 1432 1975 1436
rect 1979 1432 1980 1436
rect 1974 1431 1980 1432
rect 2062 1436 2068 1437
rect 2062 1432 2063 1436
rect 2067 1432 2068 1436
rect 2062 1431 2068 1432
rect 1094 1428 1100 1429
rect 1134 1428 1140 1429
rect 1134 1424 1135 1428
rect 1139 1424 1140 1428
rect 1134 1423 1140 1424
rect 2118 1428 2124 1429
rect 2118 1424 2119 1428
rect 2123 1424 2124 1428
rect 2118 1423 2124 1424
rect 110 1416 116 1417
rect 110 1412 111 1416
rect 115 1412 116 1416
rect 110 1411 116 1412
rect 1094 1416 1100 1417
rect 1094 1412 1095 1416
rect 1099 1412 1100 1416
rect 1094 1411 1100 1412
rect 1134 1411 1140 1412
rect 134 1408 140 1409
rect 134 1404 135 1408
rect 139 1404 140 1408
rect 134 1403 140 1404
rect 190 1408 196 1409
rect 190 1404 191 1408
rect 195 1404 196 1408
rect 190 1403 196 1404
rect 262 1408 268 1409
rect 262 1404 263 1408
rect 267 1404 268 1408
rect 262 1403 268 1404
rect 334 1408 340 1409
rect 334 1404 335 1408
rect 339 1404 340 1408
rect 334 1403 340 1404
rect 406 1408 412 1409
rect 406 1404 407 1408
rect 411 1404 412 1408
rect 406 1403 412 1404
rect 478 1408 484 1409
rect 478 1404 479 1408
rect 483 1404 484 1408
rect 478 1403 484 1404
rect 550 1408 556 1409
rect 550 1404 551 1408
rect 555 1404 556 1408
rect 550 1403 556 1404
rect 630 1408 636 1409
rect 630 1404 631 1408
rect 635 1404 636 1408
rect 630 1403 636 1404
rect 710 1408 716 1409
rect 710 1404 711 1408
rect 715 1404 716 1408
rect 710 1403 716 1404
rect 798 1408 804 1409
rect 798 1404 799 1408
rect 803 1404 804 1408
rect 798 1403 804 1404
rect 886 1408 892 1409
rect 886 1404 887 1408
rect 891 1404 892 1408
rect 886 1403 892 1404
rect 974 1408 980 1409
rect 974 1404 975 1408
rect 979 1404 980 1408
rect 974 1403 980 1404
rect 1046 1408 1052 1409
rect 1046 1404 1047 1408
rect 1051 1404 1052 1408
rect 1134 1407 1135 1411
rect 1139 1407 1140 1411
rect 2118 1411 2124 1412
rect 1134 1406 1140 1407
rect 1278 1408 1284 1409
rect 1046 1403 1052 1404
rect 1278 1404 1279 1408
rect 1283 1404 1284 1408
rect 1278 1403 1284 1404
rect 1326 1408 1332 1409
rect 1326 1404 1327 1408
rect 1331 1404 1332 1408
rect 1326 1403 1332 1404
rect 1382 1408 1388 1409
rect 1382 1404 1383 1408
rect 1387 1404 1388 1408
rect 1382 1403 1388 1404
rect 1438 1408 1444 1409
rect 1438 1404 1439 1408
rect 1443 1404 1444 1408
rect 1438 1403 1444 1404
rect 1494 1408 1500 1409
rect 1494 1404 1495 1408
rect 1499 1404 1500 1408
rect 1494 1403 1500 1404
rect 1550 1408 1556 1409
rect 1550 1404 1551 1408
rect 1555 1404 1556 1408
rect 1550 1403 1556 1404
rect 1606 1408 1612 1409
rect 1606 1404 1607 1408
rect 1611 1404 1612 1408
rect 1606 1403 1612 1404
rect 1670 1408 1676 1409
rect 1670 1404 1671 1408
rect 1675 1404 1676 1408
rect 1670 1403 1676 1404
rect 1734 1408 1740 1409
rect 1734 1404 1735 1408
rect 1739 1404 1740 1408
rect 1734 1403 1740 1404
rect 1806 1408 1812 1409
rect 1806 1404 1807 1408
rect 1811 1404 1812 1408
rect 1806 1403 1812 1404
rect 1886 1408 1892 1409
rect 1886 1404 1887 1408
rect 1891 1404 1892 1408
rect 1886 1403 1892 1404
rect 1974 1408 1980 1409
rect 1974 1404 1975 1408
rect 1979 1404 1980 1408
rect 1974 1403 1980 1404
rect 2062 1408 2068 1409
rect 2062 1404 2063 1408
rect 2067 1404 2068 1408
rect 2118 1407 2119 1411
rect 2123 1407 2124 1411
rect 2118 1406 2124 1407
rect 2062 1403 2068 1404
rect 1334 1392 1340 1393
rect 1134 1389 1140 1390
rect 1134 1385 1135 1389
rect 1139 1385 1140 1389
rect 1334 1388 1335 1392
rect 1339 1388 1340 1392
rect 1334 1387 1340 1388
rect 1374 1392 1380 1393
rect 1374 1388 1375 1392
rect 1379 1388 1380 1392
rect 1374 1387 1380 1388
rect 1414 1392 1420 1393
rect 1414 1388 1415 1392
rect 1419 1388 1420 1392
rect 1414 1387 1420 1388
rect 1454 1392 1460 1393
rect 1454 1388 1455 1392
rect 1459 1388 1460 1392
rect 1454 1387 1460 1388
rect 1494 1392 1500 1393
rect 1494 1388 1495 1392
rect 1499 1388 1500 1392
rect 1494 1387 1500 1388
rect 1534 1392 1540 1393
rect 1534 1388 1535 1392
rect 1539 1388 1540 1392
rect 1534 1387 1540 1388
rect 1582 1392 1588 1393
rect 1582 1388 1583 1392
rect 1587 1388 1588 1392
rect 1582 1387 1588 1388
rect 1646 1392 1652 1393
rect 1646 1388 1647 1392
rect 1651 1388 1652 1392
rect 1646 1387 1652 1388
rect 1718 1392 1724 1393
rect 1718 1388 1719 1392
rect 1723 1388 1724 1392
rect 1718 1387 1724 1388
rect 1806 1392 1812 1393
rect 1806 1388 1807 1392
rect 1811 1388 1812 1392
rect 1806 1387 1812 1388
rect 1894 1392 1900 1393
rect 1894 1388 1895 1392
rect 1899 1388 1900 1392
rect 1894 1387 1900 1388
rect 1990 1392 1996 1393
rect 1990 1388 1991 1392
rect 1995 1388 1996 1392
rect 1990 1387 1996 1388
rect 2070 1392 2076 1393
rect 2070 1388 2071 1392
rect 2075 1388 2076 1392
rect 2070 1387 2076 1388
rect 2118 1389 2124 1390
rect 1134 1384 1140 1385
rect 2118 1385 2119 1389
rect 2123 1385 2124 1389
rect 2118 1384 2124 1385
rect 134 1372 140 1373
rect 134 1368 135 1372
rect 139 1368 140 1372
rect 134 1367 140 1368
rect 174 1372 180 1373
rect 174 1368 175 1372
rect 179 1368 180 1372
rect 174 1367 180 1368
rect 238 1372 244 1373
rect 238 1368 239 1372
rect 243 1368 244 1372
rect 238 1367 244 1368
rect 302 1372 308 1373
rect 302 1368 303 1372
rect 307 1368 308 1372
rect 302 1367 308 1368
rect 366 1372 372 1373
rect 366 1368 367 1372
rect 371 1368 372 1372
rect 366 1367 372 1368
rect 438 1372 444 1373
rect 438 1368 439 1372
rect 443 1368 444 1372
rect 438 1367 444 1368
rect 502 1372 508 1373
rect 502 1368 503 1372
rect 507 1368 508 1372
rect 502 1367 508 1368
rect 574 1372 580 1373
rect 574 1368 575 1372
rect 579 1368 580 1372
rect 574 1367 580 1368
rect 646 1372 652 1373
rect 646 1368 647 1372
rect 651 1368 652 1372
rect 646 1367 652 1368
rect 710 1372 716 1373
rect 710 1368 711 1372
rect 715 1368 716 1372
rect 710 1367 716 1368
rect 782 1372 788 1373
rect 782 1368 783 1372
rect 787 1368 788 1372
rect 782 1367 788 1368
rect 854 1372 860 1373
rect 854 1368 855 1372
rect 859 1368 860 1372
rect 854 1367 860 1368
rect 926 1372 932 1373
rect 926 1368 927 1372
rect 931 1368 932 1372
rect 926 1367 932 1368
rect 998 1372 1004 1373
rect 998 1368 999 1372
rect 1003 1368 1004 1372
rect 998 1367 1004 1368
rect 1046 1372 1052 1373
rect 1046 1368 1047 1372
rect 1051 1368 1052 1372
rect 1046 1367 1052 1368
rect 1134 1372 1140 1373
rect 1134 1368 1135 1372
rect 1139 1368 1140 1372
rect 1134 1367 1140 1368
rect 2118 1372 2124 1373
rect 2118 1368 2119 1372
rect 2123 1368 2124 1372
rect 2118 1367 2124 1368
rect 110 1364 116 1365
rect 110 1360 111 1364
rect 115 1360 116 1364
rect 110 1359 116 1360
rect 1094 1364 1100 1365
rect 1094 1360 1095 1364
rect 1099 1360 1100 1364
rect 1094 1359 1100 1360
rect 1334 1364 1340 1365
rect 1334 1360 1335 1364
rect 1339 1360 1340 1364
rect 1334 1359 1340 1360
rect 1374 1364 1380 1365
rect 1374 1360 1375 1364
rect 1379 1360 1380 1364
rect 1374 1359 1380 1360
rect 1414 1364 1420 1365
rect 1414 1360 1415 1364
rect 1419 1360 1420 1364
rect 1414 1359 1420 1360
rect 1454 1364 1460 1365
rect 1454 1360 1455 1364
rect 1459 1360 1460 1364
rect 1454 1359 1460 1360
rect 1494 1364 1500 1365
rect 1494 1360 1495 1364
rect 1499 1360 1500 1364
rect 1494 1359 1500 1360
rect 1534 1364 1540 1365
rect 1534 1360 1535 1364
rect 1539 1360 1540 1364
rect 1534 1359 1540 1360
rect 1582 1364 1588 1365
rect 1582 1360 1583 1364
rect 1587 1360 1588 1364
rect 1582 1359 1588 1360
rect 1646 1364 1652 1365
rect 1646 1360 1647 1364
rect 1651 1360 1652 1364
rect 1646 1359 1652 1360
rect 1718 1364 1724 1365
rect 1718 1360 1719 1364
rect 1723 1360 1724 1364
rect 1718 1359 1724 1360
rect 1806 1364 1812 1365
rect 1806 1360 1807 1364
rect 1811 1360 1812 1364
rect 1806 1359 1812 1360
rect 1894 1364 1900 1365
rect 1894 1360 1895 1364
rect 1899 1360 1900 1364
rect 1894 1359 1900 1360
rect 1990 1364 1996 1365
rect 1990 1360 1991 1364
rect 1995 1360 1996 1364
rect 1990 1359 1996 1360
rect 2070 1364 2076 1365
rect 2070 1360 2071 1364
rect 2075 1360 2076 1364
rect 2070 1359 2076 1360
rect 110 1347 116 1348
rect 110 1343 111 1347
rect 115 1343 116 1347
rect 1094 1347 1100 1348
rect 110 1342 116 1343
rect 134 1344 140 1345
rect 134 1340 135 1344
rect 139 1340 140 1344
rect 134 1339 140 1340
rect 174 1344 180 1345
rect 174 1340 175 1344
rect 179 1340 180 1344
rect 174 1339 180 1340
rect 238 1344 244 1345
rect 238 1340 239 1344
rect 243 1340 244 1344
rect 238 1339 244 1340
rect 302 1344 308 1345
rect 302 1340 303 1344
rect 307 1340 308 1344
rect 302 1339 308 1340
rect 366 1344 372 1345
rect 366 1340 367 1344
rect 371 1340 372 1344
rect 366 1339 372 1340
rect 438 1344 444 1345
rect 438 1340 439 1344
rect 443 1340 444 1344
rect 438 1339 444 1340
rect 502 1344 508 1345
rect 502 1340 503 1344
rect 507 1340 508 1344
rect 502 1339 508 1340
rect 574 1344 580 1345
rect 574 1340 575 1344
rect 579 1340 580 1344
rect 574 1339 580 1340
rect 646 1344 652 1345
rect 646 1340 647 1344
rect 651 1340 652 1344
rect 646 1339 652 1340
rect 710 1344 716 1345
rect 710 1340 711 1344
rect 715 1340 716 1344
rect 710 1339 716 1340
rect 782 1344 788 1345
rect 782 1340 783 1344
rect 787 1340 788 1344
rect 782 1339 788 1340
rect 854 1344 860 1345
rect 854 1340 855 1344
rect 859 1340 860 1344
rect 854 1339 860 1340
rect 926 1344 932 1345
rect 926 1340 927 1344
rect 931 1340 932 1344
rect 926 1339 932 1340
rect 998 1344 1004 1345
rect 998 1340 999 1344
rect 1003 1340 1004 1344
rect 998 1339 1004 1340
rect 1046 1344 1052 1345
rect 1046 1340 1047 1344
rect 1051 1340 1052 1344
rect 1094 1343 1095 1347
rect 1099 1343 1100 1347
rect 1094 1342 1100 1343
rect 1046 1339 1052 1340
rect 1158 1328 1164 1329
rect 134 1324 140 1325
rect 110 1321 116 1322
rect 110 1317 111 1321
rect 115 1317 116 1321
rect 134 1320 135 1324
rect 139 1320 140 1324
rect 134 1319 140 1320
rect 174 1324 180 1325
rect 174 1320 175 1324
rect 179 1320 180 1324
rect 174 1319 180 1320
rect 214 1324 220 1325
rect 214 1320 215 1324
rect 219 1320 220 1324
rect 214 1319 220 1320
rect 254 1324 260 1325
rect 254 1320 255 1324
rect 259 1320 260 1324
rect 254 1319 260 1320
rect 318 1324 324 1325
rect 318 1320 319 1324
rect 323 1320 324 1324
rect 318 1319 324 1320
rect 390 1324 396 1325
rect 390 1320 391 1324
rect 395 1320 396 1324
rect 390 1319 396 1320
rect 462 1324 468 1325
rect 462 1320 463 1324
rect 467 1320 468 1324
rect 462 1319 468 1320
rect 542 1324 548 1325
rect 542 1320 543 1324
rect 547 1320 548 1324
rect 542 1319 548 1320
rect 622 1324 628 1325
rect 622 1320 623 1324
rect 627 1320 628 1324
rect 622 1319 628 1320
rect 702 1324 708 1325
rect 702 1320 703 1324
rect 707 1320 708 1324
rect 702 1319 708 1320
rect 782 1324 788 1325
rect 782 1320 783 1324
rect 787 1320 788 1324
rect 782 1319 788 1320
rect 862 1324 868 1325
rect 862 1320 863 1324
rect 867 1320 868 1324
rect 862 1319 868 1320
rect 942 1324 948 1325
rect 942 1320 943 1324
rect 947 1320 948 1324
rect 942 1319 948 1320
rect 1022 1324 1028 1325
rect 1022 1320 1023 1324
rect 1027 1320 1028 1324
rect 1158 1324 1159 1328
rect 1163 1324 1164 1328
rect 1158 1323 1164 1324
rect 1222 1328 1228 1329
rect 1222 1324 1223 1328
rect 1227 1324 1228 1328
rect 1222 1323 1228 1324
rect 1310 1328 1316 1329
rect 1310 1324 1311 1328
rect 1315 1324 1316 1328
rect 1310 1323 1316 1324
rect 1406 1328 1412 1329
rect 1406 1324 1407 1328
rect 1411 1324 1412 1328
rect 1406 1323 1412 1324
rect 1502 1328 1508 1329
rect 1502 1324 1503 1328
rect 1507 1324 1508 1328
rect 1502 1323 1508 1324
rect 1598 1328 1604 1329
rect 1598 1324 1599 1328
rect 1603 1324 1604 1328
rect 1598 1323 1604 1324
rect 1678 1328 1684 1329
rect 1678 1324 1679 1328
rect 1683 1324 1684 1328
rect 1678 1323 1684 1324
rect 1758 1328 1764 1329
rect 1758 1324 1759 1328
rect 1763 1324 1764 1328
rect 1758 1323 1764 1324
rect 1830 1328 1836 1329
rect 1830 1324 1831 1328
rect 1835 1324 1836 1328
rect 1830 1323 1836 1324
rect 1894 1328 1900 1329
rect 1894 1324 1895 1328
rect 1899 1324 1900 1328
rect 1894 1323 1900 1324
rect 1958 1328 1964 1329
rect 1958 1324 1959 1328
rect 1963 1324 1964 1328
rect 1958 1323 1964 1324
rect 2022 1328 2028 1329
rect 2022 1324 2023 1328
rect 2027 1324 2028 1328
rect 2022 1323 2028 1324
rect 2070 1328 2076 1329
rect 2070 1324 2071 1328
rect 2075 1324 2076 1328
rect 2070 1323 2076 1324
rect 1022 1319 1028 1320
rect 1094 1321 1100 1322
rect 110 1316 116 1317
rect 1094 1317 1095 1321
rect 1099 1317 1100 1321
rect 1094 1316 1100 1317
rect 1134 1320 1140 1321
rect 1134 1316 1135 1320
rect 1139 1316 1140 1320
rect 1134 1315 1140 1316
rect 2118 1320 2124 1321
rect 2118 1316 2119 1320
rect 2123 1316 2124 1320
rect 2118 1315 2124 1316
rect 110 1304 116 1305
rect 110 1300 111 1304
rect 115 1300 116 1304
rect 110 1299 116 1300
rect 1094 1304 1100 1305
rect 1094 1300 1095 1304
rect 1099 1300 1100 1304
rect 1094 1299 1100 1300
rect 1134 1303 1140 1304
rect 1134 1299 1135 1303
rect 1139 1299 1140 1303
rect 2118 1303 2124 1304
rect 1134 1298 1140 1299
rect 1158 1300 1164 1301
rect 134 1296 140 1297
rect 134 1292 135 1296
rect 139 1292 140 1296
rect 134 1291 140 1292
rect 174 1296 180 1297
rect 174 1292 175 1296
rect 179 1292 180 1296
rect 174 1291 180 1292
rect 214 1296 220 1297
rect 214 1292 215 1296
rect 219 1292 220 1296
rect 214 1291 220 1292
rect 254 1296 260 1297
rect 254 1292 255 1296
rect 259 1292 260 1296
rect 254 1291 260 1292
rect 318 1296 324 1297
rect 318 1292 319 1296
rect 323 1292 324 1296
rect 318 1291 324 1292
rect 390 1296 396 1297
rect 390 1292 391 1296
rect 395 1292 396 1296
rect 390 1291 396 1292
rect 462 1296 468 1297
rect 462 1292 463 1296
rect 467 1292 468 1296
rect 462 1291 468 1292
rect 542 1296 548 1297
rect 542 1292 543 1296
rect 547 1292 548 1296
rect 542 1291 548 1292
rect 622 1296 628 1297
rect 622 1292 623 1296
rect 627 1292 628 1296
rect 622 1291 628 1292
rect 702 1296 708 1297
rect 702 1292 703 1296
rect 707 1292 708 1296
rect 702 1291 708 1292
rect 782 1296 788 1297
rect 782 1292 783 1296
rect 787 1292 788 1296
rect 782 1291 788 1292
rect 862 1296 868 1297
rect 862 1292 863 1296
rect 867 1292 868 1296
rect 862 1291 868 1292
rect 942 1296 948 1297
rect 942 1292 943 1296
rect 947 1292 948 1296
rect 942 1291 948 1292
rect 1022 1296 1028 1297
rect 1022 1292 1023 1296
rect 1027 1292 1028 1296
rect 1158 1296 1159 1300
rect 1163 1296 1164 1300
rect 1158 1295 1164 1296
rect 1222 1300 1228 1301
rect 1222 1296 1223 1300
rect 1227 1296 1228 1300
rect 1222 1295 1228 1296
rect 1310 1300 1316 1301
rect 1310 1296 1311 1300
rect 1315 1296 1316 1300
rect 1310 1295 1316 1296
rect 1406 1300 1412 1301
rect 1406 1296 1407 1300
rect 1411 1296 1412 1300
rect 1406 1295 1412 1296
rect 1502 1300 1508 1301
rect 1502 1296 1503 1300
rect 1507 1296 1508 1300
rect 1502 1295 1508 1296
rect 1598 1300 1604 1301
rect 1598 1296 1599 1300
rect 1603 1296 1604 1300
rect 1598 1295 1604 1296
rect 1678 1300 1684 1301
rect 1678 1296 1679 1300
rect 1683 1296 1684 1300
rect 1678 1295 1684 1296
rect 1758 1300 1764 1301
rect 1758 1296 1759 1300
rect 1763 1296 1764 1300
rect 1758 1295 1764 1296
rect 1830 1300 1836 1301
rect 1830 1296 1831 1300
rect 1835 1296 1836 1300
rect 1830 1295 1836 1296
rect 1894 1300 1900 1301
rect 1894 1296 1895 1300
rect 1899 1296 1900 1300
rect 1894 1295 1900 1296
rect 1958 1300 1964 1301
rect 1958 1296 1959 1300
rect 1963 1296 1964 1300
rect 1958 1295 1964 1296
rect 2022 1300 2028 1301
rect 2022 1296 2023 1300
rect 2027 1296 2028 1300
rect 2022 1295 2028 1296
rect 2070 1300 2076 1301
rect 2070 1296 2071 1300
rect 2075 1296 2076 1300
rect 2118 1299 2119 1303
rect 2123 1299 2124 1303
rect 2118 1298 2124 1299
rect 2070 1295 2076 1296
rect 1022 1291 1028 1292
rect 1174 1288 1180 1289
rect 1134 1285 1140 1286
rect 1134 1281 1135 1285
rect 1139 1281 1140 1285
rect 1174 1284 1175 1288
rect 1179 1284 1180 1288
rect 1174 1283 1180 1284
rect 1230 1288 1236 1289
rect 1230 1284 1231 1288
rect 1235 1284 1236 1288
rect 1230 1283 1236 1284
rect 1302 1288 1308 1289
rect 1302 1284 1303 1288
rect 1307 1284 1308 1288
rect 1302 1283 1308 1284
rect 1390 1288 1396 1289
rect 1390 1284 1391 1288
rect 1395 1284 1396 1288
rect 1390 1283 1396 1284
rect 1478 1288 1484 1289
rect 1478 1284 1479 1288
rect 1483 1284 1484 1288
rect 1478 1283 1484 1284
rect 1566 1288 1572 1289
rect 1566 1284 1567 1288
rect 1571 1284 1572 1288
rect 1566 1283 1572 1284
rect 1654 1288 1660 1289
rect 1654 1284 1655 1288
rect 1659 1284 1660 1288
rect 1654 1283 1660 1284
rect 1742 1288 1748 1289
rect 1742 1284 1743 1288
rect 1747 1284 1748 1288
rect 1742 1283 1748 1284
rect 1830 1288 1836 1289
rect 1830 1284 1831 1288
rect 1835 1284 1836 1288
rect 1830 1283 1836 1284
rect 1918 1288 1924 1289
rect 1918 1284 1919 1288
rect 1923 1284 1924 1288
rect 1918 1283 1924 1284
rect 2006 1288 2012 1289
rect 2006 1284 2007 1288
rect 2011 1284 2012 1288
rect 2006 1283 2012 1284
rect 2070 1288 2076 1289
rect 2070 1284 2071 1288
rect 2075 1284 2076 1288
rect 2070 1283 2076 1284
rect 2118 1285 2124 1286
rect 1134 1280 1140 1281
rect 2118 1281 2119 1285
rect 2123 1281 2124 1285
rect 2118 1280 2124 1281
rect 1134 1268 1140 1269
rect 1134 1264 1135 1268
rect 1139 1264 1140 1268
rect 1134 1263 1140 1264
rect 2118 1268 2124 1269
rect 2118 1264 2119 1268
rect 2123 1264 2124 1268
rect 2118 1263 2124 1264
rect 1174 1260 1180 1261
rect 134 1256 140 1257
rect 134 1252 135 1256
rect 139 1252 140 1256
rect 134 1251 140 1252
rect 174 1256 180 1257
rect 174 1252 175 1256
rect 179 1252 180 1256
rect 174 1251 180 1252
rect 214 1256 220 1257
rect 214 1252 215 1256
rect 219 1252 220 1256
rect 214 1251 220 1252
rect 254 1256 260 1257
rect 254 1252 255 1256
rect 259 1252 260 1256
rect 254 1251 260 1252
rect 318 1256 324 1257
rect 318 1252 319 1256
rect 323 1252 324 1256
rect 318 1251 324 1252
rect 398 1256 404 1257
rect 398 1252 399 1256
rect 403 1252 404 1256
rect 398 1251 404 1252
rect 486 1256 492 1257
rect 486 1252 487 1256
rect 491 1252 492 1256
rect 486 1251 492 1252
rect 582 1256 588 1257
rect 582 1252 583 1256
rect 587 1252 588 1256
rect 582 1251 588 1252
rect 686 1256 692 1257
rect 686 1252 687 1256
rect 691 1252 692 1256
rect 686 1251 692 1252
rect 798 1256 804 1257
rect 798 1252 799 1256
rect 803 1252 804 1256
rect 798 1251 804 1252
rect 918 1256 924 1257
rect 918 1252 919 1256
rect 923 1252 924 1256
rect 918 1251 924 1252
rect 1046 1256 1052 1257
rect 1046 1252 1047 1256
rect 1051 1252 1052 1256
rect 1174 1256 1175 1260
rect 1179 1256 1180 1260
rect 1174 1255 1180 1256
rect 1230 1260 1236 1261
rect 1230 1256 1231 1260
rect 1235 1256 1236 1260
rect 1230 1255 1236 1256
rect 1302 1260 1308 1261
rect 1302 1256 1303 1260
rect 1307 1256 1308 1260
rect 1302 1255 1308 1256
rect 1390 1260 1396 1261
rect 1390 1256 1391 1260
rect 1395 1256 1396 1260
rect 1390 1255 1396 1256
rect 1478 1260 1484 1261
rect 1478 1256 1479 1260
rect 1483 1256 1484 1260
rect 1478 1255 1484 1256
rect 1566 1260 1572 1261
rect 1566 1256 1567 1260
rect 1571 1256 1572 1260
rect 1566 1255 1572 1256
rect 1654 1260 1660 1261
rect 1654 1256 1655 1260
rect 1659 1256 1660 1260
rect 1654 1255 1660 1256
rect 1742 1260 1748 1261
rect 1742 1256 1743 1260
rect 1747 1256 1748 1260
rect 1742 1255 1748 1256
rect 1830 1260 1836 1261
rect 1830 1256 1831 1260
rect 1835 1256 1836 1260
rect 1830 1255 1836 1256
rect 1918 1260 1924 1261
rect 1918 1256 1919 1260
rect 1923 1256 1924 1260
rect 1918 1255 1924 1256
rect 2006 1260 2012 1261
rect 2006 1256 2007 1260
rect 2011 1256 2012 1260
rect 2006 1255 2012 1256
rect 2070 1260 2076 1261
rect 2070 1256 2071 1260
rect 2075 1256 2076 1260
rect 2070 1255 2076 1256
rect 1046 1251 1052 1252
rect 110 1248 116 1249
rect 110 1244 111 1248
rect 115 1244 116 1248
rect 110 1243 116 1244
rect 1094 1248 1100 1249
rect 1094 1244 1095 1248
rect 1099 1244 1100 1248
rect 1094 1243 1100 1244
rect 110 1231 116 1232
rect 110 1227 111 1231
rect 115 1227 116 1231
rect 1094 1231 1100 1232
rect 110 1226 116 1227
rect 134 1228 140 1229
rect 134 1224 135 1228
rect 139 1224 140 1228
rect 134 1223 140 1224
rect 174 1228 180 1229
rect 174 1224 175 1228
rect 179 1224 180 1228
rect 174 1223 180 1224
rect 214 1228 220 1229
rect 214 1224 215 1228
rect 219 1224 220 1228
rect 214 1223 220 1224
rect 254 1228 260 1229
rect 254 1224 255 1228
rect 259 1224 260 1228
rect 254 1223 260 1224
rect 318 1228 324 1229
rect 318 1224 319 1228
rect 323 1224 324 1228
rect 318 1223 324 1224
rect 398 1228 404 1229
rect 398 1224 399 1228
rect 403 1224 404 1228
rect 398 1223 404 1224
rect 486 1228 492 1229
rect 486 1224 487 1228
rect 491 1224 492 1228
rect 486 1223 492 1224
rect 582 1228 588 1229
rect 582 1224 583 1228
rect 587 1224 588 1228
rect 582 1223 588 1224
rect 686 1228 692 1229
rect 686 1224 687 1228
rect 691 1224 692 1228
rect 686 1223 692 1224
rect 798 1228 804 1229
rect 798 1224 799 1228
rect 803 1224 804 1228
rect 798 1223 804 1224
rect 918 1228 924 1229
rect 918 1224 919 1228
rect 923 1224 924 1228
rect 918 1223 924 1224
rect 1046 1228 1052 1229
rect 1046 1224 1047 1228
rect 1051 1224 1052 1228
rect 1094 1227 1095 1231
rect 1099 1227 1100 1231
rect 1094 1226 1100 1227
rect 1046 1223 1052 1224
rect 1286 1220 1292 1221
rect 1286 1216 1287 1220
rect 1291 1216 1292 1220
rect 1286 1215 1292 1216
rect 1326 1220 1332 1221
rect 1326 1216 1327 1220
rect 1331 1216 1332 1220
rect 1326 1215 1332 1216
rect 1374 1220 1380 1221
rect 1374 1216 1375 1220
rect 1379 1216 1380 1220
rect 1374 1215 1380 1216
rect 1430 1220 1436 1221
rect 1430 1216 1431 1220
rect 1435 1216 1436 1220
rect 1430 1215 1436 1216
rect 1494 1220 1500 1221
rect 1494 1216 1495 1220
rect 1499 1216 1500 1220
rect 1494 1215 1500 1216
rect 1558 1220 1564 1221
rect 1558 1216 1559 1220
rect 1563 1216 1564 1220
rect 1558 1215 1564 1216
rect 1622 1220 1628 1221
rect 1622 1216 1623 1220
rect 1627 1216 1628 1220
rect 1622 1215 1628 1216
rect 1678 1220 1684 1221
rect 1678 1216 1679 1220
rect 1683 1216 1684 1220
rect 1678 1215 1684 1216
rect 1734 1220 1740 1221
rect 1734 1216 1735 1220
rect 1739 1216 1740 1220
rect 1734 1215 1740 1216
rect 1790 1220 1796 1221
rect 1790 1216 1791 1220
rect 1795 1216 1796 1220
rect 1790 1215 1796 1216
rect 1846 1220 1852 1221
rect 1846 1216 1847 1220
rect 1851 1216 1852 1220
rect 1846 1215 1852 1216
rect 1902 1220 1908 1221
rect 1902 1216 1903 1220
rect 1907 1216 1908 1220
rect 1902 1215 1908 1216
rect 1966 1220 1972 1221
rect 1966 1216 1967 1220
rect 1971 1216 1972 1220
rect 1966 1215 1972 1216
rect 2030 1220 2036 1221
rect 2030 1216 2031 1220
rect 2035 1216 2036 1220
rect 2030 1215 2036 1216
rect 2070 1220 2076 1221
rect 2070 1216 2071 1220
rect 2075 1216 2076 1220
rect 2070 1215 2076 1216
rect 270 1212 276 1213
rect 110 1209 116 1210
rect 110 1205 111 1209
rect 115 1205 116 1209
rect 270 1208 271 1212
rect 275 1208 276 1212
rect 270 1207 276 1208
rect 310 1212 316 1213
rect 310 1208 311 1212
rect 315 1208 316 1212
rect 310 1207 316 1208
rect 350 1212 356 1213
rect 350 1208 351 1212
rect 355 1208 356 1212
rect 350 1207 356 1208
rect 398 1212 404 1213
rect 398 1208 399 1212
rect 403 1208 404 1212
rect 398 1207 404 1208
rect 446 1212 452 1213
rect 446 1208 447 1212
rect 451 1208 452 1212
rect 446 1207 452 1208
rect 494 1212 500 1213
rect 494 1208 495 1212
rect 499 1208 500 1212
rect 494 1207 500 1208
rect 550 1212 556 1213
rect 550 1208 551 1212
rect 555 1208 556 1212
rect 550 1207 556 1208
rect 606 1212 612 1213
rect 606 1208 607 1212
rect 611 1208 612 1212
rect 606 1207 612 1208
rect 670 1212 676 1213
rect 670 1208 671 1212
rect 675 1208 676 1212
rect 670 1207 676 1208
rect 742 1212 748 1213
rect 742 1208 743 1212
rect 747 1208 748 1212
rect 742 1207 748 1208
rect 814 1212 820 1213
rect 814 1208 815 1212
rect 819 1208 820 1212
rect 814 1207 820 1208
rect 894 1212 900 1213
rect 894 1208 895 1212
rect 899 1208 900 1212
rect 894 1207 900 1208
rect 982 1212 988 1213
rect 982 1208 983 1212
rect 987 1208 988 1212
rect 1134 1212 1140 1213
rect 982 1207 988 1208
rect 1094 1209 1100 1210
rect 110 1204 116 1205
rect 1094 1205 1095 1209
rect 1099 1205 1100 1209
rect 1134 1208 1135 1212
rect 1139 1208 1140 1212
rect 1134 1207 1140 1208
rect 2118 1212 2124 1213
rect 2118 1208 2119 1212
rect 2123 1208 2124 1212
rect 2118 1207 2124 1208
rect 1094 1204 1100 1205
rect 1134 1195 1140 1196
rect 110 1192 116 1193
rect 110 1188 111 1192
rect 115 1188 116 1192
rect 110 1187 116 1188
rect 1094 1192 1100 1193
rect 1094 1188 1095 1192
rect 1099 1188 1100 1192
rect 1134 1191 1135 1195
rect 1139 1191 1140 1195
rect 2118 1195 2124 1196
rect 1134 1190 1140 1191
rect 1286 1192 1292 1193
rect 1094 1187 1100 1188
rect 1286 1188 1287 1192
rect 1291 1188 1292 1192
rect 1286 1187 1292 1188
rect 1326 1192 1332 1193
rect 1326 1188 1327 1192
rect 1331 1188 1332 1192
rect 1326 1187 1332 1188
rect 1374 1192 1380 1193
rect 1374 1188 1375 1192
rect 1379 1188 1380 1192
rect 1374 1187 1380 1188
rect 1430 1192 1436 1193
rect 1430 1188 1431 1192
rect 1435 1188 1436 1192
rect 1430 1187 1436 1188
rect 1494 1192 1500 1193
rect 1494 1188 1495 1192
rect 1499 1188 1500 1192
rect 1494 1187 1500 1188
rect 1558 1192 1564 1193
rect 1558 1188 1559 1192
rect 1563 1188 1564 1192
rect 1558 1187 1564 1188
rect 1622 1192 1628 1193
rect 1622 1188 1623 1192
rect 1627 1188 1628 1192
rect 1622 1187 1628 1188
rect 1678 1192 1684 1193
rect 1678 1188 1679 1192
rect 1683 1188 1684 1192
rect 1678 1187 1684 1188
rect 1734 1192 1740 1193
rect 1734 1188 1735 1192
rect 1739 1188 1740 1192
rect 1734 1187 1740 1188
rect 1790 1192 1796 1193
rect 1790 1188 1791 1192
rect 1795 1188 1796 1192
rect 1790 1187 1796 1188
rect 1846 1192 1852 1193
rect 1846 1188 1847 1192
rect 1851 1188 1852 1192
rect 1846 1187 1852 1188
rect 1902 1192 1908 1193
rect 1902 1188 1903 1192
rect 1907 1188 1908 1192
rect 1902 1187 1908 1188
rect 1966 1192 1972 1193
rect 1966 1188 1967 1192
rect 1971 1188 1972 1192
rect 1966 1187 1972 1188
rect 2030 1192 2036 1193
rect 2030 1188 2031 1192
rect 2035 1188 2036 1192
rect 2030 1187 2036 1188
rect 2070 1192 2076 1193
rect 2070 1188 2071 1192
rect 2075 1188 2076 1192
rect 2118 1191 2119 1195
rect 2123 1191 2124 1195
rect 2118 1190 2124 1191
rect 2070 1187 2076 1188
rect 270 1184 276 1185
rect 270 1180 271 1184
rect 275 1180 276 1184
rect 270 1179 276 1180
rect 310 1184 316 1185
rect 310 1180 311 1184
rect 315 1180 316 1184
rect 310 1179 316 1180
rect 350 1184 356 1185
rect 350 1180 351 1184
rect 355 1180 356 1184
rect 350 1179 356 1180
rect 398 1184 404 1185
rect 398 1180 399 1184
rect 403 1180 404 1184
rect 398 1179 404 1180
rect 446 1184 452 1185
rect 446 1180 447 1184
rect 451 1180 452 1184
rect 446 1179 452 1180
rect 494 1184 500 1185
rect 494 1180 495 1184
rect 499 1180 500 1184
rect 494 1179 500 1180
rect 550 1184 556 1185
rect 550 1180 551 1184
rect 555 1180 556 1184
rect 550 1179 556 1180
rect 606 1184 612 1185
rect 606 1180 607 1184
rect 611 1180 612 1184
rect 606 1179 612 1180
rect 670 1184 676 1185
rect 670 1180 671 1184
rect 675 1180 676 1184
rect 670 1179 676 1180
rect 742 1184 748 1185
rect 742 1180 743 1184
rect 747 1180 748 1184
rect 742 1179 748 1180
rect 814 1184 820 1185
rect 814 1180 815 1184
rect 819 1180 820 1184
rect 814 1179 820 1180
rect 894 1184 900 1185
rect 894 1180 895 1184
rect 899 1180 900 1184
rect 894 1179 900 1180
rect 982 1184 988 1185
rect 982 1180 983 1184
rect 987 1180 988 1184
rect 982 1179 988 1180
rect 1158 1180 1164 1181
rect 1134 1177 1140 1178
rect 1134 1173 1135 1177
rect 1139 1173 1140 1177
rect 1158 1176 1159 1180
rect 1163 1176 1164 1180
rect 1158 1175 1164 1176
rect 1206 1180 1212 1181
rect 1206 1176 1207 1180
rect 1211 1176 1212 1180
rect 1206 1175 1212 1176
rect 1278 1180 1284 1181
rect 1278 1176 1279 1180
rect 1283 1176 1284 1180
rect 1278 1175 1284 1176
rect 1350 1180 1356 1181
rect 1350 1176 1351 1180
rect 1355 1176 1356 1180
rect 1350 1175 1356 1176
rect 1422 1180 1428 1181
rect 1422 1176 1423 1180
rect 1427 1176 1428 1180
rect 1422 1175 1428 1176
rect 1486 1180 1492 1181
rect 1486 1176 1487 1180
rect 1491 1176 1492 1180
rect 1486 1175 1492 1176
rect 1558 1180 1564 1181
rect 1558 1176 1559 1180
rect 1563 1176 1564 1180
rect 1558 1175 1564 1176
rect 1630 1180 1636 1181
rect 1630 1176 1631 1180
rect 1635 1176 1636 1180
rect 1630 1175 1636 1176
rect 1710 1180 1716 1181
rect 1710 1176 1711 1180
rect 1715 1176 1716 1180
rect 1710 1175 1716 1176
rect 1798 1180 1804 1181
rect 1798 1176 1799 1180
rect 1803 1176 1804 1180
rect 1798 1175 1804 1176
rect 1886 1180 1892 1181
rect 1886 1176 1887 1180
rect 1891 1176 1892 1180
rect 1886 1175 1892 1176
rect 1982 1180 1988 1181
rect 1982 1176 1983 1180
rect 1987 1176 1988 1180
rect 1982 1175 1988 1176
rect 2070 1180 2076 1181
rect 2070 1176 2071 1180
rect 2075 1176 2076 1180
rect 2070 1175 2076 1176
rect 2118 1177 2124 1178
rect 1134 1172 1140 1173
rect 2118 1173 2119 1177
rect 2123 1173 2124 1177
rect 2118 1172 2124 1173
rect 1134 1160 1140 1161
rect 1134 1156 1135 1160
rect 1139 1156 1140 1160
rect 1134 1155 1140 1156
rect 2118 1160 2124 1161
rect 2118 1156 2119 1160
rect 2123 1156 2124 1160
rect 2118 1155 2124 1156
rect 1158 1152 1164 1153
rect 1158 1148 1159 1152
rect 1163 1148 1164 1152
rect 1158 1147 1164 1148
rect 1206 1152 1212 1153
rect 1206 1148 1207 1152
rect 1211 1148 1212 1152
rect 1206 1147 1212 1148
rect 1278 1152 1284 1153
rect 1278 1148 1279 1152
rect 1283 1148 1284 1152
rect 1278 1147 1284 1148
rect 1350 1152 1356 1153
rect 1350 1148 1351 1152
rect 1355 1148 1356 1152
rect 1350 1147 1356 1148
rect 1422 1152 1428 1153
rect 1422 1148 1423 1152
rect 1427 1148 1428 1152
rect 1422 1147 1428 1148
rect 1486 1152 1492 1153
rect 1486 1148 1487 1152
rect 1491 1148 1492 1152
rect 1486 1147 1492 1148
rect 1558 1152 1564 1153
rect 1558 1148 1559 1152
rect 1563 1148 1564 1152
rect 1558 1147 1564 1148
rect 1630 1152 1636 1153
rect 1630 1148 1631 1152
rect 1635 1148 1636 1152
rect 1630 1147 1636 1148
rect 1710 1152 1716 1153
rect 1710 1148 1711 1152
rect 1715 1148 1716 1152
rect 1710 1147 1716 1148
rect 1798 1152 1804 1153
rect 1798 1148 1799 1152
rect 1803 1148 1804 1152
rect 1798 1147 1804 1148
rect 1886 1152 1892 1153
rect 1886 1148 1887 1152
rect 1891 1148 1892 1152
rect 1886 1147 1892 1148
rect 1982 1152 1988 1153
rect 1982 1148 1983 1152
rect 1987 1148 1988 1152
rect 1982 1147 1988 1148
rect 2070 1152 2076 1153
rect 2070 1148 2071 1152
rect 2075 1148 2076 1152
rect 2070 1147 2076 1148
rect 398 1144 404 1145
rect 398 1140 399 1144
rect 403 1140 404 1144
rect 398 1139 404 1140
rect 438 1144 444 1145
rect 438 1140 439 1144
rect 443 1140 444 1144
rect 438 1139 444 1140
rect 478 1144 484 1145
rect 478 1140 479 1144
rect 483 1140 484 1144
rect 478 1139 484 1140
rect 526 1144 532 1145
rect 526 1140 527 1144
rect 531 1140 532 1144
rect 526 1139 532 1140
rect 574 1144 580 1145
rect 574 1140 575 1144
rect 579 1140 580 1144
rect 574 1139 580 1140
rect 622 1144 628 1145
rect 622 1140 623 1144
rect 627 1140 628 1144
rect 622 1139 628 1140
rect 670 1144 676 1145
rect 670 1140 671 1144
rect 675 1140 676 1144
rect 670 1139 676 1140
rect 718 1144 724 1145
rect 718 1140 719 1144
rect 723 1140 724 1144
rect 718 1139 724 1140
rect 774 1144 780 1145
rect 774 1140 775 1144
rect 779 1140 780 1144
rect 774 1139 780 1140
rect 830 1144 836 1145
rect 830 1140 831 1144
rect 835 1140 836 1144
rect 830 1139 836 1140
rect 886 1144 892 1145
rect 886 1140 887 1144
rect 891 1140 892 1144
rect 886 1139 892 1140
rect 942 1144 948 1145
rect 942 1140 943 1144
rect 947 1140 948 1144
rect 942 1139 948 1140
rect 1006 1144 1012 1145
rect 1006 1140 1007 1144
rect 1011 1140 1012 1144
rect 1006 1139 1012 1140
rect 1046 1144 1052 1145
rect 1046 1140 1047 1144
rect 1051 1140 1052 1144
rect 1046 1139 1052 1140
rect 110 1136 116 1137
rect 110 1132 111 1136
rect 115 1132 116 1136
rect 110 1131 116 1132
rect 1094 1136 1100 1137
rect 1094 1132 1095 1136
rect 1099 1132 1100 1136
rect 1094 1131 1100 1132
rect 110 1119 116 1120
rect 110 1115 111 1119
rect 115 1115 116 1119
rect 1094 1119 1100 1120
rect 110 1114 116 1115
rect 398 1116 404 1117
rect 398 1112 399 1116
rect 403 1112 404 1116
rect 398 1111 404 1112
rect 438 1116 444 1117
rect 438 1112 439 1116
rect 443 1112 444 1116
rect 438 1111 444 1112
rect 478 1116 484 1117
rect 478 1112 479 1116
rect 483 1112 484 1116
rect 478 1111 484 1112
rect 526 1116 532 1117
rect 526 1112 527 1116
rect 531 1112 532 1116
rect 526 1111 532 1112
rect 574 1116 580 1117
rect 574 1112 575 1116
rect 579 1112 580 1116
rect 574 1111 580 1112
rect 622 1116 628 1117
rect 622 1112 623 1116
rect 627 1112 628 1116
rect 622 1111 628 1112
rect 670 1116 676 1117
rect 670 1112 671 1116
rect 675 1112 676 1116
rect 670 1111 676 1112
rect 718 1116 724 1117
rect 718 1112 719 1116
rect 723 1112 724 1116
rect 718 1111 724 1112
rect 774 1116 780 1117
rect 774 1112 775 1116
rect 779 1112 780 1116
rect 774 1111 780 1112
rect 830 1116 836 1117
rect 830 1112 831 1116
rect 835 1112 836 1116
rect 830 1111 836 1112
rect 886 1116 892 1117
rect 886 1112 887 1116
rect 891 1112 892 1116
rect 886 1111 892 1112
rect 942 1116 948 1117
rect 942 1112 943 1116
rect 947 1112 948 1116
rect 942 1111 948 1112
rect 1006 1116 1012 1117
rect 1006 1112 1007 1116
rect 1011 1112 1012 1116
rect 1006 1111 1012 1112
rect 1046 1116 1052 1117
rect 1046 1112 1047 1116
rect 1051 1112 1052 1116
rect 1094 1115 1095 1119
rect 1099 1115 1100 1119
rect 1094 1114 1100 1115
rect 1046 1111 1052 1112
rect 1190 1112 1196 1113
rect 1190 1108 1191 1112
rect 1195 1108 1196 1112
rect 1190 1107 1196 1108
rect 1270 1112 1276 1113
rect 1270 1108 1271 1112
rect 1275 1108 1276 1112
rect 1270 1107 1276 1108
rect 1342 1112 1348 1113
rect 1342 1108 1343 1112
rect 1347 1108 1348 1112
rect 1342 1107 1348 1108
rect 1414 1112 1420 1113
rect 1414 1108 1415 1112
rect 1419 1108 1420 1112
rect 1414 1107 1420 1108
rect 1486 1112 1492 1113
rect 1486 1108 1487 1112
rect 1491 1108 1492 1112
rect 1486 1107 1492 1108
rect 1566 1112 1572 1113
rect 1566 1108 1567 1112
rect 1571 1108 1572 1112
rect 1566 1107 1572 1108
rect 1654 1112 1660 1113
rect 1654 1108 1655 1112
rect 1659 1108 1660 1112
rect 1654 1107 1660 1108
rect 1750 1112 1756 1113
rect 1750 1108 1751 1112
rect 1755 1108 1756 1112
rect 1750 1107 1756 1108
rect 1854 1112 1860 1113
rect 1854 1108 1855 1112
rect 1859 1108 1860 1112
rect 1854 1107 1860 1108
rect 1958 1112 1964 1113
rect 1958 1108 1959 1112
rect 1963 1108 1964 1112
rect 1958 1107 1964 1108
rect 2070 1112 2076 1113
rect 2070 1108 2071 1112
rect 2075 1108 2076 1112
rect 2070 1107 2076 1108
rect 158 1104 164 1105
rect 110 1101 116 1102
rect 110 1097 111 1101
rect 115 1097 116 1101
rect 158 1100 159 1104
rect 163 1100 164 1104
rect 158 1099 164 1100
rect 198 1104 204 1105
rect 198 1100 199 1104
rect 203 1100 204 1104
rect 198 1099 204 1100
rect 254 1104 260 1105
rect 254 1100 255 1104
rect 259 1100 260 1104
rect 254 1099 260 1100
rect 318 1104 324 1105
rect 318 1100 319 1104
rect 323 1100 324 1104
rect 318 1099 324 1100
rect 398 1104 404 1105
rect 398 1100 399 1104
rect 403 1100 404 1104
rect 398 1099 404 1100
rect 478 1104 484 1105
rect 478 1100 479 1104
rect 483 1100 484 1104
rect 478 1099 484 1100
rect 558 1104 564 1105
rect 558 1100 559 1104
rect 563 1100 564 1104
rect 558 1099 564 1100
rect 638 1104 644 1105
rect 638 1100 639 1104
rect 643 1100 644 1104
rect 638 1099 644 1100
rect 710 1104 716 1105
rect 710 1100 711 1104
rect 715 1100 716 1104
rect 710 1099 716 1100
rect 782 1104 788 1105
rect 782 1100 783 1104
rect 787 1100 788 1104
rect 782 1099 788 1100
rect 854 1104 860 1105
rect 854 1100 855 1104
rect 859 1100 860 1104
rect 854 1099 860 1100
rect 926 1104 932 1105
rect 926 1100 927 1104
rect 931 1100 932 1104
rect 926 1099 932 1100
rect 998 1104 1004 1105
rect 998 1100 999 1104
rect 1003 1100 1004 1104
rect 998 1099 1004 1100
rect 1046 1104 1052 1105
rect 1046 1100 1047 1104
rect 1051 1100 1052 1104
rect 1134 1104 1140 1105
rect 1046 1099 1052 1100
rect 1094 1101 1100 1102
rect 110 1096 116 1097
rect 1094 1097 1095 1101
rect 1099 1097 1100 1101
rect 1134 1100 1135 1104
rect 1139 1100 1140 1104
rect 1134 1099 1140 1100
rect 2118 1104 2124 1105
rect 2118 1100 2119 1104
rect 2123 1100 2124 1104
rect 2118 1099 2124 1100
rect 1094 1096 1100 1097
rect 1134 1087 1140 1088
rect 110 1084 116 1085
rect 110 1080 111 1084
rect 115 1080 116 1084
rect 110 1079 116 1080
rect 1094 1084 1100 1085
rect 1094 1080 1095 1084
rect 1099 1080 1100 1084
rect 1134 1083 1135 1087
rect 1139 1083 1140 1087
rect 2118 1087 2124 1088
rect 1134 1082 1140 1083
rect 1190 1084 1196 1085
rect 1094 1079 1100 1080
rect 1190 1080 1191 1084
rect 1195 1080 1196 1084
rect 1190 1079 1196 1080
rect 1270 1084 1276 1085
rect 1270 1080 1271 1084
rect 1275 1080 1276 1084
rect 1270 1079 1276 1080
rect 1342 1084 1348 1085
rect 1342 1080 1343 1084
rect 1347 1080 1348 1084
rect 1342 1079 1348 1080
rect 1414 1084 1420 1085
rect 1414 1080 1415 1084
rect 1419 1080 1420 1084
rect 1414 1079 1420 1080
rect 1486 1084 1492 1085
rect 1486 1080 1487 1084
rect 1491 1080 1492 1084
rect 1486 1079 1492 1080
rect 1566 1084 1572 1085
rect 1566 1080 1567 1084
rect 1571 1080 1572 1084
rect 1566 1079 1572 1080
rect 1654 1084 1660 1085
rect 1654 1080 1655 1084
rect 1659 1080 1660 1084
rect 1654 1079 1660 1080
rect 1750 1084 1756 1085
rect 1750 1080 1751 1084
rect 1755 1080 1756 1084
rect 1750 1079 1756 1080
rect 1854 1084 1860 1085
rect 1854 1080 1855 1084
rect 1859 1080 1860 1084
rect 1854 1079 1860 1080
rect 1958 1084 1964 1085
rect 1958 1080 1959 1084
rect 1963 1080 1964 1084
rect 1958 1079 1964 1080
rect 2070 1084 2076 1085
rect 2070 1080 2071 1084
rect 2075 1080 2076 1084
rect 2118 1083 2119 1087
rect 2123 1083 2124 1087
rect 2118 1082 2124 1083
rect 2070 1079 2076 1080
rect 158 1076 164 1077
rect 158 1072 159 1076
rect 163 1072 164 1076
rect 158 1071 164 1072
rect 198 1076 204 1077
rect 198 1072 199 1076
rect 203 1072 204 1076
rect 198 1071 204 1072
rect 254 1076 260 1077
rect 254 1072 255 1076
rect 259 1072 260 1076
rect 254 1071 260 1072
rect 318 1076 324 1077
rect 318 1072 319 1076
rect 323 1072 324 1076
rect 318 1071 324 1072
rect 398 1076 404 1077
rect 398 1072 399 1076
rect 403 1072 404 1076
rect 398 1071 404 1072
rect 478 1076 484 1077
rect 478 1072 479 1076
rect 483 1072 484 1076
rect 478 1071 484 1072
rect 558 1076 564 1077
rect 558 1072 559 1076
rect 563 1072 564 1076
rect 558 1071 564 1072
rect 638 1076 644 1077
rect 638 1072 639 1076
rect 643 1072 644 1076
rect 638 1071 644 1072
rect 710 1076 716 1077
rect 710 1072 711 1076
rect 715 1072 716 1076
rect 710 1071 716 1072
rect 782 1076 788 1077
rect 782 1072 783 1076
rect 787 1072 788 1076
rect 782 1071 788 1072
rect 854 1076 860 1077
rect 854 1072 855 1076
rect 859 1072 860 1076
rect 854 1071 860 1072
rect 926 1076 932 1077
rect 926 1072 927 1076
rect 931 1072 932 1076
rect 926 1071 932 1072
rect 998 1076 1004 1077
rect 998 1072 999 1076
rect 1003 1072 1004 1076
rect 998 1071 1004 1072
rect 1046 1076 1052 1077
rect 1046 1072 1047 1076
rect 1051 1072 1052 1076
rect 1046 1071 1052 1072
rect 1158 1072 1164 1073
rect 1134 1069 1140 1070
rect 1134 1065 1135 1069
rect 1139 1065 1140 1069
rect 1158 1068 1159 1072
rect 1163 1068 1164 1072
rect 1158 1067 1164 1068
rect 1198 1072 1204 1073
rect 1198 1068 1199 1072
rect 1203 1068 1204 1072
rect 1198 1067 1204 1068
rect 1246 1072 1252 1073
rect 1246 1068 1247 1072
rect 1251 1068 1252 1072
rect 1246 1067 1252 1068
rect 1302 1072 1308 1073
rect 1302 1068 1303 1072
rect 1307 1068 1308 1072
rect 1302 1067 1308 1068
rect 1350 1072 1356 1073
rect 1350 1068 1351 1072
rect 1355 1068 1356 1072
rect 1350 1067 1356 1068
rect 1398 1072 1404 1073
rect 1398 1068 1399 1072
rect 1403 1068 1404 1072
rect 1398 1067 1404 1068
rect 1454 1072 1460 1073
rect 1454 1068 1455 1072
rect 1459 1068 1460 1072
rect 1454 1067 1460 1068
rect 1510 1072 1516 1073
rect 1510 1068 1511 1072
rect 1515 1068 1516 1072
rect 1510 1067 1516 1068
rect 1582 1072 1588 1073
rect 1582 1068 1583 1072
rect 1587 1068 1588 1072
rect 1582 1067 1588 1068
rect 1662 1072 1668 1073
rect 1662 1068 1663 1072
rect 1667 1068 1668 1072
rect 1662 1067 1668 1068
rect 1758 1072 1764 1073
rect 1758 1068 1759 1072
rect 1763 1068 1764 1072
rect 1758 1067 1764 1068
rect 1862 1072 1868 1073
rect 1862 1068 1863 1072
rect 1867 1068 1868 1072
rect 1862 1067 1868 1068
rect 1966 1072 1972 1073
rect 1966 1068 1967 1072
rect 1971 1068 1972 1072
rect 1966 1067 1972 1068
rect 2070 1072 2076 1073
rect 2070 1068 2071 1072
rect 2075 1068 2076 1072
rect 2070 1067 2076 1068
rect 2118 1069 2124 1070
rect 1134 1064 1140 1065
rect 2118 1065 2119 1069
rect 2123 1065 2124 1069
rect 2118 1064 2124 1065
rect 1134 1052 1140 1053
rect 1134 1048 1135 1052
rect 1139 1048 1140 1052
rect 1134 1047 1140 1048
rect 2118 1052 2124 1053
rect 2118 1048 2119 1052
rect 2123 1048 2124 1052
rect 2118 1047 2124 1048
rect 1158 1044 1164 1045
rect 1158 1040 1159 1044
rect 1163 1040 1164 1044
rect 1158 1039 1164 1040
rect 1198 1044 1204 1045
rect 1198 1040 1199 1044
rect 1203 1040 1204 1044
rect 1198 1039 1204 1040
rect 1246 1044 1252 1045
rect 1246 1040 1247 1044
rect 1251 1040 1252 1044
rect 1246 1039 1252 1040
rect 1302 1044 1308 1045
rect 1302 1040 1303 1044
rect 1307 1040 1308 1044
rect 1302 1039 1308 1040
rect 1350 1044 1356 1045
rect 1350 1040 1351 1044
rect 1355 1040 1356 1044
rect 1350 1039 1356 1040
rect 1398 1044 1404 1045
rect 1398 1040 1399 1044
rect 1403 1040 1404 1044
rect 1398 1039 1404 1040
rect 1454 1044 1460 1045
rect 1454 1040 1455 1044
rect 1459 1040 1460 1044
rect 1454 1039 1460 1040
rect 1510 1044 1516 1045
rect 1510 1040 1511 1044
rect 1515 1040 1516 1044
rect 1510 1039 1516 1040
rect 1582 1044 1588 1045
rect 1582 1040 1583 1044
rect 1587 1040 1588 1044
rect 1582 1039 1588 1040
rect 1662 1044 1668 1045
rect 1662 1040 1663 1044
rect 1667 1040 1668 1044
rect 1662 1039 1668 1040
rect 1758 1044 1764 1045
rect 1758 1040 1759 1044
rect 1763 1040 1764 1044
rect 1758 1039 1764 1040
rect 1862 1044 1868 1045
rect 1862 1040 1863 1044
rect 1867 1040 1868 1044
rect 1862 1039 1868 1040
rect 1966 1044 1972 1045
rect 1966 1040 1967 1044
rect 1971 1040 1972 1044
rect 1966 1039 1972 1040
rect 2070 1044 2076 1045
rect 2070 1040 2071 1044
rect 2075 1040 2076 1044
rect 2070 1039 2076 1040
rect 134 1036 140 1037
rect 134 1032 135 1036
rect 139 1032 140 1036
rect 134 1031 140 1032
rect 174 1036 180 1037
rect 174 1032 175 1036
rect 179 1032 180 1036
rect 174 1031 180 1032
rect 214 1036 220 1037
rect 214 1032 215 1036
rect 219 1032 220 1036
rect 214 1031 220 1032
rect 254 1036 260 1037
rect 254 1032 255 1036
rect 259 1032 260 1036
rect 254 1031 260 1032
rect 318 1036 324 1037
rect 318 1032 319 1036
rect 323 1032 324 1036
rect 318 1031 324 1032
rect 382 1036 388 1037
rect 382 1032 383 1036
rect 387 1032 388 1036
rect 382 1031 388 1032
rect 446 1036 452 1037
rect 446 1032 447 1036
rect 451 1032 452 1036
rect 446 1031 452 1032
rect 510 1036 516 1037
rect 510 1032 511 1036
rect 515 1032 516 1036
rect 510 1031 516 1032
rect 574 1036 580 1037
rect 574 1032 575 1036
rect 579 1032 580 1036
rect 574 1031 580 1032
rect 630 1036 636 1037
rect 630 1032 631 1036
rect 635 1032 636 1036
rect 630 1031 636 1032
rect 686 1036 692 1037
rect 686 1032 687 1036
rect 691 1032 692 1036
rect 686 1031 692 1032
rect 742 1036 748 1037
rect 742 1032 743 1036
rect 747 1032 748 1036
rect 742 1031 748 1032
rect 798 1036 804 1037
rect 798 1032 799 1036
rect 803 1032 804 1036
rect 798 1031 804 1032
rect 862 1036 868 1037
rect 862 1032 863 1036
rect 867 1032 868 1036
rect 862 1031 868 1032
rect 110 1028 116 1029
rect 110 1024 111 1028
rect 115 1024 116 1028
rect 110 1023 116 1024
rect 1094 1028 1100 1029
rect 1094 1024 1095 1028
rect 1099 1024 1100 1028
rect 1094 1023 1100 1024
rect 110 1011 116 1012
rect 110 1007 111 1011
rect 115 1007 116 1011
rect 1094 1011 1100 1012
rect 110 1006 116 1007
rect 134 1008 140 1009
rect 134 1004 135 1008
rect 139 1004 140 1008
rect 134 1003 140 1004
rect 174 1008 180 1009
rect 174 1004 175 1008
rect 179 1004 180 1008
rect 174 1003 180 1004
rect 214 1008 220 1009
rect 214 1004 215 1008
rect 219 1004 220 1008
rect 214 1003 220 1004
rect 254 1008 260 1009
rect 254 1004 255 1008
rect 259 1004 260 1008
rect 254 1003 260 1004
rect 318 1008 324 1009
rect 318 1004 319 1008
rect 323 1004 324 1008
rect 318 1003 324 1004
rect 382 1008 388 1009
rect 382 1004 383 1008
rect 387 1004 388 1008
rect 382 1003 388 1004
rect 446 1008 452 1009
rect 446 1004 447 1008
rect 451 1004 452 1008
rect 446 1003 452 1004
rect 510 1008 516 1009
rect 510 1004 511 1008
rect 515 1004 516 1008
rect 510 1003 516 1004
rect 574 1008 580 1009
rect 574 1004 575 1008
rect 579 1004 580 1008
rect 574 1003 580 1004
rect 630 1008 636 1009
rect 630 1004 631 1008
rect 635 1004 636 1008
rect 630 1003 636 1004
rect 686 1008 692 1009
rect 686 1004 687 1008
rect 691 1004 692 1008
rect 686 1003 692 1004
rect 742 1008 748 1009
rect 742 1004 743 1008
rect 747 1004 748 1008
rect 742 1003 748 1004
rect 798 1008 804 1009
rect 798 1004 799 1008
rect 803 1004 804 1008
rect 798 1003 804 1004
rect 862 1008 868 1009
rect 862 1004 863 1008
rect 867 1004 868 1008
rect 1094 1007 1095 1011
rect 1099 1007 1100 1011
rect 1094 1006 1100 1007
rect 862 1003 868 1004
rect 1158 1004 1164 1005
rect 1158 1000 1159 1004
rect 1163 1000 1164 1004
rect 1158 999 1164 1000
rect 1198 1004 1204 1005
rect 1198 1000 1199 1004
rect 1203 1000 1204 1004
rect 1198 999 1204 1000
rect 1238 1004 1244 1005
rect 1238 1000 1239 1004
rect 1243 1000 1244 1004
rect 1238 999 1244 1000
rect 1294 1004 1300 1005
rect 1294 1000 1295 1004
rect 1299 1000 1300 1004
rect 1294 999 1300 1000
rect 1350 1004 1356 1005
rect 1350 1000 1351 1004
rect 1355 1000 1356 1004
rect 1350 999 1356 1000
rect 1406 1004 1412 1005
rect 1406 1000 1407 1004
rect 1411 1000 1412 1004
rect 1406 999 1412 1000
rect 1462 1004 1468 1005
rect 1462 1000 1463 1004
rect 1467 1000 1468 1004
rect 1462 999 1468 1000
rect 1518 1004 1524 1005
rect 1518 1000 1519 1004
rect 1523 1000 1524 1004
rect 1518 999 1524 1000
rect 1574 1004 1580 1005
rect 1574 1000 1575 1004
rect 1579 1000 1580 1004
rect 1574 999 1580 1000
rect 1638 1004 1644 1005
rect 1638 1000 1639 1004
rect 1643 1000 1644 1004
rect 1638 999 1644 1000
rect 1710 1004 1716 1005
rect 1710 1000 1711 1004
rect 1715 1000 1716 1004
rect 1710 999 1716 1000
rect 1790 1004 1796 1005
rect 1790 1000 1791 1004
rect 1795 1000 1796 1004
rect 1790 999 1796 1000
rect 1878 1004 1884 1005
rect 1878 1000 1879 1004
rect 1883 1000 1884 1004
rect 1878 999 1884 1000
rect 1966 1004 1972 1005
rect 1966 1000 1967 1004
rect 1971 1000 1972 1004
rect 1966 999 1972 1000
rect 2062 1004 2068 1005
rect 2062 1000 2063 1004
rect 2067 1000 2068 1004
rect 2062 999 2068 1000
rect 1134 996 1140 997
rect 134 992 140 993
rect 110 989 116 990
rect 110 985 111 989
rect 115 985 116 989
rect 134 988 135 992
rect 139 988 140 992
rect 134 987 140 988
rect 174 992 180 993
rect 174 988 175 992
rect 179 988 180 992
rect 174 987 180 988
rect 222 992 228 993
rect 222 988 223 992
rect 227 988 228 992
rect 222 987 228 988
rect 278 992 284 993
rect 278 988 279 992
rect 283 988 284 992
rect 278 987 284 988
rect 342 992 348 993
rect 342 988 343 992
rect 347 988 348 992
rect 342 987 348 988
rect 406 992 412 993
rect 406 988 407 992
rect 411 988 412 992
rect 406 987 412 988
rect 470 992 476 993
rect 470 988 471 992
rect 475 988 476 992
rect 470 987 476 988
rect 526 992 532 993
rect 526 988 527 992
rect 531 988 532 992
rect 526 987 532 988
rect 582 992 588 993
rect 582 988 583 992
rect 587 988 588 992
rect 582 987 588 988
rect 630 992 636 993
rect 630 988 631 992
rect 635 988 636 992
rect 630 987 636 988
rect 686 992 692 993
rect 686 988 687 992
rect 691 988 692 992
rect 686 987 692 988
rect 742 992 748 993
rect 742 988 743 992
rect 747 988 748 992
rect 742 987 748 988
rect 798 992 804 993
rect 798 988 799 992
rect 803 988 804 992
rect 1134 992 1135 996
rect 1139 992 1140 996
rect 1134 991 1140 992
rect 2118 996 2124 997
rect 2118 992 2119 996
rect 2123 992 2124 996
rect 2118 991 2124 992
rect 798 987 804 988
rect 1094 989 1100 990
rect 110 984 116 985
rect 1094 985 1095 989
rect 1099 985 1100 989
rect 1094 984 1100 985
rect 1134 979 1140 980
rect 1134 975 1135 979
rect 1139 975 1140 979
rect 2118 979 2124 980
rect 1134 974 1140 975
rect 1158 976 1164 977
rect 110 972 116 973
rect 110 968 111 972
rect 115 968 116 972
rect 110 967 116 968
rect 1094 972 1100 973
rect 1094 968 1095 972
rect 1099 968 1100 972
rect 1158 972 1159 976
rect 1163 972 1164 976
rect 1158 971 1164 972
rect 1198 976 1204 977
rect 1198 972 1199 976
rect 1203 972 1204 976
rect 1198 971 1204 972
rect 1238 976 1244 977
rect 1238 972 1239 976
rect 1243 972 1244 976
rect 1238 971 1244 972
rect 1294 976 1300 977
rect 1294 972 1295 976
rect 1299 972 1300 976
rect 1294 971 1300 972
rect 1350 976 1356 977
rect 1350 972 1351 976
rect 1355 972 1356 976
rect 1350 971 1356 972
rect 1406 976 1412 977
rect 1406 972 1407 976
rect 1411 972 1412 976
rect 1406 971 1412 972
rect 1462 976 1468 977
rect 1462 972 1463 976
rect 1467 972 1468 976
rect 1462 971 1468 972
rect 1518 976 1524 977
rect 1518 972 1519 976
rect 1523 972 1524 976
rect 1518 971 1524 972
rect 1574 976 1580 977
rect 1574 972 1575 976
rect 1579 972 1580 976
rect 1574 971 1580 972
rect 1638 976 1644 977
rect 1638 972 1639 976
rect 1643 972 1644 976
rect 1638 971 1644 972
rect 1710 976 1716 977
rect 1710 972 1711 976
rect 1715 972 1716 976
rect 1710 971 1716 972
rect 1790 976 1796 977
rect 1790 972 1791 976
rect 1795 972 1796 976
rect 1790 971 1796 972
rect 1878 976 1884 977
rect 1878 972 1879 976
rect 1883 972 1884 976
rect 1878 971 1884 972
rect 1966 976 1972 977
rect 1966 972 1967 976
rect 1971 972 1972 976
rect 1966 971 1972 972
rect 2062 976 2068 977
rect 2062 972 2063 976
rect 2067 972 2068 976
rect 2118 975 2119 979
rect 2123 975 2124 979
rect 2118 974 2124 975
rect 2062 971 2068 972
rect 1094 967 1100 968
rect 134 964 140 965
rect 134 960 135 964
rect 139 960 140 964
rect 134 959 140 960
rect 174 964 180 965
rect 174 960 175 964
rect 179 960 180 964
rect 174 959 180 960
rect 222 964 228 965
rect 222 960 223 964
rect 227 960 228 964
rect 222 959 228 960
rect 278 964 284 965
rect 278 960 279 964
rect 283 960 284 964
rect 278 959 284 960
rect 342 964 348 965
rect 342 960 343 964
rect 347 960 348 964
rect 342 959 348 960
rect 406 964 412 965
rect 406 960 407 964
rect 411 960 412 964
rect 406 959 412 960
rect 470 964 476 965
rect 470 960 471 964
rect 475 960 476 964
rect 470 959 476 960
rect 526 964 532 965
rect 526 960 527 964
rect 531 960 532 964
rect 526 959 532 960
rect 582 964 588 965
rect 582 960 583 964
rect 587 960 588 964
rect 582 959 588 960
rect 630 964 636 965
rect 630 960 631 964
rect 635 960 636 964
rect 630 959 636 960
rect 686 964 692 965
rect 686 960 687 964
rect 691 960 692 964
rect 686 959 692 960
rect 742 964 748 965
rect 742 960 743 964
rect 747 960 748 964
rect 742 959 748 960
rect 798 964 804 965
rect 798 960 799 964
rect 803 960 804 964
rect 798 959 804 960
rect 1158 956 1164 957
rect 1134 953 1140 954
rect 1134 949 1135 953
rect 1139 949 1140 953
rect 1158 952 1159 956
rect 1163 952 1164 956
rect 1158 951 1164 952
rect 1206 956 1212 957
rect 1206 952 1207 956
rect 1211 952 1212 956
rect 1206 951 1212 952
rect 1286 956 1292 957
rect 1286 952 1287 956
rect 1291 952 1292 956
rect 1286 951 1292 952
rect 1374 956 1380 957
rect 1374 952 1375 956
rect 1379 952 1380 956
rect 1374 951 1380 952
rect 1454 956 1460 957
rect 1454 952 1455 956
rect 1459 952 1460 956
rect 1454 951 1460 952
rect 1534 956 1540 957
rect 1534 952 1535 956
rect 1539 952 1540 956
rect 1534 951 1540 952
rect 1614 956 1620 957
rect 1614 952 1615 956
rect 1619 952 1620 956
rect 1614 951 1620 952
rect 1686 956 1692 957
rect 1686 952 1687 956
rect 1691 952 1692 956
rect 1686 951 1692 952
rect 1750 956 1756 957
rect 1750 952 1751 956
rect 1755 952 1756 956
rect 1750 951 1756 952
rect 1814 956 1820 957
rect 1814 952 1815 956
rect 1819 952 1820 956
rect 1814 951 1820 952
rect 1878 956 1884 957
rect 1878 952 1879 956
rect 1883 952 1884 956
rect 1878 951 1884 952
rect 1950 956 1956 957
rect 1950 952 1951 956
rect 1955 952 1956 956
rect 1950 951 1956 952
rect 2022 956 2028 957
rect 2022 952 2023 956
rect 2027 952 2028 956
rect 2022 951 2028 952
rect 2070 956 2076 957
rect 2070 952 2071 956
rect 2075 952 2076 956
rect 2070 951 2076 952
rect 2118 953 2124 954
rect 1134 948 1140 949
rect 2118 949 2119 953
rect 2123 949 2124 953
rect 2118 948 2124 949
rect 1134 936 1140 937
rect 1134 932 1135 936
rect 1139 932 1140 936
rect 1134 931 1140 932
rect 2118 936 2124 937
rect 2118 932 2119 936
rect 2123 932 2124 936
rect 2118 931 2124 932
rect 1158 928 1164 929
rect 262 924 268 925
rect 262 920 263 924
rect 267 920 268 924
rect 262 919 268 920
rect 302 924 308 925
rect 302 920 303 924
rect 307 920 308 924
rect 302 919 308 920
rect 350 924 356 925
rect 350 920 351 924
rect 355 920 356 924
rect 350 919 356 920
rect 398 924 404 925
rect 398 920 399 924
rect 403 920 404 924
rect 398 919 404 920
rect 454 924 460 925
rect 454 920 455 924
rect 459 920 460 924
rect 454 919 460 920
rect 510 924 516 925
rect 510 920 511 924
rect 515 920 516 924
rect 510 919 516 920
rect 566 924 572 925
rect 566 920 567 924
rect 571 920 572 924
rect 566 919 572 920
rect 622 924 628 925
rect 622 920 623 924
rect 627 920 628 924
rect 622 919 628 920
rect 686 924 692 925
rect 686 920 687 924
rect 691 920 692 924
rect 686 919 692 920
rect 750 924 756 925
rect 750 920 751 924
rect 755 920 756 924
rect 750 919 756 920
rect 814 924 820 925
rect 814 920 815 924
rect 819 920 820 924
rect 814 919 820 920
rect 878 924 884 925
rect 878 920 879 924
rect 883 920 884 924
rect 878 919 884 920
rect 942 924 948 925
rect 942 920 943 924
rect 947 920 948 924
rect 942 919 948 920
rect 1006 924 1012 925
rect 1006 920 1007 924
rect 1011 920 1012 924
rect 1006 919 1012 920
rect 1046 924 1052 925
rect 1046 920 1047 924
rect 1051 920 1052 924
rect 1158 924 1159 928
rect 1163 924 1164 928
rect 1158 923 1164 924
rect 1206 928 1212 929
rect 1206 924 1207 928
rect 1211 924 1212 928
rect 1206 923 1212 924
rect 1286 928 1292 929
rect 1286 924 1287 928
rect 1291 924 1292 928
rect 1286 923 1292 924
rect 1374 928 1380 929
rect 1374 924 1375 928
rect 1379 924 1380 928
rect 1374 923 1380 924
rect 1454 928 1460 929
rect 1454 924 1455 928
rect 1459 924 1460 928
rect 1454 923 1460 924
rect 1534 928 1540 929
rect 1534 924 1535 928
rect 1539 924 1540 928
rect 1534 923 1540 924
rect 1614 928 1620 929
rect 1614 924 1615 928
rect 1619 924 1620 928
rect 1614 923 1620 924
rect 1686 928 1692 929
rect 1686 924 1687 928
rect 1691 924 1692 928
rect 1686 923 1692 924
rect 1750 928 1756 929
rect 1750 924 1751 928
rect 1755 924 1756 928
rect 1750 923 1756 924
rect 1814 928 1820 929
rect 1814 924 1815 928
rect 1819 924 1820 928
rect 1814 923 1820 924
rect 1878 928 1884 929
rect 1878 924 1879 928
rect 1883 924 1884 928
rect 1878 923 1884 924
rect 1950 928 1956 929
rect 1950 924 1951 928
rect 1955 924 1956 928
rect 1950 923 1956 924
rect 2022 928 2028 929
rect 2022 924 2023 928
rect 2027 924 2028 928
rect 2022 923 2028 924
rect 2070 928 2076 929
rect 2070 924 2071 928
rect 2075 924 2076 928
rect 2070 923 2076 924
rect 1046 919 1052 920
rect 110 916 116 917
rect 110 912 111 916
rect 115 912 116 916
rect 110 911 116 912
rect 1094 916 1100 917
rect 1094 912 1095 916
rect 1099 912 1100 916
rect 1094 911 1100 912
rect 110 899 116 900
rect 110 895 111 899
rect 115 895 116 899
rect 1094 899 1100 900
rect 110 894 116 895
rect 262 896 268 897
rect 262 892 263 896
rect 267 892 268 896
rect 262 891 268 892
rect 302 896 308 897
rect 302 892 303 896
rect 307 892 308 896
rect 302 891 308 892
rect 350 896 356 897
rect 350 892 351 896
rect 355 892 356 896
rect 350 891 356 892
rect 398 896 404 897
rect 398 892 399 896
rect 403 892 404 896
rect 398 891 404 892
rect 454 896 460 897
rect 454 892 455 896
rect 459 892 460 896
rect 454 891 460 892
rect 510 896 516 897
rect 510 892 511 896
rect 515 892 516 896
rect 510 891 516 892
rect 566 896 572 897
rect 566 892 567 896
rect 571 892 572 896
rect 566 891 572 892
rect 622 896 628 897
rect 622 892 623 896
rect 627 892 628 896
rect 622 891 628 892
rect 686 896 692 897
rect 686 892 687 896
rect 691 892 692 896
rect 686 891 692 892
rect 750 896 756 897
rect 750 892 751 896
rect 755 892 756 896
rect 750 891 756 892
rect 814 896 820 897
rect 814 892 815 896
rect 819 892 820 896
rect 814 891 820 892
rect 878 896 884 897
rect 878 892 879 896
rect 883 892 884 896
rect 878 891 884 892
rect 942 896 948 897
rect 942 892 943 896
rect 947 892 948 896
rect 942 891 948 892
rect 1006 896 1012 897
rect 1006 892 1007 896
rect 1011 892 1012 896
rect 1006 891 1012 892
rect 1046 896 1052 897
rect 1046 892 1047 896
rect 1051 892 1052 896
rect 1094 895 1095 899
rect 1099 895 1100 899
rect 1094 894 1100 895
rect 1046 891 1052 892
rect 1238 892 1244 893
rect 1238 888 1239 892
rect 1243 888 1244 892
rect 1238 887 1244 888
rect 1318 892 1324 893
rect 1318 888 1319 892
rect 1323 888 1324 892
rect 1318 887 1324 888
rect 1406 892 1412 893
rect 1406 888 1407 892
rect 1411 888 1412 892
rect 1406 887 1412 888
rect 1494 892 1500 893
rect 1494 888 1495 892
rect 1499 888 1500 892
rect 1494 887 1500 888
rect 1582 892 1588 893
rect 1582 888 1583 892
rect 1587 888 1588 892
rect 1582 887 1588 888
rect 1662 892 1668 893
rect 1662 888 1663 892
rect 1667 888 1668 892
rect 1662 887 1668 888
rect 1742 892 1748 893
rect 1742 888 1743 892
rect 1747 888 1748 892
rect 1742 887 1748 888
rect 1814 892 1820 893
rect 1814 888 1815 892
rect 1819 888 1820 892
rect 1814 887 1820 888
rect 1886 892 1892 893
rect 1886 888 1887 892
rect 1891 888 1892 892
rect 1886 887 1892 888
rect 1950 892 1956 893
rect 1950 888 1951 892
rect 1955 888 1956 892
rect 1950 887 1956 888
rect 2022 892 2028 893
rect 2022 888 2023 892
rect 2027 888 2028 892
rect 2022 887 2028 888
rect 2070 892 2076 893
rect 2070 888 2071 892
rect 2075 888 2076 892
rect 2070 887 2076 888
rect 1134 884 1140 885
rect 302 880 308 881
rect 110 877 116 878
rect 110 873 111 877
rect 115 873 116 877
rect 302 876 303 880
rect 307 876 308 880
rect 302 875 308 876
rect 350 880 356 881
rect 350 876 351 880
rect 355 876 356 880
rect 350 875 356 876
rect 414 880 420 881
rect 414 876 415 880
rect 419 876 420 880
rect 414 875 420 876
rect 478 880 484 881
rect 478 876 479 880
rect 483 876 484 880
rect 478 875 484 876
rect 550 880 556 881
rect 550 876 551 880
rect 555 876 556 880
rect 550 875 556 876
rect 622 880 628 881
rect 622 876 623 880
rect 627 876 628 880
rect 622 875 628 876
rect 694 880 700 881
rect 694 876 695 880
rect 699 876 700 880
rect 694 875 700 876
rect 766 880 772 881
rect 766 876 767 880
rect 771 876 772 880
rect 766 875 772 876
rect 830 880 836 881
rect 830 876 831 880
rect 835 876 836 880
rect 830 875 836 876
rect 886 880 892 881
rect 886 876 887 880
rect 891 876 892 880
rect 886 875 892 876
rect 942 880 948 881
rect 942 876 943 880
rect 947 876 948 880
rect 942 875 948 876
rect 1006 880 1012 881
rect 1006 876 1007 880
rect 1011 876 1012 880
rect 1006 875 1012 876
rect 1046 880 1052 881
rect 1046 876 1047 880
rect 1051 876 1052 880
rect 1134 880 1135 884
rect 1139 880 1140 884
rect 1134 879 1140 880
rect 2118 884 2124 885
rect 2118 880 2119 884
rect 2123 880 2124 884
rect 2118 879 2124 880
rect 1046 875 1052 876
rect 1094 877 1100 878
rect 110 872 116 873
rect 1094 873 1095 877
rect 1099 873 1100 877
rect 1094 872 1100 873
rect 1134 867 1140 868
rect 1134 863 1135 867
rect 1139 863 1140 867
rect 2118 867 2124 868
rect 1134 862 1140 863
rect 1238 864 1244 865
rect 110 860 116 861
rect 110 856 111 860
rect 115 856 116 860
rect 110 855 116 856
rect 1094 860 1100 861
rect 1094 856 1095 860
rect 1099 856 1100 860
rect 1238 860 1239 864
rect 1243 860 1244 864
rect 1238 859 1244 860
rect 1318 864 1324 865
rect 1318 860 1319 864
rect 1323 860 1324 864
rect 1318 859 1324 860
rect 1406 864 1412 865
rect 1406 860 1407 864
rect 1411 860 1412 864
rect 1406 859 1412 860
rect 1494 864 1500 865
rect 1494 860 1495 864
rect 1499 860 1500 864
rect 1494 859 1500 860
rect 1582 864 1588 865
rect 1582 860 1583 864
rect 1587 860 1588 864
rect 1582 859 1588 860
rect 1662 864 1668 865
rect 1662 860 1663 864
rect 1667 860 1668 864
rect 1662 859 1668 860
rect 1742 864 1748 865
rect 1742 860 1743 864
rect 1747 860 1748 864
rect 1742 859 1748 860
rect 1814 864 1820 865
rect 1814 860 1815 864
rect 1819 860 1820 864
rect 1814 859 1820 860
rect 1886 864 1892 865
rect 1886 860 1887 864
rect 1891 860 1892 864
rect 1886 859 1892 860
rect 1950 864 1956 865
rect 1950 860 1951 864
rect 1955 860 1956 864
rect 1950 859 1956 860
rect 2022 864 2028 865
rect 2022 860 2023 864
rect 2027 860 2028 864
rect 2022 859 2028 860
rect 2070 864 2076 865
rect 2070 860 2071 864
rect 2075 860 2076 864
rect 2118 863 2119 867
rect 2123 863 2124 867
rect 2118 862 2124 863
rect 2070 859 2076 860
rect 1094 855 1100 856
rect 302 852 308 853
rect 302 848 303 852
rect 307 848 308 852
rect 302 847 308 848
rect 350 852 356 853
rect 350 848 351 852
rect 355 848 356 852
rect 350 847 356 848
rect 414 852 420 853
rect 414 848 415 852
rect 419 848 420 852
rect 414 847 420 848
rect 478 852 484 853
rect 478 848 479 852
rect 483 848 484 852
rect 478 847 484 848
rect 550 852 556 853
rect 550 848 551 852
rect 555 848 556 852
rect 550 847 556 848
rect 622 852 628 853
rect 622 848 623 852
rect 627 848 628 852
rect 622 847 628 848
rect 694 852 700 853
rect 694 848 695 852
rect 699 848 700 852
rect 694 847 700 848
rect 766 852 772 853
rect 766 848 767 852
rect 771 848 772 852
rect 766 847 772 848
rect 830 852 836 853
rect 830 848 831 852
rect 835 848 836 852
rect 830 847 836 848
rect 886 852 892 853
rect 886 848 887 852
rect 891 848 892 852
rect 886 847 892 848
rect 942 852 948 853
rect 942 848 943 852
rect 947 848 948 852
rect 942 847 948 848
rect 1006 852 1012 853
rect 1006 848 1007 852
rect 1011 848 1012 852
rect 1006 847 1012 848
rect 1046 852 1052 853
rect 1046 848 1047 852
rect 1051 848 1052 852
rect 1158 852 1164 853
rect 1046 847 1052 848
rect 1134 849 1140 850
rect 1134 845 1135 849
rect 1139 845 1140 849
rect 1158 848 1159 852
rect 1163 848 1164 852
rect 1158 847 1164 848
rect 1246 852 1252 853
rect 1246 848 1247 852
rect 1251 848 1252 852
rect 1246 847 1252 848
rect 1358 852 1364 853
rect 1358 848 1359 852
rect 1363 848 1364 852
rect 1358 847 1364 848
rect 1454 852 1460 853
rect 1454 848 1455 852
rect 1459 848 1460 852
rect 1454 847 1460 848
rect 1542 852 1548 853
rect 1542 848 1543 852
rect 1547 848 1548 852
rect 1542 847 1548 848
rect 1630 852 1636 853
rect 1630 848 1631 852
rect 1635 848 1636 852
rect 1630 847 1636 848
rect 1710 852 1716 853
rect 1710 848 1711 852
rect 1715 848 1716 852
rect 1710 847 1716 848
rect 1782 852 1788 853
rect 1782 848 1783 852
rect 1787 848 1788 852
rect 1782 847 1788 848
rect 1854 852 1860 853
rect 1854 848 1855 852
rect 1859 848 1860 852
rect 1854 847 1860 848
rect 1934 852 1940 853
rect 1934 848 1935 852
rect 1939 848 1940 852
rect 1934 847 1940 848
rect 2014 852 2020 853
rect 2014 848 2015 852
rect 2019 848 2020 852
rect 2014 847 2020 848
rect 2070 852 2076 853
rect 2070 848 2071 852
rect 2075 848 2076 852
rect 2070 847 2076 848
rect 2118 849 2124 850
rect 1134 844 1140 845
rect 2118 845 2119 849
rect 2123 845 2124 849
rect 2118 844 2124 845
rect 1134 832 1140 833
rect 1134 828 1135 832
rect 1139 828 1140 832
rect 1134 827 1140 828
rect 2118 832 2124 833
rect 2118 828 2119 832
rect 2123 828 2124 832
rect 2118 827 2124 828
rect 1158 824 1164 825
rect 1158 820 1159 824
rect 1163 820 1164 824
rect 1158 819 1164 820
rect 1246 824 1252 825
rect 1246 820 1247 824
rect 1251 820 1252 824
rect 1246 819 1252 820
rect 1358 824 1364 825
rect 1358 820 1359 824
rect 1363 820 1364 824
rect 1358 819 1364 820
rect 1454 824 1460 825
rect 1454 820 1455 824
rect 1459 820 1460 824
rect 1454 819 1460 820
rect 1542 824 1548 825
rect 1542 820 1543 824
rect 1547 820 1548 824
rect 1542 819 1548 820
rect 1630 824 1636 825
rect 1630 820 1631 824
rect 1635 820 1636 824
rect 1630 819 1636 820
rect 1710 824 1716 825
rect 1710 820 1711 824
rect 1715 820 1716 824
rect 1710 819 1716 820
rect 1782 824 1788 825
rect 1782 820 1783 824
rect 1787 820 1788 824
rect 1782 819 1788 820
rect 1854 824 1860 825
rect 1854 820 1855 824
rect 1859 820 1860 824
rect 1854 819 1860 820
rect 1934 824 1940 825
rect 1934 820 1935 824
rect 1939 820 1940 824
rect 1934 819 1940 820
rect 2014 824 2020 825
rect 2014 820 2015 824
rect 2019 820 2020 824
rect 2014 819 2020 820
rect 2070 824 2076 825
rect 2070 820 2071 824
rect 2075 820 2076 824
rect 2070 819 2076 820
rect 278 816 284 817
rect 278 812 279 816
rect 283 812 284 816
rect 278 811 284 812
rect 342 816 348 817
rect 342 812 343 816
rect 347 812 348 816
rect 342 811 348 812
rect 414 816 420 817
rect 414 812 415 816
rect 419 812 420 816
rect 414 811 420 812
rect 486 816 492 817
rect 486 812 487 816
rect 491 812 492 816
rect 486 811 492 812
rect 566 816 572 817
rect 566 812 567 816
rect 571 812 572 816
rect 566 811 572 812
rect 646 816 652 817
rect 646 812 647 816
rect 651 812 652 816
rect 646 811 652 812
rect 726 816 732 817
rect 726 812 727 816
rect 731 812 732 816
rect 726 811 732 812
rect 798 816 804 817
rect 798 812 799 816
rect 803 812 804 816
rect 798 811 804 812
rect 862 816 868 817
rect 862 812 863 816
rect 867 812 868 816
rect 862 811 868 812
rect 926 816 932 817
rect 926 812 927 816
rect 931 812 932 816
rect 926 811 932 812
rect 998 816 1004 817
rect 998 812 999 816
rect 1003 812 1004 816
rect 998 811 1004 812
rect 1046 816 1052 817
rect 1046 812 1047 816
rect 1051 812 1052 816
rect 1046 811 1052 812
rect 110 808 116 809
rect 110 804 111 808
rect 115 804 116 808
rect 110 803 116 804
rect 1094 808 1100 809
rect 1094 804 1095 808
rect 1099 804 1100 808
rect 1094 803 1100 804
rect 110 791 116 792
rect 110 787 111 791
rect 115 787 116 791
rect 1094 791 1100 792
rect 110 786 116 787
rect 278 788 284 789
rect 278 784 279 788
rect 283 784 284 788
rect 278 783 284 784
rect 342 788 348 789
rect 342 784 343 788
rect 347 784 348 788
rect 342 783 348 784
rect 414 788 420 789
rect 414 784 415 788
rect 419 784 420 788
rect 414 783 420 784
rect 486 788 492 789
rect 486 784 487 788
rect 491 784 492 788
rect 486 783 492 784
rect 566 788 572 789
rect 566 784 567 788
rect 571 784 572 788
rect 566 783 572 784
rect 646 788 652 789
rect 646 784 647 788
rect 651 784 652 788
rect 646 783 652 784
rect 726 788 732 789
rect 726 784 727 788
rect 731 784 732 788
rect 726 783 732 784
rect 798 788 804 789
rect 798 784 799 788
rect 803 784 804 788
rect 798 783 804 784
rect 862 788 868 789
rect 862 784 863 788
rect 867 784 868 788
rect 862 783 868 784
rect 926 788 932 789
rect 926 784 927 788
rect 931 784 932 788
rect 926 783 932 784
rect 998 788 1004 789
rect 998 784 999 788
rect 1003 784 1004 788
rect 998 783 1004 784
rect 1046 788 1052 789
rect 1046 784 1047 788
rect 1051 784 1052 788
rect 1094 787 1095 791
rect 1099 787 1100 791
rect 1094 786 1100 787
rect 1158 788 1164 789
rect 1046 783 1052 784
rect 1158 784 1159 788
rect 1163 784 1164 788
rect 1158 783 1164 784
rect 1278 788 1284 789
rect 1278 784 1279 788
rect 1283 784 1284 788
rect 1278 783 1284 784
rect 1406 788 1412 789
rect 1406 784 1407 788
rect 1411 784 1412 788
rect 1406 783 1412 784
rect 1518 788 1524 789
rect 1518 784 1519 788
rect 1523 784 1524 788
rect 1518 783 1524 784
rect 1622 788 1628 789
rect 1622 784 1623 788
rect 1627 784 1628 788
rect 1622 783 1628 784
rect 1718 788 1724 789
rect 1718 784 1719 788
rect 1723 784 1724 788
rect 1718 783 1724 784
rect 1814 788 1820 789
rect 1814 784 1815 788
rect 1819 784 1820 788
rect 1814 783 1820 784
rect 1902 788 1908 789
rect 1902 784 1903 788
rect 1907 784 1908 788
rect 1902 783 1908 784
rect 1998 788 2004 789
rect 1998 784 1999 788
rect 2003 784 2004 788
rect 1998 783 2004 784
rect 2070 788 2076 789
rect 2070 784 2071 788
rect 2075 784 2076 788
rect 2070 783 2076 784
rect 1134 780 1140 781
rect 214 776 220 777
rect 110 773 116 774
rect 110 769 111 773
rect 115 769 116 773
rect 214 772 215 776
rect 219 772 220 776
rect 214 771 220 772
rect 278 776 284 777
rect 278 772 279 776
rect 283 772 284 776
rect 278 771 284 772
rect 350 776 356 777
rect 350 772 351 776
rect 355 772 356 776
rect 350 771 356 772
rect 422 776 428 777
rect 422 772 423 776
rect 427 772 428 776
rect 422 771 428 772
rect 494 776 500 777
rect 494 772 495 776
rect 499 772 500 776
rect 494 771 500 772
rect 566 776 572 777
rect 566 772 567 776
rect 571 772 572 776
rect 566 771 572 772
rect 638 776 644 777
rect 638 772 639 776
rect 643 772 644 776
rect 638 771 644 772
rect 702 776 708 777
rect 702 772 703 776
rect 707 772 708 776
rect 702 771 708 772
rect 758 776 764 777
rect 758 772 759 776
rect 763 772 764 776
rect 758 771 764 772
rect 814 776 820 777
rect 814 772 815 776
rect 819 772 820 776
rect 814 771 820 772
rect 862 776 868 777
rect 862 772 863 776
rect 867 772 868 776
rect 862 771 868 772
rect 910 776 916 777
rect 910 772 911 776
rect 915 772 916 776
rect 910 771 916 772
rect 958 776 964 777
rect 958 772 959 776
rect 963 772 964 776
rect 958 771 964 772
rect 1006 776 1012 777
rect 1006 772 1007 776
rect 1011 772 1012 776
rect 1006 771 1012 772
rect 1046 776 1052 777
rect 1046 772 1047 776
rect 1051 772 1052 776
rect 1134 776 1135 780
rect 1139 776 1140 780
rect 1134 775 1140 776
rect 2118 780 2124 781
rect 2118 776 2119 780
rect 2123 776 2124 780
rect 2118 775 2124 776
rect 1046 771 1052 772
rect 1094 773 1100 774
rect 110 768 116 769
rect 1094 769 1095 773
rect 1099 769 1100 773
rect 1094 768 1100 769
rect 1134 763 1140 764
rect 1134 759 1135 763
rect 1139 759 1140 763
rect 2118 763 2124 764
rect 1134 758 1140 759
rect 1158 760 1164 761
rect 110 756 116 757
rect 110 752 111 756
rect 115 752 116 756
rect 110 751 116 752
rect 1094 756 1100 757
rect 1094 752 1095 756
rect 1099 752 1100 756
rect 1158 756 1159 760
rect 1163 756 1164 760
rect 1158 755 1164 756
rect 1278 760 1284 761
rect 1278 756 1279 760
rect 1283 756 1284 760
rect 1278 755 1284 756
rect 1406 760 1412 761
rect 1406 756 1407 760
rect 1411 756 1412 760
rect 1406 755 1412 756
rect 1518 760 1524 761
rect 1518 756 1519 760
rect 1523 756 1524 760
rect 1518 755 1524 756
rect 1622 760 1628 761
rect 1622 756 1623 760
rect 1627 756 1628 760
rect 1622 755 1628 756
rect 1718 760 1724 761
rect 1718 756 1719 760
rect 1723 756 1724 760
rect 1718 755 1724 756
rect 1814 760 1820 761
rect 1814 756 1815 760
rect 1819 756 1820 760
rect 1814 755 1820 756
rect 1902 760 1908 761
rect 1902 756 1903 760
rect 1907 756 1908 760
rect 1902 755 1908 756
rect 1998 760 2004 761
rect 1998 756 1999 760
rect 2003 756 2004 760
rect 1998 755 2004 756
rect 2070 760 2076 761
rect 2070 756 2071 760
rect 2075 756 2076 760
rect 2118 759 2119 763
rect 2123 759 2124 763
rect 2118 758 2124 759
rect 2070 755 2076 756
rect 1094 751 1100 752
rect 214 748 220 749
rect 214 744 215 748
rect 219 744 220 748
rect 214 743 220 744
rect 278 748 284 749
rect 278 744 279 748
rect 283 744 284 748
rect 278 743 284 744
rect 350 748 356 749
rect 350 744 351 748
rect 355 744 356 748
rect 350 743 356 744
rect 422 748 428 749
rect 422 744 423 748
rect 427 744 428 748
rect 422 743 428 744
rect 494 748 500 749
rect 494 744 495 748
rect 499 744 500 748
rect 494 743 500 744
rect 566 748 572 749
rect 566 744 567 748
rect 571 744 572 748
rect 566 743 572 744
rect 638 748 644 749
rect 638 744 639 748
rect 643 744 644 748
rect 638 743 644 744
rect 702 748 708 749
rect 702 744 703 748
rect 707 744 708 748
rect 702 743 708 744
rect 758 748 764 749
rect 758 744 759 748
rect 763 744 764 748
rect 758 743 764 744
rect 814 748 820 749
rect 814 744 815 748
rect 819 744 820 748
rect 814 743 820 744
rect 862 748 868 749
rect 862 744 863 748
rect 867 744 868 748
rect 862 743 868 744
rect 910 748 916 749
rect 910 744 911 748
rect 915 744 916 748
rect 910 743 916 744
rect 958 748 964 749
rect 958 744 959 748
rect 963 744 964 748
rect 958 743 964 744
rect 1006 748 1012 749
rect 1006 744 1007 748
rect 1011 744 1012 748
rect 1006 743 1012 744
rect 1046 748 1052 749
rect 1046 744 1047 748
rect 1051 744 1052 748
rect 1046 743 1052 744
rect 1334 744 1340 745
rect 1134 741 1140 742
rect 1134 737 1135 741
rect 1139 737 1140 741
rect 1334 740 1335 744
rect 1339 740 1340 744
rect 1334 739 1340 740
rect 1374 744 1380 745
rect 1374 740 1375 744
rect 1379 740 1380 744
rect 1374 739 1380 740
rect 1414 744 1420 745
rect 1414 740 1415 744
rect 1419 740 1420 744
rect 1414 739 1420 740
rect 1454 744 1460 745
rect 1454 740 1455 744
rect 1459 740 1460 744
rect 1454 739 1460 740
rect 1502 744 1508 745
rect 1502 740 1503 744
rect 1507 740 1508 744
rect 1502 739 1508 740
rect 1550 744 1556 745
rect 1550 740 1551 744
rect 1555 740 1556 744
rect 1550 739 1556 740
rect 1598 744 1604 745
rect 1598 740 1599 744
rect 1603 740 1604 744
rect 1598 739 1604 740
rect 1654 744 1660 745
rect 1654 740 1655 744
rect 1659 740 1660 744
rect 1654 739 1660 740
rect 1710 744 1716 745
rect 1710 740 1711 744
rect 1715 740 1716 744
rect 1710 739 1716 740
rect 1766 744 1772 745
rect 1766 740 1767 744
rect 1771 740 1772 744
rect 1766 739 1772 740
rect 1830 744 1836 745
rect 1830 740 1831 744
rect 1835 740 1836 744
rect 1830 739 1836 740
rect 1894 744 1900 745
rect 1894 740 1895 744
rect 1899 740 1900 744
rect 1894 739 1900 740
rect 1958 744 1964 745
rect 1958 740 1959 744
rect 1963 740 1964 744
rect 1958 739 1964 740
rect 2022 744 2028 745
rect 2022 740 2023 744
rect 2027 740 2028 744
rect 2022 739 2028 740
rect 2070 744 2076 745
rect 2070 740 2071 744
rect 2075 740 2076 744
rect 2070 739 2076 740
rect 2118 741 2124 742
rect 1134 736 1140 737
rect 2118 737 2119 741
rect 2123 737 2124 741
rect 2118 736 2124 737
rect 1134 724 1140 725
rect 1134 720 1135 724
rect 1139 720 1140 724
rect 1134 719 1140 720
rect 2118 724 2124 725
rect 2118 720 2119 724
rect 2123 720 2124 724
rect 2118 719 2124 720
rect 1334 716 1340 717
rect 174 712 180 713
rect 174 708 175 712
rect 179 708 180 712
rect 174 707 180 708
rect 238 712 244 713
rect 238 708 239 712
rect 243 708 244 712
rect 238 707 244 708
rect 310 712 316 713
rect 310 708 311 712
rect 315 708 316 712
rect 310 707 316 708
rect 390 712 396 713
rect 390 708 391 712
rect 395 708 396 712
rect 390 707 396 708
rect 470 712 476 713
rect 470 708 471 712
rect 475 708 476 712
rect 470 707 476 708
rect 542 712 548 713
rect 542 708 543 712
rect 547 708 548 712
rect 542 707 548 708
rect 614 712 620 713
rect 614 708 615 712
rect 619 708 620 712
rect 614 707 620 708
rect 678 712 684 713
rect 678 708 679 712
rect 683 708 684 712
rect 678 707 684 708
rect 734 712 740 713
rect 734 708 735 712
rect 739 708 740 712
rect 734 707 740 708
rect 798 712 804 713
rect 798 708 799 712
rect 803 708 804 712
rect 798 707 804 708
rect 862 712 868 713
rect 862 708 863 712
rect 867 708 868 712
rect 862 707 868 708
rect 926 712 932 713
rect 926 708 927 712
rect 931 708 932 712
rect 1334 712 1335 716
rect 1339 712 1340 716
rect 1334 711 1340 712
rect 1374 716 1380 717
rect 1374 712 1375 716
rect 1379 712 1380 716
rect 1374 711 1380 712
rect 1414 716 1420 717
rect 1414 712 1415 716
rect 1419 712 1420 716
rect 1414 711 1420 712
rect 1454 716 1460 717
rect 1454 712 1455 716
rect 1459 712 1460 716
rect 1454 711 1460 712
rect 1502 716 1508 717
rect 1502 712 1503 716
rect 1507 712 1508 716
rect 1502 711 1508 712
rect 1550 716 1556 717
rect 1550 712 1551 716
rect 1555 712 1556 716
rect 1550 711 1556 712
rect 1598 716 1604 717
rect 1598 712 1599 716
rect 1603 712 1604 716
rect 1598 711 1604 712
rect 1654 716 1660 717
rect 1654 712 1655 716
rect 1659 712 1660 716
rect 1654 711 1660 712
rect 1710 716 1716 717
rect 1710 712 1711 716
rect 1715 712 1716 716
rect 1710 711 1716 712
rect 1766 716 1772 717
rect 1766 712 1767 716
rect 1771 712 1772 716
rect 1766 711 1772 712
rect 1830 716 1836 717
rect 1830 712 1831 716
rect 1835 712 1836 716
rect 1830 711 1836 712
rect 1894 716 1900 717
rect 1894 712 1895 716
rect 1899 712 1900 716
rect 1894 711 1900 712
rect 1958 716 1964 717
rect 1958 712 1959 716
rect 1963 712 1964 716
rect 1958 711 1964 712
rect 2022 716 2028 717
rect 2022 712 2023 716
rect 2027 712 2028 716
rect 2022 711 2028 712
rect 2070 716 2076 717
rect 2070 712 2071 716
rect 2075 712 2076 716
rect 2070 711 2076 712
rect 926 707 932 708
rect 110 704 116 705
rect 110 700 111 704
rect 115 700 116 704
rect 110 699 116 700
rect 1094 704 1100 705
rect 1094 700 1095 704
rect 1099 700 1100 704
rect 1094 699 1100 700
rect 110 687 116 688
rect 110 683 111 687
rect 115 683 116 687
rect 1094 687 1100 688
rect 110 682 116 683
rect 174 684 180 685
rect 174 680 175 684
rect 179 680 180 684
rect 174 679 180 680
rect 238 684 244 685
rect 238 680 239 684
rect 243 680 244 684
rect 238 679 244 680
rect 310 684 316 685
rect 310 680 311 684
rect 315 680 316 684
rect 310 679 316 680
rect 390 684 396 685
rect 390 680 391 684
rect 395 680 396 684
rect 390 679 396 680
rect 470 684 476 685
rect 470 680 471 684
rect 475 680 476 684
rect 470 679 476 680
rect 542 684 548 685
rect 542 680 543 684
rect 547 680 548 684
rect 542 679 548 680
rect 614 684 620 685
rect 614 680 615 684
rect 619 680 620 684
rect 614 679 620 680
rect 678 684 684 685
rect 678 680 679 684
rect 683 680 684 684
rect 678 679 684 680
rect 734 684 740 685
rect 734 680 735 684
rect 739 680 740 684
rect 734 679 740 680
rect 798 684 804 685
rect 798 680 799 684
rect 803 680 804 684
rect 798 679 804 680
rect 862 684 868 685
rect 862 680 863 684
rect 867 680 868 684
rect 862 679 868 680
rect 926 684 932 685
rect 926 680 927 684
rect 931 680 932 684
rect 1094 683 1095 687
rect 1099 683 1100 687
rect 1094 682 1100 683
rect 926 679 932 680
rect 1246 680 1252 681
rect 1246 676 1247 680
rect 1251 676 1252 680
rect 1246 675 1252 676
rect 1286 680 1292 681
rect 1286 676 1287 680
rect 1291 676 1292 680
rect 1286 675 1292 676
rect 1334 680 1340 681
rect 1334 676 1335 680
rect 1339 676 1340 680
rect 1334 675 1340 676
rect 1390 680 1396 681
rect 1390 676 1391 680
rect 1395 676 1396 680
rect 1390 675 1396 676
rect 1446 680 1452 681
rect 1446 676 1447 680
rect 1451 676 1452 680
rect 1446 675 1452 676
rect 1510 680 1516 681
rect 1510 676 1511 680
rect 1515 676 1516 680
rect 1510 675 1516 676
rect 1582 680 1588 681
rect 1582 676 1583 680
rect 1587 676 1588 680
rect 1582 675 1588 676
rect 1654 680 1660 681
rect 1654 676 1655 680
rect 1659 676 1660 680
rect 1654 675 1660 676
rect 1734 680 1740 681
rect 1734 676 1735 680
rect 1739 676 1740 680
rect 1734 675 1740 676
rect 1822 680 1828 681
rect 1822 676 1823 680
rect 1827 676 1828 680
rect 1822 675 1828 676
rect 1910 680 1916 681
rect 1910 676 1911 680
rect 1915 676 1916 680
rect 1910 675 1916 676
rect 1998 680 2004 681
rect 1998 676 1999 680
rect 2003 676 2004 680
rect 1998 675 2004 676
rect 2070 680 2076 681
rect 2070 676 2071 680
rect 2075 676 2076 680
rect 2070 675 2076 676
rect 134 672 140 673
rect 110 669 116 670
rect 110 665 111 669
rect 115 665 116 669
rect 134 668 135 672
rect 139 668 140 672
rect 134 667 140 668
rect 174 672 180 673
rect 174 668 175 672
rect 179 668 180 672
rect 174 667 180 668
rect 214 672 220 673
rect 214 668 215 672
rect 219 668 220 672
rect 214 667 220 668
rect 270 672 276 673
rect 270 668 271 672
rect 275 668 276 672
rect 270 667 276 668
rect 334 672 340 673
rect 334 668 335 672
rect 339 668 340 672
rect 334 667 340 668
rect 398 672 404 673
rect 398 668 399 672
rect 403 668 404 672
rect 398 667 404 668
rect 462 672 468 673
rect 462 668 463 672
rect 467 668 468 672
rect 462 667 468 668
rect 526 672 532 673
rect 526 668 527 672
rect 531 668 532 672
rect 526 667 532 668
rect 590 672 596 673
rect 590 668 591 672
rect 595 668 596 672
rect 590 667 596 668
rect 646 672 652 673
rect 646 668 647 672
rect 651 668 652 672
rect 646 667 652 668
rect 702 672 708 673
rect 702 668 703 672
rect 707 668 708 672
rect 702 667 708 668
rect 758 672 764 673
rect 758 668 759 672
rect 763 668 764 672
rect 758 667 764 668
rect 822 672 828 673
rect 822 668 823 672
rect 827 668 828 672
rect 1134 672 1140 673
rect 822 667 828 668
rect 1094 669 1100 670
rect 110 664 116 665
rect 1094 665 1095 669
rect 1099 665 1100 669
rect 1134 668 1135 672
rect 1139 668 1140 672
rect 1134 667 1140 668
rect 2118 672 2124 673
rect 2118 668 2119 672
rect 2123 668 2124 672
rect 2118 667 2124 668
rect 1094 664 1100 665
rect 1134 655 1140 656
rect 110 652 116 653
rect 110 648 111 652
rect 115 648 116 652
rect 110 647 116 648
rect 1094 652 1100 653
rect 1094 648 1095 652
rect 1099 648 1100 652
rect 1134 651 1135 655
rect 1139 651 1140 655
rect 2118 655 2124 656
rect 1134 650 1140 651
rect 1246 652 1252 653
rect 1094 647 1100 648
rect 1246 648 1247 652
rect 1251 648 1252 652
rect 1246 647 1252 648
rect 1286 652 1292 653
rect 1286 648 1287 652
rect 1291 648 1292 652
rect 1286 647 1292 648
rect 1334 652 1340 653
rect 1334 648 1335 652
rect 1339 648 1340 652
rect 1334 647 1340 648
rect 1390 652 1396 653
rect 1390 648 1391 652
rect 1395 648 1396 652
rect 1390 647 1396 648
rect 1446 652 1452 653
rect 1446 648 1447 652
rect 1451 648 1452 652
rect 1446 647 1452 648
rect 1510 652 1516 653
rect 1510 648 1511 652
rect 1515 648 1516 652
rect 1510 647 1516 648
rect 1582 652 1588 653
rect 1582 648 1583 652
rect 1587 648 1588 652
rect 1582 647 1588 648
rect 1654 652 1660 653
rect 1654 648 1655 652
rect 1659 648 1660 652
rect 1654 647 1660 648
rect 1734 652 1740 653
rect 1734 648 1735 652
rect 1739 648 1740 652
rect 1734 647 1740 648
rect 1822 652 1828 653
rect 1822 648 1823 652
rect 1827 648 1828 652
rect 1822 647 1828 648
rect 1910 652 1916 653
rect 1910 648 1911 652
rect 1915 648 1916 652
rect 1910 647 1916 648
rect 1998 652 2004 653
rect 1998 648 1999 652
rect 2003 648 2004 652
rect 1998 647 2004 648
rect 2070 652 2076 653
rect 2070 648 2071 652
rect 2075 648 2076 652
rect 2118 651 2119 655
rect 2123 651 2124 655
rect 2118 650 2124 651
rect 2070 647 2076 648
rect 134 644 140 645
rect 134 640 135 644
rect 139 640 140 644
rect 134 639 140 640
rect 174 644 180 645
rect 174 640 175 644
rect 179 640 180 644
rect 174 639 180 640
rect 214 644 220 645
rect 214 640 215 644
rect 219 640 220 644
rect 214 639 220 640
rect 270 644 276 645
rect 270 640 271 644
rect 275 640 276 644
rect 270 639 276 640
rect 334 644 340 645
rect 334 640 335 644
rect 339 640 340 644
rect 334 639 340 640
rect 398 644 404 645
rect 398 640 399 644
rect 403 640 404 644
rect 398 639 404 640
rect 462 644 468 645
rect 462 640 463 644
rect 467 640 468 644
rect 462 639 468 640
rect 526 644 532 645
rect 526 640 527 644
rect 531 640 532 644
rect 526 639 532 640
rect 590 644 596 645
rect 590 640 591 644
rect 595 640 596 644
rect 590 639 596 640
rect 646 644 652 645
rect 646 640 647 644
rect 651 640 652 644
rect 646 639 652 640
rect 702 644 708 645
rect 702 640 703 644
rect 707 640 708 644
rect 702 639 708 640
rect 758 644 764 645
rect 758 640 759 644
rect 763 640 764 644
rect 758 639 764 640
rect 822 644 828 645
rect 822 640 823 644
rect 827 640 828 644
rect 822 639 828 640
rect 1158 640 1164 641
rect 1134 637 1140 638
rect 1134 633 1135 637
rect 1139 633 1140 637
rect 1158 636 1159 640
rect 1163 636 1164 640
rect 1158 635 1164 636
rect 1198 640 1204 641
rect 1198 636 1199 640
rect 1203 636 1204 640
rect 1198 635 1204 636
rect 1238 640 1244 641
rect 1238 636 1239 640
rect 1243 636 1244 640
rect 1238 635 1244 636
rect 1278 640 1284 641
rect 1278 636 1279 640
rect 1283 636 1284 640
rect 1278 635 1284 636
rect 1342 640 1348 641
rect 1342 636 1343 640
rect 1347 636 1348 640
rect 1342 635 1348 636
rect 1414 640 1420 641
rect 1414 636 1415 640
rect 1419 636 1420 640
rect 1414 635 1420 636
rect 1494 640 1500 641
rect 1494 636 1495 640
rect 1499 636 1500 640
rect 1494 635 1500 636
rect 1582 640 1588 641
rect 1582 636 1583 640
rect 1587 636 1588 640
rect 1582 635 1588 636
rect 1670 640 1676 641
rect 1670 636 1671 640
rect 1675 636 1676 640
rect 1670 635 1676 636
rect 1758 640 1764 641
rect 1758 636 1759 640
rect 1763 636 1764 640
rect 1758 635 1764 636
rect 1838 640 1844 641
rect 1838 636 1839 640
rect 1843 636 1844 640
rect 1838 635 1844 636
rect 1918 640 1924 641
rect 1918 636 1919 640
rect 1923 636 1924 640
rect 1918 635 1924 636
rect 2006 640 2012 641
rect 2006 636 2007 640
rect 2011 636 2012 640
rect 2006 635 2012 636
rect 2070 640 2076 641
rect 2070 636 2071 640
rect 2075 636 2076 640
rect 2070 635 2076 636
rect 2118 637 2124 638
rect 1134 632 1140 633
rect 2118 633 2119 637
rect 2123 633 2124 637
rect 2118 632 2124 633
rect 1134 620 1140 621
rect 1134 616 1135 620
rect 1139 616 1140 620
rect 1134 615 1140 616
rect 2118 620 2124 621
rect 2118 616 2119 620
rect 2123 616 2124 620
rect 2118 615 2124 616
rect 1158 612 1164 613
rect 1158 608 1159 612
rect 1163 608 1164 612
rect 1158 607 1164 608
rect 1198 612 1204 613
rect 1198 608 1199 612
rect 1203 608 1204 612
rect 1198 607 1204 608
rect 1238 612 1244 613
rect 1238 608 1239 612
rect 1243 608 1244 612
rect 1238 607 1244 608
rect 1278 612 1284 613
rect 1278 608 1279 612
rect 1283 608 1284 612
rect 1278 607 1284 608
rect 1342 612 1348 613
rect 1342 608 1343 612
rect 1347 608 1348 612
rect 1342 607 1348 608
rect 1414 612 1420 613
rect 1414 608 1415 612
rect 1419 608 1420 612
rect 1414 607 1420 608
rect 1494 612 1500 613
rect 1494 608 1495 612
rect 1499 608 1500 612
rect 1494 607 1500 608
rect 1582 612 1588 613
rect 1582 608 1583 612
rect 1587 608 1588 612
rect 1582 607 1588 608
rect 1670 612 1676 613
rect 1670 608 1671 612
rect 1675 608 1676 612
rect 1670 607 1676 608
rect 1758 612 1764 613
rect 1758 608 1759 612
rect 1763 608 1764 612
rect 1758 607 1764 608
rect 1838 612 1844 613
rect 1838 608 1839 612
rect 1843 608 1844 612
rect 1838 607 1844 608
rect 1918 612 1924 613
rect 1918 608 1919 612
rect 1923 608 1924 612
rect 1918 607 1924 608
rect 2006 612 2012 613
rect 2006 608 2007 612
rect 2011 608 2012 612
rect 2006 607 2012 608
rect 2070 612 2076 613
rect 2070 608 2071 612
rect 2075 608 2076 612
rect 2070 607 2076 608
rect 134 600 140 601
rect 134 596 135 600
rect 139 596 140 600
rect 134 595 140 596
rect 174 600 180 601
rect 174 596 175 600
rect 179 596 180 600
rect 174 595 180 596
rect 214 600 220 601
rect 214 596 215 600
rect 219 596 220 600
rect 214 595 220 596
rect 254 600 260 601
rect 254 596 255 600
rect 259 596 260 600
rect 254 595 260 596
rect 302 600 308 601
rect 302 596 303 600
rect 307 596 308 600
rect 302 595 308 596
rect 350 600 356 601
rect 350 596 351 600
rect 355 596 356 600
rect 350 595 356 596
rect 398 600 404 601
rect 398 596 399 600
rect 403 596 404 600
rect 398 595 404 596
rect 438 600 444 601
rect 438 596 439 600
rect 443 596 444 600
rect 438 595 444 596
rect 486 600 492 601
rect 486 596 487 600
rect 491 596 492 600
rect 486 595 492 596
rect 534 600 540 601
rect 534 596 535 600
rect 539 596 540 600
rect 534 595 540 596
rect 582 600 588 601
rect 582 596 583 600
rect 587 596 588 600
rect 582 595 588 596
rect 630 600 636 601
rect 630 596 631 600
rect 635 596 636 600
rect 630 595 636 596
rect 678 600 684 601
rect 678 596 679 600
rect 683 596 684 600
rect 678 595 684 596
rect 726 600 732 601
rect 726 596 727 600
rect 731 596 732 600
rect 726 595 732 596
rect 110 592 116 593
rect 110 588 111 592
rect 115 588 116 592
rect 110 587 116 588
rect 1094 592 1100 593
rect 1094 588 1095 592
rect 1099 588 1100 592
rect 1094 587 1100 588
rect 110 575 116 576
rect 110 571 111 575
rect 115 571 116 575
rect 1094 575 1100 576
rect 110 570 116 571
rect 134 572 140 573
rect 134 568 135 572
rect 139 568 140 572
rect 134 567 140 568
rect 174 572 180 573
rect 174 568 175 572
rect 179 568 180 572
rect 174 567 180 568
rect 214 572 220 573
rect 214 568 215 572
rect 219 568 220 572
rect 214 567 220 568
rect 254 572 260 573
rect 254 568 255 572
rect 259 568 260 572
rect 254 567 260 568
rect 302 572 308 573
rect 302 568 303 572
rect 307 568 308 572
rect 302 567 308 568
rect 350 572 356 573
rect 350 568 351 572
rect 355 568 356 572
rect 350 567 356 568
rect 398 572 404 573
rect 398 568 399 572
rect 403 568 404 572
rect 398 567 404 568
rect 438 572 444 573
rect 438 568 439 572
rect 443 568 444 572
rect 438 567 444 568
rect 486 572 492 573
rect 486 568 487 572
rect 491 568 492 572
rect 486 567 492 568
rect 534 572 540 573
rect 534 568 535 572
rect 539 568 540 572
rect 534 567 540 568
rect 582 572 588 573
rect 582 568 583 572
rect 587 568 588 572
rect 582 567 588 568
rect 630 572 636 573
rect 630 568 631 572
rect 635 568 636 572
rect 630 567 636 568
rect 678 572 684 573
rect 678 568 679 572
rect 683 568 684 572
rect 678 567 684 568
rect 726 572 732 573
rect 726 568 727 572
rect 731 568 732 572
rect 1094 571 1095 575
rect 1099 571 1100 575
rect 1094 570 1100 571
rect 1158 572 1164 573
rect 726 567 732 568
rect 1158 568 1159 572
rect 1163 568 1164 572
rect 1158 567 1164 568
rect 1198 572 1204 573
rect 1198 568 1199 572
rect 1203 568 1204 572
rect 1198 567 1204 568
rect 1238 572 1244 573
rect 1238 568 1239 572
rect 1243 568 1244 572
rect 1238 567 1244 568
rect 1278 572 1284 573
rect 1278 568 1279 572
rect 1283 568 1284 572
rect 1278 567 1284 568
rect 1318 572 1324 573
rect 1318 568 1319 572
rect 1323 568 1324 572
rect 1318 567 1324 568
rect 1358 572 1364 573
rect 1358 568 1359 572
rect 1363 568 1364 572
rect 1358 567 1364 568
rect 1414 572 1420 573
rect 1414 568 1415 572
rect 1419 568 1420 572
rect 1414 567 1420 568
rect 1486 572 1492 573
rect 1486 568 1487 572
rect 1491 568 1492 572
rect 1486 567 1492 568
rect 1566 572 1572 573
rect 1566 568 1567 572
rect 1571 568 1572 572
rect 1566 567 1572 568
rect 1654 572 1660 573
rect 1654 568 1655 572
rect 1659 568 1660 572
rect 1654 567 1660 568
rect 1750 572 1756 573
rect 1750 568 1751 572
rect 1755 568 1756 572
rect 1750 567 1756 568
rect 1854 572 1860 573
rect 1854 568 1855 572
rect 1859 568 1860 572
rect 1854 567 1860 568
rect 1966 572 1972 573
rect 1966 568 1967 572
rect 1971 568 1972 572
rect 1966 567 1972 568
rect 2070 572 2076 573
rect 2070 568 2071 572
rect 2075 568 2076 572
rect 2070 567 2076 568
rect 1134 564 1140 565
rect 1134 560 1135 564
rect 1139 560 1140 564
rect 1134 559 1140 560
rect 2118 564 2124 565
rect 2118 560 2119 564
rect 2123 560 2124 564
rect 2118 559 2124 560
rect 134 556 140 557
rect 110 553 116 554
rect 110 549 111 553
rect 115 549 116 553
rect 134 552 135 556
rect 139 552 140 556
rect 134 551 140 552
rect 174 556 180 557
rect 174 552 175 556
rect 179 552 180 556
rect 174 551 180 552
rect 222 556 228 557
rect 222 552 223 556
rect 227 552 228 556
rect 222 551 228 552
rect 278 556 284 557
rect 278 552 279 556
rect 283 552 284 556
rect 278 551 284 552
rect 326 556 332 557
rect 326 552 327 556
rect 331 552 332 556
rect 326 551 332 552
rect 374 556 380 557
rect 374 552 375 556
rect 379 552 380 556
rect 374 551 380 552
rect 422 556 428 557
rect 422 552 423 556
rect 427 552 428 556
rect 422 551 428 552
rect 462 556 468 557
rect 462 552 463 556
rect 467 552 468 556
rect 462 551 468 552
rect 510 556 516 557
rect 510 552 511 556
rect 515 552 516 556
rect 510 551 516 552
rect 558 556 564 557
rect 558 552 559 556
rect 563 552 564 556
rect 558 551 564 552
rect 606 556 612 557
rect 606 552 607 556
rect 611 552 612 556
rect 606 551 612 552
rect 654 556 660 557
rect 654 552 655 556
rect 659 552 660 556
rect 654 551 660 552
rect 702 556 708 557
rect 702 552 703 556
rect 707 552 708 556
rect 702 551 708 552
rect 750 556 756 557
rect 750 552 751 556
rect 755 552 756 556
rect 750 551 756 552
rect 1094 553 1100 554
rect 110 548 116 549
rect 1094 549 1095 553
rect 1099 549 1100 553
rect 1094 548 1100 549
rect 1134 547 1140 548
rect 1134 543 1135 547
rect 1139 543 1140 547
rect 2118 547 2124 548
rect 1134 542 1140 543
rect 1158 544 1164 545
rect 1158 540 1159 544
rect 1163 540 1164 544
rect 1158 539 1164 540
rect 1198 544 1204 545
rect 1198 540 1199 544
rect 1203 540 1204 544
rect 1198 539 1204 540
rect 1238 544 1244 545
rect 1238 540 1239 544
rect 1243 540 1244 544
rect 1238 539 1244 540
rect 1278 544 1284 545
rect 1278 540 1279 544
rect 1283 540 1284 544
rect 1278 539 1284 540
rect 1318 544 1324 545
rect 1318 540 1319 544
rect 1323 540 1324 544
rect 1318 539 1324 540
rect 1358 544 1364 545
rect 1358 540 1359 544
rect 1363 540 1364 544
rect 1358 539 1364 540
rect 1414 544 1420 545
rect 1414 540 1415 544
rect 1419 540 1420 544
rect 1414 539 1420 540
rect 1486 544 1492 545
rect 1486 540 1487 544
rect 1491 540 1492 544
rect 1486 539 1492 540
rect 1566 544 1572 545
rect 1566 540 1567 544
rect 1571 540 1572 544
rect 1566 539 1572 540
rect 1654 544 1660 545
rect 1654 540 1655 544
rect 1659 540 1660 544
rect 1654 539 1660 540
rect 1750 544 1756 545
rect 1750 540 1751 544
rect 1755 540 1756 544
rect 1750 539 1756 540
rect 1854 544 1860 545
rect 1854 540 1855 544
rect 1859 540 1860 544
rect 1854 539 1860 540
rect 1966 544 1972 545
rect 1966 540 1967 544
rect 1971 540 1972 544
rect 1966 539 1972 540
rect 2070 544 2076 545
rect 2070 540 2071 544
rect 2075 540 2076 544
rect 2118 543 2119 547
rect 2123 543 2124 547
rect 2118 542 2124 543
rect 2070 539 2076 540
rect 110 536 116 537
rect 110 532 111 536
rect 115 532 116 536
rect 110 531 116 532
rect 1094 536 1100 537
rect 1094 532 1095 536
rect 1099 532 1100 536
rect 1094 531 1100 532
rect 134 528 140 529
rect 134 524 135 528
rect 139 524 140 528
rect 134 523 140 524
rect 174 528 180 529
rect 174 524 175 528
rect 179 524 180 528
rect 174 523 180 524
rect 222 528 228 529
rect 222 524 223 528
rect 227 524 228 528
rect 222 523 228 524
rect 278 528 284 529
rect 278 524 279 528
rect 283 524 284 528
rect 278 523 284 524
rect 326 528 332 529
rect 326 524 327 528
rect 331 524 332 528
rect 326 523 332 524
rect 374 528 380 529
rect 374 524 375 528
rect 379 524 380 528
rect 374 523 380 524
rect 422 528 428 529
rect 422 524 423 528
rect 427 524 428 528
rect 422 523 428 524
rect 462 528 468 529
rect 462 524 463 528
rect 467 524 468 528
rect 462 523 468 524
rect 510 528 516 529
rect 510 524 511 528
rect 515 524 516 528
rect 510 523 516 524
rect 558 528 564 529
rect 558 524 559 528
rect 563 524 564 528
rect 558 523 564 524
rect 606 528 612 529
rect 606 524 607 528
rect 611 524 612 528
rect 606 523 612 524
rect 654 528 660 529
rect 654 524 655 528
rect 659 524 660 528
rect 654 523 660 524
rect 702 528 708 529
rect 702 524 703 528
rect 707 524 708 528
rect 702 523 708 524
rect 750 528 756 529
rect 750 524 751 528
rect 755 524 756 528
rect 1302 528 1308 529
rect 750 523 756 524
rect 1134 525 1140 526
rect 1134 521 1135 525
rect 1139 521 1140 525
rect 1302 524 1303 528
rect 1307 524 1308 528
rect 1302 523 1308 524
rect 1342 528 1348 529
rect 1342 524 1343 528
rect 1347 524 1348 528
rect 1342 523 1348 524
rect 1382 528 1388 529
rect 1382 524 1383 528
rect 1387 524 1388 528
rect 1382 523 1388 524
rect 1422 528 1428 529
rect 1422 524 1423 528
rect 1427 524 1428 528
rect 1422 523 1428 524
rect 1462 528 1468 529
rect 1462 524 1463 528
rect 1467 524 1468 528
rect 1462 523 1468 524
rect 1502 528 1508 529
rect 1502 524 1503 528
rect 1507 524 1508 528
rect 1502 523 1508 524
rect 1542 528 1548 529
rect 1542 524 1543 528
rect 1547 524 1548 528
rect 1542 523 1548 524
rect 1590 528 1596 529
rect 1590 524 1591 528
rect 1595 524 1596 528
rect 1590 523 1596 524
rect 1646 528 1652 529
rect 1646 524 1647 528
rect 1651 524 1652 528
rect 1646 523 1652 524
rect 1702 528 1708 529
rect 1702 524 1703 528
rect 1707 524 1708 528
rect 1702 523 1708 524
rect 1766 528 1772 529
rect 1766 524 1767 528
rect 1771 524 1772 528
rect 1766 523 1772 524
rect 1838 528 1844 529
rect 1838 524 1839 528
rect 1843 524 1844 528
rect 1838 523 1844 524
rect 1918 528 1924 529
rect 1918 524 1919 528
rect 1923 524 1924 528
rect 1918 523 1924 524
rect 2006 528 2012 529
rect 2006 524 2007 528
rect 2011 524 2012 528
rect 2006 523 2012 524
rect 2070 528 2076 529
rect 2070 524 2071 528
rect 2075 524 2076 528
rect 2070 523 2076 524
rect 2118 525 2124 526
rect 1134 520 1140 521
rect 2118 521 2119 525
rect 2123 521 2124 525
rect 2118 520 2124 521
rect 1134 508 1140 509
rect 1134 504 1135 508
rect 1139 504 1140 508
rect 1134 503 1140 504
rect 2118 508 2124 509
rect 2118 504 2119 508
rect 2123 504 2124 508
rect 2118 503 2124 504
rect 1302 500 1308 501
rect 1302 496 1303 500
rect 1307 496 1308 500
rect 1302 495 1308 496
rect 1342 500 1348 501
rect 1342 496 1343 500
rect 1347 496 1348 500
rect 1342 495 1348 496
rect 1382 500 1388 501
rect 1382 496 1383 500
rect 1387 496 1388 500
rect 1382 495 1388 496
rect 1422 500 1428 501
rect 1422 496 1423 500
rect 1427 496 1428 500
rect 1422 495 1428 496
rect 1462 500 1468 501
rect 1462 496 1463 500
rect 1467 496 1468 500
rect 1462 495 1468 496
rect 1502 500 1508 501
rect 1502 496 1503 500
rect 1507 496 1508 500
rect 1502 495 1508 496
rect 1542 500 1548 501
rect 1542 496 1543 500
rect 1547 496 1548 500
rect 1542 495 1548 496
rect 1590 500 1596 501
rect 1590 496 1591 500
rect 1595 496 1596 500
rect 1590 495 1596 496
rect 1646 500 1652 501
rect 1646 496 1647 500
rect 1651 496 1652 500
rect 1646 495 1652 496
rect 1702 500 1708 501
rect 1702 496 1703 500
rect 1707 496 1708 500
rect 1702 495 1708 496
rect 1766 500 1772 501
rect 1766 496 1767 500
rect 1771 496 1772 500
rect 1766 495 1772 496
rect 1838 500 1844 501
rect 1838 496 1839 500
rect 1843 496 1844 500
rect 1838 495 1844 496
rect 1918 500 1924 501
rect 1918 496 1919 500
rect 1923 496 1924 500
rect 1918 495 1924 496
rect 2006 500 2012 501
rect 2006 496 2007 500
rect 2011 496 2012 500
rect 2006 495 2012 496
rect 2070 500 2076 501
rect 2070 496 2071 500
rect 2075 496 2076 500
rect 2070 495 2076 496
rect 134 484 140 485
rect 134 480 135 484
rect 139 480 140 484
rect 134 479 140 480
rect 174 484 180 485
rect 174 480 175 484
rect 179 480 180 484
rect 174 479 180 480
rect 230 484 236 485
rect 230 480 231 484
rect 235 480 236 484
rect 230 479 236 480
rect 294 484 300 485
rect 294 480 295 484
rect 299 480 300 484
rect 294 479 300 480
rect 358 484 364 485
rect 358 480 359 484
rect 363 480 364 484
rect 358 479 364 480
rect 422 484 428 485
rect 422 480 423 484
rect 427 480 428 484
rect 422 479 428 480
rect 478 484 484 485
rect 478 480 479 484
rect 483 480 484 484
rect 478 479 484 480
rect 534 484 540 485
rect 534 480 535 484
rect 539 480 540 484
rect 534 479 540 480
rect 590 484 596 485
rect 590 480 591 484
rect 595 480 596 484
rect 590 479 596 480
rect 638 484 644 485
rect 638 480 639 484
rect 643 480 644 484
rect 638 479 644 480
rect 686 484 692 485
rect 686 480 687 484
rect 691 480 692 484
rect 686 479 692 480
rect 734 484 740 485
rect 734 480 735 484
rect 739 480 740 484
rect 734 479 740 480
rect 790 484 796 485
rect 790 480 791 484
rect 795 480 796 484
rect 790 479 796 480
rect 846 484 852 485
rect 846 480 847 484
rect 851 480 852 484
rect 846 479 852 480
rect 110 476 116 477
rect 110 472 111 476
rect 115 472 116 476
rect 110 471 116 472
rect 1094 476 1100 477
rect 1094 472 1095 476
rect 1099 472 1100 476
rect 1094 471 1100 472
rect 1294 464 1300 465
rect 1294 460 1295 464
rect 1299 460 1300 464
rect 110 459 116 460
rect 110 455 111 459
rect 115 455 116 459
rect 1094 459 1100 460
rect 1294 459 1300 460
rect 1334 464 1340 465
rect 1334 460 1335 464
rect 1339 460 1340 464
rect 1334 459 1340 460
rect 1374 464 1380 465
rect 1374 460 1375 464
rect 1379 460 1380 464
rect 1374 459 1380 460
rect 1422 464 1428 465
rect 1422 460 1423 464
rect 1427 460 1428 464
rect 1422 459 1428 460
rect 1470 464 1476 465
rect 1470 460 1471 464
rect 1475 460 1476 464
rect 1470 459 1476 460
rect 1526 464 1532 465
rect 1526 460 1527 464
rect 1531 460 1532 464
rect 1526 459 1532 460
rect 1582 464 1588 465
rect 1582 460 1583 464
rect 1587 460 1588 464
rect 1582 459 1588 460
rect 1646 464 1652 465
rect 1646 460 1647 464
rect 1651 460 1652 464
rect 1646 459 1652 460
rect 1718 464 1724 465
rect 1718 460 1719 464
rect 1723 460 1724 464
rect 1718 459 1724 460
rect 1806 464 1812 465
rect 1806 460 1807 464
rect 1811 460 1812 464
rect 1806 459 1812 460
rect 1894 464 1900 465
rect 1894 460 1895 464
rect 1899 460 1900 464
rect 1894 459 1900 460
rect 1990 464 1996 465
rect 1990 460 1991 464
rect 1995 460 1996 464
rect 1990 459 1996 460
rect 2070 464 2076 465
rect 2070 460 2071 464
rect 2075 460 2076 464
rect 2070 459 2076 460
rect 110 454 116 455
rect 134 456 140 457
rect 134 452 135 456
rect 139 452 140 456
rect 134 451 140 452
rect 174 456 180 457
rect 174 452 175 456
rect 179 452 180 456
rect 174 451 180 452
rect 230 456 236 457
rect 230 452 231 456
rect 235 452 236 456
rect 230 451 236 452
rect 294 456 300 457
rect 294 452 295 456
rect 299 452 300 456
rect 294 451 300 452
rect 358 456 364 457
rect 358 452 359 456
rect 363 452 364 456
rect 358 451 364 452
rect 422 456 428 457
rect 422 452 423 456
rect 427 452 428 456
rect 422 451 428 452
rect 478 456 484 457
rect 478 452 479 456
rect 483 452 484 456
rect 478 451 484 452
rect 534 456 540 457
rect 534 452 535 456
rect 539 452 540 456
rect 534 451 540 452
rect 590 456 596 457
rect 590 452 591 456
rect 595 452 596 456
rect 590 451 596 452
rect 638 456 644 457
rect 638 452 639 456
rect 643 452 644 456
rect 638 451 644 452
rect 686 456 692 457
rect 686 452 687 456
rect 691 452 692 456
rect 686 451 692 452
rect 734 456 740 457
rect 734 452 735 456
rect 739 452 740 456
rect 734 451 740 452
rect 790 456 796 457
rect 790 452 791 456
rect 795 452 796 456
rect 790 451 796 452
rect 846 456 852 457
rect 846 452 847 456
rect 851 452 852 456
rect 1094 455 1095 459
rect 1099 455 1100 459
rect 1094 454 1100 455
rect 1134 456 1140 457
rect 846 451 852 452
rect 1134 452 1135 456
rect 1139 452 1140 456
rect 1134 451 1140 452
rect 2118 456 2124 457
rect 2118 452 2119 456
rect 2123 452 2124 456
rect 2118 451 2124 452
rect 174 440 180 441
rect 110 437 116 438
rect 110 433 111 437
rect 115 433 116 437
rect 174 436 175 440
rect 179 436 180 440
rect 174 435 180 436
rect 214 440 220 441
rect 214 436 215 440
rect 219 436 220 440
rect 214 435 220 436
rect 262 440 268 441
rect 262 436 263 440
rect 267 436 268 440
rect 262 435 268 436
rect 326 440 332 441
rect 326 436 327 440
rect 331 436 332 440
rect 326 435 332 436
rect 390 440 396 441
rect 390 436 391 440
rect 395 436 396 440
rect 390 435 396 436
rect 462 440 468 441
rect 462 436 463 440
rect 467 436 468 440
rect 462 435 468 436
rect 534 440 540 441
rect 534 436 535 440
rect 539 436 540 440
rect 534 435 540 436
rect 606 440 612 441
rect 606 436 607 440
rect 611 436 612 440
rect 606 435 612 436
rect 678 440 684 441
rect 678 436 679 440
rect 683 436 684 440
rect 678 435 684 436
rect 742 440 748 441
rect 742 436 743 440
rect 747 436 748 440
rect 742 435 748 436
rect 806 440 812 441
rect 806 436 807 440
rect 811 436 812 440
rect 806 435 812 436
rect 870 440 876 441
rect 870 436 871 440
rect 875 436 876 440
rect 870 435 876 436
rect 942 440 948 441
rect 942 436 943 440
rect 947 436 948 440
rect 1134 439 1140 440
rect 942 435 948 436
rect 1094 437 1100 438
rect 110 432 116 433
rect 1094 433 1095 437
rect 1099 433 1100 437
rect 1134 435 1135 439
rect 1139 435 1140 439
rect 2118 439 2124 440
rect 1134 434 1140 435
rect 1294 436 1300 437
rect 1094 432 1100 433
rect 1294 432 1295 436
rect 1299 432 1300 436
rect 1294 431 1300 432
rect 1334 436 1340 437
rect 1334 432 1335 436
rect 1339 432 1340 436
rect 1334 431 1340 432
rect 1374 436 1380 437
rect 1374 432 1375 436
rect 1379 432 1380 436
rect 1374 431 1380 432
rect 1422 436 1428 437
rect 1422 432 1423 436
rect 1427 432 1428 436
rect 1422 431 1428 432
rect 1470 436 1476 437
rect 1470 432 1471 436
rect 1475 432 1476 436
rect 1470 431 1476 432
rect 1526 436 1532 437
rect 1526 432 1527 436
rect 1531 432 1532 436
rect 1526 431 1532 432
rect 1582 436 1588 437
rect 1582 432 1583 436
rect 1587 432 1588 436
rect 1582 431 1588 432
rect 1646 436 1652 437
rect 1646 432 1647 436
rect 1651 432 1652 436
rect 1646 431 1652 432
rect 1718 436 1724 437
rect 1718 432 1719 436
rect 1723 432 1724 436
rect 1718 431 1724 432
rect 1806 436 1812 437
rect 1806 432 1807 436
rect 1811 432 1812 436
rect 1806 431 1812 432
rect 1894 436 1900 437
rect 1894 432 1895 436
rect 1899 432 1900 436
rect 1894 431 1900 432
rect 1990 436 1996 437
rect 1990 432 1991 436
rect 1995 432 1996 436
rect 1990 431 1996 432
rect 2070 436 2076 437
rect 2070 432 2071 436
rect 2075 432 2076 436
rect 2118 435 2119 439
rect 2123 435 2124 439
rect 2118 434 2124 435
rect 2070 431 2076 432
rect 1158 424 1164 425
rect 1134 421 1140 422
rect 110 420 116 421
rect 110 416 111 420
rect 115 416 116 420
rect 110 415 116 416
rect 1094 420 1100 421
rect 1094 416 1095 420
rect 1099 416 1100 420
rect 1134 417 1135 421
rect 1139 417 1140 421
rect 1158 420 1159 424
rect 1163 420 1164 424
rect 1158 419 1164 420
rect 1198 424 1204 425
rect 1198 420 1199 424
rect 1203 420 1204 424
rect 1198 419 1204 420
rect 1254 424 1260 425
rect 1254 420 1255 424
rect 1259 420 1260 424
rect 1254 419 1260 420
rect 1334 424 1340 425
rect 1334 420 1335 424
rect 1339 420 1340 424
rect 1334 419 1340 420
rect 1414 424 1420 425
rect 1414 420 1415 424
rect 1419 420 1420 424
rect 1414 419 1420 420
rect 1502 424 1508 425
rect 1502 420 1503 424
rect 1507 420 1508 424
rect 1502 419 1508 420
rect 1590 424 1596 425
rect 1590 420 1591 424
rect 1595 420 1596 424
rect 1590 419 1596 420
rect 1670 424 1676 425
rect 1670 420 1671 424
rect 1675 420 1676 424
rect 1670 419 1676 420
rect 1750 424 1756 425
rect 1750 420 1751 424
rect 1755 420 1756 424
rect 1750 419 1756 420
rect 1830 424 1836 425
rect 1830 420 1831 424
rect 1835 420 1836 424
rect 1830 419 1836 420
rect 1910 424 1916 425
rect 1910 420 1911 424
rect 1915 420 1916 424
rect 1910 419 1916 420
rect 1998 424 2004 425
rect 1998 420 1999 424
rect 2003 420 2004 424
rect 1998 419 2004 420
rect 2070 424 2076 425
rect 2070 420 2071 424
rect 2075 420 2076 424
rect 2070 419 2076 420
rect 2118 421 2124 422
rect 1134 416 1140 417
rect 2118 417 2119 421
rect 2123 417 2124 421
rect 2118 416 2124 417
rect 1094 415 1100 416
rect 174 412 180 413
rect 174 408 175 412
rect 179 408 180 412
rect 174 407 180 408
rect 214 412 220 413
rect 214 408 215 412
rect 219 408 220 412
rect 214 407 220 408
rect 262 412 268 413
rect 262 408 263 412
rect 267 408 268 412
rect 262 407 268 408
rect 326 412 332 413
rect 326 408 327 412
rect 331 408 332 412
rect 326 407 332 408
rect 390 412 396 413
rect 390 408 391 412
rect 395 408 396 412
rect 390 407 396 408
rect 462 412 468 413
rect 462 408 463 412
rect 467 408 468 412
rect 462 407 468 408
rect 534 412 540 413
rect 534 408 535 412
rect 539 408 540 412
rect 534 407 540 408
rect 606 412 612 413
rect 606 408 607 412
rect 611 408 612 412
rect 606 407 612 408
rect 678 412 684 413
rect 678 408 679 412
rect 683 408 684 412
rect 678 407 684 408
rect 742 412 748 413
rect 742 408 743 412
rect 747 408 748 412
rect 742 407 748 408
rect 806 412 812 413
rect 806 408 807 412
rect 811 408 812 412
rect 806 407 812 408
rect 870 412 876 413
rect 870 408 871 412
rect 875 408 876 412
rect 870 407 876 408
rect 942 412 948 413
rect 942 408 943 412
rect 947 408 948 412
rect 942 407 948 408
rect 1134 404 1140 405
rect 1134 400 1135 404
rect 1139 400 1140 404
rect 1134 399 1140 400
rect 2118 404 2124 405
rect 2118 400 2119 404
rect 2123 400 2124 404
rect 2118 399 2124 400
rect 1158 396 1164 397
rect 1158 392 1159 396
rect 1163 392 1164 396
rect 1158 391 1164 392
rect 1198 396 1204 397
rect 1198 392 1199 396
rect 1203 392 1204 396
rect 1198 391 1204 392
rect 1254 396 1260 397
rect 1254 392 1255 396
rect 1259 392 1260 396
rect 1254 391 1260 392
rect 1334 396 1340 397
rect 1334 392 1335 396
rect 1339 392 1340 396
rect 1334 391 1340 392
rect 1414 396 1420 397
rect 1414 392 1415 396
rect 1419 392 1420 396
rect 1414 391 1420 392
rect 1502 396 1508 397
rect 1502 392 1503 396
rect 1507 392 1508 396
rect 1502 391 1508 392
rect 1590 396 1596 397
rect 1590 392 1591 396
rect 1595 392 1596 396
rect 1590 391 1596 392
rect 1670 396 1676 397
rect 1670 392 1671 396
rect 1675 392 1676 396
rect 1670 391 1676 392
rect 1750 396 1756 397
rect 1750 392 1751 396
rect 1755 392 1756 396
rect 1750 391 1756 392
rect 1830 396 1836 397
rect 1830 392 1831 396
rect 1835 392 1836 396
rect 1830 391 1836 392
rect 1910 396 1916 397
rect 1910 392 1911 396
rect 1915 392 1916 396
rect 1910 391 1916 392
rect 1998 396 2004 397
rect 1998 392 1999 396
rect 2003 392 2004 396
rect 1998 391 2004 392
rect 2070 396 2076 397
rect 2070 392 2071 396
rect 2075 392 2076 396
rect 2070 391 2076 392
rect 174 368 180 369
rect 174 364 175 368
rect 179 364 180 368
rect 174 363 180 364
rect 214 368 220 369
rect 214 364 215 368
rect 219 364 220 368
rect 214 363 220 364
rect 270 368 276 369
rect 270 364 271 368
rect 275 364 276 368
rect 270 363 276 364
rect 334 368 340 369
rect 334 364 335 368
rect 339 364 340 368
rect 334 363 340 364
rect 406 368 412 369
rect 406 364 407 368
rect 411 364 412 368
rect 406 363 412 364
rect 486 368 492 369
rect 486 364 487 368
rect 491 364 492 368
rect 486 363 492 364
rect 566 368 572 369
rect 566 364 567 368
rect 571 364 572 368
rect 566 363 572 364
rect 638 368 644 369
rect 638 364 639 368
rect 643 364 644 368
rect 638 363 644 364
rect 710 368 716 369
rect 710 364 711 368
rect 715 364 716 368
rect 710 363 716 364
rect 774 368 780 369
rect 774 364 775 368
rect 779 364 780 368
rect 774 363 780 364
rect 838 368 844 369
rect 838 364 839 368
rect 843 364 844 368
rect 838 363 844 364
rect 894 368 900 369
rect 894 364 895 368
rect 899 364 900 368
rect 894 363 900 364
rect 950 368 956 369
rect 950 364 951 368
rect 955 364 956 368
rect 950 363 956 364
rect 1006 368 1012 369
rect 1006 364 1007 368
rect 1011 364 1012 368
rect 1006 363 1012 364
rect 1046 368 1052 369
rect 1046 364 1047 368
rect 1051 364 1052 368
rect 1046 363 1052 364
rect 110 360 116 361
rect 110 356 111 360
rect 115 356 116 360
rect 110 355 116 356
rect 1094 360 1100 361
rect 1094 356 1095 360
rect 1099 356 1100 360
rect 1094 355 1100 356
rect 1158 356 1164 357
rect 1158 352 1159 356
rect 1163 352 1164 356
rect 1158 351 1164 352
rect 1246 356 1252 357
rect 1246 352 1247 356
rect 1251 352 1252 356
rect 1246 351 1252 352
rect 1358 356 1364 357
rect 1358 352 1359 356
rect 1363 352 1364 356
rect 1358 351 1364 352
rect 1462 356 1468 357
rect 1462 352 1463 356
rect 1467 352 1468 356
rect 1462 351 1468 352
rect 1558 356 1564 357
rect 1558 352 1559 356
rect 1563 352 1564 356
rect 1558 351 1564 352
rect 1646 356 1652 357
rect 1646 352 1647 356
rect 1651 352 1652 356
rect 1646 351 1652 352
rect 1726 356 1732 357
rect 1726 352 1727 356
rect 1731 352 1732 356
rect 1726 351 1732 352
rect 1798 356 1804 357
rect 1798 352 1799 356
rect 1803 352 1804 356
rect 1798 351 1804 352
rect 1862 356 1868 357
rect 1862 352 1863 356
rect 1867 352 1868 356
rect 1862 351 1868 352
rect 1918 356 1924 357
rect 1918 352 1919 356
rect 1923 352 1924 356
rect 1918 351 1924 352
rect 1974 356 1980 357
rect 1974 352 1975 356
rect 1979 352 1980 356
rect 1974 351 1980 352
rect 2030 356 2036 357
rect 2030 352 2031 356
rect 2035 352 2036 356
rect 2030 351 2036 352
rect 2070 356 2076 357
rect 2070 352 2071 356
rect 2075 352 2076 356
rect 2070 351 2076 352
rect 1134 348 1140 349
rect 1134 344 1135 348
rect 1139 344 1140 348
rect 110 343 116 344
rect 110 339 111 343
rect 115 339 116 343
rect 1094 343 1100 344
rect 1134 343 1140 344
rect 2118 348 2124 349
rect 2118 344 2119 348
rect 2123 344 2124 348
rect 2118 343 2124 344
rect 110 338 116 339
rect 174 340 180 341
rect 174 336 175 340
rect 179 336 180 340
rect 174 335 180 336
rect 214 340 220 341
rect 214 336 215 340
rect 219 336 220 340
rect 214 335 220 336
rect 270 340 276 341
rect 270 336 271 340
rect 275 336 276 340
rect 270 335 276 336
rect 334 340 340 341
rect 334 336 335 340
rect 339 336 340 340
rect 334 335 340 336
rect 406 340 412 341
rect 406 336 407 340
rect 411 336 412 340
rect 406 335 412 336
rect 486 340 492 341
rect 486 336 487 340
rect 491 336 492 340
rect 486 335 492 336
rect 566 340 572 341
rect 566 336 567 340
rect 571 336 572 340
rect 566 335 572 336
rect 638 340 644 341
rect 638 336 639 340
rect 643 336 644 340
rect 638 335 644 336
rect 710 340 716 341
rect 710 336 711 340
rect 715 336 716 340
rect 710 335 716 336
rect 774 340 780 341
rect 774 336 775 340
rect 779 336 780 340
rect 774 335 780 336
rect 838 340 844 341
rect 838 336 839 340
rect 843 336 844 340
rect 838 335 844 336
rect 894 340 900 341
rect 894 336 895 340
rect 899 336 900 340
rect 894 335 900 336
rect 950 340 956 341
rect 950 336 951 340
rect 955 336 956 340
rect 950 335 956 336
rect 1006 340 1012 341
rect 1006 336 1007 340
rect 1011 336 1012 340
rect 1006 335 1012 336
rect 1046 340 1052 341
rect 1046 336 1047 340
rect 1051 336 1052 340
rect 1094 339 1095 343
rect 1099 339 1100 343
rect 1094 338 1100 339
rect 1046 335 1052 336
rect 1134 331 1140 332
rect 1134 327 1135 331
rect 1139 327 1140 331
rect 2118 331 2124 332
rect 1134 326 1140 327
rect 1158 328 1164 329
rect 382 324 388 325
rect 110 321 116 322
rect 110 317 111 321
rect 115 317 116 321
rect 382 320 383 324
rect 387 320 388 324
rect 382 319 388 320
rect 422 324 428 325
rect 422 320 423 324
rect 427 320 428 324
rect 422 319 428 320
rect 462 324 468 325
rect 462 320 463 324
rect 467 320 468 324
rect 462 319 468 320
rect 502 324 508 325
rect 502 320 503 324
rect 507 320 508 324
rect 502 319 508 320
rect 542 324 548 325
rect 542 320 543 324
rect 547 320 548 324
rect 542 319 548 320
rect 590 324 596 325
rect 590 320 591 324
rect 595 320 596 324
rect 590 319 596 320
rect 638 324 644 325
rect 638 320 639 324
rect 643 320 644 324
rect 638 319 644 320
rect 686 324 692 325
rect 686 320 687 324
rect 691 320 692 324
rect 686 319 692 320
rect 734 324 740 325
rect 734 320 735 324
rect 739 320 740 324
rect 734 319 740 320
rect 782 324 788 325
rect 782 320 783 324
rect 787 320 788 324
rect 782 319 788 320
rect 830 324 836 325
rect 830 320 831 324
rect 835 320 836 324
rect 830 319 836 320
rect 878 324 884 325
rect 878 320 879 324
rect 883 320 884 324
rect 878 319 884 320
rect 926 324 932 325
rect 926 320 927 324
rect 931 320 932 324
rect 926 319 932 320
rect 966 324 972 325
rect 966 320 967 324
rect 971 320 972 324
rect 966 319 972 320
rect 1006 324 1012 325
rect 1006 320 1007 324
rect 1011 320 1012 324
rect 1006 319 1012 320
rect 1046 324 1052 325
rect 1046 320 1047 324
rect 1051 320 1052 324
rect 1158 324 1159 328
rect 1163 324 1164 328
rect 1158 323 1164 324
rect 1246 328 1252 329
rect 1246 324 1247 328
rect 1251 324 1252 328
rect 1246 323 1252 324
rect 1358 328 1364 329
rect 1358 324 1359 328
rect 1363 324 1364 328
rect 1358 323 1364 324
rect 1462 328 1468 329
rect 1462 324 1463 328
rect 1467 324 1468 328
rect 1462 323 1468 324
rect 1558 328 1564 329
rect 1558 324 1559 328
rect 1563 324 1564 328
rect 1558 323 1564 324
rect 1646 328 1652 329
rect 1646 324 1647 328
rect 1651 324 1652 328
rect 1646 323 1652 324
rect 1726 328 1732 329
rect 1726 324 1727 328
rect 1731 324 1732 328
rect 1726 323 1732 324
rect 1798 328 1804 329
rect 1798 324 1799 328
rect 1803 324 1804 328
rect 1798 323 1804 324
rect 1862 328 1868 329
rect 1862 324 1863 328
rect 1867 324 1868 328
rect 1862 323 1868 324
rect 1918 328 1924 329
rect 1918 324 1919 328
rect 1923 324 1924 328
rect 1918 323 1924 324
rect 1974 328 1980 329
rect 1974 324 1975 328
rect 1979 324 1980 328
rect 1974 323 1980 324
rect 2030 328 2036 329
rect 2030 324 2031 328
rect 2035 324 2036 328
rect 2030 323 2036 324
rect 2070 328 2076 329
rect 2070 324 2071 328
rect 2075 324 2076 328
rect 2118 327 2119 331
rect 2123 327 2124 331
rect 2118 326 2124 327
rect 2070 323 2076 324
rect 1046 319 1052 320
rect 1094 321 1100 322
rect 110 316 116 317
rect 1094 317 1095 321
rect 1099 317 1100 321
rect 1094 316 1100 317
rect 1350 308 1356 309
rect 1134 305 1140 306
rect 110 304 116 305
rect 110 300 111 304
rect 115 300 116 304
rect 110 299 116 300
rect 1094 304 1100 305
rect 1094 300 1095 304
rect 1099 300 1100 304
rect 1134 301 1135 305
rect 1139 301 1140 305
rect 1350 304 1351 308
rect 1355 304 1356 308
rect 1350 303 1356 304
rect 1390 308 1396 309
rect 1390 304 1391 308
rect 1395 304 1396 308
rect 1390 303 1396 304
rect 1430 308 1436 309
rect 1430 304 1431 308
rect 1435 304 1436 308
rect 1430 303 1436 304
rect 1470 308 1476 309
rect 1470 304 1471 308
rect 1475 304 1476 308
rect 1470 303 1476 304
rect 1510 308 1516 309
rect 1510 304 1511 308
rect 1515 304 1516 308
rect 1510 303 1516 304
rect 1558 308 1564 309
rect 1558 304 1559 308
rect 1563 304 1564 308
rect 1558 303 1564 304
rect 1614 308 1620 309
rect 1614 304 1615 308
rect 1619 304 1620 308
rect 1614 303 1620 304
rect 1670 308 1676 309
rect 1670 304 1671 308
rect 1675 304 1676 308
rect 1670 303 1676 304
rect 1734 308 1740 309
rect 1734 304 1735 308
rect 1739 304 1740 308
rect 1734 303 1740 304
rect 1806 308 1812 309
rect 1806 304 1807 308
rect 1811 304 1812 308
rect 1806 303 1812 304
rect 1886 308 1892 309
rect 1886 304 1887 308
rect 1891 304 1892 308
rect 1886 303 1892 304
rect 1966 308 1972 309
rect 1966 304 1967 308
rect 1971 304 1972 308
rect 1966 303 1972 304
rect 2046 308 2052 309
rect 2046 304 2047 308
rect 2051 304 2052 308
rect 2046 303 2052 304
rect 2118 305 2124 306
rect 1134 300 1140 301
rect 2118 301 2119 305
rect 2123 301 2124 305
rect 2118 300 2124 301
rect 1094 299 1100 300
rect 382 296 388 297
rect 382 292 383 296
rect 387 292 388 296
rect 382 291 388 292
rect 422 296 428 297
rect 422 292 423 296
rect 427 292 428 296
rect 422 291 428 292
rect 462 296 468 297
rect 462 292 463 296
rect 467 292 468 296
rect 462 291 468 292
rect 502 296 508 297
rect 502 292 503 296
rect 507 292 508 296
rect 502 291 508 292
rect 542 296 548 297
rect 542 292 543 296
rect 547 292 548 296
rect 542 291 548 292
rect 590 296 596 297
rect 590 292 591 296
rect 595 292 596 296
rect 590 291 596 292
rect 638 296 644 297
rect 638 292 639 296
rect 643 292 644 296
rect 638 291 644 292
rect 686 296 692 297
rect 686 292 687 296
rect 691 292 692 296
rect 686 291 692 292
rect 734 296 740 297
rect 734 292 735 296
rect 739 292 740 296
rect 734 291 740 292
rect 782 296 788 297
rect 782 292 783 296
rect 787 292 788 296
rect 782 291 788 292
rect 830 296 836 297
rect 830 292 831 296
rect 835 292 836 296
rect 830 291 836 292
rect 878 296 884 297
rect 878 292 879 296
rect 883 292 884 296
rect 878 291 884 292
rect 926 296 932 297
rect 926 292 927 296
rect 931 292 932 296
rect 926 291 932 292
rect 966 296 972 297
rect 966 292 967 296
rect 971 292 972 296
rect 966 291 972 292
rect 1006 296 1012 297
rect 1006 292 1007 296
rect 1011 292 1012 296
rect 1006 291 1012 292
rect 1046 296 1052 297
rect 1046 292 1047 296
rect 1051 292 1052 296
rect 1046 291 1052 292
rect 1134 288 1140 289
rect 1134 284 1135 288
rect 1139 284 1140 288
rect 1134 283 1140 284
rect 2118 288 2124 289
rect 2118 284 2119 288
rect 2123 284 2124 288
rect 2118 283 2124 284
rect 1350 280 1356 281
rect 1350 276 1351 280
rect 1355 276 1356 280
rect 1350 275 1356 276
rect 1390 280 1396 281
rect 1390 276 1391 280
rect 1395 276 1396 280
rect 1390 275 1396 276
rect 1430 280 1436 281
rect 1430 276 1431 280
rect 1435 276 1436 280
rect 1430 275 1436 276
rect 1470 280 1476 281
rect 1470 276 1471 280
rect 1475 276 1476 280
rect 1470 275 1476 276
rect 1510 280 1516 281
rect 1510 276 1511 280
rect 1515 276 1516 280
rect 1510 275 1516 276
rect 1558 280 1564 281
rect 1558 276 1559 280
rect 1563 276 1564 280
rect 1558 275 1564 276
rect 1614 280 1620 281
rect 1614 276 1615 280
rect 1619 276 1620 280
rect 1614 275 1620 276
rect 1670 280 1676 281
rect 1670 276 1671 280
rect 1675 276 1676 280
rect 1670 275 1676 276
rect 1734 280 1740 281
rect 1734 276 1735 280
rect 1739 276 1740 280
rect 1734 275 1740 276
rect 1806 280 1812 281
rect 1806 276 1807 280
rect 1811 276 1812 280
rect 1806 275 1812 276
rect 1886 280 1892 281
rect 1886 276 1887 280
rect 1891 276 1892 280
rect 1886 275 1892 276
rect 1966 280 1972 281
rect 1966 276 1967 280
rect 1971 276 1972 280
rect 1966 275 1972 276
rect 2046 280 2052 281
rect 2046 276 2047 280
rect 2051 276 2052 280
rect 2046 275 2052 276
rect 286 252 292 253
rect 286 248 287 252
rect 291 248 292 252
rect 286 247 292 248
rect 326 252 332 253
rect 326 248 327 252
rect 331 248 332 252
rect 326 247 332 248
rect 366 252 372 253
rect 366 248 367 252
rect 371 248 372 252
rect 366 247 372 248
rect 414 252 420 253
rect 414 248 415 252
rect 419 248 420 252
rect 414 247 420 248
rect 470 252 476 253
rect 470 248 471 252
rect 475 248 476 252
rect 470 247 476 248
rect 534 252 540 253
rect 534 248 535 252
rect 539 248 540 252
rect 534 247 540 248
rect 606 252 612 253
rect 606 248 607 252
rect 611 248 612 252
rect 606 247 612 248
rect 678 252 684 253
rect 678 248 679 252
rect 683 248 684 252
rect 678 247 684 248
rect 742 252 748 253
rect 742 248 743 252
rect 747 248 748 252
rect 742 247 748 248
rect 806 252 812 253
rect 806 248 807 252
rect 811 248 812 252
rect 806 247 812 248
rect 862 252 868 253
rect 862 248 863 252
rect 867 248 868 252
rect 862 247 868 248
rect 926 252 932 253
rect 926 248 927 252
rect 931 248 932 252
rect 926 247 932 248
rect 990 252 996 253
rect 990 248 991 252
rect 995 248 996 252
rect 990 247 996 248
rect 1046 252 1052 253
rect 1046 248 1047 252
rect 1051 248 1052 252
rect 1046 247 1052 248
rect 110 244 116 245
rect 110 240 111 244
rect 115 240 116 244
rect 110 239 116 240
rect 1094 244 1100 245
rect 1094 240 1095 244
rect 1099 240 1100 244
rect 1094 239 1100 240
rect 1262 244 1268 245
rect 1262 240 1263 244
rect 1267 240 1268 244
rect 1262 239 1268 240
rect 1302 244 1308 245
rect 1302 240 1303 244
rect 1307 240 1308 244
rect 1302 239 1308 240
rect 1342 244 1348 245
rect 1342 240 1343 244
rect 1347 240 1348 244
rect 1342 239 1348 240
rect 1382 244 1388 245
rect 1382 240 1383 244
rect 1387 240 1388 244
rect 1382 239 1388 240
rect 1422 244 1428 245
rect 1422 240 1423 244
rect 1427 240 1428 244
rect 1422 239 1428 240
rect 1462 244 1468 245
rect 1462 240 1463 244
rect 1467 240 1468 244
rect 1462 239 1468 240
rect 1502 244 1508 245
rect 1502 240 1503 244
rect 1507 240 1508 244
rect 1502 239 1508 240
rect 1542 244 1548 245
rect 1542 240 1543 244
rect 1547 240 1548 244
rect 1542 239 1548 240
rect 1598 244 1604 245
rect 1598 240 1599 244
rect 1603 240 1604 244
rect 1598 239 1604 240
rect 1670 244 1676 245
rect 1670 240 1671 244
rect 1675 240 1676 244
rect 1670 239 1676 240
rect 1758 244 1764 245
rect 1758 240 1759 244
rect 1763 240 1764 244
rect 1758 239 1764 240
rect 1862 244 1868 245
rect 1862 240 1863 244
rect 1867 240 1868 244
rect 1862 239 1868 240
rect 1974 244 1980 245
rect 1974 240 1975 244
rect 1979 240 1980 244
rect 1974 239 1980 240
rect 2070 244 2076 245
rect 2070 240 2071 244
rect 2075 240 2076 244
rect 2070 239 2076 240
rect 1134 236 1140 237
rect 1134 232 1135 236
rect 1139 232 1140 236
rect 1134 231 1140 232
rect 2118 236 2124 237
rect 2118 232 2119 236
rect 2123 232 2124 236
rect 2118 231 2124 232
rect 110 227 116 228
rect 110 223 111 227
rect 115 223 116 227
rect 1094 227 1100 228
rect 110 222 116 223
rect 286 224 292 225
rect 286 220 287 224
rect 291 220 292 224
rect 286 219 292 220
rect 326 224 332 225
rect 326 220 327 224
rect 331 220 332 224
rect 326 219 332 220
rect 366 224 372 225
rect 366 220 367 224
rect 371 220 372 224
rect 366 219 372 220
rect 414 224 420 225
rect 414 220 415 224
rect 419 220 420 224
rect 414 219 420 220
rect 470 224 476 225
rect 470 220 471 224
rect 475 220 476 224
rect 470 219 476 220
rect 534 224 540 225
rect 534 220 535 224
rect 539 220 540 224
rect 534 219 540 220
rect 606 224 612 225
rect 606 220 607 224
rect 611 220 612 224
rect 606 219 612 220
rect 678 224 684 225
rect 678 220 679 224
rect 683 220 684 224
rect 678 219 684 220
rect 742 224 748 225
rect 742 220 743 224
rect 747 220 748 224
rect 742 219 748 220
rect 806 224 812 225
rect 806 220 807 224
rect 811 220 812 224
rect 806 219 812 220
rect 862 224 868 225
rect 862 220 863 224
rect 867 220 868 224
rect 862 219 868 220
rect 926 224 932 225
rect 926 220 927 224
rect 931 220 932 224
rect 926 219 932 220
rect 990 224 996 225
rect 990 220 991 224
rect 995 220 996 224
rect 990 219 996 220
rect 1046 224 1052 225
rect 1046 220 1047 224
rect 1051 220 1052 224
rect 1094 223 1095 227
rect 1099 223 1100 227
rect 1094 222 1100 223
rect 1046 219 1052 220
rect 1134 219 1140 220
rect 1134 215 1135 219
rect 1139 215 1140 219
rect 2118 219 2124 220
rect 1134 214 1140 215
rect 1262 216 1268 217
rect 1262 212 1263 216
rect 1267 212 1268 216
rect 1262 211 1268 212
rect 1302 216 1308 217
rect 1302 212 1303 216
rect 1307 212 1308 216
rect 1302 211 1308 212
rect 1342 216 1348 217
rect 1342 212 1343 216
rect 1347 212 1348 216
rect 1342 211 1348 212
rect 1382 216 1388 217
rect 1382 212 1383 216
rect 1387 212 1388 216
rect 1382 211 1388 212
rect 1422 216 1428 217
rect 1422 212 1423 216
rect 1427 212 1428 216
rect 1422 211 1428 212
rect 1462 216 1468 217
rect 1462 212 1463 216
rect 1467 212 1468 216
rect 1462 211 1468 212
rect 1502 216 1508 217
rect 1502 212 1503 216
rect 1507 212 1508 216
rect 1502 211 1508 212
rect 1542 216 1548 217
rect 1542 212 1543 216
rect 1547 212 1548 216
rect 1542 211 1548 212
rect 1598 216 1604 217
rect 1598 212 1599 216
rect 1603 212 1604 216
rect 1598 211 1604 212
rect 1670 216 1676 217
rect 1670 212 1671 216
rect 1675 212 1676 216
rect 1670 211 1676 212
rect 1758 216 1764 217
rect 1758 212 1759 216
rect 1763 212 1764 216
rect 1758 211 1764 212
rect 1862 216 1868 217
rect 1862 212 1863 216
rect 1867 212 1868 216
rect 1862 211 1868 212
rect 1974 216 1980 217
rect 1974 212 1975 216
rect 1979 212 1980 216
rect 1974 211 1980 212
rect 2070 216 2076 217
rect 2070 212 2071 216
rect 2075 212 2076 216
rect 2118 215 2119 219
rect 2123 215 2124 219
rect 2118 214 2124 215
rect 2070 211 2076 212
rect 166 200 172 201
rect 110 197 116 198
rect 110 193 111 197
rect 115 193 116 197
rect 166 196 167 200
rect 171 196 172 200
rect 166 195 172 196
rect 206 200 212 201
rect 206 196 207 200
rect 211 196 212 200
rect 206 195 212 196
rect 246 200 252 201
rect 246 196 247 200
rect 251 196 252 200
rect 246 195 252 196
rect 294 200 300 201
rect 294 196 295 200
rect 299 196 300 200
rect 294 195 300 196
rect 342 200 348 201
rect 342 196 343 200
rect 347 196 348 200
rect 342 195 348 196
rect 398 200 404 201
rect 398 196 399 200
rect 403 196 404 200
rect 398 195 404 196
rect 462 200 468 201
rect 462 196 463 200
rect 467 196 468 200
rect 462 195 468 196
rect 526 200 532 201
rect 526 196 527 200
rect 531 196 532 200
rect 526 195 532 196
rect 598 200 604 201
rect 598 196 599 200
rect 603 196 604 200
rect 598 195 604 196
rect 670 200 676 201
rect 670 196 671 200
rect 675 196 676 200
rect 670 195 676 196
rect 750 200 756 201
rect 750 196 751 200
rect 755 196 756 200
rect 750 195 756 196
rect 830 200 836 201
rect 830 196 831 200
rect 835 196 836 200
rect 830 195 836 196
rect 910 200 916 201
rect 910 196 911 200
rect 915 196 916 200
rect 910 195 916 196
rect 990 200 996 201
rect 990 196 991 200
rect 995 196 996 200
rect 990 195 996 196
rect 1046 200 1052 201
rect 1046 196 1047 200
rect 1051 196 1052 200
rect 1182 200 1188 201
rect 1046 195 1052 196
rect 1094 197 1100 198
rect 110 192 116 193
rect 1094 193 1095 197
rect 1099 193 1100 197
rect 1094 192 1100 193
rect 1134 197 1140 198
rect 1134 193 1135 197
rect 1139 193 1140 197
rect 1182 196 1183 200
rect 1187 196 1188 200
rect 1182 195 1188 196
rect 1230 200 1236 201
rect 1230 196 1231 200
rect 1235 196 1236 200
rect 1230 195 1236 196
rect 1294 200 1300 201
rect 1294 196 1295 200
rect 1299 196 1300 200
rect 1294 195 1300 196
rect 1358 200 1364 201
rect 1358 196 1359 200
rect 1363 196 1364 200
rect 1358 195 1364 196
rect 1430 200 1436 201
rect 1430 196 1431 200
rect 1435 196 1436 200
rect 1430 195 1436 196
rect 1510 200 1516 201
rect 1510 196 1511 200
rect 1515 196 1516 200
rect 1510 195 1516 196
rect 1590 200 1596 201
rect 1590 196 1591 200
rect 1595 196 1596 200
rect 1590 195 1596 196
rect 1662 200 1668 201
rect 1662 196 1663 200
rect 1667 196 1668 200
rect 1662 195 1668 196
rect 1734 200 1740 201
rect 1734 196 1735 200
rect 1739 196 1740 200
rect 1734 195 1740 196
rect 1806 200 1812 201
rect 1806 196 1807 200
rect 1811 196 1812 200
rect 1806 195 1812 196
rect 1878 200 1884 201
rect 1878 196 1879 200
rect 1883 196 1884 200
rect 1878 195 1884 196
rect 1950 200 1956 201
rect 1950 196 1951 200
rect 1955 196 1956 200
rect 1950 195 1956 196
rect 2022 200 2028 201
rect 2022 196 2023 200
rect 2027 196 2028 200
rect 2022 195 2028 196
rect 2070 200 2076 201
rect 2070 196 2071 200
rect 2075 196 2076 200
rect 2070 195 2076 196
rect 2118 197 2124 198
rect 1134 192 1140 193
rect 2118 193 2119 197
rect 2123 193 2124 197
rect 2118 192 2124 193
rect 110 180 116 181
rect 110 176 111 180
rect 115 176 116 180
rect 110 175 116 176
rect 1094 180 1100 181
rect 1094 176 1095 180
rect 1099 176 1100 180
rect 1094 175 1100 176
rect 1134 180 1140 181
rect 1134 176 1135 180
rect 1139 176 1140 180
rect 1134 175 1140 176
rect 2118 180 2124 181
rect 2118 176 2119 180
rect 2123 176 2124 180
rect 2118 175 2124 176
rect 166 172 172 173
rect 166 168 167 172
rect 171 168 172 172
rect 166 167 172 168
rect 206 172 212 173
rect 206 168 207 172
rect 211 168 212 172
rect 206 167 212 168
rect 246 172 252 173
rect 246 168 247 172
rect 251 168 252 172
rect 246 167 252 168
rect 294 172 300 173
rect 294 168 295 172
rect 299 168 300 172
rect 294 167 300 168
rect 342 172 348 173
rect 342 168 343 172
rect 347 168 348 172
rect 342 167 348 168
rect 398 172 404 173
rect 398 168 399 172
rect 403 168 404 172
rect 398 167 404 168
rect 462 172 468 173
rect 462 168 463 172
rect 467 168 468 172
rect 462 167 468 168
rect 526 172 532 173
rect 526 168 527 172
rect 531 168 532 172
rect 526 167 532 168
rect 598 172 604 173
rect 598 168 599 172
rect 603 168 604 172
rect 598 167 604 168
rect 670 172 676 173
rect 670 168 671 172
rect 675 168 676 172
rect 670 167 676 168
rect 750 172 756 173
rect 750 168 751 172
rect 755 168 756 172
rect 750 167 756 168
rect 830 172 836 173
rect 830 168 831 172
rect 835 168 836 172
rect 830 167 836 168
rect 910 172 916 173
rect 910 168 911 172
rect 915 168 916 172
rect 910 167 916 168
rect 990 172 996 173
rect 990 168 991 172
rect 995 168 996 172
rect 990 167 996 168
rect 1046 172 1052 173
rect 1046 168 1047 172
rect 1051 168 1052 172
rect 1046 167 1052 168
rect 1182 172 1188 173
rect 1182 168 1183 172
rect 1187 168 1188 172
rect 1182 167 1188 168
rect 1230 172 1236 173
rect 1230 168 1231 172
rect 1235 168 1236 172
rect 1230 167 1236 168
rect 1294 172 1300 173
rect 1294 168 1295 172
rect 1299 168 1300 172
rect 1294 167 1300 168
rect 1358 172 1364 173
rect 1358 168 1359 172
rect 1363 168 1364 172
rect 1358 167 1364 168
rect 1430 172 1436 173
rect 1430 168 1431 172
rect 1435 168 1436 172
rect 1430 167 1436 168
rect 1510 172 1516 173
rect 1510 168 1511 172
rect 1515 168 1516 172
rect 1510 167 1516 168
rect 1590 172 1596 173
rect 1590 168 1591 172
rect 1595 168 1596 172
rect 1590 167 1596 168
rect 1662 172 1668 173
rect 1662 168 1663 172
rect 1667 168 1668 172
rect 1662 167 1668 168
rect 1734 172 1740 173
rect 1734 168 1735 172
rect 1739 168 1740 172
rect 1734 167 1740 168
rect 1806 172 1812 173
rect 1806 168 1807 172
rect 1811 168 1812 172
rect 1806 167 1812 168
rect 1878 172 1884 173
rect 1878 168 1879 172
rect 1883 168 1884 172
rect 1878 167 1884 168
rect 1950 172 1956 173
rect 1950 168 1951 172
rect 1955 168 1956 172
rect 1950 167 1956 168
rect 2022 172 2028 173
rect 2022 168 2023 172
rect 2027 168 2028 172
rect 2022 167 2028 168
rect 2070 172 2076 173
rect 2070 168 2071 172
rect 2075 168 2076 172
rect 2070 167 2076 168
rect 134 120 140 121
rect 134 116 135 120
rect 139 116 140 120
rect 134 115 140 116
rect 174 120 180 121
rect 174 116 175 120
rect 179 116 180 120
rect 174 115 180 116
rect 214 120 220 121
rect 214 116 215 120
rect 219 116 220 120
rect 214 115 220 116
rect 254 120 260 121
rect 254 116 255 120
rect 259 116 260 120
rect 254 115 260 116
rect 294 120 300 121
rect 294 116 295 120
rect 299 116 300 120
rect 294 115 300 116
rect 334 120 340 121
rect 334 116 335 120
rect 339 116 340 120
rect 334 115 340 116
rect 374 120 380 121
rect 374 116 375 120
rect 379 116 380 120
rect 374 115 380 116
rect 414 120 420 121
rect 414 116 415 120
rect 419 116 420 120
rect 414 115 420 116
rect 454 120 460 121
rect 454 116 455 120
rect 459 116 460 120
rect 454 115 460 116
rect 494 120 500 121
rect 494 116 495 120
rect 499 116 500 120
rect 494 115 500 116
rect 534 120 540 121
rect 534 116 535 120
rect 539 116 540 120
rect 534 115 540 116
rect 574 120 580 121
rect 574 116 575 120
rect 579 116 580 120
rect 574 115 580 116
rect 614 120 620 121
rect 614 116 615 120
rect 619 116 620 120
rect 614 115 620 116
rect 654 120 660 121
rect 654 116 655 120
rect 659 116 660 120
rect 654 115 660 116
rect 694 120 700 121
rect 694 116 695 120
rect 699 116 700 120
rect 694 115 700 116
rect 734 120 740 121
rect 734 116 735 120
rect 739 116 740 120
rect 734 115 740 116
rect 774 120 780 121
rect 774 116 775 120
rect 779 116 780 120
rect 774 115 780 116
rect 814 120 820 121
rect 814 116 815 120
rect 819 116 820 120
rect 814 115 820 116
rect 870 120 876 121
rect 870 116 871 120
rect 875 116 876 120
rect 870 115 876 116
rect 934 120 940 121
rect 934 116 935 120
rect 939 116 940 120
rect 934 115 940 116
rect 998 120 1004 121
rect 998 116 999 120
rect 1003 116 1004 120
rect 998 115 1004 116
rect 1046 120 1052 121
rect 1046 116 1047 120
rect 1051 116 1052 120
rect 1046 115 1052 116
rect 110 112 116 113
rect 110 108 111 112
rect 115 108 116 112
rect 110 107 116 108
rect 1094 112 1100 113
rect 1094 108 1095 112
rect 1099 108 1100 112
rect 1094 107 1100 108
rect 1158 112 1164 113
rect 1158 108 1159 112
rect 1163 108 1164 112
rect 1158 107 1164 108
rect 1198 112 1204 113
rect 1198 108 1199 112
rect 1203 108 1204 112
rect 1198 107 1204 108
rect 1238 112 1244 113
rect 1238 108 1239 112
rect 1243 108 1244 112
rect 1238 107 1244 108
rect 1278 112 1284 113
rect 1278 108 1279 112
rect 1283 108 1284 112
rect 1278 107 1284 108
rect 1318 112 1324 113
rect 1318 108 1319 112
rect 1323 108 1324 112
rect 1318 107 1324 108
rect 1366 112 1372 113
rect 1366 108 1367 112
rect 1371 108 1372 112
rect 1366 107 1372 108
rect 1430 112 1436 113
rect 1430 108 1431 112
rect 1435 108 1436 112
rect 1430 107 1436 108
rect 1494 112 1500 113
rect 1494 108 1495 112
rect 1499 108 1500 112
rect 1494 107 1500 108
rect 1558 112 1564 113
rect 1558 108 1559 112
rect 1563 108 1564 112
rect 1558 107 1564 108
rect 1614 112 1620 113
rect 1614 108 1615 112
rect 1619 108 1620 112
rect 1614 107 1620 108
rect 1670 112 1676 113
rect 1670 108 1671 112
rect 1675 108 1676 112
rect 1670 107 1676 108
rect 1718 112 1724 113
rect 1718 108 1719 112
rect 1723 108 1724 112
rect 1718 107 1724 108
rect 1766 112 1772 113
rect 1766 108 1767 112
rect 1771 108 1772 112
rect 1766 107 1772 108
rect 1806 112 1812 113
rect 1806 108 1807 112
rect 1811 108 1812 112
rect 1806 107 1812 108
rect 1854 112 1860 113
rect 1854 108 1855 112
rect 1859 108 1860 112
rect 1854 107 1860 108
rect 1902 112 1908 113
rect 1902 108 1903 112
rect 1907 108 1908 112
rect 1902 107 1908 108
rect 1950 112 1956 113
rect 1950 108 1951 112
rect 1955 108 1956 112
rect 1950 107 1956 108
rect 1990 112 1996 113
rect 1990 108 1991 112
rect 1995 108 1996 112
rect 1990 107 1996 108
rect 2030 112 2036 113
rect 2030 108 2031 112
rect 2035 108 2036 112
rect 2030 107 2036 108
rect 2070 112 2076 113
rect 2070 108 2071 112
rect 2075 108 2076 112
rect 2070 107 2076 108
rect 1134 104 1140 105
rect 1134 100 1135 104
rect 1139 100 1140 104
rect 1134 99 1140 100
rect 2118 104 2124 105
rect 2118 100 2119 104
rect 2123 100 2124 104
rect 2118 99 2124 100
rect 110 95 116 96
rect 110 91 111 95
rect 115 91 116 95
rect 1094 95 1100 96
rect 110 90 116 91
rect 134 92 140 93
rect 134 88 135 92
rect 139 88 140 92
rect 134 87 140 88
rect 174 92 180 93
rect 174 88 175 92
rect 179 88 180 92
rect 174 87 180 88
rect 214 92 220 93
rect 214 88 215 92
rect 219 88 220 92
rect 214 87 220 88
rect 254 92 260 93
rect 254 88 255 92
rect 259 88 260 92
rect 254 87 260 88
rect 294 92 300 93
rect 294 88 295 92
rect 299 88 300 92
rect 294 87 300 88
rect 334 92 340 93
rect 334 88 335 92
rect 339 88 340 92
rect 334 87 340 88
rect 374 92 380 93
rect 374 88 375 92
rect 379 88 380 92
rect 374 87 380 88
rect 414 92 420 93
rect 414 88 415 92
rect 419 88 420 92
rect 414 87 420 88
rect 454 92 460 93
rect 454 88 455 92
rect 459 88 460 92
rect 454 87 460 88
rect 494 92 500 93
rect 494 88 495 92
rect 499 88 500 92
rect 494 87 500 88
rect 534 92 540 93
rect 534 88 535 92
rect 539 88 540 92
rect 534 87 540 88
rect 574 92 580 93
rect 574 88 575 92
rect 579 88 580 92
rect 574 87 580 88
rect 614 92 620 93
rect 614 88 615 92
rect 619 88 620 92
rect 614 87 620 88
rect 654 92 660 93
rect 654 88 655 92
rect 659 88 660 92
rect 654 87 660 88
rect 694 92 700 93
rect 694 88 695 92
rect 699 88 700 92
rect 694 87 700 88
rect 734 92 740 93
rect 734 88 735 92
rect 739 88 740 92
rect 734 87 740 88
rect 774 92 780 93
rect 774 88 775 92
rect 779 88 780 92
rect 774 87 780 88
rect 814 92 820 93
rect 814 88 815 92
rect 819 88 820 92
rect 814 87 820 88
rect 870 92 876 93
rect 870 88 871 92
rect 875 88 876 92
rect 870 87 876 88
rect 934 92 940 93
rect 934 88 935 92
rect 939 88 940 92
rect 934 87 940 88
rect 998 92 1004 93
rect 998 88 999 92
rect 1003 88 1004 92
rect 998 87 1004 88
rect 1046 92 1052 93
rect 1046 88 1047 92
rect 1051 88 1052 92
rect 1094 91 1095 95
rect 1099 91 1100 95
rect 1094 90 1100 91
rect 1046 87 1052 88
rect 1134 87 1140 88
rect 1134 83 1135 87
rect 1139 83 1140 87
rect 2118 87 2124 88
rect 1134 82 1140 83
rect 1158 84 1164 85
rect 1158 80 1159 84
rect 1163 80 1164 84
rect 1158 79 1164 80
rect 1198 84 1204 85
rect 1198 80 1199 84
rect 1203 80 1204 84
rect 1198 79 1204 80
rect 1238 84 1244 85
rect 1238 80 1239 84
rect 1243 80 1244 84
rect 1238 79 1244 80
rect 1278 84 1284 85
rect 1278 80 1279 84
rect 1283 80 1284 84
rect 1278 79 1284 80
rect 1318 84 1324 85
rect 1318 80 1319 84
rect 1323 80 1324 84
rect 1318 79 1324 80
rect 1366 84 1372 85
rect 1366 80 1367 84
rect 1371 80 1372 84
rect 1366 79 1372 80
rect 1430 84 1436 85
rect 1430 80 1431 84
rect 1435 80 1436 84
rect 1430 79 1436 80
rect 1494 84 1500 85
rect 1494 80 1495 84
rect 1499 80 1500 84
rect 1494 79 1500 80
rect 1558 84 1564 85
rect 1558 80 1559 84
rect 1563 80 1564 84
rect 1558 79 1564 80
rect 1614 84 1620 85
rect 1614 80 1615 84
rect 1619 80 1620 84
rect 1614 79 1620 80
rect 1670 84 1676 85
rect 1670 80 1671 84
rect 1675 80 1676 84
rect 1670 79 1676 80
rect 1718 84 1724 85
rect 1718 80 1719 84
rect 1723 80 1724 84
rect 1718 79 1724 80
rect 1766 84 1772 85
rect 1766 80 1767 84
rect 1771 80 1772 84
rect 1766 79 1772 80
rect 1806 84 1812 85
rect 1806 80 1807 84
rect 1811 80 1812 84
rect 1806 79 1812 80
rect 1854 84 1860 85
rect 1854 80 1855 84
rect 1859 80 1860 84
rect 1854 79 1860 80
rect 1902 84 1908 85
rect 1902 80 1903 84
rect 1907 80 1908 84
rect 1902 79 1908 80
rect 1950 84 1956 85
rect 1950 80 1951 84
rect 1955 80 1956 84
rect 1950 79 1956 80
rect 1990 84 1996 85
rect 1990 80 1991 84
rect 1995 80 1996 84
rect 1990 79 1996 80
rect 2030 84 2036 85
rect 2030 80 2031 84
rect 2035 80 2036 84
rect 2030 79 2036 80
rect 2070 84 2076 85
rect 2070 80 2071 84
rect 2075 80 2076 84
rect 2118 83 2119 87
rect 2123 83 2124 87
rect 2118 82 2124 83
rect 2070 79 2076 80
<< m3c >>
rect 1343 2192 1347 2196
rect 1383 2192 1387 2196
rect 1423 2192 1427 2196
rect 1463 2192 1467 2196
rect 1503 2192 1507 2196
rect 1543 2192 1547 2196
rect 1583 2192 1587 2196
rect 1623 2192 1627 2196
rect 1663 2192 1667 2196
rect 1703 2192 1707 2196
rect 1743 2192 1747 2196
rect 1783 2192 1787 2196
rect 1823 2192 1827 2196
rect 1135 2184 1139 2188
rect 2119 2184 2123 2188
rect 1135 2167 1139 2171
rect 1343 2164 1347 2168
rect 1383 2164 1387 2168
rect 1423 2164 1427 2168
rect 1463 2164 1467 2168
rect 1503 2164 1507 2168
rect 1543 2164 1547 2168
rect 1583 2164 1587 2168
rect 1623 2164 1627 2168
rect 1663 2164 1667 2168
rect 1703 2164 1707 2168
rect 1743 2164 1747 2168
rect 1783 2164 1787 2168
rect 1823 2164 1827 2168
rect 2119 2167 2123 2171
rect 1135 2149 1139 2153
rect 1287 2152 1291 2156
rect 1327 2152 1331 2156
rect 1367 2152 1371 2156
rect 1415 2152 1419 2156
rect 1463 2152 1467 2156
rect 1519 2152 1523 2156
rect 1575 2152 1579 2156
rect 1623 2152 1627 2156
rect 1671 2152 1675 2156
rect 1719 2152 1723 2156
rect 1775 2152 1779 2156
rect 1831 2152 1835 2156
rect 1887 2152 1891 2156
rect 2119 2149 2123 2153
rect 1135 2132 1139 2136
rect 2119 2132 2123 2136
rect 1287 2124 1291 2128
rect 1327 2124 1331 2128
rect 1367 2124 1371 2128
rect 1415 2124 1419 2128
rect 1463 2124 1467 2128
rect 1519 2124 1523 2128
rect 1575 2124 1579 2128
rect 1623 2124 1627 2128
rect 1671 2124 1675 2128
rect 1719 2124 1723 2128
rect 1775 2124 1779 2128
rect 1831 2124 1835 2128
rect 1887 2124 1891 2128
rect 1223 2084 1227 2088
rect 1279 2084 1283 2088
rect 1343 2084 1347 2088
rect 1423 2084 1427 2088
rect 1503 2084 1507 2088
rect 1583 2084 1587 2088
rect 1663 2084 1667 2088
rect 1743 2084 1747 2088
rect 1831 2084 1835 2088
rect 1919 2084 1923 2088
rect 2007 2084 2011 2088
rect 2071 2084 2075 2088
rect 1135 2076 1139 2080
rect 2119 2076 2123 2080
rect 1135 2059 1139 2063
rect 1223 2056 1227 2060
rect 1279 2056 1283 2060
rect 1343 2056 1347 2060
rect 1423 2056 1427 2060
rect 1503 2056 1507 2060
rect 1583 2056 1587 2060
rect 1663 2056 1667 2060
rect 1743 2056 1747 2060
rect 1831 2056 1835 2060
rect 1919 2056 1923 2060
rect 2007 2056 2011 2060
rect 2071 2056 2075 2060
rect 2119 2059 2123 2063
rect 1135 2041 1139 2045
rect 1183 2044 1187 2048
rect 1239 2044 1243 2048
rect 1311 2044 1315 2048
rect 1399 2044 1403 2048
rect 1487 2044 1491 2048
rect 1583 2044 1587 2048
rect 1671 2044 1675 2048
rect 1759 2044 1763 2048
rect 1839 2044 1843 2048
rect 1919 2044 1923 2048
rect 2007 2044 2011 2048
rect 2071 2044 2075 2048
rect 2119 2041 2123 2045
rect 1135 2024 1139 2028
rect 2119 2024 2123 2028
rect 191 2012 195 2016
rect 231 2012 235 2016
rect 287 2012 291 2016
rect 351 2012 355 2016
rect 423 2012 427 2016
rect 495 2012 499 2016
rect 575 2012 579 2016
rect 647 2012 651 2016
rect 719 2012 723 2016
rect 783 2012 787 2016
rect 839 2012 843 2016
rect 895 2012 899 2016
rect 951 2012 955 2016
rect 1007 2012 1011 2016
rect 1047 2012 1051 2016
rect 1183 2016 1187 2020
rect 1239 2016 1243 2020
rect 1311 2016 1315 2020
rect 1399 2016 1403 2020
rect 1487 2016 1491 2020
rect 1583 2016 1587 2020
rect 1671 2016 1675 2020
rect 1759 2016 1763 2020
rect 1839 2016 1843 2020
rect 1919 2016 1923 2020
rect 2007 2016 2011 2020
rect 2071 2016 2075 2020
rect 111 2004 115 2008
rect 1095 2004 1099 2008
rect 111 1987 115 1991
rect 191 1984 195 1988
rect 231 1984 235 1988
rect 287 1984 291 1988
rect 351 1984 355 1988
rect 423 1984 427 1988
rect 495 1984 499 1988
rect 575 1984 579 1988
rect 647 1984 651 1988
rect 719 1984 723 1988
rect 783 1984 787 1988
rect 839 1984 843 1988
rect 895 1984 899 1988
rect 951 1984 955 1988
rect 1007 1984 1011 1988
rect 1047 1984 1051 1988
rect 1095 1987 1099 1991
rect 1303 1980 1307 1984
rect 1383 1980 1387 1984
rect 1463 1980 1467 1984
rect 1543 1980 1547 1984
rect 1615 1980 1619 1984
rect 1687 1980 1691 1984
rect 1751 1980 1755 1984
rect 1815 1980 1819 1984
rect 1879 1980 1883 1984
rect 1951 1980 1955 1984
rect 2023 1980 2027 1984
rect 2071 1980 2075 1984
rect 111 1969 115 1973
rect 191 1972 195 1976
rect 247 1972 251 1976
rect 311 1972 315 1976
rect 375 1972 379 1976
rect 447 1972 451 1976
rect 519 1972 523 1976
rect 591 1972 595 1976
rect 655 1972 659 1976
rect 719 1972 723 1976
rect 775 1972 779 1976
rect 823 1972 827 1976
rect 871 1972 875 1976
rect 919 1972 923 1976
rect 967 1972 971 1976
rect 1007 1972 1011 1976
rect 1047 1972 1051 1976
rect 1095 1969 1099 1973
rect 1135 1972 1139 1976
rect 2119 1972 2123 1976
rect 111 1952 115 1956
rect 1095 1952 1099 1956
rect 1135 1955 1139 1959
rect 1303 1952 1307 1956
rect 1383 1952 1387 1956
rect 1463 1952 1467 1956
rect 1543 1952 1547 1956
rect 1615 1952 1619 1956
rect 1687 1952 1691 1956
rect 1751 1952 1755 1956
rect 1815 1952 1819 1956
rect 1879 1952 1883 1956
rect 1951 1952 1955 1956
rect 2023 1952 2027 1956
rect 2071 1952 2075 1956
rect 2119 1955 2123 1959
rect 191 1944 195 1948
rect 247 1944 251 1948
rect 311 1944 315 1948
rect 375 1944 379 1948
rect 447 1944 451 1948
rect 519 1944 523 1948
rect 591 1944 595 1948
rect 655 1944 659 1948
rect 719 1944 723 1948
rect 775 1944 779 1948
rect 823 1944 827 1948
rect 871 1944 875 1948
rect 919 1944 923 1948
rect 967 1944 971 1948
rect 1007 1944 1011 1948
rect 1047 1944 1051 1948
rect 1135 1933 1139 1937
rect 1159 1936 1163 1940
rect 1223 1936 1227 1940
rect 1303 1936 1307 1940
rect 1383 1936 1387 1940
rect 1463 1936 1467 1940
rect 1535 1936 1539 1940
rect 1615 1936 1619 1940
rect 1695 1936 1699 1940
rect 1783 1936 1787 1940
rect 1879 1936 1883 1940
rect 1983 1936 1987 1940
rect 2071 1936 2075 1940
rect 2119 1933 2123 1937
rect 1135 1916 1139 1920
rect 2119 1916 2123 1920
rect 135 1908 139 1912
rect 175 1908 179 1912
rect 231 1908 235 1912
rect 295 1908 299 1912
rect 367 1908 371 1912
rect 431 1908 435 1912
rect 495 1908 499 1912
rect 559 1908 563 1912
rect 615 1908 619 1912
rect 671 1908 675 1912
rect 727 1908 731 1912
rect 783 1908 787 1912
rect 847 1908 851 1912
rect 1159 1908 1163 1912
rect 1223 1908 1227 1912
rect 1303 1908 1307 1912
rect 1383 1908 1387 1912
rect 1463 1908 1467 1912
rect 1535 1908 1539 1912
rect 1615 1908 1619 1912
rect 1695 1908 1699 1912
rect 1783 1908 1787 1912
rect 1879 1908 1883 1912
rect 1983 1908 1987 1912
rect 2071 1908 2075 1912
rect 111 1900 115 1904
rect 1095 1900 1099 1904
rect 111 1883 115 1887
rect 135 1880 139 1884
rect 175 1880 179 1884
rect 231 1880 235 1884
rect 295 1880 299 1884
rect 367 1880 371 1884
rect 431 1880 435 1884
rect 495 1880 499 1884
rect 559 1880 563 1884
rect 615 1880 619 1884
rect 671 1880 675 1884
rect 727 1880 731 1884
rect 783 1880 787 1884
rect 847 1880 851 1884
rect 1095 1883 1099 1887
rect 111 1861 115 1865
rect 135 1864 139 1868
rect 199 1864 203 1868
rect 271 1864 275 1868
rect 335 1864 339 1868
rect 399 1864 403 1868
rect 455 1864 459 1868
rect 503 1864 507 1868
rect 551 1864 555 1868
rect 599 1864 603 1868
rect 647 1864 651 1868
rect 695 1864 699 1868
rect 751 1864 755 1868
rect 1159 1868 1163 1872
rect 1199 1868 1203 1872
rect 1263 1868 1267 1872
rect 1327 1868 1331 1872
rect 1391 1868 1395 1872
rect 1447 1868 1451 1872
rect 1503 1868 1507 1872
rect 1559 1868 1563 1872
rect 1631 1868 1635 1872
rect 1711 1868 1715 1872
rect 1799 1868 1803 1872
rect 1895 1868 1899 1872
rect 1991 1868 1995 1872
rect 2071 1868 2075 1872
rect 1095 1861 1099 1865
rect 1135 1860 1139 1864
rect 2119 1860 2123 1864
rect 111 1844 115 1848
rect 1095 1844 1099 1848
rect 1135 1843 1139 1847
rect 135 1836 139 1840
rect 199 1836 203 1840
rect 271 1836 275 1840
rect 335 1836 339 1840
rect 399 1836 403 1840
rect 455 1836 459 1840
rect 503 1836 507 1840
rect 551 1836 555 1840
rect 599 1836 603 1840
rect 647 1836 651 1840
rect 695 1836 699 1840
rect 751 1836 755 1840
rect 1159 1840 1163 1844
rect 1199 1840 1203 1844
rect 1263 1840 1267 1844
rect 1327 1840 1331 1844
rect 1391 1840 1395 1844
rect 1447 1840 1451 1844
rect 1503 1840 1507 1844
rect 1559 1840 1563 1844
rect 1631 1840 1635 1844
rect 1711 1840 1715 1844
rect 1799 1840 1803 1844
rect 1895 1840 1899 1844
rect 1991 1840 1995 1844
rect 2071 1840 2075 1844
rect 2119 1843 2123 1847
rect 1135 1825 1139 1829
rect 1159 1828 1163 1832
rect 1231 1828 1235 1832
rect 1303 1828 1307 1832
rect 1383 1828 1387 1832
rect 1463 1828 1467 1832
rect 1551 1828 1555 1832
rect 1647 1828 1651 1832
rect 1751 1828 1755 1832
rect 1855 1828 1859 1832
rect 1967 1828 1971 1832
rect 2071 1828 2075 1832
rect 2119 1825 2123 1829
rect 1135 1808 1139 1812
rect 2119 1808 2123 1812
rect 1159 1800 1163 1804
rect 1231 1800 1235 1804
rect 1303 1800 1307 1804
rect 1383 1800 1387 1804
rect 1463 1800 1467 1804
rect 1551 1800 1555 1804
rect 1647 1800 1651 1804
rect 1751 1800 1755 1804
rect 1855 1800 1859 1804
rect 1967 1800 1971 1804
rect 2071 1800 2075 1804
rect 151 1792 155 1796
rect 215 1792 219 1796
rect 271 1792 275 1796
rect 327 1792 331 1796
rect 383 1792 387 1796
rect 431 1792 435 1796
rect 479 1792 483 1796
rect 527 1792 531 1796
rect 575 1792 579 1796
rect 623 1792 627 1796
rect 671 1792 675 1796
rect 727 1792 731 1796
rect 111 1784 115 1788
rect 1095 1784 1099 1788
rect 111 1767 115 1771
rect 151 1764 155 1768
rect 215 1764 219 1768
rect 271 1764 275 1768
rect 327 1764 331 1768
rect 383 1764 387 1768
rect 431 1764 435 1768
rect 479 1764 483 1768
rect 527 1764 531 1768
rect 575 1764 579 1768
rect 623 1764 627 1768
rect 671 1764 675 1768
rect 727 1764 731 1768
rect 1095 1767 1099 1771
rect 1191 1764 1195 1768
rect 1255 1764 1259 1768
rect 1319 1764 1323 1768
rect 1383 1764 1387 1768
rect 1455 1764 1459 1768
rect 1527 1764 1531 1768
rect 1607 1764 1611 1768
rect 1687 1764 1691 1768
rect 1767 1764 1771 1768
rect 1847 1764 1851 1768
rect 1927 1764 1931 1768
rect 2007 1764 2011 1768
rect 2071 1764 2075 1768
rect 111 1749 115 1753
rect 231 1752 235 1756
rect 295 1752 299 1756
rect 351 1752 355 1756
rect 415 1752 419 1756
rect 479 1752 483 1756
rect 543 1752 547 1756
rect 615 1752 619 1756
rect 687 1752 691 1756
rect 759 1752 763 1756
rect 831 1752 835 1756
rect 911 1752 915 1756
rect 991 1752 995 1756
rect 1135 1756 1139 1760
rect 2119 1756 2123 1760
rect 1095 1749 1099 1753
rect 1135 1739 1139 1743
rect 111 1732 115 1736
rect 1095 1732 1099 1736
rect 1191 1736 1195 1740
rect 1255 1736 1259 1740
rect 1319 1736 1323 1740
rect 1383 1736 1387 1740
rect 1455 1736 1459 1740
rect 1527 1736 1531 1740
rect 1607 1736 1611 1740
rect 1687 1736 1691 1740
rect 1767 1736 1771 1740
rect 1847 1736 1851 1740
rect 1927 1736 1931 1740
rect 2007 1736 2011 1740
rect 2071 1736 2075 1740
rect 2119 1739 2123 1743
rect 231 1724 235 1728
rect 295 1724 299 1728
rect 351 1724 355 1728
rect 415 1724 419 1728
rect 479 1724 483 1728
rect 543 1724 547 1728
rect 615 1724 619 1728
rect 687 1724 691 1728
rect 759 1724 763 1728
rect 831 1724 835 1728
rect 911 1724 915 1728
rect 991 1724 995 1728
rect 1135 1721 1139 1725
rect 1247 1724 1251 1728
rect 1295 1724 1299 1728
rect 1343 1724 1347 1728
rect 1399 1724 1403 1728
rect 1463 1724 1467 1728
rect 1527 1724 1531 1728
rect 1599 1724 1603 1728
rect 1671 1724 1675 1728
rect 1743 1724 1747 1728
rect 1807 1724 1811 1728
rect 1879 1724 1883 1728
rect 1951 1724 1955 1728
rect 2023 1724 2027 1728
rect 2071 1724 2075 1728
rect 2119 1721 2123 1725
rect 1135 1704 1139 1708
rect 2119 1704 2123 1708
rect 1247 1696 1251 1700
rect 1295 1696 1299 1700
rect 1343 1696 1347 1700
rect 1399 1696 1403 1700
rect 1463 1696 1467 1700
rect 1527 1696 1531 1700
rect 1599 1696 1603 1700
rect 1671 1696 1675 1700
rect 1743 1696 1747 1700
rect 1807 1696 1811 1700
rect 1879 1696 1883 1700
rect 1951 1696 1955 1700
rect 2023 1696 2027 1700
rect 2071 1696 2075 1700
rect 135 1684 139 1688
rect 199 1684 203 1688
rect 279 1684 283 1688
rect 367 1684 371 1688
rect 463 1684 467 1688
rect 551 1684 555 1688
rect 639 1684 643 1688
rect 719 1684 723 1688
rect 791 1684 795 1688
rect 855 1684 859 1688
rect 919 1684 923 1688
rect 983 1684 987 1688
rect 1047 1684 1051 1688
rect 111 1676 115 1680
rect 1095 1676 1099 1680
rect 111 1659 115 1663
rect 135 1656 139 1660
rect 199 1656 203 1660
rect 279 1656 283 1660
rect 367 1656 371 1660
rect 463 1656 467 1660
rect 551 1656 555 1660
rect 639 1656 643 1660
rect 719 1656 723 1660
rect 791 1656 795 1660
rect 855 1656 859 1660
rect 919 1656 923 1660
rect 983 1656 987 1660
rect 1047 1656 1051 1660
rect 1095 1659 1099 1663
rect 1263 1656 1267 1660
rect 1303 1656 1307 1660
rect 1343 1656 1347 1660
rect 1391 1656 1395 1660
rect 1447 1656 1451 1660
rect 1503 1656 1507 1660
rect 1567 1656 1571 1660
rect 1631 1656 1635 1660
rect 1695 1656 1699 1660
rect 1759 1656 1763 1660
rect 1831 1656 1835 1660
rect 1911 1656 1915 1660
rect 1999 1656 2003 1660
rect 2071 1656 2075 1660
rect 1135 1648 1139 1652
rect 2119 1648 2123 1652
rect 111 1637 115 1641
rect 135 1640 139 1644
rect 183 1640 187 1644
rect 263 1640 267 1644
rect 343 1640 347 1644
rect 423 1640 427 1644
rect 503 1640 507 1644
rect 583 1640 587 1644
rect 655 1640 659 1644
rect 727 1640 731 1644
rect 791 1640 795 1644
rect 847 1640 851 1644
rect 903 1640 907 1644
rect 959 1640 963 1644
rect 1007 1640 1011 1644
rect 1047 1640 1051 1644
rect 1095 1637 1099 1641
rect 1135 1631 1139 1635
rect 1263 1628 1267 1632
rect 1303 1628 1307 1632
rect 1343 1628 1347 1632
rect 1391 1628 1395 1632
rect 1447 1628 1451 1632
rect 1503 1628 1507 1632
rect 1567 1628 1571 1632
rect 1631 1628 1635 1632
rect 1695 1628 1699 1632
rect 1759 1628 1763 1632
rect 1831 1628 1835 1632
rect 1911 1628 1915 1632
rect 1999 1628 2003 1632
rect 2071 1628 2075 1632
rect 2119 1631 2123 1635
rect 111 1620 115 1624
rect 1095 1620 1099 1624
rect 135 1612 139 1616
rect 183 1612 187 1616
rect 263 1612 267 1616
rect 343 1612 347 1616
rect 423 1612 427 1616
rect 503 1612 507 1616
rect 583 1612 587 1616
rect 655 1612 659 1616
rect 727 1612 731 1616
rect 791 1612 795 1616
rect 847 1612 851 1616
rect 903 1612 907 1616
rect 959 1612 963 1616
rect 1007 1612 1011 1616
rect 1047 1612 1051 1616
rect 1135 1601 1139 1605
rect 1159 1604 1163 1608
rect 1215 1604 1219 1608
rect 1303 1604 1307 1608
rect 1383 1604 1387 1608
rect 1463 1604 1467 1608
rect 1543 1604 1547 1608
rect 1623 1604 1627 1608
rect 1711 1604 1715 1608
rect 1799 1604 1803 1608
rect 1887 1604 1891 1608
rect 1983 1604 1987 1608
rect 2071 1604 2075 1608
rect 2119 1601 2123 1605
rect 1135 1584 1139 1588
rect 2119 1584 2123 1588
rect 135 1576 139 1580
rect 175 1576 179 1580
rect 231 1576 235 1580
rect 303 1576 307 1580
rect 375 1576 379 1580
rect 455 1576 459 1580
rect 527 1576 531 1580
rect 599 1576 603 1580
rect 671 1576 675 1580
rect 743 1576 747 1580
rect 815 1576 819 1580
rect 887 1576 891 1580
rect 1159 1576 1163 1580
rect 1215 1576 1219 1580
rect 1303 1576 1307 1580
rect 1383 1576 1387 1580
rect 1463 1576 1467 1580
rect 1543 1576 1547 1580
rect 1623 1576 1627 1580
rect 1711 1576 1715 1580
rect 1799 1576 1803 1580
rect 1887 1576 1891 1580
rect 1983 1576 1987 1580
rect 2071 1576 2075 1580
rect 111 1568 115 1572
rect 1095 1568 1099 1572
rect 111 1551 115 1555
rect 135 1548 139 1552
rect 175 1548 179 1552
rect 231 1548 235 1552
rect 303 1548 307 1552
rect 375 1548 379 1552
rect 455 1548 459 1552
rect 527 1548 531 1552
rect 599 1548 603 1552
rect 671 1548 675 1552
rect 743 1548 747 1552
rect 815 1548 819 1552
rect 887 1548 891 1552
rect 1095 1551 1099 1555
rect 111 1533 115 1537
rect 135 1536 139 1540
rect 175 1536 179 1540
rect 231 1536 235 1540
rect 311 1536 315 1540
rect 391 1536 395 1540
rect 479 1536 483 1540
rect 567 1536 571 1540
rect 655 1536 659 1540
rect 743 1536 747 1540
rect 823 1536 827 1540
rect 911 1536 915 1540
rect 999 1536 1003 1540
rect 1159 1540 1163 1544
rect 1199 1540 1203 1544
rect 1247 1540 1251 1544
rect 1319 1540 1323 1544
rect 1399 1540 1403 1544
rect 1479 1540 1483 1544
rect 1559 1540 1563 1544
rect 1647 1540 1651 1544
rect 1735 1540 1739 1544
rect 1823 1540 1827 1544
rect 1911 1540 1915 1544
rect 1999 1540 2003 1544
rect 2071 1540 2075 1544
rect 1095 1533 1099 1537
rect 1135 1532 1139 1536
rect 2119 1532 2123 1536
rect 111 1516 115 1520
rect 1095 1516 1099 1520
rect 1135 1515 1139 1519
rect 135 1508 139 1512
rect 175 1508 179 1512
rect 231 1508 235 1512
rect 311 1508 315 1512
rect 391 1508 395 1512
rect 479 1508 483 1512
rect 567 1508 571 1512
rect 655 1508 659 1512
rect 743 1508 747 1512
rect 823 1508 827 1512
rect 911 1508 915 1512
rect 999 1508 1003 1512
rect 1159 1512 1163 1516
rect 1199 1512 1203 1516
rect 1247 1512 1251 1516
rect 1319 1512 1323 1516
rect 1399 1512 1403 1516
rect 1479 1512 1483 1516
rect 1559 1512 1563 1516
rect 1647 1512 1651 1516
rect 1735 1512 1739 1516
rect 1823 1512 1827 1516
rect 1911 1512 1915 1516
rect 1999 1512 2003 1516
rect 2071 1512 2075 1516
rect 2119 1515 2123 1519
rect 1135 1497 1139 1501
rect 1159 1500 1163 1504
rect 1199 1500 1203 1504
rect 1239 1500 1243 1504
rect 1303 1500 1307 1504
rect 1375 1500 1379 1504
rect 1455 1500 1459 1504
rect 1543 1500 1547 1504
rect 1623 1500 1627 1504
rect 1703 1500 1707 1504
rect 1775 1500 1779 1504
rect 1847 1500 1851 1504
rect 1919 1500 1923 1504
rect 1991 1500 1995 1504
rect 2063 1500 2067 1504
rect 2119 1497 2123 1501
rect 1135 1480 1139 1484
rect 2119 1480 2123 1484
rect 135 1472 139 1476
rect 199 1472 203 1476
rect 279 1472 283 1476
rect 359 1472 363 1476
rect 439 1472 443 1476
rect 519 1472 523 1476
rect 599 1472 603 1476
rect 679 1472 683 1476
rect 767 1472 771 1476
rect 855 1472 859 1476
rect 943 1472 947 1476
rect 1031 1472 1035 1476
rect 1159 1472 1163 1476
rect 1199 1472 1203 1476
rect 1239 1472 1243 1476
rect 1303 1472 1307 1476
rect 1375 1472 1379 1476
rect 1455 1472 1459 1476
rect 1543 1472 1547 1476
rect 1623 1472 1627 1476
rect 1703 1472 1707 1476
rect 1775 1472 1779 1476
rect 1847 1472 1851 1476
rect 1919 1472 1923 1476
rect 1991 1472 1995 1476
rect 2063 1472 2067 1476
rect 111 1464 115 1468
rect 1095 1464 1099 1468
rect 111 1447 115 1451
rect 135 1444 139 1448
rect 199 1444 203 1448
rect 279 1444 283 1448
rect 359 1444 363 1448
rect 439 1444 443 1448
rect 519 1444 523 1448
rect 599 1444 603 1448
rect 679 1444 683 1448
rect 767 1444 771 1448
rect 855 1444 859 1448
rect 943 1444 947 1448
rect 1031 1444 1035 1448
rect 1095 1447 1099 1451
rect 111 1429 115 1433
rect 135 1432 139 1436
rect 191 1432 195 1436
rect 263 1432 267 1436
rect 335 1432 339 1436
rect 407 1432 411 1436
rect 479 1432 483 1436
rect 551 1432 555 1436
rect 631 1432 635 1436
rect 711 1432 715 1436
rect 799 1432 803 1436
rect 887 1432 891 1436
rect 975 1432 979 1436
rect 1047 1432 1051 1436
rect 1095 1429 1099 1433
rect 1279 1432 1283 1436
rect 1327 1432 1331 1436
rect 1383 1432 1387 1436
rect 1439 1432 1443 1436
rect 1495 1432 1499 1436
rect 1551 1432 1555 1436
rect 1607 1432 1611 1436
rect 1671 1432 1675 1436
rect 1735 1432 1739 1436
rect 1807 1432 1811 1436
rect 1887 1432 1891 1436
rect 1975 1432 1979 1436
rect 2063 1432 2067 1436
rect 1135 1424 1139 1428
rect 2119 1424 2123 1428
rect 111 1412 115 1416
rect 1095 1412 1099 1416
rect 135 1404 139 1408
rect 191 1404 195 1408
rect 263 1404 267 1408
rect 335 1404 339 1408
rect 407 1404 411 1408
rect 479 1404 483 1408
rect 551 1404 555 1408
rect 631 1404 635 1408
rect 711 1404 715 1408
rect 799 1404 803 1408
rect 887 1404 891 1408
rect 975 1404 979 1408
rect 1047 1404 1051 1408
rect 1135 1407 1139 1411
rect 1279 1404 1283 1408
rect 1327 1404 1331 1408
rect 1383 1404 1387 1408
rect 1439 1404 1443 1408
rect 1495 1404 1499 1408
rect 1551 1404 1555 1408
rect 1607 1404 1611 1408
rect 1671 1404 1675 1408
rect 1735 1404 1739 1408
rect 1807 1404 1811 1408
rect 1887 1404 1891 1408
rect 1975 1404 1979 1408
rect 2063 1404 2067 1408
rect 2119 1407 2123 1411
rect 1135 1385 1139 1389
rect 1335 1388 1339 1392
rect 1375 1388 1379 1392
rect 1415 1388 1419 1392
rect 1455 1388 1459 1392
rect 1495 1388 1499 1392
rect 1535 1388 1539 1392
rect 1583 1388 1587 1392
rect 1647 1388 1651 1392
rect 1719 1388 1723 1392
rect 1807 1388 1811 1392
rect 1895 1388 1899 1392
rect 1991 1388 1995 1392
rect 2071 1388 2075 1392
rect 2119 1385 2123 1389
rect 135 1368 139 1372
rect 175 1368 179 1372
rect 239 1368 243 1372
rect 303 1368 307 1372
rect 367 1368 371 1372
rect 439 1368 443 1372
rect 503 1368 507 1372
rect 575 1368 579 1372
rect 647 1368 651 1372
rect 711 1368 715 1372
rect 783 1368 787 1372
rect 855 1368 859 1372
rect 927 1368 931 1372
rect 999 1368 1003 1372
rect 1047 1368 1051 1372
rect 1135 1368 1139 1372
rect 2119 1368 2123 1372
rect 111 1360 115 1364
rect 1095 1360 1099 1364
rect 1335 1360 1339 1364
rect 1375 1360 1379 1364
rect 1415 1360 1419 1364
rect 1455 1360 1459 1364
rect 1495 1360 1499 1364
rect 1535 1360 1539 1364
rect 1583 1360 1587 1364
rect 1647 1360 1651 1364
rect 1719 1360 1723 1364
rect 1807 1360 1811 1364
rect 1895 1360 1899 1364
rect 1991 1360 1995 1364
rect 2071 1360 2075 1364
rect 111 1343 115 1347
rect 135 1340 139 1344
rect 175 1340 179 1344
rect 239 1340 243 1344
rect 303 1340 307 1344
rect 367 1340 371 1344
rect 439 1340 443 1344
rect 503 1340 507 1344
rect 575 1340 579 1344
rect 647 1340 651 1344
rect 711 1340 715 1344
rect 783 1340 787 1344
rect 855 1340 859 1344
rect 927 1340 931 1344
rect 999 1340 1003 1344
rect 1047 1340 1051 1344
rect 1095 1343 1099 1347
rect 111 1317 115 1321
rect 135 1320 139 1324
rect 175 1320 179 1324
rect 215 1320 219 1324
rect 255 1320 259 1324
rect 319 1320 323 1324
rect 391 1320 395 1324
rect 463 1320 467 1324
rect 543 1320 547 1324
rect 623 1320 627 1324
rect 703 1320 707 1324
rect 783 1320 787 1324
rect 863 1320 867 1324
rect 943 1320 947 1324
rect 1023 1320 1027 1324
rect 1159 1324 1163 1328
rect 1223 1324 1227 1328
rect 1311 1324 1315 1328
rect 1407 1324 1411 1328
rect 1503 1324 1507 1328
rect 1599 1324 1603 1328
rect 1679 1324 1683 1328
rect 1759 1324 1763 1328
rect 1831 1324 1835 1328
rect 1895 1324 1899 1328
rect 1959 1324 1963 1328
rect 2023 1324 2027 1328
rect 2071 1324 2075 1328
rect 1095 1317 1099 1321
rect 1135 1316 1139 1320
rect 2119 1316 2123 1320
rect 111 1300 115 1304
rect 1095 1300 1099 1304
rect 1135 1299 1139 1303
rect 135 1292 139 1296
rect 175 1292 179 1296
rect 215 1292 219 1296
rect 255 1292 259 1296
rect 319 1292 323 1296
rect 391 1292 395 1296
rect 463 1292 467 1296
rect 543 1292 547 1296
rect 623 1292 627 1296
rect 703 1292 707 1296
rect 783 1292 787 1296
rect 863 1292 867 1296
rect 943 1292 947 1296
rect 1023 1292 1027 1296
rect 1159 1296 1163 1300
rect 1223 1296 1227 1300
rect 1311 1296 1315 1300
rect 1407 1296 1411 1300
rect 1503 1296 1507 1300
rect 1599 1296 1603 1300
rect 1679 1296 1683 1300
rect 1759 1296 1763 1300
rect 1831 1296 1835 1300
rect 1895 1296 1899 1300
rect 1959 1296 1963 1300
rect 2023 1296 2027 1300
rect 2071 1296 2075 1300
rect 2119 1299 2123 1303
rect 1135 1281 1139 1285
rect 1175 1284 1179 1288
rect 1231 1284 1235 1288
rect 1303 1284 1307 1288
rect 1391 1284 1395 1288
rect 1479 1284 1483 1288
rect 1567 1284 1571 1288
rect 1655 1284 1659 1288
rect 1743 1284 1747 1288
rect 1831 1284 1835 1288
rect 1919 1284 1923 1288
rect 2007 1284 2011 1288
rect 2071 1284 2075 1288
rect 2119 1281 2123 1285
rect 1135 1264 1139 1268
rect 2119 1264 2123 1268
rect 135 1252 139 1256
rect 175 1252 179 1256
rect 215 1252 219 1256
rect 255 1252 259 1256
rect 319 1252 323 1256
rect 399 1252 403 1256
rect 487 1252 491 1256
rect 583 1252 587 1256
rect 687 1252 691 1256
rect 799 1252 803 1256
rect 919 1252 923 1256
rect 1047 1252 1051 1256
rect 1175 1256 1179 1260
rect 1231 1256 1235 1260
rect 1303 1256 1307 1260
rect 1391 1256 1395 1260
rect 1479 1256 1483 1260
rect 1567 1256 1571 1260
rect 1655 1256 1659 1260
rect 1743 1256 1747 1260
rect 1831 1256 1835 1260
rect 1919 1256 1923 1260
rect 2007 1256 2011 1260
rect 2071 1256 2075 1260
rect 111 1244 115 1248
rect 1095 1244 1099 1248
rect 111 1227 115 1231
rect 135 1224 139 1228
rect 175 1224 179 1228
rect 215 1224 219 1228
rect 255 1224 259 1228
rect 319 1224 323 1228
rect 399 1224 403 1228
rect 487 1224 491 1228
rect 583 1224 587 1228
rect 687 1224 691 1228
rect 799 1224 803 1228
rect 919 1224 923 1228
rect 1047 1224 1051 1228
rect 1095 1227 1099 1231
rect 1287 1216 1291 1220
rect 1327 1216 1331 1220
rect 1375 1216 1379 1220
rect 1431 1216 1435 1220
rect 1495 1216 1499 1220
rect 1559 1216 1563 1220
rect 1623 1216 1627 1220
rect 1679 1216 1683 1220
rect 1735 1216 1739 1220
rect 1791 1216 1795 1220
rect 1847 1216 1851 1220
rect 1903 1216 1907 1220
rect 1967 1216 1971 1220
rect 2031 1216 2035 1220
rect 2071 1216 2075 1220
rect 111 1205 115 1209
rect 271 1208 275 1212
rect 311 1208 315 1212
rect 351 1208 355 1212
rect 399 1208 403 1212
rect 447 1208 451 1212
rect 495 1208 499 1212
rect 551 1208 555 1212
rect 607 1208 611 1212
rect 671 1208 675 1212
rect 743 1208 747 1212
rect 815 1208 819 1212
rect 895 1208 899 1212
rect 983 1208 987 1212
rect 1095 1205 1099 1209
rect 1135 1208 1139 1212
rect 2119 1208 2123 1212
rect 111 1188 115 1192
rect 1095 1188 1099 1192
rect 1135 1191 1139 1195
rect 1287 1188 1291 1192
rect 1327 1188 1331 1192
rect 1375 1188 1379 1192
rect 1431 1188 1435 1192
rect 1495 1188 1499 1192
rect 1559 1188 1563 1192
rect 1623 1188 1627 1192
rect 1679 1188 1683 1192
rect 1735 1188 1739 1192
rect 1791 1188 1795 1192
rect 1847 1188 1851 1192
rect 1903 1188 1907 1192
rect 1967 1188 1971 1192
rect 2031 1188 2035 1192
rect 2071 1188 2075 1192
rect 2119 1191 2123 1195
rect 271 1180 275 1184
rect 311 1180 315 1184
rect 351 1180 355 1184
rect 399 1180 403 1184
rect 447 1180 451 1184
rect 495 1180 499 1184
rect 551 1180 555 1184
rect 607 1180 611 1184
rect 671 1180 675 1184
rect 743 1180 747 1184
rect 815 1180 819 1184
rect 895 1180 899 1184
rect 983 1180 987 1184
rect 1135 1173 1139 1177
rect 1159 1176 1163 1180
rect 1207 1176 1211 1180
rect 1279 1176 1283 1180
rect 1351 1176 1355 1180
rect 1423 1176 1427 1180
rect 1487 1176 1491 1180
rect 1559 1176 1563 1180
rect 1631 1176 1635 1180
rect 1711 1176 1715 1180
rect 1799 1176 1803 1180
rect 1887 1176 1891 1180
rect 1983 1176 1987 1180
rect 2071 1176 2075 1180
rect 2119 1173 2123 1177
rect 1135 1156 1139 1160
rect 2119 1156 2123 1160
rect 1159 1148 1163 1152
rect 1207 1148 1211 1152
rect 1279 1148 1283 1152
rect 1351 1148 1355 1152
rect 1423 1148 1427 1152
rect 1487 1148 1491 1152
rect 1559 1148 1563 1152
rect 1631 1148 1635 1152
rect 1711 1148 1715 1152
rect 1799 1148 1803 1152
rect 1887 1148 1891 1152
rect 1983 1148 1987 1152
rect 2071 1148 2075 1152
rect 399 1140 403 1144
rect 439 1140 443 1144
rect 479 1140 483 1144
rect 527 1140 531 1144
rect 575 1140 579 1144
rect 623 1140 627 1144
rect 671 1140 675 1144
rect 719 1140 723 1144
rect 775 1140 779 1144
rect 831 1140 835 1144
rect 887 1140 891 1144
rect 943 1140 947 1144
rect 1007 1140 1011 1144
rect 1047 1140 1051 1144
rect 111 1132 115 1136
rect 1095 1132 1099 1136
rect 111 1115 115 1119
rect 399 1112 403 1116
rect 439 1112 443 1116
rect 479 1112 483 1116
rect 527 1112 531 1116
rect 575 1112 579 1116
rect 623 1112 627 1116
rect 671 1112 675 1116
rect 719 1112 723 1116
rect 775 1112 779 1116
rect 831 1112 835 1116
rect 887 1112 891 1116
rect 943 1112 947 1116
rect 1007 1112 1011 1116
rect 1047 1112 1051 1116
rect 1095 1115 1099 1119
rect 1191 1108 1195 1112
rect 1271 1108 1275 1112
rect 1343 1108 1347 1112
rect 1415 1108 1419 1112
rect 1487 1108 1491 1112
rect 1567 1108 1571 1112
rect 1655 1108 1659 1112
rect 1751 1108 1755 1112
rect 1855 1108 1859 1112
rect 1959 1108 1963 1112
rect 2071 1108 2075 1112
rect 111 1097 115 1101
rect 159 1100 163 1104
rect 199 1100 203 1104
rect 255 1100 259 1104
rect 319 1100 323 1104
rect 399 1100 403 1104
rect 479 1100 483 1104
rect 559 1100 563 1104
rect 639 1100 643 1104
rect 711 1100 715 1104
rect 783 1100 787 1104
rect 855 1100 859 1104
rect 927 1100 931 1104
rect 999 1100 1003 1104
rect 1047 1100 1051 1104
rect 1095 1097 1099 1101
rect 1135 1100 1139 1104
rect 2119 1100 2123 1104
rect 111 1080 115 1084
rect 1095 1080 1099 1084
rect 1135 1083 1139 1087
rect 1191 1080 1195 1084
rect 1271 1080 1275 1084
rect 1343 1080 1347 1084
rect 1415 1080 1419 1084
rect 1487 1080 1491 1084
rect 1567 1080 1571 1084
rect 1655 1080 1659 1084
rect 1751 1080 1755 1084
rect 1855 1080 1859 1084
rect 1959 1080 1963 1084
rect 2071 1080 2075 1084
rect 2119 1083 2123 1087
rect 159 1072 163 1076
rect 199 1072 203 1076
rect 255 1072 259 1076
rect 319 1072 323 1076
rect 399 1072 403 1076
rect 479 1072 483 1076
rect 559 1072 563 1076
rect 639 1072 643 1076
rect 711 1072 715 1076
rect 783 1072 787 1076
rect 855 1072 859 1076
rect 927 1072 931 1076
rect 999 1072 1003 1076
rect 1047 1072 1051 1076
rect 1135 1065 1139 1069
rect 1159 1068 1163 1072
rect 1199 1068 1203 1072
rect 1247 1068 1251 1072
rect 1303 1068 1307 1072
rect 1351 1068 1355 1072
rect 1399 1068 1403 1072
rect 1455 1068 1459 1072
rect 1511 1068 1515 1072
rect 1583 1068 1587 1072
rect 1663 1068 1667 1072
rect 1759 1068 1763 1072
rect 1863 1068 1867 1072
rect 1967 1068 1971 1072
rect 2071 1068 2075 1072
rect 2119 1065 2123 1069
rect 1135 1048 1139 1052
rect 2119 1048 2123 1052
rect 1159 1040 1163 1044
rect 1199 1040 1203 1044
rect 1247 1040 1251 1044
rect 1303 1040 1307 1044
rect 1351 1040 1355 1044
rect 1399 1040 1403 1044
rect 1455 1040 1459 1044
rect 1511 1040 1515 1044
rect 1583 1040 1587 1044
rect 1663 1040 1667 1044
rect 1759 1040 1763 1044
rect 1863 1040 1867 1044
rect 1967 1040 1971 1044
rect 2071 1040 2075 1044
rect 135 1032 139 1036
rect 175 1032 179 1036
rect 215 1032 219 1036
rect 255 1032 259 1036
rect 319 1032 323 1036
rect 383 1032 387 1036
rect 447 1032 451 1036
rect 511 1032 515 1036
rect 575 1032 579 1036
rect 631 1032 635 1036
rect 687 1032 691 1036
rect 743 1032 747 1036
rect 799 1032 803 1036
rect 863 1032 867 1036
rect 111 1024 115 1028
rect 1095 1024 1099 1028
rect 111 1007 115 1011
rect 135 1004 139 1008
rect 175 1004 179 1008
rect 215 1004 219 1008
rect 255 1004 259 1008
rect 319 1004 323 1008
rect 383 1004 387 1008
rect 447 1004 451 1008
rect 511 1004 515 1008
rect 575 1004 579 1008
rect 631 1004 635 1008
rect 687 1004 691 1008
rect 743 1004 747 1008
rect 799 1004 803 1008
rect 863 1004 867 1008
rect 1095 1007 1099 1011
rect 1159 1000 1163 1004
rect 1199 1000 1203 1004
rect 1239 1000 1243 1004
rect 1295 1000 1299 1004
rect 1351 1000 1355 1004
rect 1407 1000 1411 1004
rect 1463 1000 1467 1004
rect 1519 1000 1523 1004
rect 1575 1000 1579 1004
rect 1639 1000 1643 1004
rect 1711 1000 1715 1004
rect 1791 1000 1795 1004
rect 1879 1000 1883 1004
rect 1967 1000 1971 1004
rect 2063 1000 2067 1004
rect 111 985 115 989
rect 135 988 139 992
rect 175 988 179 992
rect 223 988 227 992
rect 279 988 283 992
rect 343 988 347 992
rect 407 988 411 992
rect 471 988 475 992
rect 527 988 531 992
rect 583 988 587 992
rect 631 988 635 992
rect 687 988 691 992
rect 743 988 747 992
rect 799 988 803 992
rect 1135 992 1139 996
rect 2119 992 2123 996
rect 1095 985 1099 989
rect 1135 975 1139 979
rect 111 968 115 972
rect 1095 968 1099 972
rect 1159 972 1163 976
rect 1199 972 1203 976
rect 1239 972 1243 976
rect 1295 972 1299 976
rect 1351 972 1355 976
rect 1407 972 1411 976
rect 1463 972 1467 976
rect 1519 972 1523 976
rect 1575 972 1579 976
rect 1639 972 1643 976
rect 1711 972 1715 976
rect 1791 972 1795 976
rect 1879 972 1883 976
rect 1967 972 1971 976
rect 2063 972 2067 976
rect 2119 975 2123 979
rect 135 960 139 964
rect 175 960 179 964
rect 223 960 227 964
rect 279 960 283 964
rect 343 960 347 964
rect 407 960 411 964
rect 471 960 475 964
rect 527 960 531 964
rect 583 960 587 964
rect 631 960 635 964
rect 687 960 691 964
rect 743 960 747 964
rect 799 960 803 964
rect 1135 949 1139 953
rect 1159 952 1163 956
rect 1207 952 1211 956
rect 1287 952 1291 956
rect 1375 952 1379 956
rect 1455 952 1459 956
rect 1535 952 1539 956
rect 1615 952 1619 956
rect 1687 952 1691 956
rect 1751 952 1755 956
rect 1815 952 1819 956
rect 1879 952 1883 956
rect 1951 952 1955 956
rect 2023 952 2027 956
rect 2071 952 2075 956
rect 2119 949 2123 953
rect 1135 932 1139 936
rect 2119 932 2123 936
rect 263 920 267 924
rect 303 920 307 924
rect 351 920 355 924
rect 399 920 403 924
rect 455 920 459 924
rect 511 920 515 924
rect 567 920 571 924
rect 623 920 627 924
rect 687 920 691 924
rect 751 920 755 924
rect 815 920 819 924
rect 879 920 883 924
rect 943 920 947 924
rect 1007 920 1011 924
rect 1047 920 1051 924
rect 1159 924 1163 928
rect 1207 924 1211 928
rect 1287 924 1291 928
rect 1375 924 1379 928
rect 1455 924 1459 928
rect 1535 924 1539 928
rect 1615 924 1619 928
rect 1687 924 1691 928
rect 1751 924 1755 928
rect 1815 924 1819 928
rect 1879 924 1883 928
rect 1951 924 1955 928
rect 2023 924 2027 928
rect 2071 924 2075 928
rect 111 912 115 916
rect 1095 912 1099 916
rect 111 895 115 899
rect 263 892 267 896
rect 303 892 307 896
rect 351 892 355 896
rect 399 892 403 896
rect 455 892 459 896
rect 511 892 515 896
rect 567 892 571 896
rect 623 892 627 896
rect 687 892 691 896
rect 751 892 755 896
rect 815 892 819 896
rect 879 892 883 896
rect 943 892 947 896
rect 1007 892 1011 896
rect 1047 892 1051 896
rect 1095 895 1099 899
rect 1239 888 1243 892
rect 1319 888 1323 892
rect 1407 888 1411 892
rect 1495 888 1499 892
rect 1583 888 1587 892
rect 1663 888 1667 892
rect 1743 888 1747 892
rect 1815 888 1819 892
rect 1887 888 1891 892
rect 1951 888 1955 892
rect 2023 888 2027 892
rect 2071 888 2075 892
rect 111 873 115 877
rect 303 876 307 880
rect 351 876 355 880
rect 415 876 419 880
rect 479 876 483 880
rect 551 876 555 880
rect 623 876 627 880
rect 695 876 699 880
rect 767 876 771 880
rect 831 876 835 880
rect 887 876 891 880
rect 943 876 947 880
rect 1007 876 1011 880
rect 1047 876 1051 880
rect 1135 880 1139 884
rect 2119 880 2123 884
rect 1095 873 1099 877
rect 1135 863 1139 867
rect 111 856 115 860
rect 1095 856 1099 860
rect 1239 860 1243 864
rect 1319 860 1323 864
rect 1407 860 1411 864
rect 1495 860 1499 864
rect 1583 860 1587 864
rect 1663 860 1667 864
rect 1743 860 1747 864
rect 1815 860 1819 864
rect 1887 860 1891 864
rect 1951 860 1955 864
rect 2023 860 2027 864
rect 2071 860 2075 864
rect 2119 863 2123 867
rect 303 848 307 852
rect 351 848 355 852
rect 415 848 419 852
rect 479 848 483 852
rect 551 848 555 852
rect 623 848 627 852
rect 695 848 699 852
rect 767 848 771 852
rect 831 848 835 852
rect 887 848 891 852
rect 943 848 947 852
rect 1007 848 1011 852
rect 1047 848 1051 852
rect 1135 845 1139 849
rect 1159 848 1163 852
rect 1247 848 1251 852
rect 1359 848 1363 852
rect 1455 848 1459 852
rect 1543 848 1547 852
rect 1631 848 1635 852
rect 1711 848 1715 852
rect 1783 848 1787 852
rect 1855 848 1859 852
rect 1935 848 1939 852
rect 2015 848 2019 852
rect 2071 848 2075 852
rect 2119 845 2123 849
rect 1135 828 1139 832
rect 2119 828 2123 832
rect 1159 820 1163 824
rect 1247 820 1251 824
rect 1359 820 1363 824
rect 1455 820 1459 824
rect 1543 820 1547 824
rect 1631 820 1635 824
rect 1711 820 1715 824
rect 1783 820 1787 824
rect 1855 820 1859 824
rect 1935 820 1939 824
rect 2015 820 2019 824
rect 2071 820 2075 824
rect 279 812 283 816
rect 343 812 347 816
rect 415 812 419 816
rect 487 812 491 816
rect 567 812 571 816
rect 647 812 651 816
rect 727 812 731 816
rect 799 812 803 816
rect 863 812 867 816
rect 927 812 931 816
rect 999 812 1003 816
rect 1047 812 1051 816
rect 111 804 115 808
rect 1095 804 1099 808
rect 111 787 115 791
rect 279 784 283 788
rect 343 784 347 788
rect 415 784 419 788
rect 487 784 491 788
rect 567 784 571 788
rect 647 784 651 788
rect 727 784 731 788
rect 799 784 803 788
rect 863 784 867 788
rect 927 784 931 788
rect 999 784 1003 788
rect 1047 784 1051 788
rect 1095 787 1099 791
rect 1159 784 1163 788
rect 1279 784 1283 788
rect 1407 784 1411 788
rect 1519 784 1523 788
rect 1623 784 1627 788
rect 1719 784 1723 788
rect 1815 784 1819 788
rect 1903 784 1907 788
rect 1999 784 2003 788
rect 2071 784 2075 788
rect 111 769 115 773
rect 215 772 219 776
rect 279 772 283 776
rect 351 772 355 776
rect 423 772 427 776
rect 495 772 499 776
rect 567 772 571 776
rect 639 772 643 776
rect 703 772 707 776
rect 759 772 763 776
rect 815 772 819 776
rect 863 772 867 776
rect 911 772 915 776
rect 959 772 963 776
rect 1007 772 1011 776
rect 1047 772 1051 776
rect 1135 776 1139 780
rect 2119 776 2123 780
rect 1095 769 1099 773
rect 1135 759 1139 763
rect 111 752 115 756
rect 1095 752 1099 756
rect 1159 756 1163 760
rect 1279 756 1283 760
rect 1407 756 1411 760
rect 1519 756 1523 760
rect 1623 756 1627 760
rect 1719 756 1723 760
rect 1815 756 1819 760
rect 1903 756 1907 760
rect 1999 756 2003 760
rect 2071 756 2075 760
rect 2119 759 2123 763
rect 215 744 219 748
rect 279 744 283 748
rect 351 744 355 748
rect 423 744 427 748
rect 495 744 499 748
rect 567 744 571 748
rect 639 744 643 748
rect 703 744 707 748
rect 759 744 763 748
rect 815 744 819 748
rect 863 744 867 748
rect 911 744 915 748
rect 959 744 963 748
rect 1007 744 1011 748
rect 1047 744 1051 748
rect 1135 737 1139 741
rect 1335 740 1339 744
rect 1375 740 1379 744
rect 1415 740 1419 744
rect 1455 740 1459 744
rect 1503 740 1507 744
rect 1551 740 1555 744
rect 1599 740 1603 744
rect 1655 740 1659 744
rect 1711 740 1715 744
rect 1767 740 1771 744
rect 1831 740 1835 744
rect 1895 740 1899 744
rect 1959 740 1963 744
rect 2023 740 2027 744
rect 2071 740 2075 744
rect 2119 737 2123 741
rect 1135 720 1139 724
rect 2119 720 2123 724
rect 175 708 179 712
rect 239 708 243 712
rect 311 708 315 712
rect 391 708 395 712
rect 471 708 475 712
rect 543 708 547 712
rect 615 708 619 712
rect 679 708 683 712
rect 735 708 739 712
rect 799 708 803 712
rect 863 708 867 712
rect 927 708 931 712
rect 1335 712 1339 716
rect 1375 712 1379 716
rect 1415 712 1419 716
rect 1455 712 1459 716
rect 1503 712 1507 716
rect 1551 712 1555 716
rect 1599 712 1603 716
rect 1655 712 1659 716
rect 1711 712 1715 716
rect 1767 712 1771 716
rect 1831 712 1835 716
rect 1895 712 1899 716
rect 1959 712 1963 716
rect 2023 712 2027 716
rect 2071 712 2075 716
rect 111 700 115 704
rect 1095 700 1099 704
rect 111 683 115 687
rect 175 680 179 684
rect 239 680 243 684
rect 311 680 315 684
rect 391 680 395 684
rect 471 680 475 684
rect 543 680 547 684
rect 615 680 619 684
rect 679 680 683 684
rect 735 680 739 684
rect 799 680 803 684
rect 863 680 867 684
rect 927 680 931 684
rect 1095 683 1099 687
rect 1247 676 1251 680
rect 1287 676 1291 680
rect 1335 676 1339 680
rect 1391 676 1395 680
rect 1447 676 1451 680
rect 1511 676 1515 680
rect 1583 676 1587 680
rect 1655 676 1659 680
rect 1735 676 1739 680
rect 1823 676 1827 680
rect 1911 676 1915 680
rect 1999 676 2003 680
rect 2071 676 2075 680
rect 111 665 115 669
rect 135 668 139 672
rect 175 668 179 672
rect 215 668 219 672
rect 271 668 275 672
rect 335 668 339 672
rect 399 668 403 672
rect 463 668 467 672
rect 527 668 531 672
rect 591 668 595 672
rect 647 668 651 672
rect 703 668 707 672
rect 759 668 763 672
rect 823 668 827 672
rect 1095 665 1099 669
rect 1135 668 1139 672
rect 2119 668 2123 672
rect 111 648 115 652
rect 1095 648 1099 652
rect 1135 651 1139 655
rect 1247 648 1251 652
rect 1287 648 1291 652
rect 1335 648 1339 652
rect 1391 648 1395 652
rect 1447 648 1451 652
rect 1511 648 1515 652
rect 1583 648 1587 652
rect 1655 648 1659 652
rect 1735 648 1739 652
rect 1823 648 1827 652
rect 1911 648 1915 652
rect 1999 648 2003 652
rect 2071 648 2075 652
rect 2119 651 2123 655
rect 135 640 139 644
rect 175 640 179 644
rect 215 640 219 644
rect 271 640 275 644
rect 335 640 339 644
rect 399 640 403 644
rect 463 640 467 644
rect 527 640 531 644
rect 591 640 595 644
rect 647 640 651 644
rect 703 640 707 644
rect 759 640 763 644
rect 823 640 827 644
rect 1135 633 1139 637
rect 1159 636 1163 640
rect 1199 636 1203 640
rect 1239 636 1243 640
rect 1279 636 1283 640
rect 1343 636 1347 640
rect 1415 636 1419 640
rect 1495 636 1499 640
rect 1583 636 1587 640
rect 1671 636 1675 640
rect 1759 636 1763 640
rect 1839 636 1843 640
rect 1919 636 1923 640
rect 2007 636 2011 640
rect 2071 636 2075 640
rect 2119 633 2123 637
rect 1135 616 1139 620
rect 2119 616 2123 620
rect 1159 608 1163 612
rect 1199 608 1203 612
rect 1239 608 1243 612
rect 1279 608 1283 612
rect 1343 608 1347 612
rect 1415 608 1419 612
rect 1495 608 1499 612
rect 1583 608 1587 612
rect 1671 608 1675 612
rect 1759 608 1763 612
rect 1839 608 1843 612
rect 1919 608 1923 612
rect 2007 608 2011 612
rect 2071 608 2075 612
rect 135 596 139 600
rect 175 596 179 600
rect 215 596 219 600
rect 255 596 259 600
rect 303 596 307 600
rect 351 596 355 600
rect 399 596 403 600
rect 439 596 443 600
rect 487 596 491 600
rect 535 596 539 600
rect 583 596 587 600
rect 631 596 635 600
rect 679 596 683 600
rect 727 596 731 600
rect 111 588 115 592
rect 1095 588 1099 592
rect 111 571 115 575
rect 135 568 139 572
rect 175 568 179 572
rect 215 568 219 572
rect 255 568 259 572
rect 303 568 307 572
rect 351 568 355 572
rect 399 568 403 572
rect 439 568 443 572
rect 487 568 491 572
rect 535 568 539 572
rect 583 568 587 572
rect 631 568 635 572
rect 679 568 683 572
rect 727 568 731 572
rect 1095 571 1099 575
rect 1159 568 1163 572
rect 1199 568 1203 572
rect 1239 568 1243 572
rect 1279 568 1283 572
rect 1319 568 1323 572
rect 1359 568 1363 572
rect 1415 568 1419 572
rect 1487 568 1491 572
rect 1567 568 1571 572
rect 1655 568 1659 572
rect 1751 568 1755 572
rect 1855 568 1859 572
rect 1967 568 1971 572
rect 2071 568 2075 572
rect 1135 560 1139 564
rect 2119 560 2123 564
rect 111 549 115 553
rect 135 552 139 556
rect 175 552 179 556
rect 223 552 227 556
rect 279 552 283 556
rect 327 552 331 556
rect 375 552 379 556
rect 423 552 427 556
rect 463 552 467 556
rect 511 552 515 556
rect 559 552 563 556
rect 607 552 611 556
rect 655 552 659 556
rect 703 552 707 556
rect 751 552 755 556
rect 1095 549 1099 553
rect 1135 543 1139 547
rect 1159 540 1163 544
rect 1199 540 1203 544
rect 1239 540 1243 544
rect 1279 540 1283 544
rect 1319 540 1323 544
rect 1359 540 1363 544
rect 1415 540 1419 544
rect 1487 540 1491 544
rect 1567 540 1571 544
rect 1655 540 1659 544
rect 1751 540 1755 544
rect 1855 540 1859 544
rect 1967 540 1971 544
rect 2071 540 2075 544
rect 2119 543 2123 547
rect 111 532 115 536
rect 1095 532 1099 536
rect 135 524 139 528
rect 175 524 179 528
rect 223 524 227 528
rect 279 524 283 528
rect 327 524 331 528
rect 375 524 379 528
rect 423 524 427 528
rect 463 524 467 528
rect 511 524 515 528
rect 559 524 563 528
rect 607 524 611 528
rect 655 524 659 528
rect 703 524 707 528
rect 751 524 755 528
rect 1135 521 1139 525
rect 1303 524 1307 528
rect 1343 524 1347 528
rect 1383 524 1387 528
rect 1423 524 1427 528
rect 1463 524 1467 528
rect 1503 524 1507 528
rect 1543 524 1547 528
rect 1591 524 1595 528
rect 1647 524 1651 528
rect 1703 524 1707 528
rect 1767 524 1771 528
rect 1839 524 1843 528
rect 1919 524 1923 528
rect 2007 524 2011 528
rect 2071 524 2075 528
rect 2119 521 2123 525
rect 1135 504 1139 508
rect 2119 504 2123 508
rect 1303 496 1307 500
rect 1343 496 1347 500
rect 1383 496 1387 500
rect 1423 496 1427 500
rect 1463 496 1467 500
rect 1503 496 1507 500
rect 1543 496 1547 500
rect 1591 496 1595 500
rect 1647 496 1651 500
rect 1703 496 1707 500
rect 1767 496 1771 500
rect 1839 496 1843 500
rect 1919 496 1923 500
rect 2007 496 2011 500
rect 2071 496 2075 500
rect 135 480 139 484
rect 175 480 179 484
rect 231 480 235 484
rect 295 480 299 484
rect 359 480 363 484
rect 423 480 427 484
rect 479 480 483 484
rect 535 480 539 484
rect 591 480 595 484
rect 639 480 643 484
rect 687 480 691 484
rect 735 480 739 484
rect 791 480 795 484
rect 847 480 851 484
rect 111 472 115 476
rect 1095 472 1099 476
rect 1295 460 1299 464
rect 111 455 115 459
rect 1335 460 1339 464
rect 1375 460 1379 464
rect 1423 460 1427 464
rect 1471 460 1475 464
rect 1527 460 1531 464
rect 1583 460 1587 464
rect 1647 460 1651 464
rect 1719 460 1723 464
rect 1807 460 1811 464
rect 1895 460 1899 464
rect 1991 460 1995 464
rect 2071 460 2075 464
rect 135 452 139 456
rect 175 452 179 456
rect 231 452 235 456
rect 295 452 299 456
rect 359 452 363 456
rect 423 452 427 456
rect 479 452 483 456
rect 535 452 539 456
rect 591 452 595 456
rect 639 452 643 456
rect 687 452 691 456
rect 735 452 739 456
rect 791 452 795 456
rect 847 452 851 456
rect 1095 455 1099 459
rect 1135 452 1139 456
rect 2119 452 2123 456
rect 111 433 115 437
rect 175 436 179 440
rect 215 436 219 440
rect 263 436 267 440
rect 327 436 331 440
rect 391 436 395 440
rect 463 436 467 440
rect 535 436 539 440
rect 607 436 611 440
rect 679 436 683 440
rect 743 436 747 440
rect 807 436 811 440
rect 871 436 875 440
rect 943 436 947 440
rect 1095 433 1099 437
rect 1135 435 1139 439
rect 1295 432 1299 436
rect 1335 432 1339 436
rect 1375 432 1379 436
rect 1423 432 1427 436
rect 1471 432 1475 436
rect 1527 432 1531 436
rect 1583 432 1587 436
rect 1647 432 1651 436
rect 1719 432 1723 436
rect 1807 432 1811 436
rect 1895 432 1899 436
rect 1991 432 1995 436
rect 2071 432 2075 436
rect 2119 435 2123 439
rect 111 416 115 420
rect 1095 416 1099 420
rect 1135 417 1139 421
rect 1159 420 1163 424
rect 1199 420 1203 424
rect 1255 420 1259 424
rect 1335 420 1339 424
rect 1415 420 1419 424
rect 1503 420 1507 424
rect 1591 420 1595 424
rect 1671 420 1675 424
rect 1751 420 1755 424
rect 1831 420 1835 424
rect 1911 420 1915 424
rect 1999 420 2003 424
rect 2071 420 2075 424
rect 2119 417 2123 421
rect 175 408 179 412
rect 215 408 219 412
rect 263 408 267 412
rect 327 408 331 412
rect 391 408 395 412
rect 463 408 467 412
rect 535 408 539 412
rect 607 408 611 412
rect 679 408 683 412
rect 743 408 747 412
rect 807 408 811 412
rect 871 408 875 412
rect 943 408 947 412
rect 1135 400 1139 404
rect 2119 400 2123 404
rect 1159 392 1163 396
rect 1199 392 1203 396
rect 1255 392 1259 396
rect 1335 392 1339 396
rect 1415 392 1419 396
rect 1503 392 1507 396
rect 1591 392 1595 396
rect 1671 392 1675 396
rect 1751 392 1755 396
rect 1831 392 1835 396
rect 1911 392 1915 396
rect 1999 392 2003 396
rect 2071 392 2075 396
rect 175 364 179 368
rect 215 364 219 368
rect 271 364 275 368
rect 335 364 339 368
rect 407 364 411 368
rect 487 364 491 368
rect 567 364 571 368
rect 639 364 643 368
rect 711 364 715 368
rect 775 364 779 368
rect 839 364 843 368
rect 895 364 899 368
rect 951 364 955 368
rect 1007 364 1011 368
rect 1047 364 1051 368
rect 111 356 115 360
rect 1095 356 1099 360
rect 1159 352 1163 356
rect 1247 352 1251 356
rect 1359 352 1363 356
rect 1463 352 1467 356
rect 1559 352 1563 356
rect 1647 352 1651 356
rect 1727 352 1731 356
rect 1799 352 1803 356
rect 1863 352 1867 356
rect 1919 352 1923 356
rect 1975 352 1979 356
rect 2031 352 2035 356
rect 2071 352 2075 356
rect 1135 344 1139 348
rect 111 339 115 343
rect 2119 344 2123 348
rect 175 336 179 340
rect 215 336 219 340
rect 271 336 275 340
rect 335 336 339 340
rect 407 336 411 340
rect 487 336 491 340
rect 567 336 571 340
rect 639 336 643 340
rect 711 336 715 340
rect 775 336 779 340
rect 839 336 843 340
rect 895 336 899 340
rect 951 336 955 340
rect 1007 336 1011 340
rect 1047 336 1051 340
rect 1095 339 1099 343
rect 1135 327 1139 331
rect 111 317 115 321
rect 383 320 387 324
rect 423 320 427 324
rect 463 320 467 324
rect 503 320 507 324
rect 543 320 547 324
rect 591 320 595 324
rect 639 320 643 324
rect 687 320 691 324
rect 735 320 739 324
rect 783 320 787 324
rect 831 320 835 324
rect 879 320 883 324
rect 927 320 931 324
rect 967 320 971 324
rect 1007 320 1011 324
rect 1047 320 1051 324
rect 1159 324 1163 328
rect 1247 324 1251 328
rect 1359 324 1363 328
rect 1463 324 1467 328
rect 1559 324 1563 328
rect 1647 324 1651 328
rect 1727 324 1731 328
rect 1799 324 1803 328
rect 1863 324 1867 328
rect 1919 324 1923 328
rect 1975 324 1979 328
rect 2031 324 2035 328
rect 2071 324 2075 328
rect 2119 327 2123 331
rect 1095 317 1099 321
rect 111 300 115 304
rect 1095 300 1099 304
rect 1135 301 1139 305
rect 1351 304 1355 308
rect 1391 304 1395 308
rect 1431 304 1435 308
rect 1471 304 1475 308
rect 1511 304 1515 308
rect 1559 304 1563 308
rect 1615 304 1619 308
rect 1671 304 1675 308
rect 1735 304 1739 308
rect 1807 304 1811 308
rect 1887 304 1891 308
rect 1967 304 1971 308
rect 2047 304 2051 308
rect 2119 301 2123 305
rect 383 292 387 296
rect 423 292 427 296
rect 463 292 467 296
rect 503 292 507 296
rect 543 292 547 296
rect 591 292 595 296
rect 639 292 643 296
rect 687 292 691 296
rect 735 292 739 296
rect 783 292 787 296
rect 831 292 835 296
rect 879 292 883 296
rect 927 292 931 296
rect 967 292 971 296
rect 1007 292 1011 296
rect 1047 292 1051 296
rect 1135 284 1139 288
rect 2119 284 2123 288
rect 1351 276 1355 280
rect 1391 276 1395 280
rect 1431 276 1435 280
rect 1471 276 1475 280
rect 1511 276 1515 280
rect 1559 276 1563 280
rect 1615 276 1619 280
rect 1671 276 1675 280
rect 1735 276 1739 280
rect 1807 276 1811 280
rect 1887 276 1891 280
rect 1967 276 1971 280
rect 2047 276 2051 280
rect 287 248 291 252
rect 327 248 331 252
rect 367 248 371 252
rect 415 248 419 252
rect 471 248 475 252
rect 535 248 539 252
rect 607 248 611 252
rect 679 248 683 252
rect 743 248 747 252
rect 807 248 811 252
rect 863 248 867 252
rect 927 248 931 252
rect 991 248 995 252
rect 1047 248 1051 252
rect 111 240 115 244
rect 1095 240 1099 244
rect 1263 240 1267 244
rect 1303 240 1307 244
rect 1343 240 1347 244
rect 1383 240 1387 244
rect 1423 240 1427 244
rect 1463 240 1467 244
rect 1503 240 1507 244
rect 1543 240 1547 244
rect 1599 240 1603 244
rect 1671 240 1675 244
rect 1759 240 1763 244
rect 1863 240 1867 244
rect 1975 240 1979 244
rect 2071 240 2075 244
rect 1135 232 1139 236
rect 2119 232 2123 236
rect 111 223 115 227
rect 287 220 291 224
rect 327 220 331 224
rect 367 220 371 224
rect 415 220 419 224
rect 471 220 475 224
rect 535 220 539 224
rect 607 220 611 224
rect 679 220 683 224
rect 743 220 747 224
rect 807 220 811 224
rect 863 220 867 224
rect 927 220 931 224
rect 991 220 995 224
rect 1047 220 1051 224
rect 1095 223 1099 227
rect 1135 215 1139 219
rect 1263 212 1267 216
rect 1303 212 1307 216
rect 1343 212 1347 216
rect 1383 212 1387 216
rect 1423 212 1427 216
rect 1463 212 1467 216
rect 1503 212 1507 216
rect 1543 212 1547 216
rect 1599 212 1603 216
rect 1671 212 1675 216
rect 1759 212 1763 216
rect 1863 212 1867 216
rect 1975 212 1979 216
rect 2071 212 2075 216
rect 2119 215 2123 219
rect 111 193 115 197
rect 167 196 171 200
rect 207 196 211 200
rect 247 196 251 200
rect 295 196 299 200
rect 343 196 347 200
rect 399 196 403 200
rect 463 196 467 200
rect 527 196 531 200
rect 599 196 603 200
rect 671 196 675 200
rect 751 196 755 200
rect 831 196 835 200
rect 911 196 915 200
rect 991 196 995 200
rect 1047 196 1051 200
rect 1095 193 1099 197
rect 1135 193 1139 197
rect 1183 196 1187 200
rect 1231 196 1235 200
rect 1295 196 1299 200
rect 1359 196 1363 200
rect 1431 196 1435 200
rect 1511 196 1515 200
rect 1591 196 1595 200
rect 1663 196 1667 200
rect 1735 196 1739 200
rect 1807 196 1811 200
rect 1879 196 1883 200
rect 1951 196 1955 200
rect 2023 196 2027 200
rect 2071 196 2075 200
rect 2119 193 2123 197
rect 111 176 115 180
rect 1095 176 1099 180
rect 1135 176 1139 180
rect 2119 176 2123 180
rect 167 168 171 172
rect 207 168 211 172
rect 247 168 251 172
rect 295 168 299 172
rect 343 168 347 172
rect 399 168 403 172
rect 463 168 467 172
rect 527 168 531 172
rect 599 168 603 172
rect 671 168 675 172
rect 751 168 755 172
rect 831 168 835 172
rect 911 168 915 172
rect 991 168 995 172
rect 1047 168 1051 172
rect 1183 168 1187 172
rect 1231 168 1235 172
rect 1295 168 1299 172
rect 1359 168 1363 172
rect 1431 168 1435 172
rect 1511 168 1515 172
rect 1591 168 1595 172
rect 1663 168 1667 172
rect 1735 168 1739 172
rect 1807 168 1811 172
rect 1879 168 1883 172
rect 1951 168 1955 172
rect 2023 168 2027 172
rect 2071 168 2075 172
rect 135 116 139 120
rect 175 116 179 120
rect 215 116 219 120
rect 255 116 259 120
rect 295 116 299 120
rect 335 116 339 120
rect 375 116 379 120
rect 415 116 419 120
rect 455 116 459 120
rect 495 116 499 120
rect 535 116 539 120
rect 575 116 579 120
rect 615 116 619 120
rect 655 116 659 120
rect 695 116 699 120
rect 735 116 739 120
rect 775 116 779 120
rect 815 116 819 120
rect 871 116 875 120
rect 935 116 939 120
rect 999 116 1003 120
rect 1047 116 1051 120
rect 111 108 115 112
rect 1095 108 1099 112
rect 1159 108 1163 112
rect 1199 108 1203 112
rect 1239 108 1243 112
rect 1279 108 1283 112
rect 1319 108 1323 112
rect 1367 108 1371 112
rect 1431 108 1435 112
rect 1495 108 1499 112
rect 1559 108 1563 112
rect 1615 108 1619 112
rect 1671 108 1675 112
rect 1719 108 1723 112
rect 1767 108 1771 112
rect 1807 108 1811 112
rect 1855 108 1859 112
rect 1903 108 1907 112
rect 1951 108 1955 112
rect 1991 108 1995 112
rect 2031 108 2035 112
rect 2071 108 2075 112
rect 1135 100 1139 104
rect 2119 100 2123 104
rect 111 91 115 95
rect 135 88 139 92
rect 175 88 179 92
rect 215 88 219 92
rect 255 88 259 92
rect 295 88 299 92
rect 335 88 339 92
rect 375 88 379 92
rect 415 88 419 92
rect 455 88 459 92
rect 495 88 499 92
rect 535 88 539 92
rect 575 88 579 92
rect 615 88 619 92
rect 655 88 659 92
rect 695 88 699 92
rect 735 88 739 92
rect 775 88 779 92
rect 815 88 819 92
rect 871 88 875 92
rect 935 88 939 92
rect 999 88 1003 92
rect 1047 88 1051 92
rect 1095 91 1099 95
rect 1135 83 1139 87
rect 1159 80 1163 84
rect 1199 80 1203 84
rect 1239 80 1243 84
rect 1279 80 1283 84
rect 1319 80 1323 84
rect 1367 80 1371 84
rect 1431 80 1435 84
rect 1495 80 1499 84
rect 1559 80 1563 84
rect 1615 80 1619 84
rect 1671 80 1675 84
rect 1719 80 1723 84
rect 1767 80 1771 84
rect 1807 80 1811 84
rect 1855 80 1859 84
rect 1903 80 1907 84
rect 1951 80 1955 84
rect 1991 80 1995 84
rect 2031 80 2035 84
rect 2071 80 2075 84
rect 2119 83 2123 87
<< m3 >>
rect 1135 2214 1139 2215
rect 1135 2209 1139 2210
rect 1343 2214 1347 2215
rect 1343 2209 1347 2210
rect 1383 2214 1387 2215
rect 1383 2209 1387 2210
rect 1423 2214 1427 2215
rect 1423 2209 1427 2210
rect 1463 2214 1467 2215
rect 1463 2209 1467 2210
rect 1503 2214 1507 2215
rect 1503 2209 1507 2210
rect 1543 2214 1547 2215
rect 1543 2209 1547 2210
rect 1583 2214 1587 2215
rect 1583 2209 1587 2210
rect 1623 2214 1627 2215
rect 1623 2209 1627 2210
rect 1663 2214 1667 2215
rect 1663 2209 1667 2210
rect 1703 2214 1707 2215
rect 1703 2209 1707 2210
rect 1743 2214 1747 2215
rect 1743 2209 1747 2210
rect 1783 2214 1787 2215
rect 1783 2209 1787 2210
rect 1823 2214 1827 2215
rect 1823 2209 1827 2210
rect 2119 2214 2123 2215
rect 2119 2209 2123 2210
rect 1136 2189 1138 2209
rect 1344 2197 1346 2209
rect 1384 2197 1386 2209
rect 1424 2197 1426 2209
rect 1464 2197 1466 2209
rect 1504 2197 1506 2209
rect 1544 2197 1546 2209
rect 1584 2197 1586 2209
rect 1624 2197 1626 2209
rect 1664 2197 1666 2209
rect 1704 2197 1706 2209
rect 1744 2197 1746 2209
rect 1784 2197 1786 2209
rect 1824 2197 1826 2209
rect 1342 2196 1348 2197
rect 1342 2192 1343 2196
rect 1347 2192 1348 2196
rect 1342 2191 1348 2192
rect 1382 2196 1388 2197
rect 1382 2192 1383 2196
rect 1387 2192 1388 2196
rect 1382 2191 1388 2192
rect 1422 2196 1428 2197
rect 1422 2192 1423 2196
rect 1427 2192 1428 2196
rect 1422 2191 1428 2192
rect 1462 2196 1468 2197
rect 1462 2192 1463 2196
rect 1467 2192 1468 2196
rect 1462 2191 1468 2192
rect 1502 2196 1508 2197
rect 1502 2192 1503 2196
rect 1507 2192 1508 2196
rect 1502 2191 1508 2192
rect 1542 2196 1548 2197
rect 1542 2192 1543 2196
rect 1547 2192 1548 2196
rect 1542 2191 1548 2192
rect 1582 2196 1588 2197
rect 1582 2192 1583 2196
rect 1587 2192 1588 2196
rect 1582 2191 1588 2192
rect 1622 2196 1628 2197
rect 1622 2192 1623 2196
rect 1627 2192 1628 2196
rect 1622 2191 1628 2192
rect 1662 2196 1668 2197
rect 1662 2192 1663 2196
rect 1667 2192 1668 2196
rect 1662 2191 1668 2192
rect 1702 2196 1708 2197
rect 1702 2192 1703 2196
rect 1707 2192 1708 2196
rect 1702 2191 1708 2192
rect 1742 2196 1748 2197
rect 1742 2192 1743 2196
rect 1747 2192 1748 2196
rect 1742 2191 1748 2192
rect 1782 2196 1788 2197
rect 1782 2192 1783 2196
rect 1787 2192 1788 2196
rect 1782 2191 1788 2192
rect 1822 2196 1828 2197
rect 1822 2192 1823 2196
rect 1827 2192 1828 2196
rect 1822 2191 1828 2192
rect 2120 2189 2122 2209
rect 1134 2188 1140 2189
rect 1134 2184 1135 2188
rect 1139 2184 1140 2188
rect 1134 2183 1140 2184
rect 2118 2188 2124 2189
rect 2118 2184 2119 2188
rect 2123 2184 2124 2188
rect 2118 2183 2124 2184
rect 1134 2171 1140 2172
rect 1134 2167 1135 2171
rect 1139 2167 1140 2171
rect 2118 2171 2124 2172
rect 1134 2166 1140 2167
rect 1342 2168 1348 2169
rect 1136 2163 1138 2166
rect 1342 2164 1343 2168
rect 1347 2164 1348 2168
rect 1342 2163 1348 2164
rect 1382 2168 1388 2169
rect 1382 2164 1383 2168
rect 1387 2164 1388 2168
rect 1382 2163 1388 2164
rect 1422 2168 1428 2169
rect 1422 2164 1423 2168
rect 1427 2164 1428 2168
rect 1422 2163 1428 2164
rect 1462 2168 1468 2169
rect 1462 2164 1463 2168
rect 1467 2164 1468 2168
rect 1462 2163 1468 2164
rect 1502 2168 1508 2169
rect 1502 2164 1503 2168
rect 1507 2164 1508 2168
rect 1502 2163 1508 2164
rect 1542 2168 1548 2169
rect 1542 2164 1543 2168
rect 1547 2164 1548 2168
rect 1542 2163 1548 2164
rect 1582 2168 1588 2169
rect 1582 2164 1583 2168
rect 1587 2164 1588 2168
rect 1582 2163 1588 2164
rect 1622 2168 1628 2169
rect 1622 2164 1623 2168
rect 1627 2164 1628 2168
rect 1622 2163 1628 2164
rect 1662 2168 1668 2169
rect 1662 2164 1663 2168
rect 1667 2164 1668 2168
rect 1662 2163 1668 2164
rect 1702 2168 1708 2169
rect 1702 2164 1703 2168
rect 1707 2164 1708 2168
rect 1702 2163 1708 2164
rect 1742 2168 1748 2169
rect 1742 2164 1743 2168
rect 1747 2164 1748 2168
rect 1742 2163 1748 2164
rect 1782 2168 1788 2169
rect 1782 2164 1783 2168
rect 1787 2164 1788 2168
rect 1782 2163 1788 2164
rect 1822 2168 1828 2169
rect 1822 2164 1823 2168
rect 1827 2164 1828 2168
rect 2118 2167 2119 2171
rect 2123 2167 2124 2171
rect 2118 2166 2124 2167
rect 1822 2163 1828 2164
rect 2120 2163 2122 2166
rect 1135 2162 1139 2163
rect 1135 2157 1139 2158
rect 1287 2162 1291 2163
rect 1287 2157 1291 2158
rect 1327 2162 1331 2163
rect 1327 2157 1331 2158
rect 1343 2162 1347 2163
rect 1343 2157 1347 2158
rect 1367 2162 1371 2163
rect 1367 2157 1371 2158
rect 1383 2162 1387 2163
rect 1383 2157 1387 2158
rect 1415 2162 1419 2163
rect 1415 2157 1419 2158
rect 1423 2162 1427 2163
rect 1423 2157 1427 2158
rect 1463 2162 1467 2163
rect 1463 2157 1467 2158
rect 1503 2162 1507 2163
rect 1503 2157 1507 2158
rect 1519 2162 1523 2163
rect 1519 2157 1523 2158
rect 1543 2162 1547 2163
rect 1543 2157 1547 2158
rect 1575 2162 1579 2163
rect 1575 2157 1579 2158
rect 1583 2162 1587 2163
rect 1583 2157 1587 2158
rect 1623 2162 1627 2163
rect 1623 2157 1627 2158
rect 1663 2162 1667 2163
rect 1663 2157 1667 2158
rect 1671 2162 1675 2163
rect 1671 2157 1675 2158
rect 1703 2162 1707 2163
rect 1703 2157 1707 2158
rect 1719 2162 1723 2163
rect 1719 2157 1723 2158
rect 1743 2162 1747 2163
rect 1743 2157 1747 2158
rect 1775 2162 1779 2163
rect 1775 2157 1779 2158
rect 1783 2162 1787 2163
rect 1783 2157 1787 2158
rect 1823 2162 1827 2163
rect 1823 2157 1827 2158
rect 1831 2162 1835 2163
rect 1831 2157 1835 2158
rect 1887 2162 1891 2163
rect 1887 2157 1891 2158
rect 2119 2162 2123 2163
rect 2119 2157 2123 2158
rect 1136 2154 1138 2157
rect 1286 2156 1292 2157
rect 1134 2153 1140 2154
rect 1134 2149 1135 2153
rect 1139 2149 1140 2153
rect 1286 2152 1287 2156
rect 1291 2152 1292 2156
rect 1286 2151 1292 2152
rect 1326 2156 1332 2157
rect 1326 2152 1327 2156
rect 1331 2152 1332 2156
rect 1326 2151 1332 2152
rect 1366 2156 1372 2157
rect 1366 2152 1367 2156
rect 1371 2152 1372 2156
rect 1366 2151 1372 2152
rect 1414 2156 1420 2157
rect 1414 2152 1415 2156
rect 1419 2152 1420 2156
rect 1414 2151 1420 2152
rect 1462 2156 1468 2157
rect 1462 2152 1463 2156
rect 1467 2152 1468 2156
rect 1462 2151 1468 2152
rect 1518 2156 1524 2157
rect 1518 2152 1519 2156
rect 1523 2152 1524 2156
rect 1518 2151 1524 2152
rect 1574 2156 1580 2157
rect 1574 2152 1575 2156
rect 1579 2152 1580 2156
rect 1574 2151 1580 2152
rect 1622 2156 1628 2157
rect 1622 2152 1623 2156
rect 1627 2152 1628 2156
rect 1622 2151 1628 2152
rect 1670 2156 1676 2157
rect 1670 2152 1671 2156
rect 1675 2152 1676 2156
rect 1670 2151 1676 2152
rect 1718 2156 1724 2157
rect 1718 2152 1719 2156
rect 1723 2152 1724 2156
rect 1718 2151 1724 2152
rect 1774 2156 1780 2157
rect 1774 2152 1775 2156
rect 1779 2152 1780 2156
rect 1774 2151 1780 2152
rect 1830 2156 1836 2157
rect 1830 2152 1831 2156
rect 1835 2152 1836 2156
rect 1830 2151 1836 2152
rect 1886 2156 1892 2157
rect 1886 2152 1887 2156
rect 1891 2152 1892 2156
rect 2120 2154 2122 2157
rect 1886 2151 1892 2152
rect 2118 2153 2124 2154
rect 1134 2148 1140 2149
rect 2118 2149 2119 2153
rect 2123 2149 2124 2153
rect 2118 2148 2124 2149
rect 1134 2136 1140 2137
rect 1134 2132 1135 2136
rect 1139 2132 1140 2136
rect 1134 2131 1140 2132
rect 2118 2136 2124 2137
rect 2118 2132 2119 2136
rect 2123 2132 2124 2136
rect 2118 2131 2124 2132
rect 1136 2107 1138 2131
rect 1286 2128 1292 2129
rect 1286 2124 1287 2128
rect 1291 2124 1292 2128
rect 1286 2123 1292 2124
rect 1326 2128 1332 2129
rect 1326 2124 1327 2128
rect 1331 2124 1332 2128
rect 1326 2123 1332 2124
rect 1366 2128 1372 2129
rect 1366 2124 1367 2128
rect 1371 2124 1372 2128
rect 1366 2123 1372 2124
rect 1414 2128 1420 2129
rect 1414 2124 1415 2128
rect 1419 2124 1420 2128
rect 1414 2123 1420 2124
rect 1462 2128 1468 2129
rect 1462 2124 1463 2128
rect 1467 2124 1468 2128
rect 1462 2123 1468 2124
rect 1518 2128 1524 2129
rect 1518 2124 1519 2128
rect 1523 2124 1524 2128
rect 1518 2123 1524 2124
rect 1574 2128 1580 2129
rect 1574 2124 1575 2128
rect 1579 2124 1580 2128
rect 1574 2123 1580 2124
rect 1622 2128 1628 2129
rect 1622 2124 1623 2128
rect 1627 2124 1628 2128
rect 1622 2123 1628 2124
rect 1670 2128 1676 2129
rect 1670 2124 1671 2128
rect 1675 2124 1676 2128
rect 1670 2123 1676 2124
rect 1718 2128 1724 2129
rect 1718 2124 1719 2128
rect 1723 2124 1724 2128
rect 1718 2123 1724 2124
rect 1774 2128 1780 2129
rect 1774 2124 1775 2128
rect 1779 2124 1780 2128
rect 1774 2123 1780 2124
rect 1830 2128 1836 2129
rect 1830 2124 1831 2128
rect 1835 2124 1836 2128
rect 1830 2123 1836 2124
rect 1886 2128 1892 2129
rect 1886 2124 1887 2128
rect 1891 2124 1892 2128
rect 1886 2123 1892 2124
rect 1288 2107 1290 2123
rect 1328 2107 1330 2123
rect 1368 2107 1370 2123
rect 1416 2107 1418 2123
rect 1464 2107 1466 2123
rect 1520 2107 1522 2123
rect 1576 2107 1578 2123
rect 1624 2107 1626 2123
rect 1672 2107 1674 2123
rect 1720 2107 1722 2123
rect 1776 2107 1778 2123
rect 1832 2107 1834 2123
rect 1888 2107 1890 2123
rect 2120 2107 2122 2131
rect 1135 2106 1139 2107
rect 1135 2101 1139 2102
rect 1223 2106 1227 2107
rect 1223 2101 1227 2102
rect 1279 2106 1283 2107
rect 1279 2101 1283 2102
rect 1287 2106 1291 2107
rect 1287 2101 1291 2102
rect 1327 2106 1331 2107
rect 1327 2101 1331 2102
rect 1343 2106 1347 2107
rect 1343 2101 1347 2102
rect 1367 2106 1371 2107
rect 1367 2101 1371 2102
rect 1415 2106 1419 2107
rect 1415 2101 1419 2102
rect 1423 2106 1427 2107
rect 1423 2101 1427 2102
rect 1463 2106 1467 2107
rect 1463 2101 1467 2102
rect 1503 2106 1507 2107
rect 1503 2101 1507 2102
rect 1519 2106 1523 2107
rect 1519 2101 1523 2102
rect 1575 2106 1579 2107
rect 1575 2101 1579 2102
rect 1583 2106 1587 2107
rect 1583 2101 1587 2102
rect 1623 2106 1627 2107
rect 1623 2101 1627 2102
rect 1663 2106 1667 2107
rect 1663 2101 1667 2102
rect 1671 2106 1675 2107
rect 1671 2101 1675 2102
rect 1719 2106 1723 2107
rect 1719 2101 1723 2102
rect 1743 2106 1747 2107
rect 1743 2101 1747 2102
rect 1775 2106 1779 2107
rect 1775 2101 1779 2102
rect 1831 2106 1835 2107
rect 1831 2101 1835 2102
rect 1887 2106 1891 2107
rect 1887 2101 1891 2102
rect 1919 2106 1923 2107
rect 1919 2101 1923 2102
rect 2007 2106 2011 2107
rect 2007 2101 2011 2102
rect 2071 2106 2075 2107
rect 2071 2101 2075 2102
rect 2119 2106 2123 2107
rect 2119 2101 2123 2102
rect 1136 2081 1138 2101
rect 1224 2089 1226 2101
rect 1280 2089 1282 2101
rect 1344 2089 1346 2101
rect 1424 2089 1426 2101
rect 1504 2089 1506 2101
rect 1584 2089 1586 2101
rect 1664 2089 1666 2101
rect 1744 2089 1746 2101
rect 1832 2089 1834 2101
rect 1920 2089 1922 2101
rect 2008 2089 2010 2101
rect 2072 2089 2074 2101
rect 1222 2088 1228 2089
rect 1222 2084 1223 2088
rect 1227 2084 1228 2088
rect 1222 2083 1228 2084
rect 1278 2088 1284 2089
rect 1278 2084 1279 2088
rect 1283 2084 1284 2088
rect 1278 2083 1284 2084
rect 1342 2088 1348 2089
rect 1342 2084 1343 2088
rect 1347 2084 1348 2088
rect 1342 2083 1348 2084
rect 1422 2088 1428 2089
rect 1422 2084 1423 2088
rect 1427 2084 1428 2088
rect 1422 2083 1428 2084
rect 1502 2088 1508 2089
rect 1502 2084 1503 2088
rect 1507 2084 1508 2088
rect 1502 2083 1508 2084
rect 1582 2088 1588 2089
rect 1582 2084 1583 2088
rect 1587 2084 1588 2088
rect 1582 2083 1588 2084
rect 1662 2088 1668 2089
rect 1662 2084 1663 2088
rect 1667 2084 1668 2088
rect 1662 2083 1668 2084
rect 1742 2088 1748 2089
rect 1742 2084 1743 2088
rect 1747 2084 1748 2088
rect 1742 2083 1748 2084
rect 1830 2088 1836 2089
rect 1830 2084 1831 2088
rect 1835 2084 1836 2088
rect 1830 2083 1836 2084
rect 1918 2088 1924 2089
rect 1918 2084 1919 2088
rect 1923 2084 1924 2088
rect 1918 2083 1924 2084
rect 2006 2088 2012 2089
rect 2006 2084 2007 2088
rect 2011 2084 2012 2088
rect 2006 2083 2012 2084
rect 2070 2088 2076 2089
rect 2070 2084 2071 2088
rect 2075 2084 2076 2088
rect 2070 2083 2076 2084
rect 2120 2081 2122 2101
rect 1134 2080 1140 2081
rect 1134 2076 1135 2080
rect 1139 2076 1140 2080
rect 1134 2075 1140 2076
rect 2118 2080 2124 2081
rect 2118 2076 2119 2080
rect 2123 2076 2124 2080
rect 2118 2075 2124 2076
rect 1134 2063 1140 2064
rect 1134 2059 1135 2063
rect 1139 2059 1140 2063
rect 2118 2063 2124 2064
rect 1134 2058 1140 2059
rect 1222 2060 1228 2061
rect 1136 2055 1138 2058
rect 1222 2056 1223 2060
rect 1227 2056 1228 2060
rect 1222 2055 1228 2056
rect 1278 2060 1284 2061
rect 1278 2056 1279 2060
rect 1283 2056 1284 2060
rect 1278 2055 1284 2056
rect 1342 2060 1348 2061
rect 1342 2056 1343 2060
rect 1347 2056 1348 2060
rect 1342 2055 1348 2056
rect 1422 2060 1428 2061
rect 1422 2056 1423 2060
rect 1427 2056 1428 2060
rect 1422 2055 1428 2056
rect 1502 2060 1508 2061
rect 1502 2056 1503 2060
rect 1507 2056 1508 2060
rect 1502 2055 1508 2056
rect 1582 2060 1588 2061
rect 1582 2056 1583 2060
rect 1587 2056 1588 2060
rect 1582 2055 1588 2056
rect 1662 2060 1668 2061
rect 1662 2056 1663 2060
rect 1667 2056 1668 2060
rect 1662 2055 1668 2056
rect 1742 2060 1748 2061
rect 1742 2056 1743 2060
rect 1747 2056 1748 2060
rect 1742 2055 1748 2056
rect 1830 2060 1836 2061
rect 1830 2056 1831 2060
rect 1835 2056 1836 2060
rect 1830 2055 1836 2056
rect 1918 2060 1924 2061
rect 1918 2056 1919 2060
rect 1923 2056 1924 2060
rect 1918 2055 1924 2056
rect 2006 2060 2012 2061
rect 2006 2056 2007 2060
rect 2011 2056 2012 2060
rect 2006 2055 2012 2056
rect 2070 2060 2076 2061
rect 2070 2056 2071 2060
rect 2075 2056 2076 2060
rect 2118 2059 2119 2063
rect 2123 2059 2124 2063
rect 2118 2058 2124 2059
rect 2070 2055 2076 2056
rect 2120 2055 2122 2058
rect 1135 2054 1139 2055
rect 1135 2049 1139 2050
rect 1183 2054 1187 2055
rect 1183 2049 1187 2050
rect 1223 2054 1227 2055
rect 1223 2049 1227 2050
rect 1239 2054 1243 2055
rect 1239 2049 1243 2050
rect 1279 2054 1283 2055
rect 1279 2049 1283 2050
rect 1311 2054 1315 2055
rect 1311 2049 1315 2050
rect 1343 2054 1347 2055
rect 1343 2049 1347 2050
rect 1399 2054 1403 2055
rect 1399 2049 1403 2050
rect 1423 2054 1427 2055
rect 1423 2049 1427 2050
rect 1487 2054 1491 2055
rect 1487 2049 1491 2050
rect 1503 2054 1507 2055
rect 1503 2049 1507 2050
rect 1583 2054 1587 2055
rect 1583 2049 1587 2050
rect 1663 2054 1667 2055
rect 1663 2049 1667 2050
rect 1671 2054 1675 2055
rect 1671 2049 1675 2050
rect 1743 2054 1747 2055
rect 1743 2049 1747 2050
rect 1759 2054 1763 2055
rect 1759 2049 1763 2050
rect 1831 2054 1835 2055
rect 1831 2049 1835 2050
rect 1839 2054 1843 2055
rect 1839 2049 1843 2050
rect 1919 2054 1923 2055
rect 1919 2049 1923 2050
rect 2007 2054 2011 2055
rect 2007 2049 2011 2050
rect 2071 2054 2075 2055
rect 2071 2049 2075 2050
rect 2119 2054 2123 2055
rect 2119 2049 2123 2050
rect 1136 2046 1138 2049
rect 1182 2048 1188 2049
rect 1134 2045 1140 2046
rect 1134 2041 1135 2045
rect 1139 2041 1140 2045
rect 1182 2044 1183 2048
rect 1187 2044 1188 2048
rect 1182 2043 1188 2044
rect 1238 2048 1244 2049
rect 1238 2044 1239 2048
rect 1243 2044 1244 2048
rect 1238 2043 1244 2044
rect 1310 2048 1316 2049
rect 1310 2044 1311 2048
rect 1315 2044 1316 2048
rect 1310 2043 1316 2044
rect 1398 2048 1404 2049
rect 1398 2044 1399 2048
rect 1403 2044 1404 2048
rect 1398 2043 1404 2044
rect 1486 2048 1492 2049
rect 1486 2044 1487 2048
rect 1491 2044 1492 2048
rect 1486 2043 1492 2044
rect 1582 2048 1588 2049
rect 1582 2044 1583 2048
rect 1587 2044 1588 2048
rect 1582 2043 1588 2044
rect 1670 2048 1676 2049
rect 1670 2044 1671 2048
rect 1675 2044 1676 2048
rect 1670 2043 1676 2044
rect 1758 2048 1764 2049
rect 1758 2044 1759 2048
rect 1763 2044 1764 2048
rect 1758 2043 1764 2044
rect 1838 2048 1844 2049
rect 1838 2044 1839 2048
rect 1843 2044 1844 2048
rect 1838 2043 1844 2044
rect 1918 2048 1924 2049
rect 1918 2044 1919 2048
rect 1923 2044 1924 2048
rect 1918 2043 1924 2044
rect 2006 2048 2012 2049
rect 2006 2044 2007 2048
rect 2011 2044 2012 2048
rect 2006 2043 2012 2044
rect 2070 2048 2076 2049
rect 2070 2044 2071 2048
rect 2075 2044 2076 2048
rect 2120 2046 2122 2049
rect 2070 2043 2076 2044
rect 2118 2045 2124 2046
rect 1134 2040 1140 2041
rect 2118 2041 2119 2045
rect 2123 2041 2124 2045
rect 2118 2040 2124 2041
rect 111 2034 115 2035
rect 111 2029 115 2030
rect 191 2034 195 2035
rect 191 2029 195 2030
rect 231 2034 235 2035
rect 231 2029 235 2030
rect 287 2034 291 2035
rect 287 2029 291 2030
rect 351 2034 355 2035
rect 351 2029 355 2030
rect 423 2034 427 2035
rect 423 2029 427 2030
rect 495 2034 499 2035
rect 495 2029 499 2030
rect 575 2034 579 2035
rect 575 2029 579 2030
rect 647 2034 651 2035
rect 647 2029 651 2030
rect 719 2034 723 2035
rect 719 2029 723 2030
rect 783 2034 787 2035
rect 783 2029 787 2030
rect 839 2034 843 2035
rect 839 2029 843 2030
rect 895 2034 899 2035
rect 895 2029 899 2030
rect 951 2034 955 2035
rect 951 2029 955 2030
rect 1007 2034 1011 2035
rect 1007 2029 1011 2030
rect 1047 2034 1051 2035
rect 1047 2029 1051 2030
rect 1095 2034 1099 2035
rect 1095 2029 1099 2030
rect 112 2009 114 2029
rect 192 2017 194 2029
rect 232 2017 234 2029
rect 288 2017 290 2029
rect 352 2017 354 2029
rect 424 2017 426 2029
rect 496 2017 498 2029
rect 576 2017 578 2029
rect 648 2017 650 2029
rect 720 2017 722 2029
rect 784 2017 786 2029
rect 840 2017 842 2029
rect 896 2017 898 2029
rect 952 2017 954 2029
rect 1008 2017 1010 2029
rect 1048 2017 1050 2029
rect 190 2016 196 2017
rect 190 2012 191 2016
rect 195 2012 196 2016
rect 190 2011 196 2012
rect 230 2016 236 2017
rect 230 2012 231 2016
rect 235 2012 236 2016
rect 230 2011 236 2012
rect 286 2016 292 2017
rect 286 2012 287 2016
rect 291 2012 292 2016
rect 286 2011 292 2012
rect 350 2016 356 2017
rect 350 2012 351 2016
rect 355 2012 356 2016
rect 350 2011 356 2012
rect 422 2016 428 2017
rect 422 2012 423 2016
rect 427 2012 428 2016
rect 422 2011 428 2012
rect 494 2016 500 2017
rect 494 2012 495 2016
rect 499 2012 500 2016
rect 494 2011 500 2012
rect 574 2016 580 2017
rect 574 2012 575 2016
rect 579 2012 580 2016
rect 574 2011 580 2012
rect 646 2016 652 2017
rect 646 2012 647 2016
rect 651 2012 652 2016
rect 646 2011 652 2012
rect 718 2016 724 2017
rect 718 2012 719 2016
rect 723 2012 724 2016
rect 718 2011 724 2012
rect 782 2016 788 2017
rect 782 2012 783 2016
rect 787 2012 788 2016
rect 782 2011 788 2012
rect 838 2016 844 2017
rect 838 2012 839 2016
rect 843 2012 844 2016
rect 838 2011 844 2012
rect 894 2016 900 2017
rect 894 2012 895 2016
rect 899 2012 900 2016
rect 894 2011 900 2012
rect 950 2016 956 2017
rect 950 2012 951 2016
rect 955 2012 956 2016
rect 950 2011 956 2012
rect 1006 2016 1012 2017
rect 1006 2012 1007 2016
rect 1011 2012 1012 2016
rect 1006 2011 1012 2012
rect 1046 2016 1052 2017
rect 1046 2012 1047 2016
rect 1051 2012 1052 2016
rect 1046 2011 1052 2012
rect 1096 2009 1098 2029
rect 1134 2028 1140 2029
rect 1134 2024 1135 2028
rect 1139 2024 1140 2028
rect 1134 2023 1140 2024
rect 2118 2028 2124 2029
rect 2118 2024 2119 2028
rect 2123 2024 2124 2028
rect 2118 2023 2124 2024
rect 110 2008 116 2009
rect 110 2004 111 2008
rect 115 2004 116 2008
rect 110 2003 116 2004
rect 1094 2008 1100 2009
rect 1094 2004 1095 2008
rect 1099 2004 1100 2008
rect 1094 2003 1100 2004
rect 1136 2003 1138 2023
rect 1182 2020 1188 2021
rect 1182 2016 1183 2020
rect 1187 2016 1188 2020
rect 1182 2015 1188 2016
rect 1238 2020 1244 2021
rect 1238 2016 1239 2020
rect 1243 2016 1244 2020
rect 1238 2015 1244 2016
rect 1310 2020 1316 2021
rect 1310 2016 1311 2020
rect 1315 2016 1316 2020
rect 1310 2015 1316 2016
rect 1398 2020 1404 2021
rect 1398 2016 1399 2020
rect 1403 2016 1404 2020
rect 1398 2015 1404 2016
rect 1486 2020 1492 2021
rect 1486 2016 1487 2020
rect 1491 2016 1492 2020
rect 1486 2015 1492 2016
rect 1582 2020 1588 2021
rect 1582 2016 1583 2020
rect 1587 2016 1588 2020
rect 1582 2015 1588 2016
rect 1670 2020 1676 2021
rect 1670 2016 1671 2020
rect 1675 2016 1676 2020
rect 1670 2015 1676 2016
rect 1758 2020 1764 2021
rect 1758 2016 1759 2020
rect 1763 2016 1764 2020
rect 1758 2015 1764 2016
rect 1838 2020 1844 2021
rect 1838 2016 1839 2020
rect 1843 2016 1844 2020
rect 1838 2015 1844 2016
rect 1918 2020 1924 2021
rect 1918 2016 1919 2020
rect 1923 2016 1924 2020
rect 1918 2015 1924 2016
rect 2006 2020 2012 2021
rect 2006 2016 2007 2020
rect 2011 2016 2012 2020
rect 2006 2015 2012 2016
rect 2070 2020 2076 2021
rect 2070 2016 2071 2020
rect 2075 2016 2076 2020
rect 2070 2015 2076 2016
rect 1184 2003 1186 2015
rect 1240 2003 1242 2015
rect 1312 2003 1314 2015
rect 1400 2003 1402 2015
rect 1488 2003 1490 2015
rect 1584 2003 1586 2015
rect 1672 2003 1674 2015
rect 1760 2003 1762 2015
rect 1840 2003 1842 2015
rect 1920 2003 1922 2015
rect 2008 2003 2010 2015
rect 2072 2003 2074 2015
rect 2120 2003 2122 2023
rect 1135 2002 1139 2003
rect 1135 1997 1139 1998
rect 1183 2002 1187 2003
rect 1183 1997 1187 1998
rect 1239 2002 1243 2003
rect 1239 1997 1243 1998
rect 1303 2002 1307 2003
rect 1303 1997 1307 1998
rect 1311 2002 1315 2003
rect 1311 1997 1315 1998
rect 1383 2002 1387 2003
rect 1383 1997 1387 1998
rect 1399 2002 1403 2003
rect 1399 1997 1403 1998
rect 1463 2002 1467 2003
rect 1463 1997 1467 1998
rect 1487 2002 1491 2003
rect 1487 1997 1491 1998
rect 1543 2002 1547 2003
rect 1543 1997 1547 1998
rect 1583 2002 1587 2003
rect 1583 1997 1587 1998
rect 1615 2002 1619 2003
rect 1615 1997 1619 1998
rect 1671 2002 1675 2003
rect 1671 1997 1675 1998
rect 1687 2002 1691 2003
rect 1687 1997 1691 1998
rect 1751 2002 1755 2003
rect 1751 1997 1755 1998
rect 1759 2002 1763 2003
rect 1759 1997 1763 1998
rect 1815 2002 1819 2003
rect 1815 1997 1819 1998
rect 1839 2002 1843 2003
rect 1839 1997 1843 1998
rect 1879 2002 1883 2003
rect 1879 1997 1883 1998
rect 1919 2002 1923 2003
rect 1919 1997 1923 1998
rect 1951 2002 1955 2003
rect 1951 1997 1955 1998
rect 2007 2002 2011 2003
rect 2007 1997 2011 1998
rect 2023 2002 2027 2003
rect 2023 1997 2027 1998
rect 2071 2002 2075 2003
rect 2071 1997 2075 1998
rect 2119 2002 2123 2003
rect 2119 1997 2123 1998
rect 110 1991 116 1992
rect 110 1987 111 1991
rect 115 1987 116 1991
rect 1094 1991 1100 1992
rect 110 1986 116 1987
rect 190 1988 196 1989
rect 112 1983 114 1986
rect 190 1984 191 1988
rect 195 1984 196 1988
rect 190 1983 196 1984
rect 230 1988 236 1989
rect 230 1984 231 1988
rect 235 1984 236 1988
rect 230 1983 236 1984
rect 286 1988 292 1989
rect 286 1984 287 1988
rect 291 1984 292 1988
rect 286 1983 292 1984
rect 350 1988 356 1989
rect 350 1984 351 1988
rect 355 1984 356 1988
rect 350 1983 356 1984
rect 422 1988 428 1989
rect 422 1984 423 1988
rect 427 1984 428 1988
rect 422 1983 428 1984
rect 494 1988 500 1989
rect 494 1984 495 1988
rect 499 1984 500 1988
rect 494 1983 500 1984
rect 574 1988 580 1989
rect 574 1984 575 1988
rect 579 1984 580 1988
rect 574 1983 580 1984
rect 646 1988 652 1989
rect 646 1984 647 1988
rect 651 1984 652 1988
rect 646 1983 652 1984
rect 718 1988 724 1989
rect 718 1984 719 1988
rect 723 1984 724 1988
rect 718 1983 724 1984
rect 782 1988 788 1989
rect 782 1984 783 1988
rect 787 1984 788 1988
rect 782 1983 788 1984
rect 838 1988 844 1989
rect 838 1984 839 1988
rect 843 1984 844 1988
rect 838 1983 844 1984
rect 894 1988 900 1989
rect 894 1984 895 1988
rect 899 1984 900 1988
rect 894 1983 900 1984
rect 950 1988 956 1989
rect 950 1984 951 1988
rect 955 1984 956 1988
rect 950 1983 956 1984
rect 1006 1988 1012 1989
rect 1006 1984 1007 1988
rect 1011 1984 1012 1988
rect 1006 1983 1012 1984
rect 1046 1988 1052 1989
rect 1046 1984 1047 1988
rect 1051 1984 1052 1988
rect 1094 1987 1095 1991
rect 1099 1987 1100 1991
rect 1094 1986 1100 1987
rect 1046 1983 1052 1984
rect 1096 1983 1098 1986
rect 111 1982 115 1983
rect 111 1977 115 1978
rect 191 1982 195 1983
rect 191 1977 195 1978
rect 231 1982 235 1983
rect 231 1977 235 1978
rect 247 1982 251 1983
rect 247 1977 251 1978
rect 287 1982 291 1983
rect 287 1977 291 1978
rect 311 1982 315 1983
rect 311 1977 315 1978
rect 351 1982 355 1983
rect 351 1977 355 1978
rect 375 1982 379 1983
rect 375 1977 379 1978
rect 423 1982 427 1983
rect 423 1977 427 1978
rect 447 1982 451 1983
rect 447 1977 451 1978
rect 495 1982 499 1983
rect 495 1977 499 1978
rect 519 1982 523 1983
rect 519 1977 523 1978
rect 575 1982 579 1983
rect 575 1977 579 1978
rect 591 1982 595 1983
rect 591 1977 595 1978
rect 647 1982 651 1983
rect 647 1977 651 1978
rect 655 1982 659 1983
rect 655 1977 659 1978
rect 719 1982 723 1983
rect 719 1977 723 1978
rect 775 1982 779 1983
rect 775 1977 779 1978
rect 783 1982 787 1983
rect 783 1977 787 1978
rect 823 1982 827 1983
rect 823 1977 827 1978
rect 839 1982 843 1983
rect 839 1977 843 1978
rect 871 1982 875 1983
rect 871 1977 875 1978
rect 895 1982 899 1983
rect 895 1977 899 1978
rect 919 1982 923 1983
rect 919 1977 923 1978
rect 951 1982 955 1983
rect 951 1977 955 1978
rect 967 1982 971 1983
rect 967 1977 971 1978
rect 1007 1982 1011 1983
rect 1007 1977 1011 1978
rect 1047 1982 1051 1983
rect 1047 1977 1051 1978
rect 1095 1982 1099 1983
rect 1095 1977 1099 1978
rect 1136 1977 1138 1997
rect 1304 1985 1306 1997
rect 1384 1985 1386 1997
rect 1464 1985 1466 1997
rect 1544 1985 1546 1997
rect 1616 1985 1618 1997
rect 1688 1985 1690 1997
rect 1752 1985 1754 1997
rect 1816 1985 1818 1997
rect 1880 1985 1882 1997
rect 1952 1985 1954 1997
rect 2024 1985 2026 1997
rect 2072 1985 2074 1997
rect 1302 1984 1308 1985
rect 1302 1980 1303 1984
rect 1307 1980 1308 1984
rect 1302 1979 1308 1980
rect 1382 1984 1388 1985
rect 1382 1980 1383 1984
rect 1387 1980 1388 1984
rect 1382 1979 1388 1980
rect 1462 1984 1468 1985
rect 1462 1980 1463 1984
rect 1467 1980 1468 1984
rect 1462 1979 1468 1980
rect 1542 1984 1548 1985
rect 1542 1980 1543 1984
rect 1547 1980 1548 1984
rect 1542 1979 1548 1980
rect 1614 1984 1620 1985
rect 1614 1980 1615 1984
rect 1619 1980 1620 1984
rect 1614 1979 1620 1980
rect 1686 1984 1692 1985
rect 1686 1980 1687 1984
rect 1691 1980 1692 1984
rect 1686 1979 1692 1980
rect 1750 1984 1756 1985
rect 1750 1980 1751 1984
rect 1755 1980 1756 1984
rect 1750 1979 1756 1980
rect 1814 1984 1820 1985
rect 1814 1980 1815 1984
rect 1819 1980 1820 1984
rect 1814 1979 1820 1980
rect 1878 1984 1884 1985
rect 1878 1980 1879 1984
rect 1883 1980 1884 1984
rect 1878 1979 1884 1980
rect 1950 1984 1956 1985
rect 1950 1980 1951 1984
rect 1955 1980 1956 1984
rect 1950 1979 1956 1980
rect 2022 1984 2028 1985
rect 2022 1980 2023 1984
rect 2027 1980 2028 1984
rect 2022 1979 2028 1980
rect 2070 1984 2076 1985
rect 2070 1980 2071 1984
rect 2075 1980 2076 1984
rect 2070 1979 2076 1980
rect 2120 1977 2122 1997
rect 112 1974 114 1977
rect 190 1976 196 1977
rect 110 1973 116 1974
rect 110 1969 111 1973
rect 115 1969 116 1973
rect 190 1972 191 1976
rect 195 1972 196 1976
rect 190 1971 196 1972
rect 246 1976 252 1977
rect 246 1972 247 1976
rect 251 1972 252 1976
rect 246 1971 252 1972
rect 310 1976 316 1977
rect 310 1972 311 1976
rect 315 1972 316 1976
rect 310 1971 316 1972
rect 374 1976 380 1977
rect 374 1972 375 1976
rect 379 1972 380 1976
rect 374 1971 380 1972
rect 446 1976 452 1977
rect 446 1972 447 1976
rect 451 1972 452 1976
rect 446 1971 452 1972
rect 518 1976 524 1977
rect 518 1972 519 1976
rect 523 1972 524 1976
rect 518 1971 524 1972
rect 590 1976 596 1977
rect 590 1972 591 1976
rect 595 1972 596 1976
rect 590 1971 596 1972
rect 654 1976 660 1977
rect 654 1972 655 1976
rect 659 1972 660 1976
rect 654 1971 660 1972
rect 718 1976 724 1977
rect 718 1972 719 1976
rect 723 1972 724 1976
rect 718 1971 724 1972
rect 774 1976 780 1977
rect 774 1972 775 1976
rect 779 1972 780 1976
rect 774 1971 780 1972
rect 822 1976 828 1977
rect 822 1972 823 1976
rect 827 1972 828 1976
rect 822 1971 828 1972
rect 870 1976 876 1977
rect 870 1972 871 1976
rect 875 1972 876 1976
rect 870 1971 876 1972
rect 918 1976 924 1977
rect 918 1972 919 1976
rect 923 1972 924 1976
rect 918 1971 924 1972
rect 966 1976 972 1977
rect 966 1972 967 1976
rect 971 1972 972 1976
rect 966 1971 972 1972
rect 1006 1976 1012 1977
rect 1006 1972 1007 1976
rect 1011 1972 1012 1976
rect 1006 1971 1012 1972
rect 1046 1976 1052 1977
rect 1046 1972 1047 1976
rect 1051 1972 1052 1976
rect 1096 1974 1098 1977
rect 1134 1976 1140 1977
rect 1046 1971 1052 1972
rect 1094 1973 1100 1974
rect 110 1968 116 1969
rect 1094 1969 1095 1973
rect 1099 1969 1100 1973
rect 1134 1972 1135 1976
rect 1139 1972 1140 1976
rect 1134 1971 1140 1972
rect 2118 1976 2124 1977
rect 2118 1972 2119 1976
rect 2123 1972 2124 1976
rect 2118 1971 2124 1972
rect 1094 1968 1100 1969
rect 1134 1959 1140 1960
rect 110 1956 116 1957
rect 110 1952 111 1956
rect 115 1952 116 1956
rect 110 1951 116 1952
rect 1094 1956 1100 1957
rect 1094 1952 1095 1956
rect 1099 1952 1100 1956
rect 1134 1955 1135 1959
rect 1139 1955 1140 1959
rect 2118 1959 2124 1960
rect 1134 1954 1140 1955
rect 1302 1956 1308 1957
rect 1094 1951 1100 1952
rect 112 1931 114 1951
rect 190 1948 196 1949
rect 190 1944 191 1948
rect 195 1944 196 1948
rect 190 1943 196 1944
rect 246 1948 252 1949
rect 246 1944 247 1948
rect 251 1944 252 1948
rect 246 1943 252 1944
rect 310 1948 316 1949
rect 310 1944 311 1948
rect 315 1944 316 1948
rect 310 1943 316 1944
rect 374 1948 380 1949
rect 374 1944 375 1948
rect 379 1944 380 1948
rect 374 1943 380 1944
rect 446 1948 452 1949
rect 446 1944 447 1948
rect 451 1944 452 1948
rect 446 1943 452 1944
rect 518 1948 524 1949
rect 518 1944 519 1948
rect 523 1944 524 1948
rect 518 1943 524 1944
rect 590 1948 596 1949
rect 590 1944 591 1948
rect 595 1944 596 1948
rect 590 1943 596 1944
rect 654 1948 660 1949
rect 654 1944 655 1948
rect 659 1944 660 1948
rect 654 1943 660 1944
rect 718 1948 724 1949
rect 718 1944 719 1948
rect 723 1944 724 1948
rect 718 1943 724 1944
rect 774 1948 780 1949
rect 774 1944 775 1948
rect 779 1944 780 1948
rect 774 1943 780 1944
rect 822 1948 828 1949
rect 822 1944 823 1948
rect 827 1944 828 1948
rect 822 1943 828 1944
rect 870 1948 876 1949
rect 870 1944 871 1948
rect 875 1944 876 1948
rect 870 1943 876 1944
rect 918 1948 924 1949
rect 918 1944 919 1948
rect 923 1944 924 1948
rect 918 1943 924 1944
rect 966 1948 972 1949
rect 966 1944 967 1948
rect 971 1944 972 1948
rect 966 1943 972 1944
rect 1006 1948 1012 1949
rect 1006 1944 1007 1948
rect 1011 1944 1012 1948
rect 1006 1943 1012 1944
rect 1046 1948 1052 1949
rect 1046 1944 1047 1948
rect 1051 1944 1052 1948
rect 1046 1943 1052 1944
rect 192 1931 194 1943
rect 248 1931 250 1943
rect 312 1931 314 1943
rect 376 1931 378 1943
rect 448 1931 450 1943
rect 520 1931 522 1943
rect 592 1931 594 1943
rect 656 1931 658 1943
rect 720 1931 722 1943
rect 776 1931 778 1943
rect 824 1931 826 1943
rect 872 1931 874 1943
rect 920 1931 922 1943
rect 968 1931 970 1943
rect 1008 1931 1010 1943
rect 1048 1931 1050 1943
rect 1096 1931 1098 1951
rect 1136 1947 1138 1954
rect 1302 1952 1303 1956
rect 1307 1952 1308 1956
rect 1302 1951 1308 1952
rect 1382 1956 1388 1957
rect 1382 1952 1383 1956
rect 1387 1952 1388 1956
rect 1382 1951 1388 1952
rect 1462 1956 1468 1957
rect 1462 1952 1463 1956
rect 1467 1952 1468 1956
rect 1462 1951 1468 1952
rect 1542 1956 1548 1957
rect 1542 1952 1543 1956
rect 1547 1952 1548 1956
rect 1542 1951 1548 1952
rect 1614 1956 1620 1957
rect 1614 1952 1615 1956
rect 1619 1952 1620 1956
rect 1614 1951 1620 1952
rect 1686 1956 1692 1957
rect 1686 1952 1687 1956
rect 1691 1952 1692 1956
rect 1686 1951 1692 1952
rect 1750 1956 1756 1957
rect 1750 1952 1751 1956
rect 1755 1952 1756 1956
rect 1750 1951 1756 1952
rect 1814 1956 1820 1957
rect 1814 1952 1815 1956
rect 1819 1952 1820 1956
rect 1814 1951 1820 1952
rect 1878 1956 1884 1957
rect 1878 1952 1879 1956
rect 1883 1952 1884 1956
rect 1878 1951 1884 1952
rect 1950 1956 1956 1957
rect 1950 1952 1951 1956
rect 1955 1952 1956 1956
rect 1950 1951 1956 1952
rect 2022 1956 2028 1957
rect 2022 1952 2023 1956
rect 2027 1952 2028 1956
rect 2022 1951 2028 1952
rect 2070 1956 2076 1957
rect 2070 1952 2071 1956
rect 2075 1952 2076 1956
rect 2118 1955 2119 1959
rect 2123 1955 2124 1959
rect 2118 1954 2124 1955
rect 2070 1951 2076 1952
rect 1304 1947 1306 1951
rect 1384 1947 1386 1951
rect 1464 1947 1466 1951
rect 1544 1947 1546 1951
rect 1616 1947 1618 1951
rect 1688 1947 1690 1951
rect 1752 1947 1754 1951
rect 1816 1947 1818 1951
rect 1880 1947 1882 1951
rect 1952 1947 1954 1951
rect 2024 1947 2026 1951
rect 2072 1947 2074 1951
rect 2120 1947 2122 1954
rect 1135 1946 1139 1947
rect 1135 1941 1139 1942
rect 1159 1946 1163 1947
rect 1159 1941 1163 1942
rect 1223 1946 1227 1947
rect 1223 1941 1227 1942
rect 1303 1946 1307 1947
rect 1303 1941 1307 1942
rect 1383 1946 1387 1947
rect 1383 1941 1387 1942
rect 1463 1946 1467 1947
rect 1463 1941 1467 1942
rect 1535 1946 1539 1947
rect 1535 1941 1539 1942
rect 1543 1946 1547 1947
rect 1543 1941 1547 1942
rect 1615 1946 1619 1947
rect 1615 1941 1619 1942
rect 1687 1946 1691 1947
rect 1687 1941 1691 1942
rect 1695 1946 1699 1947
rect 1695 1941 1699 1942
rect 1751 1946 1755 1947
rect 1751 1941 1755 1942
rect 1783 1946 1787 1947
rect 1783 1941 1787 1942
rect 1815 1946 1819 1947
rect 1815 1941 1819 1942
rect 1879 1946 1883 1947
rect 1879 1941 1883 1942
rect 1951 1946 1955 1947
rect 1951 1941 1955 1942
rect 1983 1946 1987 1947
rect 1983 1941 1987 1942
rect 2023 1946 2027 1947
rect 2023 1941 2027 1942
rect 2071 1946 2075 1947
rect 2071 1941 2075 1942
rect 2119 1946 2123 1947
rect 2119 1941 2123 1942
rect 1136 1938 1138 1941
rect 1158 1940 1164 1941
rect 1134 1937 1140 1938
rect 1134 1933 1135 1937
rect 1139 1933 1140 1937
rect 1158 1936 1159 1940
rect 1163 1936 1164 1940
rect 1158 1935 1164 1936
rect 1222 1940 1228 1941
rect 1222 1936 1223 1940
rect 1227 1936 1228 1940
rect 1222 1935 1228 1936
rect 1302 1940 1308 1941
rect 1302 1936 1303 1940
rect 1307 1936 1308 1940
rect 1302 1935 1308 1936
rect 1382 1940 1388 1941
rect 1382 1936 1383 1940
rect 1387 1936 1388 1940
rect 1382 1935 1388 1936
rect 1462 1940 1468 1941
rect 1462 1936 1463 1940
rect 1467 1936 1468 1940
rect 1462 1935 1468 1936
rect 1534 1940 1540 1941
rect 1534 1936 1535 1940
rect 1539 1936 1540 1940
rect 1534 1935 1540 1936
rect 1614 1940 1620 1941
rect 1614 1936 1615 1940
rect 1619 1936 1620 1940
rect 1614 1935 1620 1936
rect 1694 1940 1700 1941
rect 1694 1936 1695 1940
rect 1699 1936 1700 1940
rect 1694 1935 1700 1936
rect 1782 1940 1788 1941
rect 1782 1936 1783 1940
rect 1787 1936 1788 1940
rect 1782 1935 1788 1936
rect 1878 1940 1884 1941
rect 1878 1936 1879 1940
rect 1883 1936 1884 1940
rect 1878 1935 1884 1936
rect 1982 1940 1988 1941
rect 1982 1936 1983 1940
rect 1987 1936 1988 1940
rect 1982 1935 1988 1936
rect 2070 1940 2076 1941
rect 2070 1936 2071 1940
rect 2075 1936 2076 1940
rect 2120 1938 2122 1941
rect 2070 1935 2076 1936
rect 2118 1937 2124 1938
rect 1134 1932 1140 1933
rect 2118 1933 2119 1937
rect 2123 1933 2124 1937
rect 2118 1932 2124 1933
rect 111 1930 115 1931
rect 111 1925 115 1926
rect 135 1930 139 1931
rect 135 1925 139 1926
rect 175 1930 179 1931
rect 175 1925 179 1926
rect 191 1930 195 1931
rect 191 1925 195 1926
rect 231 1930 235 1931
rect 231 1925 235 1926
rect 247 1930 251 1931
rect 247 1925 251 1926
rect 295 1930 299 1931
rect 295 1925 299 1926
rect 311 1930 315 1931
rect 311 1925 315 1926
rect 367 1930 371 1931
rect 367 1925 371 1926
rect 375 1930 379 1931
rect 375 1925 379 1926
rect 431 1930 435 1931
rect 431 1925 435 1926
rect 447 1930 451 1931
rect 447 1925 451 1926
rect 495 1930 499 1931
rect 495 1925 499 1926
rect 519 1930 523 1931
rect 519 1925 523 1926
rect 559 1930 563 1931
rect 559 1925 563 1926
rect 591 1930 595 1931
rect 591 1925 595 1926
rect 615 1930 619 1931
rect 615 1925 619 1926
rect 655 1930 659 1931
rect 655 1925 659 1926
rect 671 1930 675 1931
rect 671 1925 675 1926
rect 719 1930 723 1931
rect 719 1925 723 1926
rect 727 1930 731 1931
rect 727 1925 731 1926
rect 775 1930 779 1931
rect 775 1925 779 1926
rect 783 1930 787 1931
rect 783 1925 787 1926
rect 823 1930 827 1931
rect 823 1925 827 1926
rect 847 1930 851 1931
rect 847 1925 851 1926
rect 871 1930 875 1931
rect 871 1925 875 1926
rect 919 1930 923 1931
rect 919 1925 923 1926
rect 967 1930 971 1931
rect 967 1925 971 1926
rect 1007 1930 1011 1931
rect 1007 1925 1011 1926
rect 1047 1930 1051 1931
rect 1047 1925 1051 1926
rect 1095 1930 1099 1931
rect 1095 1925 1099 1926
rect 112 1905 114 1925
rect 136 1913 138 1925
rect 176 1913 178 1925
rect 232 1913 234 1925
rect 296 1913 298 1925
rect 368 1913 370 1925
rect 432 1913 434 1925
rect 496 1913 498 1925
rect 560 1913 562 1925
rect 616 1913 618 1925
rect 672 1913 674 1925
rect 728 1913 730 1925
rect 784 1913 786 1925
rect 848 1913 850 1925
rect 134 1912 140 1913
rect 134 1908 135 1912
rect 139 1908 140 1912
rect 134 1907 140 1908
rect 174 1912 180 1913
rect 174 1908 175 1912
rect 179 1908 180 1912
rect 174 1907 180 1908
rect 230 1912 236 1913
rect 230 1908 231 1912
rect 235 1908 236 1912
rect 230 1907 236 1908
rect 294 1912 300 1913
rect 294 1908 295 1912
rect 299 1908 300 1912
rect 294 1907 300 1908
rect 366 1912 372 1913
rect 366 1908 367 1912
rect 371 1908 372 1912
rect 366 1907 372 1908
rect 430 1912 436 1913
rect 430 1908 431 1912
rect 435 1908 436 1912
rect 430 1907 436 1908
rect 494 1912 500 1913
rect 494 1908 495 1912
rect 499 1908 500 1912
rect 494 1907 500 1908
rect 558 1912 564 1913
rect 558 1908 559 1912
rect 563 1908 564 1912
rect 558 1907 564 1908
rect 614 1912 620 1913
rect 614 1908 615 1912
rect 619 1908 620 1912
rect 614 1907 620 1908
rect 670 1912 676 1913
rect 670 1908 671 1912
rect 675 1908 676 1912
rect 670 1907 676 1908
rect 726 1912 732 1913
rect 726 1908 727 1912
rect 731 1908 732 1912
rect 726 1907 732 1908
rect 782 1912 788 1913
rect 782 1908 783 1912
rect 787 1908 788 1912
rect 782 1907 788 1908
rect 846 1912 852 1913
rect 846 1908 847 1912
rect 851 1908 852 1912
rect 846 1907 852 1908
rect 1096 1905 1098 1925
rect 1134 1920 1140 1921
rect 1134 1916 1135 1920
rect 1139 1916 1140 1920
rect 1134 1915 1140 1916
rect 2118 1920 2124 1921
rect 2118 1916 2119 1920
rect 2123 1916 2124 1920
rect 2118 1915 2124 1916
rect 110 1904 116 1905
rect 110 1900 111 1904
rect 115 1900 116 1904
rect 110 1899 116 1900
rect 1094 1904 1100 1905
rect 1094 1900 1095 1904
rect 1099 1900 1100 1904
rect 1094 1899 1100 1900
rect 1136 1891 1138 1915
rect 1158 1912 1164 1913
rect 1158 1908 1159 1912
rect 1163 1908 1164 1912
rect 1158 1907 1164 1908
rect 1222 1912 1228 1913
rect 1222 1908 1223 1912
rect 1227 1908 1228 1912
rect 1222 1907 1228 1908
rect 1302 1912 1308 1913
rect 1302 1908 1303 1912
rect 1307 1908 1308 1912
rect 1302 1907 1308 1908
rect 1382 1912 1388 1913
rect 1382 1908 1383 1912
rect 1387 1908 1388 1912
rect 1382 1907 1388 1908
rect 1462 1912 1468 1913
rect 1462 1908 1463 1912
rect 1467 1908 1468 1912
rect 1462 1907 1468 1908
rect 1534 1912 1540 1913
rect 1534 1908 1535 1912
rect 1539 1908 1540 1912
rect 1534 1907 1540 1908
rect 1614 1912 1620 1913
rect 1614 1908 1615 1912
rect 1619 1908 1620 1912
rect 1614 1907 1620 1908
rect 1694 1912 1700 1913
rect 1694 1908 1695 1912
rect 1699 1908 1700 1912
rect 1694 1907 1700 1908
rect 1782 1912 1788 1913
rect 1782 1908 1783 1912
rect 1787 1908 1788 1912
rect 1782 1907 1788 1908
rect 1878 1912 1884 1913
rect 1878 1908 1879 1912
rect 1883 1908 1884 1912
rect 1878 1907 1884 1908
rect 1982 1912 1988 1913
rect 1982 1908 1983 1912
rect 1987 1908 1988 1912
rect 1982 1907 1988 1908
rect 2070 1912 2076 1913
rect 2070 1908 2071 1912
rect 2075 1908 2076 1912
rect 2070 1907 2076 1908
rect 1160 1891 1162 1907
rect 1224 1891 1226 1907
rect 1304 1891 1306 1907
rect 1384 1891 1386 1907
rect 1464 1891 1466 1907
rect 1536 1891 1538 1907
rect 1616 1891 1618 1907
rect 1696 1891 1698 1907
rect 1784 1891 1786 1907
rect 1880 1891 1882 1907
rect 1984 1891 1986 1907
rect 2072 1891 2074 1907
rect 2120 1891 2122 1915
rect 1135 1890 1139 1891
rect 110 1887 116 1888
rect 110 1883 111 1887
rect 115 1883 116 1887
rect 1094 1887 1100 1888
rect 110 1882 116 1883
rect 134 1884 140 1885
rect 112 1875 114 1882
rect 134 1880 135 1884
rect 139 1880 140 1884
rect 134 1879 140 1880
rect 174 1884 180 1885
rect 174 1880 175 1884
rect 179 1880 180 1884
rect 174 1879 180 1880
rect 230 1884 236 1885
rect 230 1880 231 1884
rect 235 1880 236 1884
rect 230 1879 236 1880
rect 294 1884 300 1885
rect 294 1880 295 1884
rect 299 1880 300 1884
rect 294 1879 300 1880
rect 366 1884 372 1885
rect 366 1880 367 1884
rect 371 1880 372 1884
rect 366 1879 372 1880
rect 430 1884 436 1885
rect 430 1880 431 1884
rect 435 1880 436 1884
rect 430 1879 436 1880
rect 494 1884 500 1885
rect 494 1880 495 1884
rect 499 1880 500 1884
rect 494 1879 500 1880
rect 558 1884 564 1885
rect 558 1880 559 1884
rect 563 1880 564 1884
rect 558 1879 564 1880
rect 614 1884 620 1885
rect 614 1880 615 1884
rect 619 1880 620 1884
rect 614 1879 620 1880
rect 670 1884 676 1885
rect 670 1880 671 1884
rect 675 1880 676 1884
rect 670 1879 676 1880
rect 726 1884 732 1885
rect 726 1880 727 1884
rect 731 1880 732 1884
rect 726 1879 732 1880
rect 782 1884 788 1885
rect 782 1880 783 1884
rect 787 1880 788 1884
rect 782 1879 788 1880
rect 846 1884 852 1885
rect 846 1880 847 1884
rect 851 1880 852 1884
rect 1094 1883 1095 1887
rect 1099 1883 1100 1887
rect 1135 1885 1139 1886
rect 1159 1890 1163 1891
rect 1159 1885 1163 1886
rect 1199 1890 1203 1891
rect 1199 1885 1203 1886
rect 1223 1890 1227 1891
rect 1223 1885 1227 1886
rect 1263 1890 1267 1891
rect 1263 1885 1267 1886
rect 1303 1890 1307 1891
rect 1303 1885 1307 1886
rect 1327 1890 1331 1891
rect 1327 1885 1331 1886
rect 1383 1890 1387 1891
rect 1383 1885 1387 1886
rect 1391 1890 1395 1891
rect 1391 1885 1395 1886
rect 1447 1890 1451 1891
rect 1447 1885 1451 1886
rect 1463 1890 1467 1891
rect 1463 1885 1467 1886
rect 1503 1890 1507 1891
rect 1503 1885 1507 1886
rect 1535 1890 1539 1891
rect 1535 1885 1539 1886
rect 1559 1890 1563 1891
rect 1559 1885 1563 1886
rect 1615 1890 1619 1891
rect 1615 1885 1619 1886
rect 1631 1890 1635 1891
rect 1631 1885 1635 1886
rect 1695 1890 1699 1891
rect 1695 1885 1699 1886
rect 1711 1890 1715 1891
rect 1711 1885 1715 1886
rect 1783 1890 1787 1891
rect 1783 1885 1787 1886
rect 1799 1890 1803 1891
rect 1799 1885 1803 1886
rect 1879 1890 1883 1891
rect 1879 1885 1883 1886
rect 1895 1890 1899 1891
rect 1895 1885 1899 1886
rect 1983 1890 1987 1891
rect 1983 1885 1987 1886
rect 1991 1890 1995 1891
rect 1991 1885 1995 1886
rect 2071 1890 2075 1891
rect 2071 1885 2075 1886
rect 2119 1890 2123 1891
rect 2119 1885 2123 1886
rect 1094 1882 1100 1883
rect 846 1879 852 1880
rect 136 1875 138 1879
rect 176 1875 178 1879
rect 232 1875 234 1879
rect 296 1875 298 1879
rect 368 1875 370 1879
rect 432 1875 434 1879
rect 496 1875 498 1879
rect 560 1875 562 1879
rect 616 1875 618 1879
rect 672 1875 674 1879
rect 728 1875 730 1879
rect 784 1875 786 1879
rect 848 1875 850 1879
rect 1096 1875 1098 1882
rect 111 1874 115 1875
rect 111 1869 115 1870
rect 135 1874 139 1875
rect 135 1869 139 1870
rect 175 1874 179 1875
rect 175 1869 179 1870
rect 199 1874 203 1875
rect 199 1869 203 1870
rect 231 1874 235 1875
rect 231 1869 235 1870
rect 271 1874 275 1875
rect 271 1869 275 1870
rect 295 1874 299 1875
rect 295 1869 299 1870
rect 335 1874 339 1875
rect 335 1869 339 1870
rect 367 1874 371 1875
rect 367 1869 371 1870
rect 399 1874 403 1875
rect 399 1869 403 1870
rect 431 1874 435 1875
rect 431 1869 435 1870
rect 455 1874 459 1875
rect 455 1869 459 1870
rect 495 1874 499 1875
rect 495 1869 499 1870
rect 503 1874 507 1875
rect 503 1869 507 1870
rect 551 1874 555 1875
rect 551 1869 555 1870
rect 559 1874 563 1875
rect 559 1869 563 1870
rect 599 1874 603 1875
rect 599 1869 603 1870
rect 615 1874 619 1875
rect 615 1869 619 1870
rect 647 1874 651 1875
rect 647 1869 651 1870
rect 671 1874 675 1875
rect 671 1869 675 1870
rect 695 1874 699 1875
rect 695 1869 699 1870
rect 727 1874 731 1875
rect 727 1869 731 1870
rect 751 1874 755 1875
rect 751 1869 755 1870
rect 783 1874 787 1875
rect 783 1869 787 1870
rect 847 1874 851 1875
rect 847 1869 851 1870
rect 1095 1874 1099 1875
rect 1095 1869 1099 1870
rect 112 1866 114 1869
rect 134 1868 140 1869
rect 110 1865 116 1866
rect 110 1861 111 1865
rect 115 1861 116 1865
rect 134 1864 135 1868
rect 139 1864 140 1868
rect 134 1863 140 1864
rect 198 1868 204 1869
rect 198 1864 199 1868
rect 203 1864 204 1868
rect 198 1863 204 1864
rect 270 1868 276 1869
rect 270 1864 271 1868
rect 275 1864 276 1868
rect 270 1863 276 1864
rect 334 1868 340 1869
rect 334 1864 335 1868
rect 339 1864 340 1868
rect 334 1863 340 1864
rect 398 1868 404 1869
rect 398 1864 399 1868
rect 403 1864 404 1868
rect 398 1863 404 1864
rect 454 1868 460 1869
rect 454 1864 455 1868
rect 459 1864 460 1868
rect 454 1863 460 1864
rect 502 1868 508 1869
rect 502 1864 503 1868
rect 507 1864 508 1868
rect 502 1863 508 1864
rect 550 1868 556 1869
rect 550 1864 551 1868
rect 555 1864 556 1868
rect 550 1863 556 1864
rect 598 1868 604 1869
rect 598 1864 599 1868
rect 603 1864 604 1868
rect 598 1863 604 1864
rect 646 1868 652 1869
rect 646 1864 647 1868
rect 651 1864 652 1868
rect 646 1863 652 1864
rect 694 1868 700 1869
rect 694 1864 695 1868
rect 699 1864 700 1868
rect 694 1863 700 1864
rect 750 1868 756 1869
rect 750 1864 751 1868
rect 755 1864 756 1868
rect 1096 1866 1098 1869
rect 750 1863 756 1864
rect 1094 1865 1100 1866
rect 1136 1865 1138 1885
rect 1160 1873 1162 1885
rect 1200 1873 1202 1885
rect 1264 1873 1266 1885
rect 1328 1873 1330 1885
rect 1392 1873 1394 1885
rect 1448 1873 1450 1885
rect 1504 1873 1506 1885
rect 1560 1873 1562 1885
rect 1632 1873 1634 1885
rect 1712 1873 1714 1885
rect 1800 1873 1802 1885
rect 1896 1873 1898 1885
rect 1992 1873 1994 1885
rect 2072 1873 2074 1885
rect 1158 1872 1164 1873
rect 1158 1868 1159 1872
rect 1163 1868 1164 1872
rect 1158 1867 1164 1868
rect 1198 1872 1204 1873
rect 1198 1868 1199 1872
rect 1203 1868 1204 1872
rect 1198 1867 1204 1868
rect 1262 1872 1268 1873
rect 1262 1868 1263 1872
rect 1267 1868 1268 1872
rect 1262 1867 1268 1868
rect 1326 1872 1332 1873
rect 1326 1868 1327 1872
rect 1331 1868 1332 1872
rect 1326 1867 1332 1868
rect 1390 1872 1396 1873
rect 1390 1868 1391 1872
rect 1395 1868 1396 1872
rect 1390 1867 1396 1868
rect 1446 1872 1452 1873
rect 1446 1868 1447 1872
rect 1451 1868 1452 1872
rect 1446 1867 1452 1868
rect 1502 1872 1508 1873
rect 1502 1868 1503 1872
rect 1507 1868 1508 1872
rect 1502 1867 1508 1868
rect 1558 1872 1564 1873
rect 1558 1868 1559 1872
rect 1563 1868 1564 1872
rect 1558 1867 1564 1868
rect 1630 1872 1636 1873
rect 1630 1868 1631 1872
rect 1635 1868 1636 1872
rect 1630 1867 1636 1868
rect 1710 1872 1716 1873
rect 1710 1868 1711 1872
rect 1715 1868 1716 1872
rect 1710 1867 1716 1868
rect 1798 1872 1804 1873
rect 1798 1868 1799 1872
rect 1803 1868 1804 1872
rect 1798 1867 1804 1868
rect 1894 1872 1900 1873
rect 1894 1868 1895 1872
rect 1899 1868 1900 1872
rect 1894 1867 1900 1868
rect 1990 1872 1996 1873
rect 1990 1868 1991 1872
rect 1995 1868 1996 1872
rect 1990 1867 1996 1868
rect 2070 1872 2076 1873
rect 2070 1868 2071 1872
rect 2075 1868 2076 1872
rect 2070 1867 2076 1868
rect 2120 1865 2122 1885
rect 110 1860 116 1861
rect 1094 1861 1095 1865
rect 1099 1861 1100 1865
rect 1094 1860 1100 1861
rect 1134 1864 1140 1865
rect 1134 1860 1135 1864
rect 1139 1860 1140 1864
rect 1134 1859 1140 1860
rect 2118 1864 2124 1865
rect 2118 1860 2119 1864
rect 2123 1860 2124 1864
rect 2118 1859 2124 1860
rect 110 1848 116 1849
rect 110 1844 111 1848
rect 115 1844 116 1848
rect 110 1843 116 1844
rect 1094 1848 1100 1849
rect 1094 1844 1095 1848
rect 1099 1844 1100 1848
rect 1094 1843 1100 1844
rect 1134 1847 1140 1848
rect 1134 1843 1135 1847
rect 1139 1843 1140 1847
rect 2118 1847 2124 1848
rect 112 1815 114 1843
rect 134 1840 140 1841
rect 134 1836 135 1840
rect 139 1836 140 1840
rect 134 1835 140 1836
rect 198 1840 204 1841
rect 198 1836 199 1840
rect 203 1836 204 1840
rect 198 1835 204 1836
rect 270 1840 276 1841
rect 270 1836 271 1840
rect 275 1836 276 1840
rect 270 1835 276 1836
rect 334 1840 340 1841
rect 334 1836 335 1840
rect 339 1836 340 1840
rect 334 1835 340 1836
rect 398 1840 404 1841
rect 398 1836 399 1840
rect 403 1836 404 1840
rect 398 1835 404 1836
rect 454 1840 460 1841
rect 454 1836 455 1840
rect 459 1836 460 1840
rect 454 1835 460 1836
rect 502 1840 508 1841
rect 502 1836 503 1840
rect 507 1836 508 1840
rect 502 1835 508 1836
rect 550 1840 556 1841
rect 550 1836 551 1840
rect 555 1836 556 1840
rect 550 1835 556 1836
rect 598 1840 604 1841
rect 598 1836 599 1840
rect 603 1836 604 1840
rect 598 1835 604 1836
rect 646 1840 652 1841
rect 646 1836 647 1840
rect 651 1836 652 1840
rect 646 1835 652 1836
rect 694 1840 700 1841
rect 694 1836 695 1840
rect 699 1836 700 1840
rect 694 1835 700 1836
rect 750 1840 756 1841
rect 750 1836 751 1840
rect 755 1836 756 1840
rect 750 1835 756 1836
rect 136 1815 138 1835
rect 200 1815 202 1835
rect 272 1815 274 1835
rect 336 1815 338 1835
rect 400 1815 402 1835
rect 456 1815 458 1835
rect 504 1815 506 1835
rect 552 1815 554 1835
rect 600 1815 602 1835
rect 648 1815 650 1835
rect 696 1815 698 1835
rect 752 1815 754 1835
rect 1096 1815 1098 1843
rect 1134 1842 1140 1843
rect 1158 1844 1164 1845
rect 1136 1839 1138 1842
rect 1158 1840 1159 1844
rect 1163 1840 1164 1844
rect 1158 1839 1164 1840
rect 1198 1844 1204 1845
rect 1198 1840 1199 1844
rect 1203 1840 1204 1844
rect 1198 1839 1204 1840
rect 1262 1844 1268 1845
rect 1262 1840 1263 1844
rect 1267 1840 1268 1844
rect 1262 1839 1268 1840
rect 1326 1844 1332 1845
rect 1326 1840 1327 1844
rect 1331 1840 1332 1844
rect 1326 1839 1332 1840
rect 1390 1844 1396 1845
rect 1390 1840 1391 1844
rect 1395 1840 1396 1844
rect 1390 1839 1396 1840
rect 1446 1844 1452 1845
rect 1446 1840 1447 1844
rect 1451 1840 1452 1844
rect 1446 1839 1452 1840
rect 1502 1844 1508 1845
rect 1502 1840 1503 1844
rect 1507 1840 1508 1844
rect 1502 1839 1508 1840
rect 1558 1844 1564 1845
rect 1558 1840 1559 1844
rect 1563 1840 1564 1844
rect 1558 1839 1564 1840
rect 1630 1844 1636 1845
rect 1630 1840 1631 1844
rect 1635 1840 1636 1844
rect 1630 1839 1636 1840
rect 1710 1844 1716 1845
rect 1710 1840 1711 1844
rect 1715 1840 1716 1844
rect 1710 1839 1716 1840
rect 1798 1844 1804 1845
rect 1798 1840 1799 1844
rect 1803 1840 1804 1844
rect 1798 1839 1804 1840
rect 1894 1844 1900 1845
rect 1894 1840 1895 1844
rect 1899 1840 1900 1844
rect 1894 1839 1900 1840
rect 1990 1844 1996 1845
rect 1990 1840 1991 1844
rect 1995 1840 1996 1844
rect 1990 1839 1996 1840
rect 2070 1844 2076 1845
rect 2070 1840 2071 1844
rect 2075 1840 2076 1844
rect 2118 1843 2119 1847
rect 2123 1843 2124 1847
rect 2118 1842 2124 1843
rect 2070 1839 2076 1840
rect 2120 1839 2122 1842
rect 1135 1838 1139 1839
rect 1135 1833 1139 1834
rect 1159 1838 1163 1839
rect 1159 1833 1163 1834
rect 1199 1838 1203 1839
rect 1199 1833 1203 1834
rect 1231 1838 1235 1839
rect 1231 1833 1235 1834
rect 1263 1838 1267 1839
rect 1263 1833 1267 1834
rect 1303 1838 1307 1839
rect 1303 1833 1307 1834
rect 1327 1838 1331 1839
rect 1327 1833 1331 1834
rect 1383 1838 1387 1839
rect 1383 1833 1387 1834
rect 1391 1838 1395 1839
rect 1391 1833 1395 1834
rect 1447 1838 1451 1839
rect 1447 1833 1451 1834
rect 1463 1838 1467 1839
rect 1463 1833 1467 1834
rect 1503 1838 1507 1839
rect 1503 1833 1507 1834
rect 1551 1838 1555 1839
rect 1551 1833 1555 1834
rect 1559 1838 1563 1839
rect 1559 1833 1563 1834
rect 1631 1838 1635 1839
rect 1631 1833 1635 1834
rect 1647 1838 1651 1839
rect 1647 1833 1651 1834
rect 1711 1838 1715 1839
rect 1711 1833 1715 1834
rect 1751 1838 1755 1839
rect 1751 1833 1755 1834
rect 1799 1838 1803 1839
rect 1799 1833 1803 1834
rect 1855 1838 1859 1839
rect 1855 1833 1859 1834
rect 1895 1838 1899 1839
rect 1895 1833 1899 1834
rect 1967 1838 1971 1839
rect 1967 1833 1971 1834
rect 1991 1838 1995 1839
rect 1991 1833 1995 1834
rect 2071 1838 2075 1839
rect 2071 1833 2075 1834
rect 2119 1838 2123 1839
rect 2119 1833 2123 1834
rect 1136 1830 1138 1833
rect 1158 1832 1164 1833
rect 1134 1829 1140 1830
rect 1134 1825 1135 1829
rect 1139 1825 1140 1829
rect 1158 1828 1159 1832
rect 1163 1828 1164 1832
rect 1158 1827 1164 1828
rect 1230 1832 1236 1833
rect 1230 1828 1231 1832
rect 1235 1828 1236 1832
rect 1230 1827 1236 1828
rect 1302 1832 1308 1833
rect 1302 1828 1303 1832
rect 1307 1828 1308 1832
rect 1302 1827 1308 1828
rect 1382 1832 1388 1833
rect 1382 1828 1383 1832
rect 1387 1828 1388 1832
rect 1382 1827 1388 1828
rect 1462 1832 1468 1833
rect 1462 1828 1463 1832
rect 1467 1828 1468 1832
rect 1462 1827 1468 1828
rect 1550 1832 1556 1833
rect 1550 1828 1551 1832
rect 1555 1828 1556 1832
rect 1550 1827 1556 1828
rect 1646 1832 1652 1833
rect 1646 1828 1647 1832
rect 1651 1828 1652 1832
rect 1646 1827 1652 1828
rect 1750 1832 1756 1833
rect 1750 1828 1751 1832
rect 1755 1828 1756 1832
rect 1750 1827 1756 1828
rect 1854 1832 1860 1833
rect 1854 1828 1855 1832
rect 1859 1828 1860 1832
rect 1854 1827 1860 1828
rect 1966 1832 1972 1833
rect 1966 1828 1967 1832
rect 1971 1828 1972 1832
rect 1966 1827 1972 1828
rect 2070 1832 2076 1833
rect 2070 1828 2071 1832
rect 2075 1828 2076 1832
rect 2120 1830 2122 1833
rect 2070 1827 2076 1828
rect 2118 1829 2124 1830
rect 1134 1824 1140 1825
rect 2118 1825 2119 1829
rect 2123 1825 2124 1829
rect 2118 1824 2124 1825
rect 111 1814 115 1815
rect 111 1809 115 1810
rect 135 1814 139 1815
rect 135 1809 139 1810
rect 151 1814 155 1815
rect 151 1809 155 1810
rect 199 1814 203 1815
rect 199 1809 203 1810
rect 215 1814 219 1815
rect 215 1809 219 1810
rect 271 1814 275 1815
rect 271 1809 275 1810
rect 327 1814 331 1815
rect 327 1809 331 1810
rect 335 1814 339 1815
rect 335 1809 339 1810
rect 383 1814 387 1815
rect 383 1809 387 1810
rect 399 1814 403 1815
rect 399 1809 403 1810
rect 431 1814 435 1815
rect 431 1809 435 1810
rect 455 1814 459 1815
rect 455 1809 459 1810
rect 479 1814 483 1815
rect 479 1809 483 1810
rect 503 1814 507 1815
rect 503 1809 507 1810
rect 527 1814 531 1815
rect 527 1809 531 1810
rect 551 1814 555 1815
rect 551 1809 555 1810
rect 575 1814 579 1815
rect 575 1809 579 1810
rect 599 1814 603 1815
rect 599 1809 603 1810
rect 623 1814 627 1815
rect 623 1809 627 1810
rect 647 1814 651 1815
rect 647 1809 651 1810
rect 671 1814 675 1815
rect 671 1809 675 1810
rect 695 1814 699 1815
rect 695 1809 699 1810
rect 727 1814 731 1815
rect 727 1809 731 1810
rect 751 1814 755 1815
rect 751 1809 755 1810
rect 1095 1814 1099 1815
rect 1095 1809 1099 1810
rect 1134 1812 1140 1813
rect 112 1789 114 1809
rect 152 1797 154 1809
rect 216 1797 218 1809
rect 272 1797 274 1809
rect 328 1797 330 1809
rect 384 1797 386 1809
rect 432 1797 434 1809
rect 480 1797 482 1809
rect 528 1797 530 1809
rect 576 1797 578 1809
rect 624 1797 626 1809
rect 672 1797 674 1809
rect 728 1797 730 1809
rect 150 1796 156 1797
rect 150 1792 151 1796
rect 155 1792 156 1796
rect 150 1791 156 1792
rect 214 1796 220 1797
rect 214 1792 215 1796
rect 219 1792 220 1796
rect 214 1791 220 1792
rect 270 1796 276 1797
rect 270 1792 271 1796
rect 275 1792 276 1796
rect 270 1791 276 1792
rect 326 1796 332 1797
rect 326 1792 327 1796
rect 331 1792 332 1796
rect 326 1791 332 1792
rect 382 1796 388 1797
rect 382 1792 383 1796
rect 387 1792 388 1796
rect 382 1791 388 1792
rect 430 1796 436 1797
rect 430 1792 431 1796
rect 435 1792 436 1796
rect 430 1791 436 1792
rect 478 1796 484 1797
rect 478 1792 479 1796
rect 483 1792 484 1796
rect 478 1791 484 1792
rect 526 1796 532 1797
rect 526 1792 527 1796
rect 531 1792 532 1796
rect 526 1791 532 1792
rect 574 1796 580 1797
rect 574 1792 575 1796
rect 579 1792 580 1796
rect 574 1791 580 1792
rect 622 1796 628 1797
rect 622 1792 623 1796
rect 627 1792 628 1796
rect 622 1791 628 1792
rect 670 1796 676 1797
rect 670 1792 671 1796
rect 675 1792 676 1796
rect 670 1791 676 1792
rect 726 1796 732 1797
rect 726 1792 727 1796
rect 731 1792 732 1796
rect 726 1791 732 1792
rect 1096 1789 1098 1809
rect 1134 1808 1135 1812
rect 1139 1808 1140 1812
rect 1134 1807 1140 1808
rect 2118 1812 2124 1813
rect 2118 1808 2119 1812
rect 2123 1808 2124 1812
rect 2118 1807 2124 1808
rect 110 1788 116 1789
rect 110 1784 111 1788
rect 115 1784 116 1788
rect 110 1783 116 1784
rect 1094 1788 1100 1789
rect 1094 1784 1095 1788
rect 1099 1784 1100 1788
rect 1136 1787 1138 1807
rect 1158 1804 1164 1805
rect 1158 1800 1159 1804
rect 1163 1800 1164 1804
rect 1158 1799 1164 1800
rect 1230 1804 1236 1805
rect 1230 1800 1231 1804
rect 1235 1800 1236 1804
rect 1230 1799 1236 1800
rect 1302 1804 1308 1805
rect 1302 1800 1303 1804
rect 1307 1800 1308 1804
rect 1302 1799 1308 1800
rect 1382 1804 1388 1805
rect 1382 1800 1383 1804
rect 1387 1800 1388 1804
rect 1382 1799 1388 1800
rect 1462 1804 1468 1805
rect 1462 1800 1463 1804
rect 1467 1800 1468 1804
rect 1462 1799 1468 1800
rect 1550 1804 1556 1805
rect 1550 1800 1551 1804
rect 1555 1800 1556 1804
rect 1550 1799 1556 1800
rect 1646 1804 1652 1805
rect 1646 1800 1647 1804
rect 1651 1800 1652 1804
rect 1646 1799 1652 1800
rect 1750 1804 1756 1805
rect 1750 1800 1751 1804
rect 1755 1800 1756 1804
rect 1750 1799 1756 1800
rect 1854 1804 1860 1805
rect 1854 1800 1855 1804
rect 1859 1800 1860 1804
rect 1854 1799 1860 1800
rect 1966 1804 1972 1805
rect 1966 1800 1967 1804
rect 1971 1800 1972 1804
rect 1966 1799 1972 1800
rect 2070 1804 2076 1805
rect 2070 1800 2071 1804
rect 2075 1800 2076 1804
rect 2070 1799 2076 1800
rect 1160 1787 1162 1799
rect 1232 1787 1234 1799
rect 1304 1787 1306 1799
rect 1384 1787 1386 1799
rect 1464 1787 1466 1799
rect 1552 1787 1554 1799
rect 1648 1787 1650 1799
rect 1752 1787 1754 1799
rect 1856 1787 1858 1799
rect 1968 1787 1970 1799
rect 2072 1787 2074 1799
rect 2120 1787 2122 1807
rect 1094 1783 1100 1784
rect 1135 1786 1139 1787
rect 1135 1781 1139 1782
rect 1159 1786 1163 1787
rect 1159 1781 1163 1782
rect 1191 1786 1195 1787
rect 1191 1781 1195 1782
rect 1231 1786 1235 1787
rect 1231 1781 1235 1782
rect 1255 1786 1259 1787
rect 1255 1781 1259 1782
rect 1303 1786 1307 1787
rect 1303 1781 1307 1782
rect 1319 1786 1323 1787
rect 1319 1781 1323 1782
rect 1383 1786 1387 1787
rect 1383 1781 1387 1782
rect 1455 1786 1459 1787
rect 1455 1781 1459 1782
rect 1463 1786 1467 1787
rect 1463 1781 1467 1782
rect 1527 1786 1531 1787
rect 1527 1781 1531 1782
rect 1551 1786 1555 1787
rect 1551 1781 1555 1782
rect 1607 1786 1611 1787
rect 1607 1781 1611 1782
rect 1647 1786 1651 1787
rect 1647 1781 1651 1782
rect 1687 1786 1691 1787
rect 1687 1781 1691 1782
rect 1751 1786 1755 1787
rect 1751 1781 1755 1782
rect 1767 1786 1771 1787
rect 1767 1781 1771 1782
rect 1847 1786 1851 1787
rect 1847 1781 1851 1782
rect 1855 1786 1859 1787
rect 1855 1781 1859 1782
rect 1927 1786 1931 1787
rect 1927 1781 1931 1782
rect 1967 1786 1971 1787
rect 1967 1781 1971 1782
rect 2007 1786 2011 1787
rect 2007 1781 2011 1782
rect 2071 1786 2075 1787
rect 2071 1781 2075 1782
rect 2119 1786 2123 1787
rect 2119 1781 2123 1782
rect 110 1771 116 1772
rect 110 1767 111 1771
rect 115 1767 116 1771
rect 1094 1771 1100 1772
rect 110 1766 116 1767
rect 150 1768 156 1769
rect 112 1763 114 1766
rect 150 1764 151 1768
rect 155 1764 156 1768
rect 150 1763 156 1764
rect 214 1768 220 1769
rect 214 1764 215 1768
rect 219 1764 220 1768
rect 214 1763 220 1764
rect 270 1768 276 1769
rect 270 1764 271 1768
rect 275 1764 276 1768
rect 270 1763 276 1764
rect 326 1768 332 1769
rect 326 1764 327 1768
rect 331 1764 332 1768
rect 326 1763 332 1764
rect 382 1768 388 1769
rect 382 1764 383 1768
rect 387 1764 388 1768
rect 382 1763 388 1764
rect 430 1768 436 1769
rect 430 1764 431 1768
rect 435 1764 436 1768
rect 430 1763 436 1764
rect 478 1768 484 1769
rect 478 1764 479 1768
rect 483 1764 484 1768
rect 478 1763 484 1764
rect 526 1768 532 1769
rect 526 1764 527 1768
rect 531 1764 532 1768
rect 526 1763 532 1764
rect 574 1768 580 1769
rect 574 1764 575 1768
rect 579 1764 580 1768
rect 574 1763 580 1764
rect 622 1768 628 1769
rect 622 1764 623 1768
rect 627 1764 628 1768
rect 622 1763 628 1764
rect 670 1768 676 1769
rect 670 1764 671 1768
rect 675 1764 676 1768
rect 670 1763 676 1764
rect 726 1768 732 1769
rect 726 1764 727 1768
rect 731 1764 732 1768
rect 1094 1767 1095 1771
rect 1099 1767 1100 1771
rect 1094 1766 1100 1767
rect 726 1763 732 1764
rect 1096 1763 1098 1766
rect 111 1762 115 1763
rect 111 1757 115 1758
rect 151 1762 155 1763
rect 151 1757 155 1758
rect 215 1762 219 1763
rect 215 1757 219 1758
rect 231 1762 235 1763
rect 231 1757 235 1758
rect 271 1762 275 1763
rect 271 1757 275 1758
rect 295 1762 299 1763
rect 295 1757 299 1758
rect 327 1762 331 1763
rect 327 1757 331 1758
rect 351 1762 355 1763
rect 351 1757 355 1758
rect 383 1762 387 1763
rect 383 1757 387 1758
rect 415 1762 419 1763
rect 415 1757 419 1758
rect 431 1762 435 1763
rect 431 1757 435 1758
rect 479 1762 483 1763
rect 479 1757 483 1758
rect 527 1762 531 1763
rect 527 1757 531 1758
rect 543 1762 547 1763
rect 543 1757 547 1758
rect 575 1762 579 1763
rect 575 1757 579 1758
rect 615 1762 619 1763
rect 615 1757 619 1758
rect 623 1762 627 1763
rect 623 1757 627 1758
rect 671 1762 675 1763
rect 671 1757 675 1758
rect 687 1762 691 1763
rect 687 1757 691 1758
rect 727 1762 731 1763
rect 727 1757 731 1758
rect 759 1762 763 1763
rect 759 1757 763 1758
rect 831 1762 835 1763
rect 831 1757 835 1758
rect 911 1762 915 1763
rect 911 1757 915 1758
rect 991 1762 995 1763
rect 991 1757 995 1758
rect 1095 1762 1099 1763
rect 1136 1761 1138 1781
rect 1192 1769 1194 1781
rect 1256 1769 1258 1781
rect 1320 1769 1322 1781
rect 1384 1769 1386 1781
rect 1456 1769 1458 1781
rect 1528 1769 1530 1781
rect 1608 1769 1610 1781
rect 1688 1769 1690 1781
rect 1768 1769 1770 1781
rect 1848 1769 1850 1781
rect 1928 1769 1930 1781
rect 2008 1769 2010 1781
rect 2072 1769 2074 1781
rect 1190 1768 1196 1769
rect 1190 1764 1191 1768
rect 1195 1764 1196 1768
rect 1190 1763 1196 1764
rect 1254 1768 1260 1769
rect 1254 1764 1255 1768
rect 1259 1764 1260 1768
rect 1254 1763 1260 1764
rect 1318 1768 1324 1769
rect 1318 1764 1319 1768
rect 1323 1764 1324 1768
rect 1318 1763 1324 1764
rect 1382 1768 1388 1769
rect 1382 1764 1383 1768
rect 1387 1764 1388 1768
rect 1382 1763 1388 1764
rect 1454 1768 1460 1769
rect 1454 1764 1455 1768
rect 1459 1764 1460 1768
rect 1454 1763 1460 1764
rect 1526 1768 1532 1769
rect 1526 1764 1527 1768
rect 1531 1764 1532 1768
rect 1526 1763 1532 1764
rect 1606 1768 1612 1769
rect 1606 1764 1607 1768
rect 1611 1764 1612 1768
rect 1606 1763 1612 1764
rect 1686 1768 1692 1769
rect 1686 1764 1687 1768
rect 1691 1764 1692 1768
rect 1686 1763 1692 1764
rect 1766 1768 1772 1769
rect 1766 1764 1767 1768
rect 1771 1764 1772 1768
rect 1766 1763 1772 1764
rect 1846 1768 1852 1769
rect 1846 1764 1847 1768
rect 1851 1764 1852 1768
rect 1846 1763 1852 1764
rect 1926 1768 1932 1769
rect 1926 1764 1927 1768
rect 1931 1764 1932 1768
rect 1926 1763 1932 1764
rect 2006 1768 2012 1769
rect 2006 1764 2007 1768
rect 2011 1764 2012 1768
rect 2006 1763 2012 1764
rect 2070 1768 2076 1769
rect 2070 1764 2071 1768
rect 2075 1764 2076 1768
rect 2070 1763 2076 1764
rect 2120 1761 2122 1781
rect 1095 1757 1099 1758
rect 1134 1760 1140 1761
rect 112 1754 114 1757
rect 230 1756 236 1757
rect 110 1753 116 1754
rect 110 1749 111 1753
rect 115 1749 116 1753
rect 230 1752 231 1756
rect 235 1752 236 1756
rect 230 1751 236 1752
rect 294 1756 300 1757
rect 294 1752 295 1756
rect 299 1752 300 1756
rect 294 1751 300 1752
rect 350 1756 356 1757
rect 350 1752 351 1756
rect 355 1752 356 1756
rect 350 1751 356 1752
rect 414 1756 420 1757
rect 414 1752 415 1756
rect 419 1752 420 1756
rect 414 1751 420 1752
rect 478 1756 484 1757
rect 478 1752 479 1756
rect 483 1752 484 1756
rect 478 1751 484 1752
rect 542 1756 548 1757
rect 542 1752 543 1756
rect 547 1752 548 1756
rect 542 1751 548 1752
rect 614 1756 620 1757
rect 614 1752 615 1756
rect 619 1752 620 1756
rect 614 1751 620 1752
rect 686 1756 692 1757
rect 686 1752 687 1756
rect 691 1752 692 1756
rect 686 1751 692 1752
rect 758 1756 764 1757
rect 758 1752 759 1756
rect 763 1752 764 1756
rect 758 1751 764 1752
rect 830 1756 836 1757
rect 830 1752 831 1756
rect 835 1752 836 1756
rect 830 1751 836 1752
rect 910 1756 916 1757
rect 910 1752 911 1756
rect 915 1752 916 1756
rect 910 1751 916 1752
rect 990 1756 996 1757
rect 990 1752 991 1756
rect 995 1752 996 1756
rect 1096 1754 1098 1757
rect 1134 1756 1135 1760
rect 1139 1756 1140 1760
rect 1134 1755 1140 1756
rect 2118 1760 2124 1761
rect 2118 1756 2119 1760
rect 2123 1756 2124 1760
rect 2118 1755 2124 1756
rect 990 1751 996 1752
rect 1094 1753 1100 1754
rect 110 1748 116 1749
rect 1094 1749 1095 1753
rect 1099 1749 1100 1753
rect 1094 1748 1100 1749
rect 1134 1743 1140 1744
rect 1134 1739 1135 1743
rect 1139 1739 1140 1743
rect 2118 1743 2124 1744
rect 1134 1738 1140 1739
rect 1190 1740 1196 1741
rect 110 1736 116 1737
rect 110 1732 111 1736
rect 115 1732 116 1736
rect 110 1731 116 1732
rect 1094 1736 1100 1737
rect 1094 1732 1095 1736
rect 1099 1732 1100 1736
rect 1136 1735 1138 1738
rect 1190 1736 1191 1740
rect 1195 1736 1196 1740
rect 1190 1735 1196 1736
rect 1254 1740 1260 1741
rect 1254 1736 1255 1740
rect 1259 1736 1260 1740
rect 1254 1735 1260 1736
rect 1318 1740 1324 1741
rect 1318 1736 1319 1740
rect 1323 1736 1324 1740
rect 1318 1735 1324 1736
rect 1382 1740 1388 1741
rect 1382 1736 1383 1740
rect 1387 1736 1388 1740
rect 1382 1735 1388 1736
rect 1454 1740 1460 1741
rect 1454 1736 1455 1740
rect 1459 1736 1460 1740
rect 1454 1735 1460 1736
rect 1526 1740 1532 1741
rect 1526 1736 1527 1740
rect 1531 1736 1532 1740
rect 1526 1735 1532 1736
rect 1606 1740 1612 1741
rect 1606 1736 1607 1740
rect 1611 1736 1612 1740
rect 1606 1735 1612 1736
rect 1686 1740 1692 1741
rect 1686 1736 1687 1740
rect 1691 1736 1692 1740
rect 1686 1735 1692 1736
rect 1766 1740 1772 1741
rect 1766 1736 1767 1740
rect 1771 1736 1772 1740
rect 1766 1735 1772 1736
rect 1846 1740 1852 1741
rect 1846 1736 1847 1740
rect 1851 1736 1852 1740
rect 1846 1735 1852 1736
rect 1926 1740 1932 1741
rect 1926 1736 1927 1740
rect 1931 1736 1932 1740
rect 1926 1735 1932 1736
rect 2006 1740 2012 1741
rect 2006 1736 2007 1740
rect 2011 1736 2012 1740
rect 2006 1735 2012 1736
rect 2070 1740 2076 1741
rect 2070 1736 2071 1740
rect 2075 1736 2076 1740
rect 2118 1739 2119 1743
rect 2123 1739 2124 1743
rect 2118 1738 2124 1739
rect 2070 1735 2076 1736
rect 2120 1735 2122 1738
rect 1094 1731 1100 1732
rect 1135 1734 1139 1735
rect 112 1707 114 1731
rect 230 1728 236 1729
rect 230 1724 231 1728
rect 235 1724 236 1728
rect 230 1723 236 1724
rect 294 1728 300 1729
rect 294 1724 295 1728
rect 299 1724 300 1728
rect 294 1723 300 1724
rect 350 1728 356 1729
rect 350 1724 351 1728
rect 355 1724 356 1728
rect 350 1723 356 1724
rect 414 1728 420 1729
rect 414 1724 415 1728
rect 419 1724 420 1728
rect 414 1723 420 1724
rect 478 1728 484 1729
rect 478 1724 479 1728
rect 483 1724 484 1728
rect 478 1723 484 1724
rect 542 1728 548 1729
rect 542 1724 543 1728
rect 547 1724 548 1728
rect 542 1723 548 1724
rect 614 1728 620 1729
rect 614 1724 615 1728
rect 619 1724 620 1728
rect 614 1723 620 1724
rect 686 1728 692 1729
rect 686 1724 687 1728
rect 691 1724 692 1728
rect 686 1723 692 1724
rect 758 1728 764 1729
rect 758 1724 759 1728
rect 763 1724 764 1728
rect 758 1723 764 1724
rect 830 1728 836 1729
rect 830 1724 831 1728
rect 835 1724 836 1728
rect 830 1723 836 1724
rect 910 1728 916 1729
rect 910 1724 911 1728
rect 915 1724 916 1728
rect 910 1723 916 1724
rect 990 1728 996 1729
rect 990 1724 991 1728
rect 995 1724 996 1728
rect 990 1723 996 1724
rect 232 1707 234 1723
rect 296 1707 298 1723
rect 352 1707 354 1723
rect 416 1707 418 1723
rect 480 1707 482 1723
rect 544 1707 546 1723
rect 616 1707 618 1723
rect 688 1707 690 1723
rect 760 1707 762 1723
rect 832 1707 834 1723
rect 912 1707 914 1723
rect 992 1707 994 1723
rect 1096 1707 1098 1731
rect 1135 1729 1139 1730
rect 1191 1734 1195 1735
rect 1191 1729 1195 1730
rect 1247 1734 1251 1735
rect 1247 1729 1251 1730
rect 1255 1734 1259 1735
rect 1255 1729 1259 1730
rect 1295 1734 1299 1735
rect 1295 1729 1299 1730
rect 1319 1734 1323 1735
rect 1319 1729 1323 1730
rect 1343 1734 1347 1735
rect 1343 1729 1347 1730
rect 1383 1734 1387 1735
rect 1383 1729 1387 1730
rect 1399 1734 1403 1735
rect 1399 1729 1403 1730
rect 1455 1734 1459 1735
rect 1455 1729 1459 1730
rect 1463 1734 1467 1735
rect 1463 1729 1467 1730
rect 1527 1734 1531 1735
rect 1527 1729 1531 1730
rect 1599 1734 1603 1735
rect 1599 1729 1603 1730
rect 1607 1734 1611 1735
rect 1607 1729 1611 1730
rect 1671 1734 1675 1735
rect 1671 1729 1675 1730
rect 1687 1734 1691 1735
rect 1687 1729 1691 1730
rect 1743 1734 1747 1735
rect 1743 1729 1747 1730
rect 1767 1734 1771 1735
rect 1767 1729 1771 1730
rect 1807 1734 1811 1735
rect 1807 1729 1811 1730
rect 1847 1734 1851 1735
rect 1847 1729 1851 1730
rect 1879 1734 1883 1735
rect 1879 1729 1883 1730
rect 1927 1734 1931 1735
rect 1927 1729 1931 1730
rect 1951 1734 1955 1735
rect 1951 1729 1955 1730
rect 2007 1734 2011 1735
rect 2007 1729 2011 1730
rect 2023 1734 2027 1735
rect 2023 1729 2027 1730
rect 2071 1734 2075 1735
rect 2071 1729 2075 1730
rect 2119 1734 2123 1735
rect 2119 1729 2123 1730
rect 1136 1726 1138 1729
rect 1246 1728 1252 1729
rect 1134 1725 1140 1726
rect 1134 1721 1135 1725
rect 1139 1721 1140 1725
rect 1246 1724 1247 1728
rect 1251 1724 1252 1728
rect 1246 1723 1252 1724
rect 1294 1728 1300 1729
rect 1294 1724 1295 1728
rect 1299 1724 1300 1728
rect 1294 1723 1300 1724
rect 1342 1728 1348 1729
rect 1342 1724 1343 1728
rect 1347 1724 1348 1728
rect 1342 1723 1348 1724
rect 1398 1728 1404 1729
rect 1398 1724 1399 1728
rect 1403 1724 1404 1728
rect 1398 1723 1404 1724
rect 1462 1728 1468 1729
rect 1462 1724 1463 1728
rect 1467 1724 1468 1728
rect 1462 1723 1468 1724
rect 1526 1728 1532 1729
rect 1526 1724 1527 1728
rect 1531 1724 1532 1728
rect 1526 1723 1532 1724
rect 1598 1728 1604 1729
rect 1598 1724 1599 1728
rect 1603 1724 1604 1728
rect 1598 1723 1604 1724
rect 1670 1728 1676 1729
rect 1670 1724 1671 1728
rect 1675 1724 1676 1728
rect 1670 1723 1676 1724
rect 1742 1728 1748 1729
rect 1742 1724 1743 1728
rect 1747 1724 1748 1728
rect 1742 1723 1748 1724
rect 1806 1728 1812 1729
rect 1806 1724 1807 1728
rect 1811 1724 1812 1728
rect 1806 1723 1812 1724
rect 1878 1728 1884 1729
rect 1878 1724 1879 1728
rect 1883 1724 1884 1728
rect 1878 1723 1884 1724
rect 1950 1728 1956 1729
rect 1950 1724 1951 1728
rect 1955 1724 1956 1728
rect 1950 1723 1956 1724
rect 2022 1728 2028 1729
rect 2022 1724 2023 1728
rect 2027 1724 2028 1728
rect 2022 1723 2028 1724
rect 2070 1728 2076 1729
rect 2070 1724 2071 1728
rect 2075 1724 2076 1728
rect 2120 1726 2122 1729
rect 2070 1723 2076 1724
rect 2118 1725 2124 1726
rect 1134 1720 1140 1721
rect 2118 1721 2119 1725
rect 2123 1721 2124 1725
rect 2118 1720 2124 1721
rect 1134 1708 1140 1709
rect 111 1706 115 1707
rect 111 1701 115 1702
rect 135 1706 139 1707
rect 135 1701 139 1702
rect 199 1706 203 1707
rect 199 1701 203 1702
rect 231 1706 235 1707
rect 231 1701 235 1702
rect 279 1706 283 1707
rect 279 1701 283 1702
rect 295 1706 299 1707
rect 295 1701 299 1702
rect 351 1706 355 1707
rect 351 1701 355 1702
rect 367 1706 371 1707
rect 367 1701 371 1702
rect 415 1706 419 1707
rect 415 1701 419 1702
rect 463 1706 467 1707
rect 463 1701 467 1702
rect 479 1706 483 1707
rect 479 1701 483 1702
rect 543 1706 547 1707
rect 543 1701 547 1702
rect 551 1706 555 1707
rect 551 1701 555 1702
rect 615 1706 619 1707
rect 615 1701 619 1702
rect 639 1706 643 1707
rect 639 1701 643 1702
rect 687 1706 691 1707
rect 687 1701 691 1702
rect 719 1706 723 1707
rect 719 1701 723 1702
rect 759 1706 763 1707
rect 759 1701 763 1702
rect 791 1706 795 1707
rect 791 1701 795 1702
rect 831 1706 835 1707
rect 831 1701 835 1702
rect 855 1706 859 1707
rect 855 1701 859 1702
rect 911 1706 915 1707
rect 911 1701 915 1702
rect 919 1706 923 1707
rect 919 1701 923 1702
rect 983 1706 987 1707
rect 983 1701 987 1702
rect 991 1706 995 1707
rect 991 1701 995 1702
rect 1047 1706 1051 1707
rect 1047 1701 1051 1702
rect 1095 1706 1099 1707
rect 1134 1704 1135 1708
rect 1139 1704 1140 1708
rect 1134 1703 1140 1704
rect 2118 1708 2124 1709
rect 2118 1704 2119 1708
rect 2123 1704 2124 1708
rect 2118 1703 2124 1704
rect 1095 1701 1099 1702
rect 112 1681 114 1701
rect 136 1689 138 1701
rect 200 1689 202 1701
rect 280 1689 282 1701
rect 368 1689 370 1701
rect 464 1689 466 1701
rect 552 1689 554 1701
rect 640 1689 642 1701
rect 720 1689 722 1701
rect 792 1689 794 1701
rect 856 1689 858 1701
rect 920 1689 922 1701
rect 984 1689 986 1701
rect 1048 1689 1050 1701
rect 134 1688 140 1689
rect 134 1684 135 1688
rect 139 1684 140 1688
rect 134 1683 140 1684
rect 198 1688 204 1689
rect 198 1684 199 1688
rect 203 1684 204 1688
rect 198 1683 204 1684
rect 278 1688 284 1689
rect 278 1684 279 1688
rect 283 1684 284 1688
rect 278 1683 284 1684
rect 366 1688 372 1689
rect 366 1684 367 1688
rect 371 1684 372 1688
rect 366 1683 372 1684
rect 462 1688 468 1689
rect 462 1684 463 1688
rect 467 1684 468 1688
rect 462 1683 468 1684
rect 550 1688 556 1689
rect 550 1684 551 1688
rect 555 1684 556 1688
rect 550 1683 556 1684
rect 638 1688 644 1689
rect 638 1684 639 1688
rect 643 1684 644 1688
rect 638 1683 644 1684
rect 718 1688 724 1689
rect 718 1684 719 1688
rect 723 1684 724 1688
rect 718 1683 724 1684
rect 790 1688 796 1689
rect 790 1684 791 1688
rect 795 1684 796 1688
rect 790 1683 796 1684
rect 854 1688 860 1689
rect 854 1684 855 1688
rect 859 1684 860 1688
rect 854 1683 860 1684
rect 918 1688 924 1689
rect 918 1684 919 1688
rect 923 1684 924 1688
rect 918 1683 924 1684
rect 982 1688 988 1689
rect 982 1684 983 1688
rect 987 1684 988 1688
rect 982 1683 988 1684
rect 1046 1688 1052 1689
rect 1046 1684 1047 1688
rect 1051 1684 1052 1688
rect 1046 1683 1052 1684
rect 1096 1681 1098 1701
rect 110 1680 116 1681
rect 110 1676 111 1680
rect 115 1676 116 1680
rect 110 1675 116 1676
rect 1094 1680 1100 1681
rect 1094 1676 1095 1680
rect 1099 1676 1100 1680
rect 1136 1679 1138 1703
rect 1246 1700 1252 1701
rect 1246 1696 1247 1700
rect 1251 1696 1252 1700
rect 1246 1695 1252 1696
rect 1294 1700 1300 1701
rect 1294 1696 1295 1700
rect 1299 1696 1300 1700
rect 1294 1695 1300 1696
rect 1342 1700 1348 1701
rect 1342 1696 1343 1700
rect 1347 1696 1348 1700
rect 1342 1695 1348 1696
rect 1398 1700 1404 1701
rect 1398 1696 1399 1700
rect 1403 1696 1404 1700
rect 1398 1695 1404 1696
rect 1462 1700 1468 1701
rect 1462 1696 1463 1700
rect 1467 1696 1468 1700
rect 1462 1695 1468 1696
rect 1526 1700 1532 1701
rect 1526 1696 1527 1700
rect 1531 1696 1532 1700
rect 1526 1695 1532 1696
rect 1598 1700 1604 1701
rect 1598 1696 1599 1700
rect 1603 1696 1604 1700
rect 1598 1695 1604 1696
rect 1670 1700 1676 1701
rect 1670 1696 1671 1700
rect 1675 1696 1676 1700
rect 1670 1695 1676 1696
rect 1742 1700 1748 1701
rect 1742 1696 1743 1700
rect 1747 1696 1748 1700
rect 1742 1695 1748 1696
rect 1806 1700 1812 1701
rect 1806 1696 1807 1700
rect 1811 1696 1812 1700
rect 1806 1695 1812 1696
rect 1878 1700 1884 1701
rect 1878 1696 1879 1700
rect 1883 1696 1884 1700
rect 1878 1695 1884 1696
rect 1950 1700 1956 1701
rect 1950 1696 1951 1700
rect 1955 1696 1956 1700
rect 1950 1695 1956 1696
rect 2022 1700 2028 1701
rect 2022 1696 2023 1700
rect 2027 1696 2028 1700
rect 2022 1695 2028 1696
rect 2070 1700 2076 1701
rect 2070 1696 2071 1700
rect 2075 1696 2076 1700
rect 2070 1695 2076 1696
rect 1248 1679 1250 1695
rect 1296 1679 1298 1695
rect 1344 1679 1346 1695
rect 1400 1679 1402 1695
rect 1464 1679 1466 1695
rect 1528 1679 1530 1695
rect 1600 1679 1602 1695
rect 1672 1679 1674 1695
rect 1744 1679 1746 1695
rect 1808 1679 1810 1695
rect 1880 1679 1882 1695
rect 1952 1679 1954 1695
rect 2024 1679 2026 1695
rect 2072 1679 2074 1695
rect 2120 1679 2122 1703
rect 1094 1675 1100 1676
rect 1135 1678 1139 1679
rect 1135 1673 1139 1674
rect 1247 1678 1251 1679
rect 1247 1673 1251 1674
rect 1263 1678 1267 1679
rect 1263 1673 1267 1674
rect 1295 1678 1299 1679
rect 1295 1673 1299 1674
rect 1303 1678 1307 1679
rect 1303 1673 1307 1674
rect 1343 1678 1347 1679
rect 1343 1673 1347 1674
rect 1391 1678 1395 1679
rect 1391 1673 1395 1674
rect 1399 1678 1403 1679
rect 1399 1673 1403 1674
rect 1447 1678 1451 1679
rect 1447 1673 1451 1674
rect 1463 1678 1467 1679
rect 1463 1673 1467 1674
rect 1503 1678 1507 1679
rect 1503 1673 1507 1674
rect 1527 1678 1531 1679
rect 1527 1673 1531 1674
rect 1567 1678 1571 1679
rect 1567 1673 1571 1674
rect 1599 1678 1603 1679
rect 1599 1673 1603 1674
rect 1631 1678 1635 1679
rect 1631 1673 1635 1674
rect 1671 1678 1675 1679
rect 1671 1673 1675 1674
rect 1695 1678 1699 1679
rect 1695 1673 1699 1674
rect 1743 1678 1747 1679
rect 1743 1673 1747 1674
rect 1759 1678 1763 1679
rect 1759 1673 1763 1674
rect 1807 1678 1811 1679
rect 1807 1673 1811 1674
rect 1831 1678 1835 1679
rect 1831 1673 1835 1674
rect 1879 1678 1883 1679
rect 1879 1673 1883 1674
rect 1911 1678 1915 1679
rect 1911 1673 1915 1674
rect 1951 1678 1955 1679
rect 1951 1673 1955 1674
rect 1999 1678 2003 1679
rect 1999 1673 2003 1674
rect 2023 1678 2027 1679
rect 2023 1673 2027 1674
rect 2071 1678 2075 1679
rect 2071 1673 2075 1674
rect 2119 1678 2123 1679
rect 2119 1673 2123 1674
rect 110 1663 116 1664
rect 110 1659 111 1663
rect 115 1659 116 1663
rect 1094 1663 1100 1664
rect 110 1658 116 1659
rect 134 1660 140 1661
rect 112 1651 114 1658
rect 134 1656 135 1660
rect 139 1656 140 1660
rect 134 1655 140 1656
rect 198 1660 204 1661
rect 198 1656 199 1660
rect 203 1656 204 1660
rect 198 1655 204 1656
rect 278 1660 284 1661
rect 278 1656 279 1660
rect 283 1656 284 1660
rect 278 1655 284 1656
rect 366 1660 372 1661
rect 366 1656 367 1660
rect 371 1656 372 1660
rect 366 1655 372 1656
rect 462 1660 468 1661
rect 462 1656 463 1660
rect 467 1656 468 1660
rect 462 1655 468 1656
rect 550 1660 556 1661
rect 550 1656 551 1660
rect 555 1656 556 1660
rect 550 1655 556 1656
rect 638 1660 644 1661
rect 638 1656 639 1660
rect 643 1656 644 1660
rect 638 1655 644 1656
rect 718 1660 724 1661
rect 718 1656 719 1660
rect 723 1656 724 1660
rect 718 1655 724 1656
rect 790 1660 796 1661
rect 790 1656 791 1660
rect 795 1656 796 1660
rect 790 1655 796 1656
rect 854 1660 860 1661
rect 854 1656 855 1660
rect 859 1656 860 1660
rect 854 1655 860 1656
rect 918 1660 924 1661
rect 918 1656 919 1660
rect 923 1656 924 1660
rect 918 1655 924 1656
rect 982 1660 988 1661
rect 982 1656 983 1660
rect 987 1656 988 1660
rect 982 1655 988 1656
rect 1046 1660 1052 1661
rect 1046 1656 1047 1660
rect 1051 1656 1052 1660
rect 1094 1659 1095 1663
rect 1099 1659 1100 1663
rect 1094 1658 1100 1659
rect 1046 1655 1052 1656
rect 136 1651 138 1655
rect 200 1651 202 1655
rect 280 1651 282 1655
rect 368 1651 370 1655
rect 464 1651 466 1655
rect 552 1651 554 1655
rect 640 1651 642 1655
rect 720 1651 722 1655
rect 792 1651 794 1655
rect 856 1651 858 1655
rect 920 1651 922 1655
rect 984 1651 986 1655
rect 1048 1651 1050 1655
rect 1096 1651 1098 1658
rect 1136 1653 1138 1673
rect 1264 1661 1266 1673
rect 1304 1661 1306 1673
rect 1344 1661 1346 1673
rect 1392 1661 1394 1673
rect 1448 1661 1450 1673
rect 1504 1661 1506 1673
rect 1568 1661 1570 1673
rect 1632 1661 1634 1673
rect 1696 1661 1698 1673
rect 1760 1661 1762 1673
rect 1832 1661 1834 1673
rect 1912 1661 1914 1673
rect 2000 1661 2002 1673
rect 2072 1661 2074 1673
rect 1262 1660 1268 1661
rect 1262 1656 1263 1660
rect 1267 1656 1268 1660
rect 1262 1655 1268 1656
rect 1302 1660 1308 1661
rect 1302 1656 1303 1660
rect 1307 1656 1308 1660
rect 1302 1655 1308 1656
rect 1342 1660 1348 1661
rect 1342 1656 1343 1660
rect 1347 1656 1348 1660
rect 1342 1655 1348 1656
rect 1390 1660 1396 1661
rect 1390 1656 1391 1660
rect 1395 1656 1396 1660
rect 1390 1655 1396 1656
rect 1446 1660 1452 1661
rect 1446 1656 1447 1660
rect 1451 1656 1452 1660
rect 1446 1655 1452 1656
rect 1502 1660 1508 1661
rect 1502 1656 1503 1660
rect 1507 1656 1508 1660
rect 1502 1655 1508 1656
rect 1566 1660 1572 1661
rect 1566 1656 1567 1660
rect 1571 1656 1572 1660
rect 1566 1655 1572 1656
rect 1630 1660 1636 1661
rect 1630 1656 1631 1660
rect 1635 1656 1636 1660
rect 1630 1655 1636 1656
rect 1694 1660 1700 1661
rect 1694 1656 1695 1660
rect 1699 1656 1700 1660
rect 1694 1655 1700 1656
rect 1758 1660 1764 1661
rect 1758 1656 1759 1660
rect 1763 1656 1764 1660
rect 1758 1655 1764 1656
rect 1830 1660 1836 1661
rect 1830 1656 1831 1660
rect 1835 1656 1836 1660
rect 1830 1655 1836 1656
rect 1910 1660 1916 1661
rect 1910 1656 1911 1660
rect 1915 1656 1916 1660
rect 1910 1655 1916 1656
rect 1998 1660 2004 1661
rect 1998 1656 1999 1660
rect 2003 1656 2004 1660
rect 1998 1655 2004 1656
rect 2070 1660 2076 1661
rect 2070 1656 2071 1660
rect 2075 1656 2076 1660
rect 2070 1655 2076 1656
rect 2120 1653 2122 1673
rect 1134 1652 1140 1653
rect 111 1650 115 1651
rect 111 1645 115 1646
rect 135 1650 139 1651
rect 135 1645 139 1646
rect 183 1650 187 1651
rect 183 1645 187 1646
rect 199 1650 203 1651
rect 199 1645 203 1646
rect 263 1650 267 1651
rect 263 1645 267 1646
rect 279 1650 283 1651
rect 279 1645 283 1646
rect 343 1650 347 1651
rect 343 1645 347 1646
rect 367 1650 371 1651
rect 367 1645 371 1646
rect 423 1650 427 1651
rect 423 1645 427 1646
rect 463 1650 467 1651
rect 463 1645 467 1646
rect 503 1650 507 1651
rect 503 1645 507 1646
rect 551 1650 555 1651
rect 551 1645 555 1646
rect 583 1650 587 1651
rect 583 1645 587 1646
rect 639 1650 643 1651
rect 639 1645 643 1646
rect 655 1650 659 1651
rect 655 1645 659 1646
rect 719 1650 723 1651
rect 719 1645 723 1646
rect 727 1650 731 1651
rect 727 1645 731 1646
rect 791 1650 795 1651
rect 791 1645 795 1646
rect 847 1650 851 1651
rect 847 1645 851 1646
rect 855 1650 859 1651
rect 855 1645 859 1646
rect 903 1650 907 1651
rect 903 1645 907 1646
rect 919 1650 923 1651
rect 919 1645 923 1646
rect 959 1650 963 1651
rect 959 1645 963 1646
rect 983 1650 987 1651
rect 983 1645 987 1646
rect 1007 1650 1011 1651
rect 1007 1645 1011 1646
rect 1047 1650 1051 1651
rect 1047 1645 1051 1646
rect 1095 1650 1099 1651
rect 1134 1648 1135 1652
rect 1139 1648 1140 1652
rect 1134 1647 1140 1648
rect 2118 1652 2124 1653
rect 2118 1648 2119 1652
rect 2123 1648 2124 1652
rect 2118 1647 2124 1648
rect 1095 1645 1099 1646
rect 112 1642 114 1645
rect 134 1644 140 1645
rect 110 1641 116 1642
rect 110 1637 111 1641
rect 115 1637 116 1641
rect 134 1640 135 1644
rect 139 1640 140 1644
rect 134 1639 140 1640
rect 182 1644 188 1645
rect 182 1640 183 1644
rect 187 1640 188 1644
rect 182 1639 188 1640
rect 262 1644 268 1645
rect 262 1640 263 1644
rect 267 1640 268 1644
rect 262 1639 268 1640
rect 342 1644 348 1645
rect 342 1640 343 1644
rect 347 1640 348 1644
rect 342 1639 348 1640
rect 422 1644 428 1645
rect 422 1640 423 1644
rect 427 1640 428 1644
rect 422 1639 428 1640
rect 502 1644 508 1645
rect 502 1640 503 1644
rect 507 1640 508 1644
rect 502 1639 508 1640
rect 582 1644 588 1645
rect 582 1640 583 1644
rect 587 1640 588 1644
rect 582 1639 588 1640
rect 654 1644 660 1645
rect 654 1640 655 1644
rect 659 1640 660 1644
rect 654 1639 660 1640
rect 726 1644 732 1645
rect 726 1640 727 1644
rect 731 1640 732 1644
rect 726 1639 732 1640
rect 790 1644 796 1645
rect 790 1640 791 1644
rect 795 1640 796 1644
rect 790 1639 796 1640
rect 846 1644 852 1645
rect 846 1640 847 1644
rect 851 1640 852 1644
rect 846 1639 852 1640
rect 902 1644 908 1645
rect 902 1640 903 1644
rect 907 1640 908 1644
rect 902 1639 908 1640
rect 958 1644 964 1645
rect 958 1640 959 1644
rect 963 1640 964 1644
rect 958 1639 964 1640
rect 1006 1644 1012 1645
rect 1006 1640 1007 1644
rect 1011 1640 1012 1644
rect 1006 1639 1012 1640
rect 1046 1644 1052 1645
rect 1046 1640 1047 1644
rect 1051 1640 1052 1644
rect 1096 1642 1098 1645
rect 1046 1639 1052 1640
rect 1094 1641 1100 1642
rect 110 1636 116 1637
rect 1094 1637 1095 1641
rect 1099 1637 1100 1641
rect 1094 1636 1100 1637
rect 1134 1635 1140 1636
rect 1134 1631 1135 1635
rect 1139 1631 1140 1635
rect 2118 1635 2124 1636
rect 1134 1630 1140 1631
rect 1262 1632 1268 1633
rect 110 1624 116 1625
rect 110 1620 111 1624
rect 115 1620 116 1624
rect 110 1619 116 1620
rect 1094 1624 1100 1625
rect 1094 1620 1095 1624
rect 1099 1620 1100 1624
rect 1094 1619 1100 1620
rect 112 1599 114 1619
rect 134 1616 140 1617
rect 134 1612 135 1616
rect 139 1612 140 1616
rect 134 1611 140 1612
rect 182 1616 188 1617
rect 182 1612 183 1616
rect 187 1612 188 1616
rect 182 1611 188 1612
rect 262 1616 268 1617
rect 262 1612 263 1616
rect 267 1612 268 1616
rect 262 1611 268 1612
rect 342 1616 348 1617
rect 342 1612 343 1616
rect 347 1612 348 1616
rect 342 1611 348 1612
rect 422 1616 428 1617
rect 422 1612 423 1616
rect 427 1612 428 1616
rect 422 1611 428 1612
rect 502 1616 508 1617
rect 502 1612 503 1616
rect 507 1612 508 1616
rect 502 1611 508 1612
rect 582 1616 588 1617
rect 582 1612 583 1616
rect 587 1612 588 1616
rect 582 1611 588 1612
rect 654 1616 660 1617
rect 654 1612 655 1616
rect 659 1612 660 1616
rect 654 1611 660 1612
rect 726 1616 732 1617
rect 726 1612 727 1616
rect 731 1612 732 1616
rect 726 1611 732 1612
rect 790 1616 796 1617
rect 790 1612 791 1616
rect 795 1612 796 1616
rect 790 1611 796 1612
rect 846 1616 852 1617
rect 846 1612 847 1616
rect 851 1612 852 1616
rect 846 1611 852 1612
rect 902 1616 908 1617
rect 902 1612 903 1616
rect 907 1612 908 1616
rect 902 1611 908 1612
rect 958 1616 964 1617
rect 958 1612 959 1616
rect 963 1612 964 1616
rect 958 1611 964 1612
rect 1006 1616 1012 1617
rect 1006 1612 1007 1616
rect 1011 1612 1012 1616
rect 1006 1611 1012 1612
rect 1046 1616 1052 1617
rect 1046 1612 1047 1616
rect 1051 1612 1052 1616
rect 1046 1611 1052 1612
rect 136 1599 138 1611
rect 184 1599 186 1611
rect 264 1599 266 1611
rect 344 1599 346 1611
rect 424 1599 426 1611
rect 504 1599 506 1611
rect 584 1599 586 1611
rect 656 1599 658 1611
rect 728 1599 730 1611
rect 792 1599 794 1611
rect 848 1599 850 1611
rect 904 1599 906 1611
rect 960 1599 962 1611
rect 1008 1599 1010 1611
rect 1048 1599 1050 1611
rect 1096 1599 1098 1619
rect 1136 1615 1138 1630
rect 1262 1628 1263 1632
rect 1267 1628 1268 1632
rect 1262 1627 1268 1628
rect 1302 1632 1308 1633
rect 1302 1628 1303 1632
rect 1307 1628 1308 1632
rect 1302 1627 1308 1628
rect 1342 1632 1348 1633
rect 1342 1628 1343 1632
rect 1347 1628 1348 1632
rect 1342 1627 1348 1628
rect 1390 1632 1396 1633
rect 1390 1628 1391 1632
rect 1395 1628 1396 1632
rect 1390 1627 1396 1628
rect 1446 1632 1452 1633
rect 1446 1628 1447 1632
rect 1451 1628 1452 1632
rect 1446 1627 1452 1628
rect 1502 1632 1508 1633
rect 1502 1628 1503 1632
rect 1507 1628 1508 1632
rect 1502 1627 1508 1628
rect 1566 1632 1572 1633
rect 1566 1628 1567 1632
rect 1571 1628 1572 1632
rect 1566 1627 1572 1628
rect 1630 1632 1636 1633
rect 1630 1628 1631 1632
rect 1635 1628 1636 1632
rect 1630 1627 1636 1628
rect 1694 1632 1700 1633
rect 1694 1628 1695 1632
rect 1699 1628 1700 1632
rect 1694 1627 1700 1628
rect 1758 1632 1764 1633
rect 1758 1628 1759 1632
rect 1763 1628 1764 1632
rect 1758 1627 1764 1628
rect 1830 1632 1836 1633
rect 1830 1628 1831 1632
rect 1835 1628 1836 1632
rect 1830 1627 1836 1628
rect 1910 1632 1916 1633
rect 1910 1628 1911 1632
rect 1915 1628 1916 1632
rect 1910 1627 1916 1628
rect 1998 1632 2004 1633
rect 1998 1628 1999 1632
rect 2003 1628 2004 1632
rect 1998 1627 2004 1628
rect 2070 1632 2076 1633
rect 2070 1628 2071 1632
rect 2075 1628 2076 1632
rect 2118 1631 2119 1635
rect 2123 1631 2124 1635
rect 2118 1630 2124 1631
rect 2070 1627 2076 1628
rect 1264 1615 1266 1627
rect 1304 1615 1306 1627
rect 1344 1615 1346 1627
rect 1392 1615 1394 1627
rect 1448 1615 1450 1627
rect 1504 1615 1506 1627
rect 1568 1615 1570 1627
rect 1632 1615 1634 1627
rect 1696 1615 1698 1627
rect 1760 1615 1762 1627
rect 1832 1615 1834 1627
rect 1912 1615 1914 1627
rect 2000 1615 2002 1627
rect 2072 1615 2074 1627
rect 2120 1615 2122 1630
rect 1135 1614 1139 1615
rect 1135 1609 1139 1610
rect 1159 1614 1163 1615
rect 1159 1609 1163 1610
rect 1215 1614 1219 1615
rect 1215 1609 1219 1610
rect 1263 1614 1267 1615
rect 1263 1609 1267 1610
rect 1303 1614 1307 1615
rect 1303 1609 1307 1610
rect 1343 1614 1347 1615
rect 1343 1609 1347 1610
rect 1383 1614 1387 1615
rect 1383 1609 1387 1610
rect 1391 1614 1395 1615
rect 1391 1609 1395 1610
rect 1447 1614 1451 1615
rect 1447 1609 1451 1610
rect 1463 1614 1467 1615
rect 1463 1609 1467 1610
rect 1503 1614 1507 1615
rect 1503 1609 1507 1610
rect 1543 1614 1547 1615
rect 1543 1609 1547 1610
rect 1567 1614 1571 1615
rect 1567 1609 1571 1610
rect 1623 1614 1627 1615
rect 1623 1609 1627 1610
rect 1631 1614 1635 1615
rect 1631 1609 1635 1610
rect 1695 1614 1699 1615
rect 1695 1609 1699 1610
rect 1711 1614 1715 1615
rect 1711 1609 1715 1610
rect 1759 1614 1763 1615
rect 1759 1609 1763 1610
rect 1799 1614 1803 1615
rect 1799 1609 1803 1610
rect 1831 1614 1835 1615
rect 1831 1609 1835 1610
rect 1887 1614 1891 1615
rect 1887 1609 1891 1610
rect 1911 1614 1915 1615
rect 1911 1609 1915 1610
rect 1983 1614 1987 1615
rect 1983 1609 1987 1610
rect 1999 1614 2003 1615
rect 1999 1609 2003 1610
rect 2071 1614 2075 1615
rect 2071 1609 2075 1610
rect 2119 1614 2123 1615
rect 2119 1609 2123 1610
rect 1136 1606 1138 1609
rect 1158 1608 1164 1609
rect 1134 1605 1140 1606
rect 1134 1601 1135 1605
rect 1139 1601 1140 1605
rect 1158 1604 1159 1608
rect 1163 1604 1164 1608
rect 1158 1603 1164 1604
rect 1214 1608 1220 1609
rect 1214 1604 1215 1608
rect 1219 1604 1220 1608
rect 1214 1603 1220 1604
rect 1302 1608 1308 1609
rect 1302 1604 1303 1608
rect 1307 1604 1308 1608
rect 1302 1603 1308 1604
rect 1382 1608 1388 1609
rect 1382 1604 1383 1608
rect 1387 1604 1388 1608
rect 1382 1603 1388 1604
rect 1462 1608 1468 1609
rect 1462 1604 1463 1608
rect 1467 1604 1468 1608
rect 1462 1603 1468 1604
rect 1542 1608 1548 1609
rect 1542 1604 1543 1608
rect 1547 1604 1548 1608
rect 1542 1603 1548 1604
rect 1622 1608 1628 1609
rect 1622 1604 1623 1608
rect 1627 1604 1628 1608
rect 1622 1603 1628 1604
rect 1710 1608 1716 1609
rect 1710 1604 1711 1608
rect 1715 1604 1716 1608
rect 1710 1603 1716 1604
rect 1798 1608 1804 1609
rect 1798 1604 1799 1608
rect 1803 1604 1804 1608
rect 1798 1603 1804 1604
rect 1886 1608 1892 1609
rect 1886 1604 1887 1608
rect 1891 1604 1892 1608
rect 1886 1603 1892 1604
rect 1982 1608 1988 1609
rect 1982 1604 1983 1608
rect 1987 1604 1988 1608
rect 1982 1603 1988 1604
rect 2070 1608 2076 1609
rect 2070 1604 2071 1608
rect 2075 1604 2076 1608
rect 2120 1606 2122 1609
rect 2070 1603 2076 1604
rect 2118 1605 2124 1606
rect 1134 1600 1140 1601
rect 2118 1601 2119 1605
rect 2123 1601 2124 1605
rect 2118 1600 2124 1601
rect 111 1598 115 1599
rect 111 1593 115 1594
rect 135 1598 139 1599
rect 135 1593 139 1594
rect 175 1598 179 1599
rect 175 1593 179 1594
rect 183 1598 187 1599
rect 183 1593 187 1594
rect 231 1598 235 1599
rect 231 1593 235 1594
rect 263 1598 267 1599
rect 263 1593 267 1594
rect 303 1598 307 1599
rect 303 1593 307 1594
rect 343 1598 347 1599
rect 343 1593 347 1594
rect 375 1598 379 1599
rect 375 1593 379 1594
rect 423 1598 427 1599
rect 423 1593 427 1594
rect 455 1598 459 1599
rect 455 1593 459 1594
rect 503 1598 507 1599
rect 503 1593 507 1594
rect 527 1598 531 1599
rect 527 1593 531 1594
rect 583 1598 587 1599
rect 583 1593 587 1594
rect 599 1598 603 1599
rect 599 1593 603 1594
rect 655 1598 659 1599
rect 655 1593 659 1594
rect 671 1598 675 1599
rect 671 1593 675 1594
rect 727 1598 731 1599
rect 727 1593 731 1594
rect 743 1598 747 1599
rect 743 1593 747 1594
rect 791 1598 795 1599
rect 791 1593 795 1594
rect 815 1598 819 1599
rect 815 1593 819 1594
rect 847 1598 851 1599
rect 847 1593 851 1594
rect 887 1598 891 1599
rect 887 1593 891 1594
rect 903 1598 907 1599
rect 903 1593 907 1594
rect 959 1598 963 1599
rect 959 1593 963 1594
rect 1007 1598 1011 1599
rect 1007 1593 1011 1594
rect 1047 1598 1051 1599
rect 1047 1593 1051 1594
rect 1095 1598 1099 1599
rect 1095 1593 1099 1594
rect 112 1573 114 1593
rect 136 1581 138 1593
rect 176 1581 178 1593
rect 232 1581 234 1593
rect 304 1581 306 1593
rect 376 1581 378 1593
rect 456 1581 458 1593
rect 528 1581 530 1593
rect 600 1581 602 1593
rect 672 1581 674 1593
rect 744 1581 746 1593
rect 816 1581 818 1593
rect 888 1581 890 1593
rect 134 1580 140 1581
rect 134 1576 135 1580
rect 139 1576 140 1580
rect 134 1575 140 1576
rect 174 1580 180 1581
rect 174 1576 175 1580
rect 179 1576 180 1580
rect 174 1575 180 1576
rect 230 1580 236 1581
rect 230 1576 231 1580
rect 235 1576 236 1580
rect 230 1575 236 1576
rect 302 1580 308 1581
rect 302 1576 303 1580
rect 307 1576 308 1580
rect 302 1575 308 1576
rect 374 1580 380 1581
rect 374 1576 375 1580
rect 379 1576 380 1580
rect 374 1575 380 1576
rect 454 1580 460 1581
rect 454 1576 455 1580
rect 459 1576 460 1580
rect 454 1575 460 1576
rect 526 1580 532 1581
rect 526 1576 527 1580
rect 531 1576 532 1580
rect 526 1575 532 1576
rect 598 1580 604 1581
rect 598 1576 599 1580
rect 603 1576 604 1580
rect 598 1575 604 1576
rect 670 1580 676 1581
rect 670 1576 671 1580
rect 675 1576 676 1580
rect 670 1575 676 1576
rect 742 1580 748 1581
rect 742 1576 743 1580
rect 747 1576 748 1580
rect 742 1575 748 1576
rect 814 1580 820 1581
rect 814 1576 815 1580
rect 819 1576 820 1580
rect 814 1575 820 1576
rect 886 1580 892 1581
rect 886 1576 887 1580
rect 891 1576 892 1580
rect 886 1575 892 1576
rect 1096 1573 1098 1593
rect 1134 1588 1140 1589
rect 1134 1584 1135 1588
rect 1139 1584 1140 1588
rect 1134 1583 1140 1584
rect 2118 1588 2124 1589
rect 2118 1584 2119 1588
rect 2123 1584 2124 1588
rect 2118 1583 2124 1584
rect 110 1572 116 1573
rect 110 1568 111 1572
rect 115 1568 116 1572
rect 110 1567 116 1568
rect 1094 1572 1100 1573
rect 1094 1568 1095 1572
rect 1099 1568 1100 1572
rect 1094 1567 1100 1568
rect 1136 1563 1138 1583
rect 1158 1580 1164 1581
rect 1158 1576 1159 1580
rect 1163 1576 1164 1580
rect 1158 1575 1164 1576
rect 1214 1580 1220 1581
rect 1214 1576 1215 1580
rect 1219 1576 1220 1580
rect 1214 1575 1220 1576
rect 1302 1580 1308 1581
rect 1302 1576 1303 1580
rect 1307 1576 1308 1580
rect 1302 1575 1308 1576
rect 1382 1580 1388 1581
rect 1382 1576 1383 1580
rect 1387 1576 1388 1580
rect 1382 1575 1388 1576
rect 1462 1580 1468 1581
rect 1462 1576 1463 1580
rect 1467 1576 1468 1580
rect 1462 1575 1468 1576
rect 1542 1580 1548 1581
rect 1542 1576 1543 1580
rect 1547 1576 1548 1580
rect 1542 1575 1548 1576
rect 1622 1580 1628 1581
rect 1622 1576 1623 1580
rect 1627 1576 1628 1580
rect 1622 1575 1628 1576
rect 1710 1580 1716 1581
rect 1710 1576 1711 1580
rect 1715 1576 1716 1580
rect 1710 1575 1716 1576
rect 1798 1580 1804 1581
rect 1798 1576 1799 1580
rect 1803 1576 1804 1580
rect 1798 1575 1804 1576
rect 1886 1580 1892 1581
rect 1886 1576 1887 1580
rect 1891 1576 1892 1580
rect 1886 1575 1892 1576
rect 1982 1580 1988 1581
rect 1982 1576 1983 1580
rect 1987 1576 1988 1580
rect 1982 1575 1988 1576
rect 2070 1580 2076 1581
rect 2070 1576 2071 1580
rect 2075 1576 2076 1580
rect 2070 1575 2076 1576
rect 1160 1563 1162 1575
rect 1216 1563 1218 1575
rect 1304 1563 1306 1575
rect 1384 1563 1386 1575
rect 1464 1563 1466 1575
rect 1544 1563 1546 1575
rect 1624 1563 1626 1575
rect 1712 1563 1714 1575
rect 1800 1563 1802 1575
rect 1888 1563 1890 1575
rect 1984 1563 1986 1575
rect 2072 1563 2074 1575
rect 2120 1563 2122 1583
rect 1135 1562 1139 1563
rect 1135 1557 1139 1558
rect 1159 1562 1163 1563
rect 1159 1557 1163 1558
rect 1199 1562 1203 1563
rect 1199 1557 1203 1558
rect 1215 1562 1219 1563
rect 1215 1557 1219 1558
rect 1247 1562 1251 1563
rect 1247 1557 1251 1558
rect 1303 1562 1307 1563
rect 1303 1557 1307 1558
rect 1319 1562 1323 1563
rect 1319 1557 1323 1558
rect 1383 1562 1387 1563
rect 1383 1557 1387 1558
rect 1399 1562 1403 1563
rect 1399 1557 1403 1558
rect 1463 1562 1467 1563
rect 1463 1557 1467 1558
rect 1479 1562 1483 1563
rect 1479 1557 1483 1558
rect 1543 1562 1547 1563
rect 1543 1557 1547 1558
rect 1559 1562 1563 1563
rect 1559 1557 1563 1558
rect 1623 1562 1627 1563
rect 1623 1557 1627 1558
rect 1647 1562 1651 1563
rect 1647 1557 1651 1558
rect 1711 1562 1715 1563
rect 1711 1557 1715 1558
rect 1735 1562 1739 1563
rect 1735 1557 1739 1558
rect 1799 1562 1803 1563
rect 1799 1557 1803 1558
rect 1823 1562 1827 1563
rect 1823 1557 1827 1558
rect 1887 1562 1891 1563
rect 1887 1557 1891 1558
rect 1911 1562 1915 1563
rect 1911 1557 1915 1558
rect 1983 1562 1987 1563
rect 1983 1557 1987 1558
rect 1999 1562 2003 1563
rect 1999 1557 2003 1558
rect 2071 1562 2075 1563
rect 2071 1557 2075 1558
rect 2119 1562 2123 1563
rect 2119 1557 2123 1558
rect 110 1555 116 1556
rect 110 1551 111 1555
rect 115 1551 116 1555
rect 1094 1555 1100 1556
rect 110 1550 116 1551
rect 134 1552 140 1553
rect 112 1547 114 1550
rect 134 1548 135 1552
rect 139 1548 140 1552
rect 134 1547 140 1548
rect 174 1552 180 1553
rect 174 1548 175 1552
rect 179 1548 180 1552
rect 174 1547 180 1548
rect 230 1552 236 1553
rect 230 1548 231 1552
rect 235 1548 236 1552
rect 230 1547 236 1548
rect 302 1552 308 1553
rect 302 1548 303 1552
rect 307 1548 308 1552
rect 302 1547 308 1548
rect 374 1552 380 1553
rect 374 1548 375 1552
rect 379 1548 380 1552
rect 374 1547 380 1548
rect 454 1552 460 1553
rect 454 1548 455 1552
rect 459 1548 460 1552
rect 454 1547 460 1548
rect 526 1552 532 1553
rect 526 1548 527 1552
rect 531 1548 532 1552
rect 526 1547 532 1548
rect 598 1552 604 1553
rect 598 1548 599 1552
rect 603 1548 604 1552
rect 598 1547 604 1548
rect 670 1552 676 1553
rect 670 1548 671 1552
rect 675 1548 676 1552
rect 670 1547 676 1548
rect 742 1552 748 1553
rect 742 1548 743 1552
rect 747 1548 748 1552
rect 742 1547 748 1548
rect 814 1552 820 1553
rect 814 1548 815 1552
rect 819 1548 820 1552
rect 814 1547 820 1548
rect 886 1552 892 1553
rect 886 1548 887 1552
rect 891 1548 892 1552
rect 1094 1551 1095 1555
rect 1099 1551 1100 1555
rect 1094 1550 1100 1551
rect 886 1547 892 1548
rect 1096 1547 1098 1550
rect 111 1546 115 1547
rect 111 1541 115 1542
rect 135 1546 139 1547
rect 135 1541 139 1542
rect 175 1546 179 1547
rect 175 1541 179 1542
rect 231 1546 235 1547
rect 231 1541 235 1542
rect 303 1546 307 1547
rect 303 1541 307 1542
rect 311 1546 315 1547
rect 311 1541 315 1542
rect 375 1546 379 1547
rect 375 1541 379 1542
rect 391 1546 395 1547
rect 391 1541 395 1542
rect 455 1546 459 1547
rect 455 1541 459 1542
rect 479 1546 483 1547
rect 479 1541 483 1542
rect 527 1546 531 1547
rect 527 1541 531 1542
rect 567 1546 571 1547
rect 567 1541 571 1542
rect 599 1546 603 1547
rect 599 1541 603 1542
rect 655 1546 659 1547
rect 655 1541 659 1542
rect 671 1546 675 1547
rect 671 1541 675 1542
rect 743 1546 747 1547
rect 743 1541 747 1542
rect 815 1546 819 1547
rect 815 1541 819 1542
rect 823 1546 827 1547
rect 823 1541 827 1542
rect 887 1546 891 1547
rect 887 1541 891 1542
rect 911 1546 915 1547
rect 911 1541 915 1542
rect 999 1546 1003 1547
rect 999 1541 1003 1542
rect 1095 1546 1099 1547
rect 1095 1541 1099 1542
rect 112 1538 114 1541
rect 134 1540 140 1541
rect 110 1537 116 1538
rect 110 1533 111 1537
rect 115 1533 116 1537
rect 134 1536 135 1540
rect 139 1536 140 1540
rect 134 1535 140 1536
rect 174 1540 180 1541
rect 174 1536 175 1540
rect 179 1536 180 1540
rect 174 1535 180 1536
rect 230 1540 236 1541
rect 230 1536 231 1540
rect 235 1536 236 1540
rect 230 1535 236 1536
rect 310 1540 316 1541
rect 310 1536 311 1540
rect 315 1536 316 1540
rect 310 1535 316 1536
rect 390 1540 396 1541
rect 390 1536 391 1540
rect 395 1536 396 1540
rect 390 1535 396 1536
rect 478 1540 484 1541
rect 478 1536 479 1540
rect 483 1536 484 1540
rect 478 1535 484 1536
rect 566 1540 572 1541
rect 566 1536 567 1540
rect 571 1536 572 1540
rect 566 1535 572 1536
rect 654 1540 660 1541
rect 654 1536 655 1540
rect 659 1536 660 1540
rect 654 1535 660 1536
rect 742 1540 748 1541
rect 742 1536 743 1540
rect 747 1536 748 1540
rect 742 1535 748 1536
rect 822 1540 828 1541
rect 822 1536 823 1540
rect 827 1536 828 1540
rect 822 1535 828 1536
rect 910 1540 916 1541
rect 910 1536 911 1540
rect 915 1536 916 1540
rect 910 1535 916 1536
rect 998 1540 1004 1541
rect 998 1536 999 1540
rect 1003 1536 1004 1540
rect 1096 1538 1098 1541
rect 998 1535 1004 1536
rect 1094 1537 1100 1538
rect 1136 1537 1138 1557
rect 1160 1545 1162 1557
rect 1200 1545 1202 1557
rect 1248 1545 1250 1557
rect 1320 1545 1322 1557
rect 1400 1545 1402 1557
rect 1480 1545 1482 1557
rect 1560 1545 1562 1557
rect 1648 1545 1650 1557
rect 1736 1545 1738 1557
rect 1824 1545 1826 1557
rect 1912 1545 1914 1557
rect 2000 1545 2002 1557
rect 2072 1545 2074 1557
rect 1158 1544 1164 1545
rect 1158 1540 1159 1544
rect 1163 1540 1164 1544
rect 1158 1539 1164 1540
rect 1198 1544 1204 1545
rect 1198 1540 1199 1544
rect 1203 1540 1204 1544
rect 1198 1539 1204 1540
rect 1246 1544 1252 1545
rect 1246 1540 1247 1544
rect 1251 1540 1252 1544
rect 1246 1539 1252 1540
rect 1318 1544 1324 1545
rect 1318 1540 1319 1544
rect 1323 1540 1324 1544
rect 1318 1539 1324 1540
rect 1398 1544 1404 1545
rect 1398 1540 1399 1544
rect 1403 1540 1404 1544
rect 1398 1539 1404 1540
rect 1478 1544 1484 1545
rect 1478 1540 1479 1544
rect 1483 1540 1484 1544
rect 1478 1539 1484 1540
rect 1558 1544 1564 1545
rect 1558 1540 1559 1544
rect 1563 1540 1564 1544
rect 1558 1539 1564 1540
rect 1646 1544 1652 1545
rect 1646 1540 1647 1544
rect 1651 1540 1652 1544
rect 1646 1539 1652 1540
rect 1734 1544 1740 1545
rect 1734 1540 1735 1544
rect 1739 1540 1740 1544
rect 1734 1539 1740 1540
rect 1822 1544 1828 1545
rect 1822 1540 1823 1544
rect 1827 1540 1828 1544
rect 1822 1539 1828 1540
rect 1910 1544 1916 1545
rect 1910 1540 1911 1544
rect 1915 1540 1916 1544
rect 1910 1539 1916 1540
rect 1998 1544 2004 1545
rect 1998 1540 1999 1544
rect 2003 1540 2004 1544
rect 1998 1539 2004 1540
rect 2070 1544 2076 1545
rect 2070 1540 2071 1544
rect 2075 1540 2076 1544
rect 2070 1539 2076 1540
rect 2120 1537 2122 1557
rect 110 1532 116 1533
rect 1094 1533 1095 1537
rect 1099 1533 1100 1537
rect 1094 1532 1100 1533
rect 1134 1536 1140 1537
rect 1134 1532 1135 1536
rect 1139 1532 1140 1536
rect 1134 1531 1140 1532
rect 2118 1536 2124 1537
rect 2118 1532 2119 1536
rect 2123 1532 2124 1536
rect 2118 1531 2124 1532
rect 110 1520 116 1521
rect 110 1516 111 1520
rect 115 1516 116 1520
rect 110 1515 116 1516
rect 1094 1520 1100 1521
rect 1094 1516 1095 1520
rect 1099 1516 1100 1520
rect 1094 1515 1100 1516
rect 1134 1519 1140 1520
rect 1134 1515 1135 1519
rect 1139 1515 1140 1519
rect 2118 1519 2124 1520
rect 112 1495 114 1515
rect 134 1512 140 1513
rect 134 1508 135 1512
rect 139 1508 140 1512
rect 134 1507 140 1508
rect 174 1512 180 1513
rect 174 1508 175 1512
rect 179 1508 180 1512
rect 174 1507 180 1508
rect 230 1512 236 1513
rect 230 1508 231 1512
rect 235 1508 236 1512
rect 230 1507 236 1508
rect 310 1512 316 1513
rect 310 1508 311 1512
rect 315 1508 316 1512
rect 310 1507 316 1508
rect 390 1512 396 1513
rect 390 1508 391 1512
rect 395 1508 396 1512
rect 390 1507 396 1508
rect 478 1512 484 1513
rect 478 1508 479 1512
rect 483 1508 484 1512
rect 478 1507 484 1508
rect 566 1512 572 1513
rect 566 1508 567 1512
rect 571 1508 572 1512
rect 566 1507 572 1508
rect 654 1512 660 1513
rect 654 1508 655 1512
rect 659 1508 660 1512
rect 654 1507 660 1508
rect 742 1512 748 1513
rect 742 1508 743 1512
rect 747 1508 748 1512
rect 742 1507 748 1508
rect 822 1512 828 1513
rect 822 1508 823 1512
rect 827 1508 828 1512
rect 822 1507 828 1508
rect 910 1512 916 1513
rect 910 1508 911 1512
rect 915 1508 916 1512
rect 910 1507 916 1508
rect 998 1512 1004 1513
rect 998 1508 999 1512
rect 1003 1508 1004 1512
rect 998 1507 1004 1508
rect 136 1495 138 1507
rect 176 1495 178 1507
rect 232 1495 234 1507
rect 312 1495 314 1507
rect 392 1495 394 1507
rect 480 1495 482 1507
rect 568 1495 570 1507
rect 656 1495 658 1507
rect 744 1495 746 1507
rect 824 1495 826 1507
rect 912 1495 914 1507
rect 1000 1495 1002 1507
rect 1096 1495 1098 1515
rect 1134 1514 1140 1515
rect 1158 1516 1164 1517
rect 1136 1511 1138 1514
rect 1158 1512 1159 1516
rect 1163 1512 1164 1516
rect 1158 1511 1164 1512
rect 1198 1516 1204 1517
rect 1198 1512 1199 1516
rect 1203 1512 1204 1516
rect 1198 1511 1204 1512
rect 1246 1516 1252 1517
rect 1246 1512 1247 1516
rect 1251 1512 1252 1516
rect 1246 1511 1252 1512
rect 1318 1516 1324 1517
rect 1318 1512 1319 1516
rect 1323 1512 1324 1516
rect 1318 1511 1324 1512
rect 1398 1516 1404 1517
rect 1398 1512 1399 1516
rect 1403 1512 1404 1516
rect 1398 1511 1404 1512
rect 1478 1516 1484 1517
rect 1478 1512 1479 1516
rect 1483 1512 1484 1516
rect 1478 1511 1484 1512
rect 1558 1516 1564 1517
rect 1558 1512 1559 1516
rect 1563 1512 1564 1516
rect 1558 1511 1564 1512
rect 1646 1516 1652 1517
rect 1646 1512 1647 1516
rect 1651 1512 1652 1516
rect 1646 1511 1652 1512
rect 1734 1516 1740 1517
rect 1734 1512 1735 1516
rect 1739 1512 1740 1516
rect 1734 1511 1740 1512
rect 1822 1516 1828 1517
rect 1822 1512 1823 1516
rect 1827 1512 1828 1516
rect 1822 1511 1828 1512
rect 1910 1516 1916 1517
rect 1910 1512 1911 1516
rect 1915 1512 1916 1516
rect 1910 1511 1916 1512
rect 1998 1516 2004 1517
rect 1998 1512 1999 1516
rect 2003 1512 2004 1516
rect 1998 1511 2004 1512
rect 2070 1516 2076 1517
rect 2070 1512 2071 1516
rect 2075 1512 2076 1516
rect 2118 1515 2119 1519
rect 2123 1515 2124 1519
rect 2118 1514 2124 1515
rect 2070 1511 2076 1512
rect 2120 1511 2122 1514
rect 1135 1510 1139 1511
rect 1135 1505 1139 1506
rect 1159 1510 1163 1511
rect 1159 1505 1163 1506
rect 1199 1510 1203 1511
rect 1199 1505 1203 1506
rect 1239 1510 1243 1511
rect 1239 1505 1243 1506
rect 1247 1510 1251 1511
rect 1247 1505 1251 1506
rect 1303 1510 1307 1511
rect 1303 1505 1307 1506
rect 1319 1510 1323 1511
rect 1319 1505 1323 1506
rect 1375 1510 1379 1511
rect 1375 1505 1379 1506
rect 1399 1510 1403 1511
rect 1399 1505 1403 1506
rect 1455 1510 1459 1511
rect 1455 1505 1459 1506
rect 1479 1510 1483 1511
rect 1479 1505 1483 1506
rect 1543 1510 1547 1511
rect 1543 1505 1547 1506
rect 1559 1510 1563 1511
rect 1559 1505 1563 1506
rect 1623 1510 1627 1511
rect 1623 1505 1627 1506
rect 1647 1510 1651 1511
rect 1647 1505 1651 1506
rect 1703 1510 1707 1511
rect 1703 1505 1707 1506
rect 1735 1510 1739 1511
rect 1735 1505 1739 1506
rect 1775 1510 1779 1511
rect 1775 1505 1779 1506
rect 1823 1510 1827 1511
rect 1823 1505 1827 1506
rect 1847 1510 1851 1511
rect 1847 1505 1851 1506
rect 1911 1510 1915 1511
rect 1911 1505 1915 1506
rect 1919 1510 1923 1511
rect 1919 1505 1923 1506
rect 1991 1510 1995 1511
rect 1991 1505 1995 1506
rect 1999 1510 2003 1511
rect 1999 1505 2003 1506
rect 2063 1510 2067 1511
rect 2063 1505 2067 1506
rect 2071 1510 2075 1511
rect 2071 1505 2075 1506
rect 2119 1510 2123 1511
rect 2119 1505 2123 1506
rect 1136 1502 1138 1505
rect 1158 1504 1164 1505
rect 1134 1501 1140 1502
rect 1134 1497 1135 1501
rect 1139 1497 1140 1501
rect 1158 1500 1159 1504
rect 1163 1500 1164 1504
rect 1158 1499 1164 1500
rect 1198 1504 1204 1505
rect 1198 1500 1199 1504
rect 1203 1500 1204 1504
rect 1198 1499 1204 1500
rect 1238 1504 1244 1505
rect 1238 1500 1239 1504
rect 1243 1500 1244 1504
rect 1238 1499 1244 1500
rect 1302 1504 1308 1505
rect 1302 1500 1303 1504
rect 1307 1500 1308 1504
rect 1302 1499 1308 1500
rect 1374 1504 1380 1505
rect 1374 1500 1375 1504
rect 1379 1500 1380 1504
rect 1374 1499 1380 1500
rect 1454 1504 1460 1505
rect 1454 1500 1455 1504
rect 1459 1500 1460 1504
rect 1454 1499 1460 1500
rect 1542 1504 1548 1505
rect 1542 1500 1543 1504
rect 1547 1500 1548 1504
rect 1542 1499 1548 1500
rect 1622 1504 1628 1505
rect 1622 1500 1623 1504
rect 1627 1500 1628 1504
rect 1622 1499 1628 1500
rect 1702 1504 1708 1505
rect 1702 1500 1703 1504
rect 1707 1500 1708 1504
rect 1702 1499 1708 1500
rect 1774 1504 1780 1505
rect 1774 1500 1775 1504
rect 1779 1500 1780 1504
rect 1774 1499 1780 1500
rect 1846 1504 1852 1505
rect 1846 1500 1847 1504
rect 1851 1500 1852 1504
rect 1846 1499 1852 1500
rect 1918 1504 1924 1505
rect 1918 1500 1919 1504
rect 1923 1500 1924 1504
rect 1918 1499 1924 1500
rect 1990 1504 1996 1505
rect 1990 1500 1991 1504
rect 1995 1500 1996 1504
rect 1990 1499 1996 1500
rect 2062 1504 2068 1505
rect 2062 1500 2063 1504
rect 2067 1500 2068 1504
rect 2120 1502 2122 1505
rect 2062 1499 2068 1500
rect 2118 1501 2124 1502
rect 1134 1496 1140 1497
rect 2118 1497 2119 1501
rect 2123 1497 2124 1501
rect 2118 1496 2124 1497
rect 111 1494 115 1495
rect 111 1489 115 1490
rect 135 1494 139 1495
rect 135 1489 139 1490
rect 175 1494 179 1495
rect 175 1489 179 1490
rect 199 1494 203 1495
rect 199 1489 203 1490
rect 231 1494 235 1495
rect 231 1489 235 1490
rect 279 1494 283 1495
rect 279 1489 283 1490
rect 311 1494 315 1495
rect 311 1489 315 1490
rect 359 1494 363 1495
rect 359 1489 363 1490
rect 391 1494 395 1495
rect 391 1489 395 1490
rect 439 1494 443 1495
rect 439 1489 443 1490
rect 479 1494 483 1495
rect 479 1489 483 1490
rect 519 1494 523 1495
rect 519 1489 523 1490
rect 567 1494 571 1495
rect 567 1489 571 1490
rect 599 1494 603 1495
rect 599 1489 603 1490
rect 655 1494 659 1495
rect 655 1489 659 1490
rect 679 1494 683 1495
rect 679 1489 683 1490
rect 743 1494 747 1495
rect 743 1489 747 1490
rect 767 1494 771 1495
rect 767 1489 771 1490
rect 823 1494 827 1495
rect 823 1489 827 1490
rect 855 1494 859 1495
rect 855 1489 859 1490
rect 911 1494 915 1495
rect 911 1489 915 1490
rect 943 1494 947 1495
rect 943 1489 947 1490
rect 999 1494 1003 1495
rect 999 1489 1003 1490
rect 1031 1494 1035 1495
rect 1031 1489 1035 1490
rect 1095 1494 1099 1495
rect 1095 1489 1099 1490
rect 112 1469 114 1489
rect 136 1477 138 1489
rect 200 1477 202 1489
rect 280 1477 282 1489
rect 360 1477 362 1489
rect 440 1477 442 1489
rect 520 1477 522 1489
rect 600 1477 602 1489
rect 680 1477 682 1489
rect 768 1477 770 1489
rect 856 1477 858 1489
rect 944 1477 946 1489
rect 1032 1477 1034 1489
rect 134 1476 140 1477
rect 134 1472 135 1476
rect 139 1472 140 1476
rect 134 1471 140 1472
rect 198 1476 204 1477
rect 198 1472 199 1476
rect 203 1472 204 1476
rect 198 1471 204 1472
rect 278 1476 284 1477
rect 278 1472 279 1476
rect 283 1472 284 1476
rect 278 1471 284 1472
rect 358 1476 364 1477
rect 358 1472 359 1476
rect 363 1472 364 1476
rect 358 1471 364 1472
rect 438 1476 444 1477
rect 438 1472 439 1476
rect 443 1472 444 1476
rect 438 1471 444 1472
rect 518 1476 524 1477
rect 518 1472 519 1476
rect 523 1472 524 1476
rect 518 1471 524 1472
rect 598 1476 604 1477
rect 598 1472 599 1476
rect 603 1472 604 1476
rect 598 1471 604 1472
rect 678 1476 684 1477
rect 678 1472 679 1476
rect 683 1472 684 1476
rect 678 1471 684 1472
rect 766 1476 772 1477
rect 766 1472 767 1476
rect 771 1472 772 1476
rect 766 1471 772 1472
rect 854 1476 860 1477
rect 854 1472 855 1476
rect 859 1472 860 1476
rect 854 1471 860 1472
rect 942 1476 948 1477
rect 942 1472 943 1476
rect 947 1472 948 1476
rect 942 1471 948 1472
rect 1030 1476 1036 1477
rect 1030 1472 1031 1476
rect 1035 1472 1036 1476
rect 1030 1471 1036 1472
rect 1096 1469 1098 1489
rect 1134 1484 1140 1485
rect 1134 1480 1135 1484
rect 1139 1480 1140 1484
rect 1134 1479 1140 1480
rect 2118 1484 2124 1485
rect 2118 1480 2119 1484
rect 2123 1480 2124 1484
rect 2118 1479 2124 1480
rect 110 1468 116 1469
rect 110 1464 111 1468
rect 115 1464 116 1468
rect 110 1463 116 1464
rect 1094 1468 1100 1469
rect 1094 1464 1095 1468
rect 1099 1464 1100 1468
rect 1094 1463 1100 1464
rect 1136 1455 1138 1479
rect 1158 1476 1164 1477
rect 1158 1472 1159 1476
rect 1163 1472 1164 1476
rect 1158 1471 1164 1472
rect 1198 1476 1204 1477
rect 1198 1472 1199 1476
rect 1203 1472 1204 1476
rect 1198 1471 1204 1472
rect 1238 1476 1244 1477
rect 1238 1472 1239 1476
rect 1243 1472 1244 1476
rect 1238 1471 1244 1472
rect 1302 1476 1308 1477
rect 1302 1472 1303 1476
rect 1307 1472 1308 1476
rect 1302 1471 1308 1472
rect 1374 1476 1380 1477
rect 1374 1472 1375 1476
rect 1379 1472 1380 1476
rect 1374 1471 1380 1472
rect 1454 1476 1460 1477
rect 1454 1472 1455 1476
rect 1459 1472 1460 1476
rect 1454 1471 1460 1472
rect 1542 1476 1548 1477
rect 1542 1472 1543 1476
rect 1547 1472 1548 1476
rect 1542 1471 1548 1472
rect 1622 1476 1628 1477
rect 1622 1472 1623 1476
rect 1627 1472 1628 1476
rect 1622 1471 1628 1472
rect 1702 1476 1708 1477
rect 1702 1472 1703 1476
rect 1707 1472 1708 1476
rect 1702 1471 1708 1472
rect 1774 1476 1780 1477
rect 1774 1472 1775 1476
rect 1779 1472 1780 1476
rect 1774 1471 1780 1472
rect 1846 1476 1852 1477
rect 1846 1472 1847 1476
rect 1851 1472 1852 1476
rect 1846 1471 1852 1472
rect 1918 1476 1924 1477
rect 1918 1472 1919 1476
rect 1923 1472 1924 1476
rect 1918 1471 1924 1472
rect 1990 1476 1996 1477
rect 1990 1472 1991 1476
rect 1995 1472 1996 1476
rect 1990 1471 1996 1472
rect 2062 1476 2068 1477
rect 2062 1472 2063 1476
rect 2067 1472 2068 1476
rect 2062 1471 2068 1472
rect 1160 1455 1162 1471
rect 1200 1455 1202 1471
rect 1240 1455 1242 1471
rect 1304 1455 1306 1471
rect 1376 1455 1378 1471
rect 1456 1455 1458 1471
rect 1544 1455 1546 1471
rect 1624 1455 1626 1471
rect 1704 1455 1706 1471
rect 1776 1455 1778 1471
rect 1848 1455 1850 1471
rect 1920 1455 1922 1471
rect 1992 1455 1994 1471
rect 2064 1455 2066 1471
rect 2120 1455 2122 1479
rect 1135 1454 1139 1455
rect 110 1451 116 1452
rect 110 1447 111 1451
rect 115 1447 116 1451
rect 1094 1451 1100 1452
rect 110 1446 116 1447
rect 134 1448 140 1449
rect 112 1443 114 1446
rect 134 1444 135 1448
rect 139 1444 140 1448
rect 134 1443 140 1444
rect 198 1448 204 1449
rect 198 1444 199 1448
rect 203 1444 204 1448
rect 198 1443 204 1444
rect 278 1448 284 1449
rect 278 1444 279 1448
rect 283 1444 284 1448
rect 278 1443 284 1444
rect 358 1448 364 1449
rect 358 1444 359 1448
rect 363 1444 364 1448
rect 358 1443 364 1444
rect 438 1448 444 1449
rect 438 1444 439 1448
rect 443 1444 444 1448
rect 438 1443 444 1444
rect 518 1448 524 1449
rect 518 1444 519 1448
rect 523 1444 524 1448
rect 518 1443 524 1444
rect 598 1448 604 1449
rect 598 1444 599 1448
rect 603 1444 604 1448
rect 598 1443 604 1444
rect 678 1448 684 1449
rect 678 1444 679 1448
rect 683 1444 684 1448
rect 678 1443 684 1444
rect 766 1448 772 1449
rect 766 1444 767 1448
rect 771 1444 772 1448
rect 766 1443 772 1444
rect 854 1448 860 1449
rect 854 1444 855 1448
rect 859 1444 860 1448
rect 854 1443 860 1444
rect 942 1448 948 1449
rect 942 1444 943 1448
rect 947 1444 948 1448
rect 942 1443 948 1444
rect 1030 1448 1036 1449
rect 1030 1444 1031 1448
rect 1035 1444 1036 1448
rect 1094 1447 1095 1451
rect 1099 1447 1100 1451
rect 1135 1449 1139 1450
rect 1159 1454 1163 1455
rect 1159 1449 1163 1450
rect 1199 1454 1203 1455
rect 1199 1449 1203 1450
rect 1239 1454 1243 1455
rect 1239 1449 1243 1450
rect 1279 1454 1283 1455
rect 1279 1449 1283 1450
rect 1303 1454 1307 1455
rect 1303 1449 1307 1450
rect 1327 1454 1331 1455
rect 1327 1449 1331 1450
rect 1375 1454 1379 1455
rect 1375 1449 1379 1450
rect 1383 1454 1387 1455
rect 1383 1449 1387 1450
rect 1439 1454 1443 1455
rect 1439 1449 1443 1450
rect 1455 1454 1459 1455
rect 1455 1449 1459 1450
rect 1495 1454 1499 1455
rect 1495 1449 1499 1450
rect 1543 1454 1547 1455
rect 1543 1449 1547 1450
rect 1551 1454 1555 1455
rect 1551 1449 1555 1450
rect 1607 1454 1611 1455
rect 1607 1449 1611 1450
rect 1623 1454 1627 1455
rect 1623 1449 1627 1450
rect 1671 1454 1675 1455
rect 1671 1449 1675 1450
rect 1703 1454 1707 1455
rect 1703 1449 1707 1450
rect 1735 1454 1739 1455
rect 1735 1449 1739 1450
rect 1775 1454 1779 1455
rect 1775 1449 1779 1450
rect 1807 1454 1811 1455
rect 1807 1449 1811 1450
rect 1847 1454 1851 1455
rect 1847 1449 1851 1450
rect 1887 1454 1891 1455
rect 1887 1449 1891 1450
rect 1919 1454 1923 1455
rect 1919 1449 1923 1450
rect 1975 1454 1979 1455
rect 1975 1449 1979 1450
rect 1991 1454 1995 1455
rect 1991 1449 1995 1450
rect 2063 1454 2067 1455
rect 2063 1449 2067 1450
rect 2119 1454 2123 1455
rect 2119 1449 2123 1450
rect 1094 1446 1100 1447
rect 1030 1443 1036 1444
rect 1096 1443 1098 1446
rect 111 1442 115 1443
rect 111 1437 115 1438
rect 135 1442 139 1443
rect 135 1437 139 1438
rect 191 1442 195 1443
rect 191 1437 195 1438
rect 199 1442 203 1443
rect 199 1437 203 1438
rect 263 1442 267 1443
rect 263 1437 267 1438
rect 279 1442 283 1443
rect 279 1437 283 1438
rect 335 1442 339 1443
rect 335 1437 339 1438
rect 359 1442 363 1443
rect 359 1437 363 1438
rect 407 1442 411 1443
rect 407 1437 411 1438
rect 439 1442 443 1443
rect 439 1437 443 1438
rect 479 1442 483 1443
rect 479 1437 483 1438
rect 519 1442 523 1443
rect 519 1437 523 1438
rect 551 1442 555 1443
rect 551 1437 555 1438
rect 599 1442 603 1443
rect 599 1437 603 1438
rect 631 1442 635 1443
rect 631 1437 635 1438
rect 679 1442 683 1443
rect 679 1437 683 1438
rect 711 1442 715 1443
rect 711 1437 715 1438
rect 767 1442 771 1443
rect 767 1437 771 1438
rect 799 1442 803 1443
rect 799 1437 803 1438
rect 855 1442 859 1443
rect 855 1437 859 1438
rect 887 1442 891 1443
rect 887 1437 891 1438
rect 943 1442 947 1443
rect 943 1437 947 1438
rect 975 1442 979 1443
rect 975 1437 979 1438
rect 1031 1442 1035 1443
rect 1031 1437 1035 1438
rect 1047 1442 1051 1443
rect 1047 1437 1051 1438
rect 1095 1442 1099 1443
rect 1095 1437 1099 1438
rect 112 1434 114 1437
rect 134 1436 140 1437
rect 110 1433 116 1434
rect 110 1429 111 1433
rect 115 1429 116 1433
rect 134 1432 135 1436
rect 139 1432 140 1436
rect 134 1431 140 1432
rect 190 1436 196 1437
rect 190 1432 191 1436
rect 195 1432 196 1436
rect 190 1431 196 1432
rect 262 1436 268 1437
rect 262 1432 263 1436
rect 267 1432 268 1436
rect 262 1431 268 1432
rect 334 1436 340 1437
rect 334 1432 335 1436
rect 339 1432 340 1436
rect 334 1431 340 1432
rect 406 1436 412 1437
rect 406 1432 407 1436
rect 411 1432 412 1436
rect 406 1431 412 1432
rect 478 1436 484 1437
rect 478 1432 479 1436
rect 483 1432 484 1436
rect 478 1431 484 1432
rect 550 1436 556 1437
rect 550 1432 551 1436
rect 555 1432 556 1436
rect 550 1431 556 1432
rect 630 1436 636 1437
rect 630 1432 631 1436
rect 635 1432 636 1436
rect 630 1431 636 1432
rect 710 1436 716 1437
rect 710 1432 711 1436
rect 715 1432 716 1436
rect 710 1431 716 1432
rect 798 1436 804 1437
rect 798 1432 799 1436
rect 803 1432 804 1436
rect 798 1431 804 1432
rect 886 1436 892 1437
rect 886 1432 887 1436
rect 891 1432 892 1436
rect 886 1431 892 1432
rect 974 1436 980 1437
rect 974 1432 975 1436
rect 979 1432 980 1436
rect 974 1431 980 1432
rect 1046 1436 1052 1437
rect 1046 1432 1047 1436
rect 1051 1432 1052 1436
rect 1096 1434 1098 1437
rect 1046 1431 1052 1432
rect 1094 1433 1100 1434
rect 110 1428 116 1429
rect 1094 1429 1095 1433
rect 1099 1429 1100 1433
rect 1136 1429 1138 1449
rect 1280 1437 1282 1449
rect 1328 1437 1330 1449
rect 1384 1437 1386 1449
rect 1440 1437 1442 1449
rect 1496 1437 1498 1449
rect 1552 1437 1554 1449
rect 1608 1437 1610 1449
rect 1672 1437 1674 1449
rect 1736 1437 1738 1449
rect 1808 1437 1810 1449
rect 1888 1437 1890 1449
rect 1976 1437 1978 1449
rect 2064 1437 2066 1449
rect 1278 1436 1284 1437
rect 1278 1432 1279 1436
rect 1283 1432 1284 1436
rect 1278 1431 1284 1432
rect 1326 1436 1332 1437
rect 1326 1432 1327 1436
rect 1331 1432 1332 1436
rect 1326 1431 1332 1432
rect 1382 1436 1388 1437
rect 1382 1432 1383 1436
rect 1387 1432 1388 1436
rect 1382 1431 1388 1432
rect 1438 1436 1444 1437
rect 1438 1432 1439 1436
rect 1443 1432 1444 1436
rect 1438 1431 1444 1432
rect 1494 1436 1500 1437
rect 1494 1432 1495 1436
rect 1499 1432 1500 1436
rect 1494 1431 1500 1432
rect 1550 1436 1556 1437
rect 1550 1432 1551 1436
rect 1555 1432 1556 1436
rect 1550 1431 1556 1432
rect 1606 1436 1612 1437
rect 1606 1432 1607 1436
rect 1611 1432 1612 1436
rect 1606 1431 1612 1432
rect 1670 1436 1676 1437
rect 1670 1432 1671 1436
rect 1675 1432 1676 1436
rect 1670 1431 1676 1432
rect 1734 1436 1740 1437
rect 1734 1432 1735 1436
rect 1739 1432 1740 1436
rect 1734 1431 1740 1432
rect 1806 1436 1812 1437
rect 1806 1432 1807 1436
rect 1811 1432 1812 1436
rect 1806 1431 1812 1432
rect 1886 1436 1892 1437
rect 1886 1432 1887 1436
rect 1891 1432 1892 1436
rect 1886 1431 1892 1432
rect 1974 1436 1980 1437
rect 1974 1432 1975 1436
rect 1979 1432 1980 1436
rect 1974 1431 1980 1432
rect 2062 1436 2068 1437
rect 2062 1432 2063 1436
rect 2067 1432 2068 1436
rect 2062 1431 2068 1432
rect 2120 1429 2122 1449
rect 1094 1428 1100 1429
rect 1134 1428 1140 1429
rect 1134 1424 1135 1428
rect 1139 1424 1140 1428
rect 1134 1423 1140 1424
rect 2118 1428 2124 1429
rect 2118 1424 2119 1428
rect 2123 1424 2124 1428
rect 2118 1423 2124 1424
rect 110 1416 116 1417
rect 110 1412 111 1416
rect 115 1412 116 1416
rect 110 1411 116 1412
rect 1094 1416 1100 1417
rect 1094 1412 1095 1416
rect 1099 1412 1100 1416
rect 1094 1411 1100 1412
rect 1134 1411 1140 1412
rect 112 1391 114 1411
rect 134 1408 140 1409
rect 134 1404 135 1408
rect 139 1404 140 1408
rect 134 1403 140 1404
rect 190 1408 196 1409
rect 190 1404 191 1408
rect 195 1404 196 1408
rect 190 1403 196 1404
rect 262 1408 268 1409
rect 262 1404 263 1408
rect 267 1404 268 1408
rect 262 1403 268 1404
rect 334 1408 340 1409
rect 334 1404 335 1408
rect 339 1404 340 1408
rect 334 1403 340 1404
rect 406 1408 412 1409
rect 406 1404 407 1408
rect 411 1404 412 1408
rect 406 1403 412 1404
rect 478 1408 484 1409
rect 478 1404 479 1408
rect 483 1404 484 1408
rect 478 1403 484 1404
rect 550 1408 556 1409
rect 550 1404 551 1408
rect 555 1404 556 1408
rect 550 1403 556 1404
rect 630 1408 636 1409
rect 630 1404 631 1408
rect 635 1404 636 1408
rect 630 1403 636 1404
rect 710 1408 716 1409
rect 710 1404 711 1408
rect 715 1404 716 1408
rect 710 1403 716 1404
rect 798 1408 804 1409
rect 798 1404 799 1408
rect 803 1404 804 1408
rect 798 1403 804 1404
rect 886 1408 892 1409
rect 886 1404 887 1408
rect 891 1404 892 1408
rect 886 1403 892 1404
rect 974 1408 980 1409
rect 974 1404 975 1408
rect 979 1404 980 1408
rect 974 1403 980 1404
rect 1046 1408 1052 1409
rect 1046 1404 1047 1408
rect 1051 1404 1052 1408
rect 1046 1403 1052 1404
rect 136 1391 138 1403
rect 192 1391 194 1403
rect 264 1391 266 1403
rect 336 1391 338 1403
rect 408 1391 410 1403
rect 480 1391 482 1403
rect 552 1391 554 1403
rect 632 1391 634 1403
rect 712 1391 714 1403
rect 800 1391 802 1403
rect 888 1391 890 1403
rect 976 1391 978 1403
rect 1048 1391 1050 1403
rect 1096 1391 1098 1411
rect 1134 1407 1135 1411
rect 1139 1407 1140 1411
rect 2118 1411 2124 1412
rect 1134 1406 1140 1407
rect 1278 1408 1284 1409
rect 1136 1399 1138 1406
rect 1278 1404 1279 1408
rect 1283 1404 1284 1408
rect 1278 1403 1284 1404
rect 1326 1408 1332 1409
rect 1326 1404 1327 1408
rect 1331 1404 1332 1408
rect 1326 1403 1332 1404
rect 1382 1408 1388 1409
rect 1382 1404 1383 1408
rect 1387 1404 1388 1408
rect 1382 1403 1388 1404
rect 1438 1408 1444 1409
rect 1438 1404 1439 1408
rect 1443 1404 1444 1408
rect 1438 1403 1444 1404
rect 1494 1408 1500 1409
rect 1494 1404 1495 1408
rect 1499 1404 1500 1408
rect 1494 1403 1500 1404
rect 1550 1408 1556 1409
rect 1550 1404 1551 1408
rect 1555 1404 1556 1408
rect 1550 1403 1556 1404
rect 1606 1408 1612 1409
rect 1606 1404 1607 1408
rect 1611 1404 1612 1408
rect 1606 1403 1612 1404
rect 1670 1408 1676 1409
rect 1670 1404 1671 1408
rect 1675 1404 1676 1408
rect 1670 1403 1676 1404
rect 1734 1408 1740 1409
rect 1734 1404 1735 1408
rect 1739 1404 1740 1408
rect 1734 1403 1740 1404
rect 1806 1408 1812 1409
rect 1806 1404 1807 1408
rect 1811 1404 1812 1408
rect 1806 1403 1812 1404
rect 1886 1408 1892 1409
rect 1886 1404 1887 1408
rect 1891 1404 1892 1408
rect 1886 1403 1892 1404
rect 1974 1408 1980 1409
rect 1974 1404 1975 1408
rect 1979 1404 1980 1408
rect 1974 1403 1980 1404
rect 2062 1408 2068 1409
rect 2062 1404 2063 1408
rect 2067 1404 2068 1408
rect 2118 1407 2119 1411
rect 2123 1407 2124 1411
rect 2118 1406 2124 1407
rect 2062 1403 2068 1404
rect 1280 1399 1282 1403
rect 1328 1399 1330 1403
rect 1384 1399 1386 1403
rect 1440 1399 1442 1403
rect 1496 1399 1498 1403
rect 1552 1399 1554 1403
rect 1608 1399 1610 1403
rect 1672 1399 1674 1403
rect 1736 1399 1738 1403
rect 1808 1399 1810 1403
rect 1888 1399 1890 1403
rect 1976 1399 1978 1403
rect 2064 1399 2066 1403
rect 2120 1399 2122 1406
rect 1135 1398 1139 1399
rect 1135 1393 1139 1394
rect 1279 1398 1283 1399
rect 1279 1393 1283 1394
rect 1327 1398 1331 1399
rect 1327 1393 1331 1394
rect 1335 1398 1339 1399
rect 1335 1393 1339 1394
rect 1375 1398 1379 1399
rect 1375 1393 1379 1394
rect 1383 1398 1387 1399
rect 1383 1393 1387 1394
rect 1415 1398 1419 1399
rect 1415 1393 1419 1394
rect 1439 1398 1443 1399
rect 1439 1393 1443 1394
rect 1455 1398 1459 1399
rect 1455 1393 1459 1394
rect 1495 1398 1499 1399
rect 1495 1393 1499 1394
rect 1535 1398 1539 1399
rect 1535 1393 1539 1394
rect 1551 1398 1555 1399
rect 1551 1393 1555 1394
rect 1583 1398 1587 1399
rect 1583 1393 1587 1394
rect 1607 1398 1611 1399
rect 1607 1393 1611 1394
rect 1647 1398 1651 1399
rect 1647 1393 1651 1394
rect 1671 1398 1675 1399
rect 1671 1393 1675 1394
rect 1719 1398 1723 1399
rect 1719 1393 1723 1394
rect 1735 1398 1739 1399
rect 1735 1393 1739 1394
rect 1807 1398 1811 1399
rect 1807 1393 1811 1394
rect 1887 1398 1891 1399
rect 1887 1393 1891 1394
rect 1895 1398 1899 1399
rect 1895 1393 1899 1394
rect 1975 1398 1979 1399
rect 1975 1393 1979 1394
rect 1991 1398 1995 1399
rect 1991 1393 1995 1394
rect 2063 1398 2067 1399
rect 2063 1393 2067 1394
rect 2071 1398 2075 1399
rect 2071 1393 2075 1394
rect 2119 1398 2123 1399
rect 2119 1393 2123 1394
rect 111 1390 115 1391
rect 111 1385 115 1386
rect 135 1390 139 1391
rect 135 1385 139 1386
rect 175 1390 179 1391
rect 175 1385 179 1386
rect 191 1390 195 1391
rect 191 1385 195 1386
rect 239 1390 243 1391
rect 239 1385 243 1386
rect 263 1390 267 1391
rect 263 1385 267 1386
rect 303 1390 307 1391
rect 303 1385 307 1386
rect 335 1390 339 1391
rect 335 1385 339 1386
rect 367 1390 371 1391
rect 367 1385 371 1386
rect 407 1390 411 1391
rect 407 1385 411 1386
rect 439 1390 443 1391
rect 439 1385 443 1386
rect 479 1390 483 1391
rect 479 1385 483 1386
rect 503 1390 507 1391
rect 503 1385 507 1386
rect 551 1390 555 1391
rect 551 1385 555 1386
rect 575 1390 579 1391
rect 575 1385 579 1386
rect 631 1390 635 1391
rect 631 1385 635 1386
rect 647 1390 651 1391
rect 647 1385 651 1386
rect 711 1390 715 1391
rect 711 1385 715 1386
rect 783 1390 787 1391
rect 783 1385 787 1386
rect 799 1390 803 1391
rect 799 1385 803 1386
rect 855 1390 859 1391
rect 855 1385 859 1386
rect 887 1390 891 1391
rect 887 1385 891 1386
rect 927 1390 931 1391
rect 927 1385 931 1386
rect 975 1390 979 1391
rect 975 1385 979 1386
rect 999 1390 1003 1391
rect 999 1385 1003 1386
rect 1047 1390 1051 1391
rect 1047 1385 1051 1386
rect 1095 1390 1099 1391
rect 1136 1390 1138 1393
rect 1334 1392 1340 1393
rect 1095 1385 1099 1386
rect 1134 1389 1140 1390
rect 1134 1385 1135 1389
rect 1139 1385 1140 1389
rect 1334 1388 1335 1392
rect 1339 1388 1340 1392
rect 1334 1387 1340 1388
rect 1374 1392 1380 1393
rect 1374 1388 1375 1392
rect 1379 1388 1380 1392
rect 1374 1387 1380 1388
rect 1414 1392 1420 1393
rect 1414 1388 1415 1392
rect 1419 1388 1420 1392
rect 1414 1387 1420 1388
rect 1454 1392 1460 1393
rect 1454 1388 1455 1392
rect 1459 1388 1460 1392
rect 1454 1387 1460 1388
rect 1494 1392 1500 1393
rect 1494 1388 1495 1392
rect 1499 1388 1500 1392
rect 1494 1387 1500 1388
rect 1534 1392 1540 1393
rect 1534 1388 1535 1392
rect 1539 1388 1540 1392
rect 1534 1387 1540 1388
rect 1582 1392 1588 1393
rect 1582 1388 1583 1392
rect 1587 1388 1588 1392
rect 1582 1387 1588 1388
rect 1646 1392 1652 1393
rect 1646 1388 1647 1392
rect 1651 1388 1652 1392
rect 1646 1387 1652 1388
rect 1718 1392 1724 1393
rect 1718 1388 1719 1392
rect 1723 1388 1724 1392
rect 1718 1387 1724 1388
rect 1806 1392 1812 1393
rect 1806 1388 1807 1392
rect 1811 1388 1812 1392
rect 1806 1387 1812 1388
rect 1894 1392 1900 1393
rect 1894 1388 1895 1392
rect 1899 1388 1900 1392
rect 1894 1387 1900 1388
rect 1990 1392 1996 1393
rect 1990 1388 1991 1392
rect 1995 1388 1996 1392
rect 1990 1387 1996 1388
rect 2070 1392 2076 1393
rect 2070 1388 2071 1392
rect 2075 1388 2076 1392
rect 2120 1390 2122 1393
rect 2070 1387 2076 1388
rect 2118 1389 2124 1390
rect 112 1365 114 1385
rect 136 1373 138 1385
rect 176 1373 178 1385
rect 240 1373 242 1385
rect 304 1373 306 1385
rect 368 1373 370 1385
rect 440 1373 442 1385
rect 504 1373 506 1385
rect 576 1373 578 1385
rect 648 1373 650 1385
rect 712 1373 714 1385
rect 784 1373 786 1385
rect 856 1373 858 1385
rect 928 1373 930 1385
rect 1000 1373 1002 1385
rect 1048 1373 1050 1385
rect 134 1372 140 1373
rect 134 1368 135 1372
rect 139 1368 140 1372
rect 134 1367 140 1368
rect 174 1372 180 1373
rect 174 1368 175 1372
rect 179 1368 180 1372
rect 174 1367 180 1368
rect 238 1372 244 1373
rect 238 1368 239 1372
rect 243 1368 244 1372
rect 238 1367 244 1368
rect 302 1372 308 1373
rect 302 1368 303 1372
rect 307 1368 308 1372
rect 302 1367 308 1368
rect 366 1372 372 1373
rect 366 1368 367 1372
rect 371 1368 372 1372
rect 366 1367 372 1368
rect 438 1372 444 1373
rect 438 1368 439 1372
rect 443 1368 444 1372
rect 438 1367 444 1368
rect 502 1372 508 1373
rect 502 1368 503 1372
rect 507 1368 508 1372
rect 502 1367 508 1368
rect 574 1372 580 1373
rect 574 1368 575 1372
rect 579 1368 580 1372
rect 574 1367 580 1368
rect 646 1372 652 1373
rect 646 1368 647 1372
rect 651 1368 652 1372
rect 646 1367 652 1368
rect 710 1372 716 1373
rect 710 1368 711 1372
rect 715 1368 716 1372
rect 710 1367 716 1368
rect 782 1372 788 1373
rect 782 1368 783 1372
rect 787 1368 788 1372
rect 782 1367 788 1368
rect 854 1372 860 1373
rect 854 1368 855 1372
rect 859 1368 860 1372
rect 854 1367 860 1368
rect 926 1372 932 1373
rect 926 1368 927 1372
rect 931 1368 932 1372
rect 926 1367 932 1368
rect 998 1372 1004 1373
rect 998 1368 999 1372
rect 1003 1368 1004 1372
rect 998 1367 1004 1368
rect 1046 1372 1052 1373
rect 1046 1368 1047 1372
rect 1051 1368 1052 1372
rect 1046 1367 1052 1368
rect 1096 1365 1098 1385
rect 1134 1384 1140 1385
rect 2118 1385 2119 1389
rect 2123 1385 2124 1389
rect 2118 1384 2124 1385
rect 1134 1372 1140 1373
rect 1134 1368 1135 1372
rect 1139 1368 1140 1372
rect 1134 1367 1140 1368
rect 2118 1372 2124 1373
rect 2118 1368 2119 1372
rect 2123 1368 2124 1372
rect 2118 1367 2124 1368
rect 110 1364 116 1365
rect 110 1360 111 1364
rect 115 1360 116 1364
rect 110 1359 116 1360
rect 1094 1364 1100 1365
rect 1094 1360 1095 1364
rect 1099 1360 1100 1364
rect 1094 1359 1100 1360
rect 110 1347 116 1348
rect 110 1343 111 1347
rect 115 1343 116 1347
rect 1094 1347 1100 1348
rect 1136 1347 1138 1367
rect 1334 1364 1340 1365
rect 1334 1360 1335 1364
rect 1339 1360 1340 1364
rect 1334 1359 1340 1360
rect 1374 1364 1380 1365
rect 1374 1360 1375 1364
rect 1379 1360 1380 1364
rect 1374 1359 1380 1360
rect 1414 1364 1420 1365
rect 1414 1360 1415 1364
rect 1419 1360 1420 1364
rect 1414 1359 1420 1360
rect 1454 1364 1460 1365
rect 1454 1360 1455 1364
rect 1459 1360 1460 1364
rect 1454 1359 1460 1360
rect 1494 1364 1500 1365
rect 1494 1360 1495 1364
rect 1499 1360 1500 1364
rect 1494 1359 1500 1360
rect 1534 1364 1540 1365
rect 1534 1360 1535 1364
rect 1539 1360 1540 1364
rect 1534 1359 1540 1360
rect 1582 1364 1588 1365
rect 1582 1360 1583 1364
rect 1587 1360 1588 1364
rect 1582 1359 1588 1360
rect 1646 1364 1652 1365
rect 1646 1360 1647 1364
rect 1651 1360 1652 1364
rect 1646 1359 1652 1360
rect 1718 1364 1724 1365
rect 1718 1360 1719 1364
rect 1723 1360 1724 1364
rect 1718 1359 1724 1360
rect 1806 1364 1812 1365
rect 1806 1360 1807 1364
rect 1811 1360 1812 1364
rect 1806 1359 1812 1360
rect 1894 1364 1900 1365
rect 1894 1360 1895 1364
rect 1899 1360 1900 1364
rect 1894 1359 1900 1360
rect 1990 1364 1996 1365
rect 1990 1360 1991 1364
rect 1995 1360 1996 1364
rect 1990 1359 1996 1360
rect 2070 1364 2076 1365
rect 2070 1360 2071 1364
rect 2075 1360 2076 1364
rect 2070 1359 2076 1360
rect 1336 1347 1338 1359
rect 1376 1347 1378 1359
rect 1416 1347 1418 1359
rect 1456 1347 1458 1359
rect 1496 1347 1498 1359
rect 1536 1347 1538 1359
rect 1584 1347 1586 1359
rect 1648 1347 1650 1359
rect 1720 1347 1722 1359
rect 1808 1347 1810 1359
rect 1896 1347 1898 1359
rect 1992 1347 1994 1359
rect 2072 1347 2074 1359
rect 2120 1347 2122 1367
rect 110 1342 116 1343
rect 134 1344 140 1345
rect 112 1331 114 1342
rect 134 1340 135 1344
rect 139 1340 140 1344
rect 134 1339 140 1340
rect 174 1344 180 1345
rect 174 1340 175 1344
rect 179 1340 180 1344
rect 174 1339 180 1340
rect 238 1344 244 1345
rect 238 1340 239 1344
rect 243 1340 244 1344
rect 238 1339 244 1340
rect 302 1344 308 1345
rect 302 1340 303 1344
rect 307 1340 308 1344
rect 302 1339 308 1340
rect 366 1344 372 1345
rect 366 1340 367 1344
rect 371 1340 372 1344
rect 366 1339 372 1340
rect 438 1344 444 1345
rect 438 1340 439 1344
rect 443 1340 444 1344
rect 438 1339 444 1340
rect 502 1344 508 1345
rect 502 1340 503 1344
rect 507 1340 508 1344
rect 502 1339 508 1340
rect 574 1344 580 1345
rect 574 1340 575 1344
rect 579 1340 580 1344
rect 574 1339 580 1340
rect 646 1344 652 1345
rect 646 1340 647 1344
rect 651 1340 652 1344
rect 646 1339 652 1340
rect 710 1344 716 1345
rect 710 1340 711 1344
rect 715 1340 716 1344
rect 710 1339 716 1340
rect 782 1344 788 1345
rect 782 1340 783 1344
rect 787 1340 788 1344
rect 782 1339 788 1340
rect 854 1344 860 1345
rect 854 1340 855 1344
rect 859 1340 860 1344
rect 854 1339 860 1340
rect 926 1344 932 1345
rect 926 1340 927 1344
rect 931 1340 932 1344
rect 926 1339 932 1340
rect 998 1344 1004 1345
rect 998 1340 999 1344
rect 1003 1340 1004 1344
rect 998 1339 1004 1340
rect 1046 1344 1052 1345
rect 1046 1340 1047 1344
rect 1051 1340 1052 1344
rect 1094 1343 1095 1347
rect 1099 1343 1100 1347
rect 1094 1342 1100 1343
rect 1135 1346 1139 1347
rect 1046 1339 1052 1340
rect 136 1331 138 1339
rect 176 1331 178 1339
rect 240 1331 242 1339
rect 304 1331 306 1339
rect 368 1331 370 1339
rect 440 1331 442 1339
rect 504 1331 506 1339
rect 576 1331 578 1339
rect 648 1331 650 1339
rect 712 1331 714 1339
rect 784 1331 786 1339
rect 856 1331 858 1339
rect 928 1331 930 1339
rect 1000 1331 1002 1339
rect 1048 1331 1050 1339
rect 1096 1331 1098 1342
rect 1135 1341 1139 1342
rect 1159 1346 1163 1347
rect 1159 1341 1163 1342
rect 1223 1346 1227 1347
rect 1223 1341 1227 1342
rect 1311 1346 1315 1347
rect 1311 1341 1315 1342
rect 1335 1346 1339 1347
rect 1335 1341 1339 1342
rect 1375 1346 1379 1347
rect 1375 1341 1379 1342
rect 1407 1346 1411 1347
rect 1407 1341 1411 1342
rect 1415 1346 1419 1347
rect 1415 1341 1419 1342
rect 1455 1346 1459 1347
rect 1455 1341 1459 1342
rect 1495 1346 1499 1347
rect 1495 1341 1499 1342
rect 1503 1346 1507 1347
rect 1503 1341 1507 1342
rect 1535 1346 1539 1347
rect 1535 1341 1539 1342
rect 1583 1346 1587 1347
rect 1583 1341 1587 1342
rect 1599 1346 1603 1347
rect 1599 1341 1603 1342
rect 1647 1346 1651 1347
rect 1647 1341 1651 1342
rect 1679 1346 1683 1347
rect 1679 1341 1683 1342
rect 1719 1346 1723 1347
rect 1719 1341 1723 1342
rect 1759 1346 1763 1347
rect 1759 1341 1763 1342
rect 1807 1346 1811 1347
rect 1807 1341 1811 1342
rect 1831 1346 1835 1347
rect 1831 1341 1835 1342
rect 1895 1346 1899 1347
rect 1895 1341 1899 1342
rect 1959 1346 1963 1347
rect 1959 1341 1963 1342
rect 1991 1346 1995 1347
rect 1991 1341 1995 1342
rect 2023 1346 2027 1347
rect 2023 1341 2027 1342
rect 2071 1346 2075 1347
rect 2071 1341 2075 1342
rect 2119 1346 2123 1347
rect 2119 1341 2123 1342
rect 111 1330 115 1331
rect 111 1325 115 1326
rect 135 1330 139 1331
rect 135 1325 139 1326
rect 175 1330 179 1331
rect 175 1325 179 1326
rect 215 1330 219 1331
rect 215 1325 219 1326
rect 239 1330 243 1331
rect 239 1325 243 1326
rect 255 1330 259 1331
rect 255 1325 259 1326
rect 303 1330 307 1331
rect 303 1325 307 1326
rect 319 1330 323 1331
rect 319 1325 323 1326
rect 367 1330 371 1331
rect 367 1325 371 1326
rect 391 1330 395 1331
rect 391 1325 395 1326
rect 439 1330 443 1331
rect 439 1325 443 1326
rect 463 1330 467 1331
rect 463 1325 467 1326
rect 503 1330 507 1331
rect 503 1325 507 1326
rect 543 1330 547 1331
rect 543 1325 547 1326
rect 575 1330 579 1331
rect 575 1325 579 1326
rect 623 1330 627 1331
rect 623 1325 627 1326
rect 647 1330 651 1331
rect 647 1325 651 1326
rect 703 1330 707 1331
rect 703 1325 707 1326
rect 711 1330 715 1331
rect 711 1325 715 1326
rect 783 1330 787 1331
rect 783 1325 787 1326
rect 855 1330 859 1331
rect 855 1325 859 1326
rect 863 1330 867 1331
rect 863 1325 867 1326
rect 927 1330 931 1331
rect 927 1325 931 1326
rect 943 1330 947 1331
rect 943 1325 947 1326
rect 999 1330 1003 1331
rect 999 1325 1003 1326
rect 1023 1330 1027 1331
rect 1023 1325 1027 1326
rect 1047 1330 1051 1331
rect 1047 1325 1051 1326
rect 1095 1330 1099 1331
rect 1095 1325 1099 1326
rect 112 1322 114 1325
rect 134 1324 140 1325
rect 110 1321 116 1322
rect 110 1317 111 1321
rect 115 1317 116 1321
rect 134 1320 135 1324
rect 139 1320 140 1324
rect 134 1319 140 1320
rect 174 1324 180 1325
rect 174 1320 175 1324
rect 179 1320 180 1324
rect 174 1319 180 1320
rect 214 1324 220 1325
rect 214 1320 215 1324
rect 219 1320 220 1324
rect 214 1319 220 1320
rect 254 1324 260 1325
rect 254 1320 255 1324
rect 259 1320 260 1324
rect 254 1319 260 1320
rect 318 1324 324 1325
rect 318 1320 319 1324
rect 323 1320 324 1324
rect 318 1319 324 1320
rect 390 1324 396 1325
rect 390 1320 391 1324
rect 395 1320 396 1324
rect 390 1319 396 1320
rect 462 1324 468 1325
rect 462 1320 463 1324
rect 467 1320 468 1324
rect 462 1319 468 1320
rect 542 1324 548 1325
rect 542 1320 543 1324
rect 547 1320 548 1324
rect 542 1319 548 1320
rect 622 1324 628 1325
rect 622 1320 623 1324
rect 627 1320 628 1324
rect 622 1319 628 1320
rect 702 1324 708 1325
rect 702 1320 703 1324
rect 707 1320 708 1324
rect 702 1319 708 1320
rect 782 1324 788 1325
rect 782 1320 783 1324
rect 787 1320 788 1324
rect 782 1319 788 1320
rect 862 1324 868 1325
rect 862 1320 863 1324
rect 867 1320 868 1324
rect 862 1319 868 1320
rect 942 1324 948 1325
rect 942 1320 943 1324
rect 947 1320 948 1324
rect 942 1319 948 1320
rect 1022 1324 1028 1325
rect 1022 1320 1023 1324
rect 1027 1320 1028 1324
rect 1096 1322 1098 1325
rect 1022 1319 1028 1320
rect 1094 1321 1100 1322
rect 1136 1321 1138 1341
rect 1160 1329 1162 1341
rect 1224 1329 1226 1341
rect 1312 1329 1314 1341
rect 1408 1329 1410 1341
rect 1504 1329 1506 1341
rect 1600 1329 1602 1341
rect 1680 1329 1682 1341
rect 1760 1329 1762 1341
rect 1832 1329 1834 1341
rect 1896 1329 1898 1341
rect 1960 1329 1962 1341
rect 2024 1329 2026 1341
rect 2072 1329 2074 1341
rect 1158 1328 1164 1329
rect 1158 1324 1159 1328
rect 1163 1324 1164 1328
rect 1158 1323 1164 1324
rect 1222 1328 1228 1329
rect 1222 1324 1223 1328
rect 1227 1324 1228 1328
rect 1222 1323 1228 1324
rect 1310 1328 1316 1329
rect 1310 1324 1311 1328
rect 1315 1324 1316 1328
rect 1310 1323 1316 1324
rect 1406 1328 1412 1329
rect 1406 1324 1407 1328
rect 1411 1324 1412 1328
rect 1406 1323 1412 1324
rect 1502 1328 1508 1329
rect 1502 1324 1503 1328
rect 1507 1324 1508 1328
rect 1502 1323 1508 1324
rect 1598 1328 1604 1329
rect 1598 1324 1599 1328
rect 1603 1324 1604 1328
rect 1598 1323 1604 1324
rect 1678 1328 1684 1329
rect 1678 1324 1679 1328
rect 1683 1324 1684 1328
rect 1678 1323 1684 1324
rect 1758 1328 1764 1329
rect 1758 1324 1759 1328
rect 1763 1324 1764 1328
rect 1758 1323 1764 1324
rect 1830 1328 1836 1329
rect 1830 1324 1831 1328
rect 1835 1324 1836 1328
rect 1830 1323 1836 1324
rect 1894 1328 1900 1329
rect 1894 1324 1895 1328
rect 1899 1324 1900 1328
rect 1894 1323 1900 1324
rect 1958 1328 1964 1329
rect 1958 1324 1959 1328
rect 1963 1324 1964 1328
rect 1958 1323 1964 1324
rect 2022 1328 2028 1329
rect 2022 1324 2023 1328
rect 2027 1324 2028 1328
rect 2022 1323 2028 1324
rect 2070 1328 2076 1329
rect 2070 1324 2071 1328
rect 2075 1324 2076 1328
rect 2070 1323 2076 1324
rect 2120 1321 2122 1341
rect 110 1316 116 1317
rect 1094 1317 1095 1321
rect 1099 1317 1100 1321
rect 1094 1316 1100 1317
rect 1134 1320 1140 1321
rect 1134 1316 1135 1320
rect 1139 1316 1140 1320
rect 1134 1315 1140 1316
rect 2118 1320 2124 1321
rect 2118 1316 2119 1320
rect 2123 1316 2124 1320
rect 2118 1315 2124 1316
rect 110 1304 116 1305
rect 110 1300 111 1304
rect 115 1300 116 1304
rect 110 1299 116 1300
rect 1094 1304 1100 1305
rect 1094 1300 1095 1304
rect 1099 1300 1100 1304
rect 1094 1299 1100 1300
rect 1134 1303 1140 1304
rect 1134 1299 1135 1303
rect 1139 1299 1140 1303
rect 2118 1303 2124 1304
rect 112 1275 114 1299
rect 134 1296 140 1297
rect 134 1292 135 1296
rect 139 1292 140 1296
rect 134 1291 140 1292
rect 174 1296 180 1297
rect 174 1292 175 1296
rect 179 1292 180 1296
rect 174 1291 180 1292
rect 214 1296 220 1297
rect 214 1292 215 1296
rect 219 1292 220 1296
rect 214 1291 220 1292
rect 254 1296 260 1297
rect 254 1292 255 1296
rect 259 1292 260 1296
rect 254 1291 260 1292
rect 318 1296 324 1297
rect 318 1292 319 1296
rect 323 1292 324 1296
rect 318 1291 324 1292
rect 390 1296 396 1297
rect 390 1292 391 1296
rect 395 1292 396 1296
rect 390 1291 396 1292
rect 462 1296 468 1297
rect 462 1292 463 1296
rect 467 1292 468 1296
rect 462 1291 468 1292
rect 542 1296 548 1297
rect 542 1292 543 1296
rect 547 1292 548 1296
rect 542 1291 548 1292
rect 622 1296 628 1297
rect 622 1292 623 1296
rect 627 1292 628 1296
rect 622 1291 628 1292
rect 702 1296 708 1297
rect 702 1292 703 1296
rect 707 1292 708 1296
rect 702 1291 708 1292
rect 782 1296 788 1297
rect 782 1292 783 1296
rect 787 1292 788 1296
rect 782 1291 788 1292
rect 862 1296 868 1297
rect 862 1292 863 1296
rect 867 1292 868 1296
rect 862 1291 868 1292
rect 942 1296 948 1297
rect 942 1292 943 1296
rect 947 1292 948 1296
rect 942 1291 948 1292
rect 1022 1296 1028 1297
rect 1022 1292 1023 1296
rect 1027 1292 1028 1296
rect 1022 1291 1028 1292
rect 136 1275 138 1291
rect 176 1275 178 1291
rect 216 1275 218 1291
rect 256 1275 258 1291
rect 320 1275 322 1291
rect 392 1275 394 1291
rect 464 1275 466 1291
rect 544 1275 546 1291
rect 624 1275 626 1291
rect 704 1275 706 1291
rect 784 1275 786 1291
rect 864 1275 866 1291
rect 944 1275 946 1291
rect 1024 1275 1026 1291
rect 1096 1275 1098 1299
rect 1134 1298 1140 1299
rect 1158 1300 1164 1301
rect 1136 1295 1138 1298
rect 1158 1296 1159 1300
rect 1163 1296 1164 1300
rect 1158 1295 1164 1296
rect 1222 1300 1228 1301
rect 1222 1296 1223 1300
rect 1227 1296 1228 1300
rect 1222 1295 1228 1296
rect 1310 1300 1316 1301
rect 1310 1296 1311 1300
rect 1315 1296 1316 1300
rect 1310 1295 1316 1296
rect 1406 1300 1412 1301
rect 1406 1296 1407 1300
rect 1411 1296 1412 1300
rect 1406 1295 1412 1296
rect 1502 1300 1508 1301
rect 1502 1296 1503 1300
rect 1507 1296 1508 1300
rect 1502 1295 1508 1296
rect 1598 1300 1604 1301
rect 1598 1296 1599 1300
rect 1603 1296 1604 1300
rect 1598 1295 1604 1296
rect 1678 1300 1684 1301
rect 1678 1296 1679 1300
rect 1683 1296 1684 1300
rect 1678 1295 1684 1296
rect 1758 1300 1764 1301
rect 1758 1296 1759 1300
rect 1763 1296 1764 1300
rect 1758 1295 1764 1296
rect 1830 1300 1836 1301
rect 1830 1296 1831 1300
rect 1835 1296 1836 1300
rect 1830 1295 1836 1296
rect 1894 1300 1900 1301
rect 1894 1296 1895 1300
rect 1899 1296 1900 1300
rect 1894 1295 1900 1296
rect 1958 1300 1964 1301
rect 1958 1296 1959 1300
rect 1963 1296 1964 1300
rect 1958 1295 1964 1296
rect 2022 1300 2028 1301
rect 2022 1296 2023 1300
rect 2027 1296 2028 1300
rect 2022 1295 2028 1296
rect 2070 1300 2076 1301
rect 2070 1296 2071 1300
rect 2075 1296 2076 1300
rect 2118 1299 2119 1303
rect 2123 1299 2124 1303
rect 2118 1298 2124 1299
rect 2070 1295 2076 1296
rect 2120 1295 2122 1298
rect 1135 1294 1139 1295
rect 1135 1289 1139 1290
rect 1159 1294 1163 1295
rect 1159 1289 1163 1290
rect 1175 1294 1179 1295
rect 1175 1289 1179 1290
rect 1223 1294 1227 1295
rect 1223 1289 1227 1290
rect 1231 1294 1235 1295
rect 1231 1289 1235 1290
rect 1303 1294 1307 1295
rect 1303 1289 1307 1290
rect 1311 1294 1315 1295
rect 1311 1289 1315 1290
rect 1391 1294 1395 1295
rect 1391 1289 1395 1290
rect 1407 1294 1411 1295
rect 1407 1289 1411 1290
rect 1479 1294 1483 1295
rect 1479 1289 1483 1290
rect 1503 1294 1507 1295
rect 1503 1289 1507 1290
rect 1567 1294 1571 1295
rect 1567 1289 1571 1290
rect 1599 1294 1603 1295
rect 1599 1289 1603 1290
rect 1655 1294 1659 1295
rect 1655 1289 1659 1290
rect 1679 1294 1683 1295
rect 1679 1289 1683 1290
rect 1743 1294 1747 1295
rect 1743 1289 1747 1290
rect 1759 1294 1763 1295
rect 1759 1289 1763 1290
rect 1831 1294 1835 1295
rect 1831 1289 1835 1290
rect 1895 1294 1899 1295
rect 1895 1289 1899 1290
rect 1919 1294 1923 1295
rect 1919 1289 1923 1290
rect 1959 1294 1963 1295
rect 1959 1289 1963 1290
rect 2007 1294 2011 1295
rect 2007 1289 2011 1290
rect 2023 1294 2027 1295
rect 2023 1289 2027 1290
rect 2071 1294 2075 1295
rect 2071 1289 2075 1290
rect 2119 1294 2123 1295
rect 2119 1289 2123 1290
rect 1136 1286 1138 1289
rect 1174 1288 1180 1289
rect 1134 1285 1140 1286
rect 1134 1281 1135 1285
rect 1139 1281 1140 1285
rect 1174 1284 1175 1288
rect 1179 1284 1180 1288
rect 1174 1283 1180 1284
rect 1230 1288 1236 1289
rect 1230 1284 1231 1288
rect 1235 1284 1236 1288
rect 1230 1283 1236 1284
rect 1302 1288 1308 1289
rect 1302 1284 1303 1288
rect 1307 1284 1308 1288
rect 1302 1283 1308 1284
rect 1390 1288 1396 1289
rect 1390 1284 1391 1288
rect 1395 1284 1396 1288
rect 1390 1283 1396 1284
rect 1478 1288 1484 1289
rect 1478 1284 1479 1288
rect 1483 1284 1484 1288
rect 1478 1283 1484 1284
rect 1566 1288 1572 1289
rect 1566 1284 1567 1288
rect 1571 1284 1572 1288
rect 1566 1283 1572 1284
rect 1654 1288 1660 1289
rect 1654 1284 1655 1288
rect 1659 1284 1660 1288
rect 1654 1283 1660 1284
rect 1742 1288 1748 1289
rect 1742 1284 1743 1288
rect 1747 1284 1748 1288
rect 1742 1283 1748 1284
rect 1830 1288 1836 1289
rect 1830 1284 1831 1288
rect 1835 1284 1836 1288
rect 1830 1283 1836 1284
rect 1918 1288 1924 1289
rect 1918 1284 1919 1288
rect 1923 1284 1924 1288
rect 1918 1283 1924 1284
rect 2006 1288 2012 1289
rect 2006 1284 2007 1288
rect 2011 1284 2012 1288
rect 2006 1283 2012 1284
rect 2070 1288 2076 1289
rect 2070 1284 2071 1288
rect 2075 1284 2076 1288
rect 2120 1286 2122 1289
rect 2070 1283 2076 1284
rect 2118 1285 2124 1286
rect 1134 1280 1140 1281
rect 2118 1281 2119 1285
rect 2123 1281 2124 1285
rect 2118 1280 2124 1281
rect 111 1274 115 1275
rect 111 1269 115 1270
rect 135 1274 139 1275
rect 135 1269 139 1270
rect 175 1274 179 1275
rect 175 1269 179 1270
rect 215 1274 219 1275
rect 215 1269 219 1270
rect 255 1274 259 1275
rect 255 1269 259 1270
rect 319 1274 323 1275
rect 319 1269 323 1270
rect 391 1274 395 1275
rect 391 1269 395 1270
rect 399 1274 403 1275
rect 399 1269 403 1270
rect 463 1274 467 1275
rect 463 1269 467 1270
rect 487 1274 491 1275
rect 487 1269 491 1270
rect 543 1274 547 1275
rect 543 1269 547 1270
rect 583 1274 587 1275
rect 583 1269 587 1270
rect 623 1274 627 1275
rect 623 1269 627 1270
rect 687 1274 691 1275
rect 687 1269 691 1270
rect 703 1274 707 1275
rect 703 1269 707 1270
rect 783 1274 787 1275
rect 783 1269 787 1270
rect 799 1274 803 1275
rect 799 1269 803 1270
rect 863 1274 867 1275
rect 863 1269 867 1270
rect 919 1274 923 1275
rect 919 1269 923 1270
rect 943 1274 947 1275
rect 943 1269 947 1270
rect 1023 1274 1027 1275
rect 1023 1269 1027 1270
rect 1047 1274 1051 1275
rect 1047 1269 1051 1270
rect 1095 1274 1099 1275
rect 1095 1269 1099 1270
rect 112 1249 114 1269
rect 136 1257 138 1269
rect 176 1257 178 1269
rect 216 1257 218 1269
rect 256 1257 258 1269
rect 320 1257 322 1269
rect 400 1257 402 1269
rect 488 1257 490 1269
rect 584 1257 586 1269
rect 688 1257 690 1269
rect 800 1257 802 1269
rect 920 1257 922 1269
rect 1048 1257 1050 1269
rect 134 1256 140 1257
rect 134 1252 135 1256
rect 139 1252 140 1256
rect 134 1251 140 1252
rect 174 1256 180 1257
rect 174 1252 175 1256
rect 179 1252 180 1256
rect 174 1251 180 1252
rect 214 1256 220 1257
rect 214 1252 215 1256
rect 219 1252 220 1256
rect 214 1251 220 1252
rect 254 1256 260 1257
rect 254 1252 255 1256
rect 259 1252 260 1256
rect 254 1251 260 1252
rect 318 1256 324 1257
rect 318 1252 319 1256
rect 323 1252 324 1256
rect 318 1251 324 1252
rect 398 1256 404 1257
rect 398 1252 399 1256
rect 403 1252 404 1256
rect 398 1251 404 1252
rect 486 1256 492 1257
rect 486 1252 487 1256
rect 491 1252 492 1256
rect 486 1251 492 1252
rect 582 1256 588 1257
rect 582 1252 583 1256
rect 587 1252 588 1256
rect 582 1251 588 1252
rect 686 1256 692 1257
rect 686 1252 687 1256
rect 691 1252 692 1256
rect 686 1251 692 1252
rect 798 1256 804 1257
rect 798 1252 799 1256
rect 803 1252 804 1256
rect 798 1251 804 1252
rect 918 1256 924 1257
rect 918 1252 919 1256
rect 923 1252 924 1256
rect 918 1251 924 1252
rect 1046 1256 1052 1257
rect 1046 1252 1047 1256
rect 1051 1252 1052 1256
rect 1046 1251 1052 1252
rect 1096 1249 1098 1269
rect 1134 1268 1140 1269
rect 1134 1264 1135 1268
rect 1139 1264 1140 1268
rect 1134 1263 1140 1264
rect 2118 1268 2124 1269
rect 2118 1264 2119 1268
rect 2123 1264 2124 1268
rect 2118 1263 2124 1264
rect 110 1248 116 1249
rect 110 1244 111 1248
rect 115 1244 116 1248
rect 110 1243 116 1244
rect 1094 1248 1100 1249
rect 1094 1244 1095 1248
rect 1099 1244 1100 1248
rect 1094 1243 1100 1244
rect 1136 1239 1138 1263
rect 1174 1260 1180 1261
rect 1174 1256 1175 1260
rect 1179 1256 1180 1260
rect 1174 1255 1180 1256
rect 1230 1260 1236 1261
rect 1230 1256 1231 1260
rect 1235 1256 1236 1260
rect 1230 1255 1236 1256
rect 1302 1260 1308 1261
rect 1302 1256 1303 1260
rect 1307 1256 1308 1260
rect 1302 1255 1308 1256
rect 1390 1260 1396 1261
rect 1390 1256 1391 1260
rect 1395 1256 1396 1260
rect 1390 1255 1396 1256
rect 1478 1260 1484 1261
rect 1478 1256 1479 1260
rect 1483 1256 1484 1260
rect 1478 1255 1484 1256
rect 1566 1260 1572 1261
rect 1566 1256 1567 1260
rect 1571 1256 1572 1260
rect 1566 1255 1572 1256
rect 1654 1260 1660 1261
rect 1654 1256 1655 1260
rect 1659 1256 1660 1260
rect 1654 1255 1660 1256
rect 1742 1260 1748 1261
rect 1742 1256 1743 1260
rect 1747 1256 1748 1260
rect 1742 1255 1748 1256
rect 1830 1260 1836 1261
rect 1830 1256 1831 1260
rect 1835 1256 1836 1260
rect 1830 1255 1836 1256
rect 1918 1260 1924 1261
rect 1918 1256 1919 1260
rect 1923 1256 1924 1260
rect 1918 1255 1924 1256
rect 2006 1260 2012 1261
rect 2006 1256 2007 1260
rect 2011 1256 2012 1260
rect 2006 1255 2012 1256
rect 2070 1260 2076 1261
rect 2070 1256 2071 1260
rect 2075 1256 2076 1260
rect 2070 1255 2076 1256
rect 1176 1239 1178 1255
rect 1232 1239 1234 1255
rect 1304 1239 1306 1255
rect 1392 1239 1394 1255
rect 1480 1239 1482 1255
rect 1568 1239 1570 1255
rect 1656 1239 1658 1255
rect 1744 1239 1746 1255
rect 1832 1239 1834 1255
rect 1920 1239 1922 1255
rect 2008 1239 2010 1255
rect 2072 1239 2074 1255
rect 2120 1239 2122 1263
rect 1135 1238 1139 1239
rect 1135 1233 1139 1234
rect 1175 1238 1179 1239
rect 1175 1233 1179 1234
rect 1231 1238 1235 1239
rect 1231 1233 1235 1234
rect 1287 1238 1291 1239
rect 1287 1233 1291 1234
rect 1303 1238 1307 1239
rect 1303 1233 1307 1234
rect 1327 1238 1331 1239
rect 1327 1233 1331 1234
rect 1375 1238 1379 1239
rect 1375 1233 1379 1234
rect 1391 1238 1395 1239
rect 1391 1233 1395 1234
rect 1431 1238 1435 1239
rect 1431 1233 1435 1234
rect 1479 1238 1483 1239
rect 1479 1233 1483 1234
rect 1495 1238 1499 1239
rect 1495 1233 1499 1234
rect 1559 1238 1563 1239
rect 1559 1233 1563 1234
rect 1567 1238 1571 1239
rect 1567 1233 1571 1234
rect 1623 1238 1627 1239
rect 1623 1233 1627 1234
rect 1655 1238 1659 1239
rect 1655 1233 1659 1234
rect 1679 1238 1683 1239
rect 1679 1233 1683 1234
rect 1735 1238 1739 1239
rect 1735 1233 1739 1234
rect 1743 1238 1747 1239
rect 1743 1233 1747 1234
rect 1791 1238 1795 1239
rect 1791 1233 1795 1234
rect 1831 1238 1835 1239
rect 1831 1233 1835 1234
rect 1847 1238 1851 1239
rect 1847 1233 1851 1234
rect 1903 1238 1907 1239
rect 1903 1233 1907 1234
rect 1919 1238 1923 1239
rect 1919 1233 1923 1234
rect 1967 1238 1971 1239
rect 1967 1233 1971 1234
rect 2007 1238 2011 1239
rect 2007 1233 2011 1234
rect 2031 1238 2035 1239
rect 2031 1233 2035 1234
rect 2071 1238 2075 1239
rect 2071 1233 2075 1234
rect 2119 1238 2123 1239
rect 2119 1233 2123 1234
rect 110 1231 116 1232
rect 110 1227 111 1231
rect 115 1227 116 1231
rect 1094 1231 1100 1232
rect 110 1226 116 1227
rect 134 1228 140 1229
rect 112 1219 114 1226
rect 134 1224 135 1228
rect 139 1224 140 1228
rect 134 1223 140 1224
rect 174 1228 180 1229
rect 174 1224 175 1228
rect 179 1224 180 1228
rect 174 1223 180 1224
rect 214 1228 220 1229
rect 214 1224 215 1228
rect 219 1224 220 1228
rect 214 1223 220 1224
rect 254 1228 260 1229
rect 254 1224 255 1228
rect 259 1224 260 1228
rect 254 1223 260 1224
rect 318 1228 324 1229
rect 318 1224 319 1228
rect 323 1224 324 1228
rect 318 1223 324 1224
rect 398 1228 404 1229
rect 398 1224 399 1228
rect 403 1224 404 1228
rect 398 1223 404 1224
rect 486 1228 492 1229
rect 486 1224 487 1228
rect 491 1224 492 1228
rect 486 1223 492 1224
rect 582 1228 588 1229
rect 582 1224 583 1228
rect 587 1224 588 1228
rect 582 1223 588 1224
rect 686 1228 692 1229
rect 686 1224 687 1228
rect 691 1224 692 1228
rect 686 1223 692 1224
rect 798 1228 804 1229
rect 798 1224 799 1228
rect 803 1224 804 1228
rect 798 1223 804 1224
rect 918 1228 924 1229
rect 918 1224 919 1228
rect 923 1224 924 1228
rect 918 1223 924 1224
rect 1046 1228 1052 1229
rect 1046 1224 1047 1228
rect 1051 1224 1052 1228
rect 1094 1227 1095 1231
rect 1099 1227 1100 1231
rect 1094 1226 1100 1227
rect 1046 1223 1052 1224
rect 136 1219 138 1223
rect 176 1219 178 1223
rect 216 1219 218 1223
rect 256 1219 258 1223
rect 320 1219 322 1223
rect 400 1219 402 1223
rect 488 1219 490 1223
rect 584 1219 586 1223
rect 688 1219 690 1223
rect 800 1219 802 1223
rect 920 1219 922 1223
rect 1048 1219 1050 1223
rect 1096 1219 1098 1226
rect 111 1218 115 1219
rect 111 1213 115 1214
rect 135 1218 139 1219
rect 135 1213 139 1214
rect 175 1218 179 1219
rect 175 1213 179 1214
rect 215 1218 219 1219
rect 215 1213 219 1214
rect 255 1218 259 1219
rect 255 1213 259 1214
rect 271 1218 275 1219
rect 271 1213 275 1214
rect 311 1218 315 1219
rect 311 1213 315 1214
rect 319 1218 323 1219
rect 319 1213 323 1214
rect 351 1218 355 1219
rect 351 1213 355 1214
rect 399 1218 403 1219
rect 399 1213 403 1214
rect 447 1218 451 1219
rect 447 1213 451 1214
rect 487 1218 491 1219
rect 487 1213 491 1214
rect 495 1218 499 1219
rect 495 1213 499 1214
rect 551 1218 555 1219
rect 551 1213 555 1214
rect 583 1218 587 1219
rect 583 1213 587 1214
rect 607 1218 611 1219
rect 607 1213 611 1214
rect 671 1218 675 1219
rect 671 1213 675 1214
rect 687 1218 691 1219
rect 687 1213 691 1214
rect 743 1218 747 1219
rect 743 1213 747 1214
rect 799 1218 803 1219
rect 799 1213 803 1214
rect 815 1218 819 1219
rect 815 1213 819 1214
rect 895 1218 899 1219
rect 895 1213 899 1214
rect 919 1218 923 1219
rect 919 1213 923 1214
rect 983 1218 987 1219
rect 983 1213 987 1214
rect 1047 1218 1051 1219
rect 1047 1213 1051 1214
rect 1095 1218 1099 1219
rect 1095 1213 1099 1214
rect 1136 1213 1138 1233
rect 1288 1221 1290 1233
rect 1328 1221 1330 1233
rect 1376 1221 1378 1233
rect 1432 1221 1434 1233
rect 1496 1221 1498 1233
rect 1560 1221 1562 1233
rect 1624 1221 1626 1233
rect 1680 1221 1682 1233
rect 1736 1221 1738 1233
rect 1792 1221 1794 1233
rect 1848 1221 1850 1233
rect 1904 1221 1906 1233
rect 1968 1221 1970 1233
rect 2032 1221 2034 1233
rect 2072 1221 2074 1233
rect 1286 1220 1292 1221
rect 1286 1216 1287 1220
rect 1291 1216 1292 1220
rect 1286 1215 1292 1216
rect 1326 1220 1332 1221
rect 1326 1216 1327 1220
rect 1331 1216 1332 1220
rect 1326 1215 1332 1216
rect 1374 1220 1380 1221
rect 1374 1216 1375 1220
rect 1379 1216 1380 1220
rect 1374 1215 1380 1216
rect 1430 1220 1436 1221
rect 1430 1216 1431 1220
rect 1435 1216 1436 1220
rect 1430 1215 1436 1216
rect 1494 1220 1500 1221
rect 1494 1216 1495 1220
rect 1499 1216 1500 1220
rect 1494 1215 1500 1216
rect 1558 1220 1564 1221
rect 1558 1216 1559 1220
rect 1563 1216 1564 1220
rect 1558 1215 1564 1216
rect 1622 1220 1628 1221
rect 1622 1216 1623 1220
rect 1627 1216 1628 1220
rect 1622 1215 1628 1216
rect 1678 1220 1684 1221
rect 1678 1216 1679 1220
rect 1683 1216 1684 1220
rect 1678 1215 1684 1216
rect 1734 1220 1740 1221
rect 1734 1216 1735 1220
rect 1739 1216 1740 1220
rect 1734 1215 1740 1216
rect 1790 1220 1796 1221
rect 1790 1216 1791 1220
rect 1795 1216 1796 1220
rect 1790 1215 1796 1216
rect 1846 1220 1852 1221
rect 1846 1216 1847 1220
rect 1851 1216 1852 1220
rect 1846 1215 1852 1216
rect 1902 1220 1908 1221
rect 1902 1216 1903 1220
rect 1907 1216 1908 1220
rect 1902 1215 1908 1216
rect 1966 1220 1972 1221
rect 1966 1216 1967 1220
rect 1971 1216 1972 1220
rect 1966 1215 1972 1216
rect 2030 1220 2036 1221
rect 2030 1216 2031 1220
rect 2035 1216 2036 1220
rect 2030 1215 2036 1216
rect 2070 1220 2076 1221
rect 2070 1216 2071 1220
rect 2075 1216 2076 1220
rect 2070 1215 2076 1216
rect 2120 1213 2122 1233
rect 112 1210 114 1213
rect 270 1212 276 1213
rect 110 1209 116 1210
rect 110 1205 111 1209
rect 115 1205 116 1209
rect 270 1208 271 1212
rect 275 1208 276 1212
rect 270 1207 276 1208
rect 310 1212 316 1213
rect 310 1208 311 1212
rect 315 1208 316 1212
rect 310 1207 316 1208
rect 350 1212 356 1213
rect 350 1208 351 1212
rect 355 1208 356 1212
rect 350 1207 356 1208
rect 398 1212 404 1213
rect 398 1208 399 1212
rect 403 1208 404 1212
rect 398 1207 404 1208
rect 446 1212 452 1213
rect 446 1208 447 1212
rect 451 1208 452 1212
rect 446 1207 452 1208
rect 494 1212 500 1213
rect 494 1208 495 1212
rect 499 1208 500 1212
rect 494 1207 500 1208
rect 550 1212 556 1213
rect 550 1208 551 1212
rect 555 1208 556 1212
rect 550 1207 556 1208
rect 606 1212 612 1213
rect 606 1208 607 1212
rect 611 1208 612 1212
rect 606 1207 612 1208
rect 670 1212 676 1213
rect 670 1208 671 1212
rect 675 1208 676 1212
rect 670 1207 676 1208
rect 742 1212 748 1213
rect 742 1208 743 1212
rect 747 1208 748 1212
rect 742 1207 748 1208
rect 814 1212 820 1213
rect 814 1208 815 1212
rect 819 1208 820 1212
rect 814 1207 820 1208
rect 894 1212 900 1213
rect 894 1208 895 1212
rect 899 1208 900 1212
rect 894 1207 900 1208
rect 982 1212 988 1213
rect 982 1208 983 1212
rect 987 1208 988 1212
rect 1096 1210 1098 1213
rect 1134 1212 1140 1213
rect 982 1207 988 1208
rect 1094 1209 1100 1210
rect 110 1204 116 1205
rect 1094 1205 1095 1209
rect 1099 1205 1100 1209
rect 1134 1208 1135 1212
rect 1139 1208 1140 1212
rect 1134 1207 1140 1208
rect 2118 1212 2124 1213
rect 2118 1208 2119 1212
rect 2123 1208 2124 1212
rect 2118 1207 2124 1208
rect 1094 1204 1100 1205
rect 1134 1195 1140 1196
rect 110 1192 116 1193
rect 110 1188 111 1192
rect 115 1188 116 1192
rect 110 1187 116 1188
rect 1094 1192 1100 1193
rect 1094 1188 1095 1192
rect 1099 1188 1100 1192
rect 1134 1191 1135 1195
rect 1139 1191 1140 1195
rect 2118 1195 2124 1196
rect 1134 1190 1140 1191
rect 1286 1192 1292 1193
rect 1094 1187 1100 1188
rect 1136 1187 1138 1190
rect 1286 1188 1287 1192
rect 1291 1188 1292 1192
rect 1286 1187 1292 1188
rect 1326 1192 1332 1193
rect 1326 1188 1327 1192
rect 1331 1188 1332 1192
rect 1326 1187 1332 1188
rect 1374 1192 1380 1193
rect 1374 1188 1375 1192
rect 1379 1188 1380 1192
rect 1374 1187 1380 1188
rect 1430 1192 1436 1193
rect 1430 1188 1431 1192
rect 1435 1188 1436 1192
rect 1430 1187 1436 1188
rect 1494 1192 1500 1193
rect 1494 1188 1495 1192
rect 1499 1188 1500 1192
rect 1494 1187 1500 1188
rect 1558 1192 1564 1193
rect 1558 1188 1559 1192
rect 1563 1188 1564 1192
rect 1558 1187 1564 1188
rect 1622 1192 1628 1193
rect 1622 1188 1623 1192
rect 1627 1188 1628 1192
rect 1622 1187 1628 1188
rect 1678 1192 1684 1193
rect 1678 1188 1679 1192
rect 1683 1188 1684 1192
rect 1678 1187 1684 1188
rect 1734 1192 1740 1193
rect 1734 1188 1735 1192
rect 1739 1188 1740 1192
rect 1734 1187 1740 1188
rect 1790 1192 1796 1193
rect 1790 1188 1791 1192
rect 1795 1188 1796 1192
rect 1790 1187 1796 1188
rect 1846 1192 1852 1193
rect 1846 1188 1847 1192
rect 1851 1188 1852 1192
rect 1846 1187 1852 1188
rect 1902 1192 1908 1193
rect 1902 1188 1903 1192
rect 1907 1188 1908 1192
rect 1902 1187 1908 1188
rect 1966 1192 1972 1193
rect 1966 1188 1967 1192
rect 1971 1188 1972 1192
rect 1966 1187 1972 1188
rect 2030 1192 2036 1193
rect 2030 1188 2031 1192
rect 2035 1188 2036 1192
rect 2030 1187 2036 1188
rect 2070 1192 2076 1193
rect 2070 1188 2071 1192
rect 2075 1188 2076 1192
rect 2118 1191 2119 1195
rect 2123 1191 2124 1195
rect 2118 1190 2124 1191
rect 2070 1187 2076 1188
rect 2120 1187 2122 1190
rect 112 1163 114 1187
rect 270 1184 276 1185
rect 270 1180 271 1184
rect 275 1180 276 1184
rect 270 1179 276 1180
rect 310 1184 316 1185
rect 310 1180 311 1184
rect 315 1180 316 1184
rect 310 1179 316 1180
rect 350 1184 356 1185
rect 350 1180 351 1184
rect 355 1180 356 1184
rect 350 1179 356 1180
rect 398 1184 404 1185
rect 398 1180 399 1184
rect 403 1180 404 1184
rect 398 1179 404 1180
rect 446 1184 452 1185
rect 446 1180 447 1184
rect 451 1180 452 1184
rect 446 1179 452 1180
rect 494 1184 500 1185
rect 494 1180 495 1184
rect 499 1180 500 1184
rect 494 1179 500 1180
rect 550 1184 556 1185
rect 550 1180 551 1184
rect 555 1180 556 1184
rect 550 1179 556 1180
rect 606 1184 612 1185
rect 606 1180 607 1184
rect 611 1180 612 1184
rect 606 1179 612 1180
rect 670 1184 676 1185
rect 670 1180 671 1184
rect 675 1180 676 1184
rect 670 1179 676 1180
rect 742 1184 748 1185
rect 742 1180 743 1184
rect 747 1180 748 1184
rect 742 1179 748 1180
rect 814 1184 820 1185
rect 814 1180 815 1184
rect 819 1180 820 1184
rect 814 1179 820 1180
rect 894 1184 900 1185
rect 894 1180 895 1184
rect 899 1180 900 1184
rect 894 1179 900 1180
rect 982 1184 988 1185
rect 982 1180 983 1184
rect 987 1180 988 1184
rect 982 1179 988 1180
rect 272 1163 274 1179
rect 312 1163 314 1179
rect 352 1163 354 1179
rect 400 1163 402 1179
rect 448 1163 450 1179
rect 496 1163 498 1179
rect 552 1163 554 1179
rect 608 1163 610 1179
rect 672 1163 674 1179
rect 744 1163 746 1179
rect 816 1163 818 1179
rect 896 1163 898 1179
rect 984 1163 986 1179
rect 1096 1163 1098 1187
rect 1135 1186 1139 1187
rect 1135 1181 1139 1182
rect 1159 1186 1163 1187
rect 1159 1181 1163 1182
rect 1207 1186 1211 1187
rect 1207 1181 1211 1182
rect 1279 1186 1283 1187
rect 1279 1181 1283 1182
rect 1287 1186 1291 1187
rect 1287 1181 1291 1182
rect 1327 1186 1331 1187
rect 1327 1181 1331 1182
rect 1351 1186 1355 1187
rect 1351 1181 1355 1182
rect 1375 1186 1379 1187
rect 1375 1181 1379 1182
rect 1423 1186 1427 1187
rect 1423 1181 1427 1182
rect 1431 1186 1435 1187
rect 1431 1181 1435 1182
rect 1487 1186 1491 1187
rect 1487 1181 1491 1182
rect 1495 1186 1499 1187
rect 1495 1181 1499 1182
rect 1559 1186 1563 1187
rect 1559 1181 1563 1182
rect 1623 1186 1627 1187
rect 1623 1181 1627 1182
rect 1631 1186 1635 1187
rect 1631 1181 1635 1182
rect 1679 1186 1683 1187
rect 1679 1181 1683 1182
rect 1711 1186 1715 1187
rect 1711 1181 1715 1182
rect 1735 1186 1739 1187
rect 1735 1181 1739 1182
rect 1791 1186 1795 1187
rect 1791 1181 1795 1182
rect 1799 1186 1803 1187
rect 1799 1181 1803 1182
rect 1847 1186 1851 1187
rect 1847 1181 1851 1182
rect 1887 1186 1891 1187
rect 1887 1181 1891 1182
rect 1903 1186 1907 1187
rect 1903 1181 1907 1182
rect 1967 1186 1971 1187
rect 1967 1181 1971 1182
rect 1983 1186 1987 1187
rect 1983 1181 1987 1182
rect 2031 1186 2035 1187
rect 2031 1181 2035 1182
rect 2071 1186 2075 1187
rect 2071 1181 2075 1182
rect 2119 1186 2123 1187
rect 2119 1181 2123 1182
rect 1136 1178 1138 1181
rect 1158 1180 1164 1181
rect 1134 1177 1140 1178
rect 1134 1173 1135 1177
rect 1139 1173 1140 1177
rect 1158 1176 1159 1180
rect 1163 1176 1164 1180
rect 1158 1175 1164 1176
rect 1206 1180 1212 1181
rect 1206 1176 1207 1180
rect 1211 1176 1212 1180
rect 1206 1175 1212 1176
rect 1278 1180 1284 1181
rect 1278 1176 1279 1180
rect 1283 1176 1284 1180
rect 1278 1175 1284 1176
rect 1350 1180 1356 1181
rect 1350 1176 1351 1180
rect 1355 1176 1356 1180
rect 1350 1175 1356 1176
rect 1422 1180 1428 1181
rect 1422 1176 1423 1180
rect 1427 1176 1428 1180
rect 1422 1175 1428 1176
rect 1486 1180 1492 1181
rect 1486 1176 1487 1180
rect 1491 1176 1492 1180
rect 1486 1175 1492 1176
rect 1558 1180 1564 1181
rect 1558 1176 1559 1180
rect 1563 1176 1564 1180
rect 1558 1175 1564 1176
rect 1630 1180 1636 1181
rect 1630 1176 1631 1180
rect 1635 1176 1636 1180
rect 1630 1175 1636 1176
rect 1710 1180 1716 1181
rect 1710 1176 1711 1180
rect 1715 1176 1716 1180
rect 1710 1175 1716 1176
rect 1798 1180 1804 1181
rect 1798 1176 1799 1180
rect 1803 1176 1804 1180
rect 1798 1175 1804 1176
rect 1886 1180 1892 1181
rect 1886 1176 1887 1180
rect 1891 1176 1892 1180
rect 1886 1175 1892 1176
rect 1982 1180 1988 1181
rect 1982 1176 1983 1180
rect 1987 1176 1988 1180
rect 1982 1175 1988 1176
rect 2070 1180 2076 1181
rect 2070 1176 2071 1180
rect 2075 1176 2076 1180
rect 2120 1178 2122 1181
rect 2070 1175 2076 1176
rect 2118 1177 2124 1178
rect 1134 1172 1140 1173
rect 2118 1173 2119 1177
rect 2123 1173 2124 1177
rect 2118 1172 2124 1173
rect 111 1162 115 1163
rect 111 1157 115 1158
rect 271 1162 275 1163
rect 271 1157 275 1158
rect 311 1162 315 1163
rect 311 1157 315 1158
rect 351 1162 355 1163
rect 351 1157 355 1158
rect 399 1162 403 1163
rect 399 1157 403 1158
rect 439 1162 443 1163
rect 439 1157 443 1158
rect 447 1162 451 1163
rect 447 1157 451 1158
rect 479 1162 483 1163
rect 479 1157 483 1158
rect 495 1162 499 1163
rect 495 1157 499 1158
rect 527 1162 531 1163
rect 527 1157 531 1158
rect 551 1162 555 1163
rect 551 1157 555 1158
rect 575 1162 579 1163
rect 575 1157 579 1158
rect 607 1162 611 1163
rect 607 1157 611 1158
rect 623 1162 627 1163
rect 623 1157 627 1158
rect 671 1162 675 1163
rect 671 1157 675 1158
rect 719 1162 723 1163
rect 719 1157 723 1158
rect 743 1162 747 1163
rect 743 1157 747 1158
rect 775 1162 779 1163
rect 775 1157 779 1158
rect 815 1162 819 1163
rect 815 1157 819 1158
rect 831 1162 835 1163
rect 831 1157 835 1158
rect 887 1162 891 1163
rect 887 1157 891 1158
rect 895 1162 899 1163
rect 895 1157 899 1158
rect 943 1162 947 1163
rect 943 1157 947 1158
rect 983 1162 987 1163
rect 983 1157 987 1158
rect 1007 1162 1011 1163
rect 1007 1157 1011 1158
rect 1047 1162 1051 1163
rect 1047 1157 1051 1158
rect 1095 1162 1099 1163
rect 1095 1157 1099 1158
rect 1134 1160 1140 1161
rect 112 1137 114 1157
rect 400 1145 402 1157
rect 440 1145 442 1157
rect 480 1145 482 1157
rect 528 1145 530 1157
rect 576 1145 578 1157
rect 624 1145 626 1157
rect 672 1145 674 1157
rect 720 1145 722 1157
rect 776 1145 778 1157
rect 832 1145 834 1157
rect 888 1145 890 1157
rect 944 1145 946 1157
rect 1008 1145 1010 1157
rect 1048 1145 1050 1157
rect 398 1144 404 1145
rect 398 1140 399 1144
rect 403 1140 404 1144
rect 398 1139 404 1140
rect 438 1144 444 1145
rect 438 1140 439 1144
rect 443 1140 444 1144
rect 438 1139 444 1140
rect 478 1144 484 1145
rect 478 1140 479 1144
rect 483 1140 484 1144
rect 478 1139 484 1140
rect 526 1144 532 1145
rect 526 1140 527 1144
rect 531 1140 532 1144
rect 526 1139 532 1140
rect 574 1144 580 1145
rect 574 1140 575 1144
rect 579 1140 580 1144
rect 574 1139 580 1140
rect 622 1144 628 1145
rect 622 1140 623 1144
rect 627 1140 628 1144
rect 622 1139 628 1140
rect 670 1144 676 1145
rect 670 1140 671 1144
rect 675 1140 676 1144
rect 670 1139 676 1140
rect 718 1144 724 1145
rect 718 1140 719 1144
rect 723 1140 724 1144
rect 718 1139 724 1140
rect 774 1144 780 1145
rect 774 1140 775 1144
rect 779 1140 780 1144
rect 774 1139 780 1140
rect 830 1144 836 1145
rect 830 1140 831 1144
rect 835 1140 836 1144
rect 830 1139 836 1140
rect 886 1144 892 1145
rect 886 1140 887 1144
rect 891 1140 892 1144
rect 886 1139 892 1140
rect 942 1144 948 1145
rect 942 1140 943 1144
rect 947 1140 948 1144
rect 942 1139 948 1140
rect 1006 1144 1012 1145
rect 1006 1140 1007 1144
rect 1011 1140 1012 1144
rect 1006 1139 1012 1140
rect 1046 1144 1052 1145
rect 1046 1140 1047 1144
rect 1051 1140 1052 1144
rect 1046 1139 1052 1140
rect 1096 1137 1098 1157
rect 1134 1156 1135 1160
rect 1139 1156 1140 1160
rect 1134 1155 1140 1156
rect 2118 1160 2124 1161
rect 2118 1156 2119 1160
rect 2123 1156 2124 1160
rect 2118 1155 2124 1156
rect 110 1136 116 1137
rect 110 1132 111 1136
rect 115 1132 116 1136
rect 110 1131 116 1132
rect 1094 1136 1100 1137
rect 1094 1132 1095 1136
rect 1099 1132 1100 1136
rect 1094 1131 1100 1132
rect 1136 1131 1138 1155
rect 1158 1152 1164 1153
rect 1158 1148 1159 1152
rect 1163 1148 1164 1152
rect 1158 1147 1164 1148
rect 1206 1152 1212 1153
rect 1206 1148 1207 1152
rect 1211 1148 1212 1152
rect 1206 1147 1212 1148
rect 1278 1152 1284 1153
rect 1278 1148 1279 1152
rect 1283 1148 1284 1152
rect 1278 1147 1284 1148
rect 1350 1152 1356 1153
rect 1350 1148 1351 1152
rect 1355 1148 1356 1152
rect 1350 1147 1356 1148
rect 1422 1152 1428 1153
rect 1422 1148 1423 1152
rect 1427 1148 1428 1152
rect 1422 1147 1428 1148
rect 1486 1152 1492 1153
rect 1486 1148 1487 1152
rect 1491 1148 1492 1152
rect 1486 1147 1492 1148
rect 1558 1152 1564 1153
rect 1558 1148 1559 1152
rect 1563 1148 1564 1152
rect 1558 1147 1564 1148
rect 1630 1152 1636 1153
rect 1630 1148 1631 1152
rect 1635 1148 1636 1152
rect 1630 1147 1636 1148
rect 1710 1152 1716 1153
rect 1710 1148 1711 1152
rect 1715 1148 1716 1152
rect 1710 1147 1716 1148
rect 1798 1152 1804 1153
rect 1798 1148 1799 1152
rect 1803 1148 1804 1152
rect 1798 1147 1804 1148
rect 1886 1152 1892 1153
rect 1886 1148 1887 1152
rect 1891 1148 1892 1152
rect 1886 1147 1892 1148
rect 1982 1152 1988 1153
rect 1982 1148 1983 1152
rect 1987 1148 1988 1152
rect 1982 1147 1988 1148
rect 2070 1152 2076 1153
rect 2070 1148 2071 1152
rect 2075 1148 2076 1152
rect 2070 1147 2076 1148
rect 1160 1131 1162 1147
rect 1208 1131 1210 1147
rect 1280 1131 1282 1147
rect 1352 1131 1354 1147
rect 1424 1131 1426 1147
rect 1488 1131 1490 1147
rect 1560 1131 1562 1147
rect 1632 1131 1634 1147
rect 1712 1131 1714 1147
rect 1800 1131 1802 1147
rect 1888 1131 1890 1147
rect 1984 1131 1986 1147
rect 2072 1131 2074 1147
rect 2120 1131 2122 1155
rect 1135 1130 1139 1131
rect 1135 1125 1139 1126
rect 1159 1130 1163 1131
rect 1159 1125 1163 1126
rect 1191 1130 1195 1131
rect 1191 1125 1195 1126
rect 1207 1130 1211 1131
rect 1207 1125 1211 1126
rect 1271 1130 1275 1131
rect 1271 1125 1275 1126
rect 1279 1130 1283 1131
rect 1279 1125 1283 1126
rect 1343 1130 1347 1131
rect 1343 1125 1347 1126
rect 1351 1130 1355 1131
rect 1351 1125 1355 1126
rect 1415 1130 1419 1131
rect 1415 1125 1419 1126
rect 1423 1130 1427 1131
rect 1423 1125 1427 1126
rect 1487 1130 1491 1131
rect 1487 1125 1491 1126
rect 1559 1130 1563 1131
rect 1559 1125 1563 1126
rect 1567 1130 1571 1131
rect 1567 1125 1571 1126
rect 1631 1130 1635 1131
rect 1631 1125 1635 1126
rect 1655 1130 1659 1131
rect 1655 1125 1659 1126
rect 1711 1130 1715 1131
rect 1711 1125 1715 1126
rect 1751 1130 1755 1131
rect 1751 1125 1755 1126
rect 1799 1130 1803 1131
rect 1799 1125 1803 1126
rect 1855 1130 1859 1131
rect 1855 1125 1859 1126
rect 1887 1130 1891 1131
rect 1887 1125 1891 1126
rect 1959 1130 1963 1131
rect 1959 1125 1963 1126
rect 1983 1130 1987 1131
rect 1983 1125 1987 1126
rect 2071 1130 2075 1131
rect 2071 1125 2075 1126
rect 2119 1130 2123 1131
rect 2119 1125 2123 1126
rect 110 1119 116 1120
rect 110 1115 111 1119
rect 115 1115 116 1119
rect 1094 1119 1100 1120
rect 110 1114 116 1115
rect 398 1116 404 1117
rect 112 1111 114 1114
rect 398 1112 399 1116
rect 403 1112 404 1116
rect 398 1111 404 1112
rect 438 1116 444 1117
rect 438 1112 439 1116
rect 443 1112 444 1116
rect 438 1111 444 1112
rect 478 1116 484 1117
rect 478 1112 479 1116
rect 483 1112 484 1116
rect 478 1111 484 1112
rect 526 1116 532 1117
rect 526 1112 527 1116
rect 531 1112 532 1116
rect 526 1111 532 1112
rect 574 1116 580 1117
rect 574 1112 575 1116
rect 579 1112 580 1116
rect 574 1111 580 1112
rect 622 1116 628 1117
rect 622 1112 623 1116
rect 627 1112 628 1116
rect 622 1111 628 1112
rect 670 1116 676 1117
rect 670 1112 671 1116
rect 675 1112 676 1116
rect 670 1111 676 1112
rect 718 1116 724 1117
rect 718 1112 719 1116
rect 723 1112 724 1116
rect 718 1111 724 1112
rect 774 1116 780 1117
rect 774 1112 775 1116
rect 779 1112 780 1116
rect 774 1111 780 1112
rect 830 1116 836 1117
rect 830 1112 831 1116
rect 835 1112 836 1116
rect 830 1111 836 1112
rect 886 1116 892 1117
rect 886 1112 887 1116
rect 891 1112 892 1116
rect 886 1111 892 1112
rect 942 1116 948 1117
rect 942 1112 943 1116
rect 947 1112 948 1116
rect 942 1111 948 1112
rect 1006 1116 1012 1117
rect 1006 1112 1007 1116
rect 1011 1112 1012 1116
rect 1006 1111 1012 1112
rect 1046 1116 1052 1117
rect 1046 1112 1047 1116
rect 1051 1112 1052 1116
rect 1094 1115 1095 1119
rect 1099 1115 1100 1119
rect 1094 1114 1100 1115
rect 1046 1111 1052 1112
rect 1096 1111 1098 1114
rect 111 1110 115 1111
rect 111 1105 115 1106
rect 159 1110 163 1111
rect 159 1105 163 1106
rect 199 1110 203 1111
rect 199 1105 203 1106
rect 255 1110 259 1111
rect 255 1105 259 1106
rect 319 1110 323 1111
rect 319 1105 323 1106
rect 399 1110 403 1111
rect 399 1105 403 1106
rect 439 1110 443 1111
rect 439 1105 443 1106
rect 479 1110 483 1111
rect 479 1105 483 1106
rect 527 1110 531 1111
rect 527 1105 531 1106
rect 559 1110 563 1111
rect 559 1105 563 1106
rect 575 1110 579 1111
rect 575 1105 579 1106
rect 623 1110 627 1111
rect 623 1105 627 1106
rect 639 1110 643 1111
rect 639 1105 643 1106
rect 671 1110 675 1111
rect 671 1105 675 1106
rect 711 1110 715 1111
rect 711 1105 715 1106
rect 719 1110 723 1111
rect 719 1105 723 1106
rect 775 1110 779 1111
rect 775 1105 779 1106
rect 783 1110 787 1111
rect 783 1105 787 1106
rect 831 1110 835 1111
rect 831 1105 835 1106
rect 855 1110 859 1111
rect 855 1105 859 1106
rect 887 1110 891 1111
rect 887 1105 891 1106
rect 927 1110 931 1111
rect 927 1105 931 1106
rect 943 1110 947 1111
rect 943 1105 947 1106
rect 999 1110 1003 1111
rect 999 1105 1003 1106
rect 1007 1110 1011 1111
rect 1007 1105 1011 1106
rect 1047 1110 1051 1111
rect 1047 1105 1051 1106
rect 1095 1110 1099 1111
rect 1095 1105 1099 1106
rect 1136 1105 1138 1125
rect 1192 1113 1194 1125
rect 1272 1113 1274 1125
rect 1344 1113 1346 1125
rect 1416 1113 1418 1125
rect 1488 1113 1490 1125
rect 1568 1113 1570 1125
rect 1656 1113 1658 1125
rect 1752 1113 1754 1125
rect 1856 1113 1858 1125
rect 1960 1113 1962 1125
rect 2072 1113 2074 1125
rect 1190 1112 1196 1113
rect 1190 1108 1191 1112
rect 1195 1108 1196 1112
rect 1190 1107 1196 1108
rect 1270 1112 1276 1113
rect 1270 1108 1271 1112
rect 1275 1108 1276 1112
rect 1270 1107 1276 1108
rect 1342 1112 1348 1113
rect 1342 1108 1343 1112
rect 1347 1108 1348 1112
rect 1342 1107 1348 1108
rect 1414 1112 1420 1113
rect 1414 1108 1415 1112
rect 1419 1108 1420 1112
rect 1414 1107 1420 1108
rect 1486 1112 1492 1113
rect 1486 1108 1487 1112
rect 1491 1108 1492 1112
rect 1486 1107 1492 1108
rect 1566 1112 1572 1113
rect 1566 1108 1567 1112
rect 1571 1108 1572 1112
rect 1566 1107 1572 1108
rect 1654 1112 1660 1113
rect 1654 1108 1655 1112
rect 1659 1108 1660 1112
rect 1654 1107 1660 1108
rect 1750 1112 1756 1113
rect 1750 1108 1751 1112
rect 1755 1108 1756 1112
rect 1750 1107 1756 1108
rect 1854 1112 1860 1113
rect 1854 1108 1855 1112
rect 1859 1108 1860 1112
rect 1854 1107 1860 1108
rect 1958 1112 1964 1113
rect 1958 1108 1959 1112
rect 1963 1108 1964 1112
rect 1958 1107 1964 1108
rect 2070 1112 2076 1113
rect 2070 1108 2071 1112
rect 2075 1108 2076 1112
rect 2070 1107 2076 1108
rect 2120 1105 2122 1125
rect 112 1102 114 1105
rect 158 1104 164 1105
rect 110 1101 116 1102
rect 110 1097 111 1101
rect 115 1097 116 1101
rect 158 1100 159 1104
rect 163 1100 164 1104
rect 158 1099 164 1100
rect 198 1104 204 1105
rect 198 1100 199 1104
rect 203 1100 204 1104
rect 198 1099 204 1100
rect 254 1104 260 1105
rect 254 1100 255 1104
rect 259 1100 260 1104
rect 254 1099 260 1100
rect 318 1104 324 1105
rect 318 1100 319 1104
rect 323 1100 324 1104
rect 318 1099 324 1100
rect 398 1104 404 1105
rect 398 1100 399 1104
rect 403 1100 404 1104
rect 398 1099 404 1100
rect 478 1104 484 1105
rect 478 1100 479 1104
rect 483 1100 484 1104
rect 478 1099 484 1100
rect 558 1104 564 1105
rect 558 1100 559 1104
rect 563 1100 564 1104
rect 558 1099 564 1100
rect 638 1104 644 1105
rect 638 1100 639 1104
rect 643 1100 644 1104
rect 638 1099 644 1100
rect 710 1104 716 1105
rect 710 1100 711 1104
rect 715 1100 716 1104
rect 710 1099 716 1100
rect 782 1104 788 1105
rect 782 1100 783 1104
rect 787 1100 788 1104
rect 782 1099 788 1100
rect 854 1104 860 1105
rect 854 1100 855 1104
rect 859 1100 860 1104
rect 854 1099 860 1100
rect 926 1104 932 1105
rect 926 1100 927 1104
rect 931 1100 932 1104
rect 926 1099 932 1100
rect 998 1104 1004 1105
rect 998 1100 999 1104
rect 1003 1100 1004 1104
rect 998 1099 1004 1100
rect 1046 1104 1052 1105
rect 1046 1100 1047 1104
rect 1051 1100 1052 1104
rect 1096 1102 1098 1105
rect 1134 1104 1140 1105
rect 1046 1099 1052 1100
rect 1094 1101 1100 1102
rect 110 1096 116 1097
rect 1094 1097 1095 1101
rect 1099 1097 1100 1101
rect 1134 1100 1135 1104
rect 1139 1100 1140 1104
rect 1134 1099 1140 1100
rect 2118 1104 2124 1105
rect 2118 1100 2119 1104
rect 2123 1100 2124 1104
rect 2118 1099 2124 1100
rect 1094 1096 1100 1097
rect 1134 1087 1140 1088
rect 110 1084 116 1085
rect 110 1080 111 1084
rect 115 1080 116 1084
rect 110 1079 116 1080
rect 1094 1084 1100 1085
rect 1094 1080 1095 1084
rect 1099 1080 1100 1084
rect 1134 1083 1135 1087
rect 1139 1083 1140 1087
rect 2118 1087 2124 1088
rect 1134 1082 1140 1083
rect 1190 1084 1196 1085
rect 1094 1079 1100 1080
rect 1136 1079 1138 1082
rect 1190 1080 1191 1084
rect 1195 1080 1196 1084
rect 1190 1079 1196 1080
rect 1270 1084 1276 1085
rect 1270 1080 1271 1084
rect 1275 1080 1276 1084
rect 1270 1079 1276 1080
rect 1342 1084 1348 1085
rect 1342 1080 1343 1084
rect 1347 1080 1348 1084
rect 1342 1079 1348 1080
rect 1414 1084 1420 1085
rect 1414 1080 1415 1084
rect 1419 1080 1420 1084
rect 1414 1079 1420 1080
rect 1486 1084 1492 1085
rect 1486 1080 1487 1084
rect 1491 1080 1492 1084
rect 1486 1079 1492 1080
rect 1566 1084 1572 1085
rect 1566 1080 1567 1084
rect 1571 1080 1572 1084
rect 1566 1079 1572 1080
rect 1654 1084 1660 1085
rect 1654 1080 1655 1084
rect 1659 1080 1660 1084
rect 1654 1079 1660 1080
rect 1750 1084 1756 1085
rect 1750 1080 1751 1084
rect 1755 1080 1756 1084
rect 1750 1079 1756 1080
rect 1854 1084 1860 1085
rect 1854 1080 1855 1084
rect 1859 1080 1860 1084
rect 1854 1079 1860 1080
rect 1958 1084 1964 1085
rect 1958 1080 1959 1084
rect 1963 1080 1964 1084
rect 1958 1079 1964 1080
rect 2070 1084 2076 1085
rect 2070 1080 2071 1084
rect 2075 1080 2076 1084
rect 2118 1083 2119 1087
rect 2123 1083 2124 1087
rect 2118 1082 2124 1083
rect 2070 1079 2076 1080
rect 2120 1079 2122 1082
rect 112 1055 114 1079
rect 158 1076 164 1077
rect 158 1072 159 1076
rect 163 1072 164 1076
rect 158 1071 164 1072
rect 198 1076 204 1077
rect 198 1072 199 1076
rect 203 1072 204 1076
rect 198 1071 204 1072
rect 254 1076 260 1077
rect 254 1072 255 1076
rect 259 1072 260 1076
rect 254 1071 260 1072
rect 318 1076 324 1077
rect 318 1072 319 1076
rect 323 1072 324 1076
rect 318 1071 324 1072
rect 398 1076 404 1077
rect 398 1072 399 1076
rect 403 1072 404 1076
rect 398 1071 404 1072
rect 478 1076 484 1077
rect 478 1072 479 1076
rect 483 1072 484 1076
rect 478 1071 484 1072
rect 558 1076 564 1077
rect 558 1072 559 1076
rect 563 1072 564 1076
rect 558 1071 564 1072
rect 638 1076 644 1077
rect 638 1072 639 1076
rect 643 1072 644 1076
rect 638 1071 644 1072
rect 710 1076 716 1077
rect 710 1072 711 1076
rect 715 1072 716 1076
rect 710 1071 716 1072
rect 782 1076 788 1077
rect 782 1072 783 1076
rect 787 1072 788 1076
rect 782 1071 788 1072
rect 854 1076 860 1077
rect 854 1072 855 1076
rect 859 1072 860 1076
rect 854 1071 860 1072
rect 926 1076 932 1077
rect 926 1072 927 1076
rect 931 1072 932 1076
rect 926 1071 932 1072
rect 998 1076 1004 1077
rect 998 1072 999 1076
rect 1003 1072 1004 1076
rect 998 1071 1004 1072
rect 1046 1076 1052 1077
rect 1046 1072 1047 1076
rect 1051 1072 1052 1076
rect 1046 1071 1052 1072
rect 160 1055 162 1071
rect 200 1055 202 1071
rect 256 1055 258 1071
rect 320 1055 322 1071
rect 400 1055 402 1071
rect 480 1055 482 1071
rect 560 1055 562 1071
rect 640 1055 642 1071
rect 712 1055 714 1071
rect 784 1055 786 1071
rect 856 1055 858 1071
rect 928 1055 930 1071
rect 1000 1055 1002 1071
rect 1048 1055 1050 1071
rect 1096 1055 1098 1079
rect 1135 1078 1139 1079
rect 1135 1073 1139 1074
rect 1159 1078 1163 1079
rect 1159 1073 1163 1074
rect 1191 1078 1195 1079
rect 1191 1073 1195 1074
rect 1199 1078 1203 1079
rect 1199 1073 1203 1074
rect 1247 1078 1251 1079
rect 1247 1073 1251 1074
rect 1271 1078 1275 1079
rect 1271 1073 1275 1074
rect 1303 1078 1307 1079
rect 1303 1073 1307 1074
rect 1343 1078 1347 1079
rect 1343 1073 1347 1074
rect 1351 1078 1355 1079
rect 1351 1073 1355 1074
rect 1399 1078 1403 1079
rect 1399 1073 1403 1074
rect 1415 1078 1419 1079
rect 1415 1073 1419 1074
rect 1455 1078 1459 1079
rect 1455 1073 1459 1074
rect 1487 1078 1491 1079
rect 1487 1073 1491 1074
rect 1511 1078 1515 1079
rect 1511 1073 1515 1074
rect 1567 1078 1571 1079
rect 1567 1073 1571 1074
rect 1583 1078 1587 1079
rect 1583 1073 1587 1074
rect 1655 1078 1659 1079
rect 1655 1073 1659 1074
rect 1663 1078 1667 1079
rect 1663 1073 1667 1074
rect 1751 1078 1755 1079
rect 1751 1073 1755 1074
rect 1759 1078 1763 1079
rect 1759 1073 1763 1074
rect 1855 1078 1859 1079
rect 1855 1073 1859 1074
rect 1863 1078 1867 1079
rect 1863 1073 1867 1074
rect 1959 1078 1963 1079
rect 1959 1073 1963 1074
rect 1967 1078 1971 1079
rect 1967 1073 1971 1074
rect 2071 1078 2075 1079
rect 2071 1073 2075 1074
rect 2119 1078 2123 1079
rect 2119 1073 2123 1074
rect 1136 1070 1138 1073
rect 1158 1072 1164 1073
rect 1134 1069 1140 1070
rect 1134 1065 1135 1069
rect 1139 1065 1140 1069
rect 1158 1068 1159 1072
rect 1163 1068 1164 1072
rect 1158 1067 1164 1068
rect 1198 1072 1204 1073
rect 1198 1068 1199 1072
rect 1203 1068 1204 1072
rect 1198 1067 1204 1068
rect 1246 1072 1252 1073
rect 1246 1068 1247 1072
rect 1251 1068 1252 1072
rect 1246 1067 1252 1068
rect 1302 1072 1308 1073
rect 1302 1068 1303 1072
rect 1307 1068 1308 1072
rect 1302 1067 1308 1068
rect 1350 1072 1356 1073
rect 1350 1068 1351 1072
rect 1355 1068 1356 1072
rect 1350 1067 1356 1068
rect 1398 1072 1404 1073
rect 1398 1068 1399 1072
rect 1403 1068 1404 1072
rect 1398 1067 1404 1068
rect 1454 1072 1460 1073
rect 1454 1068 1455 1072
rect 1459 1068 1460 1072
rect 1454 1067 1460 1068
rect 1510 1072 1516 1073
rect 1510 1068 1511 1072
rect 1515 1068 1516 1072
rect 1510 1067 1516 1068
rect 1582 1072 1588 1073
rect 1582 1068 1583 1072
rect 1587 1068 1588 1072
rect 1582 1067 1588 1068
rect 1662 1072 1668 1073
rect 1662 1068 1663 1072
rect 1667 1068 1668 1072
rect 1662 1067 1668 1068
rect 1758 1072 1764 1073
rect 1758 1068 1759 1072
rect 1763 1068 1764 1072
rect 1758 1067 1764 1068
rect 1862 1072 1868 1073
rect 1862 1068 1863 1072
rect 1867 1068 1868 1072
rect 1862 1067 1868 1068
rect 1966 1072 1972 1073
rect 1966 1068 1967 1072
rect 1971 1068 1972 1072
rect 1966 1067 1972 1068
rect 2070 1072 2076 1073
rect 2070 1068 2071 1072
rect 2075 1068 2076 1072
rect 2120 1070 2122 1073
rect 2070 1067 2076 1068
rect 2118 1069 2124 1070
rect 1134 1064 1140 1065
rect 2118 1065 2119 1069
rect 2123 1065 2124 1069
rect 2118 1064 2124 1065
rect 111 1054 115 1055
rect 111 1049 115 1050
rect 135 1054 139 1055
rect 135 1049 139 1050
rect 159 1054 163 1055
rect 159 1049 163 1050
rect 175 1054 179 1055
rect 175 1049 179 1050
rect 199 1054 203 1055
rect 199 1049 203 1050
rect 215 1054 219 1055
rect 215 1049 219 1050
rect 255 1054 259 1055
rect 255 1049 259 1050
rect 319 1054 323 1055
rect 319 1049 323 1050
rect 383 1054 387 1055
rect 383 1049 387 1050
rect 399 1054 403 1055
rect 399 1049 403 1050
rect 447 1054 451 1055
rect 447 1049 451 1050
rect 479 1054 483 1055
rect 479 1049 483 1050
rect 511 1054 515 1055
rect 511 1049 515 1050
rect 559 1054 563 1055
rect 559 1049 563 1050
rect 575 1054 579 1055
rect 575 1049 579 1050
rect 631 1054 635 1055
rect 631 1049 635 1050
rect 639 1054 643 1055
rect 639 1049 643 1050
rect 687 1054 691 1055
rect 687 1049 691 1050
rect 711 1054 715 1055
rect 711 1049 715 1050
rect 743 1054 747 1055
rect 743 1049 747 1050
rect 783 1054 787 1055
rect 783 1049 787 1050
rect 799 1054 803 1055
rect 799 1049 803 1050
rect 855 1054 859 1055
rect 855 1049 859 1050
rect 863 1054 867 1055
rect 863 1049 867 1050
rect 927 1054 931 1055
rect 927 1049 931 1050
rect 999 1054 1003 1055
rect 999 1049 1003 1050
rect 1047 1054 1051 1055
rect 1047 1049 1051 1050
rect 1095 1054 1099 1055
rect 1095 1049 1099 1050
rect 1134 1052 1140 1053
rect 112 1029 114 1049
rect 136 1037 138 1049
rect 176 1037 178 1049
rect 216 1037 218 1049
rect 256 1037 258 1049
rect 320 1037 322 1049
rect 384 1037 386 1049
rect 448 1037 450 1049
rect 512 1037 514 1049
rect 576 1037 578 1049
rect 632 1037 634 1049
rect 688 1037 690 1049
rect 744 1037 746 1049
rect 800 1037 802 1049
rect 864 1037 866 1049
rect 134 1036 140 1037
rect 134 1032 135 1036
rect 139 1032 140 1036
rect 134 1031 140 1032
rect 174 1036 180 1037
rect 174 1032 175 1036
rect 179 1032 180 1036
rect 174 1031 180 1032
rect 214 1036 220 1037
rect 214 1032 215 1036
rect 219 1032 220 1036
rect 214 1031 220 1032
rect 254 1036 260 1037
rect 254 1032 255 1036
rect 259 1032 260 1036
rect 254 1031 260 1032
rect 318 1036 324 1037
rect 318 1032 319 1036
rect 323 1032 324 1036
rect 318 1031 324 1032
rect 382 1036 388 1037
rect 382 1032 383 1036
rect 387 1032 388 1036
rect 382 1031 388 1032
rect 446 1036 452 1037
rect 446 1032 447 1036
rect 451 1032 452 1036
rect 446 1031 452 1032
rect 510 1036 516 1037
rect 510 1032 511 1036
rect 515 1032 516 1036
rect 510 1031 516 1032
rect 574 1036 580 1037
rect 574 1032 575 1036
rect 579 1032 580 1036
rect 574 1031 580 1032
rect 630 1036 636 1037
rect 630 1032 631 1036
rect 635 1032 636 1036
rect 630 1031 636 1032
rect 686 1036 692 1037
rect 686 1032 687 1036
rect 691 1032 692 1036
rect 686 1031 692 1032
rect 742 1036 748 1037
rect 742 1032 743 1036
rect 747 1032 748 1036
rect 742 1031 748 1032
rect 798 1036 804 1037
rect 798 1032 799 1036
rect 803 1032 804 1036
rect 798 1031 804 1032
rect 862 1036 868 1037
rect 862 1032 863 1036
rect 867 1032 868 1036
rect 862 1031 868 1032
rect 1096 1029 1098 1049
rect 1134 1048 1135 1052
rect 1139 1048 1140 1052
rect 1134 1047 1140 1048
rect 2118 1052 2124 1053
rect 2118 1048 2119 1052
rect 2123 1048 2124 1052
rect 2118 1047 2124 1048
rect 110 1028 116 1029
rect 110 1024 111 1028
rect 115 1024 116 1028
rect 110 1023 116 1024
rect 1094 1028 1100 1029
rect 1094 1024 1095 1028
rect 1099 1024 1100 1028
rect 1094 1023 1100 1024
rect 1136 1023 1138 1047
rect 1158 1044 1164 1045
rect 1158 1040 1159 1044
rect 1163 1040 1164 1044
rect 1158 1039 1164 1040
rect 1198 1044 1204 1045
rect 1198 1040 1199 1044
rect 1203 1040 1204 1044
rect 1198 1039 1204 1040
rect 1246 1044 1252 1045
rect 1246 1040 1247 1044
rect 1251 1040 1252 1044
rect 1246 1039 1252 1040
rect 1302 1044 1308 1045
rect 1302 1040 1303 1044
rect 1307 1040 1308 1044
rect 1302 1039 1308 1040
rect 1350 1044 1356 1045
rect 1350 1040 1351 1044
rect 1355 1040 1356 1044
rect 1350 1039 1356 1040
rect 1398 1044 1404 1045
rect 1398 1040 1399 1044
rect 1403 1040 1404 1044
rect 1398 1039 1404 1040
rect 1454 1044 1460 1045
rect 1454 1040 1455 1044
rect 1459 1040 1460 1044
rect 1454 1039 1460 1040
rect 1510 1044 1516 1045
rect 1510 1040 1511 1044
rect 1515 1040 1516 1044
rect 1510 1039 1516 1040
rect 1582 1044 1588 1045
rect 1582 1040 1583 1044
rect 1587 1040 1588 1044
rect 1582 1039 1588 1040
rect 1662 1044 1668 1045
rect 1662 1040 1663 1044
rect 1667 1040 1668 1044
rect 1662 1039 1668 1040
rect 1758 1044 1764 1045
rect 1758 1040 1759 1044
rect 1763 1040 1764 1044
rect 1758 1039 1764 1040
rect 1862 1044 1868 1045
rect 1862 1040 1863 1044
rect 1867 1040 1868 1044
rect 1862 1039 1868 1040
rect 1966 1044 1972 1045
rect 1966 1040 1967 1044
rect 1971 1040 1972 1044
rect 1966 1039 1972 1040
rect 2070 1044 2076 1045
rect 2070 1040 2071 1044
rect 2075 1040 2076 1044
rect 2070 1039 2076 1040
rect 1160 1023 1162 1039
rect 1200 1023 1202 1039
rect 1248 1023 1250 1039
rect 1304 1023 1306 1039
rect 1352 1023 1354 1039
rect 1400 1023 1402 1039
rect 1456 1023 1458 1039
rect 1512 1023 1514 1039
rect 1584 1023 1586 1039
rect 1664 1023 1666 1039
rect 1760 1023 1762 1039
rect 1864 1023 1866 1039
rect 1968 1023 1970 1039
rect 2072 1023 2074 1039
rect 2120 1023 2122 1047
rect 1135 1022 1139 1023
rect 1135 1017 1139 1018
rect 1159 1022 1163 1023
rect 1159 1017 1163 1018
rect 1199 1022 1203 1023
rect 1199 1017 1203 1018
rect 1239 1022 1243 1023
rect 1239 1017 1243 1018
rect 1247 1022 1251 1023
rect 1247 1017 1251 1018
rect 1295 1022 1299 1023
rect 1295 1017 1299 1018
rect 1303 1022 1307 1023
rect 1303 1017 1307 1018
rect 1351 1022 1355 1023
rect 1351 1017 1355 1018
rect 1399 1022 1403 1023
rect 1399 1017 1403 1018
rect 1407 1022 1411 1023
rect 1407 1017 1411 1018
rect 1455 1022 1459 1023
rect 1455 1017 1459 1018
rect 1463 1022 1467 1023
rect 1463 1017 1467 1018
rect 1511 1022 1515 1023
rect 1511 1017 1515 1018
rect 1519 1022 1523 1023
rect 1519 1017 1523 1018
rect 1575 1022 1579 1023
rect 1575 1017 1579 1018
rect 1583 1022 1587 1023
rect 1583 1017 1587 1018
rect 1639 1022 1643 1023
rect 1639 1017 1643 1018
rect 1663 1022 1667 1023
rect 1663 1017 1667 1018
rect 1711 1022 1715 1023
rect 1711 1017 1715 1018
rect 1759 1022 1763 1023
rect 1759 1017 1763 1018
rect 1791 1022 1795 1023
rect 1791 1017 1795 1018
rect 1863 1022 1867 1023
rect 1863 1017 1867 1018
rect 1879 1022 1883 1023
rect 1879 1017 1883 1018
rect 1967 1022 1971 1023
rect 1967 1017 1971 1018
rect 2063 1022 2067 1023
rect 2063 1017 2067 1018
rect 2071 1022 2075 1023
rect 2071 1017 2075 1018
rect 2119 1022 2123 1023
rect 2119 1017 2123 1018
rect 110 1011 116 1012
rect 110 1007 111 1011
rect 115 1007 116 1011
rect 1094 1011 1100 1012
rect 110 1006 116 1007
rect 134 1008 140 1009
rect 112 999 114 1006
rect 134 1004 135 1008
rect 139 1004 140 1008
rect 134 1003 140 1004
rect 174 1008 180 1009
rect 174 1004 175 1008
rect 179 1004 180 1008
rect 174 1003 180 1004
rect 214 1008 220 1009
rect 214 1004 215 1008
rect 219 1004 220 1008
rect 214 1003 220 1004
rect 254 1008 260 1009
rect 254 1004 255 1008
rect 259 1004 260 1008
rect 254 1003 260 1004
rect 318 1008 324 1009
rect 318 1004 319 1008
rect 323 1004 324 1008
rect 318 1003 324 1004
rect 382 1008 388 1009
rect 382 1004 383 1008
rect 387 1004 388 1008
rect 382 1003 388 1004
rect 446 1008 452 1009
rect 446 1004 447 1008
rect 451 1004 452 1008
rect 446 1003 452 1004
rect 510 1008 516 1009
rect 510 1004 511 1008
rect 515 1004 516 1008
rect 510 1003 516 1004
rect 574 1008 580 1009
rect 574 1004 575 1008
rect 579 1004 580 1008
rect 574 1003 580 1004
rect 630 1008 636 1009
rect 630 1004 631 1008
rect 635 1004 636 1008
rect 630 1003 636 1004
rect 686 1008 692 1009
rect 686 1004 687 1008
rect 691 1004 692 1008
rect 686 1003 692 1004
rect 742 1008 748 1009
rect 742 1004 743 1008
rect 747 1004 748 1008
rect 742 1003 748 1004
rect 798 1008 804 1009
rect 798 1004 799 1008
rect 803 1004 804 1008
rect 798 1003 804 1004
rect 862 1008 868 1009
rect 862 1004 863 1008
rect 867 1004 868 1008
rect 1094 1007 1095 1011
rect 1099 1007 1100 1011
rect 1094 1006 1100 1007
rect 862 1003 868 1004
rect 136 999 138 1003
rect 176 999 178 1003
rect 216 999 218 1003
rect 256 999 258 1003
rect 320 999 322 1003
rect 384 999 386 1003
rect 448 999 450 1003
rect 512 999 514 1003
rect 576 999 578 1003
rect 632 999 634 1003
rect 688 999 690 1003
rect 744 999 746 1003
rect 800 999 802 1003
rect 864 999 866 1003
rect 1096 999 1098 1006
rect 111 998 115 999
rect 111 993 115 994
rect 135 998 139 999
rect 135 993 139 994
rect 175 998 179 999
rect 175 993 179 994
rect 215 998 219 999
rect 215 993 219 994
rect 223 998 227 999
rect 223 993 227 994
rect 255 998 259 999
rect 255 993 259 994
rect 279 998 283 999
rect 279 993 283 994
rect 319 998 323 999
rect 319 993 323 994
rect 343 998 347 999
rect 343 993 347 994
rect 383 998 387 999
rect 383 993 387 994
rect 407 998 411 999
rect 407 993 411 994
rect 447 998 451 999
rect 447 993 451 994
rect 471 998 475 999
rect 471 993 475 994
rect 511 998 515 999
rect 511 993 515 994
rect 527 998 531 999
rect 527 993 531 994
rect 575 998 579 999
rect 575 993 579 994
rect 583 998 587 999
rect 583 993 587 994
rect 631 998 635 999
rect 631 993 635 994
rect 687 998 691 999
rect 687 993 691 994
rect 743 998 747 999
rect 743 993 747 994
rect 799 998 803 999
rect 799 993 803 994
rect 863 998 867 999
rect 863 993 867 994
rect 1095 998 1099 999
rect 1136 997 1138 1017
rect 1160 1005 1162 1017
rect 1200 1005 1202 1017
rect 1240 1005 1242 1017
rect 1296 1005 1298 1017
rect 1352 1005 1354 1017
rect 1408 1005 1410 1017
rect 1464 1005 1466 1017
rect 1520 1005 1522 1017
rect 1576 1005 1578 1017
rect 1640 1005 1642 1017
rect 1712 1005 1714 1017
rect 1792 1005 1794 1017
rect 1880 1005 1882 1017
rect 1968 1005 1970 1017
rect 2064 1005 2066 1017
rect 1158 1004 1164 1005
rect 1158 1000 1159 1004
rect 1163 1000 1164 1004
rect 1158 999 1164 1000
rect 1198 1004 1204 1005
rect 1198 1000 1199 1004
rect 1203 1000 1204 1004
rect 1198 999 1204 1000
rect 1238 1004 1244 1005
rect 1238 1000 1239 1004
rect 1243 1000 1244 1004
rect 1238 999 1244 1000
rect 1294 1004 1300 1005
rect 1294 1000 1295 1004
rect 1299 1000 1300 1004
rect 1294 999 1300 1000
rect 1350 1004 1356 1005
rect 1350 1000 1351 1004
rect 1355 1000 1356 1004
rect 1350 999 1356 1000
rect 1406 1004 1412 1005
rect 1406 1000 1407 1004
rect 1411 1000 1412 1004
rect 1406 999 1412 1000
rect 1462 1004 1468 1005
rect 1462 1000 1463 1004
rect 1467 1000 1468 1004
rect 1462 999 1468 1000
rect 1518 1004 1524 1005
rect 1518 1000 1519 1004
rect 1523 1000 1524 1004
rect 1518 999 1524 1000
rect 1574 1004 1580 1005
rect 1574 1000 1575 1004
rect 1579 1000 1580 1004
rect 1574 999 1580 1000
rect 1638 1004 1644 1005
rect 1638 1000 1639 1004
rect 1643 1000 1644 1004
rect 1638 999 1644 1000
rect 1710 1004 1716 1005
rect 1710 1000 1711 1004
rect 1715 1000 1716 1004
rect 1710 999 1716 1000
rect 1790 1004 1796 1005
rect 1790 1000 1791 1004
rect 1795 1000 1796 1004
rect 1790 999 1796 1000
rect 1878 1004 1884 1005
rect 1878 1000 1879 1004
rect 1883 1000 1884 1004
rect 1878 999 1884 1000
rect 1966 1004 1972 1005
rect 1966 1000 1967 1004
rect 1971 1000 1972 1004
rect 1966 999 1972 1000
rect 2062 1004 2068 1005
rect 2062 1000 2063 1004
rect 2067 1000 2068 1004
rect 2062 999 2068 1000
rect 2120 997 2122 1017
rect 1095 993 1099 994
rect 1134 996 1140 997
rect 112 990 114 993
rect 134 992 140 993
rect 110 989 116 990
rect 110 985 111 989
rect 115 985 116 989
rect 134 988 135 992
rect 139 988 140 992
rect 134 987 140 988
rect 174 992 180 993
rect 174 988 175 992
rect 179 988 180 992
rect 174 987 180 988
rect 222 992 228 993
rect 222 988 223 992
rect 227 988 228 992
rect 222 987 228 988
rect 278 992 284 993
rect 278 988 279 992
rect 283 988 284 992
rect 278 987 284 988
rect 342 992 348 993
rect 342 988 343 992
rect 347 988 348 992
rect 342 987 348 988
rect 406 992 412 993
rect 406 988 407 992
rect 411 988 412 992
rect 406 987 412 988
rect 470 992 476 993
rect 470 988 471 992
rect 475 988 476 992
rect 470 987 476 988
rect 526 992 532 993
rect 526 988 527 992
rect 531 988 532 992
rect 526 987 532 988
rect 582 992 588 993
rect 582 988 583 992
rect 587 988 588 992
rect 582 987 588 988
rect 630 992 636 993
rect 630 988 631 992
rect 635 988 636 992
rect 630 987 636 988
rect 686 992 692 993
rect 686 988 687 992
rect 691 988 692 992
rect 686 987 692 988
rect 742 992 748 993
rect 742 988 743 992
rect 747 988 748 992
rect 742 987 748 988
rect 798 992 804 993
rect 798 988 799 992
rect 803 988 804 992
rect 1096 990 1098 993
rect 1134 992 1135 996
rect 1139 992 1140 996
rect 1134 991 1140 992
rect 2118 996 2124 997
rect 2118 992 2119 996
rect 2123 992 2124 996
rect 2118 991 2124 992
rect 798 987 804 988
rect 1094 989 1100 990
rect 110 984 116 985
rect 1094 985 1095 989
rect 1099 985 1100 989
rect 1094 984 1100 985
rect 1134 979 1140 980
rect 1134 975 1135 979
rect 1139 975 1140 979
rect 2118 979 2124 980
rect 1134 974 1140 975
rect 1158 976 1164 977
rect 110 972 116 973
rect 110 968 111 972
rect 115 968 116 972
rect 110 967 116 968
rect 1094 972 1100 973
rect 1094 968 1095 972
rect 1099 968 1100 972
rect 1094 967 1100 968
rect 112 943 114 967
rect 134 964 140 965
rect 134 960 135 964
rect 139 960 140 964
rect 134 959 140 960
rect 174 964 180 965
rect 174 960 175 964
rect 179 960 180 964
rect 174 959 180 960
rect 222 964 228 965
rect 222 960 223 964
rect 227 960 228 964
rect 222 959 228 960
rect 278 964 284 965
rect 278 960 279 964
rect 283 960 284 964
rect 278 959 284 960
rect 342 964 348 965
rect 342 960 343 964
rect 347 960 348 964
rect 342 959 348 960
rect 406 964 412 965
rect 406 960 407 964
rect 411 960 412 964
rect 406 959 412 960
rect 470 964 476 965
rect 470 960 471 964
rect 475 960 476 964
rect 470 959 476 960
rect 526 964 532 965
rect 526 960 527 964
rect 531 960 532 964
rect 526 959 532 960
rect 582 964 588 965
rect 582 960 583 964
rect 587 960 588 964
rect 582 959 588 960
rect 630 964 636 965
rect 630 960 631 964
rect 635 960 636 964
rect 630 959 636 960
rect 686 964 692 965
rect 686 960 687 964
rect 691 960 692 964
rect 686 959 692 960
rect 742 964 748 965
rect 742 960 743 964
rect 747 960 748 964
rect 742 959 748 960
rect 798 964 804 965
rect 798 960 799 964
rect 803 960 804 964
rect 798 959 804 960
rect 136 943 138 959
rect 176 943 178 959
rect 224 943 226 959
rect 280 943 282 959
rect 344 943 346 959
rect 408 943 410 959
rect 472 943 474 959
rect 528 943 530 959
rect 584 943 586 959
rect 632 943 634 959
rect 688 943 690 959
rect 744 943 746 959
rect 800 943 802 959
rect 1096 943 1098 967
rect 1136 963 1138 974
rect 1158 972 1159 976
rect 1163 972 1164 976
rect 1158 971 1164 972
rect 1198 976 1204 977
rect 1198 972 1199 976
rect 1203 972 1204 976
rect 1198 971 1204 972
rect 1238 976 1244 977
rect 1238 972 1239 976
rect 1243 972 1244 976
rect 1238 971 1244 972
rect 1294 976 1300 977
rect 1294 972 1295 976
rect 1299 972 1300 976
rect 1294 971 1300 972
rect 1350 976 1356 977
rect 1350 972 1351 976
rect 1355 972 1356 976
rect 1350 971 1356 972
rect 1406 976 1412 977
rect 1406 972 1407 976
rect 1411 972 1412 976
rect 1406 971 1412 972
rect 1462 976 1468 977
rect 1462 972 1463 976
rect 1467 972 1468 976
rect 1462 971 1468 972
rect 1518 976 1524 977
rect 1518 972 1519 976
rect 1523 972 1524 976
rect 1518 971 1524 972
rect 1574 976 1580 977
rect 1574 972 1575 976
rect 1579 972 1580 976
rect 1574 971 1580 972
rect 1638 976 1644 977
rect 1638 972 1639 976
rect 1643 972 1644 976
rect 1638 971 1644 972
rect 1710 976 1716 977
rect 1710 972 1711 976
rect 1715 972 1716 976
rect 1710 971 1716 972
rect 1790 976 1796 977
rect 1790 972 1791 976
rect 1795 972 1796 976
rect 1790 971 1796 972
rect 1878 976 1884 977
rect 1878 972 1879 976
rect 1883 972 1884 976
rect 1878 971 1884 972
rect 1966 976 1972 977
rect 1966 972 1967 976
rect 1971 972 1972 976
rect 1966 971 1972 972
rect 2062 976 2068 977
rect 2062 972 2063 976
rect 2067 972 2068 976
rect 2118 975 2119 979
rect 2123 975 2124 979
rect 2118 974 2124 975
rect 2062 971 2068 972
rect 1160 963 1162 971
rect 1200 963 1202 971
rect 1240 963 1242 971
rect 1296 963 1298 971
rect 1352 963 1354 971
rect 1408 963 1410 971
rect 1464 963 1466 971
rect 1520 963 1522 971
rect 1576 963 1578 971
rect 1640 963 1642 971
rect 1712 963 1714 971
rect 1792 963 1794 971
rect 1880 963 1882 971
rect 1968 963 1970 971
rect 2064 963 2066 971
rect 2120 963 2122 974
rect 1135 962 1139 963
rect 1135 957 1139 958
rect 1159 962 1163 963
rect 1159 957 1163 958
rect 1199 962 1203 963
rect 1199 957 1203 958
rect 1207 962 1211 963
rect 1207 957 1211 958
rect 1239 962 1243 963
rect 1239 957 1243 958
rect 1287 962 1291 963
rect 1287 957 1291 958
rect 1295 962 1299 963
rect 1295 957 1299 958
rect 1351 962 1355 963
rect 1351 957 1355 958
rect 1375 962 1379 963
rect 1375 957 1379 958
rect 1407 962 1411 963
rect 1407 957 1411 958
rect 1455 962 1459 963
rect 1455 957 1459 958
rect 1463 962 1467 963
rect 1463 957 1467 958
rect 1519 962 1523 963
rect 1519 957 1523 958
rect 1535 962 1539 963
rect 1535 957 1539 958
rect 1575 962 1579 963
rect 1575 957 1579 958
rect 1615 962 1619 963
rect 1615 957 1619 958
rect 1639 962 1643 963
rect 1639 957 1643 958
rect 1687 962 1691 963
rect 1687 957 1691 958
rect 1711 962 1715 963
rect 1711 957 1715 958
rect 1751 962 1755 963
rect 1751 957 1755 958
rect 1791 962 1795 963
rect 1791 957 1795 958
rect 1815 962 1819 963
rect 1815 957 1819 958
rect 1879 962 1883 963
rect 1879 957 1883 958
rect 1951 962 1955 963
rect 1951 957 1955 958
rect 1967 962 1971 963
rect 1967 957 1971 958
rect 2023 962 2027 963
rect 2023 957 2027 958
rect 2063 962 2067 963
rect 2063 957 2067 958
rect 2071 962 2075 963
rect 2071 957 2075 958
rect 2119 962 2123 963
rect 2119 957 2123 958
rect 1136 954 1138 957
rect 1158 956 1164 957
rect 1134 953 1140 954
rect 1134 949 1135 953
rect 1139 949 1140 953
rect 1158 952 1159 956
rect 1163 952 1164 956
rect 1158 951 1164 952
rect 1206 956 1212 957
rect 1206 952 1207 956
rect 1211 952 1212 956
rect 1206 951 1212 952
rect 1286 956 1292 957
rect 1286 952 1287 956
rect 1291 952 1292 956
rect 1286 951 1292 952
rect 1374 956 1380 957
rect 1374 952 1375 956
rect 1379 952 1380 956
rect 1374 951 1380 952
rect 1454 956 1460 957
rect 1454 952 1455 956
rect 1459 952 1460 956
rect 1454 951 1460 952
rect 1534 956 1540 957
rect 1534 952 1535 956
rect 1539 952 1540 956
rect 1534 951 1540 952
rect 1614 956 1620 957
rect 1614 952 1615 956
rect 1619 952 1620 956
rect 1614 951 1620 952
rect 1686 956 1692 957
rect 1686 952 1687 956
rect 1691 952 1692 956
rect 1686 951 1692 952
rect 1750 956 1756 957
rect 1750 952 1751 956
rect 1755 952 1756 956
rect 1750 951 1756 952
rect 1814 956 1820 957
rect 1814 952 1815 956
rect 1819 952 1820 956
rect 1814 951 1820 952
rect 1878 956 1884 957
rect 1878 952 1879 956
rect 1883 952 1884 956
rect 1878 951 1884 952
rect 1950 956 1956 957
rect 1950 952 1951 956
rect 1955 952 1956 956
rect 1950 951 1956 952
rect 2022 956 2028 957
rect 2022 952 2023 956
rect 2027 952 2028 956
rect 2022 951 2028 952
rect 2070 956 2076 957
rect 2070 952 2071 956
rect 2075 952 2076 956
rect 2120 954 2122 957
rect 2070 951 2076 952
rect 2118 953 2124 954
rect 1134 948 1140 949
rect 2118 949 2119 953
rect 2123 949 2124 953
rect 2118 948 2124 949
rect 111 942 115 943
rect 111 937 115 938
rect 135 942 139 943
rect 135 937 139 938
rect 175 942 179 943
rect 175 937 179 938
rect 223 942 227 943
rect 223 937 227 938
rect 263 942 267 943
rect 263 937 267 938
rect 279 942 283 943
rect 279 937 283 938
rect 303 942 307 943
rect 303 937 307 938
rect 343 942 347 943
rect 343 937 347 938
rect 351 942 355 943
rect 351 937 355 938
rect 399 942 403 943
rect 399 937 403 938
rect 407 942 411 943
rect 407 937 411 938
rect 455 942 459 943
rect 455 937 459 938
rect 471 942 475 943
rect 471 937 475 938
rect 511 942 515 943
rect 511 937 515 938
rect 527 942 531 943
rect 527 937 531 938
rect 567 942 571 943
rect 567 937 571 938
rect 583 942 587 943
rect 583 937 587 938
rect 623 942 627 943
rect 623 937 627 938
rect 631 942 635 943
rect 631 937 635 938
rect 687 942 691 943
rect 687 937 691 938
rect 743 942 747 943
rect 743 937 747 938
rect 751 942 755 943
rect 751 937 755 938
rect 799 942 803 943
rect 799 937 803 938
rect 815 942 819 943
rect 815 937 819 938
rect 879 942 883 943
rect 879 937 883 938
rect 943 942 947 943
rect 943 937 947 938
rect 1007 942 1011 943
rect 1007 937 1011 938
rect 1047 942 1051 943
rect 1047 937 1051 938
rect 1095 942 1099 943
rect 1095 937 1099 938
rect 112 917 114 937
rect 264 925 266 937
rect 304 925 306 937
rect 352 925 354 937
rect 400 925 402 937
rect 456 925 458 937
rect 512 925 514 937
rect 568 925 570 937
rect 624 925 626 937
rect 688 925 690 937
rect 752 925 754 937
rect 816 925 818 937
rect 880 925 882 937
rect 944 925 946 937
rect 1008 925 1010 937
rect 1048 925 1050 937
rect 262 924 268 925
rect 262 920 263 924
rect 267 920 268 924
rect 262 919 268 920
rect 302 924 308 925
rect 302 920 303 924
rect 307 920 308 924
rect 302 919 308 920
rect 350 924 356 925
rect 350 920 351 924
rect 355 920 356 924
rect 350 919 356 920
rect 398 924 404 925
rect 398 920 399 924
rect 403 920 404 924
rect 398 919 404 920
rect 454 924 460 925
rect 454 920 455 924
rect 459 920 460 924
rect 454 919 460 920
rect 510 924 516 925
rect 510 920 511 924
rect 515 920 516 924
rect 510 919 516 920
rect 566 924 572 925
rect 566 920 567 924
rect 571 920 572 924
rect 566 919 572 920
rect 622 924 628 925
rect 622 920 623 924
rect 627 920 628 924
rect 622 919 628 920
rect 686 924 692 925
rect 686 920 687 924
rect 691 920 692 924
rect 686 919 692 920
rect 750 924 756 925
rect 750 920 751 924
rect 755 920 756 924
rect 750 919 756 920
rect 814 924 820 925
rect 814 920 815 924
rect 819 920 820 924
rect 814 919 820 920
rect 878 924 884 925
rect 878 920 879 924
rect 883 920 884 924
rect 878 919 884 920
rect 942 924 948 925
rect 942 920 943 924
rect 947 920 948 924
rect 942 919 948 920
rect 1006 924 1012 925
rect 1006 920 1007 924
rect 1011 920 1012 924
rect 1006 919 1012 920
rect 1046 924 1052 925
rect 1046 920 1047 924
rect 1051 920 1052 924
rect 1046 919 1052 920
rect 1096 917 1098 937
rect 1134 936 1140 937
rect 1134 932 1135 936
rect 1139 932 1140 936
rect 1134 931 1140 932
rect 2118 936 2124 937
rect 2118 932 2119 936
rect 2123 932 2124 936
rect 2118 931 2124 932
rect 110 916 116 917
rect 110 912 111 916
rect 115 912 116 916
rect 110 911 116 912
rect 1094 916 1100 917
rect 1094 912 1095 916
rect 1099 912 1100 916
rect 1094 911 1100 912
rect 1136 911 1138 931
rect 1158 928 1164 929
rect 1158 924 1159 928
rect 1163 924 1164 928
rect 1158 923 1164 924
rect 1206 928 1212 929
rect 1206 924 1207 928
rect 1211 924 1212 928
rect 1206 923 1212 924
rect 1286 928 1292 929
rect 1286 924 1287 928
rect 1291 924 1292 928
rect 1286 923 1292 924
rect 1374 928 1380 929
rect 1374 924 1375 928
rect 1379 924 1380 928
rect 1374 923 1380 924
rect 1454 928 1460 929
rect 1454 924 1455 928
rect 1459 924 1460 928
rect 1454 923 1460 924
rect 1534 928 1540 929
rect 1534 924 1535 928
rect 1539 924 1540 928
rect 1534 923 1540 924
rect 1614 928 1620 929
rect 1614 924 1615 928
rect 1619 924 1620 928
rect 1614 923 1620 924
rect 1686 928 1692 929
rect 1686 924 1687 928
rect 1691 924 1692 928
rect 1686 923 1692 924
rect 1750 928 1756 929
rect 1750 924 1751 928
rect 1755 924 1756 928
rect 1750 923 1756 924
rect 1814 928 1820 929
rect 1814 924 1815 928
rect 1819 924 1820 928
rect 1814 923 1820 924
rect 1878 928 1884 929
rect 1878 924 1879 928
rect 1883 924 1884 928
rect 1878 923 1884 924
rect 1950 928 1956 929
rect 1950 924 1951 928
rect 1955 924 1956 928
rect 1950 923 1956 924
rect 2022 928 2028 929
rect 2022 924 2023 928
rect 2027 924 2028 928
rect 2022 923 2028 924
rect 2070 928 2076 929
rect 2070 924 2071 928
rect 2075 924 2076 928
rect 2070 923 2076 924
rect 1160 911 1162 923
rect 1208 911 1210 923
rect 1288 911 1290 923
rect 1376 911 1378 923
rect 1456 911 1458 923
rect 1536 911 1538 923
rect 1616 911 1618 923
rect 1688 911 1690 923
rect 1752 911 1754 923
rect 1816 911 1818 923
rect 1880 911 1882 923
rect 1952 911 1954 923
rect 2024 911 2026 923
rect 2072 911 2074 923
rect 2120 911 2122 931
rect 1135 910 1139 911
rect 1135 905 1139 906
rect 1159 910 1163 911
rect 1159 905 1163 906
rect 1207 910 1211 911
rect 1207 905 1211 906
rect 1239 910 1243 911
rect 1239 905 1243 906
rect 1287 910 1291 911
rect 1287 905 1291 906
rect 1319 910 1323 911
rect 1319 905 1323 906
rect 1375 910 1379 911
rect 1375 905 1379 906
rect 1407 910 1411 911
rect 1407 905 1411 906
rect 1455 910 1459 911
rect 1455 905 1459 906
rect 1495 910 1499 911
rect 1495 905 1499 906
rect 1535 910 1539 911
rect 1535 905 1539 906
rect 1583 910 1587 911
rect 1583 905 1587 906
rect 1615 910 1619 911
rect 1615 905 1619 906
rect 1663 910 1667 911
rect 1663 905 1667 906
rect 1687 910 1691 911
rect 1687 905 1691 906
rect 1743 910 1747 911
rect 1743 905 1747 906
rect 1751 910 1755 911
rect 1751 905 1755 906
rect 1815 910 1819 911
rect 1815 905 1819 906
rect 1879 910 1883 911
rect 1879 905 1883 906
rect 1887 910 1891 911
rect 1887 905 1891 906
rect 1951 910 1955 911
rect 1951 905 1955 906
rect 2023 910 2027 911
rect 2023 905 2027 906
rect 2071 910 2075 911
rect 2071 905 2075 906
rect 2119 910 2123 911
rect 2119 905 2123 906
rect 110 899 116 900
rect 110 895 111 899
rect 115 895 116 899
rect 1094 899 1100 900
rect 110 894 116 895
rect 262 896 268 897
rect 112 887 114 894
rect 262 892 263 896
rect 267 892 268 896
rect 262 891 268 892
rect 302 896 308 897
rect 302 892 303 896
rect 307 892 308 896
rect 302 891 308 892
rect 350 896 356 897
rect 350 892 351 896
rect 355 892 356 896
rect 350 891 356 892
rect 398 896 404 897
rect 398 892 399 896
rect 403 892 404 896
rect 398 891 404 892
rect 454 896 460 897
rect 454 892 455 896
rect 459 892 460 896
rect 454 891 460 892
rect 510 896 516 897
rect 510 892 511 896
rect 515 892 516 896
rect 510 891 516 892
rect 566 896 572 897
rect 566 892 567 896
rect 571 892 572 896
rect 566 891 572 892
rect 622 896 628 897
rect 622 892 623 896
rect 627 892 628 896
rect 622 891 628 892
rect 686 896 692 897
rect 686 892 687 896
rect 691 892 692 896
rect 686 891 692 892
rect 750 896 756 897
rect 750 892 751 896
rect 755 892 756 896
rect 750 891 756 892
rect 814 896 820 897
rect 814 892 815 896
rect 819 892 820 896
rect 814 891 820 892
rect 878 896 884 897
rect 878 892 879 896
rect 883 892 884 896
rect 878 891 884 892
rect 942 896 948 897
rect 942 892 943 896
rect 947 892 948 896
rect 942 891 948 892
rect 1006 896 1012 897
rect 1006 892 1007 896
rect 1011 892 1012 896
rect 1006 891 1012 892
rect 1046 896 1052 897
rect 1046 892 1047 896
rect 1051 892 1052 896
rect 1094 895 1095 899
rect 1099 895 1100 899
rect 1094 894 1100 895
rect 1046 891 1052 892
rect 264 887 266 891
rect 304 887 306 891
rect 352 887 354 891
rect 400 887 402 891
rect 456 887 458 891
rect 512 887 514 891
rect 568 887 570 891
rect 624 887 626 891
rect 688 887 690 891
rect 752 887 754 891
rect 816 887 818 891
rect 880 887 882 891
rect 944 887 946 891
rect 1008 887 1010 891
rect 1048 887 1050 891
rect 1096 887 1098 894
rect 111 886 115 887
rect 111 881 115 882
rect 263 886 267 887
rect 263 881 267 882
rect 303 886 307 887
rect 303 881 307 882
rect 351 886 355 887
rect 351 881 355 882
rect 399 886 403 887
rect 399 881 403 882
rect 415 886 419 887
rect 415 881 419 882
rect 455 886 459 887
rect 455 881 459 882
rect 479 886 483 887
rect 479 881 483 882
rect 511 886 515 887
rect 511 881 515 882
rect 551 886 555 887
rect 551 881 555 882
rect 567 886 571 887
rect 567 881 571 882
rect 623 886 627 887
rect 623 881 627 882
rect 687 886 691 887
rect 687 881 691 882
rect 695 886 699 887
rect 695 881 699 882
rect 751 886 755 887
rect 751 881 755 882
rect 767 886 771 887
rect 767 881 771 882
rect 815 886 819 887
rect 815 881 819 882
rect 831 886 835 887
rect 831 881 835 882
rect 879 886 883 887
rect 879 881 883 882
rect 887 886 891 887
rect 887 881 891 882
rect 943 886 947 887
rect 943 881 947 882
rect 1007 886 1011 887
rect 1007 881 1011 882
rect 1047 886 1051 887
rect 1047 881 1051 882
rect 1095 886 1099 887
rect 1136 885 1138 905
rect 1240 893 1242 905
rect 1320 893 1322 905
rect 1408 893 1410 905
rect 1496 893 1498 905
rect 1584 893 1586 905
rect 1664 893 1666 905
rect 1744 893 1746 905
rect 1816 893 1818 905
rect 1888 893 1890 905
rect 1952 893 1954 905
rect 2024 893 2026 905
rect 2072 893 2074 905
rect 1238 892 1244 893
rect 1238 888 1239 892
rect 1243 888 1244 892
rect 1238 887 1244 888
rect 1318 892 1324 893
rect 1318 888 1319 892
rect 1323 888 1324 892
rect 1318 887 1324 888
rect 1406 892 1412 893
rect 1406 888 1407 892
rect 1411 888 1412 892
rect 1406 887 1412 888
rect 1494 892 1500 893
rect 1494 888 1495 892
rect 1499 888 1500 892
rect 1494 887 1500 888
rect 1582 892 1588 893
rect 1582 888 1583 892
rect 1587 888 1588 892
rect 1582 887 1588 888
rect 1662 892 1668 893
rect 1662 888 1663 892
rect 1667 888 1668 892
rect 1662 887 1668 888
rect 1742 892 1748 893
rect 1742 888 1743 892
rect 1747 888 1748 892
rect 1742 887 1748 888
rect 1814 892 1820 893
rect 1814 888 1815 892
rect 1819 888 1820 892
rect 1814 887 1820 888
rect 1886 892 1892 893
rect 1886 888 1887 892
rect 1891 888 1892 892
rect 1886 887 1892 888
rect 1950 892 1956 893
rect 1950 888 1951 892
rect 1955 888 1956 892
rect 1950 887 1956 888
rect 2022 892 2028 893
rect 2022 888 2023 892
rect 2027 888 2028 892
rect 2022 887 2028 888
rect 2070 892 2076 893
rect 2070 888 2071 892
rect 2075 888 2076 892
rect 2070 887 2076 888
rect 2120 885 2122 905
rect 1095 881 1099 882
rect 1134 884 1140 885
rect 112 878 114 881
rect 302 880 308 881
rect 110 877 116 878
rect 110 873 111 877
rect 115 873 116 877
rect 302 876 303 880
rect 307 876 308 880
rect 302 875 308 876
rect 350 880 356 881
rect 350 876 351 880
rect 355 876 356 880
rect 350 875 356 876
rect 414 880 420 881
rect 414 876 415 880
rect 419 876 420 880
rect 414 875 420 876
rect 478 880 484 881
rect 478 876 479 880
rect 483 876 484 880
rect 478 875 484 876
rect 550 880 556 881
rect 550 876 551 880
rect 555 876 556 880
rect 550 875 556 876
rect 622 880 628 881
rect 622 876 623 880
rect 627 876 628 880
rect 622 875 628 876
rect 694 880 700 881
rect 694 876 695 880
rect 699 876 700 880
rect 694 875 700 876
rect 766 880 772 881
rect 766 876 767 880
rect 771 876 772 880
rect 766 875 772 876
rect 830 880 836 881
rect 830 876 831 880
rect 835 876 836 880
rect 830 875 836 876
rect 886 880 892 881
rect 886 876 887 880
rect 891 876 892 880
rect 886 875 892 876
rect 942 880 948 881
rect 942 876 943 880
rect 947 876 948 880
rect 942 875 948 876
rect 1006 880 1012 881
rect 1006 876 1007 880
rect 1011 876 1012 880
rect 1006 875 1012 876
rect 1046 880 1052 881
rect 1046 876 1047 880
rect 1051 876 1052 880
rect 1096 878 1098 881
rect 1134 880 1135 884
rect 1139 880 1140 884
rect 1134 879 1140 880
rect 2118 884 2124 885
rect 2118 880 2119 884
rect 2123 880 2124 884
rect 2118 879 2124 880
rect 1046 875 1052 876
rect 1094 877 1100 878
rect 110 872 116 873
rect 1094 873 1095 877
rect 1099 873 1100 877
rect 1094 872 1100 873
rect 1134 867 1140 868
rect 1134 863 1135 867
rect 1139 863 1140 867
rect 2118 867 2124 868
rect 1134 862 1140 863
rect 1238 864 1244 865
rect 110 860 116 861
rect 110 856 111 860
rect 115 856 116 860
rect 110 855 116 856
rect 1094 860 1100 861
rect 1094 856 1095 860
rect 1099 856 1100 860
rect 1136 859 1138 862
rect 1238 860 1239 864
rect 1243 860 1244 864
rect 1238 859 1244 860
rect 1318 864 1324 865
rect 1318 860 1319 864
rect 1323 860 1324 864
rect 1318 859 1324 860
rect 1406 864 1412 865
rect 1406 860 1407 864
rect 1411 860 1412 864
rect 1406 859 1412 860
rect 1494 864 1500 865
rect 1494 860 1495 864
rect 1499 860 1500 864
rect 1494 859 1500 860
rect 1582 864 1588 865
rect 1582 860 1583 864
rect 1587 860 1588 864
rect 1582 859 1588 860
rect 1662 864 1668 865
rect 1662 860 1663 864
rect 1667 860 1668 864
rect 1662 859 1668 860
rect 1742 864 1748 865
rect 1742 860 1743 864
rect 1747 860 1748 864
rect 1742 859 1748 860
rect 1814 864 1820 865
rect 1814 860 1815 864
rect 1819 860 1820 864
rect 1814 859 1820 860
rect 1886 864 1892 865
rect 1886 860 1887 864
rect 1891 860 1892 864
rect 1886 859 1892 860
rect 1950 864 1956 865
rect 1950 860 1951 864
rect 1955 860 1956 864
rect 1950 859 1956 860
rect 2022 864 2028 865
rect 2022 860 2023 864
rect 2027 860 2028 864
rect 2022 859 2028 860
rect 2070 864 2076 865
rect 2070 860 2071 864
rect 2075 860 2076 864
rect 2118 863 2119 867
rect 2123 863 2124 867
rect 2118 862 2124 863
rect 2070 859 2076 860
rect 2120 859 2122 862
rect 1094 855 1100 856
rect 1135 858 1139 859
rect 112 835 114 855
rect 302 852 308 853
rect 302 848 303 852
rect 307 848 308 852
rect 302 847 308 848
rect 350 852 356 853
rect 350 848 351 852
rect 355 848 356 852
rect 350 847 356 848
rect 414 852 420 853
rect 414 848 415 852
rect 419 848 420 852
rect 414 847 420 848
rect 478 852 484 853
rect 478 848 479 852
rect 483 848 484 852
rect 478 847 484 848
rect 550 852 556 853
rect 550 848 551 852
rect 555 848 556 852
rect 550 847 556 848
rect 622 852 628 853
rect 622 848 623 852
rect 627 848 628 852
rect 622 847 628 848
rect 694 852 700 853
rect 694 848 695 852
rect 699 848 700 852
rect 694 847 700 848
rect 766 852 772 853
rect 766 848 767 852
rect 771 848 772 852
rect 766 847 772 848
rect 830 852 836 853
rect 830 848 831 852
rect 835 848 836 852
rect 830 847 836 848
rect 886 852 892 853
rect 886 848 887 852
rect 891 848 892 852
rect 886 847 892 848
rect 942 852 948 853
rect 942 848 943 852
rect 947 848 948 852
rect 942 847 948 848
rect 1006 852 1012 853
rect 1006 848 1007 852
rect 1011 848 1012 852
rect 1006 847 1012 848
rect 1046 852 1052 853
rect 1046 848 1047 852
rect 1051 848 1052 852
rect 1046 847 1052 848
rect 304 835 306 847
rect 352 835 354 847
rect 416 835 418 847
rect 480 835 482 847
rect 552 835 554 847
rect 624 835 626 847
rect 696 835 698 847
rect 768 835 770 847
rect 832 835 834 847
rect 888 835 890 847
rect 944 835 946 847
rect 1008 835 1010 847
rect 1048 835 1050 847
rect 1096 835 1098 855
rect 1135 853 1139 854
rect 1159 858 1163 859
rect 1159 853 1163 854
rect 1239 858 1243 859
rect 1239 853 1243 854
rect 1247 858 1251 859
rect 1247 853 1251 854
rect 1319 858 1323 859
rect 1319 853 1323 854
rect 1359 858 1363 859
rect 1359 853 1363 854
rect 1407 858 1411 859
rect 1407 853 1411 854
rect 1455 858 1459 859
rect 1455 853 1459 854
rect 1495 858 1499 859
rect 1495 853 1499 854
rect 1543 858 1547 859
rect 1543 853 1547 854
rect 1583 858 1587 859
rect 1583 853 1587 854
rect 1631 858 1635 859
rect 1631 853 1635 854
rect 1663 858 1667 859
rect 1663 853 1667 854
rect 1711 858 1715 859
rect 1711 853 1715 854
rect 1743 858 1747 859
rect 1743 853 1747 854
rect 1783 858 1787 859
rect 1783 853 1787 854
rect 1815 858 1819 859
rect 1815 853 1819 854
rect 1855 858 1859 859
rect 1855 853 1859 854
rect 1887 858 1891 859
rect 1887 853 1891 854
rect 1935 858 1939 859
rect 1935 853 1939 854
rect 1951 858 1955 859
rect 1951 853 1955 854
rect 2015 858 2019 859
rect 2015 853 2019 854
rect 2023 858 2027 859
rect 2023 853 2027 854
rect 2071 858 2075 859
rect 2071 853 2075 854
rect 2119 858 2123 859
rect 2119 853 2123 854
rect 1136 850 1138 853
rect 1158 852 1164 853
rect 1134 849 1140 850
rect 1134 845 1135 849
rect 1139 845 1140 849
rect 1158 848 1159 852
rect 1163 848 1164 852
rect 1158 847 1164 848
rect 1246 852 1252 853
rect 1246 848 1247 852
rect 1251 848 1252 852
rect 1246 847 1252 848
rect 1358 852 1364 853
rect 1358 848 1359 852
rect 1363 848 1364 852
rect 1358 847 1364 848
rect 1454 852 1460 853
rect 1454 848 1455 852
rect 1459 848 1460 852
rect 1454 847 1460 848
rect 1542 852 1548 853
rect 1542 848 1543 852
rect 1547 848 1548 852
rect 1542 847 1548 848
rect 1630 852 1636 853
rect 1630 848 1631 852
rect 1635 848 1636 852
rect 1630 847 1636 848
rect 1710 852 1716 853
rect 1710 848 1711 852
rect 1715 848 1716 852
rect 1710 847 1716 848
rect 1782 852 1788 853
rect 1782 848 1783 852
rect 1787 848 1788 852
rect 1782 847 1788 848
rect 1854 852 1860 853
rect 1854 848 1855 852
rect 1859 848 1860 852
rect 1854 847 1860 848
rect 1934 852 1940 853
rect 1934 848 1935 852
rect 1939 848 1940 852
rect 1934 847 1940 848
rect 2014 852 2020 853
rect 2014 848 2015 852
rect 2019 848 2020 852
rect 2014 847 2020 848
rect 2070 852 2076 853
rect 2070 848 2071 852
rect 2075 848 2076 852
rect 2120 850 2122 853
rect 2070 847 2076 848
rect 2118 849 2124 850
rect 1134 844 1140 845
rect 2118 845 2119 849
rect 2123 845 2124 849
rect 2118 844 2124 845
rect 111 834 115 835
rect 111 829 115 830
rect 279 834 283 835
rect 279 829 283 830
rect 303 834 307 835
rect 303 829 307 830
rect 343 834 347 835
rect 343 829 347 830
rect 351 834 355 835
rect 351 829 355 830
rect 415 834 419 835
rect 415 829 419 830
rect 479 834 483 835
rect 479 829 483 830
rect 487 834 491 835
rect 487 829 491 830
rect 551 834 555 835
rect 551 829 555 830
rect 567 834 571 835
rect 567 829 571 830
rect 623 834 627 835
rect 623 829 627 830
rect 647 834 651 835
rect 647 829 651 830
rect 695 834 699 835
rect 695 829 699 830
rect 727 834 731 835
rect 727 829 731 830
rect 767 834 771 835
rect 767 829 771 830
rect 799 834 803 835
rect 799 829 803 830
rect 831 834 835 835
rect 831 829 835 830
rect 863 834 867 835
rect 863 829 867 830
rect 887 834 891 835
rect 887 829 891 830
rect 927 834 931 835
rect 927 829 931 830
rect 943 834 947 835
rect 943 829 947 830
rect 999 834 1003 835
rect 999 829 1003 830
rect 1007 834 1011 835
rect 1007 829 1011 830
rect 1047 834 1051 835
rect 1047 829 1051 830
rect 1095 834 1099 835
rect 1095 829 1099 830
rect 1134 832 1140 833
rect 112 809 114 829
rect 280 817 282 829
rect 344 817 346 829
rect 416 817 418 829
rect 488 817 490 829
rect 568 817 570 829
rect 648 817 650 829
rect 728 817 730 829
rect 800 817 802 829
rect 864 817 866 829
rect 928 817 930 829
rect 1000 817 1002 829
rect 1048 817 1050 829
rect 278 816 284 817
rect 278 812 279 816
rect 283 812 284 816
rect 278 811 284 812
rect 342 816 348 817
rect 342 812 343 816
rect 347 812 348 816
rect 342 811 348 812
rect 414 816 420 817
rect 414 812 415 816
rect 419 812 420 816
rect 414 811 420 812
rect 486 816 492 817
rect 486 812 487 816
rect 491 812 492 816
rect 486 811 492 812
rect 566 816 572 817
rect 566 812 567 816
rect 571 812 572 816
rect 566 811 572 812
rect 646 816 652 817
rect 646 812 647 816
rect 651 812 652 816
rect 646 811 652 812
rect 726 816 732 817
rect 726 812 727 816
rect 731 812 732 816
rect 726 811 732 812
rect 798 816 804 817
rect 798 812 799 816
rect 803 812 804 816
rect 798 811 804 812
rect 862 816 868 817
rect 862 812 863 816
rect 867 812 868 816
rect 862 811 868 812
rect 926 816 932 817
rect 926 812 927 816
rect 931 812 932 816
rect 926 811 932 812
rect 998 816 1004 817
rect 998 812 999 816
rect 1003 812 1004 816
rect 998 811 1004 812
rect 1046 816 1052 817
rect 1046 812 1047 816
rect 1051 812 1052 816
rect 1046 811 1052 812
rect 1096 809 1098 829
rect 1134 828 1135 832
rect 1139 828 1140 832
rect 1134 827 1140 828
rect 2118 832 2124 833
rect 2118 828 2119 832
rect 2123 828 2124 832
rect 2118 827 2124 828
rect 110 808 116 809
rect 110 804 111 808
rect 115 804 116 808
rect 110 803 116 804
rect 1094 808 1100 809
rect 1094 804 1095 808
rect 1099 804 1100 808
rect 1136 807 1138 827
rect 1158 824 1164 825
rect 1158 820 1159 824
rect 1163 820 1164 824
rect 1158 819 1164 820
rect 1246 824 1252 825
rect 1246 820 1247 824
rect 1251 820 1252 824
rect 1246 819 1252 820
rect 1358 824 1364 825
rect 1358 820 1359 824
rect 1363 820 1364 824
rect 1358 819 1364 820
rect 1454 824 1460 825
rect 1454 820 1455 824
rect 1459 820 1460 824
rect 1454 819 1460 820
rect 1542 824 1548 825
rect 1542 820 1543 824
rect 1547 820 1548 824
rect 1542 819 1548 820
rect 1630 824 1636 825
rect 1630 820 1631 824
rect 1635 820 1636 824
rect 1630 819 1636 820
rect 1710 824 1716 825
rect 1710 820 1711 824
rect 1715 820 1716 824
rect 1710 819 1716 820
rect 1782 824 1788 825
rect 1782 820 1783 824
rect 1787 820 1788 824
rect 1782 819 1788 820
rect 1854 824 1860 825
rect 1854 820 1855 824
rect 1859 820 1860 824
rect 1854 819 1860 820
rect 1934 824 1940 825
rect 1934 820 1935 824
rect 1939 820 1940 824
rect 1934 819 1940 820
rect 2014 824 2020 825
rect 2014 820 2015 824
rect 2019 820 2020 824
rect 2014 819 2020 820
rect 2070 824 2076 825
rect 2070 820 2071 824
rect 2075 820 2076 824
rect 2070 819 2076 820
rect 1160 807 1162 819
rect 1248 807 1250 819
rect 1360 807 1362 819
rect 1456 807 1458 819
rect 1544 807 1546 819
rect 1632 807 1634 819
rect 1712 807 1714 819
rect 1784 807 1786 819
rect 1856 807 1858 819
rect 1936 807 1938 819
rect 2016 807 2018 819
rect 2072 807 2074 819
rect 2120 807 2122 827
rect 1094 803 1100 804
rect 1135 806 1139 807
rect 1135 801 1139 802
rect 1159 806 1163 807
rect 1159 801 1163 802
rect 1247 806 1251 807
rect 1247 801 1251 802
rect 1279 806 1283 807
rect 1279 801 1283 802
rect 1359 806 1363 807
rect 1359 801 1363 802
rect 1407 806 1411 807
rect 1407 801 1411 802
rect 1455 806 1459 807
rect 1455 801 1459 802
rect 1519 806 1523 807
rect 1519 801 1523 802
rect 1543 806 1547 807
rect 1543 801 1547 802
rect 1623 806 1627 807
rect 1623 801 1627 802
rect 1631 806 1635 807
rect 1631 801 1635 802
rect 1711 806 1715 807
rect 1711 801 1715 802
rect 1719 806 1723 807
rect 1719 801 1723 802
rect 1783 806 1787 807
rect 1783 801 1787 802
rect 1815 806 1819 807
rect 1815 801 1819 802
rect 1855 806 1859 807
rect 1855 801 1859 802
rect 1903 806 1907 807
rect 1903 801 1907 802
rect 1935 806 1939 807
rect 1935 801 1939 802
rect 1999 806 2003 807
rect 1999 801 2003 802
rect 2015 806 2019 807
rect 2015 801 2019 802
rect 2071 806 2075 807
rect 2071 801 2075 802
rect 2119 806 2123 807
rect 2119 801 2123 802
rect 110 791 116 792
rect 110 787 111 791
rect 115 787 116 791
rect 1094 791 1100 792
rect 110 786 116 787
rect 278 788 284 789
rect 112 783 114 786
rect 278 784 279 788
rect 283 784 284 788
rect 278 783 284 784
rect 342 788 348 789
rect 342 784 343 788
rect 347 784 348 788
rect 342 783 348 784
rect 414 788 420 789
rect 414 784 415 788
rect 419 784 420 788
rect 414 783 420 784
rect 486 788 492 789
rect 486 784 487 788
rect 491 784 492 788
rect 486 783 492 784
rect 566 788 572 789
rect 566 784 567 788
rect 571 784 572 788
rect 566 783 572 784
rect 646 788 652 789
rect 646 784 647 788
rect 651 784 652 788
rect 646 783 652 784
rect 726 788 732 789
rect 726 784 727 788
rect 731 784 732 788
rect 726 783 732 784
rect 798 788 804 789
rect 798 784 799 788
rect 803 784 804 788
rect 798 783 804 784
rect 862 788 868 789
rect 862 784 863 788
rect 867 784 868 788
rect 862 783 868 784
rect 926 788 932 789
rect 926 784 927 788
rect 931 784 932 788
rect 926 783 932 784
rect 998 788 1004 789
rect 998 784 999 788
rect 1003 784 1004 788
rect 998 783 1004 784
rect 1046 788 1052 789
rect 1046 784 1047 788
rect 1051 784 1052 788
rect 1094 787 1095 791
rect 1099 787 1100 791
rect 1094 786 1100 787
rect 1046 783 1052 784
rect 1096 783 1098 786
rect 111 782 115 783
rect 111 777 115 778
rect 215 782 219 783
rect 215 777 219 778
rect 279 782 283 783
rect 279 777 283 778
rect 343 782 347 783
rect 343 777 347 778
rect 351 782 355 783
rect 351 777 355 778
rect 415 782 419 783
rect 415 777 419 778
rect 423 782 427 783
rect 423 777 427 778
rect 487 782 491 783
rect 487 777 491 778
rect 495 782 499 783
rect 495 777 499 778
rect 567 782 571 783
rect 567 777 571 778
rect 639 782 643 783
rect 639 777 643 778
rect 647 782 651 783
rect 647 777 651 778
rect 703 782 707 783
rect 703 777 707 778
rect 727 782 731 783
rect 727 777 731 778
rect 759 782 763 783
rect 759 777 763 778
rect 799 782 803 783
rect 799 777 803 778
rect 815 782 819 783
rect 815 777 819 778
rect 863 782 867 783
rect 863 777 867 778
rect 911 782 915 783
rect 911 777 915 778
rect 927 782 931 783
rect 927 777 931 778
rect 959 782 963 783
rect 959 777 963 778
rect 999 782 1003 783
rect 999 777 1003 778
rect 1007 782 1011 783
rect 1007 777 1011 778
rect 1047 782 1051 783
rect 1047 777 1051 778
rect 1095 782 1099 783
rect 1136 781 1138 801
rect 1160 789 1162 801
rect 1280 789 1282 801
rect 1408 789 1410 801
rect 1520 789 1522 801
rect 1624 789 1626 801
rect 1720 789 1722 801
rect 1816 789 1818 801
rect 1904 789 1906 801
rect 2000 789 2002 801
rect 2072 789 2074 801
rect 1158 788 1164 789
rect 1158 784 1159 788
rect 1163 784 1164 788
rect 1158 783 1164 784
rect 1278 788 1284 789
rect 1278 784 1279 788
rect 1283 784 1284 788
rect 1278 783 1284 784
rect 1406 788 1412 789
rect 1406 784 1407 788
rect 1411 784 1412 788
rect 1406 783 1412 784
rect 1518 788 1524 789
rect 1518 784 1519 788
rect 1523 784 1524 788
rect 1518 783 1524 784
rect 1622 788 1628 789
rect 1622 784 1623 788
rect 1627 784 1628 788
rect 1622 783 1628 784
rect 1718 788 1724 789
rect 1718 784 1719 788
rect 1723 784 1724 788
rect 1718 783 1724 784
rect 1814 788 1820 789
rect 1814 784 1815 788
rect 1819 784 1820 788
rect 1814 783 1820 784
rect 1902 788 1908 789
rect 1902 784 1903 788
rect 1907 784 1908 788
rect 1902 783 1908 784
rect 1998 788 2004 789
rect 1998 784 1999 788
rect 2003 784 2004 788
rect 1998 783 2004 784
rect 2070 788 2076 789
rect 2070 784 2071 788
rect 2075 784 2076 788
rect 2070 783 2076 784
rect 2120 781 2122 801
rect 1095 777 1099 778
rect 1134 780 1140 781
rect 112 774 114 777
rect 214 776 220 777
rect 110 773 116 774
rect 110 769 111 773
rect 115 769 116 773
rect 214 772 215 776
rect 219 772 220 776
rect 214 771 220 772
rect 278 776 284 777
rect 278 772 279 776
rect 283 772 284 776
rect 278 771 284 772
rect 350 776 356 777
rect 350 772 351 776
rect 355 772 356 776
rect 350 771 356 772
rect 422 776 428 777
rect 422 772 423 776
rect 427 772 428 776
rect 422 771 428 772
rect 494 776 500 777
rect 494 772 495 776
rect 499 772 500 776
rect 494 771 500 772
rect 566 776 572 777
rect 566 772 567 776
rect 571 772 572 776
rect 566 771 572 772
rect 638 776 644 777
rect 638 772 639 776
rect 643 772 644 776
rect 638 771 644 772
rect 702 776 708 777
rect 702 772 703 776
rect 707 772 708 776
rect 702 771 708 772
rect 758 776 764 777
rect 758 772 759 776
rect 763 772 764 776
rect 758 771 764 772
rect 814 776 820 777
rect 814 772 815 776
rect 819 772 820 776
rect 814 771 820 772
rect 862 776 868 777
rect 862 772 863 776
rect 867 772 868 776
rect 862 771 868 772
rect 910 776 916 777
rect 910 772 911 776
rect 915 772 916 776
rect 910 771 916 772
rect 958 776 964 777
rect 958 772 959 776
rect 963 772 964 776
rect 958 771 964 772
rect 1006 776 1012 777
rect 1006 772 1007 776
rect 1011 772 1012 776
rect 1006 771 1012 772
rect 1046 776 1052 777
rect 1046 772 1047 776
rect 1051 772 1052 776
rect 1096 774 1098 777
rect 1134 776 1135 780
rect 1139 776 1140 780
rect 1134 775 1140 776
rect 2118 780 2124 781
rect 2118 776 2119 780
rect 2123 776 2124 780
rect 2118 775 2124 776
rect 1046 771 1052 772
rect 1094 773 1100 774
rect 110 768 116 769
rect 1094 769 1095 773
rect 1099 769 1100 773
rect 1094 768 1100 769
rect 1134 763 1140 764
rect 1134 759 1135 763
rect 1139 759 1140 763
rect 2118 763 2124 764
rect 1134 758 1140 759
rect 1158 760 1164 761
rect 110 756 116 757
rect 110 752 111 756
rect 115 752 116 756
rect 110 751 116 752
rect 1094 756 1100 757
rect 1094 752 1095 756
rect 1099 752 1100 756
rect 1094 751 1100 752
rect 1136 751 1138 758
rect 1158 756 1159 760
rect 1163 756 1164 760
rect 1158 755 1164 756
rect 1278 760 1284 761
rect 1278 756 1279 760
rect 1283 756 1284 760
rect 1278 755 1284 756
rect 1406 760 1412 761
rect 1406 756 1407 760
rect 1411 756 1412 760
rect 1406 755 1412 756
rect 1518 760 1524 761
rect 1518 756 1519 760
rect 1523 756 1524 760
rect 1518 755 1524 756
rect 1622 760 1628 761
rect 1622 756 1623 760
rect 1627 756 1628 760
rect 1622 755 1628 756
rect 1718 760 1724 761
rect 1718 756 1719 760
rect 1723 756 1724 760
rect 1718 755 1724 756
rect 1814 760 1820 761
rect 1814 756 1815 760
rect 1819 756 1820 760
rect 1814 755 1820 756
rect 1902 760 1908 761
rect 1902 756 1903 760
rect 1907 756 1908 760
rect 1902 755 1908 756
rect 1998 760 2004 761
rect 1998 756 1999 760
rect 2003 756 2004 760
rect 1998 755 2004 756
rect 2070 760 2076 761
rect 2070 756 2071 760
rect 2075 756 2076 760
rect 2118 759 2119 763
rect 2123 759 2124 763
rect 2118 758 2124 759
rect 2070 755 2076 756
rect 1160 751 1162 755
rect 1280 751 1282 755
rect 1408 751 1410 755
rect 1520 751 1522 755
rect 1624 751 1626 755
rect 1720 751 1722 755
rect 1816 751 1818 755
rect 1904 751 1906 755
rect 2000 751 2002 755
rect 2072 751 2074 755
rect 2120 751 2122 758
rect 112 731 114 751
rect 214 748 220 749
rect 214 744 215 748
rect 219 744 220 748
rect 214 743 220 744
rect 278 748 284 749
rect 278 744 279 748
rect 283 744 284 748
rect 278 743 284 744
rect 350 748 356 749
rect 350 744 351 748
rect 355 744 356 748
rect 350 743 356 744
rect 422 748 428 749
rect 422 744 423 748
rect 427 744 428 748
rect 422 743 428 744
rect 494 748 500 749
rect 494 744 495 748
rect 499 744 500 748
rect 494 743 500 744
rect 566 748 572 749
rect 566 744 567 748
rect 571 744 572 748
rect 566 743 572 744
rect 638 748 644 749
rect 638 744 639 748
rect 643 744 644 748
rect 638 743 644 744
rect 702 748 708 749
rect 702 744 703 748
rect 707 744 708 748
rect 702 743 708 744
rect 758 748 764 749
rect 758 744 759 748
rect 763 744 764 748
rect 758 743 764 744
rect 814 748 820 749
rect 814 744 815 748
rect 819 744 820 748
rect 814 743 820 744
rect 862 748 868 749
rect 862 744 863 748
rect 867 744 868 748
rect 862 743 868 744
rect 910 748 916 749
rect 910 744 911 748
rect 915 744 916 748
rect 910 743 916 744
rect 958 748 964 749
rect 958 744 959 748
rect 963 744 964 748
rect 958 743 964 744
rect 1006 748 1012 749
rect 1006 744 1007 748
rect 1011 744 1012 748
rect 1006 743 1012 744
rect 1046 748 1052 749
rect 1046 744 1047 748
rect 1051 744 1052 748
rect 1046 743 1052 744
rect 216 731 218 743
rect 280 731 282 743
rect 352 731 354 743
rect 424 731 426 743
rect 496 731 498 743
rect 568 731 570 743
rect 640 731 642 743
rect 704 731 706 743
rect 760 731 762 743
rect 816 731 818 743
rect 864 731 866 743
rect 912 731 914 743
rect 960 731 962 743
rect 1008 731 1010 743
rect 1048 731 1050 743
rect 1096 731 1098 751
rect 1135 750 1139 751
rect 1135 745 1139 746
rect 1159 750 1163 751
rect 1159 745 1163 746
rect 1279 750 1283 751
rect 1279 745 1283 746
rect 1335 750 1339 751
rect 1335 745 1339 746
rect 1375 750 1379 751
rect 1375 745 1379 746
rect 1407 750 1411 751
rect 1407 745 1411 746
rect 1415 750 1419 751
rect 1415 745 1419 746
rect 1455 750 1459 751
rect 1455 745 1459 746
rect 1503 750 1507 751
rect 1503 745 1507 746
rect 1519 750 1523 751
rect 1519 745 1523 746
rect 1551 750 1555 751
rect 1551 745 1555 746
rect 1599 750 1603 751
rect 1599 745 1603 746
rect 1623 750 1627 751
rect 1623 745 1627 746
rect 1655 750 1659 751
rect 1655 745 1659 746
rect 1711 750 1715 751
rect 1711 745 1715 746
rect 1719 750 1723 751
rect 1719 745 1723 746
rect 1767 750 1771 751
rect 1767 745 1771 746
rect 1815 750 1819 751
rect 1815 745 1819 746
rect 1831 750 1835 751
rect 1831 745 1835 746
rect 1895 750 1899 751
rect 1895 745 1899 746
rect 1903 750 1907 751
rect 1903 745 1907 746
rect 1959 750 1963 751
rect 1959 745 1963 746
rect 1999 750 2003 751
rect 1999 745 2003 746
rect 2023 750 2027 751
rect 2023 745 2027 746
rect 2071 750 2075 751
rect 2071 745 2075 746
rect 2119 750 2123 751
rect 2119 745 2123 746
rect 1136 742 1138 745
rect 1334 744 1340 745
rect 1134 741 1140 742
rect 1134 737 1135 741
rect 1139 737 1140 741
rect 1334 740 1335 744
rect 1339 740 1340 744
rect 1334 739 1340 740
rect 1374 744 1380 745
rect 1374 740 1375 744
rect 1379 740 1380 744
rect 1374 739 1380 740
rect 1414 744 1420 745
rect 1414 740 1415 744
rect 1419 740 1420 744
rect 1414 739 1420 740
rect 1454 744 1460 745
rect 1454 740 1455 744
rect 1459 740 1460 744
rect 1454 739 1460 740
rect 1502 744 1508 745
rect 1502 740 1503 744
rect 1507 740 1508 744
rect 1502 739 1508 740
rect 1550 744 1556 745
rect 1550 740 1551 744
rect 1555 740 1556 744
rect 1550 739 1556 740
rect 1598 744 1604 745
rect 1598 740 1599 744
rect 1603 740 1604 744
rect 1598 739 1604 740
rect 1654 744 1660 745
rect 1654 740 1655 744
rect 1659 740 1660 744
rect 1654 739 1660 740
rect 1710 744 1716 745
rect 1710 740 1711 744
rect 1715 740 1716 744
rect 1710 739 1716 740
rect 1766 744 1772 745
rect 1766 740 1767 744
rect 1771 740 1772 744
rect 1766 739 1772 740
rect 1830 744 1836 745
rect 1830 740 1831 744
rect 1835 740 1836 744
rect 1830 739 1836 740
rect 1894 744 1900 745
rect 1894 740 1895 744
rect 1899 740 1900 744
rect 1894 739 1900 740
rect 1958 744 1964 745
rect 1958 740 1959 744
rect 1963 740 1964 744
rect 1958 739 1964 740
rect 2022 744 2028 745
rect 2022 740 2023 744
rect 2027 740 2028 744
rect 2022 739 2028 740
rect 2070 744 2076 745
rect 2070 740 2071 744
rect 2075 740 2076 744
rect 2120 742 2122 745
rect 2070 739 2076 740
rect 2118 741 2124 742
rect 1134 736 1140 737
rect 2118 737 2119 741
rect 2123 737 2124 741
rect 2118 736 2124 737
rect 111 730 115 731
rect 111 725 115 726
rect 175 730 179 731
rect 175 725 179 726
rect 215 730 219 731
rect 215 725 219 726
rect 239 730 243 731
rect 239 725 243 726
rect 279 730 283 731
rect 279 725 283 726
rect 311 730 315 731
rect 311 725 315 726
rect 351 730 355 731
rect 351 725 355 726
rect 391 730 395 731
rect 391 725 395 726
rect 423 730 427 731
rect 423 725 427 726
rect 471 730 475 731
rect 471 725 475 726
rect 495 730 499 731
rect 495 725 499 726
rect 543 730 547 731
rect 543 725 547 726
rect 567 730 571 731
rect 567 725 571 726
rect 615 730 619 731
rect 615 725 619 726
rect 639 730 643 731
rect 639 725 643 726
rect 679 730 683 731
rect 679 725 683 726
rect 703 730 707 731
rect 703 725 707 726
rect 735 730 739 731
rect 735 725 739 726
rect 759 730 763 731
rect 759 725 763 726
rect 799 730 803 731
rect 799 725 803 726
rect 815 730 819 731
rect 815 725 819 726
rect 863 730 867 731
rect 863 725 867 726
rect 911 730 915 731
rect 911 725 915 726
rect 927 730 931 731
rect 927 725 931 726
rect 959 730 963 731
rect 959 725 963 726
rect 1007 730 1011 731
rect 1007 725 1011 726
rect 1047 730 1051 731
rect 1047 725 1051 726
rect 1095 730 1099 731
rect 1095 725 1099 726
rect 112 705 114 725
rect 176 713 178 725
rect 240 713 242 725
rect 312 713 314 725
rect 392 713 394 725
rect 472 713 474 725
rect 544 713 546 725
rect 616 713 618 725
rect 680 713 682 725
rect 736 713 738 725
rect 800 713 802 725
rect 864 713 866 725
rect 928 713 930 725
rect 174 712 180 713
rect 174 708 175 712
rect 179 708 180 712
rect 174 707 180 708
rect 238 712 244 713
rect 238 708 239 712
rect 243 708 244 712
rect 238 707 244 708
rect 310 712 316 713
rect 310 708 311 712
rect 315 708 316 712
rect 310 707 316 708
rect 390 712 396 713
rect 390 708 391 712
rect 395 708 396 712
rect 390 707 396 708
rect 470 712 476 713
rect 470 708 471 712
rect 475 708 476 712
rect 470 707 476 708
rect 542 712 548 713
rect 542 708 543 712
rect 547 708 548 712
rect 542 707 548 708
rect 614 712 620 713
rect 614 708 615 712
rect 619 708 620 712
rect 614 707 620 708
rect 678 712 684 713
rect 678 708 679 712
rect 683 708 684 712
rect 678 707 684 708
rect 734 712 740 713
rect 734 708 735 712
rect 739 708 740 712
rect 734 707 740 708
rect 798 712 804 713
rect 798 708 799 712
rect 803 708 804 712
rect 798 707 804 708
rect 862 712 868 713
rect 862 708 863 712
rect 867 708 868 712
rect 862 707 868 708
rect 926 712 932 713
rect 926 708 927 712
rect 931 708 932 712
rect 926 707 932 708
rect 1096 705 1098 725
rect 1134 724 1140 725
rect 1134 720 1135 724
rect 1139 720 1140 724
rect 1134 719 1140 720
rect 2118 724 2124 725
rect 2118 720 2119 724
rect 2123 720 2124 724
rect 2118 719 2124 720
rect 110 704 116 705
rect 110 700 111 704
rect 115 700 116 704
rect 110 699 116 700
rect 1094 704 1100 705
rect 1094 700 1095 704
rect 1099 700 1100 704
rect 1094 699 1100 700
rect 1136 699 1138 719
rect 1334 716 1340 717
rect 1334 712 1335 716
rect 1339 712 1340 716
rect 1334 711 1340 712
rect 1374 716 1380 717
rect 1374 712 1375 716
rect 1379 712 1380 716
rect 1374 711 1380 712
rect 1414 716 1420 717
rect 1414 712 1415 716
rect 1419 712 1420 716
rect 1414 711 1420 712
rect 1454 716 1460 717
rect 1454 712 1455 716
rect 1459 712 1460 716
rect 1454 711 1460 712
rect 1502 716 1508 717
rect 1502 712 1503 716
rect 1507 712 1508 716
rect 1502 711 1508 712
rect 1550 716 1556 717
rect 1550 712 1551 716
rect 1555 712 1556 716
rect 1550 711 1556 712
rect 1598 716 1604 717
rect 1598 712 1599 716
rect 1603 712 1604 716
rect 1598 711 1604 712
rect 1654 716 1660 717
rect 1654 712 1655 716
rect 1659 712 1660 716
rect 1654 711 1660 712
rect 1710 716 1716 717
rect 1710 712 1711 716
rect 1715 712 1716 716
rect 1710 711 1716 712
rect 1766 716 1772 717
rect 1766 712 1767 716
rect 1771 712 1772 716
rect 1766 711 1772 712
rect 1830 716 1836 717
rect 1830 712 1831 716
rect 1835 712 1836 716
rect 1830 711 1836 712
rect 1894 716 1900 717
rect 1894 712 1895 716
rect 1899 712 1900 716
rect 1894 711 1900 712
rect 1958 716 1964 717
rect 1958 712 1959 716
rect 1963 712 1964 716
rect 1958 711 1964 712
rect 2022 716 2028 717
rect 2022 712 2023 716
rect 2027 712 2028 716
rect 2022 711 2028 712
rect 2070 716 2076 717
rect 2070 712 2071 716
rect 2075 712 2076 716
rect 2070 711 2076 712
rect 1336 699 1338 711
rect 1376 699 1378 711
rect 1416 699 1418 711
rect 1456 699 1458 711
rect 1504 699 1506 711
rect 1552 699 1554 711
rect 1600 699 1602 711
rect 1656 699 1658 711
rect 1712 699 1714 711
rect 1768 699 1770 711
rect 1832 699 1834 711
rect 1896 699 1898 711
rect 1960 699 1962 711
rect 2024 699 2026 711
rect 2072 699 2074 711
rect 2120 699 2122 719
rect 1135 698 1139 699
rect 1135 693 1139 694
rect 1247 698 1251 699
rect 1247 693 1251 694
rect 1287 698 1291 699
rect 1287 693 1291 694
rect 1335 698 1339 699
rect 1335 693 1339 694
rect 1375 698 1379 699
rect 1375 693 1379 694
rect 1391 698 1395 699
rect 1391 693 1395 694
rect 1415 698 1419 699
rect 1415 693 1419 694
rect 1447 698 1451 699
rect 1447 693 1451 694
rect 1455 698 1459 699
rect 1455 693 1459 694
rect 1503 698 1507 699
rect 1503 693 1507 694
rect 1511 698 1515 699
rect 1511 693 1515 694
rect 1551 698 1555 699
rect 1551 693 1555 694
rect 1583 698 1587 699
rect 1583 693 1587 694
rect 1599 698 1603 699
rect 1599 693 1603 694
rect 1655 698 1659 699
rect 1655 693 1659 694
rect 1711 698 1715 699
rect 1711 693 1715 694
rect 1735 698 1739 699
rect 1735 693 1739 694
rect 1767 698 1771 699
rect 1767 693 1771 694
rect 1823 698 1827 699
rect 1823 693 1827 694
rect 1831 698 1835 699
rect 1831 693 1835 694
rect 1895 698 1899 699
rect 1895 693 1899 694
rect 1911 698 1915 699
rect 1911 693 1915 694
rect 1959 698 1963 699
rect 1959 693 1963 694
rect 1999 698 2003 699
rect 1999 693 2003 694
rect 2023 698 2027 699
rect 2023 693 2027 694
rect 2071 698 2075 699
rect 2071 693 2075 694
rect 2119 698 2123 699
rect 2119 693 2123 694
rect 110 687 116 688
rect 110 683 111 687
rect 115 683 116 687
rect 1094 687 1100 688
rect 110 682 116 683
rect 174 684 180 685
rect 112 679 114 682
rect 174 680 175 684
rect 179 680 180 684
rect 174 679 180 680
rect 238 684 244 685
rect 238 680 239 684
rect 243 680 244 684
rect 238 679 244 680
rect 310 684 316 685
rect 310 680 311 684
rect 315 680 316 684
rect 310 679 316 680
rect 390 684 396 685
rect 390 680 391 684
rect 395 680 396 684
rect 390 679 396 680
rect 470 684 476 685
rect 470 680 471 684
rect 475 680 476 684
rect 470 679 476 680
rect 542 684 548 685
rect 542 680 543 684
rect 547 680 548 684
rect 542 679 548 680
rect 614 684 620 685
rect 614 680 615 684
rect 619 680 620 684
rect 614 679 620 680
rect 678 684 684 685
rect 678 680 679 684
rect 683 680 684 684
rect 678 679 684 680
rect 734 684 740 685
rect 734 680 735 684
rect 739 680 740 684
rect 734 679 740 680
rect 798 684 804 685
rect 798 680 799 684
rect 803 680 804 684
rect 798 679 804 680
rect 862 684 868 685
rect 862 680 863 684
rect 867 680 868 684
rect 862 679 868 680
rect 926 684 932 685
rect 926 680 927 684
rect 931 680 932 684
rect 1094 683 1095 687
rect 1099 683 1100 687
rect 1094 682 1100 683
rect 926 679 932 680
rect 1096 679 1098 682
rect 111 678 115 679
rect 111 673 115 674
rect 135 678 139 679
rect 135 673 139 674
rect 175 678 179 679
rect 175 673 179 674
rect 215 678 219 679
rect 215 673 219 674
rect 239 678 243 679
rect 239 673 243 674
rect 271 678 275 679
rect 271 673 275 674
rect 311 678 315 679
rect 311 673 315 674
rect 335 678 339 679
rect 335 673 339 674
rect 391 678 395 679
rect 391 673 395 674
rect 399 678 403 679
rect 399 673 403 674
rect 463 678 467 679
rect 463 673 467 674
rect 471 678 475 679
rect 471 673 475 674
rect 527 678 531 679
rect 527 673 531 674
rect 543 678 547 679
rect 543 673 547 674
rect 591 678 595 679
rect 591 673 595 674
rect 615 678 619 679
rect 615 673 619 674
rect 647 678 651 679
rect 647 673 651 674
rect 679 678 683 679
rect 679 673 683 674
rect 703 678 707 679
rect 703 673 707 674
rect 735 678 739 679
rect 735 673 739 674
rect 759 678 763 679
rect 759 673 763 674
rect 799 678 803 679
rect 799 673 803 674
rect 823 678 827 679
rect 823 673 827 674
rect 863 678 867 679
rect 863 673 867 674
rect 927 678 931 679
rect 927 673 931 674
rect 1095 678 1099 679
rect 1095 673 1099 674
rect 1136 673 1138 693
rect 1248 681 1250 693
rect 1288 681 1290 693
rect 1336 681 1338 693
rect 1392 681 1394 693
rect 1448 681 1450 693
rect 1512 681 1514 693
rect 1584 681 1586 693
rect 1656 681 1658 693
rect 1736 681 1738 693
rect 1824 681 1826 693
rect 1912 681 1914 693
rect 2000 681 2002 693
rect 2072 681 2074 693
rect 1246 680 1252 681
rect 1246 676 1247 680
rect 1251 676 1252 680
rect 1246 675 1252 676
rect 1286 680 1292 681
rect 1286 676 1287 680
rect 1291 676 1292 680
rect 1286 675 1292 676
rect 1334 680 1340 681
rect 1334 676 1335 680
rect 1339 676 1340 680
rect 1334 675 1340 676
rect 1390 680 1396 681
rect 1390 676 1391 680
rect 1395 676 1396 680
rect 1390 675 1396 676
rect 1446 680 1452 681
rect 1446 676 1447 680
rect 1451 676 1452 680
rect 1446 675 1452 676
rect 1510 680 1516 681
rect 1510 676 1511 680
rect 1515 676 1516 680
rect 1510 675 1516 676
rect 1582 680 1588 681
rect 1582 676 1583 680
rect 1587 676 1588 680
rect 1582 675 1588 676
rect 1654 680 1660 681
rect 1654 676 1655 680
rect 1659 676 1660 680
rect 1654 675 1660 676
rect 1734 680 1740 681
rect 1734 676 1735 680
rect 1739 676 1740 680
rect 1734 675 1740 676
rect 1822 680 1828 681
rect 1822 676 1823 680
rect 1827 676 1828 680
rect 1822 675 1828 676
rect 1910 680 1916 681
rect 1910 676 1911 680
rect 1915 676 1916 680
rect 1910 675 1916 676
rect 1998 680 2004 681
rect 1998 676 1999 680
rect 2003 676 2004 680
rect 1998 675 2004 676
rect 2070 680 2076 681
rect 2070 676 2071 680
rect 2075 676 2076 680
rect 2070 675 2076 676
rect 2120 673 2122 693
rect 112 670 114 673
rect 134 672 140 673
rect 110 669 116 670
rect 110 665 111 669
rect 115 665 116 669
rect 134 668 135 672
rect 139 668 140 672
rect 134 667 140 668
rect 174 672 180 673
rect 174 668 175 672
rect 179 668 180 672
rect 174 667 180 668
rect 214 672 220 673
rect 214 668 215 672
rect 219 668 220 672
rect 214 667 220 668
rect 270 672 276 673
rect 270 668 271 672
rect 275 668 276 672
rect 270 667 276 668
rect 334 672 340 673
rect 334 668 335 672
rect 339 668 340 672
rect 334 667 340 668
rect 398 672 404 673
rect 398 668 399 672
rect 403 668 404 672
rect 398 667 404 668
rect 462 672 468 673
rect 462 668 463 672
rect 467 668 468 672
rect 462 667 468 668
rect 526 672 532 673
rect 526 668 527 672
rect 531 668 532 672
rect 526 667 532 668
rect 590 672 596 673
rect 590 668 591 672
rect 595 668 596 672
rect 590 667 596 668
rect 646 672 652 673
rect 646 668 647 672
rect 651 668 652 672
rect 646 667 652 668
rect 702 672 708 673
rect 702 668 703 672
rect 707 668 708 672
rect 702 667 708 668
rect 758 672 764 673
rect 758 668 759 672
rect 763 668 764 672
rect 758 667 764 668
rect 822 672 828 673
rect 822 668 823 672
rect 827 668 828 672
rect 1096 670 1098 673
rect 1134 672 1140 673
rect 822 667 828 668
rect 1094 669 1100 670
rect 110 664 116 665
rect 1094 665 1095 669
rect 1099 665 1100 669
rect 1134 668 1135 672
rect 1139 668 1140 672
rect 1134 667 1140 668
rect 2118 672 2124 673
rect 2118 668 2119 672
rect 2123 668 2124 672
rect 2118 667 2124 668
rect 1094 664 1100 665
rect 1134 655 1140 656
rect 110 652 116 653
rect 110 648 111 652
rect 115 648 116 652
rect 110 647 116 648
rect 1094 652 1100 653
rect 1094 648 1095 652
rect 1099 648 1100 652
rect 1134 651 1135 655
rect 1139 651 1140 655
rect 2118 655 2124 656
rect 1134 650 1140 651
rect 1246 652 1252 653
rect 1094 647 1100 648
rect 1136 647 1138 650
rect 1246 648 1247 652
rect 1251 648 1252 652
rect 1246 647 1252 648
rect 1286 652 1292 653
rect 1286 648 1287 652
rect 1291 648 1292 652
rect 1286 647 1292 648
rect 1334 652 1340 653
rect 1334 648 1335 652
rect 1339 648 1340 652
rect 1334 647 1340 648
rect 1390 652 1396 653
rect 1390 648 1391 652
rect 1395 648 1396 652
rect 1390 647 1396 648
rect 1446 652 1452 653
rect 1446 648 1447 652
rect 1451 648 1452 652
rect 1446 647 1452 648
rect 1510 652 1516 653
rect 1510 648 1511 652
rect 1515 648 1516 652
rect 1510 647 1516 648
rect 1582 652 1588 653
rect 1582 648 1583 652
rect 1587 648 1588 652
rect 1582 647 1588 648
rect 1654 652 1660 653
rect 1654 648 1655 652
rect 1659 648 1660 652
rect 1654 647 1660 648
rect 1734 652 1740 653
rect 1734 648 1735 652
rect 1739 648 1740 652
rect 1734 647 1740 648
rect 1822 652 1828 653
rect 1822 648 1823 652
rect 1827 648 1828 652
rect 1822 647 1828 648
rect 1910 652 1916 653
rect 1910 648 1911 652
rect 1915 648 1916 652
rect 1910 647 1916 648
rect 1998 652 2004 653
rect 1998 648 1999 652
rect 2003 648 2004 652
rect 1998 647 2004 648
rect 2070 652 2076 653
rect 2070 648 2071 652
rect 2075 648 2076 652
rect 2118 651 2119 655
rect 2123 651 2124 655
rect 2118 650 2124 651
rect 2070 647 2076 648
rect 2120 647 2122 650
rect 112 619 114 647
rect 134 644 140 645
rect 134 640 135 644
rect 139 640 140 644
rect 134 639 140 640
rect 174 644 180 645
rect 174 640 175 644
rect 179 640 180 644
rect 174 639 180 640
rect 214 644 220 645
rect 214 640 215 644
rect 219 640 220 644
rect 214 639 220 640
rect 270 644 276 645
rect 270 640 271 644
rect 275 640 276 644
rect 270 639 276 640
rect 334 644 340 645
rect 334 640 335 644
rect 339 640 340 644
rect 334 639 340 640
rect 398 644 404 645
rect 398 640 399 644
rect 403 640 404 644
rect 398 639 404 640
rect 462 644 468 645
rect 462 640 463 644
rect 467 640 468 644
rect 462 639 468 640
rect 526 644 532 645
rect 526 640 527 644
rect 531 640 532 644
rect 526 639 532 640
rect 590 644 596 645
rect 590 640 591 644
rect 595 640 596 644
rect 590 639 596 640
rect 646 644 652 645
rect 646 640 647 644
rect 651 640 652 644
rect 646 639 652 640
rect 702 644 708 645
rect 702 640 703 644
rect 707 640 708 644
rect 702 639 708 640
rect 758 644 764 645
rect 758 640 759 644
rect 763 640 764 644
rect 758 639 764 640
rect 822 644 828 645
rect 822 640 823 644
rect 827 640 828 644
rect 822 639 828 640
rect 136 619 138 639
rect 176 619 178 639
rect 216 619 218 639
rect 272 619 274 639
rect 336 619 338 639
rect 400 619 402 639
rect 464 619 466 639
rect 528 619 530 639
rect 592 619 594 639
rect 648 619 650 639
rect 704 619 706 639
rect 760 619 762 639
rect 824 619 826 639
rect 1096 619 1098 647
rect 1135 646 1139 647
rect 1135 641 1139 642
rect 1159 646 1163 647
rect 1159 641 1163 642
rect 1199 646 1203 647
rect 1199 641 1203 642
rect 1239 646 1243 647
rect 1239 641 1243 642
rect 1247 646 1251 647
rect 1247 641 1251 642
rect 1279 646 1283 647
rect 1279 641 1283 642
rect 1287 646 1291 647
rect 1287 641 1291 642
rect 1335 646 1339 647
rect 1335 641 1339 642
rect 1343 646 1347 647
rect 1343 641 1347 642
rect 1391 646 1395 647
rect 1391 641 1395 642
rect 1415 646 1419 647
rect 1415 641 1419 642
rect 1447 646 1451 647
rect 1447 641 1451 642
rect 1495 646 1499 647
rect 1495 641 1499 642
rect 1511 646 1515 647
rect 1511 641 1515 642
rect 1583 646 1587 647
rect 1583 641 1587 642
rect 1655 646 1659 647
rect 1655 641 1659 642
rect 1671 646 1675 647
rect 1671 641 1675 642
rect 1735 646 1739 647
rect 1735 641 1739 642
rect 1759 646 1763 647
rect 1759 641 1763 642
rect 1823 646 1827 647
rect 1823 641 1827 642
rect 1839 646 1843 647
rect 1839 641 1843 642
rect 1911 646 1915 647
rect 1911 641 1915 642
rect 1919 646 1923 647
rect 1919 641 1923 642
rect 1999 646 2003 647
rect 1999 641 2003 642
rect 2007 646 2011 647
rect 2007 641 2011 642
rect 2071 646 2075 647
rect 2071 641 2075 642
rect 2119 646 2123 647
rect 2119 641 2123 642
rect 1136 638 1138 641
rect 1158 640 1164 641
rect 1134 637 1140 638
rect 1134 633 1135 637
rect 1139 633 1140 637
rect 1158 636 1159 640
rect 1163 636 1164 640
rect 1158 635 1164 636
rect 1198 640 1204 641
rect 1198 636 1199 640
rect 1203 636 1204 640
rect 1198 635 1204 636
rect 1238 640 1244 641
rect 1238 636 1239 640
rect 1243 636 1244 640
rect 1238 635 1244 636
rect 1278 640 1284 641
rect 1278 636 1279 640
rect 1283 636 1284 640
rect 1278 635 1284 636
rect 1342 640 1348 641
rect 1342 636 1343 640
rect 1347 636 1348 640
rect 1342 635 1348 636
rect 1414 640 1420 641
rect 1414 636 1415 640
rect 1419 636 1420 640
rect 1414 635 1420 636
rect 1494 640 1500 641
rect 1494 636 1495 640
rect 1499 636 1500 640
rect 1494 635 1500 636
rect 1582 640 1588 641
rect 1582 636 1583 640
rect 1587 636 1588 640
rect 1582 635 1588 636
rect 1670 640 1676 641
rect 1670 636 1671 640
rect 1675 636 1676 640
rect 1670 635 1676 636
rect 1758 640 1764 641
rect 1758 636 1759 640
rect 1763 636 1764 640
rect 1758 635 1764 636
rect 1838 640 1844 641
rect 1838 636 1839 640
rect 1843 636 1844 640
rect 1838 635 1844 636
rect 1918 640 1924 641
rect 1918 636 1919 640
rect 1923 636 1924 640
rect 1918 635 1924 636
rect 2006 640 2012 641
rect 2006 636 2007 640
rect 2011 636 2012 640
rect 2006 635 2012 636
rect 2070 640 2076 641
rect 2070 636 2071 640
rect 2075 636 2076 640
rect 2120 638 2122 641
rect 2070 635 2076 636
rect 2118 637 2124 638
rect 1134 632 1140 633
rect 2118 633 2119 637
rect 2123 633 2124 637
rect 2118 632 2124 633
rect 1134 620 1140 621
rect 111 618 115 619
rect 111 613 115 614
rect 135 618 139 619
rect 135 613 139 614
rect 175 618 179 619
rect 175 613 179 614
rect 215 618 219 619
rect 215 613 219 614
rect 255 618 259 619
rect 255 613 259 614
rect 271 618 275 619
rect 271 613 275 614
rect 303 618 307 619
rect 303 613 307 614
rect 335 618 339 619
rect 335 613 339 614
rect 351 618 355 619
rect 351 613 355 614
rect 399 618 403 619
rect 399 613 403 614
rect 439 618 443 619
rect 439 613 443 614
rect 463 618 467 619
rect 463 613 467 614
rect 487 618 491 619
rect 487 613 491 614
rect 527 618 531 619
rect 527 613 531 614
rect 535 618 539 619
rect 535 613 539 614
rect 583 618 587 619
rect 583 613 587 614
rect 591 618 595 619
rect 591 613 595 614
rect 631 618 635 619
rect 631 613 635 614
rect 647 618 651 619
rect 647 613 651 614
rect 679 618 683 619
rect 679 613 683 614
rect 703 618 707 619
rect 703 613 707 614
rect 727 618 731 619
rect 727 613 731 614
rect 759 618 763 619
rect 759 613 763 614
rect 823 618 827 619
rect 823 613 827 614
rect 1095 618 1099 619
rect 1134 616 1135 620
rect 1139 616 1140 620
rect 1134 615 1140 616
rect 2118 620 2124 621
rect 2118 616 2119 620
rect 2123 616 2124 620
rect 2118 615 2124 616
rect 1095 613 1099 614
rect 112 593 114 613
rect 136 601 138 613
rect 176 601 178 613
rect 216 601 218 613
rect 256 601 258 613
rect 304 601 306 613
rect 352 601 354 613
rect 400 601 402 613
rect 440 601 442 613
rect 488 601 490 613
rect 536 601 538 613
rect 584 601 586 613
rect 632 601 634 613
rect 680 601 682 613
rect 728 601 730 613
rect 134 600 140 601
rect 134 596 135 600
rect 139 596 140 600
rect 134 595 140 596
rect 174 600 180 601
rect 174 596 175 600
rect 179 596 180 600
rect 174 595 180 596
rect 214 600 220 601
rect 214 596 215 600
rect 219 596 220 600
rect 214 595 220 596
rect 254 600 260 601
rect 254 596 255 600
rect 259 596 260 600
rect 254 595 260 596
rect 302 600 308 601
rect 302 596 303 600
rect 307 596 308 600
rect 302 595 308 596
rect 350 600 356 601
rect 350 596 351 600
rect 355 596 356 600
rect 350 595 356 596
rect 398 600 404 601
rect 398 596 399 600
rect 403 596 404 600
rect 398 595 404 596
rect 438 600 444 601
rect 438 596 439 600
rect 443 596 444 600
rect 438 595 444 596
rect 486 600 492 601
rect 486 596 487 600
rect 491 596 492 600
rect 486 595 492 596
rect 534 600 540 601
rect 534 596 535 600
rect 539 596 540 600
rect 534 595 540 596
rect 582 600 588 601
rect 582 596 583 600
rect 587 596 588 600
rect 582 595 588 596
rect 630 600 636 601
rect 630 596 631 600
rect 635 596 636 600
rect 630 595 636 596
rect 678 600 684 601
rect 678 596 679 600
rect 683 596 684 600
rect 678 595 684 596
rect 726 600 732 601
rect 726 596 727 600
rect 731 596 732 600
rect 726 595 732 596
rect 1096 593 1098 613
rect 110 592 116 593
rect 110 588 111 592
rect 115 588 116 592
rect 110 587 116 588
rect 1094 592 1100 593
rect 1094 588 1095 592
rect 1099 588 1100 592
rect 1136 591 1138 615
rect 1158 612 1164 613
rect 1158 608 1159 612
rect 1163 608 1164 612
rect 1158 607 1164 608
rect 1198 612 1204 613
rect 1198 608 1199 612
rect 1203 608 1204 612
rect 1198 607 1204 608
rect 1238 612 1244 613
rect 1238 608 1239 612
rect 1243 608 1244 612
rect 1238 607 1244 608
rect 1278 612 1284 613
rect 1278 608 1279 612
rect 1283 608 1284 612
rect 1278 607 1284 608
rect 1342 612 1348 613
rect 1342 608 1343 612
rect 1347 608 1348 612
rect 1342 607 1348 608
rect 1414 612 1420 613
rect 1414 608 1415 612
rect 1419 608 1420 612
rect 1414 607 1420 608
rect 1494 612 1500 613
rect 1494 608 1495 612
rect 1499 608 1500 612
rect 1494 607 1500 608
rect 1582 612 1588 613
rect 1582 608 1583 612
rect 1587 608 1588 612
rect 1582 607 1588 608
rect 1670 612 1676 613
rect 1670 608 1671 612
rect 1675 608 1676 612
rect 1670 607 1676 608
rect 1758 612 1764 613
rect 1758 608 1759 612
rect 1763 608 1764 612
rect 1758 607 1764 608
rect 1838 612 1844 613
rect 1838 608 1839 612
rect 1843 608 1844 612
rect 1838 607 1844 608
rect 1918 612 1924 613
rect 1918 608 1919 612
rect 1923 608 1924 612
rect 1918 607 1924 608
rect 2006 612 2012 613
rect 2006 608 2007 612
rect 2011 608 2012 612
rect 2006 607 2012 608
rect 2070 612 2076 613
rect 2070 608 2071 612
rect 2075 608 2076 612
rect 2070 607 2076 608
rect 1160 591 1162 607
rect 1200 591 1202 607
rect 1240 591 1242 607
rect 1280 591 1282 607
rect 1344 591 1346 607
rect 1416 591 1418 607
rect 1496 591 1498 607
rect 1584 591 1586 607
rect 1672 591 1674 607
rect 1760 591 1762 607
rect 1840 591 1842 607
rect 1920 591 1922 607
rect 2008 591 2010 607
rect 2072 591 2074 607
rect 2120 591 2122 615
rect 1094 587 1100 588
rect 1135 590 1139 591
rect 1135 585 1139 586
rect 1159 590 1163 591
rect 1159 585 1163 586
rect 1199 590 1203 591
rect 1199 585 1203 586
rect 1239 590 1243 591
rect 1239 585 1243 586
rect 1279 590 1283 591
rect 1279 585 1283 586
rect 1319 590 1323 591
rect 1319 585 1323 586
rect 1343 590 1347 591
rect 1343 585 1347 586
rect 1359 590 1363 591
rect 1359 585 1363 586
rect 1415 590 1419 591
rect 1415 585 1419 586
rect 1487 590 1491 591
rect 1487 585 1491 586
rect 1495 590 1499 591
rect 1495 585 1499 586
rect 1567 590 1571 591
rect 1567 585 1571 586
rect 1583 590 1587 591
rect 1583 585 1587 586
rect 1655 590 1659 591
rect 1655 585 1659 586
rect 1671 590 1675 591
rect 1671 585 1675 586
rect 1751 590 1755 591
rect 1751 585 1755 586
rect 1759 590 1763 591
rect 1759 585 1763 586
rect 1839 590 1843 591
rect 1839 585 1843 586
rect 1855 590 1859 591
rect 1855 585 1859 586
rect 1919 590 1923 591
rect 1919 585 1923 586
rect 1967 590 1971 591
rect 1967 585 1971 586
rect 2007 590 2011 591
rect 2007 585 2011 586
rect 2071 590 2075 591
rect 2071 585 2075 586
rect 2119 590 2123 591
rect 2119 585 2123 586
rect 110 575 116 576
rect 110 571 111 575
rect 115 571 116 575
rect 1094 575 1100 576
rect 110 570 116 571
rect 134 572 140 573
rect 112 563 114 570
rect 134 568 135 572
rect 139 568 140 572
rect 134 567 140 568
rect 174 572 180 573
rect 174 568 175 572
rect 179 568 180 572
rect 174 567 180 568
rect 214 572 220 573
rect 214 568 215 572
rect 219 568 220 572
rect 214 567 220 568
rect 254 572 260 573
rect 254 568 255 572
rect 259 568 260 572
rect 254 567 260 568
rect 302 572 308 573
rect 302 568 303 572
rect 307 568 308 572
rect 302 567 308 568
rect 350 572 356 573
rect 350 568 351 572
rect 355 568 356 572
rect 350 567 356 568
rect 398 572 404 573
rect 398 568 399 572
rect 403 568 404 572
rect 398 567 404 568
rect 438 572 444 573
rect 438 568 439 572
rect 443 568 444 572
rect 438 567 444 568
rect 486 572 492 573
rect 486 568 487 572
rect 491 568 492 572
rect 486 567 492 568
rect 534 572 540 573
rect 534 568 535 572
rect 539 568 540 572
rect 534 567 540 568
rect 582 572 588 573
rect 582 568 583 572
rect 587 568 588 572
rect 582 567 588 568
rect 630 572 636 573
rect 630 568 631 572
rect 635 568 636 572
rect 630 567 636 568
rect 678 572 684 573
rect 678 568 679 572
rect 683 568 684 572
rect 678 567 684 568
rect 726 572 732 573
rect 726 568 727 572
rect 731 568 732 572
rect 1094 571 1095 575
rect 1099 571 1100 575
rect 1094 570 1100 571
rect 726 567 732 568
rect 136 563 138 567
rect 176 563 178 567
rect 216 563 218 567
rect 256 563 258 567
rect 304 563 306 567
rect 352 563 354 567
rect 400 563 402 567
rect 440 563 442 567
rect 488 563 490 567
rect 536 563 538 567
rect 584 563 586 567
rect 632 563 634 567
rect 680 563 682 567
rect 728 563 730 567
rect 1096 563 1098 570
rect 1136 565 1138 585
rect 1160 573 1162 585
rect 1200 573 1202 585
rect 1240 573 1242 585
rect 1280 573 1282 585
rect 1320 573 1322 585
rect 1360 573 1362 585
rect 1416 573 1418 585
rect 1488 573 1490 585
rect 1568 573 1570 585
rect 1656 573 1658 585
rect 1752 573 1754 585
rect 1856 573 1858 585
rect 1968 573 1970 585
rect 2072 573 2074 585
rect 1158 572 1164 573
rect 1158 568 1159 572
rect 1163 568 1164 572
rect 1158 567 1164 568
rect 1198 572 1204 573
rect 1198 568 1199 572
rect 1203 568 1204 572
rect 1198 567 1204 568
rect 1238 572 1244 573
rect 1238 568 1239 572
rect 1243 568 1244 572
rect 1238 567 1244 568
rect 1278 572 1284 573
rect 1278 568 1279 572
rect 1283 568 1284 572
rect 1278 567 1284 568
rect 1318 572 1324 573
rect 1318 568 1319 572
rect 1323 568 1324 572
rect 1318 567 1324 568
rect 1358 572 1364 573
rect 1358 568 1359 572
rect 1363 568 1364 572
rect 1358 567 1364 568
rect 1414 572 1420 573
rect 1414 568 1415 572
rect 1419 568 1420 572
rect 1414 567 1420 568
rect 1486 572 1492 573
rect 1486 568 1487 572
rect 1491 568 1492 572
rect 1486 567 1492 568
rect 1566 572 1572 573
rect 1566 568 1567 572
rect 1571 568 1572 572
rect 1566 567 1572 568
rect 1654 572 1660 573
rect 1654 568 1655 572
rect 1659 568 1660 572
rect 1654 567 1660 568
rect 1750 572 1756 573
rect 1750 568 1751 572
rect 1755 568 1756 572
rect 1750 567 1756 568
rect 1854 572 1860 573
rect 1854 568 1855 572
rect 1859 568 1860 572
rect 1854 567 1860 568
rect 1966 572 1972 573
rect 1966 568 1967 572
rect 1971 568 1972 572
rect 1966 567 1972 568
rect 2070 572 2076 573
rect 2070 568 2071 572
rect 2075 568 2076 572
rect 2070 567 2076 568
rect 2120 565 2122 585
rect 1134 564 1140 565
rect 111 562 115 563
rect 111 557 115 558
rect 135 562 139 563
rect 135 557 139 558
rect 175 562 179 563
rect 175 557 179 558
rect 215 562 219 563
rect 215 557 219 558
rect 223 562 227 563
rect 223 557 227 558
rect 255 562 259 563
rect 255 557 259 558
rect 279 562 283 563
rect 279 557 283 558
rect 303 562 307 563
rect 303 557 307 558
rect 327 562 331 563
rect 327 557 331 558
rect 351 562 355 563
rect 351 557 355 558
rect 375 562 379 563
rect 375 557 379 558
rect 399 562 403 563
rect 399 557 403 558
rect 423 562 427 563
rect 423 557 427 558
rect 439 562 443 563
rect 439 557 443 558
rect 463 562 467 563
rect 463 557 467 558
rect 487 562 491 563
rect 487 557 491 558
rect 511 562 515 563
rect 511 557 515 558
rect 535 562 539 563
rect 535 557 539 558
rect 559 562 563 563
rect 559 557 563 558
rect 583 562 587 563
rect 583 557 587 558
rect 607 562 611 563
rect 607 557 611 558
rect 631 562 635 563
rect 631 557 635 558
rect 655 562 659 563
rect 655 557 659 558
rect 679 562 683 563
rect 679 557 683 558
rect 703 562 707 563
rect 703 557 707 558
rect 727 562 731 563
rect 727 557 731 558
rect 751 562 755 563
rect 751 557 755 558
rect 1095 562 1099 563
rect 1134 560 1135 564
rect 1139 560 1140 564
rect 1134 559 1140 560
rect 2118 564 2124 565
rect 2118 560 2119 564
rect 2123 560 2124 564
rect 2118 559 2124 560
rect 1095 557 1099 558
rect 112 554 114 557
rect 134 556 140 557
rect 110 553 116 554
rect 110 549 111 553
rect 115 549 116 553
rect 134 552 135 556
rect 139 552 140 556
rect 134 551 140 552
rect 174 556 180 557
rect 174 552 175 556
rect 179 552 180 556
rect 174 551 180 552
rect 222 556 228 557
rect 222 552 223 556
rect 227 552 228 556
rect 222 551 228 552
rect 278 556 284 557
rect 278 552 279 556
rect 283 552 284 556
rect 278 551 284 552
rect 326 556 332 557
rect 326 552 327 556
rect 331 552 332 556
rect 326 551 332 552
rect 374 556 380 557
rect 374 552 375 556
rect 379 552 380 556
rect 374 551 380 552
rect 422 556 428 557
rect 422 552 423 556
rect 427 552 428 556
rect 422 551 428 552
rect 462 556 468 557
rect 462 552 463 556
rect 467 552 468 556
rect 462 551 468 552
rect 510 556 516 557
rect 510 552 511 556
rect 515 552 516 556
rect 510 551 516 552
rect 558 556 564 557
rect 558 552 559 556
rect 563 552 564 556
rect 558 551 564 552
rect 606 556 612 557
rect 606 552 607 556
rect 611 552 612 556
rect 606 551 612 552
rect 654 556 660 557
rect 654 552 655 556
rect 659 552 660 556
rect 654 551 660 552
rect 702 556 708 557
rect 702 552 703 556
rect 707 552 708 556
rect 702 551 708 552
rect 750 556 756 557
rect 750 552 751 556
rect 755 552 756 556
rect 1096 554 1098 557
rect 750 551 756 552
rect 1094 553 1100 554
rect 110 548 116 549
rect 1094 549 1095 553
rect 1099 549 1100 553
rect 1094 548 1100 549
rect 1134 547 1140 548
rect 1134 543 1135 547
rect 1139 543 1140 547
rect 2118 547 2124 548
rect 1134 542 1140 543
rect 1158 544 1164 545
rect 110 536 116 537
rect 110 532 111 536
rect 115 532 116 536
rect 110 531 116 532
rect 1094 536 1100 537
rect 1094 532 1095 536
rect 1099 532 1100 536
rect 1136 535 1138 542
rect 1158 540 1159 544
rect 1163 540 1164 544
rect 1158 539 1164 540
rect 1198 544 1204 545
rect 1198 540 1199 544
rect 1203 540 1204 544
rect 1198 539 1204 540
rect 1238 544 1244 545
rect 1238 540 1239 544
rect 1243 540 1244 544
rect 1238 539 1244 540
rect 1278 544 1284 545
rect 1278 540 1279 544
rect 1283 540 1284 544
rect 1278 539 1284 540
rect 1318 544 1324 545
rect 1318 540 1319 544
rect 1323 540 1324 544
rect 1318 539 1324 540
rect 1358 544 1364 545
rect 1358 540 1359 544
rect 1363 540 1364 544
rect 1358 539 1364 540
rect 1414 544 1420 545
rect 1414 540 1415 544
rect 1419 540 1420 544
rect 1414 539 1420 540
rect 1486 544 1492 545
rect 1486 540 1487 544
rect 1491 540 1492 544
rect 1486 539 1492 540
rect 1566 544 1572 545
rect 1566 540 1567 544
rect 1571 540 1572 544
rect 1566 539 1572 540
rect 1654 544 1660 545
rect 1654 540 1655 544
rect 1659 540 1660 544
rect 1654 539 1660 540
rect 1750 544 1756 545
rect 1750 540 1751 544
rect 1755 540 1756 544
rect 1750 539 1756 540
rect 1854 544 1860 545
rect 1854 540 1855 544
rect 1859 540 1860 544
rect 1854 539 1860 540
rect 1966 544 1972 545
rect 1966 540 1967 544
rect 1971 540 1972 544
rect 1966 539 1972 540
rect 2070 544 2076 545
rect 2070 540 2071 544
rect 2075 540 2076 544
rect 2118 543 2119 547
rect 2123 543 2124 547
rect 2118 542 2124 543
rect 2070 539 2076 540
rect 1160 535 1162 539
rect 1200 535 1202 539
rect 1240 535 1242 539
rect 1280 535 1282 539
rect 1320 535 1322 539
rect 1360 535 1362 539
rect 1416 535 1418 539
rect 1488 535 1490 539
rect 1568 535 1570 539
rect 1656 535 1658 539
rect 1752 535 1754 539
rect 1856 535 1858 539
rect 1968 535 1970 539
rect 2072 535 2074 539
rect 2120 535 2122 542
rect 1094 531 1100 532
rect 1135 534 1139 535
rect 112 503 114 531
rect 134 528 140 529
rect 134 524 135 528
rect 139 524 140 528
rect 134 523 140 524
rect 174 528 180 529
rect 174 524 175 528
rect 179 524 180 528
rect 174 523 180 524
rect 222 528 228 529
rect 222 524 223 528
rect 227 524 228 528
rect 222 523 228 524
rect 278 528 284 529
rect 278 524 279 528
rect 283 524 284 528
rect 278 523 284 524
rect 326 528 332 529
rect 326 524 327 528
rect 331 524 332 528
rect 326 523 332 524
rect 374 528 380 529
rect 374 524 375 528
rect 379 524 380 528
rect 374 523 380 524
rect 422 528 428 529
rect 422 524 423 528
rect 427 524 428 528
rect 422 523 428 524
rect 462 528 468 529
rect 462 524 463 528
rect 467 524 468 528
rect 462 523 468 524
rect 510 528 516 529
rect 510 524 511 528
rect 515 524 516 528
rect 510 523 516 524
rect 558 528 564 529
rect 558 524 559 528
rect 563 524 564 528
rect 558 523 564 524
rect 606 528 612 529
rect 606 524 607 528
rect 611 524 612 528
rect 606 523 612 524
rect 654 528 660 529
rect 654 524 655 528
rect 659 524 660 528
rect 654 523 660 524
rect 702 528 708 529
rect 702 524 703 528
rect 707 524 708 528
rect 702 523 708 524
rect 750 528 756 529
rect 750 524 751 528
rect 755 524 756 528
rect 750 523 756 524
rect 136 503 138 523
rect 176 503 178 523
rect 224 503 226 523
rect 280 503 282 523
rect 328 503 330 523
rect 376 503 378 523
rect 424 503 426 523
rect 464 503 466 523
rect 512 503 514 523
rect 560 503 562 523
rect 608 503 610 523
rect 656 503 658 523
rect 704 503 706 523
rect 752 503 754 523
rect 1096 503 1098 531
rect 1135 529 1139 530
rect 1159 534 1163 535
rect 1159 529 1163 530
rect 1199 534 1203 535
rect 1199 529 1203 530
rect 1239 534 1243 535
rect 1239 529 1243 530
rect 1279 534 1283 535
rect 1279 529 1283 530
rect 1303 534 1307 535
rect 1303 529 1307 530
rect 1319 534 1323 535
rect 1319 529 1323 530
rect 1343 534 1347 535
rect 1343 529 1347 530
rect 1359 534 1363 535
rect 1359 529 1363 530
rect 1383 534 1387 535
rect 1383 529 1387 530
rect 1415 534 1419 535
rect 1415 529 1419 530
rect 1423 534 1427 535
rect 1423 529 1427 530
rect 1463 534 1467 535
rect 1463 529 1467 530
rect 1487 534 1491 535
rect 1487 529 1491 530
rect 1503 534 1507 535
rect 1503 529 1507 530
rect 1543 534 1547 535
rect 1543 529 1547 530
rect 1567 534 1571 535
rect 1567 529 1571 530
rect 1591 534 1595 535
rect 1591 529 1595 530
rect 1647 534 1651 535
rect 1647 529 1651 530
rect 1655 534 1659 535
rect 1655 529 1659 530
rect 1703 534 1707 535
rect 1703 529 1707 530
rect 1751 534 1755 535
rect 1751 529 1755 530
rect 1767 534 1771 535
rect 1767 529 1771 530
rect 1839 534 1843 535
rect 1839 529 1843 530
rect 1855 534 1859 535
rect 1855 529 1859 530
rect 1919 534 1923 535
rect 1919 529 1923 530
rect 1967 534 1971 535
rect 1967 529 1971 530
rect 2007 534 2011 535
rect 2007 529 2011 530
rect 2071 534 2075 535
rect 2071 529 2075 530
rect 2119 534 2123 535
rect 2119 529 2123 530
rect 1136 526 1138 529
rect 1302 528 1308 529
rect 1134 525 1140 526
rect 1134 521 1135 525
rect 1139 521 1140 525
rect 1302 524 1303 528
rect 1307 524 1308 528
rect 1302 523 1308 524
rect 1342 528 1348 529
rect 1342 524 1343 528
rect 1347 524 1348 528
rect 1342 523 1348 524
rect 1382 528 1388 529
rect 1382 524 1383 528
rect 1387 524 1388 528
rect 1382 523 1388 524
rect 1422 528 1428 529
rect 1422 524 1423 528
rect 1427 524 1428 528
rect 1422 523 1428 524
rect 1462 528 1468 529
rect 1462 524 1463 528
rect 1467 524 1468 528
rect 1462 523 1468 524
rect 1502 528 1508 529
rect 1502 524 1503 528
rect 1507 524 1508 528
rect 1502 523 1508 524
rect 1542 528 1548 529
rect 1542 524 1543 528
rect 1547 524 1548 528
rect 1542 523 1548 524
rect 1590 528 1596 529
rect 1590 524 1591 528
rect 1595 524 1596 528
rect 1590 523 1596 524
rect 1646 528 1652 529
rect 1646 524 1647 528
rect 1651 524 1652 528
rect 1646 523 1652 524
rect 1702 528 1708 529
rect 1702 524 1703 528
rect 1707 524 1708 528
rect 1702 523 1708 524
rect 1766 528 1772 529
rect 1766 524 1767 528
rect 1771 524 1772 528
rect 1766 523 1772 524
rect 1838 528 1844 529
rect 1838 524 1839 528
rect 1843 524 1844 528
rect 1838 523 1844 524
rect 1918 528 1924 529
rect 1918 524 1919 528
rect 1923 524 1924 528
rect 1918 523 1924 524
rect 2006 528 2012 529
rect 2006 524 2007 528
rect 2011 524 2012 528
rect 2006 523 2012 524
rect 2070 528 2076 529
rect 2070 524 2071 528
rect 2075 524 2076 528
rect 2120 526 2122 529
rect 2070 523 2076 524
rect 2118 525 2124 526
rect 1134 520 1140 521
rect 2118 521 2119 525
rect 2123 521 2124 525
rect 2118 520 2124 521
rect 1134 508 1140 509
rect 1134 504 1135 508
rect 1139 504 1140 508
rect 1134 503 1140 504
rect 2118 508 2124 509
rect 2118 504 2119 508
rect 2123 504 2124 508
rect 2118 503 2124 504
rect 111 502 115 503
rect 111 497 115 498
rect 135 502 139 503
rect 135 497 139 498
rect 175 502 179 503
rect 175 497 179 498
rect 223 502 227 503
rect 223 497 227 498
rect 231 502 235 503
rect 231 497 235 498
rect 279 502 283 503
rect 279 497 283 498
rect 295 502 299 503
rect 295 497 299 498
rect 327 502 331 503
rect 327 497 331 498
rect 359 502 363 503
rect 359 497 363 498
rect 375 502 379 503
rect 375 497 379 498
rect 423 502 427 503
rect 423 497 427 498
rect 463 502 467 503
rect 463 497 467 498
rect 479 502 483 503
rect 479 497 483 498
rect 511 502 515 503
rect 511 497 515 498
rect 535 502 539 503
rect 535 497 539 498
rect 559 502 563 503
rect 559 497 563 498
rect 591 502 595 503
rect 591 497 595 498
rect 607 502 611 503
rect 607 497 611 498
rect 639 502 643 503
rect 639 497 643 498
rect 655 502 659 503
rect 655 497 659 498
rect 687 502 691 503
rect 687 497 691 498
rect 703 502 707 503
rect 703 497 707 498
rect 735 502 739 503
rect 735 497 739 498
rect 751 502 755 503
rect 751 497 755 498
rect 791 502 795 503
rect 791 497 795 498
rect 847 502 851 503
rect 847 497 851 498
rect 1095 502 1099 503
rect 1095 497 1099 498
rect 112 477 114 497
rect 136 485 138 497
rect 176 485 178 497
rect 232 485 234 497
rect 296 485 298 497
rect 360 485 362 497
rect 424 485 426 497
rect 480 485 482 497
rect 536 485 538 497
rect 592 485 594 497
rect 640 485 642 497
rect 688 485 690 497
rect 736 485 738 497
rect 792 485 794 497
rect 848 485 850 497
rect 134 484 140 485
rect 134 480 135 484
rect 139 480 140 484
rect 134 479 140 480
rect 174 484 180 485
rect 174 480 175 484
rect 179 480 180 484
rect 174 479 180 480
rect 230 484 236 485
rect 230 480 231 484
rect 235 480 236 484
rect 230 479 236 480
rect 294 484 300 485
rect 294 480 295 484
rect 299 480 300 484
rect 294 479 300 480
rect 358 484 364 485
rect 358 480 359 484
rect 363 480 364 484
rect 358 479 364 480
rect 422 484 428 485
rect 422 480 423 484
rect 427 480 428 484
rect 422 479 428 480
rect 478 484 484 485
rect 478 480 479 484
rect 483 480 484 484
rect 478 479 484 480
rect 534 484 540 485
rect 534 480 535 484
rect 539 480 540 484
rect 534 479 540 480
rect 590 484 596 485
rect 590 480 591 484
rect 595 480 596 484
rect 590 479 596 480
rect 638 484 644 485
rect 638 480 639 484
rect 643 480 644 484
rect 638 479 644 480
rect 686 484 692 485
rect 686 480 687 484
rect 691 480 692 484
rect 686 479 692 480
rect 734 484 740 485
rect 734 480 735 484
rect 739 480 740 484
rect 734 479 740 480
rect 790 484 796 485
rect 790 480 791 484
rect 795 480 796 484
rect 790 479 796 480
rect 846 484 852 485
rect 846 480 847 484
rect 851 480 852 484
rect 846 479 852 480
rect 1096 477 1098 497
rect 1136 483 1138 503
rect 1302 500 1308 501
rect 1302 496 1303 500
rect 1307 496 1308 500
rect 1302 495 1308 496
rect 1342 500 1348 501
rect 1342 496 1343 500
rect 1347 496 1348 500
rect 1342 495 1348 496
rect 1382 500 1388 501
rect 1382 496 1383 500
rect 1387 496 1388 500
rect 1382 495 1388 496
rect 1422 500 1428 501
rect 1422 496 1423 500
rect 1427 496 1428 500
rect 1422 495 1428 496
rect 1462 500 1468 501
rect 1462 496 1463 500
rect 1467 496 1468 500
rect 1462 495 1468 496
rect 1502 500 1508 501
rect 1502 496 1503 500
rect 1507 496 1508 500
rect 1502 495 1508 496
rect 1542 500 1548 501
rect 1542 496 1543 500
rect 1547 496 1548 500
rect 1542 495 1548 496
rect 1590 500 1596 501
rect 1590 496 1591 500
rect 1595 496 1596 500
rect 1590 495 1596 496
rect 1646 500 1652 501
rect 1646 496 1647 500
rect 1651 496 1652 500
rect 1646 495 1652 496
rect 1702 500 1708 501
rect 1702 496 1703 500
rect 1707 496 1708 500
rect 1702 495 1708 496
rect 1766 500 1772 501
rect 1766 496 1767 500
rect 1771 496 1772 500
rect 1766 495 1772 496
rect 1838 500 1844 501
rect 1838 496 1839 500
rect 1843 496 1844 500
rect 1838 495 1844 496
rect 1918 500 1924 501
rect 1918 496 1919 500
rect 1923 496 1924 500
rect 1918 495 1924 496
rect 2006 500 2012 501
rect 2006 496 2007 500
rect 2011 496 2012 500
rect 2006 495 2012 496
rect 2070 500 2076 501
rect 2070 496 2071 500
rect 2075 496 2076 500
rect 2070 495 2076 496
rect 1304 483 1306 495
rect 1344 483 1346 495
rect 1384 483 1386 495
rect 1424 483 1426 495
rect 1464 483 1466 495
rect 1504 483 1506 495
rect 1544 483 1546 495
rect 1592 483 1594 495
rect 1648 483 1650 495
rect 1704 483 1706 495
rect 1768 483 1770 495
rect 1840 483 1842 495
rect 1920 483 1922 495
rect 2008 483 2010 495
rect 2072 483 2074 495
rect 2120 483 2122 503
rect 1135 482 1139 483
rect 1135 477 1139 478
rect 1295 482 1299 483
rect 1295 477 1299 478
rect 1303 482 1307 483
rect 1303 477 1307 478
rect 1335 482 1339 483
rect 1335 477 1339 478
rect 1343 482 1347 483
rect 1343 477 1347 478
rect 1375 482 1379 483
rect 1375 477 1379 478
rect 1383 482 1387 483
rect 1383 477 1387 478
rect 1423 482 1427 483
rect 1423 477 1427 478
rect 1463 482 1467 483
rect 1463 477 1467 478
rect 1471 482 1475 483
rect 1471 477 1475 478
rect 1503 482 1507 483
rect 1503 477 1507 478
rect 1527 482 1531 483
rect 1527 477 1531 478
rect 1543 482 1547 483
rect 1543 477 1547 478
rect 1583 482 1587 483
rect 1583 477 1587 478
rect 1591 482 1595 483
rect 1591 477 1595 478
rect 1647 482 1651 483
rect 1647 477 1651 478
rect 1703 482 1707 483
rect 1703 477 1707 478
rect 1719 482 1723 483
rect 1719 477 1723 478
rect 1767 482 1771 483
rect 1767 477 1771 478
rect 1807 482 1811 483
rect 1807 477 1811 478
rect 1839 482 1843 483
rect 1839 477 1843 478
rect 1895 482 1899 483
rect 1895 477 1899 478
rect 1919 482 1923 483
rect 1919 477 1923 478
rect 1991 482 1995 483
rect 1991 477 1995 478
rect 2007 482 2011 483
rect 2007 477 2011 478
rect 2071 482 2075 483
rect 2071 477 2075 478
rect 2119 482 2123 483
rect 2119 477 2123 478
rect 110 476 116 477
rect 110 472 111 476
rect 115 472 116 476
rect 110 471 116 472
rect 1094 476 1100 477
rect 1094 472 1095 476
rect 1099 472 1100 476
rect 1094 471 1100 472
rect 110 459 116 460
rect 110 455 111 459
rect 115 455 116 459
rect 1094 459 1100 460
rect 110 454 116 455
rect 134 456 140 457
rect 112 447 114 454
rect 134 452 135 456
rect 139 452 140 456
rect 134 451 140 452
rect 174 456 180 457
rect 174 452 175 456
rect 179 452 180 456
rect 174 451 180 452
rect 230 456 236 457
rect 230 452 231 456
rect 235 452 236 456
rect 230 451 236 452
rect 294 456 300 457
rect 294 452 295 456
rect 299 452 300 456
rect 294 451 300 452
rect 358 456 364 457
rect 358 452 359 456
rect 363 452 364 456
rect 358 451 364 452
rect 422 456 428 457
rect 422 452 423 456
rect 427 452 428 456
rect 422 451 428 452
rect 478 456 484 457
rect 478 452 479 456
rect 483 452 484 456
rect 478 451 484 452
rect 534 456 540 457
rect 534 452 535 456
rect 539 452 540 456
rect 534 451 540 452
rect 590 456 596 457
rect 590 452 591 456
rect 595 452 596 456
rect 590 451 596 452
rect 638 456 644 457
rect 638 452 639 456
rect 643 452 644 456
rect 638 451 644 452
rect 686 456 692 457
rect 686 452 687 456
rect 691 452 692 456
rect 686 451 692 452
rect 734 456 740 457
rect 734 452 735 456
rect 739 452 740 456
rect 734 451 740 452
rect 790 456 796 457
rect 790 452 791 456
rect 795 452 796 456
rect 790 451 796 452
rect 846 456 852 457
rect 846 452 847 456
rect 851 452 852 456
rect 1094 455 1095 459
rect 1099 455 1100 459
rect 1136 457 1138 477
rect 1296 465 1298 477
rect 1336 465 1338 477
rect 1376 465 1378 477
rect 1424 465 1426 477
rect 1472 465 1474 477
rect 1528 465 1530 477
rect 1584 465 1586 477
rect 1648 465 1650 477
rect 1720 465 1722 477
rect 1808 465 1810 477
rect 1896 465 1898 477
rect 1992 465 1994 477
rect 2072 465 2074 477
rect 1294 464 1300 465
rect 1294 460 1295 464
rect 1299 460 1300 464
rect 1294 459 1300 460
rect 1334 464 1340 465
rect 1334 460 1335 464
rect 1339 460 1340 464
rect 1334 459 1340 460
rect 1374 464 1380 465
rect 1374 460 1375 464
rect 1379 460 1380 464
rect 1374 459 1380 460
rect 1422 464 1428 465
rect 1422 460 1423 464
rect 1427 460 1428 464
rect 1422 459 1428 460
rect 1470 464 1476 465
rect 1470 460 1471 464
rect 1475 460 1476 464
rect 1470 459 1476 460
rect 1526 464 1532 465
rect 1526 460 1527 464
rect 1531 460 1532 464
rect 1526 459 1532 460
rect 1582 464 1588 465
rect 1582 460 1583 464
rect 1587 460 1588 464
rect 1582 459 1588 460
rect 1646 464 1652 465
rect 1646 460 1647 464
rect 1651 460 1652 464
rect 1646 459 1652 460
rect 1718 464 1724 465
rect 1718 460 1719 464
rect 1723 460 1724 464
rect 1718 459 1724 460
rect 1806 464 1812 465
rect 1806 460 1807 464
rect 1811 460 1812 464
rect 1806 459 1812 460
rect 1894 464 1900 465
rect 1894 460 1895 464
rect 1899 460 1900 464
rect 1894 459 1900 460
rect 1990 464 1996 465
rect 1990 460 1991 464
rect 1995 460 1996 464
rect 1990 459 1996 460
rect 2070 464 2076 465
rect 2070 460 2071 464
rect 2075 460 2076 464
rect 2070 459 2076 460
rect 2120 457 2122 477
rect 1094 454 1100 455
rect 1134 456 1140 457
rect 846 451 852 452
rect 136 447 138 451
rect 176 447 178 451
rect 232 447 234 451
rect 296 447 298 451
rect 360 447 362 451
rect 424 447 426 451
rect 480 447 482 451
rect 536 447 538 451
rect 592 447 594 451
rect 640 447 642 451
rect 688 447 690 451
rect 736 447 738 451
rect 792 447 794 451
rect 848 447 850 451
rect 1096 447 1098 454
rect 1134 452 1135 456
rect 1139 452 1140 456
rect 1134 451 1140 452
rect 2118 456 2124 457
rect 2118 452 2119 456
rect 2123 452 2124 456
rect 2118 451 2124 452
rect 111 446 115 447
rect 111 441 115 442
rect 135 446 139 447
rect 135 441 139 442
rect 175 446 179 447
rect 175 441 179 442
rect 215 446 219 447
rect 215 441 219 442
rect 231 446 235 447
rect 231 441 235 442
rect 263 446 267 447
rect 263 441 267 442
rect 295 446 299 447
rect 295 441 299 442
rect 327 446 331 447
rect 327 441 331 442
rect 359 446 363 447
rect 359 441 363 442
rect 391 446 395 447
rect 391 441 395 442
rect 423 446 427 447
rect 423 441 427 442
rect 463 446 467 447
rect 463 441 467 442
rect 479 446 483 447
rect 479 441 483 442
rect 535 446 539 447
rect 535 441 539 442
rect 591 446 595 447
rect 591 441 595 442
rect 607 446 611 447
rect 607 441 611 442
rect 639 446 643 447
rect 639 441 643 442
rect 679 446 683 447
rect 679 441 683 442
rect 687 446 691 447
rect 687 441 691 442
rect 735 446 739 447
rect 735 441 739 442
rect 743 446 747 447
rect 743 441 747 442
rect 791 446 795 447
rect 791 441 795 442
rect 807 446 811 447
rect 807 441 811 442
rect 847 446 851 447
rect 847 441 851 442
rect 871 446 875 447
rect 871 441 875 442
rect 943 446 947 447
rect 943 441 947 442
rect 1095 446 1099 447
rect 1095 441 1099 442
rect 112 438 114 441
rect 174 440 180 441
rect 110 437 116 438
rect 110 433 111 437
rect 115 433 116 437
rect 174 436 175 440
rect 179 436 180 440
rect 174 435 180 436
rect 214 440 220 441
rect 214 436 215 440
rect 219 436 220 440
rect 214 435 220 436
rect 262 440 268 441
rect 262 436 263 440
rect 267 436 268 440
rect 262 435 268 436
rect 326 440 332 441
rect 326 436 327 440
rect 331 436 332 440
rect 326 435 332 436
rect 390 440 396 441
rect 390 436 391 440
rect 395 436 396 440
rect 390 435 396 436
rect 462 440 468 441
rect 462 436 463 440
rect 467 436 468 440
rect 462 435 468 436
rect 534 440 540 441
rect 534 436 535 440
rect 539 436 540 440
rect 534 435 540 436
rect 606 440 612 441
rect 606 436 607 440
rect 611 436 612 440
rect 606 435 612 436
rect 678 440 684 441
rect 678 436 679 440
rect 683 436 684 440
rect 678 435 684 436
rect 742 440 748 441
rect 742 436 743 440
rect 747 436 748 440
rect 742 435 748 436
rect 806 440 812 441
rect 806 436 807 440
rect 811 436 812 440
rect 806 435 812 436
rect 870 440 876 441
rect 870 436 871 440
rect 875 436 876 440
rect 870 435 876 436
rect 942 440 948 441
rect 942 436 943 440
rect 947 436 948 440
rect 1096 438 1098 441
rect 1134 439 1140 440
rect 942 435 948 436
rect 1094 437 1100 438
rect 110 432 116 433
rect 1094 433 1095 437
rect 1099 433 1100 437
rect 1134 435 1135 439
rect 1139 435 1140 439
rect 2118 439 2124 440
rect 1134 434 1140 435
rect 1294 436 1300 437
rect 1094 432 1100 433
rect 1136 431 1138 434
rect 1294 432 1295 436
rect 1299 432 1300 436
rect 1294 431 1300 432
rect 1334 436 1340 437
rect 1334 432 1335 436
rect 1339 432 1340 436
rect 1334 431 1340 432
rect 1374 436 1380 437
rect 1374 432 1375 436
rect 1379 432 1380 436
rect 1374 431 1380 432
rect 1422 436 1428 437
rect 1422 432 1423 436
rect 1427 432 1428 436
rect 1422 431 1428 432
rect 1470 436 1476 437
rect 1470 432 1471 436
rect 1475 432 1476 436
rect 1470 431 1476 432
rect 1526 436 1532 437
rect 1526 432 1527 436
rect 1531 432 1532 436
rect 1526 431 1532 432
rect 1582 436 1588 437
rect 1582 432 1583 436
rect 1587 432 1588 436
rect 1582 431 1588 432
rect 1646 436 1652 437
rect 1646 432 1647 436
rect 1651 432 1652 436
rect 1646 431 1652 432
rect 1718 436 1724 437
rect 1718 432 1719 436
rect 1723 432 1724 436
rect 1718 431 1724 432
rect 1806 436 1812 437
rect 1806 432 1807 436
rect 1811 432 1812 436
rect 1806 431 1812 432
rect 1894 436 1900 437
rect 1894 432 1895 436
rect 1899 432 1900 436
rect 1894 431 1900 432
rect 1990 436 1996 437
rect 1990 432 1991 436
rect 1995 432 1996 436
rect 1990 431 1996 432
rect 2070 436 2076 437
rect 2070 432 2071 436
rect 2075 432 2076 436
rect 2118 435 2119 439
rect 2123 435 2124 439
rect 2118 434 2124 435
rect 2070 431 2076 432
rect 2120 431 2122 434
rect 1135 430 1139 431
rect 1135 425 1139 426
rect 1159 430 1163 431
rect 1159 425 1163 426
rect 1199 430 1203 431
rect 1199 425 1203 426
rect 1255 430 1259 431
rect 1255 425 1259 426
rect 1295 430 1299 431
rect 1295 425 1299 426
rect 1335 430 1339 431
rect 1335 425 1339 426
rect 1375 430 1379 431
rect 1375 425 1379 426
rect 1415 430 1419 431
rect 1415 425 1419 426
rect 1423 430 1427 431
rect 1423 425 1427 426
rect 1471 430 1475 431
rect 1471 425 1475 426
rect 1503 430 1507 431
rect 1503 425 1507 426
rect 1527 430 1531 431
rect 1527 425 1531 426
rect 1583 430 1587 431
rect 1583 425 1587 426
rect 1591 430 1595 431
rect 1591 425 1595 426
rect 1647 430 1651 431
rect 1647 425 1651 426
rect 1671 430 1675 431
rect 1671 425 1675 426
rect 1719 430 1723 431
rect 1719 425 1723 426
rect 1751 430 1755 431
rect 1751 425 1755 426
rect 1807 430 1811 431
rect 1807 425 1811 426
rect 1831 430 1835 431
rect 1831 425 1835 426
rect 1895 430 1899 431
rect 1895 425 1899 426
rect 1911 430 1915 431
rect 1911 425 1915 426
rect 1991 430 1995 431
rect 1991 425 1995 426
rect 1999 430 2003 431
rect 1999 425 2003 426
rect 2071 430 2075 431
rect 2071 425 2075 426
rect 2119 430 2123 431
rect 2119 425 2123 426
rect 1136 422 1138 425
rect 1158 424 1164 425
rect 1134 421 1140 422
rect 110 420 116 421
rect 110 416 111 420
rect 115 416 116 420
rect 110 415 116 416
rect 1094 420 1100 421
rect 1094 416 1095 420
rect 1099 416 1100 420
rect 1134 417 1135 421
rect 1139 417 1140 421
rect 1158 420 1159 424
rect 1163 420 1164 424
rect 1158 419 1164 420
rect 1198 424 1204 425
rect 1198 420 1199 424
rect 1203 420 1204 424
rect 1198 419 1204 420
rect 1254 424 1260 425
rect 1254 420 1255 424
rect 1259 420 1260 424
rect 1254 419 1260 420
rect 1334 424 1340 425
rect 1334 420 1335 424
rect 1339 420 1340 424
rect 1334 419 1340 420
rect 1414 424 1420 425
rect 1414 420 1415 424
rect 1419 420 1420 424
rect 1414 419 1420 420
rect 1502 424 1508 425
rect 1502 420 1503 424
rect 1507 420 1508 424
rect 1502 419 1508 420
rect 1590 424 1596 425
rect 1590 420 1591 424
rect 1595 420 1596 424
rect 1590 419 1596 420
rect 1670 424 1676 425
rect 1670 420 1671 424
rect 1675 420 1676 424
rect 1670 419 1676 420
rect 1750 424 1756 425
rect 1750 420 1751 424
rect 1755 420 1756 424
rect 1750 419 1756 420
rect 1830 424 1836 425
rect 1830 420 1831 424
rect 1835 420 1836 424
rect 1830 419 1836 420
rect 1910 424 1916 425
rect 1910 420 1911 424
rect 1915 420 1916 424
rect 1910 419 1916 420
rect 1998 424 2004 425
rect 1998 420 1999 424
rect 2003 420 2004 424
rect 1998 419 2004 420
rect 2070 424 2076 425
rect 2070 420 2071 424
rect 2075 420 2076 424
rect 2120 422 2122 425
rect 2070 419 2076 420
rect 2118 421 2124 422
rect 1134 416 1140 417
rect 2118 417 2119 421
rect 2123 417 2124 421
rect 2118 416 2124 417
rect 1094 415 1100 416
rect 112 387 114 415
rect 174 412 180 413
rect 174 408 175 412
rect 179 408 180 412
rect 174 407 180 408
rect 214 412 220 413
rect 214 408 215 412
rect 219 408 220 412
rect 214 407 220 408
rect 262 412 268 413
rect 262 408 263 412
rect 267 408 268 412
rect 262 407 268 408
rect 326 412 332 413
rect 326 408 327 412
rect 331 408 332 412
rect 326 407 332 408
rect 390 412 396 413
rect 390 408 391 412
rect 395 408 396 412
rect 390 407 396 408
rect 462 412 468 413
rect 462 408 463 412
rect 467 408 468 412
rect 462 407 468 408
rect 534 412 540 413
rect 534 408 535 412
rect 539 408 540 412
rect 534 407 540 408
rect 606 412 612 413
rect 606 408 607 412
rect 611 408 612 412
rect 606 407 612 408
rect 678 412 684 413
rect 678 408 679 412
rect 683 408 684 412
rect 678 407 684 408
rect 742 412 748 413
rect 742 408 743 412
rect 747 408 748 412
rect 742 407 748 408
rect 806 412 812 413
rect 806 408 807 412
rect 811 408 812 412
rect 806 407 812 408
rect 870 412 876 413
rect 870 408 871 412
rect 875 408 876 412
rect 870 407 876 408
rect 942 412 948 413
rect 942 408 943 412
rect 947 408 948 412
rect 942 407 948 408
rect 176 387 178 407
rect 216 387 218 407
rect 264 387 266 407
rect 328 387 330 407
rect 392 387 394 407
rect 464 387 466 407
rect 536 387 538 407
rect 608 387 610 407
rect 680 387 682 407
rect 744 387 746 407
rect 808 387 810 407
rect 872 387 874 407
rect 944 387 946 407
rect 1096 387 1098 415
rect 1134 404 1140 405
rect 1134 400 1135 404
rect 1139 400 1140 404
rect 1134 399 1140 400
rect 2118 404 2124 405
rect 2118 400 2119 404
rect 2123 400 2124 404
rect 2118 399 2124 400
rect 111 386 115 387
rect 111 381 115 382
rect 175 386 179 387
rect 175 381 179 382
rect 215 386 219 387
rect 215 381 219 382
rect 263 386 267 387
rect 263 381 267 382
rect 271 386 275 387
rect 271 381 275 382
rect 327 386 331 387
rect 327 381 331 382
rect 335 386 339 387
rect 335 381 339 382
rect 391 386 395 387
rect 391 381 395 382
rect 407 386 411 387
rect 407 381 411 382
rect 463 386 467 387
rect 463 381 467 382
rect 487 386 491 387
rect 487 381 491 382
rect 535 386 539 387
rect 535 381 539 382
rect 567 386 571 387
rect 567 381 571 382
rect 607 386 611 387
rect 607 381 611 382
rect 639 386 643 387
rect 639 381 643 382
rect 679 386 683 387
rect 679 381 683 382
rect 711 386 715 387
rect 711 381 715 382
rect 743 386 747 387
rect 743 381 747 382
rect 775 386 779 387
rect 775 381 779 382
rect 807 386 811 387
rect 807 381 811 382
rect 839 386 843 387
rect 839 381 843 382
rect 871 386 875 387
rect 871 381 875 382
rect 895 386 899 387
rect 895 381 899 382
rect 943 386 947 387
rect 943 381 947 382
rect 951 386 955 387
rect 951 381 955 382
rect 1007 386 1011 387
rect 1007 381 1011 382
rect 1047 386 1051 387
rect 1047 381 1051 382
rect 1095 386 1099 387
rect 1095 381 1099 382
rect 112 361 114 381
rect 176 369 178 381
rect 216 369 218 381
rect 272 369 274 381
rect 336 369 338 381
rect 408 369 410 381
rect 488 369 490 381
rect 568 369 570 381
rect 640 369 642 381
rect 712 369 714 381
rect 776 369 778 381
rect 840 369 842 381
rect 896 369 898 381
rect 952 369 954 381
rect 1008 369 1010 381
rect 1048 369 1050 381
rect 174 368 180 369
rect 174 364 175 368
rect 179 364 180 368
rect 174 363 180 364
rect 214 368 220 369
rect 214 364 215 368
rect 219 364 220 368
rect 214 363 220 364
rect 270 368 276 369
rect 270 364 271 368
rect 275 364 276 368
rect 270 363 276 364
rect 334 368 340 369
rect 334 364 335 368
rect 339 364 340 368
rect 334 363 340 364
rect 406 368 412 369
rect 406 364 407 368
rect 411 364 412 368
rect 406 363 412 364
rect 486 368 492 369
rect 486 364 487 368
rect 491 364 492 368
rect 486 363 492 364
rect 566 368 572 369
rect 566 364 567 368
rect 571 364 572 368
rect 566 363 572 364
rect 638 368 644 369
rect 638 364 639 368
rect 643 364 644 368
rect 638 363 644 364
rect 710 368 716 369
rect 710 364 711 368
rect 715 364 716 368
rect 710 363 716 364
rect 774 368 780 369
rect 774 364 775 368
rect 779 364 780 368
rect 774 363 780 364
rect 838 368 844 369
rect 838 364 839 368
rect 843 364 844 368
rect 838 363 844 364
rect 894 368 900 369
rect 894 364 895 368
rect 899 364 900 368
rect 894 363 900 364
rect 950 368 956 369
rect 950 364 951 368
rect 955 364 956 368
rect 950 363 956 364
rect 1006 368 1012 369
rect 1006 364 1007 368
rect 1011 364 1012 368
rect 1006 363 1012 364
rect 1046 368 1052 369
rect 1046 364 1047 368
rect 1051 364 1052 368
rect 1046 363 1052 364
rect 1096 361 1098 381
rect 1136 375 1138 399
rect 1158 396 1164 397
rect 1158 392 1159 396
rect 1163 392 1164 396
rect 1158 391 1164 392
rect 1198 396 1204 397
rect 1198 392 1199 396
rect 1203 392 1204 396
rect 1198 391 1204 392
rect 1254 396 1260 397
rect 1254 392 1255 396
rect 1259 392 1260 396
rect 1254 391 1260 392
rect 1334 396 1340 397
rect 1334 392 1335 396
rect 1339 392 1340 396
rect 1334 391 1340 392
rect 1414 396 1420 397
rect 1414 392 1415 396
rect 1419 392 1420 396
rect 1414 391 1420 392
rect 1502 396 1508 397
rect 1502 392 1503 396
rect 1507 392 1508 396
rect 1502 391 1508 392
rect 1590 396 1596 397
rect 1590 392 1591 396
rect 1595 392 1596 396
rect 1590 391 1596 392
rect 1670 396 1676 397
rect 1670 392 1671 396
rect 1675 392 1676 396
rect 1670 391 1676 392
rect 1750 396 1756 397
rect 1750 392 1751 396
rect 1755 392 1756 396
rect 1750 391 1756 392
rect 1830 396 1836 397
rect 1830 392 1831 396
rect 1835 392 1836 396
rect 1830 391 1836 392
rect 1910 396 1916 397
rect 1910 392 1911 396
rect 1915 392 1916 396
rect 1910 391 1916 392
rect 1998 396 2004 397
rect 1998 392 1999 396
rect 2003 392 2004 396
rect 1998 391 2004 392
rect 2070 396 2076 397
rect 2070 392 2071 396
rect 2075 392 2076 396
rect 2070 391 2076 392
rect 1160 375 1162 391
rect 1200 375 1202 391
rect 1256 375 1258 391
rect 1336 375 1338 391
rect 1416 375 1418 391
rect 1504 375 1506 391
rect 1592 375 1594 391
rect 1672 375 1674 391
rect 1752 375 1754 391
rect 1832 375 1834 391
rect 1912 375 1914 391
rect 2000 375 2002 391
rect 2072 375 2074 391
rect 2120 375 2122 399
rect 1135 374 1139 375
rect 1135 369 1139 370
rect 1159 374 1163 375
rect 1159 369 1163 370
rect 1199 374 1203 375
rect 1199 369 1203 370
rect 1247 374 1251 375
rect 1247 369 1251 370
rect 1255 374 1259 375
rect 1255 369 1259 370
rect 1335 374 1339 375
rect 1335 369 1339 370
rect 1359 374 1363 375
rect 1359 369 1363 370
rect 1415 374 1419 375
rect 1415 369 1419 370
rect 1463 374 1467 375
rect 1463 369 1467 370
rect 1503 374 1507 375
rect 1503 369 1507 370
rect 1559 374 1563 375
rect 1559 369 1563 370
rect 1591 374 1595 375
rect 1591 369 1595 370
rect 1647 374 1651 375
rect 1647 369 1651 370
rect 1671 374 1675 375
rect 1671 369 1675 370
rect 1727 374 1731 375
rect 1727 369 1731 370
rect 1751 374 1755 375
rect 1751 369 1755 370
rect 1799 374 1803 375
rect 1799 369 1803 370
rect 1831 374 1835 375
rect 1831 369 1835 370
rect 1863 374 1867 375
rect 1863 369 1867 370
rect 1911 374 1915 375
rect 1911 369 1915 370
rect 1919 374 1923 375
rect 1919 369 1923 370
rect 1975 374 1979 375
rect 1975 369 1979 370
rect 1999 374 2003 375
rect 1999 369 2003 370
rect 2031 374 2035 375
rect 2031 369 2035 370
rect 2071 374 2075 375
rect 2071 369 2075 370
rect 2119 374 2123 375
rect 2119 369 2123 370
rect 110 360 116 361
rect 110 356 111 360
rect 115 356 116 360
rect 110 355 116 356
rect 1094 360 1100 361
rect 1094 356 1095 360
rect 1099 356 1100 360
rect 1094 355 1100 356
rect 1136 349 1138 369
rect 1160 357 1162 369
rect 1248 357 1250 369
rect 1360 357 1362 369
rect 1464 357 1466 369
rect 1560 357 1562 369
rect 1648 357 1650 369
rect 1728 357 1730 369
rect 1800 357 1802 369
rect 1864 357 1866 369
rect 1920 357 1922 369
rect 1976 357 1978 369
rect 2032 357 2034 369
rect 2072 357 2074 369
rect 1158 356 1164 357
rect 1158 352 1159 356
rect 1163 352 1164 356
rect 1158 351 1164 352
rect 1246 356 1252 357
rect 1246 352 1247 356
rect 1251 352 1252 356
rect 1246 351 1252 352
rect 1358 356 1364 357
rect 1358 352 1359 356
rect 1363 352 1364 356
rect 1358 351 1364 352
rect 1462 356 1468 357
rect 1462 352 1463 356
rect 1467 352 1468 356
rect 1462 351 1468 352
rect 1558 356 1564 357
rect 1558 352 1559 356
rect 1563 352 1564 356
rect 1558 351 1564 352
rect 1646 356 1652 357
rect 1646 352 1647 356
rect 1651 352 1652 356
rect 1646 351 1652 352
rect 1726 356 1732 357
rect 1726 352 1727 356
rect 1731 352 1732 356
rect 1726 351 1732 352
rect 1798 356 1804 357
rect 1798 352 1799 356
rect 1803 352 1804 356
rect 1798 351 1804 352
rect 1862 356 1868 357
rect 1862 352 1863 356
rect 1867 352 1868 356
rect 1862 351 1868 352
rect 1918 356 1924 357
rect 1918 352 1919 356
rect 1923 352 1924 356
rect 1918 351 1924 352
rect 1974 356 1980 357
rect 1974 352 1975 356
rect 1979 352 1980 356
rect 1974 351 1980 352
rect 2030 356 2036 357
rect 2030 352 2031 356
rect 2035 352 2036 356
rect 2030 351 2036 352
rect 2070 356 2076 357
rect 2070 352 2071 356
rect 2075 352 2076 356
rect 2070 351 2076 352
rect 2120 349 2122 369
rect 1134 348 1140 349
rect 1134 344 1135 348
rect 1139 344 1140 348
rect 110 343 116 344
rect 110 339 111 343
rect 115 339 116 343
rect 1094 343 1100 344
rect 1134 343 1140 344
rect 2118 348 2124 349
rect 2118 344 2119 348
rect 2123 344 2124 348
rect 2118 343 2124 344
rect 110 338 116 339
rect 174 340 180 341
rect 112 331 114 338
rect 174 336 175 340
rect 179 336 180 340
rect 174 335 180 336
rect 214 340 220 341
rect 214 336 215 340
rect 219 336 220 340
rect 214 335 220 336
rect 270 340 276 341
rect 270 336 271 340
rect 275 336 276 340
rect 270 335 276 336
rect 334 340 340 341
rect 334 336 335 340
rect 339 336 340 340
rect 334 335 340 336
rect 406 340 412 341
rect 406 336 407 340
rect 411 336 412 340
rect 406 335 412 336
rect 486 340 492 341
rect 486 336 487 340
rect 491 336 492 340
rect 486 335 492 336
rect 566 340 572 341
rect 566 336 567 340
rect 571 336 572 340
rect 566 335 572 336
rect 638 340 644 341
rect 638 336 639 340
rect 643 336 644 340
rect 638 335 644 336
rect 710 340 716 341
rect 710 336 711 340
rect 715 336 716 340
rect 710 335 716 336
rect 774 340 780 341
rect 774 336 775 340
rect 779 336 780 340
rect 774 335 780 336
rect 838 340 844 341
rect 838 336 839 340
rect 843 336 844 340
rect 838 335 844 336
rect 894 340 900 341
rect 894 336 895 340
rect 899 336 900 340
rect 894 335 900 336
rect 950 340 956 341
rect 950 336 951 340
rect 955 336 956 340
rect 950 335 956 336
rect 1006 340 1012 341
rect 1006 336 1007 340
rect 1011 336 1012 340
rect 1006 335 1012 336
rect 1046 340 1052 341
rect 1046 336 1047 340
rect 1051 336 1052 340
rect 1094 339 1095 343
rect 1099 339 1100 343
rect 1094 338 1100 339
rect 1046 335 1052 336
rect 176 331 178 335
rect 216 331 218 335
rect 272 331 274 335
rect 336 331 338 335
rect 408 331 410 335
rect 488 331 490 335
rect 568 331 570 335
rect 640 331 642 335
rect 712 331 714 335
rect 776 331 778 335
rect 840 331 842 335
rect 896 331 898 335
rect 952 331 954 335
rect 1008 331 1010 335
rect 1048 331 1050 335
rect 1096 331 1098 338
rect 1134 331 1140 332
rect 111 330 115 331
rect 111 325 115 326
rect 175 330 179 331
rect 175 325 179 326
rect 215 330 219 331
rect 215 325 219 326
rect 271 330 275 331
rect 271 325 275 326
rect 335 330 339 331
rect 335 325 339 326
rect 383 330 387 331
rect 383 325 387 326
rect 407 330 411 331
rect 407 325 411 326
rect 423 330 427 331
rect 423 325 427 326
rect 463 330 467 331
rect 463 325 467 326
rect 487 330 491 331
rect 487 325 491 326
rect 503 330 507 331
rect 503 325 507 326
rect 543 330 547 331
rect 543 325 547 326
rect 567 330 571 331
rect 567 325 571 326
rect 591 330 595 331
rect 591 325 595 326
rect 639 330 643 331
rect 639 325 643 326
rect 687 330 691 331
rect 687 325 691 326
rect 711 330 715 331
rect 711 325 715 326
rect 735 330 739 331
rect 735 325 739 326
rect 775 330 779 331
rect 775 325 779 326
rect 783 330 787 331
rect 783 325 787 326
rect 831 330 835 331
rect 831 325 835 326
rect 839 330 843 331
rect 839 325 843 326
rect 879 330 883 331
rect 879 325 883 326
rect 895 330 899 331
rect 895 325 899 326
rect 927 330 931 331
rect 927 325 931 326
rect 951 330 955 331
rect 951 325 955 326
rect 967 330 971 331
rect 967 325 971 326
rect 1007 330 1011 331
rect 1007 325 1011 326
rect 1047 330 1051 331
rect 1047 325 1051 326
rect 1095 330 1099 331
rect 1134 327 1135 331
rect 1139 327 1140 331
rect 2118 331 2124 332
rect 1134 326 1140 327
rect 1158 328 1164 329
rect 1095 325 1099 326
rect 112 322 114 325
rect 382 324 388 325
rect 110 321 116 322
rect 110 317 111 321
rect 115 317 116 321
rect 382 320 383 324
rect 387 320 388 324
rect 382 319 388 320
rect 422 324 428 325
rect 422 320 423 324
rect 427 320 428 324
rect 422 319 428 320
rect 462 324 468 325
rect 462 320 463 324
rect 467 320 468 324
rect 462 319 468 320
rect 502 324 508 325
rect 502 320 503 324
rect 507 320 508 324
rect 502 319 508 320
rect 542 324 548 325
rect 542 320 543 324
rect 547 320 548 324
rect 542 319 548 320
rect 590 324 596 325
rect 590 320 591 324
rect 595 320 596 324
rect 590 319 596 320
rect 638 324 644 325
rect 638 320 639 324
rect 643 320 644 324
rect 638 319 644 320
rect 686 324 692 325
rect 686 320 687 324
rect 691 320 692 324
rect 686 319 692 320
rect 734 324 740 325
rect 734 320 735 324
rect 739 320 740 324
rect 734 319 740 320
rect 782 324 788 325
rect 782 320 783 324
rect 787 320 788 324
rect 782 319 788 320
rect 830 324 836 325
rect 830 320 831 324
rect 835 320 836 324
rect 830 319 836 320
rect 878 324 884 325
rect 878 320 879 324
rect 883 320 884 324
rect 878 319 884 320
rect 926 324 932 325
rect 926 320 927 324
rect 931 320 932 324
rect 926 319 932 320
rect 966 324 972 325
rect 966 320 967 324
rect 971 320 972 324
rect 966 319 972 320
rect 1006 324 1012 325
rect 1006 320 1007 324
rect 1011 320 1012 324
rect 1006 319 1012 320
rect 1046 324 1052 325
rect 1046 320 1047 324
rect 1051 320 1052 324
rect 1096 322 1098 325
rect 1046 319 1052 320
rect 1094 321 1100 322
rect 110 316 116 317
rect 1094 317 1095 321
rect 1099 317 1100 321
rect 1094 316 1100 317
rect 1136 315 1138 326
rect 1158 324 1159 328
rect 1163 324 1164 328
rect 1158 323 1164 324
rect 1246 328 1252 329
rect 1246 324 1247 328
rect 1251 324 1252 328
rect 1246 323 1252 324
rect 1358 328 1364 329
rect 1358 324 1359 328
rect 1363 324 1364 328
rect 1358 323 1364 324
rect 1462 328 1468 329
rect 1462 324 1463 328
rect 1467 324 1468 328
rect 1462 323 1468 324
rect 1558 328 1564 329
rect 1558 324 1559 328
rect 1563 324 1564 328
rect 1558 323 1564 324
rect 1646 328 1652 329
rect 1646 324 1647 328
rect 1651 324 1652 328
rect 1646 323 1652 324
rect 1726 328 1732 329
rect 1726 324 1727 328
rect 1731 324 1732 328
rect 1726 323 1732 324
rect 1798 328 1804 329
rect 1798 324 1799 328
rect 1803 324 1804 328
rect 1798 323 1804 324
rect 1862 328 1868 329
rect 1862 324 1863 328
rect 1867 324 1868 328
rect 1862 323 1868 324
rect 1918 328 1924 329
rect 1918 324 1919 328
rect 1923 324 1924 328
rect 1918 323 1924 324
rect 1974 328 1980 329
rect 1974 324 1975 328
rect 1979 324 1980 328
rect 1974 323 1980 324
rect 2030 328 2036 329
rect 2030 324 2031 328
rect 2035 324 2036 328
rect 2030 323 2036 324
rect 2070 328 2076 329
rect 2070 324 2071 328
rect 2075 324 2076 328
rect 2118 327 2119 331
rect 2123 327 2124 331
rect 2118 326 2124 327
rect 2070 323 2076 324
rect 1160 315 1162 323
rect 1248 315 1250 323
rect 1360 315 1362 323
rect 1464 315 1466 323
rect 1560 315 1562 323
rect 1648 315 1650 323
rect 1728 315 1730 323
rect 1800 315 1802 323
rect 1864 315 1866 323
rect 1920 315 1922 323
rect 1976 315 1978 323
rect 2032 315 2034 323
rect 2072 315 2074 323
rect 2120 315 2122 326
rect 1135 314 1139 315
rect 1135 309 1139 310
rect 1159 314 1163 315
rect 1159 309 1163 310
rect 1247 314 1251 315
rect 1247 309 1251 310
rect 1351 314 1355 315
rect 1351 309 1355 310
rect 1359 314 1363 315
rect 1359 309 1363 310
rect 1391 314 1395 315
rect 1391 309 1395 310
rect 1431 314 1435 315
rect 1431 309 1435 310
rect 1463 314 1467 315
rect 1463 309 1467 310
rect 1471 314 1475 315
rect 1471 309 1475 310
rect 1511 314 1515 315
rect 1511 309 1515 310
rect 1559 314 1563 315
rect 1559 309 1563 310
rect 1615 314 1619 315
rect 1615 309 1619 310
rect 1647 314 1651 315
rect 1647 309 1651 310
rect 1671 314 1675 315
rect 1671 309 1675 310
rect 1727 314 1731 315
rect 1727 309 1731 310
rect 1735 314 1739 315
rect 1735 309 1739 310
rect 1799 314 1803 315
rect 1799 309 1803 310
rect 1807 314 1811 315
rect 1807 309 1811 310
rect 1863 314 1867 315
rect 1863 309 1867 310
rect 1887 314 1891 315
rect 1887 309 1891 310
rect 1919 314 1923 315
rect 1919 309 1923 310
rect 1967 314 1971 315
rect 1967 309 1971 310
rect 1975 314 1979 315
rect 1975 309 1979 310
rect 2031 314 2035 315
rect 2031 309 2035 310
rect 2047 314 2051 315
rect 2047 309 2051 310
rect 2071 314 2075 315
rect 2071 309 2075 310
rect 2119 314 2123 315
rect 2119 309 2123 310
rect 1136 306 1138 309
rect 1350 308 1356 309
rect 1134 305 1140 306
rect 110 304 116 305
rect 110 300 111 304
rect 115 300 116 304
rect 110 299 116 300
rect 1094 304 1100 305
rect 1094 300 1095 304
rect 1099 300 1100 304
rect 1134 301 1135 305
rect 1139 301 1140 305
rect 1350 304 1351 308
rect 1355 304 1356 308
rect 1350 303 1356 304
rect 1390 308 1396 309
rect 1390 304 1391 308
rect 1395 304 1396 308
rect 1390 303 1396 304
rect 1430 308 1436 309
rect 1430 304 1431 308
rect 1435 304 1436 308
rect 1430 303 1436 304
rect 1470 308 1476 309
rect 1470 304 1471 308
rect 1475 304 1476 308
rect 1470 303 1476 304
rect 1510 308 1516 309
rect 1510 304 1511 308
rect 1515 304 1516 308
rect 1510 303 1516 304
rect 1558 308 1564 309
rect 1558 304 1559 308
rect 1563 304 1564 308
rect 1558 303 1564 304
rect 1614 308 1620 309
rect 1614 304 1615 308
rect 1619 304 1620 308
rect 1614 303 1620 304
rect 1670 308 1676 309
rect 1670 304 1671 308
rect 1675 304 1676 308
rect 1670 303 1676 304
rect 1734 308 1740 309
rect 1734 304 1735 308
rect 1739 304 1740 308
rect 1734 303 1740 304
rect 1806 308 1812 309
rect 1806 304 1807 308
rect 1811 304 1812 308
rect 1806 303 1812 304
rect 1886 308 1892 309
rect 1886 304 1887 308
rect 1891 304 1892 308
rect 1886 303 1892 304
rect 1966 308 1972 309
rect 1966 304 1967 308
rect 1971 304 1972 308
rect 1966 303 1972 304
rect 2046 308 2052 309
rect 2046 304 2047 308
rect 2051 304 2052 308
rect 2120 306 2122 309
rect 2046 303 2052 304
rect 2118 305 2124 306
rect 1134 300 1140 301
rect 2118 301 2119 305
rect 2123 301 2124 305
rect 2118 300 2124 301
rect 1094 299 1100 300
rect 112 271 114 299
rect 382 296 388 297
rect 382 292 383 296
rect 387 292 388 296
rect 382 291 388 292
rect 422 296 428 297
rect 422 292 423 296
rect 427 292 428 296
rect 422 291 428 292
rect 462 296 468 297
rect 462 292 463 296
rect 467 292 468 296
rect 462 291 468 292
rect 502 296 508 297
rect 502 292 503 296
rect 507 292 508 296
rect 502 291 508 292
rect 542 296 548 297
rect 542 292 543 296
rect 547 292 548 296
rect 542 291 548 292
rect 590 296 596 297
rect 590 292 591 296
rect 595 292 596 296
rect 590 291 596 292
rect 638 296 644 297
rect 638 292 639 296
rect 643 292 644 296
rect 638 291 644 292
rect 686 296 692 297
rect 686 292 687 296
rect 691 292 692 296
rect 686 291 692 292
rect 734 296 740 297
rect 734 292 735 296
rect 739 292 740 296
rect 734 291 740 292
rect 782 296 788 297
rect 782 292 783 296
rect 787 292 788 296
rect 782 291 788 292
rect 830 296 836 297
rect 830 292 831 296
rect 835 292 836 296
rect 830 291 836 292
rect 878 296 884 297
rect 878 292 879 296
rect 883 292 884 296
rect 878 291 884 292
rect 926 296 932 297
rect 926 292 927 296
rect 931 292 932 296
rect 926 291 932 292
rect 966 296 972 297
rect 966 292 967 296
rect 971 292 972 296
rect 966 291 972 292
rect 1006 296 1012 297
rect 1006 292 1007 296
rect 1011 292 1012 296
rect 1006 291 1012 292
rect 1046 296 1052 297
rect 1046 292 1047 296
rect 1051 292 1052 296
rect 1046 291 1052 292
rect 384 271 386 291
rect 424 271 426 291
rect 464 271 466 291
rect 504 271 506 291
rect 544 271 546 291
rect 592 271 594 291
rect 640 271 642 291
rect 688 271 690 291
rect 736 271 738 291
rect 784 271 786 291
rect 832 271 834 291
rect 880 271 882 291
rect 928 271 930 291
rect 968 271 970 291
rect 1008 271 1010 291
rect 1048 271 1050 291
rect 1096 271 1098 299
rect 1134 288 1140 289
rect 1134 284 1135 288
rect 1139 284 1140 288
rect 1134 283 1140 284
rect 2118 288 2124 289
rect 2118 284 2119 288
rect 2123 284 2124 288
rect 2118 283 2124 284
rect 111 270 115 271
rect 111 265 115 266
rect 287 270 291 271
rect 287 265 291 266
rect 327 270 331 271
rect 327 265 331 266
rect 367 270 371 271
rect 367 265 371 266
rect 383 270 387 271
rect 383 265 387 266
rect 415 270 419 271
rect 415 265 419 266
rect 423 270 427 271
rect 423 265 427 266
rect 463 270 467 271
rect 463 265 467 266
rect 471 270 475 271
rect 471 265 475 266
rect 503 270 507 271
rect 503 265 507 266
rect 535 270 539 271
rect 535 265 539 266
rect 543 270 547 271
rect 543 265 547 266
rect 591 270 595 271
rect 591 265 595 266
rect 607 270 611 271
rect 607 265 611 266
rect 639 270 643 271
rect 639 265 643 266
rect 679 270 683 271
rect 679 265 683 266
rect 687 270 691 271
rect 687 265 691 266
rect 735 270 739 271
rect 735 265 739 266
rect 743 270 747 271
rect 743 265 747 266
rect 783 270 787 271
rect 783 265 787 266
rect 807 270 811 271
rect 807 265 811 266
rect 831 270 835 271
rect 831 265 835 266
rect 863 270 867 271
rect 863 265 867 266
rect 879 270 883 271
rect 879 265 883 266
rect 927 270 931 271
rect 927 265 931 266
rect 967 270 971 271
rect 967 265 971 266
rect 991 270 995 271
rect 991 265 995 266
rect 1007 270 1011 271
rect 1007 265 1011 266
rect 1047 270 1051 271
rect 1047 265 1051 266
rect 1095 270 1099 271
rect 1095 265 1099 266
rect 112 245 114 265
rect 288 253 290 265
rect 328 253 330 265
rect 368 253 370 265
rect 416 253 418 265
rect 472 253 474 265
rect 536 253 538 265
rect 608 253 610 265
rect 680 253 682 265
rect 744 253 746 265
rect 808 253 810 265
rect 864 253 866 265
rect 928 253 930 265
rect 992 253 994 265
rect 1048 253 1050 265
rect 286 252 292 253
rect 286 248 287 252
rect 291 248 292 252
rect 286 247 292 248
rect 326 252 332 253
rect 326 248 327 252
rect 331 248 332 252
rect 326 247 332 248
rect 366 252 372 253
rect 366 248 367 252
rect 371 248 372 252
rect 366 247 372 248
rect 414 252 420 253
rect 414 248 415 252
rect 419 248 420 252
rect 414 247 420 248
rect 470 252 476 253
rect 470 248 471 252
rect 475 248 476 252
rect 470 247 476 248
rect 534 252 540 253
rect 534 248 535 252
rect 539 248 540 252
rect 534 247 540 248
rect 606 252 612 253
rect 606 248 607 252
rect 611 248 612 252
rect 606 247 612 248
rect 678 252 684 253
rect 678 248 679 252
rect 683 248 684 252
rect 678 247 684 248
rect 742 252 748 253
rect 742 248 743 252
rect 747 248 748 252
rect 742 247 748 248
rect 806 252 812 253
rect 806 248 807 252
rect 811 248 812 252
rect 806 247 812 248
rect 862 252 868 253
rect 862 248 863 252
rect 867 248 868 252
rect 862 247 868 248
rect 926 252 932 253
rect 926 248 927 252
rect 931 248 932 252
rect 926 247 932 248
rect 990 252 996 253
rect 990 248 991 252
rect 995 248 996 252
rect 990 247 996 248
rect 1046 252 1052 253
rect 1046 248 1047 252
rect 1051 248 1052 252
rect 1046 247 1052 248
rect 1096 245 1098 265
rect 1136 263 1138 283
rect 1350 280 1356 281
rect 1350 276 1351 280
rect 1355 276 1356 280
rect 1350 275 1356 276
rect 1390 280 1396 281
rect 1390 276 1391 280
rect 1395 276 1396 280
rect 1390 275 1396 276
rect 1430 280 1436 281
rect 1430 276 1431 280
rect 1435 276 1436 280
rect 1430 275 1436 276
rect 1470 280 1476 281
rect 1470 276 1471 280
rect 1475 276 1476 280
rect 1470 275 1476 276
rect 1510 280 1516 281
rect 1510 276 1511 280
rect 1515 276 1516 280
rect 1510 275 1516 276
rect 1558 280 1564 281
rect 1558 276 1559 280
rect 1563 276 1564 280
rect 1558 275 1564 276
rect 1614 280 1620 281
rect 1614 276 1615 280
rect 1619 276 1620 280
rect 1614 275 1620 276
rect 1670 280 1676 281
rect 1670 276 1671 280
rect 1675 276 1676 280
rect 1670 275 1676 276
rect 1734 280 1740 281
rect 1734 276 1735 280
rect 1739 276 1740 280
rect 1734 275 1740 276
rect 1806 280 1812 281
rect 1806 276 1807 280
rect 1811 276 1812 280
rect 1806 275 1812 276
rect 1886 280 1892 281
rect 1886 276 1887 280
rect 1891 276 1892 280
rect 1886 275 1892 276
rect 1966 280 1972 281
rect 1966 276 1967 280
rect 1971 276 1972 280
rect 1966 275 1972 276
rect 2046 280 2052 281
rect 2046 276 2047 280
rect 2051 276 2052 280
rect 2046 275 2052 276
rect 1352 263 1354 275
rect 1392 263 1394 275
rect 1432 263 1434 275
rect 1472 263 1474 275
rect 1512 263 1514 275
rect 1560 263 1562 275
rect 1616 263 1618 275
rect 1672 263 1674 275
rect 1736 263 1738 275
rect 1808 263 1810 275
rect 1888 263 1890 275
rect 1968 263 1970 275
rect 2048 263 2050 275
rect 2120 263 2122 283
rect 1135 262 1139 263
rect 1135 257 1139 258
rect 1263 262 1267 263
rect 1263 257 1267 258
rect 1303 262 1307 263
rect 1303 257 1307 258
rect 1343 262 1347 263
rect 1343 257 1347 258
rect 1351 262 1355 263
rect 1351 257 1355 258
rect 1383 262 1387 263
rect 1383 257 1387 258
rect 1391 262 1395 263
rect 1391 257 1395 258
rect 1423 262 1427 263
rect 1423 257 1427 258
rect 1431 262 1435 263
rect 1431 257 1435 258
rect 1463 262 1467 263
rect 1463 257 1467 258
rect 1471 262 1475 263
rect 1471 257 1475 258
rect 1503 262 1507 263
rect 1503 257 1507 258
rect 1511 262 1515 263
rect 1511 257 1515 258
rect 1543 262 1547 263
rect 1543 257 1547 258
rect 1559 262 1563 263
rect 1559 257 1563 258
rect 1599 262 1603 263
rect 1599 257 1603 258
rect 1615 262 1619 263
rect 1615 257 1619 258
rect 1671 262 1675 263
rect 1671 257 1675 258
rect 1735 262 1739 263
rect 1735 257 1739 258
rect 1759 262 1763 263
rect 1759 257 1763 258
rect 1807 262 1811 263
rect 1807 257 1811 258
rect 1863 262 1867 263
rect 1863 257 1867 258
rect 1887 262 1891 263
rect 1887 257 1891 258
rect 1967 262 1971 263
rect 1967 257 1971 258
rect 1975 262 1979 263
rect 1975 257 1979 258
rect 2047 262 2051 263
rect 2047 257 2051 258
rect 2071 262 2075 263
rect 2071 257 2075 258
rect 2119 262 2123 263
rect 2119 257 2123 258
rect 110 244 116 245
rect 110 240 111 244
rect 115 240 116 244
rect 110 239 116 240
rect 1094 244 1100 245
rect 1094 240 1095 244
rect 1099 240 1100 244
rect 1094 239 1100 240
rect 1136 237 1138 257
rect 1264 245 1266 257
rect 1304 245 1306 257
rect 1344 245 1346 257
rect 1384 245 1386 257
rect 1424 245 1426 257
rect 1464 245 1466 257
rect 1504 245 1506 257
rect 1544 245 1546 257
rect 1600 245 1602 257
rect 1672 245 1674 257
rect 1760 245 1762 257
rect 1864 245 1866 257
rect 1976 245 1978 257
rect 2072 245 2074 257
rect 1262 244 1268 245
rect 1262 240 1263 244
rect 1267 240 1268 244
rect 1262 239 1268 240
rect 1302 244 1308 245
rect 1302 240 1303 244
rect 1307 240 1308 244
rect 1302 239 1308 240
rect 1342 244 1348 245
rect 1342 240 1343 244
rect 1347 240 1348 244
rect 1342 239 1348 240
rect 1382 244 1388 245
rect 1382 240 1383 244
rect 1387 240 1388 244
rect 1382 239 1388 240
rect 1422 244 1428 245
rect 1422 240 1423 244
rect 1427 240 1428 244
rect 1422 239 1428 240
rect 1462 244 1468 245
rect 1462 240 1463 244
rect 1467 240 1468 244
rect 1462 239 1468 240
rect 1502 244 1508 245
rect 1502 240 1503 244
rect 1507 240 1508 244
rect 1502 239 1508 240
rect 1542 244 1548 245
rect 1542 240 1543 244
rect 1547 240 1548 244
rect 1542 239 1548 240
rect 1598 244 1604 245
rect 1598 240 1599 244
rect 1603 240 1604 244
rect 1598 239 1604 240
rect 1670 244 1676 245
rect 1670 240 1671 244
rect 1675 240 1676 244
rect 1670 239 1676 240
rect 1758 244 1764 245
rect 1758 240 1759 244
rect 1763 240 1764 244
rect 1758 239 1764 240
rect 1862 244 1868 245
rect 1862 240 1863 244
rect 1867 240 1868 244
rect 1862 239 1868 240
rect 1974 244 1980 245
rect 1974 240 1975 244
rect 1979 240 1980 244
rect 1974 239 1980 240
rect 2070 244 2076 245
rect 2070 240 2071 244
rect 2075 240 2076 244
rect 2070 239 2076 240
rect 2120 237 2122 257
rect 1134 236 1140 237
rect 1134 232 1135 236
rect 1139 232 1140 236
rect 1134 231 1140 232
rect 2118 236 2124 237
rect 2118 232 2119 236
rect 2123 232 2124 236
rect 2118 231 2124 232
rect 110 227 116 228
rect 110 223 111 227
rect 115 223 116 227
rect 1094 227 1100 228
rect 110 222 116 223
rect 286 224 292 225
rect 112 207 114 222
rect 286 220 287 224
rect 291 220 292 224
rect 286 219 292 220
rect 326 224 332 225
rect 326 220 327 224
rect 331 220 332 224
rect 326 219 332 220
rect 366 224 372 225
rect 366 220 367 224
rect 371 220 372 224
rect 366 219 372 220
rect 414 224 420 225
rect 414 220 415 224
rect 419 220 420 224
rect 414 219 420 220
rect 470 224 476 225
rect 470 220 471 224
rect 475 220 476 224
rect 470 219 476 220
rect 534 224 540 225
rect 534 220 535 224
rect 539 220 540 224
rect 534 219 540 220
rect 606 224 612 225
rect 606 220 607 224
rect 611 220 612 224
rect 606 219 612 220
rect 678 224 684 225
rect 678 220 679 224
rect 683 220 684 224
rect 678 219 684 220
rect 742 224 748 225
rect 742 220 743 224
rect 747 220 748 224
rect 742 219 748 220
rect 806 224 812 225
rect 806 220 807 224
rect 811 220 812 224
rect 806 219 812 220
rect 862 224 868 225
rect 862 220 863 224
rect 867 220 868 224
rect 862 219 868 220
rect 926 224 932 225
rect 926 220 927 224
rect 931 220 932 224
rect 926 219 932 220
rect 990 224 996 225
rect 990 220 991 224
rect 995 220 996 224
rect 990 219 996 220
rect 1046 224 1052 225
rect 1046 220 1047 224
rect 1051 220 1052 224
rect 1094 223 1095 227
rect 1099 223 1100 227
rect 1094 222 1100 223
rect 1046 219 1052 220
rect 288 207 290 219
rect 328 207 330 219
rect 368 207 370 219
rect 416 207 418 219
rect 472 207 474 219
rect 536 207 538 219
rect 608 207 610 219
rect 680 207 682 219
rect 744 207 746 219
rect 808 207 810 219
rect 864 207 866 219
rect 928 207 930 219
rect 992 207 994 219
rect 1048 207 1050 219
rect 1096 207 1098 222
rect 1134 219 1140 220
rect 1134 215 1135 219
rect 1139 215 1140 219
rect 2118 219 2124 220
rect 1134 214 1140 215
rect 1262 216 1268 217
rect 1136 207 1138 214
rect 1262 212 1263 216
rect 1267 212 1268 216
rect 1262 211 1268 212
rect 1302 216 1308 217
rect 1302 212 1303 216
rect 1307 212 1308 216
rect 1302 211 1308 212
rect 1342 216 1348 217
rect 1342 212 1343 216
rect 1347 212 1348 216
rect 1342 211 1348 212
rect 1382 216 1388 217
rect 1382 212 1383 216
rect 1387 212 1388 216
rect 1382 211 1388 212
rect 1422 216 1428 217
rect 1422 212 1423 216
rect 1427 212 1428 216
rect 1422 211 1428 212
rect 1462 216 1468 217
rect 1462 212 1463 216
rect 1467 212 1468 216
rect 1462 211 1468 212
rect 1502 216 1508 217
rect 1502 212 1503 216
rect 1507 212 1508 216
rect 1502 211 1508 212
rect 1542 216 1548 217
rect 1542 212 1543 216
rect 1547 212 1548 216
rect 1542 211 1548 212
rect 1598 216 1604 217
rect 1598 212 1599 216
rect 1603 212 1604 216
rect 1598 211 1604 212
rect 1670 216 1676 217
rect 1670 212 1671 216
rect 1675 212 1676 216
rect 1670 211 1676 212
rect 1758 216 1764 217
rect 1758 212 1759 216
rect 1763 212 1764 216
rect 1758 211 1764 212
rect 1862 216 1868 217
rect 1862 212 1863 216
rect 1867 212 1868 216
rect 1862 211 1868 212
rect 1974 216 1980 217
rect 1974 212 1975 216
rect 1979 212 1980 216
rect 1974 211 1980 212
rect 2070 216 2076 217
rect 2070 212 2071 216
rect 2075 212 2076 216
rect 2118 215 2119 219
rect 2123 215 2124 219
rect 2118 214 2124 215
rect 2070 211 2076 212
rect 1264 207 1266 211
rect 1304 207 1306 211
rect 1344 207 1346 211
rect 1384 207 1386 211
rect 1424 207 1426 211
rect 1464 207 1466 211
rect 1504 207 1506 211
rect 1544 207 1546 211
rect 1600 207 1602 211
rect 1672 207 1674 211
rect 1760 207 1762 211
rect 1864 207 1866 211
rect 1976 207 1978 211
rect 2072 207 2074 211
rect 2120 207 2122 214
rect 111 206 115 207
rect 111 201 115 202
rect 167 206 171 207
rect 167 201 171 202
rect 207 206 211 207
rect 207 201 211 202
rect 247 206 251 207
rect 247 201 251 202
rect 287 206 291 207
rect 287 201 291 202
rect 295 206 299 207
rect 295 201 299 202
rect 327 206 331 207
rect 327 201 331 202
rect 343 206 347 207
rect 343 201 347 202
rect 367 206 371 207
rect 367 201 371 202
rect 399 206 403 207
rect 399 201 403 202
rect 415 206 419 207
rect 415 201 419 202
rect 463 206 467 207
rect 463 201 467 202
rect 471 206 475 207
rect 471 201 475 202
rect 527 206 531 207
rect 527 201 531 202
rect 535 206 539 207
rect 535 201 539 202
rect 599 206 603 207
rect 599 201 603 202
rect 607 206 611 207
rect 607 201 611 202
rect 671 206 675 207
rect 671 201 675 202
rect 679 206 683 207
rect 679 201 683 202
rect 743 206 747 207
rect 743 201 747 202
rect 751 206 755 207
rect 751 201 755 202
rect 807 206 811 207
rect 807 201 811 202
rect 831 206 835 207
rect 831 201 835 202
rect 863 206 867 207
rect 863 201 867 202
rect 911 206 915 207
rect 911 201 915 202
rect 927 206 931 207
rect 927 201 931 202
rect 991 206 995 207
rect 991 201 995 202
rect 1047 206 1051 207
rect 1047 201 1051 202
rect 1095 206 1099 207
rect 1095 201 1099 202
rect 1135 206 1139 207
rect 1135 201 1139 202
rect 1183 206 1187 207
rect 1183 201 1187 202
rect 1231 206 1235 207
rect 1231 201 1235 202
rect 1263 206 1267 207
rect 1263 201 1267 202
rect 1295 206 1299 207
rect 1295 201 1299 202
rect 1303 206 1307 207
rect 1303 201 1307 202
rect 1343 206 1347 207
rect 1343 201 1347 202
rect 1359 206 1363 207
rect 1359 201 1363 202
rect 1383 206 1387 207
rect 1383 201 1387 202
rect 1423 206 1427 207
rect 1423 201 1427 202
rect 1431 206 1435 207
rect 1431 201 1435 202
rect 1463 206 1467 207
rect 1463 201 1467 202
rect 1503 206 1507 207
rect 1503 201 1507 202
rect 1511 206 1515 207
rect 1511 201 1515 202
rect 1543 206 1547 207
rect 1543 201 1547 202
rect 1591 206 1595 207
rect 1591 201 1595 202
rect 1599 206 1603 207
rect 1599 201 1603 202
rect 1663 206 1667 207
rect 1663 201 1667 202
rect 1671 206 1675 207
rect 1671 201 1675 202
rect 1735 206 1739 207
rect 1735 201 1739 202
rect 1759 206 1763 207
rect 1759 201 1763 202
rect 1807 206 1811 207
rect 1807 201 1811 202
rect 1863 206 1867 207
rect 1863 201 1867 202
rect 1879 206 1883 207
rect 1879 201 1883 202
rect 1951 206 1955 207
rect 1951 201 1955 202
rect 1975 206 1979 207
rect 1975 201 1979 202
rect 2023 206 2027 207
rect 2023 201 2027 202
rect 2071 206 2075 207
rect 2071 201 2075 202
rect 2119 206 2123 207
rect 2119 201 2123 202
rect 112 198 114 201
rect 166 200 172 201
rect 110 197 116 198
rect 110 193 111 197
rect 115 193 116 197
rect 166 196 167 200
rect 171 196 172 200
rect 166 195 172 196
rect 206 200 212 201
rect 206 196 207 200
rect 211 196 212 200
rect 206 195 212 196
rect 246 200 252 201
rect 246 196 247 200
rect 251 196 252 200
rect 246 195 252 196
rect 294 200 300 201
rect 294 196 295 200
rect 299 196 300 200
rect 294 195 300 196
rect 342 200 348 201
rect 342 196 343 200
rect 347 196 348 200
rect 342 195 348 196
rect 398 200 404 201
rect 398 196 399 200
rect 403 196 404 200
rect 398 195 404 196
rect 462 200 468 201
rect 462 196 463 200
rect 467 196 468 200
rect 462 195 468 196
rect 526 200 532 201
rect 526 196 527 200
rect 531 196 532 200
rect 526 195 532 196
rect 598 200 604 201
rect 598 196 599 200
rect 603 196 604 200
rect 598 195 604 196
rect 670 200 676 201
rect 670 196 671 200
rect 675 196 676 200
rect 670 195 676 196
rect 750 200 756 201
rect 750 196 751 200
rect 755 196 756 200
rect 750 195 756 196
rect 830 200 836 201
rect 830 196 831 200
rect 835 196 836 200
rect 830 195 836 196
rect 910 200 916 201
rect 910 196 911 200
rect 915 196 916 200
rect 910 195 916 196
rect 990 200 996 201
rect 990 196 991 200
rect 995 196 996 200
rect 990 195 996 196
rect 1046 200 1052 201
rect 1046 196 1047 200
rect 1051 196 1052 200
rect 1096 198 1098 201
rect 1136 198 1138 201
rect 1182 200 1188 201
rect 1046 195 1052 196
rect 1094 197 1100 198
rect 110 192 116 193
rect 1094 193 1095 197
rect 1099 193 1100 197
rect 1094 192 1100 193
rect 1134 197 1140 198
rect 1134 193 1135 197
rect 1139 193 1140 197
rect 1182 196 1183 200
rect 1187 196 1188 200
rect 1182 195 1188 196
rect 1230 200 1236 201
rect 1230 196 1231 200
rect 1235 196 1236 200
rect 1230 195 1236 196
rect 1294 200 1300 201
rect 1294 196 1295 200
rect 1299 196 1300 200
rect 1294 195 1300 196
rect 1358 200 1364 201
rect 1358 196 1359 200
rect 1363 196 1364 200
rect 1358 195 1364 196
rect 1430 200 1436 201
rect 1430 196 1431 200
rect 1435 196 1436 200
rect 1430 195 1436 196
rect 1510 200 1516 201
rect 1510 196 1511 200
rect 1515 196 1516 200
rect 1510 195 1516 196
rect 1590 200 1596 201
rect 1590 196 1591 200
rect 1595 196 1596 200
rect 1590 195 1596 196
rect 1662 200 1668 201
rect 1662 196 1663 200
rect 1667 196 1668 200
rect 1662 195 1668 196
rect 1734 200 1740 201
rect 1734 196 1735 200
rect 1739 196 1740 200
rect 1734 195 1740 196
rect 1806 200 1812 201
rect 1806 196 1807 200
rect 1811 196 1812 200
rect 1806 195 1812 196
rect 1878 200 1884 201
rect 1878 196 1879 200
rect 1883 196 1884 200
rect 1878 195 1884 196
rect 1950 200 1956 201
rect 1950 196 1951 200
rect 1955 196 1956 200
rect 1950 195 1956 196
rect 2022 200 2028 201
rect 2022 196 2023 200
rect 2027 196 2028 200
rect 2022 195 2028 196
rect 2070 200 2076 201
rect 2070 196 2071 200
rect 2075 196 2076 200
rect 2120 198 2122 201
rect 2070 195 2076 196
rect 2118 197 2124 198
rect 1134 192 1140 193
rect 2118 193 2119 197
rect 2123 193 2124 197
rect 2118 192 2124 193
rect 110 180 116 181
rect 110 176 111 180
rect 115 176 116 180
rect 110 175 116 176
rect 1094 180 1100 181
rect 1094 176 1095 180
rect 1099 176 1100 180
rect 1094 175 1100 176
rect 1134 180 1140 181
rect 1134 176 1135 180
rect 1139 176 1140 180
rect 1134 175 1140 176
rect 2118 180 2124 181
rect 2118 176 2119 180
rect 2123 176 2124 180
rect 2118 175 2124 176
rect 112 139 114 175
rect 166 172 172 173
rect 166 168 167 172
rect 171 168 172 172
rect 166 167 172 168
rect 206 172 212 173
rect 206 168 207 172
rect 211 168 212 172
rect 206 167 212 168
rect 246 172 252 173
rect 246 168 247 172
rect 251 168 252 172
rect 246 167 252 168
rect 294 172 300 173
rect 294 168 295 172
rect 299 168 300 172
rect 294 167 300 168
rect 342 172 348 173
rect 342 168 343 172
rect 347 168 348 172
rect 342 167 348 168
rect 398 172 404 173
rect 398 168 399 172
rect 403 168 404 172
rect 398 167 404 168
rect 462 172 468 173
rect 462 168 463 172
rect 467 168 468 172
rect 462 167 468 168
rect 526 172 532 173
rect 526 168 527 172
rect 531 168 532 172
rect 526 167 532 168
rect 598 172 604 173
rect 598 168 599 172
rect 603 168 604 172
rect 598 167 604 168
rect 670 172 676 173
rect 670 168 671 172
rect 675 168 676 172
rect 670 167 676 168
rect 750 172 756 173
rect 750 168 751 172
rect 755 168 756 172
rect 750 167 756 168
rect 830 172 836 173
rect 830 168 831 172
rect 835 168 836 172
rect 830 167 836 168
rect 910 172 916 173
rect 910 168 911 172
rect 915 168 916 172
rect 910 167 916 168
rect 990 172 996 173
rect 990 168 991 172
rect 995 168 996 172
rect 990 167 996 168
rect 1046 172 1052 173
rect 1046 168 1047 172
rect 1051 168 1052 172
rect 1046 167 1052 168
rect 168 139 170 167
rect 208 139 210 167
rect 248 139 250 167
rect 296 139 298 167
rect 344 139 346 167
rect 400 139 402 167
rect 464 139 466 167
rect 528 139 530 167
rect 600 139 602 167
rect 672 139 674 167
rect 752 139 754 167
rect 832 139 834 167
rect 912 139 914 167
rect 992 139 994 167
rect 1048 139 1050 167
rect 1096 139 1098 175
rect 111 138 115 139
rect 111 133 115 134
rect 135 138 139 139
rect 135 133 139 134
rect 167 138 171 139
rect 167 133 171 134
rect 175 138 179 139
rect 175 133 179 134
rect 207 138 211 139
rect 207 133 211 134
rect 215 138 219 139
rect 215 133 219 134
rect 247 138 251 139
rect 247 133 251 134
rect 255 138 259 139
rect 255 133 259 134
rect 295 138 299 139
rect 295 133 299 134
rect 335 138 339 139
rect 335 133 339 134
rect 343 138 347 139
rect 343 133 347 134
rect 375 138 379 139
rect 375 133 379 134
rect 399 138 403 139
rect 399 133 403 134
rect 415 138 419 139
rect 415 133 419 134
rect 455 138 459 139
rect 455 133 459 134
rect 463 138 467 139
rect 463 133 467 134
rect 495 138 499 139
rect 495 133 499 134
rect 527 138 531 139
rect 527 133 531 134
rect 535 138 539 139
rect 535 133 539 134
rect 575 138 579 139
rect 575 133 579 134
rect 599 138 603 139
rect 599 133 603 134
rect 615 138 619 139
rect 615 133 619 134
rect 655 138 659 139
rect 655 133 659 134
rect 671 138 675 139
rect 671 133 675 134
rect 695 138 699 139
rect 695 133 699 134
rect 735 138 739 139
rect 735 133 739 134
rect 751 138 755 139
rect 751 133 755 134
rect 775 138 779 139
rect 775 133 779 134
rect 815 138 819 139
rect 815 133 819 134
rect 831 138 835 139
rect 831 133 835 134
rect 871 138 875 139
rect 871 133 875 134
rect 911 138 915 139
rect 911 133 915 134
rect 935 138 939 139
rect 935 133 939 134
rect 991 138 995 139
rect 991 133 995 134
rect 999 138 1003 139
rect 999 133 1003 134
rect 1047 138 1051 139
rect 1047 133 1051 134
rect 1095 138 1099 139
rect 1095 133 1099 134
rect 112 113 114 133
rect 136 121 138 133
rect 176 121 178 133
rect 216 121 218 133
rect 256 121 258 133
rect 296 121 298 133
rect 336 121 338 133
rect 376 121 378 133
rect 416 121 418 133
rect 456 121 458 133
rect 496 121 498 133
rect 536 121 538 133
rect 576 121 578 133
rect 616 121 618 133
rect 656 121 658 133
rect 696 121 698 133
rect 736 121 738 133
rect 776 121 778 133
rect 816 121 818 133
rect 872 121 874 133
rect 936 121 938 133
rect 1000 121 1002 133
rect 1048 121 1050 133
rect 134 120 140 121
rect 134 116 135 120
rect 139 116 140 120
rect 134 115 140 116
rect 174 120 180 121
rect 174 116 175 120
rect 179 116 180 120
rect 174 115 180 116
rect 214 120 220 121
rect 214 116 215 120
rect 219 116 220 120
rect 214 115 220 116
rect 254 120 260 121
rect 254 116 255 120
rect 259 116 260 120
rect 254 115 260 116
rect 294 120 300 121
rect 294 116 295 120
rect 299 116 300 120
rect 294 115 300 116
rect 334 120 340 121
rect 334 116 335 120
rect 339 116 340 120
rect 334 115 340 116
rect 374 120 380 121
rect 374 116 375 120
rect 379 116 380 120
rect 374 115 380 116
rect 414 120 420 121
rect 414 116 415 120
rect 419 116 420 120
rect 414 115 420 116
rect 454 120 460 121
rect 454 116 455 120
rect 459 116 460 120
rect 454 115 460 116
rect 494 120 500 121
rect 494 116 495 120
rect 499 116 500 120
rect 494 115 500 116
rect 534 120 540 121
rect 534 116 535 120
rect 539 116 540 120
rect 534 115 540 116
rect 574 120 580 121
rect 574 116 575 120
rect 579 116 580 120
rect 574 115 580 116
rect 614 120 620 121
rect 614 116 615 120
rect 619 116 620 120
rect 614 115 620 116
rect 654 120 660 121
rect 654 116 655 120
rect 659 116 660 120
rect 654 115 660 116
rect 694 120 700 121
rect 694 116 695 120
rect 699 116 700 120
rect 694 115 700 116
rect 734 120 740 121
rect 734 116 735 120
rect 739 116 740 120
rect 734 115 740 116
rect 774 120 780 121
rect 774 116 775 120
rect 779 116 780 120
rect 774 115 780 116
rect 814 120 820 121
rect 814 116 815 120
rect 819 116 820 120
rect 814 115 820 116
rect 870 120 876 121
rect 870 116 871 120
rect 875 116 876 120
rect 870 115 876 116
rect 934 120 940 121
rect 934 116 935 120
rect 939 116 940 120
rect 934 115 940 116
rect 998 120 1004 121
rect 998 116 999 120
rect 1003 116 1004 120
rect 998 115 1004 116
rect 1046 120 1052 121
rect 1046 116 1047 120
rect 1051 116 1052 120
rect 1046 115 1052 116
rect 1096 113 1098 133
rect 1136 131 1138 175
rect 1182 172 1188 173
rect 1182 168 1183 172
rect 1187 168 1188 172
rect 1182 167 1188 168
rect 1230 172 1236 173
rect 1230 168 1231 172
rect 1235 168 1236 172
rect 1230 167 1236 168
rect 1294 172 1300 173
rect 1294 168 1295 172
rect 1299 168 1300 172
rect 1294 167 1300 168
rect 1358 172 1364 173
rect 1358 168 1359 172
rect 1363 168 1364 172
rect 1358 167 1364 168
rect 1430 172 1436 173
rect 1430 168 1431 172
rect 1435 168 1436 172
rect 1430 167 1436 168
rect 1510 172 1516 173
rect 1510 168 1511 172
rect 1515 168 1516 172
rect 1510 167 1516 168
rect 1590 172 1596 173
rect 1590 168 1591 172
rect 1595 168 1596 172
rect 1590 167 1596 168
rect 1662 172 1668 173
rect 1662 168 1663 172
rect 1667 168 1668 172
rect 1662 167 1668 168
rect 1734 172 1740 173
rect 1734 168 1735 172
rect 1739 168 1740 172
rect 1734 167 1740 168
rect 1806 172 1812 173
rect 1806 168 1807 172
rect 1811 168 1812 172
rect 1806 167 1812 168
rect 1878 172 1884 173
rect 1878 168 1879 172
rect 1883 168 1884 172
rect 1878 167 1884 168
rect 1950 172 1956 173
rect 1950 168 1951 172
rect 1955 168 1956 172
rect 1950 167 1956 168
rect 2022 172 2028 173
rect 2022 168 2023 172
rect 2027 168 2028 172
rect 2022 167 2028 168
rect 2070 172 2076 173
rect 2070 168 2071 172
rect 2075 168 2076 172
rect 2070 167 2076 168
rect 1184 131 1186 167
rect 1232 131 1234 167
rect 1296 131 1298 167
rect 1360 131 1362 167
rect 1432 131 1434 167
rect 1512 131 1514 167
rect 1592 131 1594 167
rect 1664 131 1666 167
rect 1736 131 1738 167
rect 1808 131 1810 167
rect 1880 131 1882 167
rect 1952 131 1954 167
rect 2024 131 2026 167
rect 2072 131 2074 167
rect 2120 131 2122 175
rect 1135 130 1139 131
rect 1135 125 1139 126
rect 1159 130 1163 131
rect 1159 125 1163 126
rect 1183 130 1187 131
rect 1183 125 1187 126
rect 1199 130 1203 131
rect 1199 125 1203 126
rect 1231 130 1235 131
rect 1231 125 1235 126
rect 1239 130 1243 131
rect 1239 125 1243 126
rect 1279 130 1283 131
rect 1279 125 1283 126
rect 1295 130 1299 131
rect 1295 125 1299 126
rect 1319 130 1323 131
rect 1319 125 1323 126
rect 1359 130 1363 131
rect 1359 125 1363 126
rect 1367 130 1371 131
rect 1367 125 1371 126
rect 1431 130 1435 131
rect 1431 125 1435 126
rect 1495 130 1499 131
rect 1495 125 1499 126
rect 1511 130 1515 131
rect 1511 125 1515 126
rect 1559 130 1563 131
rect 1559 125 1563 126
rect 1591 130 1595 131
rect 1591 125 1595 126
rect 1615 130 1619 131
rect 1615 125 1619 126
rect 1663 130 1667 131
rect 1663 125 1667 126
rect 1671 130 1675 131
rect 1671 125 1675 126
rect 1719 130 1723 131
rect 1719 125 1723 126
rect 1735 130 1739 131
rect 1735 125 1739 126
rect 1767 130 1771 131
rect 1767 125 1771 126
rect 1807 130 1811 131
rect 1807 125 1811 126
rect 1855 130 1859 131
rect 1855 125 1859 126
rect 1879 130 1883 131
rect 1879 125 1883 126
rect 1903 130 1907 131
rect 1903 125 1907 126
rect 1951 130 1955 131
rect 1951 125 1955 126
rect 1991 130 1995 131
rect 1991 125 1995 126
rect 2023 130 2027 131
rect 2023 125 2027 126
rect 2031 130 2035 131
rect 2031 125 2035 126
rect 2071 130 2075 131
rect 2071 125 2075 126
rect 2119 130 2123 131
rect 2119 125 2123 126
rect 110 112 116 113
rect 110 108 111 112
rect 115 108 116 112
rect 110 107 116 108
rect 1094 112 1100 113
rect 1094 108 1095 112
rect 1099 108 1100 112
rect 1094 107 1100 108
rect 1136 105 1138 125
rect 1160 113 1162 125
rect 1200 113 1202 125
rect 1240 113 1242 125
rect 1280 113 1282 125
rect 1320 113 1322 125
rect 1368 113 1370 125
rect 1432 113 1434 125
rect 1496 113 1498 125
rect 1560 113 1562 125
rect 1616 113 1618 125
rect 1672 113 1674 125
rect 1720 113 1722 125
rect 1768 113 1770 125
rect 1808 113 1810 125
rect 1856 113 1858 125
rect 1904 113 1906 125
rect 1952 113 1954 125
rect 1992 113 1994 125
rect 2032 113 2034 125
rect 2072 113 2074 125
rect 1158 112 1164 113
rect 1158 108 1159 112
rect 1163 108 1164 112
rect 1158 107 1164 108
rect 1198 112 1204 113
rect 1198 108 1199 112
rect 1203 108 1204 112
rect 1198 107 1204 108
rect 1238 112 1244 113
rect 1238 108 1239 112
rect 1243 108 1244 112
rect 1238 107 1244 108
rect 1278 112 1284 113
rect 1278 108 1279 112
rect 1283 108 1284 112
rect 1278 107 1284 108
rect 1318 112 1324 113
rect 1318 108 1319 112
rect 1323 108 1324 112
rect 1318 107 1324 108
rect 1366 112 1372 113
rect 1366 108 1367 112
rect 1371 108 1372 112
rect 1366 107 1372 108
rect 1430 112 1436 113
rect 1430 108 1431 112
rect 1435 108 1436 112
rect 1430 107 1436 108
rect 1494 112 1500 113
rect 1494 108 1495 112
rect 1499 108 1500 112
rect 1494 107 1500 108
rect 1558 112 1564 113
rect 1558 108 1559 112
rect 1563 108 1564 112
rect 1558 107 1564 108
rect 1614 112 1620 113
rect 1614 108 1615 112
rect 1619 108 1620 112
rect 1614 107 1620 108
rect 1670 112 1676 113
rect 1670 108 1671 112
rect 1675 108 1676 112
rect 1670 107 1676 108
rect 1718 112 1724 113
rect 1718 108 1719 112
rect 1723 108 1724 112
rect 1718 107 1724 108
rect 1766 112 1772 113
rect 1766 108 1767 112
rect 1771 108 1772 112
rect 1766 107 1772 108
rect 1806 112 1812 113
rect 1806 108 1807 112
rect 1811 108 1812 112
rect 1806 107 1812 108
rect 1854 112 1860 113
rect 1854 108 1855 112
rect 1859 108 1860 112
rect 1854 107 1860 108
rect 1902 112 1908 113
rect 1902 108 1903 112
rect 1907 108 1908 112
rect 1902 107 1908 108
rect 1950 112 1956 113
rect 1950 108 1951 112
rect 1955 108 1956 112
rect 1950 107 1956 108
rect 1990 112 1996 113
rect 1990 108 1991 112
rect 1995 108 1996 112
rect 1990 107 1996 108
rect 2030 112 2036 113
rect 2030 108 2031 112
rect 2035 108 2036 112
rect 2030 107 2036 108
rect 2070 112 2076 113
rect 2070 108 2071 112
rect 2075 108 2076 112
rect 2070 107 2076 108
rect 2120 105 2122 125
rect 1134 104 1140 105
rect 1134 100 1135 104
rect 1139 100 1140 104
rect 1134 99 1140 100
rect 2118 104 2124 105
rect 2118 100 2119 104
rect 2123 100 2124 104
rect 2118 99 2124 100
rect 110 95 116 96
rect 110 91 111 95
rect 115 91 116 95
rect 1094 95 1100 96
rect 110 90 116 91
rect 134 92 140 93
rect 112 87 114 90
rect 134 88 135 92
rect 139 88 140 92
rect 134 87 140 88
rect 174 92 180 93
rect 174 88 175 92
rect 179 88 180 92
rect 174 87 180 88
rect 214 92 220 93
rect 214 88 215 92
rect 219 88 220 92
rect 214 87 220 88
rect 254 92 260 93
rect 254 88 255 92
rect 259 88 260 92
rect 254 87 260 88
rect 294 92 300 93
rect 294 88 295 92
rect 299 88 300 92
rect 294 87 300 88
rect 334 92 340 93
rect 334 88 335 92
rect 339 88 340 92
rect 334 87 340 88
rect 374 92 380 93
rect 374 88 375 92
rect 379 88 380 92
rect 374 87 380 88
rect 414 92 420 93
rect 414 88 415 92
rect 419 88 420 92
rect 414 87 420 88
rect 454 92 460 93
rect 454 88 455 92
rect 459 88 460 92
rect 454 87 460 88
rect 494 92 500 93
rect 494 88 495 92
rect 499 88 500 92
rect 494 87 500 88
rect 534 92 540 93
rect 534 88 535 92
rect 539 88 540 92
rect 534 87 540 88
rect 574 92 580 93
rect 574 88 575 92
rect 579 88 580 92
rect 574 87 580 88
rect 614 92 620 93
rect 614 88 615 92
rect 619 88 620 92
rect 614 87 620 88
rect 654 92 660 93
rect 654 88 655 92
rect 659 88 660 92
rect 654 87 660 88
rect 694 92 700 93
rect 694 88 695 92
rect 699 88 700 92
rect 694 87 700 88
rect 734 92 740 93
rect 734 88 735 92
rect 739 88 740 92
rect 734 87 740 88
rect 774 92 780 93
rect 774 88 775 92
rect 779 88 780 92
rect 774 87 780 88
rect 814 92 820 93
rect 814 88 815 92
rect 819 88 820 92
rect 814 87 820 88
rect 870 92 876 93
rect 870 88 871 92
rect 875 88 876 92
rect 870 87 876 88
rect 934 92 940 93
rect 934 88 935 92
rect 939 88 940 92
rect 934 87 940 88
rect 998 92 1004 93
rect 998 88 999 92
rect 1003 88 1004 92
rect 998 87 1004 88
rect 1046 92 1052 93
rect 1046 88 1047 92
rect 1051 88 1052 92
rect 1094 91 1095 95
rect 1099 91 1100 95
rect 1094 90 1100 91
rect 1046 87 1052 88
rect 1096 87 1098 90
rect 1134 87 1140 88
rect 111 86 115 87
rect 111 81 115 82
rect 135 86 139 87
rect 135 81 139 82
rect 175 86 179 87
rect 175 81 179 82
rect 215 86 219 87
rect 215 81 219 82
rect 255 86 259 87
rect 255 81 259 82
rect 295 86 299 87
rect 295 81 299 82
rect 335 86 339 87
rect 335 81 339 82
rect 375 86 379 87
rect 375 81 379 82
rect 415 86 419 87
rect 415 81 419 82
rect 455 86 459 87
rect 455 81 459 82
rect 495 86 499 87
rect 495 81 499 82
rect 535 86 539 87
rect 535 81 539 82
rect 575 86 579 87
rect 575 81 579 82
rect 615 86 619 87
rect 615 81 619 82
rect 655 86 659 87
rect 655 81 659 82
rect 695 86 699 87
rect 695 81 699 82
rect 735 86 739 87
rect 735 81 739 82
rect 775 86 779 87
rect 775 81 779 82
rect 815 86 819 87
rect 815 81 819 82
rect 871 86 875 87
rect 871 81 875 82
rect 935 86 939 87
rect 935 81 939 82
rect 999 86 1003 87
rect 999 81 1003 82
rect 1047 86 1051 87
rect 1047 81 1051 82
rect 1095 86 1099 87
rect 1134 83 1135 87
rect 1139 83 1140 87
rect 2118 87 2124 88
rect 1134 82 1140 83
rect 1158 84 1164 85
rect 1095 81 1099 82
rect 1136 79 1138 82
rect 1158 80 1159 84
rect 1163 80 1164 84
rect 1158 79 1164 80
rect 1198 84 1204 85
rect 1198 80 1199 84
rect 1203 80 1204 84
rect 1198 79 1204 80
rect 1238 84 1244 85
rect 1238 80 1239 84
rect 1243 80 1244 84
rect 1238 79 1244 80
rect 1278 84 1284 85
rect 1278 80 1279 84
rect 1283 80 1284 84
rect 1278 79 1284 80
rect 1318 84 1324 85
rect 1318 80 1319 84
rect 1323 80 1324 84
rect 1318 79 1324 80
rect 1366 84 1372 85
rect 1366 80 1367 84
rect 1371 80 1372 84
rect 1366 79 1372 80
rect 1430 84 1436 85
rect 1430 80 1431 84
rect 1435 80 1436 84
rect 1430 79 1436 80
rect 1494 84 1500 85
rect 1494 80 1495 84
rect 1499 80 1500 84
rect 1494 79 1500 80
rect 1558 84 1564 85
rect 1558 80 1559 84
rect 1563 80 1564 84
rect 1558 79 1564 80
rect 1614 84 1620 85
rect 1614 80 1615 84
rect 1619 80 1620 84
rect 1614 79 1620 80
rect 1670 84 1676 85
rect 1670 80 1671 84
rect 1675 80 1676 84
rect 1670 79 1676 80
rect 1718 84 1724 85
rect 1718 80 1719 84
rect 1723 80 1724 84
rect 1718 79 1724 80
rect 1766 84 1772 85
rect 1766 80 1767 84
rect 1771 80 1772 84
rect 1766 79 1772 80
rect 1806 84 1812 85
rect 1806 80 1807 84
rect 1811 80 1812 84
rect 1806 79 1812 80
rect 1854 84 1860 85
rect 1854 80 1855 84
rect 1859 80 1860 84
rect 1854 79 1860 80
rect 1902 84 1908 85
rect 1902 80 1903 84
rect 1907 80 1908 84
rect 1902 79 1908 80
rect 1950 84 1956 85
rect 1950 80 1951 84
rect 1955 80 1956 84
rect 1950 79 1956 80
rect 1990 84 1996 85
rect 1990 80 1991 84
rect 1995 80 1996 84
rect 1990 79 1996 80
rect 2030 84 2036 85
rect 2030 80 2031 84
rect 2035 80 2036 84
rect 2030 79 2036 80
rect 2070 84 2076 85
rect 2070 80 2071 84
rect 2075 80 2076 84
rect 2118 83 2119 87
rect 2123 83 2124 87
rect 2118 82 2124 83
rect 2070 79 2076 80
rect 2120 79 2122 82
rect 1135 78 1139 79
rect 1135 73 1139 74
rect 1159 78 1163 79
rect 1159 73 1163 74
rect 1199 78 1203 79
rect 1199 73 1203 74
rect 1239 78 1243 79
rect 1239 73 1243 74
rect 1279 78 1283 79
rect 1279 73 1283 74
rect 1319 78 1323 79
rect 1319 73 1323 74
rect 1367 78 1371 79
rect 1367 73 1371 74
rect 1431 78 1435 79
rect 1431 73 1435 74
rect 1495 78 1499 79
rect 1495 73 1499 74
rect 1559 78 1563 79
rect 1559 73 1563 74
rect 1615 78 1619 79
rect 1615 73 1619 74
rect 1671 78 1675 79
rect 1671 73 1675 74
rect 1719 78 1723 79
rect 1719 73 1723 74
rect 1767 78 1771 79
rect 1767 73 1771 74
rect 1807 78 1811 79
rect 1807 73 1811 74
rect 1855 78 1859 79
rect 1855 73 1859 74
rect 1903 78 1907 79
rect 1903 73 1907 74
rect 1951 78 1955 79
rect 1951 73 1955 74
rect 1991 78 1995 79
rect 1991 73 1995 74
rect 2031 78 2035 79
rect 2031 73 2035 74
rect 2071 78 2075 79
rect 2071 73 2075 74
rect 2119 78 2123 79
rect 2119 73 2123 74
<< m4c >>
rect 1135 2210 1139 2214
rect 1343 2210 1347 2214
rect 1383 2210 1387 2214
rect 1423 2210 1427 2214
rect 1463 2210 1467 2214
rect 1503 2210 1507 2214
rect 1543 2210 1547 2214
rect 1583 2210 1587 2214
rect 1623 2210 1627 2214
rect 1663 2210 1667 2214
rect 1703 2210 1707 2214
rect 1743 2210 1747 2214
rect 1783 2210 1787 2214
rect 1823 2210 1827 2214
rect 2119 2210 2123 2214
rect 1135 2158 1139 2162
rect 1287 2158 1291 2162
rect 1327 2158 1331 2162
rect 1343 2158 1347 2162
rect 1367 2158 1371 2162
rect 1383 2158 1387 2162
rect 1415 2158 1419 2162
rect 1423 2158 1427 2162
rect 1463 2158 1467 2162
rect 1503 2158 1507 2162
rect 1519 2158 1523 2162
rect 1543 2158 1547 2162
rect 1575 2158 1579 2162
rect 1583 2158 1587 2162
rect 1623 2158 1627 2162
rect 1663 2158 1667 2162
rect 1671 2158 1675 2162
rect 1703 2158 1707 2162
rect 1719 2158 1723 2162
rect 1743 2158 1747 2162
rect 1775 2158 1779 2162
rect 1783 2158 1787 2162
rect 1823 2158 1827 2162
rect 1831 2158 1835 2162
rect 1887 2158 1891 2162
rect 2119 2158 2123 2162
rect 1135 2102 1139 2106
rect 1223 2102 1227 2106
rect 1279 2102 1283 2106
rect 1287 2102 1291 2106
rect 1327 2102 1331 2106
rect 1343 2102 1347 2106
rect 1367 2102 1371 2106
rect 1415 2102 1419 2106
rect 1423 2102 1427 2106
rect 1463 2102 1467 2106
rect 1503 2102 1507 2106
rect 1519 2102 1523 2106
rect 1575 2102 1579 2106
rect 1583 2102 1587 2106
rect 1623 2102 1627 2106
rect 1663 2102 1667 2106
rect 1671 2102 1675 2106
rect 1719 2102 1723 2106
rect 1743 2102 1747 2106
rect 1775 2102 1779 2106
rect 1831 2102 1835 2106
rect 1887 2102 1891 2106
rect 1919 2102 1923 2106
rect 2007 2102 2011 2106
rect 2071 2102 2075 2106
rect 2119 2102 2123 2106
rect 1135 2050 1139 2054
rect 1183 2050 1187 2054
rect 1223 2050 1227 2054
rect 1239 2050 1243 2054
rect 1279 2050 1283 2054
rect 1311 2050 1315 2054
rect 1343 2050 1347 2054
rect 1399 2050 1403 2054
rect 1423 2050 1427 2054
rect 1487 2050 1491 2054
rect 1503 2050 1507 2054
rect 1583 2050 1587 2054
rect 1663 2050 1667 2054
rect 1671 2050 1675 2054
rect 1743 2050 1747 2054
rect 1759 2050 1763 2054
rect 1831 2050 1835 2054
rect 1839 2050 1843 2054
rect 1919 2050 1923 2054
rect 2007 2050 2011 2054
rect 2071 2050 2075 2054
rect 2119 2050 2123 2054
rect 111 2030 115 2034
rect 191 2030 195 2034
rect 231 2030 235 2034
rect 287 2030 291 2034
rect 351 2030 355 2034
rect 423 2030 427 2034
rect 495 2030 499 2034
rect 575 2030 579 2034
rect 647 2030 651 2034
rect 719 2030 723 2034
rect 783 2030 787 2034
rect 839 2030 843 2034
rect 895 2030 899 2034
rect 951 2030 955 2034
rect 1007 2030 1011 2034
rect 1047 2030 1051 2034
rect 1095 2030 1099 2034
rect 1135 1998 1139 2002
rect 1183 1998 1187 2002
rect 1239 1998 1243 2002
rect 1303 1998 1307 2002
rect 1311 1998 1315 2002
rect 1383 1998 1387 2002
rect 1399 1998 1403 2002
rect 1463 1998 1467 2002
rect 1487 1998 1491 2002
rect 1543 1998 1547 2002
rect 1583 1998 1587 2002
rect 1615 1998 1619 2002
rect 1671 1998 1675 2002
rect 1687 1998 1691 2002
rect 1751 1998 1755 2002
rect 1759 1998 1763 2002
rect 1815 1998 1819 2002
rect 1839 1998 1843 2002
rect 1879 1998 1883 2002
rect 1919 1998 1923 2002
rect 1951 1998 1955 2002
rect 2007 1998 2011 2002
rect 2023 1998 2027 2002
rect 2071 1998 2075 2002
rect 2119 1998 2123 2002
rect 111 1978 115 1982
rect 191 1978 195 1982
rect 231 1978 235 1982
rect 247 1978 251 1982
rect 287 1978 291 1982
rect 311 1978 315 1982
rect 351 1978 355 1982
rect 375 1978 379 1982
rect 423 1978 427 1982
rect 447 1978 451 1982
rect 495 1978 499 1982
rect 519 1978 523 1982
rect 575 1978 579 1982
rect 591 1978 595 1982
rect 647 1978 651 1982
rect 655 1978 659 1982
rect 719 1978 723 1982
rect 775 1978 779 1982
rect 783 1978 787 1982
rect 823 1978 827 1982
rect 839 1978 843 1982
rect 871 1978 875 1982
rect 895 1978 899 1982
rect 919 1978 923 1982
rect 951 1978 955 1982
rect 967 1978 971 1982
rect 1007 1978 1011 1982
rect 1047 1978 1051 1982
rect 1095 1978 1099 1982
rect 1135 1942 1139 1946
rect 1159 1942 1163 1946
rect 1223 1942 1227 1946
rect 1303 1942 1307 1946
rect 1383 1942 1387 1946
rect 1463 1942 1467 1946
rect 1535 1942 1539 1946
rect 1543 1942 1547 1946
rect 1615 1942 1619 1946
rect 1687 1942 1691 1946
rect 1695 1942 1699 1946
rect 1751 1942 1755 1946
rect 1783 1942 1787 1946
rect 1815 1942 1819 1946
rect 1879 1942 1883 1946
rect 1951 1942 1955 1946
rect 1983 1942 1987 1946
rect 2023 1942 2027 1946
rect 2071 1942 2075 1946
rect 2119 1942 2123 1946
rect 111 1926 115 1930
rect 135 1926 139 1930
rect 175 1926 179 1930
rect 191 1926 195 1930
rect 231 1926 235 1930
rect 247 1926 251 1930
rect 295 1926 299 1930
rect 311 1926 315 1930
rect 367 1926 371 1930
rect 375 1926 379 1930
rect 431 1926 435 1930
rect 447 1926 451 1930
rect 495 1926 499 1930
rect 519 1926 523 1930
rect 559 1926 563 1930
rect 591 1926 595 1930
rect 615 1926 619 1930
rect 655 1926 659 1930
rect 671 1926 675 1930
rect 719 1926 723 1930
rect 727 1926 731 1930
rect 775 1926 779 1930
rect 783 1926 787 1930
rect 823 1926 827 1930
rect 847 1926 851 1930
rect 871 1926 875 1930
rect 919 1926 923 1930
rect 967 1926 971 1930
rect 1007 1926 1011 1930
rect 1047 1926 1051 1930
rect 1095 1926 1099 1930
rect 1135 1886 1139 1890
rect 1159 1886 1163 1890
rect 1199 1886 1203 1890
rect 1223 1886 1227 1890
rect 1263 1886 1267 1890
rect 1303 1886 1307 1890
rect 1327 1886 1331 1890
rect 1383 1886 1387 1890
rect 1391 1886 1395 1890
rect 1447 1886 1451 1890
rect 1463 1886 1467 1890
rect 1503 1886 1507 1890
rect 1535 1886 1539 1890
rect 1559 1886 1563 1890
rect 1615 1886 1619 1890
rect 1631 1886 1635 1890
rect 1695 1886 1699 1890
rect 1711 1886 1715 1890
rect 1783 1886 1787 1890
rect 1799 1886 1803 1890
rect 1879 1886 1883 1890
rect 1895 1886 1899 1890
rect 1983 1886 1987 1890
rect 1991 1886 1995 1890
rect 2071 1886 2075 1890
rect 2119 1886 2123 1890
rect 111 1870 115 1874
rect 135 1870 139 1874
rect 175 1870 179 1874
rect 199 1870 203 1874
rect 231 1870 235 1874
rect 271 1870 275 1874
rect 295 1870 299 1874
rect 335 1870 339 1874
rect 367 1870 371 1874
rect 399 1870 403 1874
rect 431 1870 435 1874
rect 455 1870 459 1874
rect 495 1870 499 1874
rect 503 1870 507 1874
rect 551 1870 555 1874
rect 559 1870 563 1874
rect 599 1870 603 1874
rect 615 1870 619 1874
rect 647 1870 651 1874
rect 671 1870 675 1874
rect 695 1870 699 1874
rect 727 1870 731 1874
rect 751 1870 755 1874
rect 783 1870 787 1874
rect 847 1870 851 1874
rect 1095 1870 1099 1874
rect 1135 1834 1139 1838
rect 1159 1834 1163 1838
rect 1199 1834 1203 1838
rect 1231 1834 1235 1838
rect 1263 1834 1267 1838
rect 1303 1834 1307 1838
rect 1327 1834 1331 1838
rect 1383 1834 1387 1838
rect 1391 1834 1395 1838
rect 1447 1834 1451 1838
rect 1463 1834 1467 1838
rect 1503 1834 1507 1838
rect 1551 1834 1555 1838
rect 1559 1834 1563 1838
rect 1631 1834 1635 1838
rect 1647 1834 1651 1838
rect 1711 1834 1715 1838
rect 1751 1834 1755 1838
rect 1799 1834 1803 1838
rect 1855 1834 1859 1838
rect 1895 1834 1899 1838
rect 1967 1834 1971 1838
rect 1991 1834 1995 1838
rect 2071 1834 2075 1838
rect 2119 1834 2123 1838
rect 111 1810 115 1814
rect 135 1810 139 1814
rect 151 1810 155 1814
rect 199 1810 203 1814
rect 215 1810 219 1814
rect 271 1810 275 1814
rect 327 1810 331 1814
rect 335 1810 339 1814
rect 383 1810 387 1814
rect 399 1810 403 1814
rect 431 1810 435 1814
rect 455 1810 459 1814
rect 479 1810 483 1814
rect 503 1810 507 1814
rect 527 1810 531 1814
rect 551 1810 555 1814
rect 575 1810 579 1814
rect 599 1810 603 1814
rect 623 1810 627 1814
rect 647 1810 651 1814
rect 671 1810 675 1814
rect 695 1810 699 1814
rect 727 1810 731 1814
rect 751 1810 755 1814
rect 1095 1810 1099 1814
rect 1135 1782 1139 1786
rect 1159 1782 1163 1786
rect 1191 1782 1195 1786
rect 1231 1782 1235 1786
rect 1255 1782 1259 1786
rect 1303 1782 1307 1786
rect 1319 1782 1323 1786
rect 1383 1782 1387 1786
rect 1455 1782 1459 1786
rect 1463 1782 1467 1786
rect 1527 1782 1531 1786
rect 1551 1782 1555 1786
rect 1607 1782 1611 1786
rect 1647 1782 1651 1786
rect 1687 1782 1691 1786
rect 1751 1782 1755 1786
rect 1767 1782 1771 1786
rect 1847 1782 1851 1786
rect 1855 1782 1859 1786
rect 1927 1782 1931 1786
rect 1967 1782 1971 1786
rect 2007 1782 2011 1786
rect 2071 1782 2075 1786
rect 2119 1782 2123 1786
rect 111 1758 115 1762
rect 151 1758 155 1762
rect 215 1758 219 1762
rect 231 1758 235 1762
rect 271 1758 275 1762
rect 295 1758 299 1762
rect 327 1758 331 1762
rect 351 1758 355 1762
rect 383 1758 387 1762
rect 415 1758 419 1762
rect 431 1758 435 1762
rect 479 1758 483 1762
rect 527 1758 531 1762
rect 543 1758 547 1762
rect 575 1758 579 1762
rect 615 1758 619 1762
rect 623 1758 627 1762
rect 671 1758 675 1762
rect 687 1758 691 1762
rect 727 1758 731 1762
rect 759 1758 763 1762
rect 831 1758 835 1762
rect 911 1758 915 1762
rect 991 1758 995 1762
rect 1095 1758 1099 1762
rect 1135 1730 1139 1734
rect 1191 1730 1195 1734
rect 1247 1730 1251 1734
rect 1255 1730 1259 1734
rect 1295 1730 1299 1734
rect 1319 1730 1323 1734
rect 1343 1730 1347 1734
rect 1383 1730 1387 1734
rect 1399 1730 1403 1734
rect 1455 1730 1459 1734
rect 1463 1730 1467 1734
rect 1527 1730 1531 1734
rect 1599 1730 1603 1734
rect 1607 1730 1611 1734
rect 1671 1730 1675 1734
rect 1687 1730 1691 1734
rect 1743 1730 1747 1734
rect 1767 1730 1771 1734
rect 1807 1730 1811 1734
rect 1847 1730 1851 1734
rect 1879 1730 1883 1734
rect 1927 1730 1931 1734
rect 1951 1730 1955 1734
rect 2007 1730 2011 1734
rect 2023 1730 2027 1734
rect 2071 1730 2075 1734
rect 2119 1730 2123 1734
rect 111 1702 115 1706
rect 135 1702 139 1706
rect 199 1702 203 1706
rect 231 1702 235 1706
rect 279 1702 283 1706
rect 295 1702 299 1706
rect 351 1702 355 1706
rect 367 1702 371 1706
rect 415 1702 419 1706
rect 463 1702 467 1706
rect 479 1702 483 1706
rect 543 1702 547 1706
rect 551 1702 555 1706
rect 615 1702 619 1706
rect 639 1702 643 1706
rect 687 1702 691 1706
rect 719 1702 723 1706
rect 759 1702 763 1706
rect 791 1702 795 1706
rect 831 1702 835 1706
rect 855 1702 859 1706
rect 911 1702 915 1706
rect 919 1702 923 1706
rect 983 1702 987 1706
rect 991 1702 995 1706
rect 1047 1702 1051 1706
rect 1095 1702 1099 1706
rect 1135 1674 1139 1678
rect 1247 1674 1251 1678
rect 1263 1674 1267 1678
rect 1295 1674 1299 1678
rect 1303 1674 1307 1678
rect 1343 1674 1347 1678
rect 1391 1674 1395 1678
rect 1399 1674 1403 1678
rect 1447 1674 1451 1678
rect 1463 1674 1467 1678
rect 1503 1674 1507 1678
rect 1527 1674 1531 1678
rect 1567 1674 1571 1678
rect 1599 1674 1603 1678
rect 1631 1674 1635 1678
rect 1671 1674 1675 1678
rect 1695 1674 1699 1678
rect 1743 1674 1747 1678
rect 1759 1674 1763 1678
rect 1807 1674 1811 1678
rect 1831 1674 1835 1678
rect 1879 1674 1883 1678
rect 1911 1674 1915 1678
rect 1951 1674 1955 1678
rect 1999 1674 2003 1678
rect 2023 1674 2027 1678
rect 2071 1674 2075 1678
rect 2119 1674 2123 1678
rect 111 1646 115 1650
rect 135 1646 139 1650
rect 183 1646 187 1650
rect 199 1646 203 1650
rect 263 1646 267 1650
rect 279 1646 283 1650
rect 343 1646 347 1650
rect 367 1646 371 1650
rect 423 1646 427 1650
rect 463 1646 467 1650
rect 503 1646 507 1650
rect 551 1646 555 1650
rect 583 1646 587 1650
rect 639 1646 643 1650
rect 655 1646 659 1650
rect 719 1646 723 1650
rect 727 1646 731 1650
rect 791 1646 795 1650
rect 847 1646 851 1650
rect 855 1646 859 1650
rect 903 1646 907 1650
rect 919 1646 923 1650
rect 959 1646 963 1650
rect 983 1646 987 1650
rect 1007 1646 1011 1650
rect 1047 1646 1051 1650
rect 1095 1646 1099 1650
rect 1135 1610 1139 1614
rect 1159 1610 1163 1614
rect 1215 1610 1219 1614
rect 1263 1610 1267 1614
rect 1303 1610 1307 1614
rect 1343 1610 1347 1614
rect 1383 1610 1387 1614
rect 1391 1610 1395 1614
rect 1447 1610 1451 1614
rect 1463 1610 1467 1614
rect 1503 1610 1507 1614
rect 1543 1610 1547 1614
rect 1567 1610 1571 1614
rect 1623 1610 1627 1614
rect 1631 1610 1635 1614
rect 1695 1610 1699 1614
rect 1711 1610 1715 1614
rect 1759 1610 1763 1614
rect 1799 1610 1803 1614
rect 1831 1610 1835 1614
rect 1887 1610 1891 1614
rect 1911 1610 1915 1614
rect 1983 1610 1987 1614
rect 1999 1610 2003 1614
rect 2071 1610 2075 1614
rect 2119 1610 2123 1614
rect 111 1594 115 1598
rect 135 1594 139 1598
rect 175 1594 179 1598
rect 183 1594 187 1598
rect 231 1594 235 1598
rect 263 1594 267 1598
rect 303 1594 307 1598
rect 343 1594 347 1598
rect 375 1594 379 1598
rect 423 1594 427 1598
rect 455 1594 459 1598
rect 503 1594 507 1598
rect 527 1594 531 1598
rect 583 1594 587 1598
rect 599 1594 603 1598
rect 655 1594 659 1598
rect 671 1594 675 1598
rect 727 1594 731 1598
rect 743 1594 747 1598
rect 791 1594 795 1598
rect 815 1594 819 1598
rect 847 1594 851 1598
rect 887 1594 891 1598
rect 903 1594 907 1598
rect 959 1594 963 1598
rect 1007 1594 1011 1598
rect 1047 1594 1051 1598
rect 1095 1594 1099 1598
rect 1135 1558 1139 1562
rect 1159 1558 1163 1562
rect 1199 1558 1203 1562
rect 1215 1558 1219 1562
rect 1247 1558 1251 1562
rect 1303 1558 1307 1562
rect 1319 1558 1323 1562
rect 1383 1558 1387 1562
rect 1399 1558 1403 1562
rect 1463 1558 1467 1562
rect 1479 1558 1483 1562
rect 1543 1558 1547 1562
rect 1559 1558 1563 1562
rect 1623 1558 1627 1562
rect 1647 1558 1651 1562
rect 1711 1558 1715 1562
rect 1735 1558 1739 1562
rect 1799 1558 1803 1562
rect 1823 1558 1827 1562
rect 1887 1558 1891 1562
rect 1911 1558 1915 1562
rect 1983 1558 1987 1562
rect 1999 1558 2003 1562
rect 2071 1558 2075 1562
rect 2119 1558 2123 1562
rect 111 1542 115 1546
rect 135 1542 139 1546
rect 175 1542 179 1546
rect 231 1542 235 1546
rect 303 1542 307 1546
rect 311 1542 315 1546
rect 375 1542 379 1546
rect 391 1542 395 1546
rect 455 1542 459 1546
rect 479 1542 483 1546
rect 527 1542 531 1546
rect 567 1542 571 1546
rect 599 1542 603 1546
rect 655 1542 659 1546
rect 671 1542 675 1546
rect 743 1542 747 1546
rect 815 1542 819 1546
rect 823 1542 827 1546
rect 887 1542 891 1546
rect 911 1542 915 1546
rect 999 1542 1003 1546
rect 1095 1542 1099 1546
rect 1135 1506 1139 1510
rect 1159 1506 1163 1510
rect 1199 1506 1203 1510
rect 1239 1506 1243 1510
rect 1247 1506 1251 1510
rect 1303 1506 1307 1510
rect 1319 1506 1323 1510
rect 1375 1506 1379 1510
rect 1399 1506 1403 1510
rect 1455 1506 1459 1510
rect 1479 1506 1483 1510
rect 1543 1506 1547 1510
rect 1559 1506 1563 1510
rect 1623 1506 1627 1510
rect 1647 1506 1651 1510
rect 1703 1506 1707 1510
rect 1735 1506 1739 1510
rect 1775 1506 1779 1510
rect 1823 1506 1827 1510
rect 1847 1506 1851 1510
rect 1911 1506 1915 1510
rect 1919 1506 1923 1510
rect 1991 1506 1995 1510
rect 1999 1506 2003 1510
rect 2063 1506 2067 1510
rect 2071 1506 2075 1510
rect 2119 1506 2123 1510
rect 111 1490 115 1494
rect 135 1490 139 1494
rect 175 1490 179 1494
rect 199 1490 203 1494
rect 231 1490 235 1494
rect 279 1490 283 1494
rect 311 1490 315 1494
rect 359 1490 363 1494
rect 391 1490 395 1494
rect 439 1490 443 1494
rect 479 1490 483 1494
rect 519 1490 523 1494
rect 567 1490 571 1494
rect 599 1490 603 1494
rect 655 1490 659 1494
rect 679 1490 683 1494
rect 743 1490 747 1494
rect 767 1490 771 1494
rect 823 1490 827 1494
rect 855 1490 859 1494
rect 911 1490 915 1494
rect 943 1490 947 1494
rect 999 1490 1003 1494
rect 1031 1490 1035 1494
rect 1095 1490 1099 1494
rect 1135 1450 1139 1454
rect 1159 1450 1163 1454
rect 1199 1450 1203 1454
rect 1239 1450 1243 1454
rect 1279 1450 1283 1454
rect 1303 1450 1307 1454
rect 1327 1450 1331 1454
rect 1375 1450 1379 1454
rect 1383 1450 1387 1454
rect 1439 1450 1443 1454
rect 1455 1450 1459 1454
rect 1495 1450 1499 1454
rect 1543 1450 1547 1454
rect 1551 1450 1555 1454
rect 1607 1450 1611 1454
rect 1623 1450 1627 1454
rect 1671 1450 1675 1454
rect 1703 1450 1707 1454
rect 1735 1450 1739 1454
rect 1775 1450 1779 1454
rect 1807 1450 1811 1454
rect 1847 1450 1851 1454
rect 1887 1450 1891 1454
rect 1919 1450 1923 1454
rect 1975 1450 1979 1454
rect 1991 1450 1995 1454
rect 2063 1450 2067 1454
rect 2119 1450 2123 1454
rect 111 1438 115 1442
rect 135 1438 139 1442
rect 191 1438 195 1442
rect 199 1438 203 1442
rect 263 1438 267 1442
rect 279 1438 283 1442
rect 335 1438 339 1442
rect 359 1438 363 1442
rect 407 1438 411 1442
rect 439 1438 443 1442
rect 479 1438 483 1442
rect 519 1438 523 1442
rect 551 1438 555 1442
rect 599 1438 603 1442
rect 631 1438 635 1442
rect 679 1438 683 1442
rect 711 1438 715 1442
rect 767 1438 771 1442
rect 799 1438 803 1442
rect 855 1438 859 1442
rect 887 1438 891 1442
rect 943 1438 947 1442
rect 975 1438 979 1442
rect 1031 1438 1035 1442
rect 1047 1438 1051 1442
rect 1095 1438 1099 1442
rect 1135 1394 1139 1398
rect 1279 1394 1283 1398
rect 1327 1394 1331 1398
rect 1335 1394 1339 1398
rect 1375 1394 1379 1398
rect 1383 1394 1387 1398
rect 1415 1394 1419 1398
rect 1439 1394 1443 1398
rect 1455 1394 1459 1398
rect 1495 1394 1499 1398
rect 1535 1394 1539 1398
rect 1551 1394 1555 1398
rect 1583 1394 1587 1398
rect 1607 1394 1611 1398
rect 1647 1394 1651 1398
rect 1671 1394 1675 1398
rect 1719 1394 1723 1398
rect 1735 1394 1739 1398
rect 1807 1394 1811 1398
rect 1887 1394 1891 1398
rect 1895 1394 1899 1398
rect 1975 1394 1979 1398
rect 1991 1394 1995 1398
rect 2063 1394 2067 1398
rect 2071 1394 2075 1398
rect 2119 1394 2123 1398
rect 111 1386 115 1390
rect 135 1386 139 1390
rect 175 1386 179 1390
rect 191 1386 195 1390
rect 239 1386 243 1390
rect 263 1386 267 1390
rect 303 1386 307 1390
rect 335 1386 339 1390
rect 367 1386 371 1390
rect 407 1386 411 1390
rect 439 1386 443 1390
rect 479 1386 483 1390
rect 503 1386 507 1390
rect 551 1386 555 1390
rect 575 1386 579 1390
rect 631 1386 635 1390
rect 647 1386 651 1390
rect 711 1386 715 1390
rect 783 1386 787 1390
rect 799 1386 803 1390
rect 855 1386 859 1390
rect 887 1386 891 1390
rect 927 1386 931 1390
rect 975 1386 979 1390
rect 999 1386 1003 1390
rect 1047 1386 1051 1390
rect 1095 1386 1099 1390
rect 1135 1342 1139 1346
rect 1159 1342 1163 1346
rect 1223 1342 1227 1346
rect 1311 1342 1315 1346
rect 1335 1342 1339 1346
rect 1375 1342 1379 1346
rect 1407 1342 1411 1346
rect 1415 1342 1419 1346
rect 1455 1342 1459 1346
rect 1495 1342 1499 1346
rect 1503 1342 1507 1346
rect 1535 1342 1539 1346
rect 1583 1342 1587 1346
rect 1599 1342 1603 1346
rect 1647 1342 1651 1346
rect 1679 1342 1683 1346
rect 1719 1342 1723 1346
rect 1759 1342 1763 1346
rect 1807 1342 1811 1346
rect 1831 1342 1835 1346
rect 1895 1342 1899 1346
rect 1959 1342 1963 1346
rect 1991 1342 1995 1346
rect 2023 1342 2027 1346
rect 2071 1342 2075 1346
rect 2119 1342 2123 1346
rect 111 1326 115 1330
rect 135 1326 139 1330
rect 175 1326 179 1330
rect 215 1326 219 1330
rect 239 1326 243 1330
rect 255 1326 259 1330
rect 303 1326 307 1330
rect 319 1326 323 1330
rect 367 1326 371 1330
rect 391 1326 395 1330
rect 439 1326 443 1330
rect 463 1326 467 1330
rect 503 1326 507 1330
rect 543 1326 547 1330
rect 575 1326 579 1330
rect 623 1326 627 1330
rect 647 1326 651 1330
rect 703 1326 707 1330
rect 711 1326 715 1330
rect 783 1326 787 1330
rect 855 1326 859 1330
rect 863 1326 867 1330
rect 927 1326 931 1330
rect 943 1326 947 1330
rect 999 1326 1003 1330
rect 1023 1326 1027 1330
rect 1047 1326 1051 1330
rect 1095 1326 1099 1330
rect 1135 1290 1139 1294
rect 1159 1290 1163 1294
rect 1175 1290 1179 1294
rect 1223 1290 1227 1294
rect 1231 1290 1235 1294
rect 1303 1290 1307 1294
rect 1311 1290 1315 1294
rect 1391 1290 1395 1294
rect 1407 1290 1411 1294
rect 1479 1290 1483 1294
rect 1503 1290 1507 1294
rect 1567 1290 1571 1294
rect 1599 1290 1603 1294
rect 1655 1290 1659 1294
rect 1679 1290 1683 1294
rect 1743 1290 1747 1294
rect 1759 1290 1763 1294
rect 1831 1290 1835 1294
rect 1895 1290 1899 1294
rect 1919 1290 1923 1294
rect 1959 1290 1963 1294
rect 2007 1290 2011 1294
rect 2023 1290 2027 1294
rect 2071 1290 2075 1294
rect 2119 1290 2123 1294
rect 111 1270 115 1274
rect 135 1270 139 1274
rect 175 1270 179 1274
rect 215 1270 219 1274
rect 255 1270 259 1274
rect 319 1270 323 1274
rect 391 1270 395 1274
rect 399 1270 403 1274
rect 463 1270 467 1274
rect 487 1270 491 1274
rect 543 1270 547 1274
rect 583 1270 587 1274
rect 623 1270 627 1274
rect 687 1270 691 1274
rect 703 1270 707 1274
rect 783 1270 787 1274
rect 799 1270 803 1274
rect 863 1270 867 1274
rect 919 1270 923 1274
rect 943 1270 947 1274
rect 1023 1270 1027 1274
rect 1047 1270 1051 1274
rect 1095 1270 1099 1274
rect 1135 1234 1139 1238
rect 1175 1234 1179 1238
rect 1231 1234 1235 1238
rect 1287 1234 1291 1238
rect 1303 1234 1307 1238
rect 1327 1234 1331 1238
rect 1375 1234 1379 1238
rect 1391 1234 1395 1238
rect 1431 1234 1435 1238
rect 1479 1234 1483 1238
rect 1495 1234 1499 1238
rect 1559 1234 1563 1238
rect 1567 1234 1571 1238
rect 1623 1234 1627 1238
rect 1655 1234 1659 1238
rect 1679 1234 1683 1238
rect 1735 1234 1739 1238
rect 1743 1234 1747 1238
rect 1791 1234 1795 1238
rect 1831 1234 1835 1238
rect 1847 1234 1851 1238
rect 1903 1234 1907 1238
rect 1919 1234 1923 1238
rect 1967 1234 1971 1238
rect 2007 1234 2011 1238
rect 2031 1234 2035 1238
rect 2071 1234 2075 1238
rect 2119 1234 2123 1238
rect 111 1214 115 1218
rect 135 1214 139 1218
rect 175 1214 179 1218
rect 215 1214 219 1218
rect 255 1214 259 1218
rect 271 1214 275 1218
rect 311 1214 315 1218
rect 319 1214 323 1218
rect 351 1214 355 1218
rect 399 1214 403 1218
rect 447 1214 451 1218
rect 487 1214 491 1218
rect 495 1214 499 1218
rect 551 1214 555 1218
rect 583 1214 587 1218
rect 607 1214 611 1218
rect 671 1214 675 1218
rect 687 1214 691 1218
rect 743 1214 747 1218
rect 799 1214 803 1218
rect 815 1214 819 1218
rect 895 1214 899 1218
rect 919 1214 923 1218
rect 983 1214 987 1218
rect 1047 1214 1051 1218
rect 1095 1214 1099 1218
rect 1135 1182 1139 1186
rect 1159 1182 1163 1186
rect 1207 1182 1211 1186
rect 1279 1182 1283 1186
rect 1287 1182 1291 1186
rect 1327 1182 1331 1186
rect 1351 1182 1355 1186
rect 1375 1182 1379 1186
rect 1423 1182 1427 1186
rect 1431 1182 1435 1186
rect 1487 1182 1491 1186
rect 1495 1182 1499 1186
rect 1559 1182 1563 1186
rect 1623 1182 1627 1186
rect 1631 1182 1635 1186
rect 1679 1182 1683 1186
rect 1711 1182 1715 1186
rect 1735 1182 1739 1186
rect 1791 1182 1795 1186
rect 1799 1182 1803 1186
rect 1847 1182 1851 1186
rect 1887 1182 1891 1186
rect 1903 1182 1907 1186
rect 1967 1182 1971 1186
rect 1983 1182 1987 1186
rect 2031 1182 2035 1186
rect 2071 1182 2075 1186
rect 2119 1182 2123 1186
rect 111 1158 115 1162
rect 271 1158 275 1162
rect 311 1158 315 1162
rect 351 1158 355 1162
rect 399 1158 403 1162
rect 439 1158 443 1162
rect 447 1158 451 1162
rect 479 1158 483 1162
rect 495 1158 499 1162
rect 527 1158 531 1162
rect 551 1158 555 1162
rect 575 1158 579 1162
rect 607 1158 611 1162
rect 623 1158 627 1162
rect 671 1158 675 1162
rect 719 1158 723 1162
rect 743 1158 747 1162
rect 775 1158 779 1162
rect 815 1158 819 1162
rect 831 1158 835 1162
rect 887 1158 891 1162
rect 895 1158 899 1162
rect 943 1158 947 1162
rect 983 1158 987 1162
rect 1007 1158 1011 1162
rect 1047 1158 1051 1162
rect 1095 1158 1099 1162
rect 1135 1126 1139 1130
rect 1159 1126 1163 1130
rect 1191 1126 1195 1130
rect 1207 1126 1211 1130
rect 1271 1126 1275 1130
rect 1279 1126 1283 1130
rect 1343 1126 1347 1130
rect 1351 1126 1355 1130
rect 1415 1126 1419 1130
rect 1423 1126 1427 1130
rect 1487 1126 1491 1130
rect 1559 1126 1563 1130
rect 1567 1126 1571 1130
rect 1631 1126 1635 1130
rect 1655 1126 1659 1130
rect 1711 1126 1715 1130
rect 1751 1126 1755 1130
rect 1799 1126 1803 1130
rect 1855 1126 1859 1130
rect 1887 1126 1891 1130
rect 1959 1126 1963 1130
rect 1983 1126 1987 1130
rect 2071 1126 2075 1130
rect 2119 1126 2123 1130
rect 111 1106 115 1110
rect 159 1106 163 1110
rect 199 1106 203 1110
rect 255 1106 259 1110
rect 319 1106 323 1110
rect 399 1106 403 1110
rect 439 1106 443 1110
rect 479 1106 483 1110
rect 527 1106 531 1110
rect 559 1106 563 1110
rect 575 1106 579 1110
rect 623 1106 627 1110
rect 639 1106 643 1110
rect 671 1106 675 1110
rect 711 1106 715 1110
rect 719 1106 723 1110
rect 775 1106 779 1110
rect 783 1106 787 1110
rect 831 1106 835 1110
rect 855 1106 859 1110
rect 887 1106 891 1110
rect 927 1106 931 1110
rect 943 1106 947 1110
rect 999 1106 1003 1110
rect 1007 1106 1011 1110
rect 1047 1106 1051 1110
rect 1095 1106 1099 1110
rect 1135 1074 1139 1078
rect 1159 1074 1163 1078
rect 1191 1074 1195 1078
rect 1199 1074 1203 1078
rect 1247 1074 1251 1078
rect 1271 1074 1275 1078
rect 1303 1074 1307 1078
rect 1343 1074 1347 1078
rect 1351 1074 1355 1078
rect 1399 1074 1403 1078
rect 1415 1074 1419 1078
rect 1455 1074 1459 1078
rect 1487 1074 1491 1078
rect 1511 1074 1515 1078
rect 1567 1074 1571 1078
rect 1583 1074 1587 1078
rect 1655 1074 1659 1078
rect 1663 1074 1667 1078
rect 1751 1074 1755 1078
rect 1759 1074 1763 1078
rect 1855 1074 1859 1078
rect 1863 1074 1867 1078
rect 1959 1074 1963 1078
rect 1967 1074 1971 1078
rect 2071 1074 2075 1078
rect 2119 1074 2123 1078
rect 111 1050 115 1054
rect 135 1050 139 1054
rect 159 1050 163 1054
rect 175 1050 179 1054
rect 199 1050 203 1054
rect 215 1050 219 1054
rect 255 1050 259 1054
rect 319 1050 323 1054
rect 383 1050 387 1054
rect 399 1050 403 1054
rect 447 1050 451 1054
rect 479 1050 483 1054
rect 511 1050 515 1054
rect 559 1050 563 1054
rect 575 1050 579 1054
rect 631 1050 635 1054
rect 639 1050 643 1054
rect 687 1050 691 1054
rect 711 1050 715 1054
rect 743 1050 747 1054
rect 783 1050 787 1054
rect 799 1050 803 1054
rect 855 1050 859 1054
rect 863 1050 867 1054
rect 927 1050 931 1054
rect 999 1050 1003 1054
rect 1047 1050 1051 1054
rect 1095 1050 1099 1054
rect 1135 1018 1139 1022
rect 1159 1018 1163 1022
rect 1199 1018 1203 1022
rect 1239 1018 1243 1022
rect 1247 1018 1251 1022
rect 1295 1018 1299 1022
rect 1303 1018 1307 1022
rect 1351 1018 1355 1022
rect 1399 1018 1403 1022
rect 1407 1018 1411 1022
rect 1455 1018 1459 1022
rect 1463 1018 1467 1022
rect 1511 1018 1515 1022
rect 1519 1018 1523 1022
rect 1575 1018 1579 1022
rect 1583 1018 1587 1022
rect 1639 1018 1643 1022
rect 1663 1018 1667 1022
rect 1711 1018 1715 1022
rect 1759 1018 1763 1022
rect 1791 1018 1795 1022
rect 1863 1018 1867 1022
rect 1879 1018 1883 1022
rect 1967 1018 1971 1022
rect 2063 1018 2067 1022
rect 2071 1018 2075 1022
rect 2119 1018 2123 1022
rect 111 994 115 998
rect 135 994 139 998
rect 175 994 179 998
rect 215 994 219 998
rect 223 994 227 998
rect 255 994 259 998
rect 279 994 283 998
rect 319 994 323 998
rect 343 994 347 998
rect 383 994 387 998
rect 407 994 411 998
rect 447 994 451 998
rect 471 994 475 998
rect 511 994 515 998
rect 527 994 531 998
rect 575 994 579 998
rect 583 994 587 998
rect 631 994 635 998
rect 687 994 691 998
rect 743 994 747 998
rect 799 994 803 998
rect 863 994 867 998
rect 1095 994 1099 998
rect 1135 958 1139 962
rect 1159 958 1163 962
rect 1199 958 1203 962
rect 1207 958 1211 962
rect 1239 958 1243 962
rect 1287 958 1291 962
rect 1295 958 1299 962
rect 1351 958 1355 962
rect 1375 958 1379 962
rect 1407 958 1411 962
rect 1455 958 1459 962
rect 1463 958 1467 962
rect 1519 958 1523 962
rect 1535 958 1539 962
rect 1575 958 1579 962
rect 1615 958 1619 962
rect 1639 958 1643 962
rect 1687 958 1691 962
rect 1711 958 1715 962
rect 1751 958 1755 962
rect 1791 958 1795 962
rect 1815 958 1819 962
rect 1879 958 1883 962
rect 1951 958 1955 962
rect 1967 958 1971 962
rect 2023 958 2027 962
rect 2063 958 2067 962
rect 2071 958 2075 962
rect 2119 958 2123 962
rect 111 938 115 942
rect 135 938 139 942
rect 175 938 179 942
rect 223 938 227 942
rect 263 938 267 942
rect 279 938 283 942
rect 303 938 307 942
rect 343 938 347 942
rect 351 938 355 942
rect 399 938 403 942
rect 407 938 411 942
rect 455 938 459 942
rect 471 938 475 942
rect 511 938 515 942
rect 527 938 531 942
rect 567 938 571 942
rect 583 938 587 942
rect 623 938 627 942
rect 631 938 635 942
rect 687 938 691 942
rect 743 938 747 942
rect 751 938 755 942
rect 799 938 803 942
rect 815 938 819 942
rect 879 938 883 942
rect 943 938 947 942
rect 1007 938 1011 942
rect 1047 938 1051 942
rect 1095 938 1099 942
rect 1135 906 1139 910
rect 1159 906 1163 910
rect 1207 906 1211 910
rect 1239 906 1243 910
rect 1287 906 1291 910
rect 1319 906 1323 910
rect 1375 906 1379 910
rect 1407 906 1411 910
rect 1455 906 1459 910
rect 1495 906 1499 910
rect 1535 906 1539 910
rect 1583 906 1587 910
rect 1615 906 1619 910
rect 1663 906 1667 910
rect 1687 906 1691 910
rect 1743 906 1747 910
rect 1751 906 1755 910
rect 1815 906 1819 910
rect 1879 906 1883 910
rect 1887 906 1891 910
rect 1951 906 1955 910
rect 2023 906 2027 910
rect 2071 906 2075 910
rect 2119 906 2123 910
rect 111 882 115 886
rect 263 882 267 886
rect 303 882 307 886
rect 351 882 355 886
rect 399 882 403 886
rect 415 882 419 886
rect 455 882 459 886
rect 479 882 483 886
rect 511 882 515 886
rect 551 882 555 886
rect 567 882 571 886
rect 623 882 627 886
rect 687 882 691 886
rect 695 882 699 886
rect 751 882 755 886
rect 767 882 771 886
rect 815 882 819 886
rect 831 882 835 886
rect 879 882 883 886
rect 887 882 891 886
rect 943 882 947 886
rect 1007 882 1011 886
rect 1047 882 1051 886
rect 1095 882 1099 886
rect 1135 854 1139 858
rect 1159 854 1163 858
rect 1239 854 1243 858
rect 1247 854 1251 858
rect 1319 854 1323 858
rect 1359 854 1363 858
rect 1407 854 1411 858
rect 1455 854 1459 858
rect 1495 854 1499 858
rect 1543 854 1547 858
rect 1583 854 1587 858
rect 1631 854 1635 858
rect 1663 854 1667 858
rect 1711 854 1715 858
rect 1743 854 1747 858
rect 1783 854 1787 858
rect 1815 854 1819 858
rect 1855 854 1859 858
rect 1887 854 1891 858
rect 1935 854 1939 858
rect 1951 854 1955 858
rect 2015 854 2019 858
rect 2023 854 2027 858
rect 2071 854 2075 858
rect 2119 854 2123 858
rect 111 830 115 834
rect 279 830 283 834
rect 303 830 307 834
rect 343 830 347 834
rect 351 830 355 834
rect 415 830 419 834
rect 479 830 483 834
rect 487 830 491 834
rect 551 830 555 834
rect 567 830 571 834
rect 623 830 627 834
rect 647 830 651 834
rect 695 830 699 834
rect 727 830 731 834
rect 767 830 771 834
rect 799 830 803 834
rect 831 830 835 834
rect 863 830 867 834
rect 887 830 891 834
rect 927 830 931 834
rect 943 830 947 834
rect 999 830 1003 834
rect 1007 830 1011 834
rect 1047 830 1051 834
rect 1095 830 1099 834
rect 1135 802 1139 806
rect 1159 802 1163 806
rect 1247 802 1251 806
rect 1279 802 1283 806
rect 1359 802 1363 806
rect 1407 802 1411 806
rect 1455 802 1459 806
rect 1519 802 1523 806
rect 1543 802 1547 806
rect 1623 802 1627 806
rect 1631 802 1635 806
rect 1711 802 1715 806
rect 1719 802 1723 806
rect 1783 802 1787 806
rect 1815 802 1819 806
rect 1855 802 1859 806
rect 1903 802 1907 806
rect 1935 802 1939 806
rect 1999 802 2003 806
rect 2015 802 2019 806
rect 2071 802 2075 806
rect 2119 802 2123 806
rect 111 778 115 782
rect 215 778 219 782
rect 279 778 283 782
rect 343 778 347 782
rect 351 778 355 782
rect 415 778 419 782
rect 423 778 427 782
rect 487 778 491 782
rect 495 778 499 782
rect 567 778 571 782
rect 639 778 643 782
rect 647 778 651 782
rect 703 778 707 782
rect 727 778 731 782
rect 759 778 763 782
rect 799 778 803 782
rect 815 778 819 782
rect 863 778 867 782
rect 911 778 915 782
rect 927 778 931 782
rect 959 778 963 782
rect 999 778 1003 782
rect 1007 778 1011 782
rect 1047 778 1051 782
rect 1095 778 1099 782
rect 1135 746 1139 750
rect 1159 746 1163 750
rect 1279 746 1283 750
rect 1335 746 1339 750
rect 1375 746 1379 750
rect 1407 746 1411 750
rect 1415 746 1419 750
rect 1455 746 1459 750
rect 1503 746 1507 750
rect 1519 746 1523 750
rect 1551 746 1555 750
rect 1599 746 1603 750
rect 1623 746 1627 750
rect 1655 746 1659 750
rect 1711 746 1715 750
rect 1719 746 1723 750
rect 1767 746 1771 750
rect 1815 746 1819 750
rect 1831 746 1835 750
rect 1895 746 1899 750
rect 1903 746 1907 750
rect 1959 746 1963 750
rect 1999 746 2003 750
rect 2023 746 2027 750
rect 2071 746 2075 750
rect 2119 746 2123 750
rect 111 726 115 730
rect 175 726 179 730
rect 215 726 219 730
rect 239 726 243 730
rect 279 726 283 730
rect 311 726 315 730
rect 351 726 355 730
rect 391 726 395 730
rect 423 726 427 730
rect 471 726 475 730
rect 495 726 499 730
rect 543 726 547 730
rect 567 726 571 730
rect 615 726 619 730
rect 639 726 643 730
rect 679 726 683 730
rect 703 726 707 730
rect 735 726 739 730
rect 759 726 763 730
rect 799 726 803 730
rect 815 726 819 730
rect 863 726 867 730
rect 911 726 915 730
rect 927 726 931 730
rect 959 726 963 730
rect 1007 726 1011 730
rect 1047 726 1051 730
rect 1095 726 1099 730
rect 1135 694 1139 698
rect 1247 694 1251 698
rect 1287 694 1291 698
rect 1335 694 1339 698
rect 1375 694 1379 698
rect 1391 694 1395 698
rect 1415 694 1419 698
rect 1447 694 1451 698
rect 1455 694 1459 698
rect 1503 694 1507 698
rect 1511 694 1515 698
rect 1551 694 1555 698
rect 1583 694 1587 698
rect 1599 694 1603 698
rect 1655 694 1659 698
rect 1711 694 1715 698
rect 1735 694 1739 698
rect 1767 694 1771 698
rect 1823 694 1827 698
rect 1831 694 1835 698
rect 1895 694 1899 698
rect 1911 694 1915 698
rect 1959 694 1963 698
rect 1999 694 2003 698
rect 2023 694 2027 698
rect 2071 694 2075 698
rect 2119 694 2123 698
rect 111 674 115 678
rect 135 674 139 678
rect 175 674 179 678
rect 215 674 219 678
rect 239 674 243 678
rect 271 674 275 678
rect 311 674 315 678
rect 335 674 339 678
rect 391 674 395 678
rect 399 674 403 678
rect 463 674 467 678
rect 471 674 475 678
rect 527 674 531 678
rect 543 674 547 678
rect 591 674 595 678
rect 615 674 619 678
rect 647 674 651 678
rect 679 674 683 678
rect 703 674 707 678
rect 735 674 739 678
rect 759 674 763 678
rect 799 674 803 678
rect 823 674 827 678
rect 863 674 867 678
rect 927 674 931 678
rect 1095 674 1099 678
rect 1135 642 1139 646
rect 1159 642 1163 646
rect 1199 642 1203 646
rect 1239 642 1243 646
rect 1247 642 1251 646
rect 1279 642 1283 646
rect 1287 642 1291 646
rect 1335 642 1339 646
rect 1343 642 1347 646
rect 1391 642 1395 646
rect 1415 642 1419 646
rect 1447 642 1451 646
rect 1495 642 1499 646
rect 1511 642 1515 646
rect 1583 642 1587 646
rect 1655 642 1659 646
rect 1671 642 1675 646
rect 1735 642 1739 646
rect 1759 642 1763 646
rect 1823 642 1827 646
rect 1839 642 1843 646
rect 1911 642 1915 646
rect 1919 642 1923 646
rect 1999 642 2003 646
rect 2007 642 2011 646
rect 2071 642 2075 646
rect 2119 642 2123 646
rect 111 614 115 618
rect 135 614 139 618
rect 175 614 179 618
rect 215 614 219 618
rect 255 614 259 618
rect 271 614 275 618
rect 303 614 307 618
rect 335 614 339 618
rect 351 614 355 618
rect 399 614 403 618
rect 439 614 443 618
rect 463 614 467 618
rect 487 614 491 618
rect 527 614 531 618
rect 535 614 539 618
rect 583 614 587 618
rect 591 614 595 618
rect 631 614 635 618
rect 647 614 651 618
rect 679 614 683 618
rect 703 614 707 618
rect 727 614 731 618
rect 759 614 763 618
rect 823 614 827 618
rect 1095 614 1099 618
rect 1135 586 1139 590
rect 1159 586 1163 590
rect 1199 586 1203 590
rect 1239 586 1243 590
rect 1279 586 1283 590
rect 1319 586 1323 590
rect 1343 586 1347 590
rect 1359 586 1363 590
rect 1415 586 1419 590
rect 1487 586 1491 590
rect 1495 586 1499 590
rect 1567 586 1571 590
rect 1583 586 1587 590
rect 1655 586 1659 590
rect 1671 586 1675 590
rect 1751 586 1755 590
rect 1759 586 1763 590
rect 1839 586 1843 590
rect 1855 586 1859 590
rect 1919 586 1923 590
rect 1967 586 1971 590
rect 2007 586 2011 590
rect 2071 586 2075 590
rect 2119 586 2123 590
rect 111 558 115 562
rect 135 558 139 562
rect 175 558 179 562
rect 215 558 219 562
rect 223 558 227 562
rect 255 558 259 562
rect 279 558 283 562
rect 303 558 307 562
rect 327 558 331 562
rect 351 558 355 562
rect 375 558 379 562
rect 399 558 403 562
rect 423 558 427 562
rect 439 558 443 562
rect 463 558 467 562
rect 487 558 491 562
rect 511 558 515 562
rect 535 558 539 562
rect 559 558 563 562
rect 583 558 587 562
rect 607 558 611 562
rect 631 558 635 562
rect 655 558 659 562
rect 679 558 683 562
rect 703 558 707 562
rect 727 558 731 562
rect 751 558 755 562
rect 1095 558 1099 562
rect 1135 530 1139 534
rect 1159 530 1163 534
rect 1199 530 1203 534
rect 1239 530 1243 534
rect 1279 530 1283 534
rect 1303 530 1307 534
rect 1319 530 1323 534
rect 1343 530 1347 534
rect 1359 530 1363 534
rect 1383 530 1387 534
rect 1415 530 1419 534
rect 1423 530 1427 534
rect 1463 530 1467 534
rect 1487 530 1491 534
rect 1503 530 1507 534
rect 1543 530 1547 534
rect 1567 530 1571 534
rect 1591 530 1595 534
rect 1647 530 1651 534
rect 1655 530 1659 534
rect 1703 530 1707 534
rect 1751 530 1755 534
rect 1767 530 1771 534
rect 1839 530 1843 534
rect 1855 530 1859 534
rect 1919 530 1923 534
rect 1967 530 1971 534
rect 2007 530 2011 534
rect 2071 530 2075 534
rect 2119 530 2123 534
rect 111 498 115 502
rect 135 498 139 502
rect 175 498 179 502
rect 223 498 227 502
rect 231 498 235 502
rect 279 498 283 502
rect 295 498 299 502
rect 327 498 331 502
rect 359 498 363 502
rect 375 498 379 502
rect 423 498 427 502
rect 463 498 467 502
rect 479 498 483 502
rect 511 498 515 502
rect 535 498 539 502
rect 559 498 563 502
rect 591 498 595 502
rect 607 498 611 502
rect 639 498 643 502
rect 655 498 659 502
rect 687 498 691 502
rect 703 498 707 502
rect 735 498 739 502
rect 751 498 755 502
rect 791 498 795 502
rect 847 498 851 502
rect 1095 498 1099 502
rect 1135 478 1139 482
rect 1295 478 1299 482
rect 1303 478 1307 482
rect 1335 478 1339 482
rect 1343 478 1347 482
rect 1375 478 1379 482
rect 1383 478 1387 482
rect 1423 478 1427 482
rect 1463 478 1467 482
rect 1471 478 1475 482
rect 1503 478 1507 482
rect 1527 478 1531 482
rect 1543 478 1547 482
rect 1583 478 1587 482
rect 1591 478 1595 482
rect 1647 478 1651 482
rect 1703 478 1707 482
rect 1719 478 1723 482
rect 1767 478 1771 482
rect 1807 478 1811 482
rect 1839 478 1843 482
rect 1895 478 1899 482
rect 1919 478 1923 482
rect 1991 478 1995 482
rect 2007 478 2011 482
rect 2071 478 2075 482
rect 2119 478 2123 482
rect 111 442 115 446
rect 135 442 139 446
rect 175 442 179 446
rect 215 442 219 446
rect 231 442 235 446
rect 263 442 267 446
rect 295 442 299 446
rect 327 442 331 446
rect 359 442 363 446
rect 391 442 395 446
rect 423 442 427 446
rect 463 442 467 446
rect 479 442 483 446
rect 535 442 539 446
rect 591 442 595 446
rect 607 442 611 446
rect 639 442 643 446
rect 679 442 683 446
rect 687 442 691 446
rect 735 442 739 446
rect 743 442 747 446
rect 791 442 795 446
rect 807 442 811 446
rect 847 442 851 446
rect 871 442 875 446
rect 943 442 947 446
rect 1095 442 1099 446
rect 1135 426 1139 430
rect 1159 426 1163 430
rect 1199 426 1203 430
rect 1255 426 1259 430
rect 1295 426 1299 430
rect 1335 426 1339 430
rect 1375 426 1379 430
rect 1415 426 1419 430
rect 1423 426 1427 430
rect 1471 426 1475 430
rect 1503 426 1507 430
rect 1527 426 1531 430
rect 1583 426 1587 430
rect 1591 426 1595 430
rect 1647 426 1651 430
rect 1671 426 1675 430
rect 1719 426 1723 430
rect 1751 426 1755 430
rect 1807 426 1811 430
rect 1831 426 1835 430
rect 1895 426 1899 430
rect 1911 426 1915 430
rect 1991 426 1995 430
rect 1999 426 2003 430
rect 2071 426 2075 430
rect 2119 426 2123 430
rect 111 382 115 386
rect 175 382 179 386
rect 215 382 219 386
rect 263 382 267 386
rect 271 382 275 386
rect 327 382 331 386
rect 335 382 339 386
rect 391 382 395 386
rect 407 382 411 386
rect 463 382 467 386
rect 487 382 491 386
rect 535 382 539 386
rect 567 382 571 386
rect 607 382 611 386
rect 639 382 643 386
rect 679 382 683 386
rect 711 382 715 386
rect 743 382 747 386
rect 775 382 779 386
rect 807 382 811 386
rect 839 382 843 386
rect 871 382 875 386
rect 895 382 899 386
rect 943 382 947 386
rect 951 382 955 386
rect 1007 382 1011 386
rect 1047 382 1051 386
rect 1095 382 1099 386
rect 1135 370 1139 374
rect 1159 370 1163 374
rect 1199 370 1203 374
rect 1247 370 1251 374
rect 1255 370 1259 374
rect 1335 370 1339 374
rect 1359 370 1363 374
rect 1415 370 1419 374
rect 1463 370 1467 374
rect 1503 370 1507 374
rect 1559 370 1563 374
rect 1591 370 1595 374
rect 1647 370 1651 374
rect 1671 370 1675 374
rect 1727 370 1731 374
rect 1751 370 1755 374
rect 1799 370 1803 374
rect 1831 370 1835 374
rect 1863 370 1867 374
rect 1911 370 1915 374
rect 1919 370 1923 374
rect 1975 370 1979 374
rect 1999 370 2003 374
rect 2031 370 2035 374
rect 2071 370 2075 374
rect 2119 370 2123 374
rect 111 326 115 330
rect 175 326 179 330
rect 215 326 219 330
rect 271 326 275 330
rect 335 326 339 330
rect 383 326 387 330
rect 407 326 411 330
rect 423 326 427 330
rect 463 326 467 330
rect 487 326 491 330
rect 503 326 507 330
rect 543 326 547 330
rect 567 326 571 330
rect 591 326 595 330
rect 639 326 643 330
rect 687 326 691 330
rect 711 326 715 330
rect 735 326 739 330
rect 775 326 779 330
rect 783 326 787 330
rect 831 326 835 330
rect 839 326 843 330
rect 879 326 883 330
rect 895 326 899 330
rect 927 326 931 330
rect 951 326 955 330
rect 967 326 971 330
rect 1007 326 1011 330
rect 1047 326 1051 330
rect 1095 326 1099 330
rect 1135 310 1139 314
rect 1159 310 1163 314
rect 1247 310 1251 314
rect 1351 310 1355 314
rect 1359 310 1363 314
rect 1391 310 1395 314
rect 1431 310 1435 314
rect 1463 310 1467 314
rect 1471 310 1475 314
rect 1511 310 1515 314
rect 1559 310 1563 314
rect 1615 310 1619 314
rect 1647 310 1651 314
rect 1671 310 1675 314
rect 1727 310 1731 314
rect 1735 310 1739 314
rect 1799 310 1803 314
rect 1807 310 1811 314
rect 1863 310 1867 314
rect 1887 310 1891 314
rect 1919 310 1923 314
rect 1967 310 1971 314
rect 1975 310 1979 314
rect 2031 310 2035 314
rect 2047 310 2051 314
rect 2071 310 2075 314
rect 2119 310 2123 314
rect 111 266 115 270
rect 287 266 291 270
rect 327 266 331 270
rect 367 266 371 270
rect 383 266 387 270
rect 415 266 419 270
rect 423 266 427 270
rect 463 266 467 270
rect 471 266 475 270
rect 503 266 507 270
rect 535 266 539 270
rect 543 266 547 270
rect 591 266 595 270
rect 607 266 611 270
rect 639 266 643 270
rect 679 266 683 270
rect 687 266 691 270
rect 735 266 739 270
rect 743 266 747 270
rect 783 266 787 270
rect 807 266 811 270
rect 831 266 835 270
rect 863 266 867 270
rect 879 266 883 270
rect 927 266 931 270
rect 967 266 971 270
rect 991 266 995 270
rect 1007 266 1011 270
rect 1047 266 1051 270
rect 1095 266 1099 270
rect 1135 258 1139 262
rect 1263 258 1267 262
rect 1303 258 1307 262
rect 1343 258 1347 262
rect 1351 258 1355 262
rect 1383 258 1387 262
rect 1391 258 1395 262
rect 1423 258 1427 262
rect 1431 258 1435 262
rect 1463 258 1467 262
rect 1471 258 1475 262
rect 1503 258 1507 262
rect 1511 258 1515 262
rect 1543 258 1547 262
rect 1559 258 1563 262
rect 1599 258 1603 262
rect 1615 258 1619 262
rect 1671 258 1675 262
rect 1735 258 1739 262
rect 1759 258 1763 262
rect 1807 258 1811 262
rect 1863 258 1867 262
rect 1887 258 1891 262
rect 1967 258 1971 262
rect 1975 258 1979 262
rect 2047 258 2051 262
rect 2071 258 2075 262
rect 2119 258 2123 262
rect 111 202 115 206
rect 167 202 171 206
rect 207 202 211 206
rect 247 202 251 206
rect 287 202 291 206
rect 295 202 299 206
rect 327 202 331 206
rect 343 202 347 206
rect 367 202 371 206
rect 399 202 403 206
rect 415 202 419 206
rect 463 202 467 206
rect 471 202 475 206
rect 527 202 531 206
rect 535 202 539 206
rect 599 202 603 206
rect 607 202 611 206
rect 671 202 675 206
rect 679 202 683 206
rect 743 202 747 206
rect 751 202 755 206
rect 807 202 811 206
rect 831 202 835 206
rect 863 202 867 206
rect 911 202 915 206
rect 927 202 931 206
rect 991 202 995 206
rect 1047 202 1051 206
rect 1095 202 1099 206
rect 1135 202 1139 206
rect 1183 202 1187 206
rect 1231 202 1235 206
rect 1263 202 1267 206
rect 1295 202 1299 206
rect 1303 202 1307 206
rect 1343 202 1347 206
rect 1359 202 1363 206
rect 1383 202 1387 206
rect 1423 202 1427 206
rect 1431 202 1435 206
rect 1463 202 1467 206
rect 1503 202 1507 206
rect 1511 202 1515 206
rect 1543 202 1547 206
rect 1591 202 1595 206
rect 1599 202 1603 206
rect 1663 202 1667 206
rect 1671 202 1675 206
rect 1735 202 1739 206
rect 1759 202 1763 206
rect 1807 202 1811 206
rect 1863 202 1867 206
rect 1879 202 1883 206
rect 1951 202 1955 206
rect 1975 202 1979 206
rect 2023 202 2027 206
rect 2071 202 2075 206
rect 2119 202 2123 206
rect 111 134 115 138
rect 135 134 139 138
rect 167 134 171 138
rect 175 134 179 138
rect 207 134 211 138
rect 215 134 219 138
rect 247 134 251 138
rect 255 134 259 138
rect 295 134 299 138
rect 335 134 339 138
rect 343 134 347 138
rect 375 134 379 138
rect 399 134 403 138
rect 415 134 419 138
rect 455 134 459 138
rect 463 134 467 138
rect 495 134 499 138
rect 527 134 531 138
rect 535 134 539 138
rect 575 134 579 138
rect 599 134 603 138
rect 615 134 619 138
rect 655 134 659 138
rect 671 134 675 138
rect 695 134 699 138
rect 735 134 739 138
rect 751 134 755 138
rect 775 134 779 138
rect 815 134 819 138
rect 831 134 835 138
rect 871 134 875 138
rect 911 134 915 138
rect 935 134 939 138
rect 991 134 995 138
rect 999 134 1003 138
rect 1047 134 1051 138
rect 1095 134 1099 138
rect 1135 126 1139 130
rect 1159 126 1163 130
rect 1183 126 1187 130
rect 1199 126 1203 130
rect 1231 126 1235 130
rect 1239 126 1243 130
rect 1279 126 1283 130
rect 1295 126 1299 130
rect 1319 126 1323 130
rect 1359 126 1363 130
rect 1367 126 1371 130
rect 1431 126 1435 130
rect 1495 126 1499 130
rect 1511 126 1515 130
rect 1559 126 1563 130
rect 1591 126 1595 130
rect 1615 126 1619 130
rect 1663 126 1667 130
rect 1671 126 1675 130
rect 1719 126 1723 130
rect 1735 126 1739 130
rect 1767 126 1771 130
rect 1807 126 1811 130
rect 1855 126 1859 130
rect 1879 126 1883 130
rect 1903 126 1907 130
rect 1951 126 1955 130
rect 1991 126 1995 130
rect 2023 126 2027 130
rect 2031 126 2035 130
rect 2071 126 2075 130
rect 2119 126 2123 130
rect 111 82 115 86
rect 135 82 139 86
rect 175 82 179 86
rect 215 82 219 86
rect 255 82 259 86
rect 295 82 299 86
rect 335 82 339 86
rect 375 82 379 86
rect 415 82 419 86
rect 455 82 459 86
rect 495 82 499 86
rect 535 82 539 86
rect 575 82 579 86
rect 615 82 619 86
rect 655 82 659 86
rect 695 82 699 86
rect 735 82 739 86
rect 775 82 779 86
rect 815 82 819 86
rect 871 82 875 86
rect 935 82 939 86
rect 999 82 1003 86
rect 1047 82 1051 86
rect 1095 82 1099 86
rect 1135 74 1139 78
rect 1159 74 1163 78
rect 1199 74 1203 78
rect 1239 74 1243 78
rect 1279 74 1283 78
rect 1319 74 1323 78
rect 1367 74 1371 78
rect 1431 74 1435 78
rect 1495 74 1499 78
rect 1559 74 1563 78
rect 1615 74 1619 78
rect 1671 74 1675 78
rect 1719 74 1723 78
rect 1767 74 1771 78
rect 1807 74 1811 78
rect 1855 74 1859 78
rect 1903 74 1907 78
rect 1951 74 1955 78
rect 1991 74 1995 78
rect 2031 74 2035 78
rect 2071 74 2075 78
rect 2119 74 2123 78
<< m4 >>
rect 1118 2209 1119 2215
rect 1125 2214 2155 2215
rect 1125 2210 1135 2214
rect 1139 2210 1343 2214
rect 1347 2210 1383 2214
rect 1387 2210 1423 2214
rect 1427 2210 1463 2214
rect 1467 2210 1503 2214
rect 1507 2210 1543 2214
rect 1547 2210 1583 2214
rect 1587 2210 1623 2214
rect 1627 2210 1663 2214
rect 1667 2210 1703 2214
rect 1707 2210 1743 2214
rect 1747 2210 1783 2214
rect 1787 2210 1823 2214
rect 1827 2210 2119 2214
rect 2123 2210 2155 2214
rect 1125 2209 2155 2210
rect 2161 2209 2162 2215
rect 1106 2157 1107 2163
rect 1113 2162 2143 2163
rect 1113 2158 1135 2162
rect 1139 2158 1287 2162
rect 1291 2158 1327 2162
rect 1331 2158 1343 2162
rect 1347 2158 1367 2162
rect 1371 2158 1383 2162
rect 1387 2158 1415 2162
rect 1419 2158 1423 2162
rect 1427 2158 1463 2162
rect 1467 2158 1503 2162
rect 1507 2158 1519 2162
rect 1523 2158 1543 2162
rect 1547 2158 1575 2162
rect 1579 2158 1583 2162
rect 1587 2158 1623 2162
rect 1627 2158 1663 2162
rect 1667 2158 1671 2162
rect 1675 2158 1703 2162
rect 1707 2158 1719 2162
rect 1723 2158 1743 2162
rect 1747 2158 1775 2162
rect 1779 2158 1783 2162
rect 1787 2158 1823 2162
rect 1827 2158 1831 2162
rect 1835 2158 1887 2162
rect 1891 2158 2119 2162
rect 2123 2158 2143 2162
rect 1113 2157 2143 2158
rect 2149 2157 2150 2163
rect 1118 2101 1119 2107
rect 1125 2106 2155 2107
rect 1125 2102 1135 2106
rect 1139 2102 1223 2106
rect 1227 2102 1279 2106
rect 1283 2102 1287 2106
rect 1291 2102 1327 2106
rect 1331 2102 1343 2106
rect 1347 2102 1367 2106
rect 1371 2102 1415 2106
rect 1419 2102 1423 2106
rect 1427 2102 1463 2106
rect 1467 2102 1503 2106
rect 1507 2102 1519 2106
rect 1523 2102 1575 2106
rect 1579 2102 1583 2106
rect 1587 2102 1623 2106
rect 1627 2102 1663 2106
rect 1667 2102 1671 2106
rect 1675 2102 1719 2106
rect 1723 2102 1743 2106
rect 1747 2102 1775 2106
rect 1779 2102 1831 2106
rect 1835 2102 1887 2106
rect 1891 2102 1919 2106
rect 1923 2102 2007 2106
rect 2011 2102 2071 2106
rect 2075 2102 2119 2106
rect 2123 2102 2155 2106
rect 1125 2101 2155 2102
rect 2161 2101 2162 2107
rect 1106 2049 1107 2055
rect 1113 2054 2143 2055
rect 1113 2050 1135 2054
rect 1139 2050 1183 2054
rect 1187 2050 1223 2054
rect 1227 2050 1239 2054
rect 1243 2050 1279 2054
rect 1283 2050 1311 2054
rect 1315 2050 1343 2054
rect 1347 2050 1399 2054
rect 1403 2050 1423 2054
rect 1427 2050 1487 2054
rect 1491 2050 1503 2054
rect 1507 2050 1583 2054
rect 1587 2050 1663 2054
rect 1667 2050 1671 2054
rect 1675 2050 1743 2054
rect 1747 2050 1759 2054
rect 1763 2050 1831 2054
rect 1835 2050 1839 2054
rect 1843 2050 1919 2054
rect 1923 2050 2007 2054
rect 2011 2050 2071 2054
rect 2075 2050 2119 2054
rect 2123 2050 2143 2054
rect 1113 2049 2143 2050
rect 2149 2049 2150 2055
rect 96 2029 97 2035
rect 103 2034 1119 2035
rect 103 2030 111 2034
rect 115 2030 191 2034
rect 195 2030 231 2034
rect 235 2030 287 2034
rect 291 2030 351 2034
rect 355 2030 423 2034
rect 427 2030 495 2034
rect 499 2030 575 2034
rect 579 2030 647 2034
rect 651 2030 719 2034
rect 723 2030 783 2034
rect 787 2030 839 2034
rect 843 2030 895 2034
rect 899 2030 951 2034
rect 955 2030 1007 2034
rect 1011 2030 1047 2034
rect 1051 2030 1095 2034
rect 1099 2030 1119 2034
rect 103 2029 1119 2030
rect 1125 2029 1126 2035
rect 1118 1997 1119 2003
rect 1125 2002 2155 2003
rect 1125 1998 1135 2002
rect 1139 1998 1183 2002
rect 1187 1998 1239 2002
rect 1243 1998 1303 2002
rect 1307 1998 1311 2002
rect 1315 1998 1383 2002
rect 1387 1998 1399 2002
rect 1403 1998 1463 2002
rect 1467 1998 1487 2002
rect 1491 1998 1543 2002
rect 1547 1998 1583 2002
rect 1587 1998 1615 2002
rect 1619 1998 1671 2002
rect 1675 1998 1687 2002
rect 1691 1998 1751 2002
rect 1755 1998 1759 2002
rect 1763 1998 1815 2002
rect 1819 1998 1839 2002
rect 1843 1998 1879 2002
rect 1883 1998 1919 2002
rect 1923 1998 1951 2002
rect 1955 1998 2007 2002
rect 2011 1998 2023 2002
rect 2027 1998 2071 2002
rect 2075 1998 2119 2002
rect 2123 1998 2155 2002
rect 1125 1997 2155 1998
rect 2161 1997 2162 2003
rect 84 1977 85 1983
rect 91 1982 1107 1983
rect 91 1978 111 1982
rect 115 1978 191 1982
rect 195 1978 231 1982
rect 235 1978 247 1982
rect 251 1978 287 1982
rect 291 1978 311 1982
rect 315 1978 351 1982
rect 355 1978 375 1982
rect 379 1978 423 1982
rect 427 1978 447 1982
rect 451 1978 495 1982
rect 499 1978 519 1982
rect 523 1978 575 1982
rect 579 1978 591 1982
rect 595 1978 647 1982
rect 651 1978 655 1982
rect 659 1978 719 1982
rect 723 1978 775 1982
rect 779 1978 783 1982
rect 787 1978 823 1982
rect 827 1978 839 1982
rect 843 1978 871 1982
rect 875 1978 895 1982
rect 899 1978 919 1982
rect 923 1978 951 1982
rect 955 1978 967 1982
rect 971 1978 1007 1982
rect 1011 1978 1047 1982
rect 1051 1978 1095 1982
rect 1099 1978 1107 1982
rect 91 1977 1107 1978
rect 1113 1977 1114 1983
rect 1106 1941 1107 1947
rect 1113 1946 2143 1947
rect 1113 1942 1135 1946
rect 1139 1942 1159 1946
rect 1163 1942 1223 1946
rect 1227 1942 1303 1946
rect 1307 1942 1383 1946
rect 1387 1942 1463 1946
rect 1467 1942 1535 1946
rect 1539 1942 1543 1946
rect 1547 1942 1615 1946
rect 1619 1942 1687 1946
rect 1691 1942 1695 1946
rect 1699 1942 1751 1946
rect 1755 1942 1783 1946
rect 1787 1942 1815 1946
rect 1819 1942 1879 1946
rect 1883 1942 1951 1946
rect 1955 1942 1983 1946
rect 1987 1942 2023 1946
rect 2027 1942 2071 1946
rect 2075 1942 2119 1946
rect 2123 1942 2143 1946
rect 1113 1941 2143 1942
rect 2149 1941 2150 1947
rect 96 1925 97 1931
rect 103 1930 1119 1931
rect 103 1926 111 1930
rect 115 1926 135 1930
rect 139 1926 175 1930
rect 179 1926 191 1930
rect 195 1926 231 1930
rect 235 1926 247 1930
rect 251 1926 295 1930
rect 299 1926 311 1930
rect 315 1926 367 1930
rect 371 1926 375 1930
rect 379 1926 431 1930
rect 435 1926 447 1930
rect 451 1926 495 1930
rect 499 1926 519 1930
rect 523 1926 559 1930
rect 563 1926 591 1930
rect 595 1926 615 1930
rect 619 1926 655 1930
rect 659 1926 671 1930
rect 675 1926 719 1930
rect 723 1926 727 1930
rect 731 1926 775 1930
rect 779 1926 783 1930
rect 787 1926 823 1930
rect 827 1926 847 1930
rect 851 1926 871 1930
rect 875 1926 919 1930
rect 923 1926 967 1930
rect 971 1926 1007 1930
rect 1011 1926 1047 1930
rect 1051 1926 1095 1930
rect 1099 1926 1119 1930
rect 103 1925 1119 1926
rect 1125 1925 1126 1931
rect 1118 1885 1119 1891
rect 1125 1890 2155 1891
rect 1125 1886 1135 1890
rect 1139 1886 1159 1890
rect 1163 1886 1199 1890
rect 1203 1886 1223 1890
rect 1227 1886 1263 1890
rect 1267 1886 1303 1890
rect 1307 1886 1327 1890
rect 1331 1886 1383 1890
rect 1387 1886 1391 1890
rect 1395 1886 1447 1890
rect 1451 1886 1463 1890
rect 1467 1886 1503 1890
rect 1507 1886 1535 1890
rect 1539 1886 1559 1890
rect 1563 1886 1615 1890
rect 1619 1886 1631 1890
rect 1635 1886 1695 1890
rect 1699 1886 1711 1890
rect 1715 1886 1783 1890
rect 1787 1886 1799 1890
rect 1803 1886 1879 1890
rect 1883 1886 1895 1890
rect 1899 1886 1983 1890
rect 1987 1886 1991 1890
rect 1995 1886 2071 1890
rect 2075 1886 2119 1890
rect 2123 1886 2155 1890
rect 1125 1885 2155 1886
rect 2161 1885 2162 1891
rect 84 1869 85 1875
rect 91 1874 1107 1875
rect 91 1870 111 1874
rect 115 1870 135 1874
rect 139 1870 175 1874
rect 179 1870 199 1874
rect 203 1870 231 1874
rect 235 1870 271 1874
rect 275 1870 295 1874
rect 299 1870 335 1874
rect 339 1870 367 1874
rect 371 1870 399 1874
rect 403 1870 431 1874
rect 435 1870 455 1874
rect 459 1870 495 1874
rect 499 1870 503 1874
rect 507 1870 551 1874
rect 555 1870 559 1874
rect 563 1870 599 1874
rect 603 1870 615 1874
rect 619 1870 647 1874
rect 651 1870 671 1874
rect 675 1870 695 1874
rect 699 1870 727 1874
rect 731 1870 751 1874
rect 755 1870 783 1874
rect 787 1870 847 1874
rect 851 1870 1095 1874
rect 1099 1870 1107 1874
rect 91 1869 1107 1870
rect 1113 1869 1114 1875
rect 1106 1833 1107 1839
rect 1113 1838 2143 1839
rect 1113 1834 1135 1838
rect 1139 1834 1159 1838
rect 1163 1834 1199 1838
rect 1203 1834 1231 1838
rect 1235 1834 1263 1838
rect 1267 1834 1303 1838
rect 1307 1834 1327 1838
rect 1331 1834 1383 1838
rect 1387 1834 1391 1838
rect 1395 1834 1447 1838
rect 1451 1834 1463 1838
rect 1467 1834 1503 1838
rect 1507 1834 1551 1838
rect 1555 1834 1559 1838
rect 1563 1834 1631 1838
rect 1635 1834 1647 1838
rect 1651 1834 1711 1838
rect 1715 1834 1751 1838
rect 1755 1834 1799 1838
rect 1803 1834 1855 1838
rect 1859 1834 1895 1838
rect 1899 1834 1967 1838
rect 1971 1834 1991 1838
rect 1995 1834 2071 1838
rect 2075 1834 2119 1838
rect 2123 1834 2143 1838
rect 1113 1833 2143 1834
rect 2149 1833 2150 1839
rect 96 1809 97 1815
rect 103 1814 1119 1815
rect 103 1810 111 1814
rect 115 1810 135 1814
rect 139 1810 151 1814
rect 155 1810 199 1814
rect 203 1810 215 1814
rect 219 1810 271 1814
rect 275 1810 327 1814
rect 331 1810 335 1814
rect 339 1810 383 1814
rect 387 1810 399 1814
rect 403 1810 431 1814
rect 435 1810 455 1814
rect 459 1810 479 1814
rect 483 1810 503 1814
rect 507 1810 527 1814
rect 531 1810 551 1814
rect 555 1810 575 1814
rect 579 1810 599 1814
rect 603 1810 623 1814
rect 627 1810 647 1814
rect 651 1810 671 1814
rect 675 1810 695 1814
rect 699 1810 727 1814
rect 731 1810 751 1814
rect 755 1810 1095 1814
rect 1099 1810 1119 1814
rect 103 1809 1119 1810
rect 1125 1809 1126 1815
rect 1118 1781 1119 1787
rect 1125 1786 2155 1787
rect 1125 1782 1135 1786
rect 1139 1782 1159 1786
rect 1163 1782 1191 1786
rect 1195 1782 1231 1786
rect 1235 1782 1255 1786
rect 1259 1782 1303 1786
rect 1307 1782 1319 1786
rect 1323 1782 1383 1786
rect 1387 1782 1455 1786
rect 1459 1782 1463 1786
rect 1467 1782 1527 1786
rect 1531 1782 1551 1786
rect 1555 1782 1607 1786
rect 1611 1782 1647 1786
rect 1651 1782 1687 1786
rect 1691 1782 1751 1786
rect 1755 1782 1767 1786
rect 1771 1782 1847 1786
rect 1851 1782 1855 1786
rect 1859 1782 1927 1786
rect 1931 1782 1967 1786
rect 1971 1782 2007 1786
rect 2011 1782 2071 1786
rect 2075 1782 2119 1786
rect 2123 1782 2155 1786
rect 1125 1781 2155 1782
rect 2161 1781 2162 1787
rect 84 1757 85 1763
rect 91 1762 1107 1763
rect 91 1758 111 1762
rect 115 1758 151 1762
rect 155 1758 215 1762
rect 219 1758 231 1762
rect 235 1758 271 1762
rect 275 1758 295 1762
rect 299 1758 327 1762
rect 331 1758 351 1762
rect 355 1758 383 1762
rect 387 1758 415 1762
rect 419 1758 431 1762
rect 435 1758 479 1762
rect 483 1758 527 1762
rect 531 1758 543 1762
rect 547 1758 575 1762
rect 579 1758 615 1762
rect 619 1758 623 1762
rect 627 1758 671 1762
rect 675 1758 687 1762
rect 691 1758 727 1762
rect 731 1758 759 1762
rect 763 1758 831 1762
rect 835 1758 911 1762
rect 915 1758 991 1762
rect 995 1758 1095 1762
rect 1099 1758 1107 1762
rect 91 1757 1107 1758
rect 1113 1757 1114 1763
rect 1106 1729 1107 1735
rect 1113 1734 2143 1735
rect 1113 1730 1135 1734
rect 1139 1730 1191 1734
rect 1195 1730 1247 1734
rect 1251 1730 1255 1734
rect 1259 1730 1295 1734
rect 1299 1730 1319 1734
rect 1323 1730 1343 1734
rect 1347 1730 1383 1734
rect 1387 1730 1399 1734
rect 1403 1730 1455 1734
rect 1459 1730 1463 1734
rect 1467 1730 1527 1734
rect 1531 1730 1599 1734
rect 1603 1730 1607 1734
rect 1611 1730 1671 1734
rect 1675 1730 1687 1734
rect 1691 1730 1743 1734
rect 1747 1730 1767 1734
rect 1771 1730 1807 1734
rect 1811 1730 1847 1734
rect 1851 1730 1879 1734
rect 1883 1730 1927 1734
rect 1931 1730 1951 1734
rect 1955 1730 2007 1734
rect 2011 1730 2023 1734
rect 2027 1730 2071 1734
rect 2075 1730 2119 1734
rect 2123 1730 2143 1734
rect 1113 1729 2143 1730
rect 2149 1729 2150 1735
rect 96 1701 97 1707
rect 103 1706 1119 1707
rect 103 1702 111 1706
rect 115 1702 135 1706
rect 139 1702 199 1706
rect 203 1702 231 1706
rect 235 1702 279 1706
rect 283 1702 295 1706
rect 299 1702 351 1706
rect 355 1702 367 1706
rect 371 1702 415 1706
rect 419 1702 463 1706
rect 467 1702 479 1706
rect 483 1702 543 1706
rect 547 1702 551 1706
rect 555 1702 615 1706
rect 619 1702 639 1706
rect 643 1702 687 1706
rect 691 1702 719 1706
rect 723 1702 759 1706
rect 763 1702 791 1706
rect 795 1702 831 1706
rect 835 1702 855 1706
rect 859 1702 911 1706
rect 915 1702 919 1706
rect 923 1702 983 1706
rect 987 1702 991 1706
rect 995 1702 1047 1706
rect 1051 1702 1095 1706
rect 1099 1702 1119 1706
rect 103 1701 1119 1702
rect 1125 1701 1126 1707
rect 1118 1673 1119 1679
rect 1125 1678 2155 1679
rect 1125 1674 1135 1678
rect 1139 1674 1247 1678
rect 1251 1674 1263 1678
rect 1267 1674 1295 1678
rect 1299 1674 1303 1678
rect 1307 1674 1343 1678
rect 1347 1674 1391 1678
rect 1395 1674 1399 1678
rect 1403 1674 1447 1678
rect 1451 1674 1463 1678
rect 1467 1674 1503 1678
rect 1507 1674 1527 1678
rect 1531 1674 1567 1678
rect 1571 1674 1599 1678
rect 1603 1674 1631 1678
rect 1635 1674 1671 1678
rect 1675 1674 1695 1678
rect 1699 1674 1743 1678
rect 1747 1674 1759 1678
rect 1763 1674 1807 1678
rect 1811 1674 1831 1678
rect 1835 1674 1879 1678
rect 1883 1674 1911 1678
rect 1915 1674 1951 1678
rect 1955 1674 1999 1678
rect 2003 1674 2023 1678
rect 2027 1674 2071 1678
rect 2075 1674 2119 1678
rect 2123 1674 2155 1678
rect 1125 1673 2155 1674
rect 2161 1673 2162 1679
rect 84 1645 85 1651
rect 91 1650 1107 1651
rect 91 1646 111 1650
rect 115 1646 135 1650
rect 139 1646 183 1650
rect 187 1646 199 1650
rect 203 1646 263 1650
rect 267 1646 279 1650
rect 283 1646 343 1650
rect 347 1646 367 1650
rect 371 1646 423 1650
rect 427 1646 463 1650
rect 467 1646 503 1650
rect 507 1646 551 1650
rect 555 1646 583 1650
rect 587 1646 639 1650
rect 643 1646 655 1650
rect 659 1646 719 1650
rect 723 1646 727 1650
rect 731 1646 791 1650
rect 795 1646 847 1650
rect 851 1646 855 1650
rect 859 1646 903 1650
rect 907 1646 919 1650
rect 923 1646 959 1650
rect 963 1646 983 1650
rect 987 1646 1007 1650
rect 1011 1646 1047 1650
rect 1051 1646 1095 1650
rect 1099 1646 1107 1650
rect 91 1645 1107 1646
rect 1113 1645 1114 1651
rect 1106 1609 1107 1615
rect 1113 1614 2143 1615
rect 1113 1610 1135 1614
rect 1139 1610 1159 1614
rect 1163 1610 1215 1614
rect 1219 1610 1263 1614
rect 1267 1610 1303 1614
rect 1307 1610 1343 1614
rect 1347 1610 1383 1614
rect 1387 1610 1391 1614
rect 1395 1610 1447 1614
rect 1451 1610 1463 1614
rect 1467 1610 1503 1614
rect 1507 1610 1543 1614
rect 1547 1610 1567 1614
rect 1571 1610 1623 1614
rect 1627 1610 1631 1614
rect 1635 1610 1695 1614
rect 1699 1610 1711 1614
rect 1715 1610 1759 1614
rect 1763 1610 1799 1614
rect 1803 1610 1831 1614
rect 1835 1610 1887 1614
rect 1891 1610 1911 1614
rect 1915 1610 1983 1614
rect 1987 1610 1999 1614
rect 2003 1610 2071 1614
rect 2075 1610 2119 1614
rect 2123 1610 2143 1614
rect 1113 1609 2143 1610
rect 2149 1609 2150 1615
rect 96 1593 97 1599
rect 103 1598 1119 1599
rect 103 1594 111 1598
rect 115 1594 135 1598
rect 139 1594 175 1598
rect 179 1594 183 1598
rect 187 1594 231 1598
rect 235 1594 263 1598
rect 267 1594 303 1598
rect 307 1594 343 1598
rect 347 1594 375 1598
rect 379 1594 423 1598
rect 427 1594 455 1598
rect 459 1594 503 1598
rect 507 1594 527 1598
rect 531 1594 583 1598
rect 587 1594 599 1598
rect 603 1594 655 1598
rect 659 1594 671 1598
rect 675 1594 727 1598
rect 731 1594 743 1598
rect 747 1594 791 1598
rect 795 1594 815 1598
rect 819 1594 847 1598
rect 851 1594 887 1598
rect 891 1594 903 1598
rect 907 1594 959 1598
rect 963 1594 1007 1598
rect 1011 1594 1047 1598
rect 1051 1594 1095 1598
rect 1099 1594 1119 1598
rect 103 1593 1119 1594
rect 1125 1593 1126 1599
rect 1118 1557 1119 1563
rect 1125 1562 2155 1563
rect 1125 1558 1135 1562
rect 1139 1558 1159 1562
rect 1163 1558 1199 1562
rect 1203 1558 1215 1562
rect 1219 1558 1247 1562
rect 1251 1558 1303 1562
rect 1307 1558 1319 1562
rect 1323 1558 1383 1562
rect 1387 1558 1399 1562
rect 1403 1558 1463 1562
rect 1467 1558 1479 1562
rect 1483 1558 1543 1562
rect 1547 1558 1559 1562
rect 1563 1558 1623 1562
rect 1627 1558 1647 1562
rect 1651 1558 1711 1562
rect 1715 1558 1735 1562
rect 1739 1558 1799 1562
rect 1803 1558 1823 1562
rect 1827 1558 1887 1562
rect 1891 1558 1911 1562
rect 1915 1558 1983 1562
rect 1987 1558 1999 1562
rect 2003 1558 2071 1562
rect 2075 1558 2119 1562
rect 2123 1558 2155 1562
rect 1125 1557 2155 1558
rect 2161 1557 2162 1563
rect 84 1541 85 1547
rect 91 1546 1107 1547
rect 91 1542 111 1546
rect 115 1542 135 1546
rect 139 1542 175 1546
rect 179 1542 231 1546
rect 235 1542 303 1546
rect 307 1542 311 1546
rect 315 1542 375 1546
rect 379 1542 391 1546
rect 395 1542 455 1546
rect 459 1542 479 1546
rect 483 1542 527 1546
rect 531 1542 567 1546
rect 571 1542 599 1546
rect 603 1542 655 1546
rect 659 1542 671 1546
rect 675 1542 743 1546
rect 747 1542 815 1546
rect 819 1542 823 1546
rect 827 1542 887 1546
rect 891 1542 911 1546
rect 915 1542 999 1546
rect 1003 1542 1095 1546
rect 1099 1542 1107 1546
rect 91 1541 1107 1542
rect 1113 1541 1114 1547
rect 1106 1505 1107 1511
rect 1113 1510 2143 1511
rect 1113 1506 1135 1510
rect 1139 1506 1159 1510
rect 1163 1506 1199 1510
rect 1203 1506 1239 1510
rect 1243 1506 1247 1510
rect 1251 1506 1303 1510
rect 1307 1506 1319 1510
rect 1323 1506 1375 1510
rect 1379 1506 1399 1510
rect 1403 1506 1455 1510
rect 1459 1506 1479 1510
rect 1483 1506 1543 1510
rect 1547 1506 1559 1510
rect 1563 1506 1623 1510
rect 1627 1506 1647 1510
rect 1651 1506 1703 1510
rect 1707 1506 1735 1510
rect 1739 1506 1775 1510
rect 1779 1506 1823 1510
rect 1827 1506 1847 1510
rect 1851 1506 1911 1510
rect 1915 1506 1919 1510
rect 1923 1506 1991 1510
rect 1995 1506 1999 1510
rect 2003 1506 2063 1510
rect 2067 1506 2071 1510
rect 2075 1506 2119 1510
rect 2123 1506 2143 1510
rect 1113 1505 2143 1506
rect 2149 1505 2150 1511
rect 96 1489 97 1495
rect 103 1494 1119 1495
rect 103 1490 111 1494
rect 115 1490 135 1494
rect 139 1490 175 1494
rect 179 1490 199 1494
rect 203 1490 231 1494
rect 235 1490 279 1494
rect 283 1490 311 1494
rect 315 1490 359 1494
rect 363 1490 391 1494
rect 395 1490 439 1494
rect 443 1490 479 1494
rect 483 1490 519 1494
rect 523 1490 567 1494
rect 571 1490 599 1494
rect 603 1490 655 1494
rect 659 1490 679 1494
rect 683 1490 743 1494
rect 747 1490 767 1494
rect 771 1490 823 1494
rect 827 1490 855 1494
rect 859 1490 911 1494
rect 915 1490 943 1494
rect 947 1490 999 1494
rect 1003 1490 1031 1494
rect 1035 1490 1095 1494
rect 1099 1490 1119 1494
rect 103 1489 1119 1490
rect 1125 1489 1126 1495
rect 1118 1449 1119 1455
rect 1125 1454 2155 1455
rect 1125 1450 1135 1454
rect 1139 1450 1159 1454
rect 1163 1450 1199 1454
rect 1203 1450 1239 1454
rect 1243 1450 1279 1454
rect 1283 1450 1303 1454
rect 1307 1450 1327 1454
rect 1331 1450 1375 1454
rect 1379 1450 1383 1454
rect 1387 1450 1439 1454
rect 1443 1450 1455 1454
rect 1459 1450 1495 1454
rect 1499 1450 1543 1454
rect 1547 1450 1551 1454
rect 1555 1450 1607 1454
rect 1611 1450 1623 1454
rect 1627 1450 1671 1454
rect 1675 1450 1703 1454
rect 1707 1450 1735 1454
rect 1739 1450 1775 1454
rect 1779 1450 1807 1454
rect 1811 1450 1847 1454
rect 1851 1450 1887 1454
rect 1891 1450 1919 1454
rect 1923 1450 1975 1454
rect 1979 1450 1991 1454
rect 1995 1450 2063 1454
rect 2067 1450 2119 1454
rect 2123 1450 2155 1454
rect 1125 1449 2155 1450
rect 2161 1449 2162 1455
rect 84 1437 85 1443
rect 91 1442 1107 1443
rect 91 1438 111 1442
rect 115 1438 135 1442
rect 139 1438 191 1442
rect 195 1438 199 1442
rect 203 1438 263 1442
rect 267 1438 279 1442
rect 283 1438 335 1442
rect 339 1438 359 1442
rect 363 1438 407 1442
rect 411 1438 439 1442
rect 443 1438 479 1442
rect 483 1438 519 1442
rect 523 1438 551 1442
rect 555 1438 599 1442
rect 603 1438 631 1442
rect 635 1438 679 1442
rect 683 1438 711 1442
rect 715 1438 767 1442
rect 771 1438 799 1442
rect 803 1438 855 1442
rect 859 1438 887 1442
rect 891 1438 943 1442
rect 947 1438 975 1442
rect 979 1438 1031 1442
rect 1035 1438 1047 1442
rect 1051 1438 1095 1442
rect 1099 1438 1107 1442
rect 91 1437 1107 1438
rect 1113 1437 1114 1443
rect 1106 1395 1107 1401
rect 1113 1399 1138 1401
rect 1113 1398 2143 1399
rect 1113 1395 1135 1398
rect 1132 1394 1135 1395
rect 1139 1394 1279 1398
rect 1283 1394 1327 1398
rect 1331 1394 1335 1398
rect 1339 1394 1375 1398
rect 1379 1394 1383 1398
rect 1387 1394 1415 1398
rect 1419 1394 1439 1398
rect 1443 1394 1455 1398
rect 1459 1394 1495 1398
rect 1499 1394 1535 1398
rect 1539 1394 1551 1398
rect 1555 1394 1583 1398
rect 1587 1394 1607 1398
rect 1611 1394 1647 1398
rect 1651 1394 1671 1398
rect 1675 1394 1719 1398
rect 1723 1394 1735 1398
rect 1739 1394 1807 1398
rect 1811 1394 1887 1398
rect 1891 1394 1895 1398
rect 1899 1394 1975 1398
rect 1979 1394 1991 1398
rect 1995 1394 2063 1398
rect 2067 1394 2071 1398
rect 2075 1394 2119 1398
rect 2123 1394 2143 1398
rect 1132 1393 2143 1394
rect 2149 1393 2150 1399
rect 96 1385 97 1391
rect 103 1390 1119 1391
rect 103 1386 111 1390
rect 115 1386 135 1390
rect 139 1386 175 1390
rect 179 1386 191 1390
rect 195 1386 239 1390
rect 243 1386 263 1390
rect 267 1386 303 1390
rect 307 1386 335 1390
rect 339 1386 367 1390
rect 371 1386 407 1390
rect 411 1386 439 1390
rect 443 1386 479 1390
rect 483 1386 503 1390
rect 507 1386 551 1390
rect 555 1386 575 1390
rect 579 1386 631 1390
rect 635 1386 647 1390
rect 651 1386 711 1390
rect 715 1386 783 1390
rect 787 1386 799 1390
rect 803 1386 855 1390
rect 859 1386 887 1390
rect 891 1386 927 1390
rect 931 1386 975 1390
rect 979 1386 999 1390
rect 1003 1386 1047 1390
rect 1051 1386 1095 1390
rect 1099 1386 1119 1390
rect 103 1385 1119 1386
rect 1125 1385 1126 1391
rect 1118 1341 1119 1347
rect 1125 1346 2155 1347
rect 1125 1342 1135 1346
rect 1139 1342 1159 1346
rect 1163 1342 1223 1346
rect 1227 1342 1311 1346
rect 1315 1342 1335 1346
rect 1339 1342 1375 1346
rect 1379 1342 1407 1346
rect 1411 1342 1415 1346
rect 1419 1342 1455 1346
rect 1459 1342 1495 1346
rect 1499 1342 1503 1346
rect 1507 1342 1535 1346
rect 1539 1342 1583 1346
rect 1587 1342 1599 1346
rect 1603 1342 1647 1346
rect 1651 1342 1679 1346
rect 1683 1342 1719 1346
rect 1723 1342 1759 1346
rect 1763 1342 1807 1346
rect 1811 1342 1831 1346
rect 1835 1342 1895 1346
rect 1899 1342 1959 1346
rect 1963 1342 1991 1346
rect 1995 1342 2023 1346
rect 2027 1342 2071 1346
rect 2075 1342 2119 1346
rect 2123 1342 2155 1346
rect 1125 1341 2155 1342
rect 2161 1341 2162 1347
rect 84 1325 85 1331
rect 91 1330 1107 1331
rect 91 1326 111 1330
rect 115 1326 135 1330
rect 139 1326 175 1330
rect 179 1326 215 1330
rect 219 1326 239 1330
rect 243 1326 255 1330
rect 259 1326 303 1330
rect 307 1326 319 1330
rect 323 1326 367 1330
rect 371 1326 391 1330
rect 395 1326 439 1330
rect 443 1326 463 1330
rect 467 1326 503 1330
rect 507 1326 543 1330
rect 547 1326 575 1330
rect 579 1326 623 1330
rect 627 1326 647 1330
rect 651 1326 703 1330
rect 707 1326 711 1330
rect 715 1326 783 1330
rect 787 1326 855 1330
rect 859 1326 863 1330
rect 867 1326 927 1330
rect 931 1326 943 1330
rect 947 1326 999 1330
rect 1003 1326 1023 1330
rect 1027 1326 1047 1330
rect 1051 1326 1095 1330
rect 1099 1326 1107 1330
rect 91 1325 1107 1326
rect 1113 1325 1114 1331
rect 1106 1289 1107 1295
rect 1113 1294 2143 1295
rect 1113 1290 1135 1294
rect 1139 1290 1159 1294
rect 1163 1290 1175 1294
rect 1179 1290 1223 1294
rect 1227 1290 1231 1294
rect 1235 1290 1303 1294
rect 1307 1290 1311 1294
rect 1315 1290 1391 1294
rect 1395 1290 1407 1294
rect 1411 1290 1479 1294
rect 1483 1290 1503 1294
rect 1507 1290 1567 1294
rect 1571 1290 1599 1294
rect 1603 1290 1655 1294
rect 1659 1290 1679 1294
rect 1683 1290 1743 1294
rect 1747 1290 1759 1294
rect 1763 1290 1831 1294
rect 1835 1290 1895 1294
rect 1899 1290 1919 1294
rect 1923 1290 1959 1294
rect 1963 1290 2007 1294
rect 2011 1290 2023 1294
rect 2027 1290 2071 1294
rect 2075 1290 2119 1294
rect 2123 1290 2143 1294
rect 1113 1289 2143 1290
rect 2149 1289 2150 1295
rect 96 1269 97 1275
rect 103 1274 1119 1275
rect 103 1270 111 1274
rect 115 1270 135 1274
rect 139 1270 175 1274
rect 179 1270 215 1274
rect 219 1270 255 1274
rect 259 1270 319 1274
rect 323 1270 391 1274
rect 395 1270 399 1274
rect 403 1270 463 1274
rect 467 1270 487 1274
rect 491 1270 543 1274
rect 547 1270 583 1274
rect 587 1270 623 1274
rect 627 1270 687 1274
rect 691 1270 703 1274
rect 707 1270 783 1274
rect 787 1270 799 1274
rect 803 1270 863 1274
rect 867 1270 919 1274
rect 923 1270 943 1274
rect 947 1270 1023 1274
rect 1027 1270 1047 1274
rect 1051 1270 1095 1274
rect 1099 1270 1119 1274
rect 103 1269 1119 1270
rect 1125 1269 1126 1275
rect 1118 1233 1119 1239
rect 1125 1238 2155 1239
rect 1125 1234 1135 1238
rect 1139 1234 1175 1238
rect 1179 1234 1231 1238
rect 1235 1234 1287 1238
rect 1291 1234 1303 1238
rect 1307 1234 1327 1238
rect 1331 1234 1375 1238
rect 1379 1234 1391 1238
rect 1395 1234 1431 1238
rect 1435 1234 1479 1238
rect 1483 1234 1495 1238
rect 1499 1234 1559 1238
rect 1563 1234 1567 1238
rect 1571 1234 1623 1238
rect 1627 1234 1655 1238
rect 1659 1234 1679 1238
rect 1683 1234 1735 1238
rect 1739 1234 1743 1238
rect 1747 1234 1791 1238
rect 1795 1234 1831 1238
rect 1835 1234 1847 1238
rect 1851 1234 1903 1238
rect 1907 1234 1919 1238
rect 1923 1234 1967 1238
rect 1971 1234 2007 1238
rect 2011 1234 2031 1238
rect 2035 1234 2071 1238
rect 2075 1234 2119 1238
rect 2123 1234 2155 1238
rect 1125 1233 2155 1234
rect 2161 1233 2162 1239
rect 84 1213 85 1219
rect 91 1218 1107 1219
rect 91 1214 111 1218
rect 115 1214 135 1218
rect 139 1214 175 1218
rect 179 1214 215 1218
rect 219 1214 255 1218
rect 259 1214 271 1218
rect 275 1214 311 1218
rect 315 1214 319 1218
rect 323 1214 351 1218
rect 355 1214 399 1218
rect 403 1214 447 1218
rect 451 1214 487 1218
rect 491 1214 495 1218
rect 499 1214 551 1218
rect 555 1214 583 1218
rect 587 1214 607 1218
rect 611 1214 671 1218
rect 675 1214 687 1218
rect 691 1214 743 1218
rect 747 1214 799 1218
rect 803 1214 815 1218
rect 819 1214 895 1218
rect 899 1214 919 1218
rect 923 1214 983 1218
rect 987 1214 1047 1218
rect 1051 1214 1095 1218
rect 1099 1214 1107 1218
rect 91 1213 1107 1214
rect 1113 1213 1114 1219
rect 1106 1181 1107 1187
rect 1113 1186 2143 1187
rect 1113 1182 1135 1186
rect 1139 1182 1159 1186
rect 1163 1182 1207 1186
rect 1211 1182 1279 1186
rect 1283 1182 1287 1186
rect 1291 1182 1327 1186
rect 1331 1182 1351 1186
rect 1355 1182 1375 1186
rect 1379 1182 1423 1186
rect 1427 1182 1431 1186
rect 1435 1182 1487 1186
rect 1491 1182 1495 1186
rect 1499 1182 1559 1186
rect 1563 1182 1623 1186
rect 1627 1182 1631 1186
rect 1635 1182 1679 1186
rect 1683 1182 1711 1186
rect 1715 1182 1735 1186
rect 1739 1182 1791 1186
rect 1795 1182 1799 1186
rect 1803 1182 1847 1186
rect 1851 1182 1887 1186
rect 1891 1182 1903 1186
rect 1907 1182 1967 1186
rect 1971 1182 1983 1186
rect 1987 1182 2031 1186
rect 2035 1182 2071 1186
rect 2075 1182 2119 1186
rect 2123 1182 2143 1186
rect 1113 1181 2143 1182
rect 2149 1181 2150 1187
rect 96 1157 97 1163
rect 103 1162 1119 1163
rect 103 1158 111 1162
rect 115 1158 271 1162
rect 275 1158 311 1162
rect 315 1158 351 1162
rect 355 1158 399 1162
rect 403 1158 439 1162
rect 443 1158 447 1162
rect 451 1158 479 1162
rect 483 1158 495 1162
rect 499 1158 527 1162
rect 531 1158 551 1162
rect 555 1158 575 1162
rect 579 1158 607 1162
rect 611 1158 623 1162
rect 627 1158 671 1162
rect 675 1158 719 1162
rect 723 1158 743 1162
rect 747 1158 775 1162
rect 779 1158 815 1162
rect 819 1158 831 1162
rect 835 1158 887 1162
rect 891 1158 895 1162
rect 899 1158 943 1162
rect 947 1158 983 1162
rect 987 1158 1007 1162
rect 1011 1158 1047 1162
rect 1051 1158 1095 1162
rect 1099 1158 1119 1162
rect 103 1157 1119 1158
rect 1125 1157 1126 1163
rect 1118 1125 1119 1131
rect 1125 1130 2155 1131
rect 1125 1126 1135 1130
rect 1139 1126 1159 1130
rect 1163 1126 1191 1130
rect 1195 1126 1207 1130
rect 1211 1126 1271 1130
rect 1275 1126 1279 1130
rect 1283 1126 1343 1130
rect 1347 1126 1351 1130
rect 1355 1126 1415 1130
rect 1419 1126 1423 1130
rect 1427 1126 1487 1130
rect 1491 1126 1559 1130
rect 1563 1126 1567 1130
rect 1571 1126 1631 1130
rect 1635 1126 1655 1130
rect 1659 1126 1711 1130
rect 1715 1126 1751 1130
rect 1755 1126 1799 1130
rect 1803 1126 1855 1130
rect 1859 1126 1887 1130
rect 1891 1126 1959 1130
rect 1963 1126 1983 1130
rect 1987 1126 2071 1130
rect 2075 1126 2119 1130
rect 2123 1126 2155 1130
rect 1125 1125 2155 1126
rect 2161 1125 2162 1131
rect 84 1105 85 1111
rect 91 1110 1107 1111
rect 91 1106 111 1110
rect 115 1106 159 1110
rect 163 1106 199 1110
rect 203 1106 255 1110
rect 259 1106 319 1110
rect 323 1106 399 1110
rect 403 1106 439 1110
rect 443 1106 479 1110
rect 483 1106 527 1110
rect 531 1106 559 1110
rect 563 1106 575 1110
rect 579 1106 623 1110
rect 627 1106 639 1110
rect 643 1106 671 1110
rect 675 1106 711 1110
rect 715 1106 719 1110
rect 723 1106 775 1110
rect 779 1106 783 1110
rect 787 1106 831 1110
rect 835 1106 855 1110
rect 859 1106 887 1110
rect 891 1106 927 1110
rect 931 1106 943 1110
rect 947 1106 999 1110
rect 1003 1106 1007 1110
rect 1011 1106 1047 1110
rect 1051 1106 1095 1110
rect 1099 1106 1107 1110
rect 91 1105 1107 1106
rect 1113 1105 1114 1111
rect 1106 1073 1107 1079
rect 1113 1078 2143 1079
rect 1113 1074 1135 1078
rect 1139 1074 1159 1078
rect 1163 1074 1191 1078
rect 1195 1074 1199 1078
rect 1203 1074 1247 1078
rect 1251 1074 1271 1078
rect 1275 1074 1303 1078
rect 1307 1074 1343 1078
rect 1347 1074 1351 1078
rect 1355 1074 1399 1078
rect 1403 1074 1415 1078
rect 1419 1074 1455 1078
rect 1459 1074 1487 1078
rect 1491 1074 1511 1078
rect 1515 1074 1567 1078
rect 1571 1074 1583 1078
rect 1587 1074 1655 1078
rect 1659 1074 1663 1078
rect 1667 1074 1751 1078
rect 1755 1074 1759 1078
rect 1763 1074 1855 1078
rect 1859 1074 1863 1078
rect 1867 1074 1959 1078
rect 1963 1074 1967 1078
rect 1971 1074 2071 1078
rect 2075 1074 2119 1078
rect 2123 1074 2143 1078
rect 1113 1073 2143 1074
rect 2149 1073 2150 1079
rect 96 1049 97 1055
rect 103 1054 1119 1055
rect 103 1050 111 1054
rect 115 1050 135 1054
rect 139 1050 159 1054
rect 163 1050 175 1054
rect 179 1050 199 1054
rect 203 1050 215 1054
rect 219 1050 255 1054
rect 259 1050 319 1054
rect 323 1050 383 1054
rect 387 1050 399 1054
rect 403 1050 447 1054
rect 451 1050 479 1054
rect 483 1050 511 1054
rect 515 1050 559 1054
rect 563 1050 575 1054
rect 579 1050 631 1054
rect 635 1050 639 1054
rect 643 1050 687 1054
rect 691 1050 711 1054
rect 715 1050 743 1054
rect 747 1050 783 1054
rect 787 1050 799 1054
rect 803 1050 855 1054
rect 859 1050 863 1054
rect 867 1050 927 1054
rect 931 1050 999 1054
rect 1003 1050 1047 1054
rect 1051 1050 1095 1054
rect 1099 1050 1119 1054
rect 103 1049 1119 1050
rect 1125 1049 1126 1055
rect 1118 1017 1119 1023
rect 1125 1022 2155 1023
rect 1125 1018 1135 1022
rect 1139 1018 1159 1022
rect 1163 1018 1199 1022
rect 1203 1018 1239 1022
rect 1243 1018 1247 1022
rect 1251 1018 1295 1022
rect 1299 1018 1303 1022
rect 1307 1018 1351 1022
rect 1355 1018 1399 1022
rect 1403 1018 1407 1022
rect 1411 1018 1455 1022
rect 1459 1018 1463 1022
rect 1467 1018 1511 1022
rect 1515 1018 1519 1022
rect 1523 1018 1575 1022
rect 1579 1018 1583 1022
rect 1587 1018 1639 1022
rect 1643 1018 1663 1022
rect 1667 1018 1711 1022
rect 1715 1018 1759 1022
rect 1763 1018 1791 1022
rect 1795 1018 1863 1022
rect 1867 1018 1879 1022
rect 1883 1018 1967 1022
rect 1971 1018 2063 1022
rect 2067 1018 2071 1022
rect 2075 1018 2119 1022
rect 2123 1018 2155 1022
rect 1125 1017 2155 1018
rect 2161 1017 2162 1023
rect 84 993 85 999
rect 91 998 1107 999
rect 91 994 111 998
rect 115 994 135 998
rect 139 994 175 998
rect 179 994 215 998
rect 219 994 223 998
rect 227 994 255 998
rect 259 994 279 998
rect 283 994 319 998
rect 323 994 343 998
rect 347 994 383 998
rect 387 994 407 998
rect 411 994 447 998
rect 451 994 471 998
rect 475 994 511 998
rect 515 994 527 998
rect 531 994 575 998
rect 579 994 583 998
rect 587 994 631 998
rect 635 994 687 998
rect 691 994 743 998
rect 747 994 799 998
rect 803 994 863 998
rect 867 994 1095 998
rect 1099 994 1107 998
rect 91 993 1107 994
rect 1113 993 1114 999
rect 1106 957 1107 963
rect 1113 962 2143 963
rect 1113 958 1135 962
rect 1139 958 1159 962
rect 1163 958 1199 962
rect 1203 958 1207 962
rect 1211 958 1239 962
rect 1243 958 1287 962
rect 1291 958 1295 962
rect 1299 958 1351 962
rect 1355 958 1375 962
rect 1379 958 1407 962
rect 1411 958 1455 962
rect 1459 958 1463 962
rect 1467 958 1519 962
rect 1523 958 1535 962
rect 1539 958 1575 962
rect 1579 958 1615 962
rect 1619 958 1639 962
rect 1643 958 1687 962
rect 1691 958 1711 962
rect 1715 958 1751 962
rect 1755 958 1791 962
rect 1795 958 1815 962
rect 1819 958 1879 962
rect 1883 958 1951 962
rect 1955 958 1967 962
rect 1971 958 2023 962
rect 2027 958 2063 962
rect 2067 958 2071 962
rect 2075 958 2119 962
rect 2123 958 2143 962
rect 1113 957 2143 958
rect 2149 957 2150 963
rect 96 937 97 943
rect 103 942 1119 943
rect 103 938 111 942
rect 115 938 135 942
rect 139 938 175 942
rect 179 938 223 942
rect 227 938 263 942
rect 267 938 279 942
rect 283 938 303 942
rect 307 938 343 942
rect 347 938 351 942
rect 355 938 399 942
rect 403 938 407 942
rect 411 938 455 942
rect 459 938 471 942
rect 475 938 511 942
rect 515 938 527 942
rect 531 938 567 942
rect 571 938 583 942
rect 587 938 623 942
rect 627 938 631 942
rect 635 938 687 942
rect 691 938 743 942
rect 747 938 751 942
rect 755 938 799 942
rect 803 938 815 942
rect 819 938 879 942
rect 883 938 943 942
rect 947 938 1007 942
rect 1011 938 1047 942
rect 1051 938 1095 942
rect 1099 938 1119 942
rect 103 937 1119 938
rect 1125 937 1126 943
rect 1118 905 1119 911
rect 1125 910 2155 911
rect 1125 906 1135 910
rect 1139 906 1159 910
rect 1163 906 1207 910
rect 1211 906 1239 910
rect 1243 906 1287 910
rect 1291 906 1319 910
rect 1323 906 1375 910
rect 1379 906 1407 910
rect 1411 906 1455 910
rect 1459 906 1495 910
rect 1499 906 1535 910
rect 1539 906 1583 910
rect 1587 906 1615 910
rect 1619 906 1663 910
rect 1667 906 1687 910
rect 1691 906 1743 910
rect 1747 906 1751 910
rect 1755 906 1815 910
rect 1819 906 1879 910
rect 1883 906 1887 910
rect 1891 906 1951 910
rect 1955 906 2023 910
rect 2027 906 2071 910
rect 2075 906 2119 910
rect 2123 906 2155 910
rect 1125 905 2155 906
rect 2161 905 2162 911
rect 84 881 85 887
rect 91 886 1107 887
rect 91 882 111 886
rect 115 882 263 886
rect 267 882 303 886
rect 307 882 351 886
rect 355 882 399 886
rect 403 882 415 886
rect 419 882 455 886
rect 459 882 479 886
rect 483 882 511 886
rect 515 882 551 886
rect 555 882 567 886
rect 571 882 623 886
rect 627 882 687 886
rect 691 882 695 886
rect 699 882 751 886
rect 755 882 767 886
rect 771 882 815 886
rect 819 882 831 886
rect 835 882 879 886
rect 883 882 887 886
rect 891 882 943 886
rect 947 882 1007 886
rect 1011 882 1047 886
rect 1051 882 1095 886
rect 1099 882 1107 886
rect 91 881 1107 882
rect 1113 881 1114 887
rect 1106 853 1107 859
rect 1113 858 2143 859
rect 1113 854 1135 858
rect 1139 854 1159 858
rect 1163 854 1239 858
rect 1243 854 1247 858
rect 1251 854 1319 858
rect 1323 854 1359 858
rect 1363 854 1407 858
rect 1411 854 1455 858
rect 1459 854 1495 858
rect 1499 854 1543 858
rect 1547 854 1583 858
rect 1587 854 1631 858
rect 1635 854 1663 858
rect 1667 854 1711 858
rect 1715 854 1743 858
rect 1747 854 1783 858
rect 1787 854 1815 858
rect 1819 854 1855 858
rect 1859 854 1887 858
rect 1891 854 1935 858
rect 1939 854 1951 858
rect 1955 854 2015 858
rect 2019 854 2023 858
rect 2027 854 2071 858
rect 2075 854 2119 858
rect 2123 854 2143 858
rect 1113 853 2143 854
rect 2149 853 2150 859
rect 96 829 97 835
rect 103 834 1119 835
rect 103 830 111 834
rect 115 830 279 834
rect 283 830 303 834
rect 307 830 343 834
rect 347 830 351 834
rect 355 830 415 834
rect 419 830 479 834
rect 483 830 487 834
rect 491 830 551 834
rect 555 830 567 834
rect 571 830 623 834
rect 627 830 647 834
rect 651 830 695 834
rect 699 830 727 834
rect 731 830 767 834
rect 771 830 799 834
rect 803 830 831 834
rect 835 830 863 834
rect 867 830 887 834
rect 891 830 927 834
rect 931 830 943 834
rect 947 830 999 834
rect 1003 830 1007 834
rect 1011 830 1047 834
rect 1051 830 1095 834
rect 1099 830 1119 834
rect 103 829 1119 830
rect 1125 829 1126 835
rect 1118 801 1119 807
rect 1125 806 2155 807
rect 1125 802 1135 806
rect 1139 802 1159 806
rect 1163 802 1247 806
rect 1251 802 1279 806
rect 1283 802 1359 806
rect 1363 802 1407 806
rect 1411 802 1455 806
rect 1459 802 1519 806
rect 1523 802 1543 806
rect 1547 802 1623 806
rect 1627 802 1631 806
rect 1635 802 1711 806
rect 1715 802 1719 806
rect 1723 802 1783 806
rect 1787 802 1815 806
rect 1819 802 1855 806
rect 1859 802 1903 806
rect 1907 802 1935 806
rect 1939 802 1999 806
rect 2003 802 2015 806
rect 2019 802 2071 806
rect 2075 802 2119 806
rect 2123 802 2155 806
rect 1125 801 2155 802
rect 2161 801 2162 807
rect 84 777 85 783
rect 91 782 1107 783
rect 91 778 111 782
rect 115 778 215 782
rect 219 778 279 782
rect 283 778 343 782
rect 347 778 351 782
rect 355 778 415 782
rect 419 778 423 782
rect 427 778 487 782
rect 491 778 495 782
rect 499 778 567 782
rect 571 778 639 782
rect 643 778 647 782
rect 651 778 703 782
rect 707 778 727 782
rect 731 778 759 782
rect 763 778 799 782
rect 803 778 815 782
rect 819 778 863 782
rect 867 778 911 782
rect 915 778 927 782
rect 931 778 959 782
rect 963 778 999 782
rect 1003 778 1007 782
rect 1011 778 1047 782
rect 1051 778 1095 782
rect 1099 778 1107 782
rect 91 777 1107 778
rect 1113 777 1114 783
rect 1106 745 1107 751
rect 1113 750 2143 751
rect 1113 746 1135 750
rect 1139 746 1159 750
rect 1163 746 1279 750
rect 1283 746 1335 750
rect 1339 746 1375 750
rect 1379 746 1407 750
rect 1411 746 1415 750
rect 1419 746 1455 750
rect 1459 746 1503 750
rect 1507 746 1519 750
rect 1523 746 1551 750
rect 1555 746 1599 750
rect 1603 746 1623 750
rect 1627 746 1655 750
rect 1659 746 1711 750
rect 1715 746 1719 750
rect 1723 746 1767 750
rect 1771 746 1815 750
rect 1819 746 1831 750
rect 1835 746 1895 750
rect 1899 746 1903 750
rect 1907 746 1959 750
rect 1963 746 1999 750
rect 2003 746 2023 750
rect 2027 746 2071 750
rect 2075 746 2119 750
rect 2123 746 2143 750
rect 1113 745 2143 746
rect 2149 745 2150 751
rect 96 725 97 731
rect 103 730 1119 731
rect 103 726 111 730
rect 115 726 175 730
rect 179 726 215 730
rect 219 726 239 730
rect 243 726 279 730
rect 283 726 311 730
rect 315 726 351 730
rect 355 726 391 730
rect 395 726 423 730
rect 427 726 471 730
rect 475 726 495 730
rect 499 726 543 730
rect 547 726 567 730
rect 571 726 615 730
rect 619 726 639 730
rect 643 726 679 730
rect 683 726 703 730
rect 707 726 735 730
rect 739 726 759 730
rect 763 726 799 730
rect 803 726 815 730
rect 819 726 863 730
rect 867 726 911 730
rect 915 726 927 730
rect 931 726 959 730
rect 963 726 1007 730
rect 1011 726 1047 730
rect 1051 726 1095 730
rect 1099 726 1119 730
rect 103 725 1119 726
rect 1125 725 1126 731
rect 1118 693 1119 699
rect 1125 698 2155 699
rect 1125 694 1135 698
rect 1139 694 1247 698
rect 1251 694 1287 698
rect 1291 694 1335 698
rect 1339 694 1375 698
rect 1379 694 1391 698
rect 1395 694 1415 698
rect 1419 694 1447 698
rect 1451 694 1455 698
rect 1459 694 1503 698
rect 1507 694 1511 698
rect 1515 694 1551 698
rect 1555 694 1583 698
rect 1587 694 1599 698
rect 1603 694 1655 698
rect 1659 694 1711 698
rect 1715 694 1735 698
rect 1739 694 1767 698
rect 1771 694 1823 698
rect 1827 694 1831 698
rect 1835 694 1895 698
rect 1899 694 1911 698
rect 1915 694 1959 698
rect 1963 694 1999 698
rect 2003 694 2023 698
rect 2027 694 2071 698
rect 2075 694 2119 698
rect 2123 694 2155 698
rect 1125 693 2155 694
rect 2161 693 2162 699
rect 84 673 85 679
rect 91 678 1107 679
rect 91 674 111 678
rect 115 674 135 678
rect 139 674 175 678
rect 179 674 215 678
rect 219 674 239 678
rect 243 674 271 678
rect 275 674 311 678
rect 315 674 335 678
rect 339 674 391 678
rect 395 674 399 678
rect 403 674 463 678
rect 467 674 471 678
rect 475 674 527 678
rect 531 674 543 678
rect 547 674 591 678
rect 595 674 615 678
rect 619 674 647 678
rect 651 674 679 678
rect 683 674 703 678
rect 707 674 735 678
rect 739 674 759 678
rect 763 674 799 678
rect 803 674 823 678
rect 827 674 863 678
rect 867 674 927 678
rect 931 674 1095 678
rect 1099 674 1107 678
rect 91 673 1107 674
rect 1113 673 1114 679
rect 1106 641 1107 647
rect 1113 646 2143 647
rect 1113 642 1135 646
rect 1139 642 1159 646
rect 1163 642 1199 646
rect 1203 642 1239 646
rect 1243 642 1247 646
rect 1251 642 1279 646
rect 1283 642 1287 646
rect 1291 642 1335 646
rect 1339 642 1343 646
rect 1347 642 1391 646
rect 1395 642 1415 646
rect 1419 642 1447 646
rect 1451 642 1495 646
rect 1499 642 1511 646
rect 1515 642 1583 646
rect 1587 642 1655 646
rect 1659 642 1671 646
rect 1675 642 1735 646
rect 1739 642 1759 646
rect 1763 642 1823 646
rect 1827 642 1839 646
rect 1843 642 1911 646
rect 1915 642 1919 646
rect 1923 642 1999 646
rect 2003 642 2007 646
rect 2011 642 2071 646
rect 2075 642 2119 646
rect 2123 642 2143 646
rect 1113 641 2143 642
rect 2149 641 2150 647
rect 96 613 97 619
rect 103 618 1119 619
rect 103 614 111 618
rect 115 614 135 618
rect 139 614 175 618
rect 179 614 215 618
rect 219 614 255 618
rect 259 614 271 618
rect 275 614 303 618
rect 307 614 335 618
rect 339 614 351 618
rect 355 614 399 618
rect 403 614 439 618
rect 443 614 463 618
rect 467 614 487 618
rect 491 614 527 618
rect 531 614 535 618
rect 539 614 583 618
rect 587 614 591 618
rect 595 614 631 618
rect 635 614 647 618
rect 651 614 679 618
rect 683 614 703 618
rect 707 614 727 618
rect 731 614 759 618
rect 763 614 823 618
rect 827 614 1095 618
rect 1099 614 1119 618
rect 103 613 1119 614
rect 1125 613 1126 619
rect 1118 585 1119 591
rect 1125 590 2155 591
rect 1125 586 1135 590
rect 1139 586 1159 590
rect 1163 586 1199 590
rect 1203 586 1239 590
rect 1243 586 1279 590
rect 1283 586 1319 590
rect 1323 586 1343 590
rect 1347 586 1359 590
rect 1363 586 1415 590
rect 1419 586 1487 590
rect 1491 586 1495 590
rect 1499 586 1567 590
rect 1571 586 1583 590
rect 1587 586 1655 590
rect 1659 586 1671 590
rect 1675 586 1751 590
rect 1755 586 1759 590
rect 1763 586 1839 590
rect 1843 586 1855 590
rect 1859 586 1919 590
rect 1923 586 1967 590
rect 1971 586 2007 590
rect 2011 586 2071 590
rect 2075 586 2119 590
rect 2123 586 2155 590
rect 1125 585 2155 586
rect 2161 585 2162 591
rect 84 557 85 563
rect 91 562 1107 563
rect 91 558 111 562
rect 115 558 135 562
rect 139 558 175 562
rect 179 558 215 562
rect 219 558 223 562
rect 227 558 255 562
rect 259 558 279 562
rect 283 558 303 562
rect 307 558 327 562
rect 331 558 351 562
rect 355 558 375 562
rect 379 558 399 562
rect 403 558 423 562
rect 427 558 439 562
rect 443 558 463 562
rect 467 558 487 562
rect 491 558 511 562
rect 515 558 535 562
rect 539 558 559 562
rect 563 558 583 562
rect 587 558 607 562
rect 611 558 631 562
rect 635 558 655 562
rect 659 558 679 562
rect 683 558 703 562
rect 707 558 727 562
rect 731 558 751 562
rect 755 558 1095 562
rect 1099 558 1107 562
rect 91 557 1107 558
rect 1113 557 1114 563
rect 1106 529 1107 535
rect 1113 534 2143 535
rect 1113 530 1135 534
rect 1139 530 1159 534
rect 1163 530 1199 534
rect 1203 530 1239 534
rect 1243 530 1279 534
rect 1283 530 1303 534
rect 1307 530 1319 534
rect 1323 530 1343 534
rect 1347 530 1359 534
rect 1363 530 1383 534
rect 1387 530 1415 534
rect 1419 530 1423 534
rect 1427 530 1463 534
rect 1467 530 1487 534
rect 1491 530 1503 534
rect 1507 530 1543 534
rect 1547 530 1567 534
rect 1571 530 1591 534
rect 1595 530 1647 534
rect 1651 530 1655 534
rect 1659 530 1703 534
rect 1707 530 1751 534
rect 1755 530 1767 534
rect 1771 530 1839 534
rect 1843 530 1855 534
rect 1859 530 1919 534
rect 1923 530 1967 534
rect 1971 530 2007 534
rect 2011 530 2071 534
rect 2075 530 2119 534
rect 2123 530 2143 534
rect 1113 529 2143 530
rect 2149 529 2150 535
rect 96 497 97 503
rect 103 502 1119 503
rect 103 498 111 502
rect 115 498 135 502
rect 139 498 175 502
rect 179 498 223 502
rect 227 498 231 502
rect 235 498 279 502
rect 283 498 295 502
rect 299 498 327 502
rect 331 498 359 502
rect 363 498 375 502
rect 379 498 423 502
rect 427 498 463 502
rect 467 498 479 502
rect 483 498 511 502
rect 515 498 535 502
rect 539 498 559 502
rect 563 498 591 502
rect 595 498 607 502
rect 611 498 639 502
rect 643 498 655 502
rect 659 498 687 502
rect 691 498 703 502
rect 707 498 735 502
rect 739 498 751 502
rect 755 498 791 502
rect 795 498 847 502
rect 851 498 1095 502
rect 1099 498 1119 502
rect 103 497 1119 498
rect 1125 497 1126 503
rect 1118 477 1119 483
rect 1125 482 2155 483
rect 1125 478 1135 482
rect 1139 478 1295 482
rect 1299 478 1303 482
rect 1307 478 1335 482
rect 1339 478 1343 482
rect 1347 478 1375 482
rect 1379 478 1383 482
rect 1387 478 1423 482
rect 1427 478 1463 482
rect 1467 478 1471 482
rect 1475 478 1503 482
rect 1507 478 1527 482
rect 1531 478 1543 482
rect 1547 478 1583 482
rect 1587 478 1591 482
rect 1595 478 1647 482
rect 1651 478 1703 482
rect 1707 478 1719 482
rect 1723 478 1767 482
rect 1771 478 1807 482
rect 1811 478 1839 482
rect 1843 478 1895 482
rect 1899 478 1919 482
rect 1923 478 1991 482
rect 1995 478 2007 482
rect 2011 478 2071 482
rect 2075 478 2119 482
rect 2123 478 2155 482
rect 1125 477 2155 478
rect 2161 477 2162 483
rect 84 441 85 447
rect 91 446 1107 447
rect 91 442 111 446
rect 115 442 135 446
rect 139 442 175 446
rect 179 442 215 446
rect 219 442 231 446
rect 235 442 263 446
rect 267 442 295 446
rect 299 442 327 446
rect 331 442 359 446
rect 363 442 391 446
rect 395 442 423 446
rect 427 442 463 446
rect 467 442 479 446
rect 483 442 535 446
rect 539 442 591 446
rect 595 442 607 446
rect 611 442 639 446
rect 643 442 679 446
rect 683 442 687 446
rect 691 442 735 446
rect 739 442 743 446
rect 747 442 791 446
rect 795 442 807 446
rect 811 442 847 446
rect 851 442 871 446
rect 875 442 943 446
rect 947 442 1095 446
rect 1099 442 1107 446
rect 91 441 1107 442
rect 1113 441 1114 447
rect 1106 425 1107 431
rect 1113 430 2143 431
rect 1113 426 1135 430
rect 1139 426 1159 430
rect 1163 426 1199 430
rect 1203 426 1255 430
rect 1259 426 1295 430
rect 1299 426 1335 430
rect 1339 426 1375 430
rect 1379 426 1415 430
rect 1419 426 1423 430
rect 1427 426 1471 430
rect 1475 426 1503 430
rect 1507 426 1527 430
rect 1531 426 1583 430
rect 1587 426 1591 430
rect 1595 426 1647 430
rect 1651 426 1671 430
rect 1675 426 1719 430
rect 1723 426 1751 430
rect 1755 426 1807 430
rect 1811 426 1831 430
rect 1835 426 1895 430
rect 1899 426 1911 430
rect 1915 426 1991 430
rect 1995 426 1999 430
rect 2003 426 2071 430
rect 2075 426 2119 430
rect 2123 426 2143 430
rect 1113 425 2143 426
rect 2149 425 2150 431
rect 96 381 97 387
rect 103 386 1119 387
rect 103 382 111 386
rect 115 382 175 386
rect 179 382 215 386
rect 219 382 263 386
rect 267 382 271 386
rect 275 382 327 386
rect 331 382 335 386
rect 339 382 391 386
rect 395 382 407 386
rect 411 382 463 386
rect 467 382 487 386
rect 491 382 535 386
rect 539 382 567 386
rect 571 382 607 386
rect 611 382 639 386
rect 643 382 679 386
rect 683 382 711 386
rect 715 382 743 386
rect 747 382 775 386
rect 779 382 807 386
rect 811 382 839 386
rect 843 382 871 386
rect 875 382 895 386
rect 899 382 943 386
rect 947 382 951 386
rect 955 382 1007 386
rect 1011 382 1047 386
rect 1051 382 1095 386
rect 1099 382 1119 386
rect 103 381 1119 382
rect 1125 381 1126 387
rect 1118 369 1119 375
rect 1125 374 2155 375
rect 1125 370 1135 374
rect 1139 370 1159 374
rect 1163 370 1199 374
rect 1203 370 1247 374
rect 1251 370 1255 374
rect 1259 370 1335 374
rect 1339 370 1359 374
rect 1363 370 1415 374
rect 1419 370 1463 374
rect 1467 370 1503 374
rect 1507 370 1559 374
rect 1563 370 1591 374
rect 1595 370 1647 374
rect 1651 370 1671 374
rect 1675 370 1727 374
rect 1731 370 1751 374
rect 1755 370 1799 374
rect 1803 370 1831 374
rect 1835 370 1863 374
rect 1867 370 1911 374
rect 1915 370 1919 374
rect 1923 370 1975 374
rect 1979 370 1999 374
rect 2003 370 2031 374
rect 2035 370 2071 374
rect 2075 370 2119 374
rect 2123 370 2155 374
rect 1125 369 2155 370
rect 2161 369 2162 375
rect 84 325 85 331
rect 91 330 1107 331
rect 91 326 111 330
rect 115 326 175 330
rect 179 326 215 330
rect 219 326 271 330
rect 275 326 335 330
rect 339 326 383 330
rect 387 326 407 330
rect 411 326 423 330
rect 427 326 463 330
rect 467 326 487 330
rect 491 326 503 330
rect 507 326 543 330
rect 547 326 567 330
rect 571 326 591 330
rect 595 326 639 330
rect 643 326 687 330
rect 691 326 711 330
rect 715 326 735 330
rect 739 326 775 330
rect 779 326 783 330
rect 787 326 831 330
rect 835 326 839 330
rect 843 326 879 330
rect 883 326 895 330
rect 899 326 927 330
rect 931 326 951 330
rect 955 326 967 330
rect 971 326 1007 330
rect 1011 326 1047 330
rect 1051 326 1095 330
rect 1099 326 1107 330
rect 91 325 1107 326
rect 1113 325 1114 331
rect 1106 309 1107 315
rect 1113 314 2143 315
rect 1113 310 1135 314
rect 1139 310 1159 314
rect 1163 310 1247 314
rect 1251 310 1351 314
rect 1355 310 1359 314
rect 1363 310 1391 314
rect 1395 310 1431 314
rect 1435 310 1463 314
rect 1467 310 1471 314
rect 1475 310 1511 314
rect 1515 310 1559 314
rect 1563 310 1615 314
rect 1619 310 1647 314
rect 1651 310 1671 314
rect 1675 310 1727 314
rect 1731 310 1735 314
rect 1739 310 1799 314
rect 1803 310 1807 314
rect 1811 310 1863 314
rect 1867 310 1887 314
rect 1891 310 1919 314
rect 1923 310 1967 314
rect 1971 310 1975 314
rect 1979 310 2031 314
rect 2035 310 2047 314
rect 2051 310 2071 314
rect 2075 310 2119 314
rect 2123 310 2143 314
rect 1113 309 2143 310
rect 2149 309 2150 315
rect 96 265 97 271
rect 103 270 1119 271
rect 103 266 111 270
rect 115 266 287 270
rect 291 266 327 270
rect 331 266 367 270
rect 371 266 383 270
rect 387 266 415 270
rect 419 266 423 270
rect 427 266 463 270
rect 467 266 471 270
rect 475 266 503 270
rect 507 266 535 270
rect 539 266 543 270
rect 547 266 591 270
rect 595 266 607 270
rect 611 266 639 270
rect 643 266 679 270
rect 683 266 687 270
rect 691 266 735 270
rect 739 266 743 270
rect 747 266 783 270
rect 787 266 807 270
rect 811 266 831 270
rect 835 266 863 270
rect 867 266 879 270
rect 883 266 927 270
rect 931 266 967 270
rect 971 266 991 270
rect 995 266 1007 270
rect 1011 266 1047 270
rect 1051 266 1095 270
rect 1099 266 1119 270
rect 103 265 1119 266
rect 1125 265 1126 271
rect 1118 263 1126 265
rect 1118 257 1119 263
rect 1125 262 2155 263
rect 1125 258 1135 262
rect 1139 258 1263 262
rect 1267 258 1303 262
rect 1307 258 1343 262
rect 1347 258 1351 262
rect 1355 258 1383 262
rect 1387 258 1391 262
rect 1395 258 1423 262
rect 1427 258 1431 262
rect 1435 258 1463 262
rect 1467 258 1471 262
rect 1475 258 1503 262
rect 1507 258 1511 262
rect 1515 258 1543 262
rect 1547 258 1559 262
rect 1563 258 1599 262
rect 1603 258 1615 262
rect 1619 258 1671 262
rect 1675 258 1735 262
rect 1739 258 1759 262
rect 1763 258 1807 262
rect 1811 258 1863 262
rect 1867 258 1887 262
rect 1891 258 1967 262
rect 1971 258 1975 262
rect 1979 258 2047 262
rect 2051 258 2071 262
rect 2075 258 2119 262
rect 2123 258 2155 262
rect 1125 257 2155 258
rect 2161 257 2162 263
rect 84 201 85 207
rect 91 206 1107 207
rect 91 202 111 206
rect 115 202 167 206
rect 171 202 207 206
rect 211 202 247 206
rect 251 202 287 206
rect 291 202 295 206
rect 299 202 327 206
rect 331 202 343 206
rect 347 202 367 206
rect 371 202 399 206
rect 403 202 415 206
rect 419 202 463 206
rect 467 202 471 206
rect 475 202 527 206
rect 531 202 535 206
rect 539 202 599 206
rect 603 202 607 206
rect 611 202 671 206
rect 675 202 679 206
rect 683 202 743 206
rect 747 202 751 206
rect 755 202 807 206
rect 811 202 831 206
rect 835 202 863 206
rect 867 202 911 206
rect 915 202 927 206
rect 931 202 991 206
rect 995 202 1047 206
rect 1051 202 1095 206
rect 1099 202 1107 206
rect 91 201 1107 202
rect 1113 206 2150 207
rect 1113 202 1135 206
rect 1139 202 1183 206
rect 1187 202 1231 206
rect 1235 202 1263 206
rect 1267 202 1295 206
rect 1299 202 1303 206
rect 1307 202 1343 206
rect 1347 202 1359 206
rect 1363 202 1383 206
rect 1387 202 1423 206
rect 1427 202 1431 206
rect 1435 202 1463 206
rect 1467 202 1503 206
rect 1507 202 1511 206
rect 1515 202 1543 206
rect 1547 202 1591 206
rect 1595 202 1599 206
rect 1603 202 1663 206
rect 1667 202 1671 206
rect 1675 202 1735 206
rect 1739 202 1759 206
rect 1763 202 1807 206
rect 1811 202 1863 206
rect 1867 202 1879 206
rect 1883 202 1951 206
rect 1955 202 1975 206
rect 1979 202 2023 206
rect 2027 202 2071 206
rect 2075 202 2119 206
rect 2123 202 2150 206
rect 1113 201 2150 202
rect 96 133 97 139
rect 103 138 1119 139
rect 103 134 111 138
rect 115 134 135 138
rect 139 134 167 138
rect 171 134 175 138
rect 179 134 207 138
rect 211 134 215 138
rect 219 134 247 138
rect 251 134 255 138
rect 259 134 295 138
rect 299 134 335 138
rect 339 134 343 138
rect 347 134 375 138
rect 379 134 399 138
rect 403 134 415 138
rect 419 134 455 138
rect 459 134 463 138
rect 467 134 495 138
rect 499 134 527 138
rect 531 134 535 138
rect 539 134 575 138
rect 579 134 599 138
rect 603 134 615 138
rect 619 134 655 138
rect 659 134 671 138
rect 675 134 695 138
rect 699 134 735 138
rect 739 134 751 138
rect 755 134 775 138
rect 779 134 815 138
rect 819 134 831 138
rect 835 134 871 138
rect 875 134 911 138
rect 915 134 935 138
rect 939 134 991 138
rect 995 134 999 138
rect 1003 134 1047 138
rect 1051 134 1095 138
rect 1099 134 1119 138
rect 103 133 1119 134
rect 1125 133 1126 139
rect 1118 131 1126 133
rect 1118 125 1119 131
rect 1125 130 2155 131
rect 1125 126 1135 130
rect 1139 126 1159 130
rect 1163 126 1183 130
rect 1187 126 1199 130
rect 1203 126 1231 130
rect 1235 126 1239 130
rect 1243 126 1279 130
rect 1283 126 1295 130
rect 1299 126 1319 130
rect 1323 126 1359 130
rect 1363 126 1367 130
rect 1371 126 1431 130
rect 1435 126 1495 130
rect 1499 126 1511 130
rect 1515 126 1559 130
rect 1563 126 1591 130
rect 1595 126 1615 130
rect 1619 126 1663 130
rect 1667 126 1671 130
rect 1675 126 1719 130
rect 1723 126 1735 130
rect 1739 126 1767 130
rect 1771 126 1807 130
rect 1811 126 1855 130
rect 1859 126 1879 130
rect 1883 126 1903 130
rect 1907 126 1951 130
rect 1955 126 1991 130
rect 1995 126 2023 130
rect 2027 126 2031 130
rect 2035 126 2071 130
rect 2075 126 2119 130
rect 2123 126 2155 130
rect 1125 125 2155 126
rect 2161 125 2162 131
rect 84 81 85 87
rect 91 86 1107 87
rect 91 82 111 86
rect 115 82 135 86
rect 139 82 175 86
rect 179 82 215 86
rect 219 82 255 86
rect 259 82 295 86
rect 299 82 335 86
rect 339 82 375 86
rect 379 82 415 86
rect 419 82 455 86
rect 459 82 495 86
rect 499 82 535 86
rect 539 82 575 86
rect 579 82 615 86
rect 619 82 655 86
rect 659 82 695 86
rect 699 82 735 86
rect 739 82 775 86
rect 779 82 815 86
rect 819 82 871 86
rect 875 82 935 86
rect 939 82 999 86
rect 1003 82 1047 86
rect 1051 82 1095 86
rect 1099 82 1107 86
rect 91 81 1107 82
rect 1113 81 1114 87
rect 1106 79 1114 81
rect 1106 73 1107 79
rect 1113 78 2143 79
rect 1113 74 1135 78
rect 1139 74 1159 78
rect 1163 74 1199 78
rect 1203 74 1239 78
rect 1243 74 1279 78
rect 1283 74 1319 78
rect 1323 74 1367 78
rect 1371 74 1431 78
rect 1435 74 1495 78
rect 1499 74 1559 78
rect 1563 74 1615 78
rect 1619 74 1671 78
rect 1675 74 1719 78
rect 1723 74 1767 78
rect 1771 74 1807 78
rect 1811 74 1855 78
rect 1859 74 1903 78
rect 1907 74 1951 78
rect 1955 74 1991 78
rect 1995 74 2031 78
rect 2035 74 2071 78
rect 2075 74 2119 78
rect 2123 74 2143 78
rect 1113 73 2143 74
rect 2149 73 2150 79
<< m5c >>
rect 1119 2209 1125 2215
rect 2155 2209 2161 2215
rect 1107 2157 1113 2163
rect 2143 2157 2149 2163
rect 1119 2101 1125 2107
rect 2155 2101 2161 2107
rect 1107 2049 1113 2055
rect 2143 2049 2149 2055
rect 97 2029 103 2035
rect 1119 2029 1125 2035
rect 1119 1997 1125 2003
rect 2155 1997 2161 2003
rect 85 1977 91 1983
rect 1107 1977 1113 1983
rect 1107 1941 1113 1947
rect 2143 1941 2149 1947
rect 97 1925 103 1931
rect 1119 1925 1125 1931
rect 1119 1885 1125 1891
rect 2155 1885 2161 1891
rect 85 1869 91 1875
rect 1107 1869 1113 1875
rect 1107 1833 1113 1839
rect 2143 1833 2149 1839
rect 97 1809 103 1815
rect 1119 1809 1125 1815
rect 1119 1781 1125 1787
rect 2155 1781 2161 1787
rect 85 1757 91 1763
rect 1107 1757 1113 1763
rect 1107 1729 1113 1735
rect 2143 1729 2149 1735
rect 97 1701 103 1707
rect 1119 1701 1125 1707
rect 1119 1673 1125 1679
rect 2155 1673 2161 1679
rect 85 1645 91 1651
rect 1107 1645 1113 1651
rect 1107 1609 1113 1615
rect 2143 1609 2149 1615
rect 97 1593 103 1599
rect 1119 1593 1125 1599
rect 1119 1557 1125 1563
rect 2155 1557 2161 1563
rect 85 1541 91 1547
rect 1107 1541 1113 1547
rect 1107 1505 1113 1511
rect 2143 1505 2149 1511
rect 97 1489 103 1495
rect 1119 1489 1125 1495
rect 1119 1449 1125 1455
rect 2155 1449 2161 1455
rect 85 1437 91 1443
rect 1107 1437 1113 1443
rect 1107 1395 1113 1401
rect 2143 1393 2149 1399
rect 97 1385 103 1391
rect 1119 1385 1125 1391
rect 1119 1341 1125 1347
rect 2155 1341 2161 1347
rect 85 1325 91 1331
rect 1107 1325 1113 1331
rect 1107 1289 1113 1295
rect 2143 1289 2149 1295
rect 97 1269 103 1275
rect 1119 1269 1125 1275
rect 1119 1233 1125 1239
rect 2155 1233 2161 1239
rect 85 1213 91 1219
rect 1107 1213 1113 1219
rect 1107 1181 1113 1187
rect 2143 1181 2149 1187
rect 97 1157 103 1163
rect 1119 1157 1125 1163
rect 1119 1125 1125 1131
rect 2155 1125 2161 1131
rect 85 1105 91 1111
rect 1107 1105 1113 1111
rect 1107 1073 1113 1079
rect 2143 1073 2149 1079
rect 97 1049 103 1055
rect 1119 1049 1125 1055
rect 1119 1017 1125 1023
rect 2155 1017 2161 1023
rect 85 993 91 999
rect 1107 993 1113 999
rect 1107 957 1113 963
rect 2143 957 2149 963
rect 97 937 103 943
rect 1119 937 1125 943
rect 1119 905 1125 911
rect 2155 905 2161 911
rect 85 881 91 887
rect 1107 881 1113 887
rect 1107 853 1113 859
rect 2143 853 2149 859
rect 97 829 103 835
rect 1119 829 1125 835
rect 1119 801 1125 807
rect 2155 801 2161 807
rect 85 777 91 783
rect 1107 777 1113 783
rect 1107 745 1113 751
rect 2143 745 2149 751
rect 97 725 103 731
rect 1119 725 1125 731
rect 1119 693 1125 699
rect 2155 693 2161 699
rect 85 673 91 679
rect 1107 673 1113 679
rect 1107 641 1113 647
rect 2143 641 2149 647
rect 97 613 103 619
rect 1119 613 1125 619
rect 1119 585 1125 591
rect 2155 585 2161 591
rect 85 557 91 563
rect 1107 557 1113 563
rect 1107 529 1113 535
rect 2143 529 2149 535
rect 97 497 103 503
rect 1119 497 1125 503
rect 1119 477 1125 483
rect 2155 477 2161 483
rect 85 441 91 447
rect 1107 441 1113 447
rect 1107 425 1113 431
rect 2143 425 2149 431
rect 97 381 103 387
rect 1119 381 1125 387
rect 1119 369 1125 375
rect 2155 369 2161 375
rect 85 325 91 331
rect 1107 325 1113 331
rect 1107 309 1113 315
rect 2143 309 2149 315
rect 97 265 103 271
rect 1119 265 1125 271
rect 1119 257 1125 263
rect 2155 257 2161 263
rect 85 201 91 207
rect 1107 201 1113 207
rect 97 133 103 139
rect 1119 133 1125 139
rect 1119 125 1125 131
rect 2155 125 2161 131
rect 85 81 91 87
rect 1107 81 1113 87
rect 1107 73 1113 79
rect 2143 73 2149 79
<< m5 >>
rect 84 1983 92 2232
rect 84 1977 85 1983
rect 91 1977 92 1983
rect 84 1875 92 1977
rect 84 1869 85 1875
rect 91 1869 92 1875
rect 84 1763 92 1869
rect 84 1757 85 1763
rect 91 1757 92 1763
rect 84 1651 92 1757
rect 84 1645 85 1651
rect 91 1645 92 1651
rect 84 1547 92 1645
rect 84 1541 85 1547
rect 91 1541 92 1547
rect 84 1443 92 1541
rect 84 1437 85 1443
rect 91 1437 92 1443
rect 84 1331 92 1437
rect 84 1325 85 1331
rect 91 1325 92 1331
rect 84 1219 92 1325
rect 84 1213 85 1219
rect 91 1213 92 1219
rect 84 1111 92 1213
rect 84 1105 85 1111
rect 91 1105 92 1111
rect 84 999 92 1105
rect 84 993 85 999
rect 91 993 92 999
rect 84 887 92 993
rect 84 881 85 887
rect 91 881 92 887
rect 84 783 92 881
rect 84 777 85 783
rect 91 777 92 783
rect 84 679 92 777
rect 84 673 85 679
rect 91 673 92 679
rect 84 563 92 673
rect 84 557 85 563
rect 91 557 92 563
rect 84 447 92 557
rect 84 441 85 447
rect 91 441 92 447
rect 84 331 92 441
rect 84 325 85 331
rect 91 325 92 331
rect 84 207 92 325
rect 84 201 85 207
rect 91 201 92 207
rect 84 87 92 201
rect 84 81 85 87
rect 91 81 92 87
rect 84 72 92 81
rect 96 2035 104 2232
rect 96 2029 97 2035
rect 103 2029 104 2035
rect 96 1931 104 2029
rect 96 1925 97 1931
rect 103 1925 104 1931
rect 96 1815 104 1925
rect 96 1809 97 1815
rect 103 1809 104 1815
rect 96 1707 104 1809
rect 96 1701 97 1707
rect 103 1701 104 1707
rect 96 1599 104 1701
rect 96 1593 97 1599
rect 103 1593 104 1599
rect 96 1495 104 1593
rect 96 1489 97 1495
rect 103 1489 104 1495
rect 96 1391 104 1489
rect 96 1385 97 1391
rect 103 1385 104 1391
rect 96 1275 104 1385
rect 96 1269 97 1275
rect 103 1269 104 1275
rect 96 1163 104 1269
rect 96 1157 97 1163
rect 103 1157 104 1163
rect 96 1055 104 1157
rect 96 1049 97 1055
rect 103 1049 104 1055
rect 96 943 104 1049
rect 96 937 97 943
rect 103 937 104 943
rect 96 835 104 937
rect 96 829 97 835
rect 103 829 104 835
rect 96 731 104 829
rect 96 725 97 731
rect 103 725 104 731
rect 96 619 104 725
rect 96 613 97 619
rect 103 613 104 619
rect 96 503 104 613
rect 96 497 97 503
rect 103 497 104 503
rect 96 387 104 497
rect 96 381 97 387
rect 103 381 104 387
rect 96 271 104 381
rect 96 265 97 271
rect 103 265 104 271
rect 96 139 104 265
rect 96 133 97 139
rect 103 133 104 139
rect 96 72 104 133
rect 1106 2163 1114 2232
rect 1106 2157 1107 2163
rect 1113 2157 1114 2163
rect 1106 2055 1114 2157
rect 1106 2049 1107 2055
rect 1113 2049 1114 2055
rect 1106 1983 1114 2049
rect 1106 1977 1107 1983
rect 1113 1977 1114 1983
rect 1106 1947 1114 1977
rect 1106 1941 1107 1947
rect 1113 1941 1114 1947
rect 1106 1875 1114 1941
rect 1106 1869 1107 1875
rect 1113 1869 1114 1875
rect 1106 1839 1114 1869
rect 1106 1833 1107 1839
rect 1113 1833 1114 1839
rect 1106 1763 1114 1833
rect 1106 1757 1107 1763
rect 1113 1757 1114 1763
rect 1106 1735 1114 1757
rect 1106 1729 1107 1735
rect 1113 1729 1114 1735
rect 1106 1651 1114 1729
rect 1106 1645 1107 1651
rect 1113 1645 1114 1651
rect 1106 1615 1114 1645
rect 1106 1609 1107 1615
rect 1113 1609 1114 1615
rect 1106 1547 1114 1609
rect 1106 1541 1107 1547
rect 1113 1541 1114 1547
rect 1106 1511 1114 1541
rect 1106 1505 1107 1511
rect 1113 1505 1114 1511
rect 1106 1443 1114 1505
rect 1106 1437 1107 1443
rect 1113 1437 1114 1443
rect 1106 1401 1114 1437
rect 1106 1395 1107 1401
rect 1113 1395 1114 1401
rect 1106 1331 1114 1395
rect 1106 1325 1107 1331
rect 1113 1325 1114 1331
rect 1106 1295 1114 1325
rect 1106 1289 1107 1295
rect 1113 1289 1114 1295
rect 1106 1219 1114 1289
rect 1106 1213 1107 1219
rect 1113 1213 1114 1219
rect 1106 1187 1114 1213
rect 1106 1181 1107 1187
rect 1113 1181 1114 1187
rect 1106 1111 1114 1181
rect 1106 1105 1107 1111
rect 1113 1105 1114 1111
rect 1106 1079 1114 1105
rect 1106 1073 1107 1079
rect 1113 1073 1114 1079
rect 1106 999 1114 1073
rect 1106 993 1107 999
rect 1113 993 1114 999
rect 1106 963 1114 993
rect 1106 957 1107 963
rect 1113 957 1114 963
rect 1106 887 1114 957
rect 1106 881 1107 887
rect 1113 881 1114 887
rect 1106 859 1114 881
rect 1106 853 1107 859
rect 1113 853 1114 859
rect 1106 783 1114 853
rect 1106 777 1107 783
rect 1113 777 1114 783
rect 1106 751 1114 777
rect 1106 745 1107 751
rect 1113 745 1114 751
rect 1106 679 1114 745
rect 1106 673 1107 679
rect 1113 673 1114 679
rect 1106 647 1114 673
rect 1106 641 1107 647
rect 1113 641 1114 647
rect 1106 563 1114 641
rect 1106 557 1107 563
rect 1113 557 1114 563
rect 1106 535 1114 557
rect 1106 529 1107 535
rect 1113 529 1114 535
rect 1106 447 1114 529
rect 1106 441 1107 447
rect 1113 441 1114 447
rect 1106 431 1114 441
rect 1106 425 1107 431
rect 1113 425 1114 431
rect 1106 331 1114 425
rect 1106 325 1107 331
rect 1113 325 1114 331
rect 1106 315 1114 325
rect 1106 309 1107 315
rect 1113 309 1114 315
rect 1106 207 1114 309
rect 1106 201 1107 207
rect 1113 201 1114 207
rect 1106 87 1114 201
rect 1106 81 1107 87
rect 1113 81 1114 87
rect 1106 79 1114 81
rect 1106 73 1107 79
rect 1113 73 1114 79
rect 1106 72 1114 73
rect 1118 2215 1126 2232
rect 1118 2209 1119 2215
rect 1125 2209 1126 2215
rect 1118 2107 1126 2209
rect 1118 2101 1119 2107
rect 1125 2101 1126 2107
rect 1118 2035 1126 2101
rect 1118 2029 1119 2035
rect 1125 2029 1126 2035
rect 1118 2003 1126 2029
rect 1118 1997 1119 2003
rect 1125 1997 1126 2003
rect 1118 1931 1126 1997
rect 1118 1925 1119 1931
rect 1125 1925 1126 1931
rect 1118 1891 1126 1925
rect 1118 1885 1119 1891
rect 1125 1885 1126 1891
rect 1118 1815 1126 1885
rect 1118 1809 1119 1815
rect 1125 1809 1126 1815
rect 1118 1787 1126 1809
rect 1118 1781 1119 1787
rect 1125 1781 1126 1787
rect 1118 1707 1126 1781
rect 1118 1701 1119 1707
rect 1125 1701 1126 1707
rect 1118 1679 1126 1701
rect 1118 1673 1119 1679
rect 1125 1673 1126 1679
rect 1118 1599 1126 1673
rect 1118 1593 1119 1599
rect 1125 1593 1126 1599
rect 1118 1563 1126 1593
rect 1118 1557 1119 1563
rect 1125 1557 1126 1563
rect 1118 1495 1126 1557
rect 1118 1489 1119 1495
rect 1125 1489 1126 1495
rect 1118 1455 1126 1489
rect 1118 1449 1119 1455
rect 1125 1449 1126 1455
rect 1118 1391 1126 1449
rect 1118 1385 1119 1391
rect 1125 1385 1126 1391
rect 1118 1347 1126 1385
rect 1118 1341 1119 1347
rect 1125 1341 1126 1347
rect 1118 1275 1126 1341
rect 1118 1269 1119 1275
rect 1125 1269 1126 1275
rect 1118 1239 1126 1269
rect 1118 1233 1119 1239
rect 1125 1233 1126 1239
rect 1118 1163 1126 1233
rect 1118 1157 1119 1163
rect 1125 1157 1126 1163
rect 1118 1131 1126 1157
rect 1118 1125 1119 1131
rect 1125 1125 1126 1131
rect 1118 1055 1126 1125
rect 1118 1049 1119 1055
rect 1125 1049 1126 1055
rect 1118 1023 1126 1049
rect 1118 1017 1119 1023
rect 1125 1017 1126 1023
rect 1118 943 1126 1017
rect 1118 937 1119 943
rect 1125 937 1126 943
rect 1118 911 1126 937
rect 1118 905 1119 911
rect 1125 905 1126 911
rect 1118 835 1126 905
rect 1118 829 1119 835
rect 1125 829 1126 835
rect 1118 807 1126 829
rect 1118 801 1119 807
rect 1125 801 1126 807
rect 1118 731 1126 801
rect 1118 725 1119 731
rect 1125 725 1126 731
rect 1118 699 1126 725
rect 1118 693 1119 699
rect 1125 693 1126 699
rect 1118 619 1126 693
rect 1118 613 1119 619
rect 1125 613 1126 619
rect 1118 591 1126 613
rect 1118 585 1119 591
rect 1125 585 1126 591
rect 1118 503 1126 585
rect 1118 497 1119 503
rect 1125 497 1126 503
rect 1118 483 1126 497
rect 1118 477 1119 483
rect 1125 477 1126 483
rect 1118 387 1126 477
rect 1118 381 1119 387
rect 1125 381 1126 387
rect 1118 375 1126 381
rect 1118 369 1119 375
rect 1125 369 1126 375
rect 1118 271 1126 369
rect 1118 265 1119 271
rect 1125 265 1126 271
rect 1118 263 1126 265
rect 1118 257 1119 263
rect 1125 257 1126 263
rect 1118 139 1126 257
rect 1118 133 1119 139
rect 1125 133 1126 139
rect 1118 131 1126 133
rect 1118 125 1119 131
rect 1125 125 1126 131
rect 1118 72 1126 125
rect 2142 2163 2150 2232
rect 2142 2157 2143 2163
rect 2149 2157 2150 2163
rect 2142 2055 2150 2157
rect 2142 2049 2143 2055
rect 2149 2049 2150 2055
rect 2142 1947 2150 2049
rect 2142 1941 2143 1947
rect 2149 1941 2150 1947
rect 2142 1839 2150 1941
rect 2142 1833 2143 1839
rect 2149 1833 2150 1839
rect 2142 1735 2150 1833
rect 2142 1729 2143 1735
rect 2149 1729 2150 1735
rect 2142 1615 2150 1729
rect 2142 1609 2143 1615
rect 2149 1609 2150 1615
rect 2142 1511 2150 1609
rect 2142 1505 2143 1511
rect 2149 1505 2150 1511
rect 2142 1399 2150 1505
rect 2142 1393 2143 1399
rect 2149 1393 2150 1399
rect 2142 1295 2150 1393
rect 2142 1289 2143 1295
rect 2149 1289 2150 1295
rect 2142 1187 2150 1289
rect 2142 1181 2143 1187
rect 2149 1181 2150 1187
rect 2142 1079 2150 1181
rect 2142 1073 2143 1079
rect 2149 1073 2150 1079
rect 2142 963 2150 1073
rect 2142 957 2143 963
rect 2149 957 2150 963
rect 2142 859 2150 957
rect 2142 853 2143 859
rect 2149 853 2150 859
rect 2142 751 2150 853
rect 2142 745 2143 751
rect 2149 745 2150 751
rect 2142 647 2150 745
rect 2142 641 2143 647
rect 2149 641 2150 647
rect 2142 535 2150 641
rect 2142 529 2143 535
rect 2149 529 2150 535
rect 2142 431 2150 529
rect 2142 425 2143 431
rect 2149 425 2150 431
rect 2142 315 2150 425
rect 2142 309 2143 315
rect 2149 309 2150 315
rect 2142 79 2150 309
rect 2142 73 2143 79
rect 2149 73 2150 79
rect 2142 72 2150 73
rect 2154 2215 2162 2232
rect 2154 2209 2155 2215
rect 2161 2209 2162 2215
rect 2154 2107 2162 2209
rect 2154 2101 2155 2107
rect 2161 2101 2162 2107
rect 2154 2003 2162 2101
rect 2154 1997 2155 2003
rect 2161 1997 2162 2003
rect 2154 1891 2162 1997
rect 2154 1885 2155 1891
rect 2161 1885 2162 1891
rect 2154 1787 2162 1885
rect 2154 1781 2155 1787
rect 2161 1781 2162 1787
rect 2154 1679 2162 1781
rect 2154 1673 2155 1679
rect 2161 1673 2162 1679
rect 2154 1563 2162 1673
rect 2154 1557 2155 1563
rect 2161 1557 2162 1563
rect 2154 1455 2162 1557
rect 2154 1449 2155 1455
rect 2161 1449 2162 1455
rect 2154 1347 2162 1449
rect 2154 1341 2155 1347
rect 2161 1341 2162 1347
rect 2154 1239 2162 1341
rect 2154 1233 2155 1239
rect 2161 1233 2162 1239
rect 2154 1131 2162 1233
rect 2154 1125 2155 1131
rect 2161 1125 2162 1131
rect 2154 1023 2162 1125
rect 2154 1017 2155 1023
rect 2161 1017 2162 1023
rect 2154 911 2162 1017
rect 2154 905 2155 911
rect 2161 905 2162 911
rect 2154 807 2162 905
rect 2154 801 2155 807
rect 2161 801 2162 807
rect 2154 699 2162 801
rect 2154 693 2155 699
rect 2161 693 2162 699
rect 2154 591 2162 693
rect 2154 585 2155 591
rect 2161 585 2162 591
rect 2154 483 2162 585
rect 2154 477 2155 483
rect 2161 477 2162 483
rect 2154 375 2162 477
rect 2154 369 2155 375
rect 2161 369 2162 375
rect 2154 263 2162 369
rect 2154 257 2155 263
rect 2161 257 2162 263
rect 2154 131 2162 257
rect 2154 125 2155 131
rect 2161 125 2162 131
rect 2154 72 2162 125
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__147
timestamp 1731220619
transform 1 0 2112 0 1 2164
box 7 3 12 24
use welltap_svt  __well_tap__146
timestamp 1731220619
transform 1 0 1128 0 1 2164
box 7 3 12 24
use welltap_svt  __well_tap__145
timestamp 1731220619
transform 1 0 2112 0 -1 2156
box 7 3 12 24
use welltap_svt  __well_tap__144
timestamp 1731220619
transform 1 0 1128 0 -1 2156
box 7 3 12 24
use welltap_svt  __well_tap__143
timestamp 1731220619
transform 1 0 2112 0 1 2056
box 7 3 12 24
use welltap_svt  __well_tap__142
timestamp 1731220619
transform 1 0 1128 0 1 2056
box 7 3 12 24
use welltap_svt  __well_tap__141
timestamp 1731220619
transform 1 0 2112 0 -1 2048
box 7 3 12 24
use welltap_svt  __well_tap__140
timestamp 1731220619
transform 1 0 1128 0 -1 2048
box 7 3 12 24
use welltap_svt  __well_tap__139
timestamp 1731220619
transform 1 0 2112 0 1 1952
box 7 3 12 24
use welltap_svt  __well_tap__138
timestamp 1731220619
transform 1 0 1128 0 1 1952
box 7 3 12 24
use welltap_svt  __well_tap__137
timestamp 1731220619
transform 1 0 2112 0 -1 1940
box 7 3 12 24
use welltap_svt  __well_tap__136
timestamp 1731220619
transform 1 0 1128 0 -1 1940
box 7 3 12 24
use welltap_svt  __well_tap__135
timestamp 1731220619
transform 1 0 2112 0 1 1840
box 7 3 12 24
use welltap_svt  __well_tap__134
timestamp 1731220619
transform 1 0 1128 0 1 1840
box 7 3 12 24
use welltap_svt  __well_tap__133
timestamp 1731220619
transform 1 0 2112 0 -1 1832
box 7 3 12 24
use welltap_svt  __well_tap__132
timestamp 1731220619
transform 1 0 1128 0 -1 1832
box 7 3 12 24
use welltap_svt  __well_tap__131
timestamp 1731220619
transform 1 0 2112 0 1 1736
box 7 3 12 24
use welltap_svt  __well_tap__130
timestamp 1731220619
transform 1 0 1128 0 1 1736
box 7 3 12 24
use welltap_svt  __well_tap__129
timestamp 1731220619
transform 1 0 2112 0 -1 1728
box 7 3 12 24
use welltap_svt  __well_tap__128
timestamp 1731220619
transform 1 0 1128 0 -1 1728
box 7 3 12 24
use welltap_svt  __well_tap__127
timestamp 1731220619
transform 1 0 2112 0 1 1628
box 7 3 12 24
use welltap_svt  __well_tap__126
timestamp 1731220619
transform 1 0 1128 0 1 1628
box 7 3 12 24
use welltap_svt  __well_tap__125
timestamp 1731220619
transform 1 0 2112 0 -1 1608
box 7 3 12 24
use welltap_svt  __well_tap__124
timestamp 1731220619
transform 1 0 1128 0 -1 1608
box 7 3 12 24
use welltap_svt  __well_tap__123
timestamp 1731220619
transform 1 0 2112 0 1 1512
box 7 3 12 24
use welltap_svt  __well_tap__122
timestamp 1731220619
transform 1 0 1128 0 1 1512
box 7 3 12 24
use welltap_svt  __well_tap__121
timestamp 1731220619
transform 1 0 2112 0 -1 1504
box 7 3 12 24
use welltap_svt  __well_tap__120
timestamp 1731220619
transform 1 0 1128 0 -1 1504
box 7 3 12 24
use welltap_svt  __well_tap__119
timestamp 1731220619
transform 1 0 2112 0 1 1404
box 7 3 12 24
use welltap_svt  __well_tap__118
timestamp 1731220619
transform 1 0 1128 0 1 1404
box 7 3 12 24
use welltap_svt  __well_tap__117
timestamp 1731220619
transform 1 0 2112 0 -1 1392
box 7 3 12 24
use welltap_svt  __well_tap__116
timestamp 1731220619
transform 1 0 1128 0 -1 1392
box 7 3 12 24
use welltap_svt  __well_tap__115
timestamp 1731220619
transform 1 0 2112 0 1 1296
box 7 3 12 24
use welltap_svt  __well_tap__114
timestamp 1731220619
transform 1 0 1128 0 1 1296
box 7 3 12 24
use welltap_svt  __well_tap__113
timestamp 1731220619
transform 1 0 2112 0 -1 1288
box 7 3 12 24
use welltap_svt  __well_tap__112
timestamp 1731220619
transform 1 0 1128 0 -1 1288
box 7 3 12 24
use welltap_svt  __well_tap__111
timestamp 1731220619
transform 1 0 2112 0 1 1188
box 7 3 12 24
use welltap_svt  __well_tap__110
timestamp 1731220619
transform 1 0 1128 0 1 1188
box 7 3 12 24
use welltap_svt  __well_tap__109
timestamp 1731220619
transform 1 0 2112 0 -1 1180
box 7 3 12 24
use welltap_svt  __well_tap__108
timestamp 1731220619
transform 1 0 1128 0 -1 1180
box 7 3 12 24
use welltap_svt  __well_tap__107
timestamp 1731220619
transform 1 0 2112 0 1 1080
box 7 3 12 24
use welltap_svt  __well_tap__106
timestamp 1731220619
transform 1 0 1128 0 1 1080
box 7 3 12 24
use welltap_svt  __well_tap__105
timestamp 1731220619
transform 1 0 2112 0 -1 1072
box 7 3 12 24
use welltap_svt  __well_tap__104
timestamp 1731220619
transform 1 0 1128 0 -1 1072
box 7 3 12 24
use welltap_svt  __well_tap__103
timestamp 1731220619
transform 1 0 2112 0 1 972
box 7 3 12 24
use welltap_svt  __well_tap__102
timestamp 1731220619
transform 1 0 1128 0 1 972
box 7 3 12 24
use welltap_svt  __well_tap__101
timestamp 1731220619
transform 1 0 2112 0 -1 956
box 7 3 12 24
use welltap_svt  __well_tap__100
timestamp 1731220619
transform 1 0 1128 0 -1 956
box 7 3 12 24
use welltap_svt  __well_tap__99
timestamp 1731220619
transform 1 0 2112 0 1 860
box 7 3 12 24
use welltap_svt  __well_tap__98
timestamp 1731220619
transform 1 0 1128 0 1 860
box 7 3 12 24
use welltap_svt  __well_tap__97
timestamp 1731220619
transform 1 0 2112 0 -1 852
box 7 3 12 24
use welltap_svt  __well_tap__96
timestamp 1731220619
transform 1 0 1128 0 -1 852
box 7 3 12 24
use welltap_svt  __well_tap__95
timestamp 1731220619
transform 1 0 2112 0 1 756
box 7 3 12 24
use welltap_svt  __well_tap__94
timestamp 1731220619
transform 1 0 1128 0 1 756
box 7 3 12 24
use welltap_svt  __well_tap__93
timestamp 1731220619
transform 1 0 2112 0 -1 744
box 7 3 12 24
use welltap_svt  __well_tap__92
timestamp 1731220619
transform 1 0 1128 0 -1 744
box 7 3 12 24
use welltap_svt  __well_tap__91
timestamp 1731220619
transform 1 0 2112 0 1 648
box 7 3 12 24
use welltap_svt  __well_tap__90
timestamp 1731220619
transform 1 0 1128 0 1 648
box 7 3 12 24
use welltap_svt  __well_tap__89
timestamp 1731220619
transform 1 0 2112 0 -1 640
box 7 3 12 24
use welltap_svt  __well_tap__88
timestamp 1731220619
transform 1 0 1128 0 -1 640
box 7 3 12 24
use welltap_svt  __well_tap__87
timestamp 1731220619
transform 1 0 2112 0 1 540
box 7 3 12 24
use welltap_svt  __well_tap__86
timestamp 1731220619
transform 1 0 1128 0 1 540
box 7 3 12 24
use welltap_svt  __well_tap__85
timestamp 1731220619
transform 1 0 2112 0 -1 528
box 7 3 12 24
use welltap_svt  __well_tap__84
timestamp 1731220619
transform 1 0 1128 0 -1 528
box 7 3 12 24
use welltap_svt  __well_tap__83
timestamp 1731220619
transform 1 0 2112 0 1 432
box 7 3 12 24
use welltap_svt  __well_tap__82
timestamp 1731220619
transform 1 0 1128 0 1 432
box 7 3 12 24
use welltap_svt  __well_tap__81
timestamp 1731220619
transform 1 0 2112 0 -1 424
box 7 3 12 24
use welltap_svt  __well_tap__80
timestamp 1731220619
transform 1 0 1128 0 -1 424
box 7 3 12 24
use welltap_svt  __well_tap__79
timestamp 1731220619
transform 1 0 2112 0 1 324
box 7 3 12 24
use welltap_svt  __well_tap__78
timestamp 1731220619
transform 1 0 1128 0 1 324
box 7 3 12 24
use welltap_svt  __well_tap__77
timestamp 1731220619
transform 1 0 2112 0 -1 308
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220619
transform 1 0 1128 0 -1 308
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220619
transform 1 0 2112 0 1 212
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220619
transform 1 0 1128 0 1 212
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220619
transform 1 0 2112 0 -1 200
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220619
transform 1 0 1128 0 -1 200
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220619
transform 1 0 2112 0 1 80
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220619
transform 1 0 1128 0 1 80
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220619
transform 1 0 1088 0 1 1984
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220619
transform 1 0 104 0 1 1984
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220619
transform 1 0 1088 0 -1 1976
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220619
transform 1 0 104 0 -1 1976
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220619
transform 1 0 1088 0 1 1880
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220619
transform 1 0 104 0 1 1880
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220619
transform 1 0 1088 0 -1 1868
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220619
transform 1 0 104 0 -1 1868
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220619
transform 1 0 1088 0 1 1764
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220619
transform 1 0 104 0 1 1764
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220619
transform 1 0 1088 0 -1 1756
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220619
transform 1 0 104 0 -1 1756
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220619
transform 1 0 1088 0 1 1656
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220619
transform 1 0 104 0 1 1656
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220619
transform 1 0 1088 0 -1 1644
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220619
transform 1 0 104 0 -1 1644
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220619
transform 1 0 1088 0 1 1548
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220619
transform 1 0 104 0 1 1548
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220619
transform 1 0 1088 0 -1 1540
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220619
transform 1 0 104 0 -1 1540
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220619
transform 1 0 1088 0 1 1444
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220619
transform 1 0 104 0 1 1444
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220619
transform 1 0 1088 0 -1 1436
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220619
transform 1 0 104 0 -1 1436
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220619
transform 1 0 1088 0 1 1340
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220619
transform 1 0 104 0 1 1340
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220619
transform 1 0 1088 0 -1 1324
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220619
transform 1 0 104 0 -1 1324
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220619
transform 1 0 1088 0 1 1224
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220619
transform 1 0 104 0 1 1224
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220619
transform 1 0 1088 0 -1 1212
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220619
transform 1 0 104 0 -1 1212
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220619
transform 1 0 1088 0 1 1112
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220619
transform 1 0 104 0 1 1112
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220619
transform 1 0 1088 0 -1 1104
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220619
transform 1 0 104 0 -1 1104
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220619
transform 1 0 1088 0 1 1004
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220619
transform 1 0 104 0 1 1004
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220619
transform 1 0 1088 0 -1 992
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220619
transform 1 0 104 0 -1 992
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220619
transform 1 0 1088 0 1 892
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220619
transform 1 0 104 0 1 892
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220619
transform 1 0 1088 0 -1 880
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220619
transform 1 0 104 0 -1 880
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220619
transform 1 0 1088 0 1 784
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220619
transform 1 0 104 0 1 784
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220619
transform 1 0 1088 0 -1 776
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220619
transform 1 0 104 0 -1 776
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220619
transform 1 0 1088 0 1 680
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220619
transform 1 0 104 0 1 680
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220619
transform 1 0 1088 0 -1 672
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220619
transform 1 0 104 0 -1 672
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220619
transform 1 0 1088 0 1 568
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220619
transform 1 0 104 0 1 568
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220619
transform 1 0 1088 0 -1 556
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220619
transform 1 0 104 0 -1 556
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220619
transform 1 0 1088 0 1 452
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220619
transform 1 0 104 0 1 452
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220619
transform 1 0 1088 0 -1 440
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220619
transform 1 0 104 0 -1 440
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220619
transform 1 0 1088 0 1 336
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220619
transform 1 0 104 0 1 336
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220619
transform 1 0 1088 0 -1 324
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220619
transform 1 0 104 0 -1 324
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220619
transform 1 0 1088 0 1 220
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220619
transform 1 0 104 0 1 220
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220619
transform 1 0 1088 0 -1 200
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220619
transform 1 0 104 0 -1 200
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220619
transform 1 0 1088 0 1 88
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220619
transform 1 0 104 0 1 88
box 7 3 12 24
use _0_0std_0_0cells_0_0NOR2X1  tst_5999_6
timestamp 1731220619
transform 1 0 128 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5998_6
timestamp 1731220619
transform 1 0 168 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5997_6
timestamp 1731220619
transform 1 0 208 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5996_6
timestamp 1731220619
transform 1 0 248 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5995_6
timestamp 1731220619
transform 1 0 288 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5994_6
timestamp 1731220619
transform 1 0 328 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5993_6
timestamp 1731220619
transform 1 0 368 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5992_6
timestamp 1731220619
transform 1 0 408 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5991_6
timestamp 1731220619
transform 1 0 448 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5990_6
timestamp 1731220619
transform 1 0 488 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5989_6
timestamp 1731220619
transform 1 0 160 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5988_6
timestamp 1731220619
transform 1 0 200 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5987_6
timestamp 1731220619
transform 1 0 240 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5986_6
timestamp 1731220619
transform 1 0 288 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5985_6
timestamp 1731220619
transform 1 0 336 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5984_6
timestamp 1731220619
transform 1 0 392 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5983_6
timestamp 1731220619
transform 1 0 456 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5982_6
timestamp 1731220619
transform 1 0 280 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5981_6
timestamp 1731220619
transform 1 0 320 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5980_6
timestamp 1731220619
transform 1 0 360 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5979_6
timestamp 1731220619
transform 1 0 408 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5978_6
timestamp 1731220619
transform 1 0 464 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5977_6
timestamp 1731220619
transform 1 0 528 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5976_6
timestamp 1731220619
transform 1 0 600 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5975_6
timestamp 1731220619
transform 1 0 376 0 -1 328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5974_6
timestamp 1731220619
transform 1 0 416 0 -1 328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5973_6
timestamp 1731220619
transform 1 0 456 0 -1 328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5972_6
timestamp 1731220619
transform 1 0 496 0 -1 328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5971_6
timestamp 1731220619
transform 1 0 536 0 -1 328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5970_6
timestamp 1731220619
transform 1 0 584 0 -1 328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5969_6
timestamp 1731220619
transform 1 0 632 0 -1 328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5968_6
timestamp 1731220619
transform 1 0 680 0 -1 328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5967_6
timestamp 1731220619
transform 1 0 672 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5966_6
timestamp 1731220619
transform 1 0 664 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5965_6
timestamp 1731220619
transform 1 0 592 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5964_6
timestamp 1731220619
transform 1 0 520 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5963_6
timestamp 1731220619
transform 1 0 528 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5962_6
timestamp 1731220619
transform 1 0 568 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5961_6
timestamp 1731220619
transform 1 0 608 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5960_6
timestamp 1731220619
transform 1 0 648 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5959_6
timestamp 1731220619
transform 1 0 688 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5958_6
timestamp 1731220619
transform 1 0 728 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5957_6
timestamp 1731220619
transform 1 0 768 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5956_6
timestamp 1731220619
transform 1 0 808 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5955_6
timestamp 1731220619
transform 1 0 864 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5954_6
timestamp 1731220619
transform 1 0 928 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5953_6
timestamp 1731220619
transform 1 0 904 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5952_6
timestamp 1731220619
transform 1 0 824 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5951_6
timestamp 1731220619
transform 1 0 744 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5950_6
timestamp 1731220619
transform 1 0 800 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5949_6
timestamp 1731220619
transform 1 0 736 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5948_6
timestamp 1731220619
transform 1 0 728 0 -1 328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5947_6
timestamp 1731220619
transform 1 0 776 0 -1 328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5946_6
timestamp 1731220619
transform 1 0 824 0 -1 328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5945_6
timestamp 1731220619
transform 1 0 872 0 -1 328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5944_6
timestamp 1731220619
transform 1 0 856 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5943_6
timestamp 1731220619
transform 1 0 920 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5942_6
timestamp 1731220619
transform 1 0 984 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5941_6
timestamp 1731220619
transform 1 0 1040 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5940_6
timestamp 1731220619
transform 1 0 1040 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5939_6
timestamp 1731220619
transform 1 0 984 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5938_6
timestamp 1731220619
transform 1 0 992 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5937_6
timestamp 1731220619
transform 1 0 1040 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5936_6
timestamp 1731220619
transform 1 0 1152 0 1 76
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5935_6
timestamp 1731220619
transform 1 0 1192 0 1 76
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5934_6
timestamp 1731220619
transform 1 0 1232 0 1 76
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5933_6
timestamp 1731220619
transform 1 0 1272 0 1 76
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5932_6
timestamp 1731220619
transform 1 0 1312 0 1 76
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5931_6
timestamp 1731220619
transform 1 0 1360 0 1 76
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5930_6
timestamp 1731220619
transform 1 0 1424 0 1 76
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5929_6
timestamp 1731220619
transform 1 0 1488 0 1 76
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5928_6
timestamp 1731220619
transform 1 0 1176 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5927_6
timestamp 1731220619
transform 1 0 1224 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5926_6
timestamp 1731220619
transform 1 0 1288 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5925_6
timestamp 1731220619
transform 1 0 1352 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5924_6
timestamp 1731220619
transform 1 0 1424 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5923_6
timestamp 1731220619
transform 1 0 1504 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5922_6
timestamp 1731220619
transform 1 0 1256 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5921_6
timestamp 1731220619
transform 1 0 1296 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5920_6
timestamp 1731220619
transform 1 0 1336 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5919_6
timestamp 1731220619
transform 1 0 1376 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5918_6
timestamp 1731220619
transform 1 0 1416 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5917_6
timestamp 1731220619
transform 1 0 1456 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5916_6
timestamp 1731220619
transform 1 0 1496 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5915_6
timestamp 1731220619
transform 1 0 1344 0 -1 312
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5914_6
timestamp 1731220619
transform 1 0 1384 0 -1 312
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5913_6
timestamp 1731220619
transform 1 0 1424 0 -1 312
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5912_6
timestamp 1731220619
transform 1 0 1464 0 -1 312
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5911_6
timestamp 1731220619
transform 1 0 1504 0 -1 312
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5910_6
timestamp 1731220619
transform 1 0 1552 0 -1 312
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5909_6
timestamp 1731220619
transform 1 0 1608 0 -1 312
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5908_6
timestamp 1731220619
transform 1 0 1664 0 -1 312
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5907_6
timestamp 1731220619
transform 1 0 1728 0 -1 312
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5906_6
timestamp 1731220619
transform 1 0 1800 0 -1 312
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5905_6
timestamp 1731220619
transform 1 0 1536 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5904_6
timestamp 1731220619
transform 1 0 1592 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5903_6
timestamp 1731220619
transform 1 0 1664 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5902_6
timestamp 1731220619
transform 1 0 1752 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5901_6
timestamp 1731220619
transform 1 0 1856 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5900_6
timestamp 1731220619
transform 1 0 1968 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5899_6
timestamp 1731220619
transform 1 0 1584 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5898_6
timestamp 1731220619
transform 1 0 1656 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5897_6
timestamp 1731220619
transform 1 0 1728 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5896_6
timestamp 1731220619
transform 1 0 1800 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5895_6
timestamp 1731220619
transform 1 0 1552 0 1 76
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5894_6
timestamp 1731220619
transform 1 0 1608 0 1 76
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5893_6
timestamp 1731220619
transform 1 0 1664 0 1 76
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5892_6
timestamp 1731220619
transform 1 0 1712 0 1 76
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5891_6
timestamp 1731220619
transform 1 0 1760 0 1 76
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5890_6
timestamp 1731220619
transform 1 0 1800 0 1 76
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5889_6
timestamp 1731220619
transform 1 0 1848 0 1 76
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5888_6
timestamp 1731220619
transform 1 0 1896 0 1 76
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5887_6
timestamp 1731220619
transform 1 0 1944 0 1 76
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5886_6
timestamp 1731220619
transform 1 0 1872 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5885_6
timestamp 1731220619
transform 1 0 1944 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5884_6
timestamp 1731220619
transform 1 0 1984 0 1 76
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5883_6
timestamp 1731220619
transform 1 0 2024 0 1 76
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5882_6
timestamp 1731220619
transform 1 0 2064 0 1 76
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5881_6
timestamp 1731220619
transform 1 0 2064 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5880_6
timestamp 1731220619
transform 1 0 2016 0 -1 204
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5879_6
timestamp 1731220619
transform 1 0 2064 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5878_6
timestamp 1731220619
transform 1 0 2040 0 -1 312
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5877_6
timestamp 1731220619
transform 1 0 1960 0 -1 312
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5876_6
timestamp 1731220619
transform 1 0 1880 0 -1 312
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5875_6
timestamp 1731220619
transform 1 0 1856 0 1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5874_6
timestamp 1731220619
transform 1 0 1792 0 1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5873_6
timestamp 1731220619
transform 1 0 1720 0 1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5872_6
timestamp 1731220619
transform 1 0 1552 0 1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5871_6
timestamp 1731220619
transform 1 0 1640 0 1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5870_6
timestamp 1731220619
transform 1 0 1664 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5869_6
timestamp 1731220619
transform 1 0 1744 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5868_6
timestamp 1731220619
transform 1 0 1824 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5867_6
timestamp 1731220619
transform 1 0 1584 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5866_6
timestamp 1731220619
transform 1 0 1576 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5865_6
timestamp 1731220619
transform 1 0 1640 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5864_6
timestamp 1731220619
transform 1 0 1712 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5863_6
timestamp 1731220619
transform 1 0 1800 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5862_6
timestamp 1731220619
transform 1 0 1888 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5861_6
timestamp 1731220619
transform 1 0 1832 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5860_6
timestamp 1731220619
transform 1 0 1760 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5859_6
timestamp 1731220619
transform 1 0 1696 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5858_6
timestamp 1731220619
transform 1 0 1640 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5857_6
timestamp 1731220619
transform 1 0 1584 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5856_6
timestamp 1731220619
transform 1 0 1480 0 1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5855_6
timestamp 1731220619
transform 1 0 1560 0 1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5854_6
timestamp 1731220619
transform 1 0 1648 0 1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5853_6
timestamp 1731220619
transform 1 0 1744 0 1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5852_6
timestamp 1731220619
transform 1 0 1488 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5851_6
timestamp 1731220619
transform 1 0 1576 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5850_6
timestamp 1731220619
transform 1 0 1664 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5849_6
timestamp 1731220619
transform 1 0 1752 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5848_6
timestamp 1731220619
transform 1 0 1576 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5847_6
timestamp 1731220619
transform 1 0 1648 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5846_6
timestamp 1731220619
transform 1 0 1728 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5845_6
timestamp 1731220619
transform 1 0 1816 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5844_6
timestamp 1731220619
transform 1 0 1648 0 -1 748
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5843_6
timestamp 1731220619
transform 1 0 1704 0 -1 748
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5842_6
timestamp 1731220619
transform 1 0 1760 0 -1 748
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5841_6
timestamp 1731220619
transform 1 0 1824 0 -1 748
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5840_6
timestamp 1731220619
transform 1 0 1712 0 1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5839_6
timestamp 1731220619
transform 1 0 1616 0 1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5838_6
timestamp 1731220619
transform 1 0 1512 0 1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5837_6
timestamp 1731220619
transform 1 0 1536 0 -1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5836_6
timestamp 1731220619
transform 1 0 1624 0 -1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5835_6
timestamp 1731220619
transform 1 0 1704 0 -1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5834_6
timestamp 1731220619
transform 1 0 1656 0 1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5833_6
timestamp 1731220619
transform 1 0 1736 0 1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5832_6
timestamp 1731220619
transform 1 0 1776 0 -1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5831_6
timestamp 1731220619
transform 1 0 1848 0 -1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5830_6
timestamp 1731220619
transform 1 0 1928 0 -1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5829_6
timestamp 1731220619
transform 1 0 1808 0 1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5828_6
timestamp 1731220619
transform 1 0 1896 0 1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5827_6
timestamp 1731220619
transform 1 0 1992 0 1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5826_6
timestamp 1731220619
transform 1 0 1952 0 -1 748
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5825_6
timestamp 1731220619
transform 1 0 1888 0 -1 748
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5824_6
timestamp 1731220619
transform 1 0 1904 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5823_6
timestamp 1731220619
transform 1 0 1992 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5822_6
timestamp 1731220619
transform 1 0 1912 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5821_6
timestamp 1731220619
transform 1 0 1832 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5820_6
timestamp 1731220619
transform 1 0 1848 0 1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5819_6
timestamp 1731220619
transform 1 0 1960 0 1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5818_6
timestamp 1731220619
transform 1 0 1912 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5817_6
timestamp 1731220619
transform 1 0 1984 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5816_6
timestamp 1731220619
transform 1 0 1992 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5815_6
timestamp 1731220619
transform 1 0 1904 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5814_6
timestamp 1731220619
transform 1 0 1912 0 1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5813_6
timestamp 1731220619
transform 1 0 1968 0 1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5812_6
timestamp 1731220619
transform 1 0 2024 0 1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5811_6
timestamp 1731220619
transform 1 0 2064 0 1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5810_6
timestamp 1731220619
transform 1 0 2064 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5809_6
timestamp 1731220619
transform 1 0 2064 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5808_6
timestamp 1731220619
transform 1 0 2064 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5807_6
timestamp 1731220619
transform 1 0 2000 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5806_6
timestamp 1731220619
transform 1 0 2064 0 1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5805_6
timestamp 1731220619
transform 1 0 2000 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5804_6
timestamp 1731220619
transform 1 0 2064 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5803_6
timestamp 1731220619
transform 1 0 2064 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5802_6
timestamp 1731220619
transform 1 0 2016 0 -1 748
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5801_6
timestamp 1731220619
transform 1 0 2064 0 -1 748
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5800_6
timestamp 1731220619
transform 1 0 2064 0 1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5799_6
timestamp 1731220619
transform 1 0 2064 0 -1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5798_6
timestamp 1731220619
transform 1 0 2064 0 1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5797_6
timestamp 1731220619
transform 1 0 2064 0 -1 960
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5796_6
timestamp 1731220619
transform 1 0 2008 0 -1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5795_6
timestamp 1731220619
transform 1 0 1808 0 1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5794_6
timestamp 1731220619
transform 1 0 1880 0 1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5793_6
timestamp 1731220619
transform 1 0 1944 0 1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5792_6
timestamp 1731220619
transform 1 0 2016 0 1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5791_6
timestamp 1731220619
transform 1 0 2016 0 -1 960
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5790_6
timestamp 1731220619
transform 1 0 1944 0 -1 960
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5789_6
timestamp 1731220619
transform 1 0 1872 0 -1 960
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5788_6
timestamp 1731220619
transform 1 0 1808 0 -1 960
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5787_6
timestamp 1731220619
transform 1 0 1608 0 -1 960
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5786_6
timestamp 1731220619
transform 1 0 1680 0 -1 960
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5785_6
timestamp 1731220619
transform 1 0 1744 0 -1 960
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5784_6
timestamp 1731220619
transform 1 0 1784 0 1 968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5783_6
timestamp 1731220619
transform 1 0 1872 0 1 968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5782_6
timestamp 1731220619
transform 1 0 1704 0 1 968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5781_6
timestamp 1731220619
transform 1 0 1512 0 1 968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5780_6
timestamp 1731220619
transform 1 0 1568 0 1 968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5779_6
timestamp 1731220619
transform 1 0 1632 0 1 968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5778_6
timestamp 1731220619
transform 1 0 1656 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5777_6
timestamp 1731220619
transform 1 0 1752 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5776_6
timestamp 1731220619
transform 1 0 1856 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5775_6
timestamp 1731220619
transform 1 0 1576 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5774_6
timestamp 1731220619
transform 1 0 1504 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5773_6
timestamp 1731220619
transform 1 0 1408 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5772_6
timestamp 1731220619
transform 1 0 1448 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5771_6
timestamp 1731220619
transform 1 0 1480 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5770_6
timestamp 1731220619
transform 1 0 1560 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5769_6
timestamp 1731220619
transform 1 0 1648 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5768_6
timestamp 1731220619
transform 1 0 1744 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5767_6
timestamp 1731220619
transform 1 0 1848 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5766_6
timestamp 1731220619
transform 1 0 1552 0 -1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5765_6
timestamp 1731220619
transform 1 0 1624 0 -1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5764_6
timestamp 1731220619
transform 1 0 1704 0 -1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5763_6
timestamp 1731220619
transform 1 0 1792 0 -1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5762_6
timestamp 1731220619
transform 1 0 1880 0 -1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5761_6
timestamp 1731220619
transform 1 0 1616 0 1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5760_6
timestamp 1731220619
transform 1 0 1672 0 1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5759_6
timestamp 1731220619
transform 1 0 1728 0 1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5758_6
timestamp 1731220619
transform 1 0 1784 0 1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5757_6
timestamp 1731220619
transform 1 0 1840 0 1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5756_6
timestamp 1731220619
transform 1 0 1896 0 1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5755_6
timestamp 1731220619
transform 1 0 1648 0 -1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5754_6
timestamp 1731220619
transform 1 0 1736 0 -1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5753_6
timestamp 1731220619
transform 1 0 1824 0 -1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5752_6
timestamp 1731220619
transform 1 0 1912 0 -1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5751_6
timestamp 1731220619
transform 1 0 1672 0 1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5750_6
timestamp 1731220619
transform 1 0 1752 0 1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5749_6
timestamp 1731220619
transform 1 0 1824 0 1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5748_6
timestamp 1731220619
transform 1 0 1888 0 1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5747_6
timestamp 1731220619
transform 1 0 1952 0 1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5746_6
timestamp 1731220619
transform 1 0 2016 0 1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5745_6
timestamp 1731220619
transform 1 0 2000 0 -1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5744_6
timestamp 1731220619
transform 1 0 1960 0 1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5743_6
timestamp 1731220619
transform 1 0 1976 0 -1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5742_6
timestamp 1731220619
transform 1 0 1952 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5741_6
timestamp 1731220619
transform 1 0 1960 0 1 968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5740_6
timestamp 1731220619
transform 1 0 2056 0 1 968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5739_6
timestamp 1731220619
transform 1 0 1960 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5738_6
timestamp 1731220619
transform 1 0 2064 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5737_6
timestamp 1731220619
transform 1 0 2064 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5736_6
timestamp 1731220619
transform 1 0 2064 0 -1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5735_6
timestamp 1731220619
transform 1 0 2024 0 1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5734_6
timestamp 1731220619
transform 1 0 2064 0 1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5733_6
timestamp 1731220619
transform 1 0 2064 0 -1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5732_6
timestamp 1731220619
transform 1 0 2064 0 1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5731_6
timestamp 1731220619
transform 1 0 2064 0 -1 1396
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5730_6
timestamp 1731220619
transform 1 0 1984 0 -1 1396
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5729_6
timestamp 1731220619
transform 1 0 1968 0 1 1400
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5728_6
timestamp 1731220619
transform 1 0 2056 0 1 1400
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5727_6
timestamp 1731220619
transform 1 0 2056 0 -1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5726_6
timestamp 1731220619
transform 1 0 1984 0 -1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5725_6
timestamp 1731220619
transform 1 0 1992 0 1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5724_6
timestamp 1731220619
transform 1 0 1904 0 1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5723_6
timestamp 1731220619
transform 1 0 1816 0 1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5722_6
timestamp 1731220619
transform 1 0 1616 0 -1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5721_6
timestamp 1731220619
transform 1 0 1696 0 -1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5720_6
timestamp 1731220619
transform 1 0 1768 0 -1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5719_6
timestamp 1731220619
transform 1 0 1840 0 -1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5718_6
timestamp 1731220619
transform 1 0 1880 0 1 1400
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5717_6
timestamp 1731220619
transform 1 0 1800 0 1 1400
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5716_6
timestamp 1731220619
transform 1 0 1728 0 1 1400
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5715_6
timestamp 1731220619
transform 1 0 1544 0 1 1400
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5714_6
timestamp 1731220619
transform 1 0 1600 0 1 1400
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5713_6
timestamp 1731220619
transform 1 0 1664 0 1 1400
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5712_6
timestamp 1731220619
transform 1 0 1712 0 -1 1396
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5711_6
timestamp 1731220619
transform 1 0 1800 0 -1 1396
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5710_6
timestamp 1731220619
transform 1 0 1888 0 -1 1396
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5709_6
timestamp 1731220619
transform 1 0 1640 0 -1 1396
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5708_6
timestamp 1731220619
transform 1 0 1576 0 -1 1396
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5707_6
timestamp 1731220619
transform 1 0 1448 0 -1 1396
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5706_6
timestamp 1731220619
transform 1 0 1488 0 -1 1396
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5705_6
timestamp 1731220619
transform 1 0 1528 0 -1 1396
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5704_6
timestamp 1731220619
transform 1 0 1592 0 1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5703_6
timestamp 1731220619
transform 1 0 1496 0 1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5702_6
timestamp 1731220619
transform 1 0 1400 0 1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5701_6
timestamp 1731220619
transform 1 0 1408 0 -1 1396
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5700_6
timestamp 1731220619
transform 1 0 1368 0 -1 1396
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5699_6
timestamp 1731220619
transform 1 0 1328 0 -1 1396
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5698_6
timestamp 1731220619
transform 1 0 1272 0 1 1400
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5697_6
timestamp 1731220619
transform 1 0 1320 0 1 1400
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5696_6
timestamp 1731220619
transform 1 0 1376 0 1 1400
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5695_6
timestamp 1731220619
transform 1 0 1432 0 1 1400
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5694_6
timestamp 1731220619
transform 1 0 1488 0 1 1400
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5693_6
timestamp 1731220619
transform 1 0 1536 0 -1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5692_6
timestamp 1731220619
transform 1 0 1448 0 -1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5691_6
timestamp 1731220619
transform 1 0 1368 0 -1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5690_6
timestamp 1731220619
transform 1 0 1296 0 -1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5689_6
timestamp 1731220619
transform 1 0 1232 0 -1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5688_6
timestamp 1731220619
transform 1 0 1192 0 -1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5687_6
timestamp 1731220619
transform 1 0 1152 0 -1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5686_6
timestamp 1731220619
transform 1 0 1152 0 1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5685_6
timestamp 1731220619
transform 1 0 1192 0 1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5684_6
timestamp 1731220619
transform 1 0 1240 0 1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5683_6
timestamp 1731220619
transform 1 0 1312 0 1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5682_6
timestamp 1731220619
transform 1 0 1392 0 1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5681_6
timestamp 1731220619
transform 1 0 1472 0 1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5680_6
timestamp 1731220619
transform 1 0 1376 0 -1 1612
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5679_6
timestamp 1731220619
transform 1 0 1296 0 -1 1612
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5678_6
timestamp 1731220619
transform 1 0 1208 0 -1 1612
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5677_6
timestamp 1731220619
transform 1 0 1152 0 -1 1612
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5676_6
timestamp 1731220619
transform 1 0 1040 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5675_6
timestamp 1731220619
transform 1 0 896 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5674_6
timestamp 1731220619
transform 1 0 952 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5673_6
timestamp 1731220619
transform 1 0 1000 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5672_6
timestamp 1731220619
transform 1 0 1040 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5671_6
timestamp 1731220619
transform 1 0 912 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5670_6
timestamp 1731220619
transform 1 0 976 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5669_6
timestamp 1731220619
transform 1 0 984 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5668_6
timestamp 1731220619
transform 1 0 904 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5667_6
timestamp 1731220619
transform 1 0 824 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5666_6
timestamp 1731220619
transform 1 0 712 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5665_6
timestamp 1731220619
transform 1 0 784 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5664_6
timestamp 1731220619
transform 1 0 848 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5663_6
timestamp 1731220619
transform 1 0 840 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5662_6
timestamp 1731220619
transform 1 0 784 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5661_6
timestamp 1731220619
transform 1 0 720 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5660_6
timestamp 1731220619
transform 1 0 736 0 1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5659_6
timestamp 1731220619
transform 1 0 664 0 1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5658_6
timestamp 1731220619
transform 1 0 592 0 1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5657_6
timestamp 1731220619
transform 1 0 520 0 1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5656_6
timestamp 1731220619
transform 1 0 560 0 -1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5655_6
timestamp 1731220619
transform 1 0 648 0 -1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5654_6
timestamp 1731220619
transform 1 0 736 0 -1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5653_6
timestamp 1731220619
transform 1 0 672 0 1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5652_6
timestamp 1731220619
transform 1 0 760 0 1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5651_6
timestamp 1731220619
transform 1 0 848 0 1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5650_6
timestamp 1731220619
transform 1 0 792 0 -1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5649_6
timestamp 1731220619
transform 1 0 880 0 -1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5648_6
timestamp 1731220619
transform 1 0 920 0 1 1336
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5647_6
timestamp 1731220619
transform 1 0 848 0 1 1336
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5646_6
timestamp 1731220619
transform 1 0 776 0 1 1336
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5645_6
timestamp 1731220619
transform 1 0 776 0 -1 1328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5644_6
timestamp 1731220619
transform 1 0 856 0 -1 1328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5643_6
timestamp 1731220619
transform 1 0 936 0 -1 1328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5642_6
timestamp 1731220619
transform 1 0 1016 0 -1 1328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5641_6
timestamp 1731220619
transform 1 0 1040 0 1 1220
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5640_6
timestamp 1731220619
transform 1 0 912 0 1 1220
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5639_6
timestamp 1731220619
transform 1 0 976 0 -1 1216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5638_6
timestamp 1731220619
transform 1 0 936 0 1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5637_6
timestamp 1731220619
transform 1 0 992 0 -1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5636_6
timestamp 1731220619
transform 1 0 920 0 -1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5635_6
timestamp 1731220619
transform 1 0 568 0 1 1000
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5634_6
timestamp 1731220619
transform 1 0 504 0 1 1000
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5633_6
timestamp 1731220619
transform 1 0 520 0 -1 996
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5632_6
timestamp 1731220619
transform 1 0 464 0 -1 996
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5631_6
timestamp 1731220619
transform 1 0 448 0 1 888
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5630_6
timestamp 1731220619
transform 1 0 504 0 1 888
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5629_6
timestamp 1731220619
transform 1 0 560 0 1 888
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5628_6
timestamp 1731220619
transform 1 0 616 0 1 888
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5627_6
timestamp 1731220619
transform 1 0 616 0 -1 884
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5626_6
timestamp 1731220619
transform 1 0 544 0 -1 884
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5625_6
timestamp 1731220619
transform 1 0 472 0 -1 884
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5624_6
timestamp 1731220619
transform 1 0 480 0 1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5623_6
timestamp 1731220619
transform 1 0 560 0 1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5622_6
timestamp 1731220619
transform 1 0 640 0 1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5621_6
timestamp 1731220619
transform 1 0 560 0 -1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5620_6
timestamp 1731220619
transform 1 0 488 0 -1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5619_6
timestamp 1731220619
transform 1 0 536 0 1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5618_6
timestamp 1731220619
transform 1 0 464 0 1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5617_6
timestamp 1731220619
transform 1 0 384 0 1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5616_6
timestamp 1731220619
transform 1 0 392 0 -1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5615_6
timestamp 1731220619
transform 1 0 456 0 -1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5614_6
timestamp 1731220619
transform 1 0 328 0 -1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5613_6
timestamp 1731220619
transform 1 0 296 0 1 564
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5612_6
timestamp 1731220619
transform 1 0 344 0 1 564
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5611_6
timestamp 1731220619
transform 1 0 392 0 1 564
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5610_6
timestamp 1731220619
transform 1 0 416 0 -1 560
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5609_6
timestamp 1731220619
transform 1 0 368 0 -1 560
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5608_6
timestamp 1731220619
transform 1 0 320 0 -1 560
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5607_6
timestamp 1731220619
transform 1 0 352 0 1 448
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5606_6
timestamp 1731220619
transform 1 0 416 0 1 448
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5605_6
timestamp 1731220619
transform 1 0 472 0 1 448
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5604_6
timestamp 1731220619
transform 1 0 528 0 -1 444
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5603_6
timestamp 1731220619
transform 1 0 456 0 -1 444
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5602_6
timestamp 1731220619
transform 1 0 320 0 -1 444
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5601_6
timestamp 1731220619
transform 1 0 384 0 -1 444
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5600_6
timestamp 1731220619
transform 1 0 400 0 1 332
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5599_6
timestamp 1731220619
transform 1 0 480 0 1 332
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5598_6
timestamp 1731220619
transform 1 0 560 0 1 332
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5597_6
timestamp 1731220619
transform 1 0 328 0 1 332
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5596_6
timestamp 1731220619
transform 1 0 264 0 1 332
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5595_6
timestamp 1731220619
transform 1 0 208 0 1 332
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5594_6
timestamp 1731220619
transform 1 0 168 0 1 332
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5593_6
timestamp 1731220619
transform 1 0 168 0 -1 444
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5592_6
timestamp 1731220619
transform 1 0 208 0 -1 444
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5591_6
timestamp 1731220619
transform 1 0 256 0 -1 444
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5590_6
timestamp 1731220619
transform 1 0 128 0 1 448
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5589_6
timestamp 1731220619
transform 1 0 168 0 1 448
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5588_6
timestamp 1731220619
transform 1 0 224 0 1 448
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5587_6
timestamp 1731220619
transform 1 0 288 0 1 448
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5586_6
timestamp 1731220619
transform 1 0 272 0 -1 560
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5585_6
timestamp 1731220619
transform 1 0 216 0 -1 560
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5584_6
timestamp 1731220619
transform 1 0 168 0 -1 560
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5583_6
timestamp 1731220619
transform 1 0 128 0 -1 560
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5582_6
timestamp 1731220619
transform 1 0 128 0 1 564
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5581_6
timestamp 1731220619
transform 1 0 168 0 1 564
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5580_6
timestamp 1731220619
transform 1 0 208 0 1 564
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5579_6
timestamp 1731220619
transform 1 0 248 0 1 564
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5578_6
timestamp 1731220619
transform 1 0 128 0 -1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5577_6
timestamp 1731220619
transform 1 0 168 0 -1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5576_6
timestamp 1731220619
transform 1 0 208 0 -1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5575_6
timestamp 1731220619
transform 1 0 264 0 -1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5574_6
timestamp 1731220619
transform 1 0 304 0 1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5573_6
timestamp 1731220619
transform 1 0 232 0 1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5572_6
timestamp 1731220619
transform 1 0 168 0 1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5571_6
timestamp 1731220619
transform 1 0 208 0 -1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5570_6
timestamp 1731220619
transform 1 0 272 0 -1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5569_6
timestamp 1731220619
transform 1 0 344 0 -1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5568_6
timestamp 1731220619
transform 1 0 416 0 -1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5567_6
timestamp 1731220619
transform 1 0 408 0 1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5566_6
timestamp 1731220619
transform 1 0 336 0 1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5565_6
timestamp 1731220619
transform 1 0 272 0 1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5564_6
timestamp 1731220619
transform 1 0 296 0 -1 884
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5563_6
timestamp 1731220619
transform 1 0 344 0 -1 884
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5562_6
timestamp 1731220619
transform 1 0 408 0 -1 884
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5561_6
timestamp 1731220619
transform 1 0 256 0 1 888
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5560_6
timestamp 1731220619
transform 1 0 296 0 1 888
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5559_6
timestamp 1731220619
transform 1 0 344 0 1 888
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5558_6
timestamp 1731220619
transform 1 0 392 0 1 888
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5557_6
timestamp 1731220619
transform 1 0 400 0 -1 996
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5556_6
timestamp 1731220619
transform 1 0 336 0 -1 996
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5555_6
timestamp 1731220619
transform 1 0 272 0 -1 996
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5554_6
timestamp 1731220619
transform 1 0 128 0 -1 996
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5553_6
timestamp 1731220619
transform 1 0 168 0 -1 996
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5552_6
timestamp 1731220619
transform 1 0 216 0 -1 996
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5551_6
timestamp 1731220619
transform 1 0 312 0 1 1000
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5550_6
timestamp 1731220619
transform 1 0 376 0 1 1000
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5549_6
timestamp 1731220619
transform 1 0 440 0 1 1000
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5548_6
timestamp 1731220619
transform 1 0 128 0 1 1000
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5547_6
timestamp 1731220619
transform 1 0 168 0 1 1000
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5546_6
timestamp 1731220619
transform 1 0 208 0 1 1000
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5545_6
timestamp 1731220619
transform 1 0 248 0 1 1000
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5544_6
timestamp 1731220619
transform 1 0 152 0 -1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5543_6
timestamp 1731220619
transform 1 0 192 0 -1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5542_6
timestamp 1731220619
transform 1 0 248 0 -1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5541_6
timestamp 1731220619
transform 1 0 312 0 -1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5540_6
timestamp 1731220619
transform 1 0 392 0 -1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5539_6
timestamp 1731220619
transform 1 0 472 0 -1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5538_6
timestamp 1731220619
transform 1 0 552 0 -1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5537_6
timestamp 1731220619
transform 1 0 392 0 1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5536_6
timestamp 1731220619
transform 1 0 432 0 1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5535_6
timestamp 1731220619
transform 1 0 472 0 1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5534_6
timestamp 1731220619
transform 1 0 520 0 1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5533_6
timestamp 1731220619
transform 1 0 568 0 1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5532_6
timestamp 1731220619
transform 1 0 616 0 1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5531_6
timestamp 1731220619
transform 1 0 488 0 -1 1216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5530_6
timestamp 1731220619
transform 1 0 440 0 -1 1216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5529_6
timestamp 1731220619
transform 1 0 392 0 -1 1216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5528_6
timestamp 1731220619
transform 1 0 264 0 -1 1216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5527_6
timestamp 1731220619
transform 1 0 304 0 -1 1216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5526_6
timestamp 1731220619
transform 1 0 344 0 -1 1216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5525_6
timestamp 1731220619
transform 1 0 392 0 1 1220
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5524_6
timestamp 1731220619
transform 1 0 312 0 1 1220
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5523_6
timestamp 1731220619
transform 1 0 248 0 1 1220
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5522_6
timestamp 1731220619
transform 1 0 128 0 1 1220
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5521_6
timestamp 1731220619
transform 1 0 168 0 1 1220
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5520_6
timestamp 1731220619
transform 1 0 208 0 1 1220
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5519_6
timestamp 1731220619
transform 1 0 248 0 -1 1328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5518_6
timestamp 1731220619
transform 1 0 312 0 -1 1328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5517_6
timestamp 1731220619
transform 1 0 208 0 -1 1328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5516_6
timestamp 1731220619
transform 1 0 168 0 -1 1328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5515_6
timestamp 1731220619
transform 1 0 128 0 -1 1328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5514_6
timestamp 1731220619
transform 1 0 128 0 1 1336
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5513_6
timestamp 1731220619
transform 1 0 128 0 -1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5512_6
timestamp 1731220619
transform 1 0 128 0 1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5511_6
timestamp 1731220619
transform 1 0 192 0 1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5510_6
timestamp 1731220619
transform 1 0 128 0 -1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5509_6
timestamp 1731220619
transform 1 0 168 0 -1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5508_6
timestamp 1731220619
transform 1 0 224 0 1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5507_6
timestamp 1731220619
transform 1 0 168 0 1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5506_6
timestamp 1731220619
transform 1 0 128 0 1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5505_6
timestamp 1731220619
transform 1 0 128 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5504_6
timestamp 1731220619
transform 1 0 176 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5503_6
timestamp 1731220619
transform 1 0 128 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5502_6
timestamp 1731220619
transform 1 0 192 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5501_6
timestamp 1731220619
transform 1 0 272 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5500_6
timestamp 1731220619
transform 1 0 288 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5499_6
timestamp 1731220619
transform 1 0 224 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5498_6
timestamp 1731220619
transform 1 0 264 0 1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5497_6
timestamp 1731220619
transform 1 0 208 0 1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5496_6
timestamp 1731220619
transform 1 0 144 0 1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5495_6
timestamp 1731220619
transform 1 0 192 0 -1 1872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5494_6
timestamp 1731220619
transform 1 0 264 0 -1 1872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5493_6
timestamp 1731220619
transform 1 0 128 0 -1 1872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5492_6
timestamp 1731220619
transform 1 0 128 0 1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5491_6
timestamp 1731220619
transform 1 0 168 0 1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5490_6
timestamp 1731220619
transform 1 0 224 0 1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5489_6
timestamp 1731220619
transform 1 0 288 0 1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5488_6
timestamp 1731220619
transform 1 0 304 0 -1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5487_6
timestamp 1731220619
transform 1 0 240 0 -1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5486_6
timestamp 1731220619
transform 1 0 184 0 -1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5485_6
timestamp 1731220619
transform 1 0 184 0 1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5484_6
timestamp 1731220619
transform 1 0 224 0 1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5483_6
timestamp 1731220619
transform 1 0 280 0 1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5482_6
timestamp 1731220619
transform 1 0 344 0 1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5481_6
timestamp 1731220619
transform 1 0 416 0 1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5480_6
timestamp 1731220619
transform 1 0 488 0 1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5479_6
timestamp 1731220619
transform 1 0 568 0 1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5478_6
timestamp 1731220619
transform 1 0 512 0 -1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5477_6
timestamp 1731220619
transform 1 0 440 0 -1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5476_6
timestamp 1731220619
transform 1 0 368 0 -1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5475_6
timestamp 1731220619
transform 1 0 360 0 1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5474_6
timestamp 1731220619
transform 1 0 424 0 1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5473_6
timestamp 1731220619
transform 1 0 488 0 1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5472_6
timestamp 1731220619
transform 1 0 448 0 -1 1872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5471_6
timestamp 1731220619
transform 1 0 328 0 -1 1872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5470_6
timestamp 1731220619
transform 1 0 392 0 -1 1872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5469_6
timestamp 1731220619
transform 1 0 424 0 1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5468_6
timestamp 1731220619
transform 1 0 376 0 1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5467_6
timestamp 1731220619
transform 1 0 320 0 1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5466_6
timestamp 1731220619
transform 1 0 344 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5465_6
timestamp 1731220619
transform 1 0 408 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5464_6
timestamp 1731220619
transform 1 0 472 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5463_6
timestamp 1731220619
transform 1 0 536 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5462_6
timestamp 1731220619
transform 1 0 544 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5461_6
timestamp 1731220619
transform 1 0 456 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5460_6
timestamp 1731220619
transform 1 0 360 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5459_6
timestamp 1731220619
transform 1 0 256 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5458_6
timestamp 1731220619
transform 1 0 336 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5457_6
timestamp 1731220619
transform 1 0 416 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5456_6
timestamp 1731220619
transform 1 0 496 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5455_6
timestamp 1731220619
transform 1 0 448 0 1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5454_6
timestamp 1731220619
transform 1 0 368 0 1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5453_6
timestamp 1731220619
transform 1 0 296 0 1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5452_6
timestamp 1731220619
transform 1 0 224 0 -1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5451_6
timestamp 1731220619
transform 1 0 304 0 -1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5450_6
timestamp 1731220619
transform 1 0 384 0 -1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5449_6
timestamp 1731220619
transform 1 0 472 0 -1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5448_6
timestamp 1731220619
transform 1 0 352 0 1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5447_6
timestamp 1731220619
transform 1 0 272 0 1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5446_6
timestamp 1731220619
transform 1 0 256 0 -1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5445_6
timestamp 1731220619
transform 1 0 184 0 -1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5444_6
timestamp 1731220619
transform 1 0 168 0 1 1336
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5443_6
timestamp 1731220619
transform 1 0 232 0 1 1336
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5442_6
timestamp 1731220619
transform 1 0 384 0 -1 1328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5441_6
timestamp 1731220619
transform 1 0 456 0 -1 1328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5440_6
timestamp 1731220619
transform 1 0 296 0 1 1336
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5439_6
timestamp 1731220619
transform 1 0 360 0 1 1336
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5438_6
timestamp 1731220619
transform 1 0 432 0 1 1336
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5437_6
timestamp 1731220619
transform 1 0 496 0 1 1336
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5436_6
timestamp 1731220619
transform 1 0 472 0 -1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5435_6
timestamp 1731220619
transform 1 0 328 0 -1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5434_6
timestamp 1731220619
transform 1 0 400 0 -1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5433_6
timestamp 1731220619
transform 1 0 432 0 1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5432_6
timestamp 1731220619
transform 1 0 512 0 1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5431_6
timestamp 1731220619
transform 1 0 592 0 1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5430_6
timestamp 1731220619
transform 1 0 624 0 -1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5429_6
timestamp 1731220619
transform 1 0 704 0 -1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5428_6
timestamp 1731220619
transform 1 0 544 0 -1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5427_6
timestamp 1731220619
transform 1 0 568 0 1 1336
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5426_6
timestamp 1731220619
transform 1 0 640 0 1 1336
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5425_6
timestamp 1731220619
transform 1 0 704 0 1 1336
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5424_6
timestamp 1731220619
transform 1 0 696 0 -1 1328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5423_6
timestamp 1731220619
transform 1 0 616 0 -1 1328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5422_6
timestamp 1731220619
transform 1 0 536 0 -1 1328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5421_6
timestamp 1731220619
transform 1 0 480 0 1 1220
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5420_6
timestamp 1731220619
transform 1 0 576 0 1 1220
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5419_6
timestamp 1731220619
transform 1 0 680 0 1 1220
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5418_6
timestamp 1731220619
transform 1 0 792 0 1 1220
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5417_6
timestamp 1731220619
transform 1 0 544 0 -1 1216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5416_6
timestamp 1731220619
transform 1 0 600 0 -1 1216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5415_6
timestamp 1731220619
transform 1 0 664 0 -1 1216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5414_6
timestamp 1731220619
transform 1 0 736 0 -1 1216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5413_6
timestamp 1731220619
transform 1 0 808 0 -1 1216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5412_6
timestamp 1731220619
transform 1 0 888 0 -1 1216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5411_6
timestamp 1731220619
transform 1 0 664 0 1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5410_6
timestamp 1731220619
transform 1 0 712 0 1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5409_6
timestamp 1731220619
transform 1 0 768 0 1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5408_6
timestamp 1731220619
transform 1 0 824 0 1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5407_6
timestamp 1731220619
transform 1 0 880 0 1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5406_6
timestamp 1731220619
transform 1 0 632 0 -1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5405_6
timestamp 1731220619
transform 1 0 704 0 -1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5404_6
timestamp 1731220619
transform 1 0 776 0 -1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5403_6
timestamp 1731220619
transform 1 0 848 0 -1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5402_6
timestamp 1731220619
transform 1 0 856 0 1 1000
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5401_6
timestamp 1731220619
transform 1 0 792 0 1 1000
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5400_6
timestamp 1731220619
transform 1 0 736 0 1 1000
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5399_6
timestamp 1731220619
transform 1 0 680 0 1 1000
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5398_6
timestamp 1731220619
transform 1 0 624 0 1 1000
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5397_6
timestamp 1731220619
transform 1 0 576 0 -1 996
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5396_6
timestamp 1731220619
transform 1 0 624 0 -1 996
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5395_6
timestamp 1731220619
transform 1 0 680 0 -1 996
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5394_6
timestamp 1731220619
transform 1 0 736 0 -1 996
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5393_6
timestamp 1731220619
transform 1 0 792 0 -1 996
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5392_6
timestamp 1731220619
transform 1 0 680 0 1 888
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5391_6
timestamp 1731220619
transform 1 0 744 0 1 888
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5390_6
timestamp 1731220619
transform 1 0 808 0 1 888
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5389_6
timestamp 1731220619
transform 1 0 872 0 1 888
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5388_6
timestamp 1731220619
transform 1 0 936 0 1 888
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5387_6
timestamp 1731220619
transform 1 0 688 0 -1 884
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5386_6
timestamp 1731220619
transform 1 0 760 0 -1 884
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5385_6
timestamp 1731220619
transform 1 0 824 0 -1 884
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5384_6
timestamp 1731220619
transform 1 0 880 0 -1 884
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5383_6
timestamp 1731220619
transform 1 0 720 0 1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5382_6
timestamp 1731220619
transform 1 0 792 0 1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5381_6
timestamp 1731220619
transform 1 0 936 0 -1 884
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5380_6
timestamp 1731220619
transform 1 0 1000 0 -1 884
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5379_6
timestamp 1731220619
transform 1 0 1040 0 -1 884
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5378_6
timestamp 1731220619
transform 1 0 1000 0 1 888
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5377_6
timestamp 1731220619
transform 1 0 1040 0 1 888
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5376_6
timestamp 1731220619
transform 1 0 1152 0 -1 960
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5375_6
timestamp 1731220619
transform 1 0 1200 0 -1 960
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5374_6
timestamp 1731220619
transform 1 0 1152 0 1 968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5373_6
timestamp 1731220619
transform 1 0 1192 0 1 968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5372_6
timestamp 1731220619
transform 1 0 1192 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5371_6
timestamp 1731220619
transform 1 0 1152 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5370_6
timestamp 1731220619
transform 1 0 1040 0 -1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5369_6
timestamp 1731220619
transform 1 0 1000 0 1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5368_6
timestamp 1731220619
transform 1 0 1040 0 1 1108
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5367_6
timestamp 1731220619
transform 1 0 1152 0 -1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5366_6
timestamp 1731220619
transform 1 0 1200 0 -1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5365_6
timestamp 1731220619
transform 1 0 1272 0 -1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5364_6
timestamp 1731220619
transform 1 0 1184 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5363_6
timestamp 1731220619
transform 1 0 1264 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5362_6
timestamp 1731220619
transform 1 0 1296 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5361_6
timestamp 1731220619
transform 1 0 1240 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5360_6
timestamp 1731220619
transform 1 0 1232 0 1 968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5359_6
timestamp 1731220619
transform 1 0 1288 0 1 968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5358_6
timestamp 1731220619
transform 1 0 1344 0 1 968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5357_6
timestamp 1731220619
transform 1 0 1368 0 -1 960
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5356_6
timestamp 1731220619
transform 1 0 1280 0 -1 960
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5355_6
timestamp 1731220619
transform 1 0 1232 0 1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5354_6
timestamp 1731220619
transform 1 0 1312 0 1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5353_6
timestamp 1731220619
transform 1 0 1400 0 1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5352_6
timestamp 1731220619
transform 1 0 1352 0 -1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5351_6
timestamp 1731220619
transform 1 0 1240 0 -1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5350_6
timestamp 1731220619
transform 1 0 1152 0 -1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5349_6
timestamp 1731220619
transform 1 0 1152 0 1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5348_6
timestamp 1731220619
transform 1 0 1040 0 1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5347_6
timestamp 1731220619
transform 1 0 1040 0 -1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5346_6
timestamp 1731220619
transform 1 0 1000 0 -1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5345_6
timestamp 1731220619
transform 1 0 952 0 -1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5344_6
timestamp 1731220619
transform 1 0 992 0 1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5343_6
timestamp 1731220619
transform 1 0 920 0 1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5342_6
timestamp 1731220619
transform 1 0 856 0 1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5341_6
timestamp 1731220619
transform 1 0 904 0 -1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5340_6
timestamp 1731220619
transform 1 0 856 0 -1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5339_6
timestamp 1731220619
transform 1 0 808 0 -1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5338_6
timestamp 1731220619
transform 1 0 632 0 -1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5337_6
timestamp 1731220619
transform 1 0 696 0 -1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5336_6
timestamp 1731220619
transform 1 0 752 0 -1 780
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5335_6
timestamp 1731220619
transform 1 0 792 0 1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5334_6
timestamp 1731220619
transform 1 0 856 0 1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5333_6
timestamp 1731220619
transform 1 0 920 0 1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5332_6
timestamp 1731220619
transform 1 0 728 0 1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5331_6
timestamp 1731220619
transform 1 0 608 0 1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5330_6
timestamp 1731220619
transform 1 0 672 0 1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5329_6
timestamp 1731220619
transform 1 0 696 0 -1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5328_6
timestamp 1731220619
transform 1 0 752 0 -1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5327_6
timestamp 1731220619
transform 1 0 816 0 -1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5326_6
timestamp 1731220619
transform 1 0 640 0 -1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5325_6
timestamp 1731220619
transform 1 0 520 0 -1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5324_6
timestamp 1731220619
transform 1 0 584 0 -1 676
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5323_6
timestamp 1731220619
transform 1 0 624 0 1 564
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5322_6
timestamp 1731220619
transform 1 0 672 0 1 564
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5321_6
timestamp 1731220619
transform 1 0 720 0 1 564
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5320_6
timestamp 1731220619
transform 1 0 576 0 1 564
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5319_6
timestamp 1731220619
transform 1 0 528 0 1 564
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5318_6
timestamp 1731220619
transform 1 0 480 0 1 564
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5317_6
timestamp 1731220619
transform 1 0 432 0 1 564
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5316_6
timestamp 1731220619
transform 1 0 456 0 -1 560
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5315_6
timestamp 1731220619
transform 1 0 504 0 -1 560
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5314_6
timestamp 1731220619
transform 1 0 552 0 -1 560
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5313_6
timestamp 1731220619
transform 1 0 600 0 -1 560
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5312_6
timestamp 1731220619
transform 1 0 648 0 -1 560
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5311_6
timestamp 1731220619
transform 1 0 696 0 -1 560
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5310_6
timestamp 1731220619
transform 1 0 744 0 -1 560
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5309_6
timestamp 1731220619
transform 1 0 528 0 1 448
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5308_6
timestamp 1731220619
transform 1 0 584 0 1 448
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5307_6
timestamp 1731220619
transform 1 0 632 0 1 448
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5306_6
timestamp 1731220619
transform 1 0 680 0 1 448
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5305_6
timestamp 1731220619
transform 1 0 728 0 1 448
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5304_6
timestamp 1731220619
transform 1 0 784 0 1 448
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5303_6
timestamp 1731220619
transform 1 0 840 0 1 448
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5302_6
timestamp 1731220619
transform 1 0 600 0 -1 444
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5301_6
timestamp 1731220619
transform 1 0 672 0 -1 444
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5300_6
timestamp 1731220619
transform 1 0 736 0 -1 444
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5299_6
timestamp 1731220619
transform 1 0 800 0 -1 444
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5298_6
timestamp 1731220619
transform 1 0 864 0 -1 444
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5297_6
timestamp 1731220619
transform 1 0 936 0 -1 444
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5296_6
timestamp 1731220619
transform 1 0 632 0 1 332
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5295_6
timestamp 1731220619
transform 1 0 704 0 1 332
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5294_6
timestamp 1731220619
transform 1 0 768 0 1 332
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5293_6
timestamp 1731220619
transform 1 0 832 0 1 332
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5292_6
timestamp 1731220619
transform 1 0 888 0 1 332
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5291_6
timestamp 1731220619
transform 1 0 944 0 1 332
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5290_6
timestamp 1731220619
transform 1 0 1000 0 1 332
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5289_6
timestamp 1731220619
transform 1 0 920 0 -1 328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5288_6
timestamp 1731220619
transform 1 0 960 0 -1 328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5287_6
timestamp 1731220619
transform 1 0 1000 0 -1 328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5286_6
timestamp 1731220619
transform 1 0 1040 0 -1 328
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5285_6
timestamp 1731220619
transform 1 0 1040 0 1 332
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5284_6
timestamp 1731220619
transform 1 0 1152 0 1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5283_6
timestamp 1731220619
transform 1 0 1240 0 1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5282_6
timestamp 1731220619
transform 1 0 1352 0 1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5281_6
timestamp 1731220619
transform 1 0 1456 0 1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5280_6
timestamp 1731220619
transform 1 0 1152 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5279_6
timestamp 1731220619
transform 1 0 1192 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5278_6
timestamp 1731220619
transform 1 0 1248 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5277_6
timestamp 1731220619
transform 1 0 1328 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5276_6
timestamp 1731220619
transform 1 0 1408 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5275_6
timestamp 1731220619
transform 1 0 1496 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5274_6
timestamp 1731220619
transform 1 0 1288 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5273_6
timestamp 1731220619
transform 1 0 1328 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5272_6
timestamp 1731220619
transform 1 0 1368 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5271_6
timestamp 1731220619
transform 1 0 1416 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5270_6
timestamp 1731220619
transform 1 0 1464 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5269_6
timestamp 1731220619
transform 1 0 1520 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5268_6
timestamp 1731220619
transform 1 0 1536 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5267_6
timestamp 1731220619
transform 1 0 1496 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5266_6
timestamp 1731220619
transform 1 0 1456 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5265_6
timestamp 1731220619
transform 1 0 1416 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5264_6
timestamp 1731220619
transform 1 0 1296 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5263_6
timestamp 1731220619
transform 1 0 1336 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5262_6
timestamp 1731220619
transform 1 0 1376 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5261_6
timestamp 1731220619
transform 1 0 1408 0 1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5260_6
timestamp 1731220619
transform 1 0 1352 0 1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5259_6
timestamp 1731220619
transform 1 0 1312 0 1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5258_6
timestamp 1731220619
transform 1 0 1272 0 1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5257_6
timestamp 1731220619
transform 1 0 1232 0 1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5256_6
timestamp 1731220619
transform 1 0 1192 0 1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5255_6
timestamp 1731220619
transform 1 0 1152 0 1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5254_6
timestamp 1731220619
transform 1 0 1152 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5253_6
timestamp 1731220619
transform 1 0 1192 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5252_6
timestamp 1731220619
transform 1 0 1232 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5251_6
timestamp 1731220619
transform 1 0 1272 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5250_6
timestamp 1731220619
transform 1 0 1336 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5249_6
timestamp 1731220619
transform 1 0 1408 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5248_6
timestamp 1731220619
transform 1 0 1240 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5247_6
timestamp 1731220619
transform 1 0 1280 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5246_6
timestamp 1731220619
transform 1 0 1328 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5245_6
timestamp 1731220619
transform 1 0 1384 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5244_6
timestamp 1731220619
transform 1 0 1440 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5243_6
timestamp 1731220619
transform 1 0 1504 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5242_6
timestamp 1731220619
transform 1 0 1328 0 -1 748
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5241_6
timestamp 1731220619
transform 1 0 1368 0 -1 748
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5240_6
timestamp 1731220619
transform 1 0 1408 0 -1 748
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5239_6
timestamp 1731220619
transform 1 0 1448 0 -1 748
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5238_6
timestamp 1731220619
transform 1 0 1496 0 -1 748
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5237_6
timestamp 1731220619
transform 1 0 1544 0 -1 748
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5236_6
timestamp 1731220619
transform 1 0 1592 0 -1 748
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5235_6
timestamp 1731220619
transform 1 0 1272 0 1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5234_6
timestamp 1731220619
transform 1 0 1400 0 1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5233_6
timestamp 1731220619
transform 1 0 1448 0 -1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5232_6
timestamp 1731220619
transform 1 0 1488 0 1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5231_6
timestamp 1731220619
transform 1 0 1576 0 1 856
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5230_6
timestamp 1731220619
transform 1 0 1528 0 -1 960
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5229_6
timestamp 1731220619
transform 1 0 1448 0 -1 960
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5228_6
timestamp 1731220619
transform 1 0 1456 0 1 968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5227_6
timestamp 1731220619
transform 1 0 1400 0 1 968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5226_6
timestamp 1731220619
transform 1 0 1392 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5225_6
timestamp 1731220619
transform 1 0 1344 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5224_6
timestamp 1731220619
transform 1 0 1336 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5223_6
timestamp 1731220619
transform 1 0 1344 0 -1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5222_6
timestamp 1731220619
transform 1 0 1416 0 -1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5221_6
timestamp 1731220619
transform 1 0 1480 0 -1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5220_6
timestamp 1731220619
transform 1 0 1488 0 1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5219_6
timestamp 1731220619
transform 1 0 1552 0 1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5218_6
timestamp 1731220619
transform 1 0 1424 0 1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5217_6
timestamp 1731220619
transform 1 0 1280 0 1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5216_6
timestamp 1731220619
transform 1 0 1320 0 1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5215_6
timestamp 1731220619
transform 1 0 1368 0 1 1184
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5214_6
timestamp 1731220619
transform 1 0 1384 0 -1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5213_6
timestamp 1731220619
transform 1 0 1472 0 -1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5212_6
timestamp 1731220619
transform 1 0 1560 0 -1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5211_6
timestamp 1731220619
transform 1 0 1168 0 -1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5210_6
timestamp 1731220619
transform 1 0 1224 0 -1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5209_6
timestamp 1731220619
transform 1 0 1296 0 -1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5208_6
timestamp 1731220619
transform 1 0 1304 0 1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5207_6
timestamp 1731220619
transform 1 0 1216 0 1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5206_6
timestamp 1731220619
transform 1 0 1152 0 1 1292
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5205_6
timestamp 1731220619
transform 1 0 1040 0 1 1336
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5204_6
timestamp 1731220619
transform 1 0 992 0 1 1336
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5203_6
timestamp 1731220619
transform 1 0 968 0 -1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5202_6
timestamp 1731220619
transform 1 0 1040 0 -1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5201_6
timestamp 1731220619
transform 1 0 1024 0 1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5200_6
timestamp 1731220619
transform 1 0 936 0 1 1440
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5199_6
timestamp 1731220619
transform 1 0 992 0 -1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5198_6
timestamp 1731220619
transform 1 0 904 0 -1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5197_6
timestamp 1731220619
transform 1 0 816 0 -1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5196_6
timestamp 1731220619
transform 1 0 880 0 1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5195_6
timestamp 1731220619
transform 1 0 808 0 1 1544
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5194_6
timestamp 1731220619
transform 1 0 648 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5193_6
timestamp 1731220619
transform 1 0 576 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5192_6
timestamp 1731220619
transform 1 0 632 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5191_6
timestamp 1731220619
transform 1 0 608 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5190_6
timestamp 1731220619
transform 1 0 680 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5189_6
timestamp 1731220619
transform 1 0 752 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5188_6
timestamp 1731220619
transform 1 0 720 0 1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5187_6
timestamp 1731220619
transform 1 0 664 0 1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5186_6
timestamp 1731220619
transform 1 0 472 0 1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5185_6
timestamp 1731220619
transform 1 0 520 0 1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5184_6
timestamp 1731220619
transform 1 0 568 0 1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5183_6
timestamp 1731220619
transform 1 0 616 0 1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5182_6
timestamp 1731220619
transform 1 0 496 0 -1 1872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5181_6
timestamp 1731220619
transform 1 0 544 0 -1 1872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5180_6
timestamp 1731220619
transform 1 0 592 0 -1 1872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5179_6
timestamp 1731220619
transform 1 0 640 0 -1 1872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5178_6
timestamp 1731220619
transform 1 0 688 0 -1 1872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5177_6
timestamp 1731220619
transform 1 0 744 0 -1 1872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5176_6
timestamp 1731220619
transform 1 0 552 0 1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5175_6
timestamp 1731220619
transform 1 0 608 0 1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5174_6
timestamp 1731220619
transform 1 0 664 0 1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5173_6
timestamp 1731220619
transform 1 0 720 0 1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5172_6
timestamp 1731220619
transform 1 0 776 0 1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5171_6
timestamp 1731220619
transform 1 0 840 0 1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5170_6
timestamp 1731220619
transform 1 0 584 0 -1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5169_6
timestamp 1731220619
transform 1 0 648 0 -1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5168_6
timestamp 1731220619
transform 1 0 712 0 -1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5167_6
timestamp 1731220619
transform 1 0 768 0 -1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5166_6
timestamp 1731220619
transform 1 0 816 0 -1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5165_6
timestamp 1731220619
transform 1 0 864 0 -1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5164_6
timestamp 1731220619
transform 1 0 640 0 1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5163_6
timestamp 1731220619
transform 1 0 712 0 1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5162_6
timestamp 1731220619
transform 1 0 776 0 1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5161_6
timestamp 1731220619
transform 1 0 832 0 1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5160_6
timestamp 1731220619
transform 1 0 888 0 1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5159_6
timestamp 1731220619
transform 1 0 944 0 1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5158_6
timestamp 1731220619
transform 1 0 1000 0 1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5157_6
timestamp 1731220619
transform 1 0 1040 0 1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5156_6
timestamp 1731220619
transform 1 0 912 0 -1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5155_6
timestamp 1731220619
transform 1 0 960 0 -1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5154_6
timestamp 1731220619
transform 1 0 1000 0 -1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5153_6
timestamp 1731220619
transform 1 0 1040 0 -1 1980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5152_6
timestamp 1731220619
transform 1 0 1152 0 -1 1944
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5151_6
timestamp 1731220619
transform 1 0 1216 0 -1 1944
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5150_6
timestamp 1731220619
transform 1 0 1152 0 1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5149_6
timestamp 1731220619
transform 1 0 1192 0 1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5148_6
timestamp 1731220619
transform 1 0 1256 0 1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5147_6
timestamp 1731220619
transform 1 0 1296 0 -1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5146_6
timestamp 1731220619
transform 1 0 1224 0 -1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5145_6
timestamp 1731220619
transform 1 0 1152 0 -1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5144_6
timestamp 1731220619
transform 1 0 1184 0 1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5143_6
timestamp 1731220619
transform 1 0 1248 0 1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5142_6
timestamp 1731220619
transform 1 0 1312 0 1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5141_6
timestamp 1731220619
transform 1 0 1336 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5140_6
timestamp 1731220619
transform 1 0 1288 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5139_6
timestamp 1731220619
transform 1 0 1240 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5138_6
timestamp 1731220619
transform 1 0 1256 0 1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5137_6
timestamp 1731220619
transform 1 0 1296 0 1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5136_6
timestamp 1731220619
transform 1 0 1336 0 1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5135_6
timestamp 1731220619
transform 1 0 1384 0 1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5134_6
timestamp 1731220619
transform 1 0 1440 0 1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5133_6
timestamp 1731220619
transform 1 0 1496 0 1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5132_6
timestamp 1731220619
transform 1 0 1520 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5131_6
timestamp 1731220619
transform 1 0 1456 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5130_6
timestamp 1731220619
transform 1 0 1392 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5129_6
timestamp 1731220619
transform 1 0 1376 0 1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5128_6
timestamp 1731220619
transform 1 0 1448 0 1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5127_6
timestamp 1731220619
transform 1 0 1520 0 1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5126_6
timestamp 1731220619
transform 1 0 1544 0 -1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5125_6
timestamp 1731220619
transform 1 0 1456 0 -1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5124_6
timestamp 1731220619
transform 1 0 1376 0 -1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5123_6
timestamp 1731220619
transform 1 0 1320 0 1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5122_6
timestamp 1731220619
transform 1 0 1384 0 1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5121_6
timestamp 1731220619
transform 1 0 1440 0 1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5120_6
timestamp 1731220619
transform 1 0 1456 0 -1 1944
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5119_6
timestamp 1731220619
transform 1 0 1376 0 -1 1944
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5118_6
timestamp 1731220619
transform 1 0 1296 0 -1 1944
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5117_6
timestamp 1731220619
transform 1 0 1296 0 1 1948
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5116_6
timestamp 1731220619
transform 1 0 1376 0 1 1948
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5115_6
timestamp 1731220619
transform 1 0 1456 0 1 1948
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5114_6
timestamp 1731220619
transform 1 0 1536 0 1 1948
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5113_6
timestamp 1731220619
transform 1 0 1576 0 -1 2052
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5112_6
timestamp 1731220619
transform 1 0 1480 0 -1 2052
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5111_6
timestamp 1731220619
transform 1 0 1392 0 -1 2052
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5110_6
timestamp 1731220619
transform 1 0 1304 0 -1 2052
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5109_6
timestamp 1731220619
transform 1 0 1232 0 -1 2052
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5108_6
timestamp 1731220619
transform 1 0 1176 0 -1 2052
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5107_6
timestamp 1731220619
transform 1 0 1216 0 1 2052
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5106_6
timestamp 1731220619
transform 1 0 1272 0 1 2052
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5105_6
timestamp 1731220619
transform 1 0 1336 0 1 2052
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5104_6
timestamp 1731220619
transform 1 0 1416 0 1 2052
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5103_6
timestamp 1731220619
transform 1 0 1496 0 1 2052
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5102_6
timestamp 1731220619
transform 1 0 1576 0 1 2052
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5101_6
timestamp 1731220619
transform 1 0 1280 0 -1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5100_6
timestamp 1731220619
transform 1 0 1320 0 -1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_599_6
timestamp 1731220619
transform 1 0 1360 0 -1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_598_6
timestamp 1731220619
transform 1 0 1408 0 -1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_597_6
timestamp 1731220619
transform 1 0 1456 0 -1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_596_6
timestamp 1731220619
transform 1 0 1512 0 -1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_595_6
timestamp 1731220619
transform 1 0 1568 0 -1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_594_6
timestamp 1731220619
transform 1 0 1336 0 1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_593_6
timestamp 1731220619
transform 1 0 1376 0 1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_592_6
timestamp 1731220619
transform 1 0 1416 0 1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_591_6
timestamp 1731220619
transform 1 0 1456 0 1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_590_6
timestamp 1731220619
transform 1 0 1496 0 1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_589_6
timestamp 1731220619
transform 1 0 1536 0 1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_588_6
timestamp 1731220619
transform 1 0 1576 0 1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_587_6
timestamp 1731220619
transform 1 0 1616 0 1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_586_6
timestamp 1731220619
transform 1 0 1656 0 1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_585_6
timestamp 1731220619
transform 1 0 1696 0 1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_584_6
timestamp 1731220619
transform 1 0 1736 0 1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_583_6
timestamp 1731220619
transform 1 0 1776 0 1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_582_6
timestamp 1731220619
transform 1 0 1816 0 1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_581_6
timestamp 1731220619
transform 1 0 1616 0 -1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_580_6
timestamp 1731220619
transform 1 0 1664 0 -1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_579_6
timestamp 1731220619
transform 1 0 1712 0 -1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_578_6
timestamp 1731220619
transform 1 0 1768 0 -1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_577_6
timestamp 1731220619
transform 1 0 1824 0 -1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_576_6
timestamp 1731220619
transform 1 0 1880 0 -1 2160
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_575_6
timestamp 1731220619
transform 1 0 1656 0 1 2052
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_574_6
timestamp 1731220619
transform 1 0 1736 0 1 2052
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_573_6
timestamp 1731220619
transform 1 0 1824 0 1 2052
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_572_6
timestamp 1731220619
transform 1 0 1912 0 1 2052
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_571_6
timestamp 1731220619
transform 1 0 2000 0 1 2052
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_570_6
timestamp 1731220619
transform 1 0 2000 0 -1 2052
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_569_6
timestamp 1731220619
transform 1 0 1912 0 -1 2052
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_568_6
timestamp 1731220619
transform 1 0 1832 0 -1 2052
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_567_6
timestamp 1731220619
transform 1 0 1664 0 -1 2052
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_566_6
timestamp 1731220619
transform 1 0 1752 0 -1 2052
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_565_6
timestamp 1731220619
transform 1 0 1808 0 1 1948
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_564_6
timestamp 1731220619
transform 1 0 1872 0 1 1948
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_563_6
timestamp 1731220619
transform 1 0 1944 0 1 1948
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_562_6
timestamp 1731220619
transform 1 0 1608 0 1 1948
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_561_6
timestamp 1731220619
transform 1 0 1680 0 1 1948
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_560_6
timestamp 1731220619
transform 1 0 1744 0 1 1948
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_559_6
timestamp 1731220619
transform 1 0 1776 0 -1 1944
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_558_6
timestamp 1731220619
transform 1 0 1872 0 -1 1944
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_557_6
timestamp 1731220619
transform 1 0 1976 0 -1 1944
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_556_6
timestamp 1731220619
transform 1 0 1528 0 -1 1944
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_555_6
timestamp 1731220619
transform 1 0 1608 0 -1 1944
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_554_6
timestamp 1731220619
transform 1 0 1688 0 -1 1944
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_553_6
timestamp 1731220619
transform 1 0 1704 0 1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_552_6
timestamp 1731220619
transform 1 0 1792 0 1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_551_6
timestamp 1731220619
transform 1 0 1888 0 1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_550_6
timestamp 1731220619
transform 1 0 1496 0 1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_549_6
timestamp 1731220619
transform 1 0 1552 0 1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_548_6
timestamp 1731220619
transform 1 0 1624 0 1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_547_6
timestamp 1731220619
transform 1 0 1640 0 -1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_546_6
timestamp 1731220619
transform 1 0 1744 0 -1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_545_6
timestamp 1731220619
transform 1 0 1680 0 1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_544_6
timestamp 1731220619
transform 1 0 1600 0 1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_543_6
timestamp 1731220619
transform 1 0 1664 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_542_6
timestamp 1731220619
transform 1 0 1592 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_541_6
timestamp 1731220619
transform 1 0 1560 0 1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_540_6
timestamp 1731220619
transform 1 0 1624 0 1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_539_6
timestamp 1731220619
transform 1 0 1616 0 -1 1612
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_538_6
timestamp 1731220619
transform 1 0 1456 0 -1 1612
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_537_6
timestamp 1731220619
transform 1 0 1536 0 -1 1612
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_536_6
timestamp 1731220619
transform 1 0 1552 0 1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_535_6
timestamp 1731220619
transform 1 0 1640 0 1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_534_6
timestamp 1731220619
transform 1 0 1728 0 1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_533_6
timestamp 1731220619
transform 1 0 1792 0 -1 1612
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_532_6
timestamp 1731220619
transform 1 0 1880 0 -1 1612
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_531_6
timestamp 1731220619
transform 1 0 1704 0 -1 1612
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_530_6
timestamp 1731220619
transform 1 0 1688 0 1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_529_6
timestamp 1731220619
transform 1 0 1752 0 1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_528_6
timestamp 1731220619
transform 1 0 1824 0 1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_527_6
timestamp 1731220619
transform 1 0 1904 0 1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_526_6
timestamp 1731220619
transform 1 0 1872 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_525_6
timestamp 1731220619
transform 1 0 1800 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_524_6
timestamp 1731220619
transform 1 0 1736 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_523_6
timestamp 1731220619
transform 1 0 1760 0 1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_522_6
timestamp 1731220619
transform 1 0 1840 0 1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_521_6
timestamp 1731220619
transform 1 0 1920 0 1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_520_6
timestamp 1731220619
transform 1 0 1848 0 -1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_519_6
timestamp 1731220619
transform 1 0 1960 0 -1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_518_6
timestamp 1731220619
transform 1 0 2000 0 1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_517_6
timestamp 1731220619
transform 1 0 1944 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_516_6
timestamp 1731220619
transform 1 0 1992 0 1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_515_6
timestamp 1731220619
transform 1 0 1976 0 -1 1612
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_514_6
timestamp 1731220619
transform 1 0 1912 0 -1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_513_6
timestamp 1731220619
transform 1 0 2064 0 1 1508
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_512_6
timestamp 1731220619
transform 1 0 2064 0 -1 1612
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_511_6
timestamp 1731220619
transform 1 0 2064 0 1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_510_6
timestamp 1731220619
transform 1 0 2016 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_59_6
timestamp 1731220619
transform 1 0 2064 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_58_6
timestamp 1731220619
transform 1 0 2064 0 1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_57_6
timestamp 1731220619
transform 1 0 2064 0 -1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_56_6
timestamp 1731220619
transform 1 0 1984 0 1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_55_6
timestamp 1731220619
transform 1 0 2064 0 1 1836
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_54_6
timestamp 1731220619
transform 1 0 2064 0 -1 1944
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_53_6
timestamp 1731220619
transform 1 0 2016 0 1 1948
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_52_6
timestamp 1731220619
transform 1 0 2064 0 1 1948
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_51_6
timestamp 1731220619
transform 1 0 2064 0 -1 2052
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_50_6
timestamp 1731220619
transform 1 0 2064 0 1 2052
box 4 6 36 48
<< end >>
