magic
tech sky130l
timestamp 1731220323
<< m2 >>
rect 110 3484 116 3485
rect 1766 3484 1772 3485
rect 110 3480 111 3484
rect 115 3480 116 3484
rect 110 3479 116 3480
rect 134 3483 140 3484
rect 134 3479 135 3483
rect 139 3479 140 3483
rect 134 3478 140 3479
rect 270 3483 276 3484
rect 270 3479 271 3483
rect 275 3479 276 3483
rect 270 3478 276 3479
rect 438 3483 444 3484
rect 438 3479 439 3483
rect 443 3479 444 3483
rect 438 3478 444 3479
rect 614 3483 620 3484
rect 614 3479 615 3483
rect 619 3479 620 3483
rect 614 3478 620 3479
rect 790 3483 796 3484
rect 790 3479 791 3483
rect 795 3479 796 3483
rect 790 3478 796 3479
rect 958 3483 964 3484
rect 958 3479 959 3483
rect 963 3479 964 3483
rect 958 3478 964 3479
rect 1118 3483 1124 3484
rect 1118 3479 1119 3483
rect 1123 3479 1124 3483
rect 1118 3478 1124 3479
rect 1262 3483 1268 3484
rect 1262 3479 1263 3483
rect 1267 3479 1268 3483
rect 1262 3478 1268 3479
rect 1406 3483 1412 3484
rect 1406 3479 1407 3483
rect 1411 3479 1412 3483
rect 1406 3478 1412 3479
rect 1550 3483 1556 3484
rect 1550 3479 1551 3483
rect 1555 3479 1556 3483
rect 1550 3478 1556 3479
rect 1670 3483 1676 3484
rect 1670 3479 1671 3483
rect 1675 3479 1676 3483
rect 1766 3480 1767 3484
rect 1771 3480 1772 3484
rect 1766 3479 1772 3480
rect 1670 3478 1676 3479
rect 1806 3472 1812 3473
rect 3462 3472 3468 3473
rect 1806 3468 1807 3472
rect 1811 3468 1812 3472
rect 110 3467 116 3468
rect 110 3463 111 3467
rect 115 3463 116 3467
rect 1766 3467 1772 3468
rect 1806 3467 1812 3468
rect 1830 3471 1836 3472
rect 1830 3467 1831 3471
rect 1835 3467 1836 3471
rect 110 3462 116 3463
rect 134 3464 140 3465
rect 134 3460 135 3464
rect 139 3460 140 3464
rect 134 3459 140 3460
rect 270 3464 276 3465
rect 270 3460 271 3464
rect 275 3460 276 3464
rect 270 3459 276 3460
rect 438 3464 444 3465
rect 438 3460 439 3464
rect 443 3460 444 3464
rect 438 3459 444 3460
rect 614 3464 620 3465
rect 614 3460 615 3464
rect 619 3460 620 3464
rect 614 3459 620 3460
rect 790 3464 796 3465
rect 790 3460 791 3464
rect 795 3460 796 3464
rect 790 3459 796 3460
rect 958 3464 964 3465
rect 958 3460 959 3464
rect 963 3460 964 3464
rect 958 3459 964 3460
rect 1118 3464 1124 3465
rect 1118 3460 1119 3464
rect 1123 3460 1124 3464
rect 1118 3459 1124 3460
rect 1262 3464 1268 3465
rect 1262 3460 1263 3464
rect 1267 3460 1268 3464
rect 1262 3459 1268 3460
rect 1406 3464 1412 3465
rect 1406 3460 1407 3464
rect 1411 3460 1412 3464
rect 1406 3459 1412 3460
rect 1550 3464 1556 3465
rect 1550 3460 1551 3464
rect 1555 3460 1556 3464
rect 1550 3459 1556 3460
rect 1670 3464 1676 3465
rect 1670 3460 1671 3464
rect 1675 3460 1676 3464
rect 1766 3463 1767 3467
rect 1771 3463 1772 3467
rect 1830 3466 1836 3467
rect 1974 3471 1980 3472
rect 1974 3467 1975 3471
rect 1979 3467 1980 3471
rect 1974 3466 1980 3467
rect 2142 3471 2148 3472
rect 2142 3467 2143 3471
rect 2147 3467 2148 3471
rect 2142 3466 2148 3467
rect 2310 3471 2316 3472
rect 2310 3467 2311 3471
rect 2315 3467 2316 3471
rect 2310 3466 2316 3467
rect 2478 3471 2484 3472
rect 2478 3467 2479 3471
rect 2483 3467 2484 3471
rect 2478 3466 2484 3467
rect 2638 3471 2644 3472
rect 2638 3467 2639 3471
rect 2643 3467 2644 3471
rect 2638 3466 2644 3467
rect 2798 3471 2804 3472
rect 2798 3467 2799 3471
rect 2803 3467 2804 3471
rect 2798 3466 2804 3467
rect 2966 3471 2972 3472
rect 2966 3467 2967 3471
rect 2971 3467 2972 3471
rect 3462 3468 3463 3472
rect 3467 3468 3468 3472
rect 3462 3467 3468 3468
rect 2966 3466 2972 3467
rect 1766 3462 1772 3463
rect 1670 3459 1676 3460
rect 1806 3455 1812 3456
rect 1806 3451 1807 3455
rect 1811 3451 1812 3455
rect 3462 3455 3468 3456
rect 1806 3450 1812 3451
rect 1830 3452 1836 3453
rect 1830 3448 1831 3452
rect 1835 3448 1836 3452
rect 1830 3447 1836 3448
rect 1974 3452 1980 3453
rect 1974 3448 1975 3452
rect 1979 3448 1980 3452
rect 1974 3447 1980 3448
rect 2142 3452 2148 3453
rect 2142 3448 2143 3452
rect 2147 3448 2148 3452
rect 2142 3447 2148 3448
rect 2310 3452 2316 3453
rect 2310 3448 2311 3452
rect 2315 3448 2316 3452
rect 2310 3447 2316 3448
rect 2478 3452 2484 3453
rect 2478 3448 2479 3452
rect 2483 3448 2484 3452
rect 2478 3447 2484 3448
rect 2638 3452 2644 3453
rect 2638 3448 2639 3452
rect 2643 3448 2644 3452
rect 2638 3447 2644 3448
rect 2798 3452 2804 3453
rect 2798 3448 2799 3452
rect 2803 3448 2804 3452
rect 2798 3447 2804 3448
rect 2966 3452 2972 3453
rect 2966 3448 2967 3452
rect 2971 3448 2972 3452
rect 3462 3451 3463 3455
rect 3467 3451 3468 3455
rect 3462 3450 3468 3451
rect 2966 3447 2972 3448
rect 134 3416 140 3417
rect 110 3413 116 3414
rect 110 3409 111 3413
rect 115 3409 116 3413
rect 134 3412 135 3416
rect 139 3412 140 3416
rect 134 3411 140 3412
rect 254 3416 260 3417
rect 254 3412 255 3416
rect 259 3412 260 3416
rect 254 3411 260 3412
rect 414 3416 420 3417
rect 414 3412 415 3416
rect 419 3412 420 3416
rect 414 3411 420 3412
rect 574 3416 580 3417
rect 574 3412 575 3416
rect 579 3412 580 3416
rect 574 3411 580 3412
rect 734 3416 740 3417
rect 734 3412 735 3416
rect 739 3412 740 3416
rect 734 3411 740 3412
rect 894 3416 900 3417
rect 894 3412 895 3416
rect 899 3412 900 3416
rect 894 3411 900 3412
rect 1062 3416 1068 3417
rect 1062 3412 1063 3416
rect 1067 3412 1068 3416
rect 1062 3411 1068 3412
rect 1230 3416 1236 3417
rect 1230 3412 1231 3416
rect 1235 3412 1236 3416
rect 1230 3411 1236 3412
rect 1398 3416 1404 3417
rect 1398 3412 1399 3416
rect 1403 3412 1404 3416
rect 1398 3411 1404 3412
rect 1766 3413 1772 3414
rect 110 3408 116 3409
rect 1766 3409 1767 3413
rect 1771 3409 1772 3413
rect 1766 3408 1772 3409
rect 2030 3408 2036 3409
rect 1806 3405 1812 3406
rect 1806 3401 1807 3405
rect 1811 3401 1812 3405
rect 2030 3404 2031 3408
rect 2035 3404 2036 3408
rect 2030 3403 2036 3404
rect 2150 3408 2156 3409
rect 2150 3404 2151 3408
rect 2155 3404 2156 3408
rect 2150 3403 2156 3404
rect 2270 3408 2276 3409
rect 2270 3404 2271 3408
rect 2275 3404 2276 3408
rect 2270 3403 2276 3404
rect 2390 3408 2396 3409
rect 2390 3404 2391 3408
rect 2395 3404 2396 3408
rect 2390 3403 2396 3404
rect 2510 3408 2516 3409
rect 2510 3404 2511 3408
rect 2515 3404 2516 3408
rect 2510 3403 2516 3404
rect 2622 3408 2628 3409
rect 2622 3404 2623 3408
rect 2627 3404 2628 3408
rect 2622 3403 2628 3404
rect 2726 3408 2732 3409
rect 2726 3404 2727 3408
rect 2731 3404 2732 3408
rect 2726 3403 2732 3404
rect 2830 3408 2836 3409
rect 2830 3404 2831 3408
rect 2835 3404 2836 3408
rect 2830 3403 2836 3404
rect 2934 3408 2940 3409
rect 2934 3404 2935 3408
rect 2939 3404 2940 3408
rect 2934 3403 2940 3404
rect 3038 3408 3044 3409
rect 3038 3404 3039 3408
rect 3043 3404 3044 3408
rect 3038 3403 3044 3404
rect 3150 3408 3156 3409
rect 3150 3404 3151 3408
rect 3155 3404 3156 3408
rect 3150 3403 3156 3404
rect 3462 3405 3468 3406
rect 1806 3400 1812 3401
rect 3462 3401 3463 3405
rect 3467 3401 3468 3405
rect 3462 3400 3468 3401
rect 134 3397 140 3398
rect 110 3396 116 3397
rect 110 3392 111 3396
rect 115 3392 116 3396
rect 134 3393 135 3397
rect 139 3393 140 3397
rect 134 3392 140 3393
rect 254 3397 260 3398
rect 254 3393 255 3397
rect 259 3393 260 3397
rect 254 3392 260 3393
rect 414 3397 420 3398
rect 414 3393 415 3397
rect 419 3393 420 3397
rect 414 3392 420 3393
rect 574 3397 580 3398
rect 574 3393 575 3397
rect 579 3393 580 3397
rect 574 3392 580 3393
rect 734 3397 740 3398
rect 734 3393 735 3397
rect 739 3393 740 3397
rect 734 3392 740 3393
rect 894 3397 900 3398
rect 894 3393 895 3397
rect 899 3393 900 3397
rect 894 3392 900 3393
rect 1062 3397 1068 3398
rect 1062 3393 1063 3397
rect 1067 3393 1068 3397
rect 1062 3392 1068 3393
rect 1230 3397 1236 3398
rect 1230 3393 1231 3397
rect 1235 3393 1236 3397
rect 1230 3392 1236 3393
rect 1398 3397 1404 3398
rect 1398 3393 1399 3397
rect 1403 3393 1404 3397
rect 1398 3392 1404 3393
rect 1766 3396 1772 3397
rect 1766 3392 1767 3396
rect 1771 3392 1772 3396
rect 110 3391 116 3392
rect 1766 3391 1772 3392
rect 2030 3389 2036 3390
rect 1806 3388 1812 3389
rect 1806 3384 1807 3388
rect 1811 3384 1812 3388
rect 2030 3385 2031 3389
rect 2035 3385 2036 3389
rect 2030 3384 2036 3385
rect 2150 3389 2156 3390
rect 2150 3385 2151 3389
rect 2155 3385 2156 3389
rect 2150 3384 2156 3385
rect 2270 3389 2276 3390
rect 2270 3385 2271 3389
rect 2275 3385 2276 3389
rect 2270 3384 2276 3385
rect 2390 3389 2396 3390
rect 2390 3385 2391 3389
rect 2395 3385 2396 3389
rect 2390 3384 2396 3385
rect 2510 3389 2516 3390
rect 2510 3385 2511 3389
rect 2515 3385 2516 3389
rect 2510 3384 2516 3385
rect 2622 3389 2628 3390
rect 2622 3385 2623 3389
rect 2627 3385 2628 3389
rect 2622 3384 2628 3385
rect 2726 3389 2732 3390
rect 2726 3385 2727 3389
rect 2731 3385 2732 3389
rect 2726 3384 2732 3385
rect 2830 3389 2836 3390
rect 2830 3385 2831 3389
rect 2835 3385 2836 3389
rect 2830 3384 2836 3385
rect 2934 3389 2940 3390
rect 2934 3385 2935 3389
rect 2939 3385 2940 3389
rect 2934 3384 2940 3385
rect 3038 3389 3044 3390
rect 3038 3385 3039 3389
rect 3043 3385 3044 3389
rect 3038 3384 3044 3385
rect 3150 3389 3156 3390
rect 3150 3385 3151 3389
rect 3155 3385 3156 3389
rect 3150 3384 3156 3385
rect 3462 3388 3468 3389
rect 3462 3384 3463 3388
rect 3467 3384 3468 3388
rect 1806 3383 1812 3384
rect 3462 3383 3468 3384
rect 110 3344 116 3345
rect 1766 3344 1772 3345
rect 110 3340 111 3344
rect 115 3340 116 3344
rect 110 3339 116 3340
rect 134 3343 140 3344
rect 134 3339 135 3343
rect 139 3339 140 3343
rect 134 3338 140 3339
rect 326 3343 332 3344
rect 326 3339 327 3343
rect 331 3339 332 3343
rect 326 3338 332 3339
rect 534 3343 540 3344
rect 534 3339 535 3343
rect 539 3339 540 3343
rect 534 3338 540 3339
rect 742 3343 748 3344
rect 742 3339 743 3343
rect 747 3339 748 3343
rect 742 3338 748 3339
rect 934 3343 940 3344
rect 934 3339 935 3343
rect 939 3339 940 3343
rect 934 3338 940 3339
rect 1118 3343 1124 3344
rect 1118 3339 1119 3343
rect 1123 3339 1124 3343
rect 1118 3338 1124 3339
rect 1294 3343 1300 3344
rect 1294 3339 1295 3343
rect 1299 3339 1300 3343
rect 1294 3338 1300 3339
rect 1462 3343 1468 3344
rect 1462 3339 1463 3343
rect 1467 3339 1468 3343
rect 1462 3338 1468 3339
rect 1638 3343 1644 3344
rect 1638 3339 1639 3343
rect 1643 3339 1644 3343
rect 1766 3340 1767 3344
rect 1771 3340 1772 3344
rect 1766 3339 1772 3340
rect 1806 3340 1812 3341
rect 3462 3340 3468 3341
rect 1638 3338 1644 3339
rect 1806 3336 1807 3340
rect 1811 3336 1812 3340
rect 1806 3335 1812 3336
rect 2158 3339 2164 3340
rect 2158 3335 2159 3339
rect 2163 3335 2164 3339
rect 2158 3334 2164 3335
rect 2294 3339 2300 3340
rect 2294 3335 2295 3339
rect 2299 3335 2300 3339
rect 2294 3334 2300 3335
rect 2430 3339 2436 3340
rect 2430 3335 2431 3339
rect 2435 3335 2436 3339
rect 2430 3334 2436 3335
rect 2566 3339 2572 3340
rect 2566 3335 2567 3339
rect 2571 3335 2572 3339
rect 2566 3334 2572 3335
rect 2702 3339 2708 3340
rect 2702 3335 2703 3339
rect 2707 3335 2708 3339
rect 2702 3334 2708 3335
rect 2838 3339 2844 3340
rect 2838 3335 2839 3339
rect 2843 3335 2844 3339
rect 2838 3334 2844 3335
rect 2974 3339 2980 3340
rect 2974 3335 2975 3339
rect 2979 3335 2980 3339
rect 2974 3334 2980 3335
rect 3118 3339 3124 3340
rect 3118 3335 3119 3339
rect 3123 3335 3124 3339
rect 3462 3336 3463 3340
rect 3467 3336 3468 3340
rect 3462 3335 3468 3336
rect 3118 3334 3124 3335
rect 110 3327 116 3328
rect 110 3323 111 3327
rect 115 3323 116 3327
rect 1766 3327 1772 3328
rect 110 3322 116 3323
rect 134 3324 140 3325
rect 134 3320 135 3324
rect 139 3320 140 3324
rect 134 3319 140 3320
rect 326 3324 332 3325
rect 326 3320 327 3324
rect 331 3320 332 3324
rect 326 3319 332 3320
rect 534 3324 540 3325
rect 534 3320 535 3324
rect 539 3320 540 3324
rect 534 3319 540 3320
rect 742 3324 748 3325
rect 742 3320 743 3324
rect 747 3320 748 3324
rect 742 3319 748 3320
rect 934 3324 940 3325
rect 934 3320 935 3324
rect 939 3320 940 3324
rect 934 3319 940 3320
rect 1118 3324 1124 3325
rect 1118 3320 1119 3324
rect 1123 3320 1124 3324
rect 1118 3319 1124 3320
rect 1294 3324 1300 3325
rect 1294 3320 1295 3324
rect 1299 3320 1300 3324
rect 1294 3319 1300 3320
rect 1462 3324 1468 3325
rect 1462 3320 1463 3324
rect 1467 3320 1468 3324
rect 1462 3319 1468 3320
rect 1638 3324 1644 3325
rect 1638 3320 1639 3324
rect 1643 3320 1644 3324
rect 1766 3323 1767 3327
rect 1771 3323 1772 3327
rect 1766 3322 1772 3323
rect 1806 3323 1812 3324
rect 1638 3319 1644 3320
rect 1806 3319 1807 3323
rect 1811 3319 1812 3323
rect 3462 3323 3468 3324
rect 1806 3318 1812 3319
rect 2158 3320 2164 3321
rect 2158 3316 2159 3320
rect 2163 3316 2164 3320
rect 2158 3315 2164 3316
rect 2294 3320 2300 3321
rect 2294 3316 2295 3320
rect 2299 3316 2300 3320
rect 2294 3315 2300 3316
rect 2430 3320 2436 3321
rect 2430 3316 2431 3320
rect 2435 3316 2436 3320
rect 2430 3315 2436 3316
rect 2566 3320 2572 3321
rect 2566 3316 2567 3320
rect 2571 3316 2572 3320
rect 2566 3315 2572 3316
rect 2702 3320 2708 3321
rect 2702 3316 2703 3320
rect 2707 3316 2708 3320
rect 2702 3315 2708 3316
rect 2838 3320 2844 3321
rect 2838 3316 2839 3320
rect 2843 3316 2844 3320
rect 2838 3315 2844 3316
rect 2974 3320 2980 3321
rect 2974 3316 2975 3320
rect 2979 3316 2980 3320
rect 2974 3315 2980 3316
rect 3118 3320 3124 3321
rect 3118 3316 3119 3320
rect 3123 3316 3124 3320
rect 3462 3319 3463 3323
rect 3467 3319 3468 3323
rect 3462 3318 3468 3319
rect 3118 3315 3124 3316
rect 2086 3276 2092 3277
rect 1806 3273 1812 3274
rect 134 3272 140 3273
rect 110 3269 116 3270
rect 110 3265 111 3269
rect 115 3265 116 3269
rect 134 3268 135 3272
rect 139 3268 140 3272
rect 134 3267 140 3268
rect 278 3272 284 3273
rect 278 3268 279 3272
rect 283 3268 284 3272
rect 278 3267 284 3268
rect 462 3272 468 3273
rect 462 3268 463 3272
rect 467 3268 468 3272
rect 462 3267 468 3268
rect 646 3272 652 3273
rect 646 3268 647 3272
rect 651 3268 652 3272
rect 646 3267 652 3268
rect 830 3272 836 3273
rect 830 3268 831 3272
rect 835 3268 836 3272
rect 830 3267 836 3268
rect 1006 3272 1012 3273
rect 1006 3268 1007 3272
rect 1011 3268 1012 3272
rect 1006 3267 1012 3268
rect 1174 3272 1180 3273
rect 1174 3268 1175 3272
rect 1179 3268 1180 3272
rect 1174 3267 1180 3268
rect 1342 3272 1348 3273
rect 1342 3268 1343 3272
rect 1347 3268 1348 3272
rect 1342 3267 1348 3268
rect 1502 3272 1508 3273
rect 1502 3268 1503 3272
rect 1507 3268 1508 3272
rect 1502 3267 1508 3268
rect 1670 3272 1676 3273
rect 1670 3268 1671 3272
rect 1675 3268 1676 3272
rect 1670 3267 1676 3268
rect 1766 3269 1772 3270
rect 110 3264 116 3265
rect 1766 3265 1767 3269
rect 1771 3265 1772 3269
rect 1806 3269 1807 3273
rect 1811 3269 1812 3273
rect 2086 3272 2087 3276
rect 2091 3272 2092 3276
rect 2086 3271 2092 3272
rect 2238 3276 2244 3277
rect 2238 3272 2239 3276
rect 2243 3272 2244 3276
rect 2238 3271 2244 3272
rect 2398 3276 2404 3277
rect 2398 3272 2399 3276
rect 2403 3272 2404 3276
rect 2398 3271 2404 3272
rect 2558 3276 2564 3277
rect 2558 3272 2559 3276
rect 2563 3272 2564 3276
rect 2558 3271 2564 3272
rect 2718 3276 2724 3277
rect 2718 3272 2719 3276
rect 2723 3272 2724 3276
rect 2718 3271 2724 3272
rect 2878 3276 2884 3277
rect 2878 3272 2879 3276
rect 2883 3272 2884 3276
rect 2878 3271 2884 3272
rect 3038 3276 3044 3277
rect 3038 3272 3039 3276
rect 3043 3272 3044 3276
rect 3038 3271 3044 3272
rect 3198 3276 3204 3277
rect 3198 3272 3199 3276
rect 3203 3272 3204 3276
rect 3198 3271 3204 3272
rect 3462 3273 3468 3274
rect 1806 3268 1812 3269
rect 3462 3269 3463 3273
rect 3467 3269 3468 3273
rect 3462 3268 3468 3269
rect 1766 3264 1772 3265
rect 2086 3257 2092 3258
rect 1806 3256 1812 3257
rect 134 3253 140 3254
rect 110 3252 116 3253
rect 110 3248 111 3252
rect 115 3248 116 3252
rect 134 3249 135 3253
rect 139 3249 140 3253
rect 134 3248 140 3249
rect 278 3253 284 3254
rect 278 3249 279 3253
rect 283 3249 284 3253
rect 278 3248 284 3249
rect 462 3253 468 3254
rect 462 3249 463 3253
rect 467 3249 468 3253
rect 462 3248 468 3249
rect 646 3253 652 3254
rect 646 3249 647 3253
rect 651 3249 652 3253
rect 646 3248 652 3249
rect 830 3253 836 3254
rect 830 3249 831 3253
rect 835 3249 836 3253
rect 830 3248 836 3249
rect 1006 3253 1012 3254
rect 1006 3249 1007 3253
rect 1011 3249 1012 3253
rect 1006 3248 1012 3249
rect 1174 3253 1180 3254
rect 1174 3249 1175 3253
rect 1179 3249 1180 3253
rect 1174 3248 1180 3249
rect 1342 3253 1348 3254
rect 1342 3249 1343 3253
rect 1347 3249 1348 3253
rect 1342 3248 1348 3249
rect 1502 3253 1508 3254
rect 1502 3249 1503 3253
rect 1507 3249 1508 3253
rect 1502 3248 1508 3249
rect 1670 3253 1676 3254
rect 1670 3249 1671 3253
rect 1675 3249 1676 3253
rect 1670 3248 1676 3249
rect 1766 3252 1772 3253
rect 1766 3248 1767 3252
rect 1771 3248 1772 3252
rect 1806 3252 1807 3256
rect 1811 3252 1812 3256
rect 2086 3253 2087 3257
rect 2091 3253 2092 3257
rect 2086 3252 2092 3253
rect 2238 3257 2244 3258
rect 2238 3253 2239 3257
rect 2243 3253 2244 3257
rect 2238 3252 2244 3253
rect 2398 3257 2404 3258
rect 2398 3253 2399 3257
rect 2403 3253 2404 3257
rect 2398 3252 2404 3253
rect 2558 3257 2564 3258
rect 2558 3253 2559 3257
rect 2563 3253 2564 3257
rect 2558 3252 2564 3253
rect 2718 3257 2724 3258
rect 2718 3253 2719 3257
rect 2723 3253 2724 3257
rect 2718 3252 2724 3253
rect 2878 3257 2884 3258
rect 2878 3253 2879 3257
rect 2883 3253 2884 3257
rect 2878 3252 2884 3253
rect 3038 3257 3044 3258
rect 3038 3253 3039 3257
rect 3043 3253 3044 3257
rect 3038 3252 3044 3253
rect 3198 3257 3204 3258
rect 3198 3253 3199 3257
rect 3203 3253 3204 3257
rect 3198 3252 3204 3253
rect 3462 3256 3468 3257
rect 3462 3252 3463 3256
rect 3467 3252 3468 3256
rect 1806 3251 1812 3252
rect 3462 3251 3468 3252
rect 110 3247 116 3248
rect 1766 3247 1772 3248
rect 1806 3208 1812 3209
rect 3462 3208 3468 3209
rect 1806 3204 1807 3208
rect 1811 3204 1812 3208
rect 1806 3203 1812 3204
rect 1910 3207 1916 3208
rect 1910 3203 1911 3207
rect 1915 3203 1916 3207
rect 1910 3202 1916 3203
rect 2046 3207 2052 3208
rect 2046 3203 2047 3207
rect 2051 3203 2052 3207
rect 2046 3202 2052 3203
rect 2198 3207 2204 3208
rect 2198 3203 2199 3207
rect 2203 3203 2204 3207
rect 2198 3202 2204 3203
rect 2358 3207 2364 3208
rect 2358 3203 2359 3207
rect 2363 3203 2364 3207
rect 2358 3202 2364 3203
rect 2526 3207 2532 3208
rect 2526 3203 2527 3207
rect 2531 3203 2532 3207
rect 2526 3202 2532 3203
rect 2686 3207 2692 3208
rect 2686 3203 2687 3207
rect 2691 3203 2692 3207
rect 2686 3202 2692 3203
rect 2846 3207 2852 3208
rect 2846 3203 2847 3207
rect 2851 3203 2852 3207
rect 2846 3202 2852 3203
rect 3006 3207 3012 3208
rect 3006 3203 3007 3207
rect 3011 3203 3012 3207
rect 3006 3202 3012 3203
rect 3166 3207 3172 3208
rect 3166 3203 3167 3207
rect 3171 3203 3172 3207
rect 3166 3202 3172 3203
rect 3334 3207 3340 3208
rect 3334 3203 3335 3207
rect 3339 3203 3340 3207
rect 3462 3204 3463 3208
rect 3467 3204 3468 3208
rect 3462 3203 3468 3204
rect 3334 3202 3340 3203
rect 110 3200 116 3201
rect 1766 3200 1772 3201
rect 110 3196 111 3200
rect 115 3196 116 3200
rect 110 3195 116 3196
rect 182 3199 188 3200
rect 182 3195 183 3199
rect 187 3195 188 3199
rect 182 3194 188 3195
rect 326 3199 332 3200
rect 326 3195 327 3199
rect 331 3195 332 3199
rect 326 3194 332 3195
rect 486 3199 492 3200
rect 486 3195 487 3199
rect 491 3195 492 3199
rect 486 3194 492 3195
rect 646 3199 652 3200
rect 646 3195 647 3199
rect 651 3195 652 3199
rect 646 3194 652 3195
rect 806 3199 812 3200
rect 806 3195 807 3199
rect 811 3195 812 3199
rect 806 3194 812 3195
rect 966 3199 972 3200
rect 966 3195 967 3199
rect 971 3195 972 3199
rect 966 3194 972 3195
rect 1134 3199 1140 3200
rect 1134 3195 1135 3199
rect 1139 3195 1140 3199
rect 1134 3194 1140 3195
rect 1302 3199 1308 3200
rect 1302 3195 1303 3199
rect 1307 3195 1308 3199
rect 1302 3194 1308 3195
rect 1470 3199 1476 3200
rect 1470 3195 1471 3199
rect 1475 3195 1476 3199
rect 1766 3196 1767 3200
rect 1771 3196 1772 3200
rect 1766 3195 1772 3196
rect 1470 3194 1476 3195
rect 1806 3191 1812 3192
rect 1806 3187 1807 3191
rect 1811 3187 1812 3191
rect 3462 3191 3468 3192
rect 1806 3186 1812 3187
rect 1910 3188 1916 3189
rect 1910 3184 1911 3188
rect 1915 3184 1916 3188
rect 110 3183 116 3184
rect 110 3179 111 3183
rect 115 3179 116 3183
rect 1766 3183 1772 3184
rect 1910 3183 1916 3184
rect 2046 3188 2052 3189
rect 2046 3184 2047 3188
rect 2051 3184 2052 3188
rect 2046 3183 2052 3184
rect 2198 3188 2204 3189
rect 2198 3184 2199 3188
rect 2203 3184 2204 3188
rect 2198 3183 2204 3184
rect 2358 3188 2364 3189
rect 2358 3184 2359 3188
rect 2363 3184 2364 3188
rect 2358 3183 2364 3184
rect 2526 3188 2532 3189
rect 2526 3184 2527 3188
rect 2531 3184 2532 3188
rect 2526 3183 2532 3184
rect 2686 3188 2692 3189
rect 2686 3184 2687 3188
rect 2691 3184 2692 3188
rect 2686 3183 2692 3184
rect 2846 3188 2852 3189
rect 2846 3184 2847 3188
rect 2851 3184 2852 3188
rect 2846 3183 2852 3184
rect 3006 3188 3012 3189
rect 3006 3184 3007 3188
rect 3011 3184 3012 3188
rect 3006 3183 3012 3184
rect 3166 3188 3172 3189
rect 3166 3184 3167 3188
rect 3171 3184 3172 3188
rect 3166 3183 3172 3184
rect 3334 3188 3340 3189
rect 3334 3184 3335 3188
rect 3339 3184 3340 3188
rect 3462 3187 3463 3191
rect 3467 3187 3468 3191
rect 3462 3186 3468 3187
rect 3334 3183 3340 3184
rect 110 3178 116 3179
rect 182 3180 188 3181
rect 182 3176 183 3180
rect 187 3176 188 3180
rect 182 3175 188 3176
rect 326 3180 332 3181
rect 326 3176 327 3180
rect 331 3176 332 3180
rect 326 3175 332 3176
rect 486 3180 492 3181
rect 486 3176 487 3180
rect 491 3176 492 3180
rect 486 3175 492 3176
rect 646 3180 652 3181
rect 646 3176 647 3180
rect 651 3176 652 3180
rect 646 3175 652 3176
rect 806 3180 812 3181
rect 806 3176 807 3180
rect 811 3176 812 3180
rect 806 3175 812 3176
rect 966 3180 972 3181
rect 966 3176 967 3180
rect 971 3176 972 3180
rect 966 3175 972 3176
rect 1134 3180 1140 3181
rect 1134 3176 1135 3180
rect 1139 3176 1140 3180
rect 1134 3175 1140 3176
rect 1302 3180 1308 3181
rect 1302 3176 1303 3180
rect 1307 3176 1308 3180
rect 1302 3175 1308 3176
rect 1470 3180 1476 3181
rect 1470 3176 1471 3180
rect 1475 3176 1476 3180
rect 1766 3179 1767 3183
rect 1771 3179 1772 3183
rect 1766 3178 1772 3179
rect 1470 3175 1476 3176
rect 1830 3144 1836 3145
rect 1806 3141 1812 3142
rect 1806 3137 1807 3141
rect 1811 3137 1812 3141
rect 1830 3140 1831 3144
rect 1835 3140 1836 3144
rect 1830 3139 1836 3140
rect 2006 3144 2012 3145
rect 2006 3140 2007 3144
rect 2011 3140 2012 3144
rect 2006 3139 2012 3140
rect 2206 3144 2212 3145
rect 2206 3140 2207 3144
rect 2211 3140 2212 3144
rect 2206 3139 2212 3140
rect 2398 3144 2404 3145
rect 2398 3140 2399 3144
rect 2403 3140 2404 3144
rect 2398 3139 2404 3140
rect 2582 3144 2588 3145
rect 2582 3140 2583 3144
rect 2587 3140 2588 3144
rect 2582 3139 2588 3140
rect 2758 3144 2764 3145
rect 2758 3140 2759 3144
rect 2763 3140 2764 3144
rect 2758 3139 2764 3140
rect 2918 3144 2924 3145
rect 2918 3140 2919 3144
rect 2923 3140 2924 3144
rect 2918 3139 2924 3140
rect 3078 3144 3084 3145
rect 3078 3140 3079 3144
rect 3083 3140 3084 3144
rect 3078 3139 3084 3140
rect 3230 3144 3236 3145
rect 3230 3140 3231 3144
rect 3235 3140 3236 3144
rect 3230 3139 3236 3140
rect 3366 3144 3372 3145
rect 3366 3140 3367 3144
rect 3371 3140 3372 3144
rect 3366 3139 3372 3140
rect 3462 3141 3468 3142
rect 366 3136 372 3137
rect 110 3133 116 3134
rect 110 3129 111 3133
rect 115 3129 116 3133
rect 366 3132 367 3136
rect 371 3132 372 3136
rect 366 3131 372 3132
rect 486 3136 492 3137
rect 486 3132 487 3136
rect 491 3132 492 3136
rect 486 3131 492 3132
rect 606 3136 612 3137
rect 606 3132 607 3136
rect 611 3132 612 3136
rect 606 3131 612 3132
rect 726 3136 732 3137
rect 726 3132 727 3136
rect 731 3132 732 3136
rect 726 3131 732 3132
rect 846 3136 852 3137
rect 846 3132 847 3136
rect 851 3132 852 3136
rect 846 3131 852 3132
rect 966 3136 972 3137
rect 966 3132 967 3136
rect 971 3132 972 3136
rect 966 3131 972 3132
rect 1078 3136 1084 3137
rect 1078 3132 1079 3136
rect 1083 3132 1084 3136
rect 1078 3131 1084 3132
rect 1198 3136 1204 3137
rect 1198 3132 1199 3136
rect 1203 3132 1204 3136
rect 1198 3131 1204 3132
rect 1318 3136 1324 3137
rect 1806 3136 1812 3137
rect 3462 3137 3463 3141
rect 3467 3137 3468 3141
rect 3462 3136 3468 3137
rect 1318 3132 1319 3136
rect 1323 3132 1324 3136
rect 1318 3131 1324 3132
rect 1766 3133 1772 3134
rect 110 3128 116 3129
rect 1766 3129 1767 3133
rect 1771 3129 1772 3133
rect 1766 3128 1772 3129
rect 1830 3125 1836 3126
rect 1806 3124 1812 3125
rect 1806 3120 1807 3124
rect 1811 3120 1812 3124
rect 1830 3121 1831 3125
rect 1835 3121 1836 3125
rect 1830 3120 1836 3121
rect 2006 3125 2012 3126
rect 2006 3121 2007 3125
rect 2011 3121 2012 3125
rect 2006 3120 2012 3121
rect 2206 3125 2212 3126
rect 2206 3121 2207 3125
rect 2211 3121 2212 3125
rect 2206 3120 2212 3121
rect 2398 3125 2404 3126
rect 2398 3121 2399 3125
rect 2403 3121 2404 3125
rect 2398 3120 2404 3121
rect 2582 3125 2588 3126
rect 2582 3121 2583 3125
rect 2587 3121 2588 3125
rect 2582 3120 2588 3121
rect 2758 3125 2764 3126
rect 2758 3121 2759 3125
rect 2763 3121 2764 3125
rect 2758 3120 2764 3121
rect 2918 3125 2924 3126
rect 2918 3121 2919 3125
rect 2923 3121 2924 3125
rect 2918 3120 2924 3121
rect 3078 3125 3084 3126
rect 3078 3121 3079 3125
rect 3083 3121 3084 3125
rect 3078 3120 3084 3121
rect 3230 3125 3236 3126
rect 3230 3121 3231 3125
rect 3235 3121 3236 3125
rect 3230 3120 3236 3121
rect 3366 3125 3372 3126
rect 3366 3121 3367 3125
rect 3371 3121 3372 3125
rect 3366 3120 3372 3121
rect 3462 3124 3468 3125
rect 3462 3120 3463 3124
rect 3467 3120 3468 3124
rect 1806 3119 1812 3120
rect 3462 3119 3468 3120
rect 366 3117 372 3118
rect 110 3116 116 3117
rect 110 3112 111 3116
rect 115 3112 116 3116
rect 366 3113 367 3117
rect 371 3113 372 3117
rect 366 3112 372 3113
rect 486 3117 492 3118
rect 486 3113 487 3117
rect 491 3113 492 3117
rect 486 3112 492 3113
rect 606 3117 612 3118
rect 606 3113 607 3117
rect 611 3113 612 3117
rect 606 3112 612 3113
rect 726 3117 732 3118
rect 726 3113 727 3117
rect 731 3113 732 3117
rect 726 3112 732 3113
rect 846 3117 852 3118
rect 846 3113 847 3117
rect 851 3113 852 3117
rect 846 3112 852 3113
rect 966 3117 972 3118
rect 966 3113 967 3117
rect 971 3113 972 3117
rect 966 3112 972 3113
rect 1078 3117 1084 3118
rect 1078 3113 1079 3117
rect 1083 3113 1084 3117
rect 1078 3112 1084 3113
rect 1198 3117 1204 3118
rect 1198 3113 1199 3117
rect 1203 3113 1204 3117
rect 1198 3112 1204 3113
rect 1318 3117 1324 3118
rect 1318 3113 1319 3117
rect 1323 3113 1324 3117
rect 1318 3112 1324 3113
rect 1766 3116 1772 3117
rect 1766 3112 1767 3116
rect 1771 3112 1772 3116
rect 110 3111 116 3112
rect 1766 3111 1772 3112
rect 1806 3072 1812 3073
rect 3462 3072 3468 3073
rect 110 3068 116 3069
rect 1766 3068 1772 3069
rect 110 3064 111 3068
rect 115 3064 116 3068
rect 110 3063 116 3064
rect 438 3067 444 3068
rect 438 3063 439 3067
rect 443 3063 444 3067
rect 438 3062 444 3063
rect 526 3067 532 3068
rect 526 3063 527 3067
rect 531 3063 532 3067
rect 526 3062 532 3063
rect 614 3067 620 3068
rect 614 3063 615 3067
rect 619 3063 620 3067
rect 614 3062 620 3063
rect 702 3067 708 3068
rect 702 3063 703 3067
rect 707 3063 708 3067
rect 702 3062 708 3063
rect 790 3067 796 3068
rect 790 3063 791 3067
rect 795 3063 796 3067
rect 790 3062 796 3063
rect 878 3067 884 3068
rect 878 3063 879 3067
rect 883 3063 884 3067
rect 878 3062 884 3063
rect 966 3067 972 3068
rect 966 3063 967 3067
rect 971 3063 972 3067
rect 966 3062 972 3063
rect 1054 3067 1060 3068
rect 1054 3063 1055 3067
rect 1059 3063 1060 3067
rect 1054 3062 1060 3063
rect 1142 3067 1148 3068
rect 1142 3063 1143 3067
rect 1147 3063 1148 3067
rect 1766 3064 1767 3068
rect 1771 3064 1772 3068
rect 1806 3068 1807 3072
rect 1811 3068 1812 3072
rect 1806 3067 1812 3068
rect 1830 3071 1836 3072
rect 1830 3067 1831 3071
rect 1835 3067 1836 3071
rect 1830 3066 1836 3067
rect 1958 3071 1964 3072
rect 1958 3067 1959 3071
rect 1963 3067 1964 3071
rect 1958 3066 1964 3067
rect 2118 3071 2124 3072
rect 2118 3067 2119 3071
rect 2123 3067 2124 3071
rect 2118 3066 2124 3067
rect 2294 3071 2300 3072
rect 2294 3067 2295 3071
rect 2299 3067 2300 3071
rect 2294 3066 2300 3067
rect 2486 3071 2492 3072
rect 2486 3067 2487 3071
rect 2491 3067 2492 3071
rect 2486 3066 2492 3067
rect 2694 3071 2700 3072
rect 2694 3067 2695 3071
rect 2699 3067 2700 3071
rect 2694 3066 2700 3067
rect 2918 3071 2924 3072
rect 2918 3067 2919 3071
rect 2923 3067 2924 3071
rect 2918 3066 2924 3067
rect 3150 3071 3156 3072
rect 3150 3067 3151 3071
rect 3155 3067 3156 3071
rect 3150 3066 3156 3067
rect 3366 3071 3372 3072
rect 3366 3067 3367 3071
rect 3371 3067 3372 3071
rect 3462 3068 3463 3072
rect 3467 3068 3468 3072
rect 3462 3067 3468 3068
rect 3366 3066 3372 3067
rect 1766 3063 1772 3064
rect 1142 3062 1148 3063
rect 1806 3055 1812 3056
rect 110 3051 116 3052
rect 110 3047 111 3051
rect 115 3047 116 3051
rect 1766 3051 1772 3052
rect 110 3046 116 3047
rect 438 3048 444 3049
rect 438 3044 439 3048
rect 443 3044 444 3048
rect 438 3043 444 3044
rect 526 3048 532 3049
rect 526 3044 527 3048
rect 531 3044 532 3048
rect 526 3043 532 3044
rect 614 3048 620 3049
rect 614 3044 615 3048
rect 619 3044 620 3048
rect 614 3043 620 3044
rect 702 3048 708 3049
rect 702 3044 703 3048
rect 707 3044 708 3048
rect 702 3043 708 3044
rect 790 3048 796 3049
rect 790 3044 791 3048
rect 795 3044 796 3048
rect 790 3043 796 3044
rect 878 3048 884 3049
rect 878 3044 879 3048
rect 883 3044 884 3048
rect 878 3043 884 3044
rect 966 3048 972 3049
rect 966 3044 967 3048
rect 971 3044 972 3048
rect 966 3043 972 3044
rect 1054 3048 1060 3049
rect 1054 3044 1055 3048
rect 1059 3044 1060 3048
rect 1054 3043 1060 3044
rect 1142 3048 1148 3049
rect 1142 3044 1143 3048
rect 1147 3044 1148 3048
rect 1766 3047 1767 3051
rect 1771 3047 1772 3051
rect 1806 3051 1807 3055
rect 1811 3051 1812 3055
rect 3462 3055 3468 3056
rect 1806 3050 1812 3051
rect 1830 3052 1836 3053
rect 1830 3048 1831 3052
rect 1835 3048 1836 3052
rect 1830 3047 1836 3048
rect 1958 3052 1964 3053
rect 1958 3048 1959 3052
rect 1963 3048 1964 3052
rect 1958 3047 1964 3048
rect 2118 3052 2124 3053
rect 2118 3048 2119 3052
rect 2123 3048 2124 3052
rect 2118 3047 2124 3048
rect 2294 3052 2300 3053
rect 2294 3048 2295 3052
rect 2299 3048 2300 3052
rect 2294 3047 2300 3048
rect 2486 3052 2492 3053
rect 2486 3048 2487 3052
rect 2491 3048 2492 3052
rect 2486 3047 2492 3048
rect 2694 3052 2700 3053
rect 2694 3048 2695 3052
rect 2699 3048 2700 3052
rect 2694 3047 2700 3048
rect 2918 3052 2924 3053
rect 2918 3048 2919 3052
rect 2923 3048 2924 3052
rect 2918 3047 2924 3048
rect 3150 3052 3156 3053
rect 3150 3048 3151 3052
rect 3155 3048 3156 3052
rect 3150 3047 3156 3048
rect 3366 3052 3372 3053
rect 3366 3048 3367 3052
rect 3371 3048 3372 3052
rect 3462 3051 3463 3055
rect 3467 3051 3468 3055
rect 3462 3050 3468 3051
rect 3366 3047 3372 3048
rect 1766 3046 1772 3047
rect 1142 3043 1148 3044
rect 502 2996 508 2997
rect 110 2993 116 2994
rect 110 2989 111 2993
rect 115 2989 116 2993
rect 502 2992 503 2996
rect 507 2992 508 2996
rect 502 2991 508 2992
rect 590 2996 596 2997
rect 590 2992 591 2996
rect 595 2992 596 2996
rect 590 2991 596 2992
rect 678 2996 684 2997
rect 678 2992 679 2996
rect 683 2992 684 2996
rect 678 2991 684 2992
rect 766 2996 772 2997
rect 766 2992 767 2996
rect 771 2992 772 2996
rect 766 2991 772 2992
rect 854 2996 860 2997
rect 854 2992 855 2996
rect 859 2992 860 2996
rect 854 2991 860 2992
rect 942 2996 948 2997
rect 942 2992 943 2996
rect 947 2992 948 2996
rect 942 2991 948 2992
rect 1030 2996 1036 2997
rect 1030 2992 1031 2996
rect 1035 2992 1036 2996
rect 1030 2991 1036 2992
rect 1118 2996 1124 2997
rect 1118 2992 1119 2996
rect 1123 2992 1124 2996
rect 1118 2991 1124 2992
rect 1206 2996 1212 2997
rect 1206 2992 1207 2996
rect 1211 2992 1212 2996
rect 1206 2991 1212 2992
rect 1294 2996 1300 2997
rect 1294 2992 1295 2996
rect 1299 2992 1300 2996
rect 1294 2991 1300 2992
rect 1766 2993 1772 2994
rect 110 2988 116 2989
rect 1766 2989 1767 2993
rect 1771 2989 1772 2993
rect 1830 2992 1836 2993
rect 1766 2988 1772 2989
rect 1806 2989 1812 2990
rect 1806 2985 1807 2989
rect 1811 2985 1812 2989
rect 1830 2988 1831 2992
rect 1835 2988 1836 2992
rect 1830 2987 1836 2988
rect 1918 2992 1924 2993
rect 1918 2988 1919 2992
rect 1923 2988 1924 2992
rect 1918 2987 1924 2988
rect 2030 2992 2036 2993
rect 2030 2988 2031 2992
rect 2035 2988 2036 2992
rect 2030 2987 2036 2988
rect 2142 2992 2148 2993
rect 2142 2988 2143 2992
rect 2147 2988 2148 2992
rect 2142 2987 2148 2988
rect 2246 2992 2252 2993
rect 2246 2988 2247 2992
rect 2251 2988 2252 2992
rect 2246 2987 2252 2988
rect 2358 2992 2364 2993
rect 2358 2988 2359 2992
rect 2363 2988 2364 2992
rect 2358 2987 2364 2988
rect 2478 2992 2484 2993
rect 2478 2988 2479 2992
rect 2483 2988 2484 2992
rect 2478 2987 2484 2988
rect 2622 2992 2628 2993
rect 2622 2988 2623 2992
rect 2627 2988 2628 2992
rect 2622 2987 2628 2988
rect 2790 2992 2796 2993
rect 2790 2988 2791 2992
rect 2795 2988 2796 2992
rect 2790 2987 2796 2988
rect 2982 2992 2988 2993
rect 2982 2988 2983 2992
rect 2987 2988 2988 2992
rect 2982 2987 2988 2988
rect 3182 2992 3188 2993
rect 3182 2988 3183 2992
rect 3187 2988 3188 2992
rect 3182 2987 3188 2988
rect 3366 2992 3372 2993
rect 3366 2988 3367 2992
rect 3371 2988 3372 2992
rect 3366 2987 3372 2988
rect 3462 2989 3468 2990
rect 1806 2984 1812 2985
rect 3462 2985 3463 2989
rect 3467 2985 3468 2989
rect 3462 2984 3468 2985
rect 502 2977 508 2978
rect 110 2976 116 2977
rect 110 2972 111 2976
rect 115 2972 116 2976
rect 502 2973 503 2977
rect 507 2973 508 2977
rect 502 2972 508 2973
rect 590 2977 596 2978
rect 590 2973 591 2977
rect 595 2973 596 2977
rect 590 2972 596 2973
rect 678 2977 684 2978
rect 678 2973 679 2977
rect 683 2973 684 2977
rect 678 2972 684 2973
rect 766 2977 772 2978
rect 766 2973 767 2977
rect 771 2973 772 2977
rect 766 2972 772 2973
rect 854 2977 860 2978
rect 854 2973 855 2977
rect 859 2973 860 2977
rect 854 2972 860 2973
rect 942 2977 948 2978
rect 942 2973 943 2977
rect 947 2973 948 2977
rect 942 2972 948 2973
rect 1030 2977 1036 2978
rect 1030 2973 1031 2977
rect 1035 2973 1036 2977
rect 1030 2972 1036 2973
rect 1118 2977 1124 2978
rect 1118 2973 1119 2977
rect 1123 2973 1124 2977
rect 1118 2972 1124 2973
rect 1206 2977 1212 2978
rect 1206 2973 1207 2977
rect 1211 2973 1212 2977
rect 1206 2972 1212 2973
rect 1294 2977 1300 2978
rect 1294 2973 1295 2977
rect 1299 2973 1300 2977
rect 1294 2972 1300 2973
rect 1766 2976 1772 2977
rect 1766 2972 1767 2976
rect 1771 2972 1772 2976
rect 1830 2973 1836 2974
rect 110 2971 116 2972
rect 1766 2971 1772 2972
rect 1806 2972 1812 2973
rect 1806 2968 1807 2972
rect 1811 2968 1812 2972
rect 1830 2969 1831 2973
rect 1835 2969 1836 2973
rect 1830 2968 1836 2969
rect 1918 2973 1924 2974
rect 1918 2969 1919 2973
rect 1923 2969 1924 2973
rect 1918 2968 1924 2969
rect 2030 2973 2036 2974
rect 2030 2969 2031 2973
rect 2035 2969 2036 2973
rect 2030 2968 2036 2969
rect 2142 2973 2148 2974
rect 2142 2969 2143 2973
rect 2147 2969 2148 2973
rect 2142 2968 2148 2969
rect 2246 2973 2252 2974
rect 2246 2969 2247 2973
rect 2251 2969 2252 2973
rect 2246 2968 2252 2969
rect 2358 2973 2364 2974
rect 2358 2969 2359 2973
rect 2363 2969 2364 2973
rect 2358 2968 2364 2969
rect 2478 2973 2484 2974
rect 2478 2969 2479 2973
rect 2483 2969 2484 2973
rect 2478 2968 2484 2969
rect 2622 2973 2628 2974
rect 2622 2969 2623 2973
rect 2627 2969 2628 2973
rect 2622 2968 2628 2969
rect 2790 2973 2796 2974
rect 2790 2969 2791 2973
rect 2795 2969 2796 2973
rect 2790 2968 2796 2969
rect 2982 2973 2988 2974
rect 2982 2969 2983 2973
rect 2987 2969 2988 2973
rect 2982 2968 2988 2969
rect 3182 2973 3188 2974
rect 3182 2969 3183 2973
rect 3187 2969 3188 2973
rect 3182 2968 3188 2969
rect 3366 2973 3372 2974
rect 3366 2969 3367 2973
rect 3371 2969 3372 2973
rect 3366 2968 3372 2969
rect 3462 2972 3468 2973
rect 3462 2968 3463 2972
rect 3467 2968 3468 2972
rect 1806 2967 1812 2968
rect 3462 2967 3468 2968
rect 110 2920 116 2921
rect 1766 2920 1772 2921
rect 110 2916 111 2920
rect 115 2916 116 2920
rect 110 2915 116 2916
rect 326 2919 332 2920
rect 326 2915 327 2919
rect 331 2915 332 2919
rect 326 2914 332 2915
rect 446 2919 452 2920
rect 446 2915 447 2919
rect 451 2915 452 2919
rect 446 2914 452 2915
rect 574 2919 580 2920
rect 574 2915 575 2919
rect 579 2915 580 2919
rect 574 2914 580 2915
rect 710 2919 716 2920
rect 710 2915 711 2919
rect 715 2915 716 2919
rect 710 2914 716 2915
rect 846 2919 852 2920
rect 846 2915 847 2919
rect 851 2915 852 2919
rect 846 2914 852 2915
rect 974 2919 980 2920
rect 974 2915 975 2919
rect 979 2915 980 2919
rect 974 2914 980 2915
rect 1102 2919 1108 2920
rect 1102 2915 1103 2919
rect 1107 2915 1108 2919
rect 1102 2914 1108 2915
rect 1230 2919 1236 2920
rect 1230 2915 1231 2919
rect 1235 2915 1236 2919
rect 1230 2914 1236 2915
rect 1358 2919 1364 2920
rect 1358 2915 1359 2919
rect 1363 2915 1364 2919
rect 1358 2914 1364 2915
rect 1494 2919 1500 2920
rect 1494 2915 1495 2919
rect 1499 2915 1500 2919
rect 1766 2916 1767 2920
rect 1771 2916 1772 2920
rect 1766 2915 1772 2916
rect 1806 2916 1812 2917
rect 3462 2916 3468 2917
rect 1494 2914 1500 2915
rect 1806 2912 1807 2916
rect 1811 2912 1812 2916
rect 1806 2911 1812 2912
rect 1830 2915 1836 2916
rect 1830 2911 1831 2915
rect 1835 2911 1836 2915
rect 1830 2910 1836 2911
rect 2014 2915 2020 2916
rect 2014 2911 2015 2915
rect 2019 2911 2020 2915
rect 2014 2910 2020 2911
rect 2214 2915 2220 2916
rect 2214 2911 2215 2915
rect 2219 2911 2220 2915
rect 2214 2910 2220 2911
rect 2406 2915 2412 2916
rect 2406 2911 2407 2915
rect 2411 2911 2412 2915
rect 2406 2910 2412 2911
rect 2590 2915 2596 2916
rect 2590 2911 2591 2915
rect 2595 2911 2596 2915
rect 2590 2910 2596 2911
rect 2758 2915 2764 2916
rect 2758 2911 2759 2915
rect 2763 2911 2764 2915
rect 2758 2910 2764 2911
rect 2910 2915 2916 2916
rect 2910 2911 2911 2915
rect 2915 2911 2916 2915
rect 2910 2910 2916 2911
rect 3062 2915 3068 2916
rect 3062 2911 3063 2915
rect 3067 2911 3068 2915
rect 3062 2910 3068 2911
rect 3206 2915 3212 2916
rect 3206 2911 3207 2915
rect 3211 2911 3212 2915
rect 3206 2910 3212 2911
rect 3358 2915 3364 2916
rect 3358 2911 3359 2915
rect 3363 2911 3364 2915
rect 3462 2912 3463 2916
rect 3467 2912 3468 2916
rect 3462 2911 3468 2912
rect 3358 2910 3364 2911
rect 110 2903 116 2904
rect 110 2899 111 2903
rect 115 2899 116 2903
rect 1766 2903 1772 2904
rect 110 2898 116 2899
rect 326 2900 332 2901
rect 326 2896 327 2900
rect 331 2896 332 2900
rect 326 2895 332 2896
rect 446 2900 452 2901
rect 446 2896 447 2900
rect 451 2896 452 2900
rect 446 2895 452 2896
rect 574 2900 580 2901
rect 574 2896 575 2900
rect 579 2896 580 2900
rect 574 2895 580 2896
rect 710 2900 716 2901
rect 710 2896 711 2900
rect 715 2896 716 2900
rect 710 2895 716 2896
rect 846 2900 852 2901
rect 846 2896 847 2900
rect 851 2896 852 2900
rect 846 2895 852 2896
rect 974 2900 980 2901
rect 974 2896 975 2900
rect 979 2896 980 2900
rect 974 2895 980 2896
rect 1102 2900 1108 2901
rect 1102 2896 1103 2900
rect 1107 2896 1108 2900
rect 1102 2895 1108 2896
rect 1230 2900 1236 2901
rect 1230 2896 1231 2900
rect 1235 2896 1236 2900
rect 1230 2895 1236 2896
rect 1358 2900 1364 2901
rect 1358 2896 1359 2900
rect 1363 2896 1364 2900
rect 1358 2895 1364 2896
rect 1494 2900 1500 2901
rect 1494 2896 1495 2900
rect 1499 2896 1500 2900
rect 1766 2899 1767 2903
rect 1771 2899 1772 2903
rect 1766 2898 1772 2899
rect 1806 2899 1812 2900
rect 1494 2895 1500 2896
rect 1806 2895 1807 2899
rect 1811 2895 1812 2899
rect 3462 2899 3468 2900
rect 1806 2894 1812 2895
rect 1830 2896 1836 2897
rect 1830 2892 1831 2896
rect 1835 2892 1836 2896
rect 1830 2891 1836 2892
rect 2014 2896 2020 2897
rect 2014 2892 2015 2896
rect 2019 2892 2020 2896
rect 2014 2891 2020 2892
rect 2214 2896 2220 2897
rect 2214 2892 2215 2896
rect 2219 2892 2220 2896
rect 2214 2891 2220 2892
rect 2406 2896 2412 2897
rect 2406 2892 2407 2896
rect 2411 2892 2412 2896
rect 2406 2891 2412 2892
rect 2590 2896 2596 2897
rect 2590 2892 2591 2896
rect 2595 2892 2596 2896
rect 2590 2891 2596 2892
rect 2758 2896 2764 2897
rect 2758 2892 2759 2896
rect 2763 2892 2764 2896
rect 2758 2891 2764 2892
rect 2910 2896 2916 2897
rect 2910 2892 2911 2896
rect 2915 2892 2916 2896
rect 2910 2891 2916 2892
rect 3062 2896 3068 2897
rect 3062 2892 3063 2896
rect 3067 2892 3068 2896
rect 3062 2891 3068 2892
rect 3206 2896 3212 2897
rect 3206 2892 3207 2896
rect 3211 2892 3212 2896
rect 3206 2891 3212 2892
rect 3358 2896 3364 2897
rect 3358 2892 3359 2896
rect 3363 2892 3364 2896
rect 3462 2895 3463 2899
rect 3467 2895 3468 2899
rect 3462 2894 3468 2895
rect 3358 2891 3364 2892
rect 1830 2852 1836 2853
rect 1806 2849 1812 2850
rect 134 2848 140 2849
rect 110 2845 116 2846
rect 110 2841 111 2845
rect 115 2841 116 2845
rect 134 2844 135 2848
rect 139 2844 140 2848
rect 134 2843 140 2844
rect 254 2848 260 2849
rect 254 2844 255 2848
rect 259 2844 260 2848
rect 254 2843 260 2844
rect 414 2848 420 2849
rect 414 2844 415 2848
rect 419 2844 420 2848
rect 414 2843 420 2844
rect 574 2848 580 2849
rect 574 2844 575 2848
rect 579 2844 580 2848
rect 574 2843 580 2844
rect 734 2848 740 2849
rect 734 2844 735 2848
rect 739 2844 740 2848
rect 734 2843 740 2844
rect 894 2848 900 2849
rect 894 2844 895 2848
rect 899 2844 900 2848
rect 894 2843 900 2844
rect 1046 2848 1052 2849
rect 1046 2844 1047 2848
rect 1051 2844 1052 2848
rect 1046 2843 1052 2844
rect 1190 2848 1196 2849
rect 1190 2844 1191 2848
rect 1195 2844 1196 2848
rect 1190 2843 1196 2844
rect 1342 2848 1348 2849
rect 1342 2844 1343 2848
rect 1347 2844 1348 2848
rect 1342 2843 1348 2844
rect 1494 2848 1500 2849
rect 1494 2844 1495 2848
rect 1499 2844 1500 2848
rect 1494 2843 1500 2844
rect 1766 2845 1772 2846
rect 110 2840 116 2841
rect 1766 2841 1767 2845
rect 1771 2841 1772 2845
rect 1806 2845 1807 2849
rect 1811 2845 1812 2849
rect 1830 2848 1831 2852
rect 1835 2848 1836 2852
rect 1830 2847 1836 2848
rect 1998 2852 2004 2853
rect 1998 2848 1999 2852
rect 2003 2848 2004 2852
rect 1998 2847 2004 2848
rect 2190 2852 2196 2853
rect 2190 2848 2191 2852
rect 2195 2848 2196 2852
rect 2190 2847 2196 2848
rect 2382 2852 2388 2853
rect 2382 2848 2383 2852
rect 2387 2848 2388 2852
rect 2382 2847 2388 2848
rect 2566 2852 2572 2853
rect 2566 2848 2567 2852
rect 2571 2848 2572 2852
rect 2566 2847 2572 2848
rect 2734 2852 2740 2853
rect 2734 2848 2735 2852
rect 2739 2848 2740 2852
rect 2734 2847 2740 2848
rect 2902 2852 2908 2853
rect 2902 2848 2903 2852
rect 2907 2848 2908 2852
rect 2902 2847 2908 2848
rect 3062 2852 3068 2853
rect 3062 2848 3063 2852
rect 3067 2848 3068 2852
rect 3062 2847 3068 2848
rect 3222 2852 3228 2853
rect 3222 2848 3223 2852
rect 3227 2848 3228 2852
rect 3222 2847 3228 2848
rect 3366 2852 3372 2853
rect 3366 2848 3367 2852
rect 3371 2848 3372 2852
rect 3366 2847 3372 2848
rect 3462 2849 3468 2850
rect 1806 2844 1812 2845
rect 3462 2845 3463 2849
rect 3467 2845 3468 2849
rect 3462 2844 3468 2845
rect 1766 2840 1772 2841
rect 1830 2833 1836 2834
rect 1806 2832 1812 2833
rect 134 2829 140 2830
rect 110 2828 116 2829
rect 110 2824 111 2828
rect 115 2824 116 2828
rect 134 2825 135 2829
rect 139 2825 140 2829
rect 134 2824 140 2825
rect 254 2829 260 2830
rect 254 2825 255 2829
rect 259 2825 260 2829
rect 254 2824 260 2825
rect 414 2829 420 2830
rect 414 2825 415 2829
rect 419 2825 420 2829
rect 414 2824 420 2825
rect 574 2829 580 2830
rect 574 2825 575 2829
rect 579 2825 580 2829
rect 574 2824 580 2825
rect 734 2829 740 2830
rect 734 2825 735 2829
rect 739 2825 740 2829
rect 734 2824 740 2825
rect 894 2829 900 2830
rect 894 2825 895 2829
rect 899 2825 900 2829
rect 894 2824 900 2825
rect 1046 2829 1052 2830
rect 1046 2825 1047 2829
rect 1051 2825 1052 2829
rect 1046 2824 1052 2825
rect 1190 2829 1196 2830
rect 1190 2825 1191 2829
rect 1195 2825 1196 2829
rect 1190 2824 1196 2825
rect 1342 2829 1348 2830
rect 1342 2825 1343 2829
rect 1347 2825 1348 2829
rect 1342 2824 1348 2825
rect 1494 2829 1500 2830
rect 1494 2825 1495 2829
rect 1499 2825 1500 2829
rect 1494 2824 1500 2825
rect 1766 2828 1772 2829
rect 1766 2824 1767 2828
rect 1771 2824 1772 2828
rect 1806 2828 1807 2832
rect 1811 2828 1812 2832
rect 1830 2829 1831 2833
rect 1835 2829 1836 2833
rect 1830 2828 1836 2829
rect 1998 2833 2004 2834
rect 1998 2829 1999 2833
rect 2003 2829 2004 2833
rect 1998 2828 2004 2829
rect 2190 2833 2196 2834
rect 2190 2829 2191 2833
rect 2195 2829 2196 2833
rect 2190 2828 2196 2829
rect 2382 2833 2388 2834
rect 2382 2829 2383 2833
rect 2387 2829 2388 2833
rect 2382 2828 2388 2829
rect 2566 2833 2572 2834
rect 2566 2829 2567 2833
rect 2571 2829 2572 2833
rect 2566 2828 2572 2829
rect 2734 2833 2740 2834
rect 2734 2829 2735 2833
rect 2739 2829 2740 2833
rect 2734 2828 2740 2829
rect 2902 2833 2908 2834
rect 2902 2829 2903 2833
rect 2907 2829 2908 2833
rect 2902 2828 2908 2829
rect 3062 2833 3068 2834
rect 3062 2829 3063 2833
rect 3067 2829 3068 2833
rect 3062 2828 3068 2829
rect 3222 2833 3228 2834
rect 3222 2829 3223 2833
rect 3227 2829 3228 2833
rect 3222 2828 3228 2829
rect 3366 2833 3372 2834
rect 3366 2829 3367 2833
rect 3371 2829 3372 2833
rect 3366 2828 3372 2829
rect 3462 2832 3468 2833
rect 3462 2828 3463 2832
rect 3467 2828 3468 2832
rect 1806 2827 1812 2828
rect 3462 2827 3468 2828
rect 110 2823 116 2824
rect 1766 2823 1772 2824
rect 1806 2784 1812 2785
rect 3462 2784 3468 2785
rect 1806 2780 1807 2784
rect 1811 2780 1812 2784
rect 1806 2779 1812 2780
rect 1830 2783 1836 2784
rect 1830 2779 1831 2783
rect 1835 2779 1836 2783
rect 1830 2778 1836 2779
rect 2014 2783 2020 2784
rect 2014 2779 2015 2783
rect 2019 2779 2020 2783
rect 2014 2778 2020 2779
rect 2214 2783 2220 2784
rect 2214 2779 2215 2783
rect 2219 2779 2220 2783
rect 2214 2778 2220 2779
rect 2406 2783 2412 2784
rect 2406 2779 2407 2783
rect 2411 2779 2412 2783
rect 2406 2778 2412 2779
rect 2582 2783 2588 2784
rect 2582 2779 2583 2783
rect 2587 2779 2588 2783
rect 2582 2778 2588 2779
rect 2750 2783 2756 2784
rect 2750 2779 2751 2783
rect 2755 2779 2756 2783
rect 2750 2778 2756 2779
rect 2910 2783 2916 2784
rect 2910 2779 2911 2783
rect 2915 2779 2916 2783
rect 2910 2778 2916 2779
rect 3070 2783 3076 2784
rect 3070 2779 3071 2783
rect 3075 2779 3076 2783
rect 3070 2778 3076 2779
rect 3230 2783 3236 2784
rect 3230 2779 3231 2783
rect 3235 2779 3236 2783
rect 3230 2778 3236 2779
rect 3366 2783 3372 2784
rect 3366 2779 3367 2783
rect 3371 2779 3372 2783
rect 3462 2780 3463 2784
rect 3467 2780 3468 2784
rect 3462 2779 3468 2780
rect 3366 2778 3372 2779
rect 110 2772 116 2773
rect 1766 2772 1772 2773
rect 110 2768 111 2772
rect 115 2768 116 2772
rect 110 2767 116 2768
rect 134 2771 140 2772
rect 134 2767 135 2771
rect 139 2767 140 2771
rect 134 2766 140 2767
rect 246 2771 252 2772
rect 246 2767 247 2771
rect 251 2767 252 2771
rect 246 2766 252 2767
rect 390 2771 396 2772
rect 390 2767 391 2771
rect 395 2767 396 2771
rect 390 2766 396 2767
rect 542 2771 548 2772
rect 542 2767 543 2771
rect 547 2767 548 2771
rect 542 2766 548 2767
rect 694 2771 700 2772
rect 694 2767 695 2771
rect 699 2767 700 2771
rect 694 2766 700 2767
rect 854 2771 860 2772
rect 854 2767 855 2771
rect 859 2767 860 2771
rect 854 2766 860 2767
rect 1022 2771 1028 2772
rect 1022 2767 1023 2771
rect 1027 2767 1028 2771
rect 1022 2766 1028 2767
rect 1190 2771 1196 2772
rect 1190 2767 1191 2771
rect 1195 2767 1196 2771
rect 1190 2766 1196 2767
rect 1358 2771 1364 2772
rect 1358 2767 1359 2771
rect 1363 2767 1364 2771
rect 1358 2766 1364 2767
rect 1526 2771 1532 2772
rect 1526 2767 1527 2771
rect 1531 2767 1532 2771
rect 1526 2766 1532 2767
rect 1670 2771 1676 2772
rect 1670 2767 1671 2771
rect 1675 2767 1676 2771
rect 1766 2768 1767 2772
rect 1771 2768 1772 2772
rect 1766 2767 1772 2768
rect 1806 2767 1812 2768
rect 1670 2766 1676 2767
rect 1806 2763 1807 2767
rect 1811 2763 1812 2767
rect 3462 2767 3468 2768
rect 1806 2762 1812 2763
rect 1830 2764 1836 2765
rect 1830 2760 1831 2764
rect 1835 2760 1836 2764
rect 1830 2759 1836 2760
rect 2014 2764 2020 2765
rect 2014 2760 2015 2764
rect 2019 2760 2020 2764
rect 2014 2759 2020 2760
rect 2214 2764 2220 2765
rect 2214 2760 2215 2764
rect 2219 2760 2220 2764
rect 2214 2759 2220 2760
rect 2406 2764 2412 2765
rect 2406 2760 2407 2764
rect 2411 2760 2412 2764
rect 2406 2759 2412 2760
rect 2582 2764 2588 2765
rect 2582 2760 2583 2764
rect 2587 2760 2588 2764
rect 2582 2759 2588 2760
rect 2750 2764 2756 2765
rect 2750 2760 2751 2764
rect 2755 2760 2756 2764
rect 2750 2759 2756 2760
rect 2910 2764 2916 2765
rect 2910 2760 2911 2764
rect 2915 2760 2916 2764
rect 2910 2759 2916 2760
rect 3070 2764 3076 2765
rect 3070 2760 3071 2764
rect 3075 2760 3076 2764
rect 3070 2759 3076 2760
rect 3230 2764 3236 2765
rect 3230 2760 3231 2764
rect 3235 2760 3236 2764
rect 3230 2759 3236 2760
rect 3366 2764 3372 2765
rect 3366 2760 3367 2764
rect 3371 2760 3372 2764
rect 3462 2763 3463 2767
rect 3467 2763 3468 2767
rect 3462 2762 3468 2763
rect 3366 2759 3372 2760
rect 110 2755 116 2756
rect 110 2751 111 2755
rect 115 2751 116 2755
rect 1766 2755 1772 2756
rect 110 2750 116 2751
rect 134 2752 140 2753
rect 134 2748 135 2752
rect 139 2748 140 2752
rect 134 2747 140 2748
rect 246 2752 252 2753
rect 246 2748 247 2752
rect 251 2748 252 2752
rect 246 2747 252 2748
rect 390 2752 396 2753
rect 390 2748 391 2752
rect 395 2748 396 2752
rect 390 2747 396 2748
rect 542 2752 548 2753
rect 542 2748 543 2752
rect 547 2748 548 2752
rect 542 2747 548 2748
rect 694 2752 700 2753
rect 694 2748 695 2752
rect 699 2748 700 2752
rect 694 2747 700 2748
rect 854 2752 860 2753
rect 854 2748 855 2752
rect 859 2748 860 2752
rect 854 2747 860 2748
rect 1022 2752 1028 2753
rect 1022 2748 1023 2752
rect 1027 2748 1028 2752
rect 1022 2747 1028 2748
rect 1190 2752 1196 2753
rect 1190 2748 1191 2752
rect 1195 2748 1196 2752
rect 1190 2747 1196 2748
rect 1358 2752 1364 2753
rect 1358 2748 1359 2752
rect 1363 2748 1364 2752
rect 1358 2747 1364 2748
rect 1526 2752 1532 2753
rect 1526 2748 1527 2752
rect 1531 2748 1532 2752
rect 1526 2747 1532 2748
rect 1670 2752 1676 2753
rect 1670 2748 1671 2752
rect 1675 2748 1676 2752
rect 1766 2751 1767 2755
rect 1771 2751 1772 2755
rect 1766 2750 1772 2751
rect 1670 2747 1676 2748
rect 2038 2704 2044 2705
rect 1806 2701 1812 2702
rect 246 2700 252 2701
rect 110 2697 116 2698
rect 110 2693 111 2697
rect 115 2693 116 2697
rect 246 2696 247 2700
rect 251 2696 252 2700
rect 246 2695 252 2696
rect 358 2700 364 2701
rect 358 2696 359 2700
rect 363 2696 364 2700
rect 358 2695 364 2696
rect 478 2700 484 2701
rect 478 2696 479 2700
rect 483 2696 484 2700
rect 478 2695 484 2696
rect 614 2700 620 2701
rect 614 2696 615 2700
rect 619 2696 620 2700
rect 614 2695 620 2696
rect 758 2700 764 2701
rect 758 2696 759 2700
rect 763 2696 764 2700
rect 758 2695 764 2696
rect 910 2700 916 2701
rect 910 2696 911 2700
rect 915 2696 916 2700
rect 910 2695 916 2696
rect 1062 2700 1068 2701
rect 1062 2696 1063 2700
rect 1067 2696 1068 2700
rect 1062 2695 1068 2696
rect 1214 2700 1220 2701
rect 1214 2696 1215 2700
rect 1219 2696 1220 2700
rect 1214 2695 1220 2696
rect 1374 2700 1380 2701
rect 1374 2696 1375 2700
rect 1379 2696 1380 2700
rect 1374 2695 1380 2696
rect 1534 2700 1540 2701
rect 1534 2696 1535 2700
rect 1539 2696 1540 2700
rect 1534 2695 1540 2696
rect 1670 2700 1676 2701
rect 1670 2696 1671 2700
rect 1675 2696 1676 2700
rect 1670 2695 1676 2696
rect 1766 2697 1772 2698
rect 110 2692 116 2693
rect 1766 2693 1767 2697
rect 1771 2693 1772 2697
rect 1806 2697 1807 2701
rect 1811 2697 1812 2701
rect 2038 2700 2039 2704
rect 2043 2700 2044 2704
rect 2038 2699 2044 2700
rect 2158 2704 2164 2705
rect 2158 2700 2159 2704
rect 2163 2700 2164 2704
rect 2158 2699 2164 2700
rect 2278 2704 2284 2705
rect 2278 2700 2279 2704
rect 2283 2700 2284 2704
rect 2278 2699 2284 2700
rect 2406 2704 2412 2705
rect 2406 2700 2407 2704
rect 2411 2700 2412 2704
rect 2406 2699 2412 2700
rect 2542 2704 2548 2705
rect 2542 2700 2543 2704
rect 2547 2700 2548 2704
rect 2542 2699 2548 2700
rect 2686 2704 2692 2705
rect 2686 2700 2687 2704
rect 2691 2700 2692 2704
rect 2686 2699 2692 2700
rect 2846 2704 2852 2705
rect 2846 2700 2847 2704
rect 2851 2700 2852 2704
rect 2846 2699 2852 2700
rect 3022 2704 3028 2705
rect 3022 2700 3023 2704
rect 3027 2700 3028 2704
rect 3022 2699 3028 2700
rect 3206 2704 3212 2705
rect 3206 2700 3207 2704
rect 3211 2700 3212 2704
rect 3206 2699 3212 2700
rect 3366 2704 3372 2705
rect 3366 2700 3367 2704
rect 3371 2700 3372 2704
rect 3366 2699 3372 2700
rect 3462 2701 3468 2702
rect 1806 2696 1812 2697
rect 3462 2697 3463 2701
rect 3467 2697 3468 2701
rect 3462 2696 3468 2697
rect 1766 2692 1772 2693
rect 2038 2685 2044 2686
rect 1806 2684 1812 2685
rect 246 2681 252 2682
rect 110 2680 116 2681
rect 110 2676 111 2680
rect 115 2676 116 2680
rect 246 2677 247 2681
rect 251 2677 252 2681
rect 246 2676 252 2677
rect 358 2681 364 2682
rect 358 2677 359 2681
rect 363 2677 364 2681
rect 358 2676 364 2677
rect 478 2681 484 2682
rect 478 2677 479 2681
rect 483 2677 484 2681
rect 478 2676 484 2677
rect 614 2681 620 2682
rect 614 2677 615 2681
rect 619 2677 620 2681
rect 614 2676 620 2677
rect 758 2681 764 2682
rect 758 2677 759 2681
rect 763 2677 764 2681
rect 758 2676 764 2677
rect 910 2681 916 2682
rect 910 2677 911 2681
rect 915 2677 916 2681
rect 910 2676 916 2677
rect 1062 2681 1068 2682
rect 1062 2677 1063 2681
rect 1067 2677 1068 2681
rect 1062 2676 1068 2677
rect 1214 2681 1220 2682
rect 1214 2677 1215 2681
rect 1219 2677 1220 2681
rect 1214 2676 1220 2677
rect 1374 2681 1380 2682
rect 1374 2677 1375 2681
rect 1379 2677 1380 2681
rect 1374 2676 1380 2677
rect 1534 2681 1540 2682
rect 1534 2677 1535 2681
rect 1539 2677 1540 2681
rect 1534 2676 1540 2677
rect 1670 2681 1676 2682
rect 1670 2677 1671 2681
rect 1675 2677 1676 2681
rect 1670 2676 1676 2677
rect 1766 2680 1772 2681
rect 1766 2676 1767 2680
rect 1771 2676 1772 2680
rect 1806 2680 1807 2684
rect 1811 2680 1812 2684
rect 2038 2681 2039 2685
rect 2043 2681 2044 2685
rect 2038 2680 2044 2681
rect 2158 2685 2164 2686
rect 2158 2681 2159 2685
rect 2163 2681 2164 2685
rect 2158 2680 2164 2681
rect 2278 2685 2284 2686
rect 2278 2681 2279 2685
rect 2283 2681 2284 2685
rect 2278 2680 2284 2681
rect 2406 2685 2412 2686
rect 2406 2681 2407 2685
rect 2411 2681 2412 2685
rect 2406 2680 2412 2681
rect 2542 2685 2548 2686
rect 2542 2681 2543 2685
rect 2547 2681 2548 2685
rect 2542 2680 2548 2681
rect 2686 2685 2692 2686
rect 2686 2681 2687 2685
rect 2691 2681 2692 2685
rect 2686 2680 2692 2681
rect 2846 2685 2852 2686
rect 2846 2681 2847 2685
rect 2851 2681 2852 2685
rect 2846 2680 2852 2681
rect 3022 2685 3028 2686
rect 3022 2681 3023 2685
rect 3027 2681 3028 2685
rect 3022 2680 3028 2681
rect 3206 2685 3212 2686
rect 3206 2681 3207 2685
rect 3211 2681 3212 2685
rect 3206 2680 3212 2681
rect 3366 2685 3372 2686
rect 3366 2681 3367 2685
rect 3371 2681 3372 2685
rect 3366 2680 3372 2681
rect 3462 2684 3468 2685
rect 3462 2680 3463 2684
rect 3467 2680 3468 2684
rect 1806 2679 1812 2680
rect 3462 2679 3468 2680
rect 110 2675 116 2676
rect 1766 2675 1772 2676
rect 110 2628 116 2629
rect 1766 2628 1772 2629
rect 110 2624 111 2628
rect 115 2624 116 2628
rect 110 2623 116 2624
rect 462 2627 468 2628
rect 462 2623 463 2627
rect 467 2623 468 2627
rect 462 2622 468 2623
rect 550 2627 556 2628
rect 550 2623 551 2627
rect 555 2623 556 2627
rect 550 2622 556 2623
rect 638 2627 644 2628
rect 638 2623 639 2627
rect 643 2623 644 2627
rect 638 2622 644 2623
rect 742 2627 748 2628
rect 742 2623 743 2627
rect 747 2623 748 2627
rect 742 2622 748 2623
rect 854 2627 860 2628
rect 854 2623 855 2627
rect 859 2623 860 2627
rect 854 2622 860 2623
rect 982 2627 988 2628
rect 982 2623 983 2627
rect 987 2623 988 2627
rect 982 2622 988 2623
rect 1126 2627 1132 2628
rect 1126 2623 1127 2627
rect 1131 2623 1132 2627
rect 1126 2622 1132 2623
rect 1278 2627 1284 2628
rect 1278 2623 1279 2627
rect 1283 2623 1284 2627
rect 1278 2622 1284 2623
rect 1438 2627 1444 2628
rect 1438 2623 1439 2627
rect 1443 2623 1444 2627
rect 1438 2622 1444 2623
rect 1606 2627 1612 2628
rect 1606 2623 1607 2627
rect 1611 2623 1612 2627
rect 1766 2624 1767 2628
rect 1771 2624 1772 2628
rect 1766 2623 1772 2624
rect 1806 2628 1812 2629
rect 3462 2628 3468 2629
rect 1806 2624 1807 2628
rect 1811 2624 1812 2628
rect 1806 2623 1812 2624
rect 1870 2627 1876 2628
rect 1870 2623 1871 2627
rect 1875 2623 1876 2627
rect 1606 2622 1612 2623
rect 1870 2622 1876 2623
rect 1966 2627 1972 2628
rect 1966 2623 1967 2627
rect 1971 2623 1972 2627
rect 1966 2622 1972 2623
rect 2070 2627 2076 2628
rect 2070 2623 2071 2627
rect 2075 2623 2076 2627
rect 2070 2622 2076 2623
rect 2182 2627 2188 2628
rect 2182 2623 2183 2627
rect 2187 2623 2188 2627
rect 2182 2622 2188 2623
rect 2294 2627 2300 2628
rect 2294 2623 2295 2627
rect 2299 2623 2300 2627
rect 2294 2622 2300 2623
rect 2430 2627 2436 2628
rect 2430 2623 2431 2627
rect 2435 2623 2436 2627
rect 2430 2622 2436 2623
rect 2582 2627 2588 2628
rect 2582 2623 2583 2627
rect 2587 2623 2588 2627
rect 2582 2622 2588 2623
rect 2758 2627 2764 2628
rect 2758 2623 2759 2627
rect 2763 2623 2764 2627
rect 2758 2622 2764 2623
rect 2958 2627 2964 2628
rect 2958 2623 2959 2627
rect 2963 2623 2964 2627
rect 2958 2622 2964 2623
rect 3166 2627 3172 2628
rect 3166 2623 3167 2627
rect 3171 2623 3172 2627
rect 3166 2622 3172 2623
rect 3366 2627 3372 2628
rect 3366 2623 3367 2627
rect 3371 2623 3372 2627
rect 3462 2624 3463 2628
rect 3467 2624 3468 2628
rect 3462 2623 3468 2624
rect 3366 2622 3372 2623
rect 110 2611 116 2612
rect 110 2607 111 2611
rect 115 2607 116 2611
rect 1766 2611 1772 2612
rect 110 2606 116 2607
rect 462 2608 468 2609
rect 462 2604 463 2608
rect 467 2604 468 2608
rect 462 2603 468 2604
rect 550 2608 556 2609
rect 550 2604 551 2608
rect 555 2604 556 2608
rect 550 2603 556 2604
rect 638 2608 644 2609
rect 638 2604 639 2608
rect 643 2604 644 2608
rect 638 2603 644 2604
rect 742 2608 748 2609
rect 742 2604 743 2608
rect 747 2604 748 2608
rect 742 2603 748 2604
rect 854 2608 860 2609
rect 854 2604 855 2608
rect 859 2604 860 2608
rect 854 2603 860 2604
rect 982 2608 988 2609
rect 982 2604 983 2608
rect 987 2604 988 2608
rect 982 2603 988 2604
rect 1126 2608 1132 2609
rect 1126 2604 1127 2608
rect 1131 2604 1132 2608
rect 1126 2603 1132 2604
rect 1278 2608 1284 2609
rect 1278 2604 1279 2608
rect 1283 2604 1284 2608
rect 1278 2603 1284 2604
rect 1438 2608 1444 2609
rect 1438 2604 1439 2608
rect 1443 2604 1444 2608
rect 1438 2603 1444 2604
rect 1606 2608 1612 2609
rect 1606 2604 1607 2608
rect 1611 2604 1612 2608
rect 1766 2607 1767 2611
rect 1771 2607 1772 2611
rect 1766 2606 1772 2607
rect 1806 2611 1812 2612
rect 1806 2607 1807 2611
rect 1811 2607 1812 2611
rect 3462 2611 3468 2612
rect 1806 2606 1812 2607
rect 1870 2608 1876 2609
rect 1606 2603 1612 2604
rect 1870 2604 1871 2608
rect 1875 2604 1876 2608
rect 1870 2603 1876 2604
rect 1966 2608 1972 2609
rect 1966 2604 1967 2608
rect 1971 2604 1972 2608
rect 1966 2603 1972 2604
rect 2070 2608 2076 2609
rect 2070 2604 2071 2608
rect 2075 2604 2076 2608
rect 2070 2603 2076 2604
rect 2182 2608 2188 2609
rect 2182 2604 2183 2608
rect 2187 2604 2188 2608
rect 2182 2603 2188 2604
rect 2294 2608 2300 2609
rect 2294 2604 2295 2608
rect 2299 2604 2300 2608
rect 2294 2603 2300 2604
rect 2430 2608 2436 2609
rect 2430 2604 2431 2608
rect 2435 2604 2436 2608
rect 2430 2603 2436 2604
rect 2582 2608 2588 2609
rect 2582 2604 2583 2608
rect 2587 2604 2588 2608
rect 2582 2603 2588 2604
rect 2758 2608 2764 2609
rect 2758 2604 2759 2608
rect 2763 2604 2764 2608
rect 2758 2603 2764 2604
rect 2958 2608 2964 2609
rect 2958 2604 2959 2608
rect 2963 2604 2964 2608
rect 2958 2603 2964 2604
rect 3166 2608 3172 2609
rect 3166 2604 3167 2608
rect 3171 2604 3172 2608
rect 3166 2603 3172 2604
rect 3366 2608 3372 2609
rect 3366 2604 3367 2608
rect 3371 2604 3372 2608
rect 3462 2607 3463 2611
rect 3467 2607 3468 2611
rect 3462 2606 3468 2607
rect 3366 2603 3372 2604
rect 502 2556 508 2557
rect 110 2553 116 2554
rect 110 2549 111 2553
rect 115 2549 116 2553
rect 502 2552 503 2556
rect 507 2552 508 2556
rect 502 2551 508 2552
rect 590 2556 596 2557
rect 590 2552 591 2556
rect 595 2552 596 2556
rect 590 2551 596 2552
rect 678 2556 684 2557
rect 678 2552 679 2556
rect 683 2552 684 2556
rect 678 2551 684 2552
rect 774 2556 780 2557
rect 774 2552 775 2556
rect 779 2552 780 2556
rect 774 2551 780 2552
rect 878 2556 884 2557
rect 878 2552 879 2556
rect 883 2552 884 2556
rect 878 2551 884 2552
rect 990 2556 996 2557
rect 990 2552 991 2556
rect 995 2552 996 2556
rect 990 2551 996 2552
rect 1102 2556 1108 2557
rect 1102 2552 1103 2556
rect 1107 2552 1108 2556
rect 1102 2551 1108 2552
rect 1222 2556 1228 2557
rect 1222 2552 1223 2556
rect 1227 2552 1228 2556
rect 1222 2551 1228 2552
rect 1350 2556 1356 2557
rect 1350 2552 1351 2556
rect 1355 2552 1356 2556
rect 1350 2551 1356 2552
rect 1478 2556 1484 2557
rect 1478 2552 1479 2556
rect 1483 2552 1484 2556
rect 1478 2551 1484 2552
rect 1606 2556 1612 2557
rect 1606 2552 1607 2556
rect 1611 2552 1612 2556
rect 1606 2551 1612 2552
rect 1766 2553 1772 2554
rect 110 2548 116 2549
rect 1766 2549 1767 2553
rect 1771 2549 1772 2553
rect 1830 2552 1836 2553
rect 1766 2548 1772 2549
rect 1806 2549 1812 2550
rect 1806 2545 1807 2549
rect 1811 2545 1812 2549
rect 1830 2548 1831 2552
rect 1835 2548 1836 2552
rect 1830 2547 1836 2548
rect 1918 2552 1924 2553
rect 1918 2548 1919 2552
rect 1923 2548 1924 2552
rect 1918 2547 1924 2548
rect 2006 2552 2012 2553
rect 2006 2548 2007 2552
rect 2011 2548 2012 2552
rect 2006 2547 2012 2548
rect 2110 2552 2116 2553
rect 2110 2548 2111 2552
rect 2115 2548 2116 2552
rect 2110 2547 2116 2548
rect 2222 2552 2228 2553
rect 2222 2548 2223 2552
rect 2227 2548 2228 2552
rect 2222 2547 2228 2548
rect 2342 2552 2348 2553
rect 2342 2548 2343 2552
rect 2347 2548 2348 2552
rect 2342 2547 2348 2548
rect 2486 2552 2492 2553
rect 2486 2548 2487 2552
rect 2491 2548 2492 2552
rect 2486 2547 2492 2548
rect 2646 2552 2652 2553
rect 2646 2548 2647 2552
rect 2651 2548 2652 2552
rect 2646 2547 2652 2548
rect 2814 2552 2820 2553
rect 2814 2548 2815 2552
rect 2819 2548 2820 2552
rect 2814 2547 2820 2548
rect 2998 2552 3004 2553
rect 2998 2548 2999 2552
rect 3003 2548 3004 2552
rect 2998 2547 3004 2548
rect 3190 2552 3196 2553
rect 3190 2548 3191 2552
rect 3195 2548 3196 2552
rect 3190 2547 3196 2548
rect 3366 2552 3372 2553
rect 3366 2548 3367 2552
rect 3371 2548 3372 2552
rect 3366 2547 3372 2548
rect 3462 2549 3468 2550
rect 1806 2544 1812 2545
rect 3462 2545 3463 2549
rect 3467 2545 3468 2549
rect 3462 2544 3468 2545
rect 502 2537 508 2538
rect 110 2536 116 2537
rect 110 2532 111 2536
rect 115 2532 116 2536
rect 502 2533 503 2537
rect 507 2533 508 2537
rect 502 2532 508 2533
rect 590 2537 596 2538
rect 590 2533 591 2537
rect 595 2533 596 2537
rect 590 2532 596 2533
rect 678 2537 684 2538
rect 678 2533 679 2537
rect 683 2533 684 2537
rect 678 2532 684 2533
rect 774 2537 780 2538
rect 774 2533 775 2537
rect 779 2533 780 2537
rect 774 2532 780 2533
rect 878 2537 884 2538
rect 878 2533 879 2537
rect 883 2533 884 2537
rect 878 2532 884 2533
rect 990 2537 996 2538
rect 990 2533 991 2537
rect 995 2533 996 2537
rect 990 2532 996 2533
rect 1102 2537 1108 2538
rect 1102 2533 1103 2537
rect 1107 2533 1108 2537
rect 1102 2532 1108 2533
rect 1222 2537 1228 2538
rect 1222 2533 1223 2537
rect 1227 2533 1228 2537
rect 1222 2532 1228 2533
rect 1350 2537 1356 2538
rect 1350 2533 1351 2537
rect 1355 2533 1356 2537
rect 1350 2532 1356 2533
rect 1478 2537 1484 2538
rect 1478 2533 1479 2537
rect 1483 2533 1484 2537
rect 1478 2532 1484 2533
rect 1606 2537 1612 2538
rect 1606 2533 1607 2537
rect 1611 2533 1612 2537
rect 1606 2532 1612 2533
rect 1766 2536 1772 2537
rect 1766 2532 1767 2536
rect 1771 2532 1772 2536
rect 1830 2533 1836 2534
rect 110 2531 116 2532
rect 1766 2531 1772 2532
rect 1806 2532 1812 2533
rect 1806 2528 1807 2532
rect 1811 2528 1812 2532
rect 1830 2529 1831 2533
rect 1835 2529 1836 2533
rect 1830 2528 1836 2529
rect 1918 2533 1924 2534
rect 1918 2529 1919 2533
rect 1923 2529 1924 2533
rect 1918 2528 1924 2529
rect 2006 2533 2012 2534
rect 2006 2529 2007 2533
rect 2011 2529 2012 2533
rect 2006 2528 2012 2529
rect 2110 2533 2116 2534
rect 2110 2529 2111 2533
rect 2115 2529 2116 2533
rect 2110 2528 2116 2529
rect 2222 2533 2228 2534
rect 2222 2529 2223 2533
rect 2227 2529 2228 2533
rect 2222 2528 2228 2529
rect 2342 2533 2348 2534
rect 2342 2529 2343 2533
rect 2347 2529 2348 2533
rect 2342 2528 2348 2529
rect 2486 2533 2492 2534
rect 2486 2529 2487 2533
rect 2491 2529 2492 2533
rect 2486 2528 2492 2529
rect 2646 2533 2652 2534
rect 2646 2529 2647 2533
rect 2651 2529 2652 2533
rect 2646 2528 2652 2529
rect 2814 2533 2820 2534
rect 2814 2529 2815 2533
rect 2819 2529 2820 2533
rect 2814 2528 2820 2529
rect 2998 2533 3004 2534
rect 2998 2529 2999 2533
rect 3003 2529 3004 2533
rect 2998 2528 3004 2529
rect 3190 2533 3196 2534
rect 3190 2529 3191 2533
rect 3195 2529 3196 2533
rect 3190 2528 3196 2529
rect 3366 2533 3372 2534
rect 3366 2529 3367 2533
rect 3371 2529 3372 2533
rect 3366 2528 3372 2529
rect 3462 2532 3468 2533
rect 3462 2528 3463 2532
rect 3467 2528 3468 2532
rect 1806 2527 1812 2528
rect 3462 2527 3468 2528
rect 1806 2488 1812 2489
rect 3462 2488 3468 2489
rect 110 2484 116 2485
rect 1766 2484 1772 2485
rect 110 2480 111 2484
rect 115 2480 116 2484
rect 110 2479 116 2480
rect 550 2483 556 2484
rect 550 2479 551 2483
rect 555 2479 556 2483
rect 550 2478 556 2479
rect 734 2483 740 2484
rect 734 2479 735 2483
rect 739 2479 740 2483
rect 734 2478 740 2479
rect 910 2483 916 2484
rect 910 2479 911 2483
rect 915 2479 916 2483
rect 910 2478 916 2479
rect 1078 2483 1084 2484
rect 1078 2479 1079 2483
rect 1083 2479 1084 2483
rect 1078 2478 1084 2479
rect 1238 2483 1244 2484
rect 1238 2479 1239 2483
rect 1243 2479 1244 2483
rect 1238 2478 1244 2479
rect 1398 2483 1404 2484
rect 1398 2479 1399 2483
rect 1403 2479 1404 2483
rect 1398 2478 1404 2479
rect 1566 2483 1572 2484
rect 1566 2479 1567 2483
rect 1571 2479 1572 2483
rect 1766 2480 1767 2484
rect 1771 2480 1772 2484
rect 1806 2484 1807 2488
rect 1811 2484 1812 2488
rect 1806 2483 1812 2484
rect 1950 2487 1956 2488
rect 1950 2483 1951 2487
rect 1955 2483 1956 2487
rect 1950 2482 1956 2483
rect 2038 2487 2044 2488
rect 2038 2483 2039 2487
rect 2043 2483 2044 2487
rect 2038 2482 2044 2483
rect 2134 2487 2140 2488
rect 2134 2483 2135 2487
rect 2139 2483 2140 2487
rect 2134 2482 2140 2483
rect 2238 2487 2244 2488
rect 2238 2483 2239 2487
rect 2243 2483 2244 2487
rect 2238 2482 2244 2483
rect 2366 2487 2372 2488
rect 2366 2483 2367 2487
rect 2371 2483 2372 2487
rect 2366 2482 2372 2483
rect 2526 2487 2532 2488
rect 2526 2483 2527 2487
rect 2531 2483 2532 2487
rect 2526 2482 2532 2483
rect 2710 2487 2716 2488
rect 2710 2483 2711 2487
rect 2715 2483 2716 2487
rect 2710 2482 2716 2483
rect 2918 2487 2924 2488
rect 2918 2483 2919 2487
rect 2923 2483 2924 2487
rect 2918 2482 2924 2483
rect 3142 2487 3148 2488
rect 3142 2483 3143 2487
rect 3147 2483 3148 2487
rect 3142 2482 3148 2483
rect 3366 2487 3372 2488
rect 3366 2483 3367 2487
rect 3371 2483 3372 2487
rect 3462 2484 3463 2488
rect 3467 2484 3468 2488
rect 3462 2483 3468 2484
rect 3366 2482 3372 2483
rect 1766 2479 1772 2480
rect 1566 2478 1572 2479
rect 1806 2471 1812 2472
rect 110 2467 116 2468
rect 110 2463 111 2467
rect 115 2463 116 2467
rect 1766 2467 1772 2468
rect 110 2462 116 2463
rect 550 2464 556 2465
rect 550 2460 551 2464
rect 555 2460 556 2464
rect 550 2459 556 2460
rect 734 2464 740 2465
rect 734 2460 735 2464
rect 739 2460 740 2464
rect 734 2459 740 2460
rect 910 2464 916 2465
rect 910 2460 911 2464
rect 915 2460 916 2464
rect 910 2459 916 2460
rect 1078 2464 1084 2465
rect 1078 2460 1079 2464
rect 1083 2460 1084 2464
rect 1078 2459 1084 2460
rect 1238 2464 1244 2465
rect 1238 2460 1239 2464
rect 1243 2460 1244 2464
rect 1238 2459 1244 2460
rect 1398 2464 1404 2465
rect 1398 2460 1399 2464
rect 1403 2460 1404 2464
rect 1398 2459 1404 2460
rect 1566 2464 1572 2465
rect 1566 2460 1567 2464
rect 1571 2460 1572 2464
rect 1766 2463 1767 2467
rect 1771 2463 1772 2467
rect 1806 2467 1807 2471
rect 1811 2467 1812 2471
rect 3462 2471 3468 2472
rect 1806 2466 1812 2467
rect 1950 2468 1956 2469
rect 1950 2464 1951 2468
rect 1955 2464 1956 2468
rect 1950 2463 1956 2464
rect 2038 2468 2044 2469
rect 2038 2464 2039 2468
rect 2043 2464 2044 2468
rect 2038 2463 2044 2464
rect 2134 2468 2140 2469
rect 2134 2464 2135 2468
rect 2139 2464 2140 2468
rect 2134 2463 2140 2464
rect 2238 2468 2244 2469
rect 2238 2464 2239 2468
rect 2243 2464 2244 2468
rect 2238 2463 2244 2464
rect 2366 2468 2372 2469
rect 2366 2464 2367 2468
rect 2371 2464 2372 2468
rect 2366 2463 2372 2464
rect 2526 2468 2532 2469
rect 2526 2464 2527 2468
rect 2531 2464 2532 2468
rect 2526 2463 2532 2464
rect 2710 2468 2716 2469
rect 2710 2464 2711 2468
rect 2715 2464 2716 2468
rect 2710 2463 2716 2464
rect 2918 2468 2924 2469
rect 2918 2464 2919 2468
rect 2923 2464 2924 2468
rect 2918 2463 2924 2464
rect 3142 2468 3148 2469
rect 3142 2464 3143 2468
rect 3147 2464 3148 2468
rect 3142 2463 3148 2464
rect 3366 2468 3372 2469
rect 3366 2464 3367 2468
rect 3371 2464 3372 2468
rect 3462 2467 3463 2471
rect 3467 2467 3468 2471
rect 3462 2466 3468 2467
rect 3366 2463 3372 2464
rect 1766 2462 1772 2463
rect 1566 2459 1572 2460
rect 414 2420 420 2421
rect 110 2417 116 2418
rect 110 2413 111 2417
rect 115 2413 116 2417
rect 414 2416 415 2420
rect 419 2416 420 2420
rect 414 2415 420 2416
rect 502 2420 508 2421
rect 502 2416 503 2420
rect 507 2416 508 2420
rect 502 2415 508 2416
rect 598 2420 604 2421
rect 598 2416 599 2420
rect 603 2416 604 2420
rect 598 2415 604 2416
rect 702 2420 708 2421
rect 702 2416 703 2420
rect 707 2416 708 2420
rect 702 2415 708 2416
rect 806 2420 812 2421
rect 806 2416 807 2420
rect 811 2416 812 2420
rect 806 2415 812 2416
rect 918 2420 924 2421
rect 918 2416 919 2420
rect 923 2416 924 2420
rect 918 2415 924 2416
rect 1038 2420 1044 2421
rect 1038 2416 1039 2420
rect 1043 2416 1044 2420
rect 1038 2415 1044 2416
rect 1166 2420 1172 2421
rect 1166 2416 1167 2420
rect 1171 2416 1172 2420
rect 1166 2415 1172 2416
rect 1294 2420 1300 2421
rect 1294 2416 1295 2420
rect 1299 2416 1300 2420
rect 1294 2415 1300 2416
rect 1422 2420 1428 2421
rect 1422 2416 1423 2420
rect 1427 2416 1428 2420
rect 1422 2415 1428 2416
rect 1766 2417 1772 2418
rect 110 2412 116 2413
rect 1766 2413 1767 2417
rect 1771 2413 1772 2417
rect 2214 2416 2220 2417
rect 1766 2412 1772 2413
rect 1806 2413 1812 2414
rect 1806 2409 1807 2413
rect 1811 2409 1812 2413
rect 2214 2412 2215 2416
rect 2219 2412 2220 2416
rect 2214 2411 2220 2412
rect 2302 2416 2308 2417
rect 2302 2412 2303 2416
rect 2307 2412 2308 2416
rect 2302 2411 2308 2412
rect 2390 2416 2396 2417
rect 2390 2412 2391 2416
rect 2395 2412 2396 2416
rect 2390 2411 2396 2412
rect 2478 2416 2484 2417
rect 2478 2412 2479 2416
rect 2483 2412 2484 2416
rect 2478 2411 2484 2412
rect 2566 2416 2572 2417
rect 2566 2412 2567 2416
rect 2571 2412 2572 2416
rect 2566 2411 2572 2412
rect 2654 2416 2660 2417
rect 2654 2412 2655 2416
rect 2659 2412 2660 2416
rect 2654 2411 2660 2412
rect 2742 2416 2748 2417
rect 2742 2412 2743 2416
rect 2747 2412 2748 2416
rect 2742 2411 2748 2412
rect 2838 2416 2844 2417
rect 2838 2412 2839 2416
rect 2843 2412 2844 2416
rect 2838 2411 2844 2412
rect 2934 2416 2940 2417
rect 2934 2412 2935 2416
rect 2939 2412 2940 2416
rect 2934 2411 2940 2412
rect 3462 2413 3468 2414
rect 1806 2408 1812 2409
rect 3462 2409 3463 2413
rect 3467 2409 3468 2413
rect 3462 2408 3468 2409
rect 414 2401 420 2402
rect 110 2400 116 2401
rect 110 2396 111 2400
rect 115 2396 116 2400
rect 414 2397 415 2401
rect 419 2397 420 2401
rect 414 2396 420 2397
rect 502 2401 508 2402
rect 502 2397 503 2401
rect 507 2397 508 2401
rect 502 2396 508 2397
rect 598 2401 604 2402
rect 598 2397 599 2401
rect 603 2397 604 2401
rect 598 2396 604 2397
rect 702 2401 708 2402
rect 702 2397 703 2401
rect 707 2397 708 2401
rect 702 2396 708 2397
rect 806 2401 812 2402
rect 806 2397 807 2401
rect 811 2397 812 2401
rect 806 2396 812 2397
rect 918 2401 924 2402
rect 918 2397 919 2401
rect 923 2397 924 2401
rect 918 2396 924 2397
rect 1038 2401 1044 2402
rect 1038 2397 1039 2401
rect 1043 2397 1044 2401
rect 1038 2396 1044 2397
rect 1166 2401 1172 2402
rect 1166 2397 1167 2401
rect 1171 2397 1172 2401
rect 1166 2396 1172 2397
rect 1294 2401 1300 2402
rect 1294 2397 1295 2401
rect 1299 2397 1300 2401
rect 1294 2396 1300 2397
rect 1422 2401 1428 2402
rect 1422 2397 1423 2401
rect 1427 2397 1428 2401
rect 1422 2396 1428 2397
rect 1766 2400 1772 2401
rect 1766 2396 1767 2400
rect 1771 2396 1772 2400
rect 2214 2397 2220 2398
rect 110 2395 116 2396
rect 1766 2395 1772 2396
rect 1806 2396 1812 2397
rect 1806 2392 1807 2396
rect 1811 2392 1812 2396
rect 2214 2393 2215 2397
rect 2219 2393 2220 2397
rect 2214 2392 2220 2393
rect 2302 2397 2308 2398
rect 2302 2393 2303 2397
rect 2307 2393 2308 2397
rect 2302 2392 2308 2393
rect 2390 2397 2396 2398
rect 2390 2393 2391 2397
rect 2395 2393 2396 2397
rect 2390 2392 2396 2393
rect 2478 2397 2484 2398
rect 2478 2393 2479 2397
rect 2483 2393 2484 2397
rect 2478 2392 2484 2393
rect 2566 2397 2572 2398
rect 2566 2393 2567 2397
rect 2571 2393 2572 2397
rect 2566 2392 2572 2393
rect 2654 2397 2660 2398
rect 2654 2393 2655 2397
rect 2659 2393 2660 2397
rect 2654 2392 2660 2393
rect 2742 2397 2748 2398
rect 2742 2393 2743 2397
rect 2747 2393 2748 2397
rect 2742 2392 2748 2393
rect 2838 2397 2844 2398
rect 2838 2393 2839 2397
rect 2843 2393 2844 2397
rect 2838 2392 2844 2393
rect 2934 2397 2940 2398
rect 2934 2393 2935 2397
rect 2939 2393 2940 2397
rect 2934 2392 2940 2393
rect 3462 2396 3468 2397
rect 3462 2392 3463 2396
rect 3467 2392 3468 2396
rect 1806 2391 1812 2392
rect 3462 2391 3468 2392
rect 110 2352 116 2353
rect 1766 2352 1772 2353
rect 110 2348 111 2352
rect 115 2348 116 2352
rect 110 2347 116 2348
rect 318 2351 324 2352
rect 318 2347 319 2351
rect 323 2347 324 2351
rect 318 2346 324 2347
rect 430 2351 436 2352
rect 430 2347 431 2351
rect 435 2347 436 2351
rect 430 2346 436 2347
rect 542 2351 548 2352
rect 542 2347 543 2351
rect 547 2347 548 2351
rect 542 2346 548 2347
rect 654 2351 660 2352
rect 654 2347 655 2351
rect 659 2347 660 2351
rect 654 2346 660 2347
rect 766 2351 772 2352
rect 766 2347 767 2351
rect 771 2347 772 2351
rect 766 2346 772 2347
rect 878 2351 884 2352
rect 878 2347 879 2351
rect 883 2347 884 2351
rect 878 2346 884 2347
rect 990 2351 996 2352
rect 990 2347 991 2351
rect 995 2347 996 2351
rect 990 2346 996 2347
rect 1102 2351 1108 2352
rect 1102 2347 1103 2351
rect 1107 2347 1108 2351
rect 1102 2346 1108 2347
rect 1214 2351 1220 2352
rect 1214 2347 1215 2351
rect 1219 2347 1220 2351
rect 1214 2346 1220 2347
rect 1334 2351 1340 2352
rect 1334 2347 1335 2351
rect 1339 2347 1340 2351
rect 1766 2348 1767 2352
rect 1771 2348 1772 2352
rect 1766 2347 1772 2348
rect 1806 2352 1812 2353
rect 3462 2352 3468 2353
rect 1806 2348 1807 2352
rect 1811 2348 1812 2352
rect 1806 2347 1812 2348
rect 2166 2351 2172 2352
rect 2166 2347 2167 2351
rect 2171 2347 2172 2351
rect 1334 2346 1340 2347
rect 2166 2346 2172 2347
rect 2262 2351 2268 2352
rect 2262 2347 2263 2351
rect 2267 2347 2268 2351
rect 2262 2346 2268 2347
rect 2366 2351 2372 2352
rect 2366 2347 2367 2351
rect 2371 2347 2372 2351
rect 2366 2346 2372 2347
rect 2470 2351 2476 2352
rect 2470 2347 2471 2351
rect 2475 2347 2476 2351
rect 2470 2346 2476 2347
rect 2574 2351 2580 2352
rect 2574 2347 2575 2351
rect 2579 2347 2580 2351
rect 2574 2346 2580 2347
rect 2686 2351 2692 2352
rect 2686 2347 2687 2351
rect 2691 2347 2692 2351
rect 2686 2346 2692 2347
rect 2798 2351 2804 2352
rect 2798 2347 2799 2351
rect 2803 2347 2804 2351
rect 2798 2346 2804 2347
rect 2910 2351 2916 2352
rect 2910 2347 2911 2351
rect 2915 2347 2916 2351
rect 2910 2346 2916 2347
rect 3022 2351 3028 2352
rect 3022 2347 3023 2351
rect 3027 2347 3028 2351
rect 3462 2348 3463 2352
rect 3467 2348 3468 2352
rect 3462 2347 3468 2348
rect 3022 2346 3028 2347
rect 110 2335 116 2336
rect 110 2331 111 2335
rect 115 2331 116 2335
rect 1766 2335 1772 2336
rect 110 2330 116 2331
rect 318 2332 324 2333
rect 318 2328 319 2332
rect 323 2328 324 2332
rect 318 2327 324 2328
rect 430 2332 436 2333
rect 430 2328 431 2332
rect 435 2328 436 2332
rect 430 2327 436 2328
rect 542 2332 548 2333
rect 542 2328 543 2332
rect 547 2328 548 2332
rect 542 2327 548 2328
rect 654 2332 660 2333
rect 654 2328 655 2332
rect 659 2328 660 2332
rect 654 2327 660 2328
rect 766 2332 772 2333
rect 766 2328 767 2332
rect 771 2328 772 2332
rect 766 2327 772 2328
rect 878 2332 884 2333
rect 878 2328 879 2332
rect 883 2328 884 2332
rect 878 2327 884 2328
rect 990 2332 996 2333
rect 990 2328 991 2332
rect 995 2328 996 2332
rect 990 2327 996 2328
rect 1102 2332 1108 2333
rect 1102 2328 1103 2332
rect 1107 2328 1108 2332
rect 1102 2327 1108 2328
rect 1214 2332 1220 2333
rect 1214 2328 1215 2332
rect 1219 2328 1220 2332
rect 1214 2327 1220 2328
rect 1334 2332 1340 2333
rect 1334 2328 1335 2332
rect 1339 2328 1340 2332
rect 1766 2331 1767 2335
rect 1771 2331 1772 2335
rect 1766 2330 1772 2331
rect 1806 2335 1812 2336
rect 1806 2331 1807 2335
rect 1811 2331 1812 2335
rect 3462 2335 3468 2336
rect 1806 2330 1812 2331
rect 2166 2332 2172 2333
rect 1334 2327 1340 2328
rect 2166 2328 2167 2332
rect 2171 2328 2172 2332
rect 2166 2327 2172 2328
rect 2262 2332 2268 2333
rect 2262 2328 2263 2332
rect 2267 2328 2268 2332
rect 2262 2327 2268 2328
rect 2366 2332 2372 2333
rect 2366 2328 2367 2332
rect 2371 2328 2372 2332
rect 2366 2327 2372 2328
rect 2470 2332 2476 2333
rect 2470 2328 2471 2332
rect 2475 2328 2476 2332
rect 2470 2327 2476 2328
rect 2574 2332 2580 2333
rect 2574 2328 2575 2332
rect 2579 2328 2580 2332
rect 2574 2327 2580 2328
rect 2686 2332 2692 2333
rect 2686 2328 2687 2332
rect 2691 2328 2692 2332
rect 2686 2327 2692 2328
rect 2798 2332 2804 2333
rect 2798 2328 2799 2332
rect 2803 2328 2804 2332
rect 2798 2327 2804 2328
rect 2910 2332 2916 2333
rect 2910 2328 2911 2332
rect 2915 2328 2916 2332
rect 2910 2327 2916 2328
rect 3022 2332 3028 2333
rect 3022 2328 3023 2332
rect 3027 2328 3028 2332
rect 3462 2331 3463 2335
rect 3467 2331 3468 2335
rect 3462 2330 3468 2331
rect 3022 2327 3028 2328
rect 150 2280 156 2281
rect 110 2277 116 2278
rect 110 2273 111 2277
rect 115 2273 116 2277
rect 150 2276 151 2280
rect 155 2276 156 2280
rect 150 2275 156 2276
rect 270 2280 276 2281
rect 270 2276 271 2280
rect 275 2276 276 2280
rect 270 2275 276 2276
rect 390 2280 396 2281
rect 390 2276 391 2280
rect 395 2276 396 2280
rect 390 2275 396 2276
rect 518 2280 524 2281
rect 518 2276 519 2280
rect 523 2276 524 2280
rect 518 2275 524 2276
rect 646 2280 652 2281
rect 646 2276 647 2280
rect 651 2276 652 2280
rect 646 2275 652 2276
rect 774 2280 780 2281
rect 774 2276 775 2280
rect 779 2276 780 2280
rect 774 2275 780 2276
rect 894 2280 900 2281
rect 894 2276 895 2280
rect 899 2276 900 2280
rect 894 2275 900 2276
rect 1014 2280 1020 2281
rect 1014 2276 1015 2280
rect 1019 2276 1020 2280
rect 1014 2275 1020 2276
rect 1142 2280 1148 2281
rect 1142 2276 1143 2280
rect 1147 2276 1148 2280
rect 1142 2275 1148 2276
rect 1270 2280 1276 2281
rect 1270 2276 1271 2280
rect 1275 2276 1276 2280
rect 1886 2280 1892 2281
rect 1270 2275 1276 2276
rect 1766 2277 1772 2278
rect 110 2272 116 2273
rect 1766 2273 1767 2277
rect 1771 2273 1772 2277
rect 1766 2272 1772 2273
rect 1806 2277 1812 2278
rect 1806 2273 1807 2277
rect 1811 2273 1812 2277
rect 1886 2276 1887 2280
rect 1891 2276 1892 2280
rect 1886 2275 1892 2276
rect 2038 2280 2044 2281
rect 2038 2276 2039 2280
rect 2043 2276 2044 2280
rect 2038 2275 2044 2276
rect 2198 2280 2204 2281
rect 2198 2276 2199 2280
rect 2203 2276 2204 2280
rect 2198 2275 2204 2276
rect 2374 2280 2380 2281
rect 2374 2276 2375 2280
rect 2379 2276 2380 2280
rect 2374 2275 2380 2276
rect 2550 2280 2556 2281
rect 2550 2276 2551 2280
rect 2555 2276 2556 2280
rect 2550 2275 2556 2276
rect 2718 2280 2724 2281
rect 2718 2276 2719 2280
rect 2723 2276 2724 2280
rect 2718 2275 2724 2276
rect 2886 2280 2892 2281
rect 2886 2276 2887 2280
rect 2891 2276 2892 2280
rect 2886 2275 2892 2276
rect 3054 2280 3060 2281
rect 3054 2276 3055 2280
rect 3059 2276 3060 2280
rect 3054 2275 3060 2276
rect 3222 2280 3228 2281
rect 3222 2276 3223 2280
rect 3227 2276 3228 2280
rect 3222 2275 3228 2276
rect 3366 2280 3372 2281
rect 3366 2276 3367 2280
rect 3371 2276 3372 2280
rect 3366 2275 3372 2276
rect 3462 2277 3468 2278
rect 1806 2272 1812 2273
rect 3462 2273 3463 2277
rect 3467 2273 3468 2277
rect 3462 2272 3468 2273
rect 150 2261 156 2262
rect 110 2260 116 2261
rect 110 2256 111 2260
rect 115 2256 116 2260
rect 150 2257 151 2261
rect 155 2257 156 2261
rect 150 2256 156 2257
rect 270 2261 276 2262
rect 270 2257 271 2261
rect 275 2257 276 2261
rect 270 2256 276 2257
rect 390 2261 396 2262
rect 390 2257 391 2261
rect 395 2257 396 2261
rect 390 2256 396 2257
rect 518 2261 524 2262
rect 518 2257 519 2261
rect 523 2257 524 2261
rect 518 2256 524 2257
rect 646 2261 652 2262
rect 646 2257 647 2261
rect 651 2257 652 2261
rect 646 2256 652 2257
rect 774 2261 780 2262
rect 774 2257 775 2261
rect 779 2257 780 2261
rect 774 2256 780 2257
rect 894 2261 900 2262
rect 894 2257 895 2261
rect 899 2257 900 2261
rect 894 2256 900 2257
rect 1014 2261 1020 2262
rect 1014 2257 1015 2261
rect 1019 2257 1020 2261
rect 1014 2256 1020 2257
rect 1142 2261 1148 2262
rect 1142 2257 1143 2261
rect 1147 2257 1148 2261
rect 1142 2256 1148 2257
rect 1270 2261 1276 2262
rect 1886 2261 1892 2262
rect 1270 2257 1271 2261
rect 1275 2257 1276 2261
rect 1270 2256 1276 2257
rect 1766 2260 1772 2261
rect 1766 2256 1767 2260
rect 1771 2256 1772 2260
rect 110 2255 116 2256
rect 1766 2255 1772 2256
rect 1806 2260 1812 2261
rect 1806 2256 1807 2260
rect 1811 2256 1812 2260
rect 1886 2257 1887 2261
rect 1891 2257 1892 2261
rect 1886 2256 1892 2257
rect 2038 2261 2044 2262
rect 2038 2257 2039 2261
rect 2043 2257 2044 2261
rect 2038 2256 2044 2257
rect 2198 2261 2204 2262
rect 2198 2257 2199 2261
rect 2203 2257 2204 2261
rect 2198 2256 2204 2257
rect 2374 2261 2380 2262
rect 2374 2257 2375 2261
rect 2379 2257 2380 2261
rect 2374 2256 2380 2257
rect 2550 2261 2556 2262
rect 2550 2257 2551 2261
rect 2555 2257 2556 2261
rect 2550 2256 2556 2257
rect 2718 2261 2724 2262
rect 2718 2257 2719 2261
rect 2723 2257 2724 2261
rect 2718 2256 2724 2257
rect 2886 2261 2892 2262
rect 2886 2257 2887 2261
rect 2891 2257 2892 2261
rect 2886 2256 2892 2257
rect 3054 2261 3060 2262
rect 3054 2257 3055 2261
rect 3059 2257 3060 2261
rect 3054 2256 3060 2257
rect 3222 2261 3228 2262
rect 3222 2257 3223 2261
rect 3227 2257 3228 2261
rect 3222 2256 3228 2257
rect 3366 2261 3372 2262
rect 3366 2257 3367 2261
rect 3371 2257 3372 2261
rect 3366 2256 3372 2257
rect 3462 2260 3468 2261
rect 3462 2256 3463 2260
rect 3467 2256 3468 2260
rect 1806 2255 1812 2256
rect 3462 2255 3468 2256
rect 1806 2216 1812 2217
rect 3462 2216 3468 2217
rect 110 2212 116 2213
rect 1766 2212 1772 2213
rect 110 2208 111 2212
rect 115 2208 116 2212
rect 110 2207 116 2208
rect 134 2211 140 2212
rect 134 2207 135 2211
rect 139 2207 140 2211
rect 134 2206 140 2207
rect 246 2211 252 2212
rect 246 2207 247 2211
rect 251 2207 252 2211
rect 246 2206 252 2207
rect 406 2211 412 2212
rect 406 2207 407 2211
rect 411 2207 412 2211
rect 406 2206 412 2207
rect 582 2211 588 2212
rect 582 2207 583 2211
rect 587 2207 588 2211
rect 582 2206 588 2207
rect 766 2211 772 2212
rect 766 2207 767 2211
rect 771 2207 772 2211
rect 766 2206 772 2207
rect 950 2211 956 2212
rect 950 2207 951 2211
rect 955 2207 956 2211
rect 950 2206 956 2207
rect 1134 2211 1140 2212
rect 1134 2207 1135 2211
rect 1139 2207 1140 2211
rect 1134 2206 1140 2207
rect 1318 2211 1324 2212
rect 1318 2207 1319 2211
rect 1323 2207 1324 2211
rect 1318 2206 1324 2207
rect 1502 2211 1508 2212
rect 1502 2207 1503 2211
rect 1507 2207 1508 2211
rect 1502 2206 1508 2207
rect 1670 2211 1676 2212
rect 1670 2207 1671 2211
rect 1675 2207 1676 2211
rect 1766 2208 1767 2212
rect 1771 2208 1772 2212
rect 1806 2212 1807 2216
rect 1811 2212 1812 2216
rect 1806 2211 1812 2212
rect 1830 2215 1836 2216
rect 1830 2211 1831 2215
rect 1835 2211 1836 2215
rect 1830 2210 1836 2211
rect 1966 2215 1972 2216
rect 1966 2211 1967 2215
rect 1971 2211 1972 2215
rect 1966 2210 1972 2211
rect 2134 2215 2140 2216
rect 2134 2211 2135 2215
rect 2139 2211 2140 2215
rect 2134 2210 2140 2211
rect 2310 2215 2316 2216
rect 2310 2211 2311 2215
rect 2315 2211 2316 2215
rect 2310 2210 2316 2211
rect 2486 2215 2492 2216
rect 2486 2211 2487 2215
rect 2491 2211 2492 2215
rect 2486 2210 2492 2211
rect 2654 2215 2660 2216
rect 2654 2211 2655 2215
rect 2659 2211 2660 2215
rect 2654 2210 2660 2211
rect 2814 2215 2820 2216
rect 2814 2211 2815 2215
rect 2819 2211 2820 2215
rect 2814 2210 2820 2211
rect 2958 2215 2964 2216
rect 2958 2211 2959 2215
rect 2963 2211 2964 2215
rect 2958 2210 2964 2211
rect 3102 2215 3108 2216
rect 3102 2211 3103 2215
rect 3107 2211 3108 2215
rect 3102 2210 3108 2211
rect 3246 2215 3252 2216
rect 3246 2211 3247 2215
rect 3251 2211 3252 2215
rect 3246 2210 3252 2211
rect 3366 2215 3372 2216
rect 3366 2211 3367 2215
rect 3371 2211 3372 2215
rect 3462 2212 3463 2216
rect 3467 2212 3468 2216
rect 3462 2211 3468 2212
rect 3366 2210 3372 2211
rect 1766 2207 1772 2208
rect 1670 2206 1676 2207
rect 1806 2199 1812 2200
rect 110 2195 116 2196
rect 110 2191 111 2195
rect 115 2191 116 2195
rect 1766 2195 1772 2196
rect 110 2190 116 2191
rect 134 2192 140 2193
rect 134 2188 135 2192
rect 139 2188 140 2192
rect 134 2187 140 2188
rect 246 2192 252 2193
rect 246 2188 247 2192
rect 251 2188 252 2192
rect 246 2187 252 2188
rect 406 2192 412 2193
rect 406 2188 407 2192
rect 411 2188 412 2192
rect 406 2187 412 2188
rect 582 2192 588 2193
rect 582 2188 583 2192
rect 587 2188 588 2192
rect 582 2187 588 2188
rect 766 2192 772 2193
rect 766 2188 767 2192
rect 771 2188 772 2192
rect 766 2187 772 2188
rect 950 2192 956 2193
rect 950 2188 951 2192
rect 955 2188 956 2192
rect 950 2187 956 2188
rect 1134 2192 1140 2193
rect 1134 2188 1135 2192
rect 1139 2188 1140 2192
rect 1134 2187 1140 2188
rect 1318 2192 1324 2193
rect 1318 2188 1319 2192
rect 1323 2188 1324 2192
rect 1318 2187 1324 2188
rect 1502 2192 1508 2193
rect 1502 2188 1503 2192
rect 1507 2188 1508 2192
rect 1502 2187 1508 2188
rect 1670 2192 1676 2193
rect 1670 2188 1671 2192
rect 1675 2188 1676 2192
rect 1766 2191 1767 2195
rect 1771 2191 1772 2195
rect 1806 2195 1807 2199
rect 1811 2195 1812 2199
rect 3462 2199 3468 2200
rect 1806 2194 1812 2195
rect 1830 2196 1836 2197
rect 1830 2192 1831 2196
rect 1835 2192 1836 2196
rect 1830 2191 1836 2192
rect 1966 2196 1972 2197
rect 1966 2192 1967 2196
rect 1971 2192 1972 2196
rect 1966 2191 1972 2192
rect 2134 2196 2140 2197
rect 2134 2192 2135 2196
rect 2139 2192 2140 2196
rect 2134 2191 2140 2192
rect 2310 2196 2316 2197
rect 2310 2192 2311 2196
rect 2315 2192 2316 2196
rect 2310 2191 2316 2192
rect 2486 2196 2492 2197
rect 2486 2192 2487 2196
rect 2491 2192 2492 2196
rect 2486 2191 2492 2192
rect 2654 2196 2660 2197
rect 2654 2192 2655 2196
rect 2659 2192 2660 2196
rect 2654 2191 2660 2192
rect 2814 2196 2820 2197
rect 2814 2192 2815 2196
rect 2819 2192 2820 2196
rect 2814 2191 2820 2192
rect 2958 2196 2964 2197
rect 2958 2192 2959 2196
rect 2963 2192 2964 2196
rect 2958 2191 2964 2192
rect 3102 2196 3108 2197
rect 3102 2192 3103 2196
rect 3107 2192 3108 2196
rect 3102 2191 3108 2192
rect 3246 2196 3252 2197
rect 3246 2192 3247 2196
rect 3251 2192 3252 2196
rect 3246 2191 3252 2192
rect 3366 2196 3372 2197
rect 3366 2192 3367 2196
rect 3371 2192 3372 2196
rect 3462 2195 3463 2199
rect 3467 2195 3468 2199
rect 3462 2194 3468 2195
rect 3366 2191 3372 2192
rect 1766 2190 1772 2191
rect 1670 2187 1676 2188
rect 2926 2152 2932 2153
rect 1806 2149 1812 2150
rect 1806 2145 1807 2149
rect 1811 2145 1812 2149
rect 2926 2148 2927 2152
rect 2931 2148 2932 2152
rect 2926 2147 2932 2148
rect 3014 2152 3020 2153
rect 3014 2148 3015 2152
rect 3019 2148 3020 2152
rect 3014 2147 3020 2148
rect 3102 2152 3108 2153
rect 3102 2148 3103 2152
rect 3107 2148 3108 2152
rect 3102 2147 3108 2148
rect 3190 2152 3196 2153
rect 3190 2148 3191 2152
rect 3195 2148 3196 2152
rect 3190 2147 3196 2148
rect 3278 2152 3284 2153
rect 3278 2148 3279 2152
rect 3283 2148 3284 2152
rect 3278 2147 3284 2148
rect 3366 2152 3372 2153
rect 3366 2148 3367 2152
rect 3371 2148 3372 2152
rect 3366 2147 3372 2148
rect 3462 2149 3468 2150
rect 1806 2144 1812 2145
rect 3462 2145 3463 2149
rect 3467 2145 3468 2149
rect 3462 2144 3468 2145
rect 134 2140 140 2141
rect 110 2137 116 2138
rect 110 2133 111 2137
rect 115 2133 116 2137
rect 134 2136 135 2140
rect 139 2136 140 2140
rect 134 2135 140 2136
rect 246 2140 252 2141
rect 246 2136 247 2140
rect 251 2136 252 2140
rect 246 2135 252 2136
rect 390 2140 396 2141
rect 390 2136 391 2140
rect 395 2136 396 2140
rect 390 2135 396 2136
rect 542 2140 548 2141
rect 542 2136 543 2140
rect 547 2136 548 2140
rect 542 2135 548 2136
rect 694 2140 700 2141
rect 694 2136 695 2140
rect 699 2136 700 2140
rect 694 2135 700 2136
rect 838 2140 844 2141
rect 838 2136 839 2140
rect 843 2136 844 2140
rect 838 2135 844 2136
rect 974 2140 980 2141
rect 974 2136 975 2140
rect 979 2136 980 2140
rect 974 2135 980 2136
rect 1102 2140 1108 2141
rect 1102 2136 1103 2140
rect 1107 2136 1108 2140
rect 1102 2135 1108 2136
rect 1230 2140 1236 2141
rect 1230 2136 1231 2140
rect 1235 2136 1236 2140
rect 1230 2135 1236 2136
rect 1350 2140 1356 2141
rect 1350 2136 1351 2140
rect 1355 2136 1356 2140
rect 1350 2135 1356 2136
rect 1462 2140 1468 2141
rect 1462 2136 1463 2140
rect 1467 2136 1468 2140
rect 1462 2135 1468 2136
rect 1574 2140 1580 2141
rect 1574 2136 1575 2140
rect 1579 2136 1580 2140
rect 1574 2135 1580 2136
rect 1670 2140 1676 2141
rect 1670 2136 1671 2140
rect 1675 2136 1676 2140
rect 1670 2135 1676 2136
rect 1766 2137 1772 2138
rect 110 2132 116 2133
rect 1766 2133 1767 2137
rect 1771 2133 1772 2137
rect 2926 2133 2932 2134
rect 1766 2132 1772 2133
rect 1806 2132 1812 2133
rect 1806 2128 1807 2132
rect 1811 2128 1812 2132
rect 2926 2129 2927 2133
rect 2931 2129 2932 2133
rect 2926 2128 2932 2129
rect 3014 2133 3020 2134
rect 3014 2129 3015 2133
rect 3019 2129 3020 2133
rect 3014 2128 3020 2129
rect 3102 2133 3108 2134
rect 3102 2129 3103 2133
rect 3107 2129 3108 2133
rect 3102 2128 3108 2129
rect 3190 2133 3196 2134
rect 3190 2129 3191 2133
rect 3195 2129 3196 2133
rect 3190 2128 3196 2129
rect 3278 2133 3284 2134
rect 3278 2129 3279 2133
rect 3283 2129 3284 2133
rect 3278 2128 3284 2129
rect 3366 2133 3372 2134
rect 3366 2129 3367 2133
rect 3371 2129 3372 2133
rect 3366 2128 3372 2129
rect 3462 2132 3468 2133
rect 3462 2128 3463 2132
rect 3467 2128 3468 2132
rect 1806 2127 1812 2128
rect 3462 2127 3468 2128
rect 134 2121 140 2122
rect 110 2120 116 2121
rect 110 2116 111 2120
rect 115 2116 116 2120
rect 134 2117 135 2121
rect 139 2117 140 2121
rect 134 2116 140 2117
rect 246 2121 252 2122
rect 246 2117 247 2121
rect 251 2117 252 2121
rect 246 2116 252 2117
rect 390 2121 396 2122
rect 390 2117 391 2121
rect 395 2117 396 2121
rect 390 2116 396 2117
rect 542 2121 548 2122
rect 542 2117 543 2121
rect 547 2117 548 2121
rect 542 2116 548 2117
rect 694 2121 700 2122
rect 694 2117 695 2121
rect 699 2117 700 2121
rect 694 2116 700 2117
rect 838 2121 844 2122
rect 838 2117 839 2121
rect 843 2117 844 2121
rect 838 2116 844 2117
rect 974 2121 980 2122
rect 974 2117 975 2121
rect 979 2117 980 2121
rect 974 2116 980 2117
rect 1102 2121 1108 2122
rect 1102 2117 1103 2121
rect 1107 2117 1108 2121
rect 1102 2116 1108 2117
rect 1230 2121 1236 2122
rect 1230 2117 1231 2121
rect 1235 2117 1236 2121
rect 1230 2116 1236 2117
rect 1350 2121 1356 2122
rect 1350 2117 1351 2121
rect 1355 2117 1356 2121
rect 1350 2116 1356 2117
rect 1462 2121 1468 2122
rect 1462 2117 1463 2121
rect 1467 2117 1468 2121
rect 1462 2116 1468 2117
rect 1574 2121 1580 2122
rect 1574 2117 1575 2121
rect 1579 2117 1580 2121
rect 1574 2116 1580 2117
rect 1670 2121 1676 2122
rect 1670 2117 1671 2121
rect 1675 2117 1676 2121
rect 1670 2116 1676 2117
rect 1766 2120 1772 2121
rect 1766 2116 1767 2120
rect 1771 2116 1772 2120
rect 110 2115 116 2116
rect 1766 2115 1772 2116
rect 1806 2080 1812 2081
rect 3462 2080 3468 2081
rect 1806 2076 1807 2080
rect 1811 2076 1812 2080
rect 1806 2075 1812 2076
rect 1830 2079 1836 2080
rect 1830 2075 1831 2079
rect 1835 2075 1836 2079
rect 1830 2074 1836 2075
rect 1990 2079 1996 2080
rect 1990 2075 1991 2079
rect 1995 2075 1996 2079
rect 1990 2074 1996 2075
rect 2166 2079 2172 2080
rect 2166 2075 2167 2079
rect 2171 2075 2172 2079
rect 2166 2074 2172 2075
rect 2342 2079 2348 2080
rect 2342 2075 2343 2079
rect 2347 2075 2348 2079
rect 2342 2074 2348 2075
rect 2502 2079 2508 2080
rect 2502 2075 2503 2079
rect 2507 2075 2508 2079
rect 2502 2074 2508 2075
rect 2654 2079 2660 2080
rect 2654 2075 2655 2079
rect 2659 2075 2660 2079
rect 2654 2074 2660 2075
rect 2790 2079 2796 2080
rect 2790 2075 2791 2079
rect 2795 2075 2796 2079
rect 2790 2074 2796 2075
rect 2918 2079 2924 2080
rect 2918 2075 2919 2079
rect 2923 2075 2924 2079
rect 2918 2074 2924 2075
rect 3038 2079 3044 2080
rect 3038 2075 3039 2079
rect 3043 2075 3044 2079
rect 3038 2074 3044 2075
rect 3158 2079 3164 2080
rect 3158 2075 3159 2079
rect 3163 2075 3164 2079
rect 3158 2074 3164 2075
rect 3270 2079 3276 2080
rect 3270 2075 3271 2079
rect 3275 2075 3276 2079
rect 3270 2074 3276 2075
rect 3366 2079 3372 2080
rect 3366 2075 3367 2079
rect 3371 2075 3372 2079
rect 3462 2076 3463 2080
rect 3467 2076 3468 2080
rect 3462 2075 3468 2076
rect 3366 2074 3372 2075
rect 110 2072 116 2073
rect 1766 2072 1772 2073
rect 110 2068 111 2072
rect 115 2068 116 2072
rect 110 2067 116 2068
rect 134 2071 140 2072
rect 134 2067 135 2071
rect 139 2067 140 2071
rect 134 2066 140 2067
rect 222 2071 228 2072
rect 222 2067 223 2071
rect 227 2067 228 2071
rect 222 2066 228 2067
rect 342 2071 348 2072
rect 342 2067 343 2071
rect 347 2067 348 2071
rect 342 2066 348 2067
rect 462 2071 468 2072
rect 462 2067 463 2071
rect 467 2067 468 2071
rect 462 2066 468 2067
rect 582 2071 588 2072
rect 582 2067 583 2071
rect 587 2067 588 2071
rect 582 2066 588 2067
rect 702 2071 708 2072
rect 702 2067 703 2071
rect 707 2067 708 2071
rect 702 2066 708 2067
rect 822 2071 828 2072
rect 822 2067 823 2071
rect 827 2067 828 2071
rect 822 2066 828 2067
rect 934 2071 940 2072
rect 934 2067 935 2071
rect 939 2067 940 2071
rect 934 2066 940 2067
rect 1046 2071 1052 2072
rect 1046 2067 1047 2071
rect 1051 2067 1052 2071
rect 1046 2066 1052 2067
rect 1158 2071 1164 2072
rect 1158 2067 1159 2071
rect 1163 2067 1164 2071
rect 1158 2066 1164 2067
rect 1278 2071 1284 2072
rect 1278 2067 1279 2071
rect 1283 2067 1284 2071
rect 1766 2068 1767 2072
rect 1771 2068 1772 2072
rect 1766 2067 1772 2068
rect 1278 2066 1284 2067
rect 1806 2063 1812 2064
rect 1806 2059 1807 2063
rect 1811 2059 1812 2063
rect 3462 2063 3468 2064
rect 1806 2058 1812 2059
rect 1830 2060 1836 2061
rect 1830 2056 1831 2060
rect 1835 2056 1836 2060
rect 110 2055 116 2056
rect 110 2051 111 2055
rect 115 2051 116 2055
rect 1766 2055 1772 2056
rect 1830 2055 1836 2056
rect 1990 2060 1996 2061
rect 1990 2056 1991 2060
rect 1995 2056 1996 2060
rect 1990 2055 1996 2056
rect 2166 2060 2172 2061
rect 2166 2056 2167 2060
rect 2171 2056 2172 2060
rect 2166 2055 2172 2056
rect 2342 2060 2348 2061
rect 2342 2056 2343 2060
rect 2347 2056 2348 2060
rect 2342 2055 2348 2056
rect 2502 2060 2508 2061
rect 2502 2056 2503 2060
rect 2507 2056 2508 2060
rect 2502 2055 2508 2056
rect 2654 2060 2660 2061
rect 2654 2056 2655 2060
rect 2659 2056 2660 2060
rect 2654 2055 2660 2056
rect 2790 2060 2796 2061
rect 2790 2056 2791 2060
rect 2795 2056 2796 2060
rect 2790 2055 2796 2056
rect 2918 2060 2924 2061
rect 2918 2056 2919 2060
rect 2923 2056 2924 2060
rect 2918 2055 2924 2056
rect 3038 2060 3044 2061
rect 3038 2056 3039 2060
rect 3043 2056 3044 2060
rect 3038 2055 3044 2056
rect 3158 2060 3164 2061
rect 3158 2056 3159 2060
rect 3163 2056 3164 2060
rect 3158 2055 3164 2056
rect 3270 2060 3276 2061
rect 3270 2056 3271 2060
rect 3275 2056 3276 2060
rect 3270 2055 3276 2056
rect 3366 2060 3372 2061
rect 3366 2056 3367 2060
rect 3371 2056 3372 2060
rect 3462 2059 3463 2063
rect 3467 2059 3468 2063
rect 3462 2058 3468 2059
rect 3366 2055 3372 2056
rect 110 2050 116 2051
rect 134 2052 140 2053
rect 134 2048 135 2052
rect 139 2048 140 2052
rect 134 2047 140 2048
rect 222 2052 228 2053
rect 222 2048 223 2052
rect 227 2048 228 2052
rect 222 2047 228 2048
rect 342 2052 348 2053
rect 342 2048 343 2052
rect 347 2048 348 2052
rect 342 2047 348 2048
rect 462 2052 468 2053
rect 462 2048 463 2052
rect 467 2048 468 2052
rect 462 2047 468 2048
rect 582 2052 588 2053
rect 582 2048 583 2052
rect 587 2048 588 2052
rect 582 2047 588 2048
rect 702 2052 708 2053
rect 702 2048 703 2052
rect 707 2048 708 2052
rect 702 2047 708 2048
rect 822 2052 828 2053
rect 822 2048 823 2052
rect 827 2048 828 2052
rect 822 2047 828 2048
rect 934 2052 940 2053
rect 934 2048 935 2052
rect 939 2048 940 2052
rect 934 2047 940 2048
rect 1046 2052 1052 2053
rect 1046 2048 1047 2052
rect 1051 2048 1052 2052
rect 1046 2047 1052 2048
rect 1158 2052 1164 2053
rect 1158 2048 1159 2052
rect 1163 2048 1164 2052
rect 1158 2047 1164 2048
rect 1278 2052 1284 2053
rect 1278 2048 1279 2052
rect 1283 2048 1284 2052
rect 1766 2051 1767 2055
rect 1771 2051 1772 2055
rect 1766 2050 1772 2051
rect 1278 2047 1284 2048
rect 1830 2012 1836 2013
rect 1806 2009 1812 2010
rect 1806 2005 1807 2009
rect 1811 2005 1812 2009
rect 1830 2008 1831 2012
rect 1835 2008 1836 2012
rect 1830 2007 1836 2008
rect 2014 2012 2020 2013
rect 2014 2008 2015 2012
rect 2019 2008 2020 2012
rect 2014 2007 2020 2008
rect 2222 2012 2228 2013
rect 2222 2008 2223 2012
rect 2227 2008 2228 2012
rect 2222 2007 2228 2008
rect 2430 2012 2436 2013
rect 2430 2008 2431 2012
rect 2435 2008 2436 2012
rect 2430 2007 2436 2008
rect 2630 2012 2636 2013
rect 2630 2008 2631 2012
rect 2635 2008 2636 2012
rect 2630 2007 2636 2008
rect 2822 2012 2828 2013
rect 2822 2008 2823 2012
rect 2827 2008 2828 2012
rect 2822 2007 2828 2008
rect 3006 2012 3012 2013
rect 3006 2008 3007 2012
rect 3011 2008 3012 2012
rect 3006 2007 3012 2008
rect 3198 2012 3204 2013
rect 3198 2008 3199 2012
rect 3203 2008 3204 2012
rect 3198 2007 3204 2008
rect 3366 2012 3372 2013
rect 3366 2008 3367 2012
rect 3371 2008 3372 2012
rect 3366 2007 3372 2008
rect 3462 2009 3468 2010
rect 1806 2004 1812 2005
rect 3462 2005 3463 2009
rect 3467 2005 3468 2009
rect 3462 2004 3468 2005
rect 134 2000 140 2001
rect 110 1997 116 1998
rect 110 1993 111 1997
rect 115 1993 116 1997
rect 134 1996 135 2000
rect 139 1996 140 2000
rect 134 1995 140 1996
rect 238 2000 244 2001
rect 238 1996 239 2000
rect 243 1996 244 2000
rect 238 1995 244 1996
rect 366 2000 372 2001
rect 366 1996 367 2000
rect 371 1996 372 2000
rect 366 1995 372 1996
rect 502 2000 508 2001
rect 502 1996 503 2000
rect 507 1996 508 2000
rect 502 1995 508 1996
rect 638 2000 644 2001
rect 638 1996 639 2000
rect 643 1996 644 2000
rect 638 1995 644 1996
rect 774 2000 780 2001
rect 774 1996 775 2000
rect 779 1996 780 2000
rect 774 1995 780 1996
rect 910 2000 916 2001
rect 910 1996 911 2000
rect 915 1996 916 2000
rect 910 1995 916 1996
rect 1046 2000 1052 2001
rect 1046 1996 1047 2000
rect 1051 1996 1052 2000
rect 1046 1995 1052 1996
rect 1182 2000 1188 2001
rect 1182 1996 1183 2000
rect 1187 1996 1188 2000
rect 1182 1995 1188 1996
rect 1326 2000 1332 2001
rect 1326 1996 1327 2000
rect 1331 1996 1332 2000
rect 1326 1995 1332 1996
rect 1766 1997 1772 1998
rect 110 1992 116 1993
rect 1766 1993 1767 1997
rect 1771 1993 1772 1997
rect 1830 1993 1836 1994
rect 1766 1992 1772 1993
rect 1806 1992 1812 1993
rect 1806 1988 1807 1992
rect 1811 1988 1812 1992
rect 1830 1989 1831 1993
rect 1835 1989 1836 1993
rect 1830 1988 1836 1989
rect 2014 1993 2020 1994
rect 2014 1989 2015 1993
rect 2019 1989 2020 1993
rect 2014 1988 2020 1989
rect 2222 1993 2228 1994
rect 2222 1989 2223 1993
rect 2227 1989 2228 1993
rect 2222 1988 2228 1989
rect 2430 1993 2436 1994
rect 2430 1989 2431 1993
rect 2435 1989 2436 1993
rect 2430 1988 2436 1989
rect 2630 1993 2636 1994
rect 2630 1989 2631 1993
rect 2635 1989 2636 1993
rect 2630 1988 2636 1989
rect 2822 1993 2828 1994
rect 2822 1989 2823 1993
rect 2827 1989 2828 1993
rect 2822 1988 2828 1989
rect 3006 1993 3012 1994
rect 3006 1989 3007 1993
rect 3011 1989 3012 1993
rect 3006 1988 3012 1989
rect 3198 1993 3204 1994
rect 3198 1989 3199 1993
rect 3203 1989 3204 1993
rect 3198 1988 3204 1989
rect 3366 1993 3372 1994
rect 3366 1989 3367 1993
rect 3371 1989 3372 1993
rect 3366 1988 3372 1989
rect 3462 1992 3468 1993
rect 3462 1988 3463 1992
rect 3467 1988 3468 1992
rect 1806 1987 1812 1988
rect 3462 1987 3468 1988
rect 134 1981 140 1982
rect 110 1980 116 1981
rect 110 1976 111 1980
rect 115 1976 116 1980
rect 134 1977 135 1981
rect 139 1977 140 1981
rect 134 1976 140 1977
rect 238 1981 244 1982
rect 238 1977 239 1981
rect 243 1977 244 1981
rect 238 1976 244 1977
rect 366 1981 372 1982
rect 366 1977 367 1981
rect 371 1977 372 1981
rect 366 1976 372 1977
rect 502 1981 508 1982
rect 502 1977 503 1981
rect 507 1977 508 1981
rect 502 1976 508 1977
rect 638 1981 644 1982
rect 638 1977 639 1981
rect 643 1977 644 1981
rect 638 1976 644 1977
rect 774 1981 780 1982
rect 774 1977 775 1981
rect 779 1977 780 1981
rect 774 1976 780 1977
rect 910 1981 916 1982
rect 910 1977 911 1981
rect 915 1977 916 1981
rect 910 1976 916 1977
rect 1046 1981 1052 1982
rect 1046 1977 1047 1981
rect 1051 1977 1052 1981
rect 1046 1976 1052 1977
rect 1182 1981 1188 1982
rect 1182 1977 1183 1981
rect 1187 1977 1188 1981
rect 1182 1976 1188 1977
rect 1326 1981 1332 1982
rect 1326 1977 1327 1981
rect 1331 1977 1332 1981
rect 1326 1976 1332 1977
rect 1766 1980 1772 1981
rect 1766 1976 1767 1980
rect 1771 1976 1772 1980
rect 110 1975 116 1976
rect 1766 1975 1772 1976
rect 1806 1944 1812 1945
rect 3462 1944 3468 1945
rect 1806 1940 1807 1944
rect 1811 1940 1812 1944
rect 1806 1939 1812 1940
rect 1862 1943 1868 1944
rect 1862 1939 1863 1943
rect 1867 1939 1868 1943
rect 1862 1938 1868 1939
rect 1998 1943 2004 1944
rect 1998 1939 1999 1943
rect 2003 1939 2004 1943
rect 1998 1938 2004 1939
rect 2142 1943 2148 1944
rect 2142 1939 2143 1943
rect 2147 1939 2148 1943
rect 2142 1938 2148 1939
rect 2286 1943 2292 1944
rect 2286 1939 2287 1943
rect 2291 1939 2292 1943
rect 2286 1938 2292 1939
rect 2430 1943 2436 1944
rect 2430 1939 2431 1943
rect 2435 1939 2436 1943
rect 2430 1938 2436 1939
rect 2574 1943 2580 1944
rect 2574 1939 2575 1943
rect 2579 1939 2580 1943
rect 2574 1938 2580 1939
rect 2710 1943 2716 1944
rect 2710 1939 2711 1943
rect 2715 1939 2716 1943
rect 2710 1938 2716 1939
rect 2830 1943 2836 1944
rect 2830 1939 2831 1943
rect 2835 1939 2836 1943
rect 2830 1938 2836 1939
rect 2950 1943 2956 1944
rect 2950 1939 2951 1943
rect 2955 1939 2956 1943
rect 2950 1938 2956 1939
rect 3062 1943 3068 1944
rect 3062 1939 3063 1943
rect 3067 1939 3068 1943
rect 3062 1938 3068 1939
rect 3166 1943 3172 1944
rect 3166 1939 3167 1943
rect 3171 1939 3172 1943
rect 3166 1938 3172 1939
rect 3278 1943 3284 1944
rect 3278 1939 3279 1943
rect 3283 1939 3284 1943
rect 3278 1938 3284 1939
rect 3366 1943 3372 1944
rect 3366 1939 3367 1943
rect 3371 1939 3372 1943
rect 3462 1940 3463 1944
rect 3467 1940 3468 1944
rect 3462 1939 3468 1940
rect 3366 1938 3372 1939
rect 110 1932 116 1933
rect 1766 1932 1772 1933
rect 110 1928 111 1932
rect 115 1928 116 1932
rect 110 1927 116 1928
rect 294 1931 300 1932
rect 294 1927 295 1931
rect 299 1927 300 1931
rect 294 1926 300 1927
rect 422 1931 428 1932
rect 422 1927 423 1931
rect 427 1927 428 1931
rect 422 1926 428 1927
rect 558 1931 564 1932
rect 558 1927 559 1931
rect 563 1927 564 1931
rect 558 1926 564 1927
rect 702 1931 708 1932
rect 702 1927 703 1931
rect 707 1927 708 1931
rect 702 1926 708 1927
rect 854 1931 860 1932
rect 854 1927 855 1931
rect 859 1927 860 1931
rect 854 1926 860 1927
rect 1006 1931 1012 1932
rect 1006 1927 1007 1931
rect 1011 1927 1012 1931
rect 1006 1926 1012 1927
rect 1158 1931 1164 1932
rect 1158 1927 1159 1931
rect 1163 1927 1164 1931
rect 1158 1926 1164 1927
rect 1310 1931 1316 1932
rect 1310 1927 1311 1931
rect 1315 1927 1316 1931
rect 1310 1926 1316 1927
rect 1470 1931 1476 1932
rect 1470 1927 1471 1931
rect 1475 1927 1476 1931
rect 1766 1928 1767 1932
rect 1771 1928 1772 1932
rect 1766 1927 1772 1928
rect 1806 1927 1812 1928
rect 1470 1926 1476 1927
rect 1806 1923 1807 1927
rect 1811 1923 1812 1927
rect 3462 1927 3468 1928
rect 1806 1922 1812 1923
rect 1862 1924 1868 1925
rect 1862 1920 1863 1924
rect 1867 1920 1868 1924
rect 1862 1919 1868 1920
rect 1998 1924 2004 1925
rect 1998 1920 1999 1924
rect 2003 1920 2004 1924
rect 1998 1919 2004 1920
rect 2142 1924 2148 1925
rect 2142 1920 2143 1924
rect 2147 1920 2148 1924
rect 2142 1919 2148 1920
rect 2286 1924 2292 1925
rect 2286 1920 2287 1924
rect 2291 1920 2292 1924
rect 2286 1919 2292 1920
rect 2430 1924 2436 1925
rect 2430 1920 2431 1924
rect 2435 1920 2436 1924
rect 2430 1919 2436 1920
rect 2574 1924 2580 1925
rect 2574 1920 2575 1924
rect 2579 1920 2580 1924
rect 2574 1919 2580 1920
rect 2710 1924 2716 1925
rect 2710 1920 2711 1924
rect 2715 1920 2716 1924
rect 2710 1919 2716 1920
rect 2830 1924 2836 1925
rect 2830 1920 2831 1924
rect 2835 1920 2836 1924
rect 2830 1919 2836 1920
rect 2950 1924 2956 1925
rect 2950 1920 2951 1924
rect 2955 1920 2956 1924
rect 2950 1919 2956 1920
rect 3062 1924 3068 1925
rect 3062 1920 3063 1924
rect 3067 1920 3068 1924
rect 3062 1919 3068 1920
rect 3166 1924 3172 1925
rect 3166 1920 3167 1924
rect 3171 1920 3172 1924
rect 3166 1919 3172 1920
rect 3278 1924 3284 1925
rect 3278 1920 3279 1924
rect 3283 1920 3284 1924
rect 3278 1919 3284 1920
rect 3366 1924 3372 1925
rect 3366 1920 3367 1924
rect 3371 1920 3372 1924
rect 3462 1923 3463 1927
rect 3467 1923 3468 1927
rect 3462 1922 3468 1923
rect 3366 1919 3372 1920
rect 110 1915 116 1916
rect 110 1911 111 1915
rect 115 1911 116 1915
rect 1766 1915 1772 1916
rect 110 1910 116 1911
rect 294 1912 300 1913
rect 294 1908 295 1912
rect 299 1908 300 1912
rect 294 1907 300 1908
rect 422 1912 428 1913
rect 422 1908 423 1912
rect 427 1908 428 1912
rect 422 1907 428 1908
rect 558 1912 564 1913
rect 558 1908 559 1912
rect 563 1908 564 1912
rect 558 1907 564 1908
rect 702 1912 708 1913
rect 702 1908 703 1912
rect 707 1908 708 1912
rect 702 1907 708 1908
rect 854 1912 860 1913
rect 854 1908 855 1912
rect 859 1908 860 1912
rect 854 1907 860 1908
rect 1006 1912 1012 1913
rect 1006 1908 1007 1912
rect 1011 1908 1012 1912
rect 1006 1907 1012 1908
rect 1158 1912 1164 1913
rect 1158 1908 1159 1912
rect 1163 1908 1164 1912
rect 1158 1907 1164 1908
rect 1310 1912 1316 1913
rect 1310 1908 1311 1912
rect 1315 1908 1316 1912
rect 1310 1907 1316 1908
rect 1470 1912 1476 1913
rect 1470 1908 1471 1912
rect 1475 1908 1476 1912
rect 1766 1911 1767 1915
rect 1771 1911 1772 1915
rect 1766 1910 1772 1911
rect 1470 1907 1476 1908
rect 2014 1876 2020 1877
rect 1806 1873 1812 1874
rect 1806 1869 1807 1873
rect 1811 1869 1812 1873
rect 2014 1872 2015 1876
rect 2019 1872 2020 1876
rect 2014 1871 2020 1872
rect 2110 1876 2116 1877
rect 2110 1872 2111 1876
rect 2115 1872 2116 1876
rect 2110 1871 2116 1872
rect 2214 1876 2220 1877
rect 2214 1872 2215 1876
rect 2219 1872 2220 1876
rect 2214 1871 2220 1872
rect 2326 1876 2332 1877
rect 2326 1872 2327 1876
rect 2331 1872 2332 1876
rect 2326 1871 2332 1872
rect 2438 1876 2444 1877
rect 2438 1872 2439 1876
rect 2443 1872 2444 1876
rect 2438 1871 2444 1872
rect 2542 1876 2548 1877
rect 2542 1872 2543 1876
rect 2547 1872 2548 1876
rect 2542 1871 2548 1872
rect 2646 1876 2652 1877
rect 2646 1872 2647 1876
rect 2651 1872 2652 1876
rect 2646 1871 2652 1872
rect 2758 1876 2764 1877
rect 2758 1872 2759 1876
rect 2763 1872 2764 1876
rect 2758 1871 2764 1872
rect 2870 1876 2876 1877
rect 2870 1872 2871 1876
rect 2875 1872 2876 1876
rect 2870 1871 2876 1872
rect 2982 1876 2988 1877
rect 2982 1872 2983 1876
rect 2987 1872 2988 1876
rect 2982 1871 2988 1872
rect 3462 1873 3468 1874
rect 430 1868 436 1869
rect 110 1865 116 1866
rect 110 1861 111 1865
rect 115 1861 116 1865
rect 430 1864 431 1868
rect 435 1864 436 1868
rect 430 1863 436 1864
rect 574 1868 580 1869
rect 574 1864 575 1868
rect 579 1864 580 1868
rect 574 1863 580 1864
rect 726 1868 732 1869
rect 726 1864 727 1868
rect 731 1864 732 1868
rect 726 1863 732 1864
rect 886 1868 892 1869
rect 886 1864 887 1868
rect 891 1864 892 1868
rect 886 1863 892 1864
rect 1046 1868 1052 1869
rect 1046 1864 1047 1868
rect 1051 1864 1052 1868
rect 1046 1863 1052 1864
rect 1198 1868 1204 1869
rect 1198 1864 1199 1868
rect 1203 1864 1204 1868
rect 1198 1863 1204 1864
rect 1350 1868 1356 1869
rect 1350 1864 1351 1868
rect 1355 1864 1356 1868
rect 1350 1863 1356 1864
rect 1510 1868 1516 1869
rect 1510 1864 1511 1868
rect 1515 1864 1516 1868
rect 1510 1863 1516 1864
rect 1670 1868 1676 1869
rect 1806 1868 1812 1869
rect 3462 1869 3463 1873
rect 3467 1869 3468 1873
rect 3462 1868 3468 1869
rect 1670 1864 1671 1868
rect 1675 1864 1676 1868
rect 1670 1863 1676 1864
rect 1766 1865 1772 1866
rect 110 1860 116 1861
rect 1766 1861 1767 1865
rect 1771 1861 1772 1865
rect 1766 1860 1772 1861
rect 2014 1857 2020 1858
rect 1806 1856 1812 1857
rect 1806 1852 1807 1856
rect 1811 1852 1812 1856
rect 2014 1853 2015 1857
rect 2019 1853 2020 1857
rect 2014 1852 2020 1853
rect 2110 1857 2116 1858
rect 2110 1853 2111 1857
rect 2115 1853 2116 1857
rect 2110 1852 2116 1853
rect 2214 1857 2220 1858
rect 2214 1853 2215 1857
rect 2219 1853 2220 1857
rect 2214 1852 2220 1853
rect 2326 1857 2332 1858
rect 2326 1853 2327 1857
rect 2331 1853 2332 1857
rect 2326 1852 2332 1853
rect 2438 1857 2444 1858
rect 2438 1853 2439 1857
rect 2443 1853 2444 1857
rect 2438 1852 2444 1853
rect 2542 1857 2548 1858
rect 2542 1853 2543 1857
rect 2547 1853 2548 1857
rect 2542 1852 2548 1853
rect 2646 1857 2652 1858
rect 2646 1853 2647 1857
rect 2651 1853 2652 1857
rect 2646 1852 2652 1853
rect 2758 1857 2764 1858
rect 2758 1853 2759 1857
rect 2763 1853 2764 1857
rect 2758 1852 2764 1853
rect 2870 1857 2876 1858
rect 2870 1853 2871 1857
rect 2875 1853 2876 1857
rect 2870 1852 2876 1853
rect 2982 1857 2988 1858
rect 2982 1853 2983 1857
rect 2987 1853 2988 1857
rect 2982 1852 2988 1853
rect 3462 1856 3468 1857
rect 3462 1852 3463 1856
rect 3467 1852 3468 1856
rect 1806 1851 1812 1852
rect 3462 1851 3468 1852
rect 430 1849 436 1850
rect 110 1848 116 1849
rect 110 1844 111 1848
rect 115 1844 116 1848
rect 430 1845 431 1849
rect 435 1845 436 1849
rect 430 1844 436 1845
rect 574 1849 580 1850
rect 574 1845 575 1849
rect 579 1845 580 1849
rect 574 1844 580 1845
rect 726 1849 732 1850
rect 726 1845 727 1849
rect 731 1845 732 1849
rect 726 1844 732 1845
rect 886 1849 892 1850
rect 886 1845 887 1849
rect 891 1845 892 1849
rect 886 1844 892 1845
rect 1046 1849 1052 1850
rect 1046 1845 1047 1849
rect 1051 1845 1052 1849
rect 1046 1844 1052 1845
rect 1198 1849 1204 1850
rect 1198 1845 1199 1849
rect 1203 1845 1204 1849
rect 1198 1844 1204 1845
rect 1350 1849 1356 1850
rect 1350 1845 1351 1849
rect 1355 1845 1356 1849
rect 1350 1844 1356 1845
rect 1510 1849 1516 1850
rect 1510 1845 1511 1849
rect 1515 1845 1516 1849
rect 1510 1844 1516 1845
rect 1670 1849 1676 1850
rect 1670 1845 1671 1849
rect 1675 1845 1676 1849
rect 1670 1844 1676 1845
rect 1766 1848 1772 1849
rect 1766 1844 1767 1848
rect 1771 1844 1772 1848
rect 110 1843 116 1844
rect 1766 1843 1772 1844
rect 1806 1804 1812 1805
rect 3462 1804 3468 1805
rect 110 1800 116 1801
rect 1766 1800 1772 1801
rect 110 1796 111 1800
rect 115 1796 116 1800
rect 110 1795 116 1796
rect 510 1799 516 1800
rect 510 1795 511 1799
rect 515 1795 516 1799
rect 510 1794 516 1795
rect 630 1799 636 1800
rect 630 1795 631 1799
rect 635 1795 636 1799
rect 630 1794 636 1795
rect 758 1799 764 1800
rect 758 1795 759 1799
rect 763 1795 764 1799
rect 758 1794 764 1795
rect 886 1799 892 1800
rect 886 1795 887 1799
rect 891 1795 892 1799
rect 886 1794 892 1795
rect 1022 1799 1028 1800
rect 1022 1795 1023 1799
rect 1027 1795 1028 1799
rect 1022 1794 1028 1795
rect 1150 1799 1156 1800
rect 1150 1795 1151 1799
rect 1155 1795 1156 1799
rect 1150 1794 1156 1795
rect 1278 1799 1284 1800
rect 1278 1795 1279 1799
rect 1283 1795 1284 1799
rect 1278 1794 1284 1795
rect 1406 1799 1412 1800
rect 1406 1795 1407 1799
rect 1411 1795 1412 1799
rect 1406 1794 1412 1795
rect 1534 1799 1540 1800
rect 1534 1795 1535 1799
rect 1539 1795 1540 1799
rect 1534 1794 1540 1795
rect 1670 1799 1676 1800
rect 1670 1795 1671 1799
rect 1675 1795 1676 1799
rect 1766 1796 1767 1800
rect 1771 1796 1772 1800
rect 1806 1800 1807 1804
rect 1811 1800 1812 1804
rect 1806 1799 1812 1800
rect 2102 1803 2108 1804
rect 2102 1799 2103 1803
rect 2107 1799 2108 1803
rect 2102 1798 2108 1799
rect 2190 1803 2196 1804
rect 2190 1799 2191 1803
rect 2195 1799 2196 1803
rect 2190 1798 2196 1799
rect 2278 1803 2284 1804
rect 2278 1799 2279 1803
rect 2283 1799 2284 1803
rect 2278 1798 2284 1799
rect 2366 1803 2372 1804
rect 2366 1799 2367 1803
rect 2371 1799 2372 1803
rect 2366 1798 2372 1799
rect 2454 1803 2460 1804
rect 2454 1799 2455 1803
rect 2459 1799 2460 1803
rect 2454 1798 2460 1799
rect 2542 1803 2548 1804
rect 2542 1799 2543 1803
rect 2547 1799 2548 1803
rect 2542 1798 2548 1799
rect 2630 1803 2636 1804
rect 2630 1799 2631 1803
rect 2635 1799 2636 1803
rect 2630 1798 2636 1799
rect 2718 1803 2724 1804
rect 2718 1799 2719 1803
rect 2723 1799 2724 1803
rect 2718 1798 2724 1799
rect 2806 1803 2812 1804
rect 2806 1799 2807 1803
rect 2811 1799 2812 1803
rect 2806 1798 2812 1799
rect 2894 1803 2900 1804
rect 2894 1799 2895 1803
rect 2899 1799 2900 1803
rect 3462 1800 3463 1804
rect 3467 1800 3468 1804
rect 3462 1799 3468 1800
rect 2894 1798 2900 1799
rect 1766 1795 1772 1796
rect 1670 1794 1676 1795
rect 1806 1787 1812 1788
rect 110 1783 116 1784
rect 110 1779 111 1783
rect 115 1779 116 1783
rect 1766 1783 1772 1784
rect 110 1778 116 1779
rect 510 1780 516 1781
rect 510 1776 511 1780
rect 515 1776 516 1780
rect 510 1775 516 1776
rect 630 1780 636 1781
rect 630 1776 631 1780
rect 635 1776 636 1780
rect 630 1775 636 1776
rect 758 1780 764 1781
rect 758 1776 759 1780
rect 763 1776 764 1780
rect 758 1775 764 1776
rect 886 1780 892 1781
rect 886 1776 887 1780
rect 891 1776 892 1780
rect 886 1775 892 1776
rect 1022 1780 1028 1781
rect 1022 1776 1023 1780
rect 1027 1776 1028 1780
rect 1022 1775 1028 1776
rect 1150 1780 1156 1781
rect 1150 1776 1151 1780
rect 1155 1776 1156 1780
rect 1150 1775 1156 1776
rect 1278 1780 1284 1781
rect 1278 1776 1279 1780
rect 1283 1776 1284 1780
rect 1278 1775 1284 1776
rect 1406 1780 1412 1781
rect 1406 1776 1407 1780
rect 1411 1776 1412 1780
rect 1406 1775 1412 1776
rect 1534 1780 1540 1781
rect 1534 1776 1535 1780
rect 1539 1776 1540 1780
rect 1534 1775 1540 1776
rect 1670 1780 1676 1781
rect 1670 1776 1671 1780
rect 1675 1776 1676 1780
rect 1766 1779 1767 1783
rect 1771 1779 1772 1783
rect 1806 1783 1807 1787
rect 1811 1783 1812 1787
rect 3462 1787 3468 1788
rect 1806 1782 1812 1783
rect 2102 1784 2108 1785
rect 2102 1780 2103 1784
rect 2107 1780 2108 1784
rect 2102 1779 2108 1780
rect 2190 1784 2196 1785
rect 2190 1780 2191 1784
rect 2195 1780 2196 1784
rect 2190 1779 2196 1780
rect 2278 1784 2284 1785
rect 2278 1780 2279 1784
rect 2283 1780 2284 1784
rect 2278 1779 2284 1780
rect 2366 1784 2372 1785
rect 2366 1780 2367 1784
rect 2371 1780 2372 1784
rect 2366 1779 2372 1780
rect 2454 1784 2460 1785
rect 2454 1780 2455 1784
rect 2459 1780 2460 1784
rect 2454 1779 2460 1780
rect 2542 1784 2548 1785
rect 2542 1780 2543 1784
rect 2547 1780 2548 1784
rect 2542 1779 2548 1780
rect 2630 1784 2636 1785
rect 2630 1780 2631 1784
rect 2635 1780 2636 1784
rect 2630 1779 2636 1780
rect 2718 1784 2724 1785
rect 2718 1780 2719 1784
rect 2723 1780 2724 1784
rect 2718 1779 2724 1780
rect 2806 1784 2812 1785
rect 2806 1780 2807 1784
rect 2811 1780 2812 1784
rect 2806 1779 2812 1780
rect 2894 1784 2900 1785
rect 2894 1780 2895 1784
rect 2899 1780 2900 1784
rect 3462 1783 3463 1787
rect 3467 1783 3468 1787
rect 3462 1782 3468 1783
rect 2894 1779 2900 1780
rect 1766 1778 1772 1779
rect 1670 1775 1676 1776
rect 438 1732 444 1733
rect 110 1729 116 1730
rect 110 1725 111 1729
rect 115 1725 116 1729
rect 438 1728 439 1732
rect 443 1728 444 1732
rect 438 1727 444 1728
rect 534 1732 540 1733
rect 534 1728 535 1732
rect 539 1728 540 1732
rect 534 1727 540 1728
rect 638 1732 644 1733
rect 638 1728 639 1732
rect 643 1728 644 1732
rect 638 1727 644 1728
rect 742 1732 748 1733
rect 742 1728 743 1732
rect 747 1728 748 1732
rect 742 1727 748 1728
rect 846 1732 852 1733
rect 846 1728 847 1732
rect 851 1728 852 1732
rect 846 1727 852 1728
rect 950 1732 956 1733
rect 950 1728 951 1732
rect 955 1728 956 1732
rect 950 1727 956 1728
rect 1054 1732 1060 1733
rect 1054 1728 1055 1732
rect 1059 1728 1060 1732
rect 1054 1727 1060 1728
rect 1158 1732 1164 1733
rect 1158 1728 1159 1732
rect 1163 1728 1164 1732
rect 1158 1727 1164 1728
rect 1270 1732 1276 1733
rect 1270 1728 1271 1732
rect 1275 1728 1276 1732
rect 1270 1727 1276 1728
rect 1382 1732 1388 1733
rect 1382 1728 1383 1732
rect 1387 1728 1388 1732
rect 1382 1727 1388 1728
rect 1766 1729 1772 1730
rect 110 1724 116 1725
rect 1766 1725 1767 1729
rect 1771 1725 1772 1729
rect 2142 1728 2148 1729
rect 1766 1724 1772 1725
rect 1806 1725 1812 1726
rect 1806 1721 1807 1725
rect 1811 1721 1812 1725
rect 2142 1724 2143 1728
rect 2147 1724 2148 1728
rect 2142 1723 2148 1724
rect 2230 1728 2236 1729
rect 2230 1724 2231 1728
rect 2235 1724 2236 1728
rect 2230 1723 2236 1724
rect 2318 1728 2324 1729
rect 2318 1724 2319 1728
rect 2323 1724 2324 1728
rect 2318 1723 2324 1724
rect 2406 1728 2412 1729
rect 2406 1724 2407 1728
rect 2411 1724 2412 1728
rect 2406 1723 2412 1724
rect 2494 1728 2500 1729
rect 2494 1724 2495 1728
rect 2499 1724 2500 1728
rect 2494 1723 2500 1724
rect 2582 1728 2588 1729
rect 2582 1724 2583 1728
rect 2587 1724 2588 1728
rect 2582 1723 2588 1724
rect 2670 1728 2676 1729
rect 2670 1724 2671 1728
rect 2675 1724 2676 1728
rect 2670 1723 2676 1724
rect 2758 1728 2764 1729
rect 2758 1724 2759 1728
rect 2763 1724 2764 1728
rect 2758 1723 2764 1724
rect 2846 1728 2852 1729
rect 2846 1724 2847 1728
rect 2851 1724 2852 1728
rect 2846 1723 2852 1724
rect 3462 1725 3468 1726
rect 1806 1720 1812 1721
rect 3462 1721 3463 1725
rect 3467 1721 3468 1725
rect 3462 1720 3468 1721
rect 438 1713 444 1714
rect 110 1712 116 1713
rect 110 1708 111 1712
rect 115 1708 116 1712
rect 438 1709 439 1713
rect 443 1709 444 1713
rect 438 1708 444 1709
rect 534 1713 540 1714
rect 534 1709 535 1713
rect 539 1709 540 1713
rect 534 1708 540 1709
rect 638 1713 644 1714
rect 638 1709 639 1713
rect 643 1709 644 1713
rect 638 1708 644 1709
rect 742 1713 748 1714
rect 742 1709 743 1713
rect 747 1709 748 1713
rect 742 1708 748 1709
rect 846 1713 852 1714
rect 846 1709 847 1713
rect 851 1709 852 1713
rect 846 1708 852 1709
rect 950 1713 956 1714
rect 950 1709 951 1713
rect 955 1709 956 1713
rect 950 1708 956 1709
rect 1054 1713 1060 1714
rect 1054 1709 1055 1713
rect 1059 1709 1060 1713
rect 1054 1708 1060 1709
rect 1158 1713 1164 1714
rect 1158 1709 1159 1713
rect 1163 1709 1164 1713
rect 1158 1708 1164 1709
rect 1270 1713 1276 1714
rect 1270 1709 1271 1713
rect 1275 1709 1276 1713
rect 1270 1708 1276 1709
rect 1382 1713 1388 1714
rect 1382 1709 1383 1713
rect 1387 1709 1388 1713
rect 1382 1708 1388 1709
rect 1766 1712 1772 1713
rect 1766 1708 1767 1712
rect 1771 1708 1772 1712
rect 2142 1709 2148 1710
rect 110 1707 116 1708
rect 1766 1707 1772 1708
rect 1806 1708 1812 1709
rect 1806 1704 1807 1708
rect 1811 1704 1812 1708
rect 2142 1705 2143 1709
rect 2147 1705 2148 1709
rect 2142 1704 2148 1705
rect 2230 1709 2236 1710
rect 2230 1705 2231 1709
rect 2235 1705 2236 1709
rect 2230 1704 2236 1705
rect 2318 1709 2324 1710
rect 2318 1705 2319 1709
rect 2323 1705 2324 1709
rect 2318 1704 2324 1705
rect 2406 1709 2412 1710
rect 2406 1705 2407 1709
rect 2411 1705 2412 1709
rect 2406 1704 2412 1705
rect 2494 1709 2500 1710
rect 2494 1705 2495 1709
rect 2499 1705 2500 1709
rect 2494 1704 2500 1705
rect 2582 1709 2588 1710
rect 2582 1705 2583 1709
rect 2587 1705 2588 1709
rect 2582 1704 2588 1705
rect 2670 1709 2676 1710
rect 2670 1705 2671 1709
rect 2675 1705 2676 1709
rect 2670 1704 2676 1705
rect 2758 1709 2764 1710
rect 2758 1705 2759 1709
rect 2763 1705 2764 1709
rect 2758 1704 2764 1705
rect 2846 1709 2852 1710
rect 2846 1705 2847 1709
rect 2851 1705 2852 1709
rect 2846 1704 2852 1705
rect 3462 1708 3468 1709
rect 3462 1704 3463 1708
rect 3467 1704 3468 1708
rect 1806 1703 1812 1704
rect 3462 1703 3468 1704
rect 110 1664 116 1665
rect 1766 1664 1772 1665
rect 110 1660 111 1664
rect 115 1660 116 1664
rect 110 1659 116 1660
rect 398 1663 404 1664
rect 398 1659 399 1663
rect 403 1659 404 1663
rect 398 1658 404 1659
rect 486 1663 492 1664
rect 486 1659 487 1663
rect 491 1659 492 1663
rect 486 1658 492 1659
rect 574 1663 580 1664
rect 574 1659 575 1663
rect 579 1659 580 1663
rect 574 1658 580 1659
rect 662 1663 668 1664
rect 662 1659 663 1663
rect 667 1659 668 1663
rect 662 1658 668 1659
rect 758 1663 764 1664
rect 758 1659 759 1663
rect 763 1659 764 1663
rect 758 1658 764 1659
rect 854 1663 860 1664
rect 854 1659 855 1663
rect 859 1659 860 1663
rect 854 1658 860 1659
rect 950 1663 956 1664
rect 950 1659 951 1663
rect 955 1659 956 1663
rect 950 1658 956 1659
rect 1046 1663 1052 1664
rect 1046 1659 1047 1663
rect 1051 1659 1052 1663
rect 1046 1658 1052 1659
rect 1142 1663 1148 1664
rect 1142 1659 1143 1663
rect 1147 1659 1148 1663
rect 1766 1660 1767 1664
rect 1771 1660 1772 1664
rect 1766 1659 1772 1660
rect 1806 1660 1812 1661
rect 3462 1660 3468 1661
rect 1142 1658 1148 1659
rect 1806 1656 1807 1660
rect 1811 1656 1812 1660
rect 1806 1655 1812 1656
rect 2102 1659 2108 1660
rect 2102 1655 2103 1659
rect 2107 1655 2108 1659
rect 2102 1654 2108 1655
rect 2190 1659 2196 1660
rect 2190 1655 2191 1659
rect 2195 1655 2196 1659
rect 2190 1654 2196 1655
rect 2278 1659 2284 1660
rect 2278 1655 2279 1659
rect 2283 1655 2284 1659
rect 2278 1654 2284 1655
rect 2366 1659 2372 1660
rect 2366 1655 2367 1659
rect 2371 1655 2372 1659
rect 2366 1654 2372 1655
rect 2454 1659 2460 1660
rect 2454 1655 2455 1659
rect 2459 1655 2460 1659
rect 2454 1654 2460 1655
rect 2542 1659 2548 1660
rect 2542 1655 2543 1659
rect 2547 1655 2548 1659
rect 2542 1654 2548 1655
rect 2630 1659 2636 1660
rect 2630 1655 2631 1659
rect 2635 1655 2636 1659
rect 2630 1654 2636 1655
rect 2718 1659 2724 1660
rect 2718 1655 2719 1659
rect 2723 1655 2724 1659
rect 2718 1654 2724 1655
rect 2806 1659 2812 1660
rect 2806 1655 2807 1659
rect 2811 1655 2812 1659
rect 2806 1654 2812 1655
rect 2894 1659 2900 1660
rect 2894 1655 2895 1659
rect 2899 1655 2900 1659
rect 3462 1656 3463 1660
rect 3467 1656 3468 1660
rect 3462 1655 3468 1656
rect 2894 1654 2900 1655
rect 110 1647 116 1648
rect 110 1643 111 1647
rect 115 1643 116 1647
rect 1766 1647 1772 1648
rect 110 1642 116 1643
rect 398 1644 404 1645
rect 398 1640 399 1644
rect 403 1640 404 1644
rect 398 1639 404 1640
rect 486 1644 492 1645
rect 486 1640 487 1644
rect 491 1640 492 1644
rect 486 1639 492 1640
rect 574 1644 580 1645
rect 574 1640 575 1644
rect 579 1640 580 1644
rect 574 1639 580 1640
rect 662 1644 668 1645
rect 662 1640 663 1644
rect 667 1640 668 1644
rect 662 1639 668 1640
rect 758 1644 764 1645
rect 758 1640 759 1644
rect 763 1640 764 1644
rect 758 1639 764 1640
rect 854 1644 860 1645
rect 854 1640 855 1644
rect 859 1640 860 1644
rect 854 1639 860 1640
rect 950 1644 956 1645
rect 950 1640 951 1644
rect 955 1640 956 1644
rect 950 1639 956 1640
rect 1046 1644 1052 1645
rect 1046 1640 1047 1644
rect 1051 1640 1052 1644
rect 1046 1639 1052 1640
rect 1142 1644 1148 1645
rect 1142 1640 1143 1644
rect 1147 1640 1148 1644
rect 1766 1643 1767 1647
rect 1771 1643 1772 1647
rect 1766 1642 1772 1643
rect 1806 1643 1812 1644
rect 1142 1639 1148 1640
rect 1806 1639 1807 1643
rect 1811 1639 1812 1643
rect 3462 1643 3468 1644
rect 1806 1638 1812 1639
rect 2102 1640 2108 1641
rect 2102 1636 2103 1640
rect 2107 1636 2108 1640
rect 2102 1635 2108 1636
rect 2190 1640 2196 1641
rect 2190 1636 2191 1640
rect 2195 1636 2196 1640
rect 2190 1635 2196 1636
rect 2278 1640 2284 1641
rect 2278 1636 2279 1640
rect 2283 1636 2284 1640
rect 2278 1635 2284 1636
rect 2366 1640 2372 1641
rect 2366 1636 2367 1640
rect 2371 1636 2372 1640
rect 2366 1635 2372 1636
rect 2454 1640 2460 1641
rect 2454 1636 2455 1640
rect 2459 1636 2460 1640
rect 2454 1635 2460 1636
rect 2542 1640 2548 1641
rect 2542 1636 2543 1640
rect 2547 1636 2548 1640
rect 2542 1635 2548 1636
rect 2630 1640 2636 1641
rect 2630 1636 2631 1640
rect 2635 1636 2636 1640
rect 2630 1635 2636 1636
rect 2718 1640 2724 1641
rect 2718 1636 2719 1640
rect 2723 1636 2724 1640
rect 2718 1635 2724 1636
rect 2806 1640 2812 1641
rect 2806 1636 2807 1640
rect 2811 1636 2812 1640
rect 2806 1635 2812 1636
rect 2894 1640 2900 1641
rect 2894 1636 2895 1640
rect 2899 1636 2900 1640
rect 3462 1639 3463 1643
rect 3467 1639 3468 1643
rect 3462 1638 3468 1639
rect 2894 1635 2900 1636
rect 278 1596 284 1597
rect 110 1593 116 1594
rect 110 1589 111 1593
rect 115 1589 116 1593
rect 278 1592 279 1596
rect 283 1592 284 1596
rect 278 1591 284 1592
rect 382 1596 388 1597
rect 382 1592 383 1596
rect 387 1592 388 1596
rect 382 1591 388 1592
rect 494 1596 500 1597
rect 494 1592 495 1596
rect 499 1592 500 1596
rect 494 1591 500 1592
rect 606 1596 612 1597
rect 606 1592 607 1596
rect 611 1592 612 1596
rect 606 1591 612 1592
rect 718 1596 724 1597
rect 718 1592 719 1596
rect 723 1592 724 1596
rect 718 1591 724 1592
rect 830 1596 836 1597
rect 830 1592 831 1596
rect 835 1592 836 1596
rect 830 1591 836 1592
rect 942 1596 948 1597
rect 942 1592 943 1596
rect 947 1592 948 1596
rect 942 1591 948 1592
rect 1054 1596 1060 1597
rect 1054 1592 1055 1596
rect 1059 1592 1060 1596
rect 1054 1591 1060 1592
rect 1166 1596 1172 1597
rect 1166 1592 1167 1596
rect 1171 1592 1172 1596
rect 1166 1591 1172 1592
rect 1278 1596 1284 1597
rect 1278 1592 1279 1596
rect 1283 1592 1284 1596
rect 1278 1591 1284 1592
rect 1766 1593 1772 1594
rect 110 1588 116 1589
rect 1766 1589 1767 1593
rect 1771 1589 1772 1593
rect 2062 1592 2068 1593
rect 1766 1588 1772 1589
rect 1806 1589 1812 1590
rect 1806 1585 1807 1589
rect 1811 1585 1812 1589
rect 2062 1588 2063 1592
rect 2067 1588 2068 1592
rect 2062 1587 2068 1588
rect 2158 1592 2164 1593
rect 2158 1588 2159 1592
rect 2163 1588 2164 1592
rect 2158 1587 2164 1588
rect 2254 1592 2260 1593
rect 2254 1588 2255 1592
rect 2259 1588 2260 1592
rect 2254 1587 2260 1588
rect 2358 1592 2364 1593
rect 2358 1588 2359 1592
rect 2363 1588 2364 1592
rect 2358 1587 2364 1588
rect 2462 1592 2468 1593
rect 2462 1588 2463 1592
rect 2467 1588 2468 1592
rect 2462 1587 2468 1588
rect 2566 1592 2572 1593
rect 2566 1588 2567 1592
rect 2571 1588 2572 1592
rect 2566 1587 2572 1588
rect 2670 1592 2676 1593
rect 2670 1588 2671 1592
rect 2675 1588 2676 1592
rect 2670 1587 2676 1588
rect 2774 1592 2780 1593
rect 2774 1588 2775 1592
rect 2779 1588 2780 1592
rect 2774 1587 2780 1588
rect 2886 1592 2892 1593
rect 2886 1588 2887 1592
rect 2891 1588 2892 1592
rect 2886 1587 2892 1588
rect 3462 1589 3468 1590
rect 1806 1584 1812 1585
rect 3462 1585 3463 1589
rect 3467 1585 3468 1589
rect 3462 1584 3468 1585
rect 278 1577 284 1578
rect 110 1576 116 1577
rect 110 1572 111 1576
rect 115 1572 116 1576
rect 278 1573 279 1577
rect 283 1573 284 1577
rect 278 1572 284 1573
rect 382 1577 388 1578
rect 382 1573 383 1577
rect 387 1573 388 1577
rect 382 1572 388 1573
rect 494 1577 500 1578
rect 494 1573 495 1577
rect 499 1573 500 1577
rect 494 1572 500 1573
rect 606 1577 612 1578
rect 606 1573 607 1577
rect 611 1573 612 1577
rect 606 1572 612 1573
rect 718 1577 724 1578
rect 718 1573 719 1577
rect 723 1573 724 1577
rect 718 1572 724 1573
rect 830 1577 836 1578
rect 830 1573 831 1577
rect 835 1573 836 1577
rect 830 1572 836 1573
rect 942 1577 948 1578
rect 942 1573 943 1577
rect 947 1573 948 1577
rect 942 1572 948 1573
rect 1054 1577 1060 1578
rect 1054 1573 1055 1577
rect 1059 1573 1060 1577
rect 1054 1572 1060 1573
rect 1166 1577 1172 1578
rect 1166 1573 1167 1577
rect 1171 1573 1172 1577
rect 1166 1572 1172 1573
rect 1278 1577 1284 1578
rect 1278 1573 1279 1577
rect 1283 1573 1284 1577
rect 1278 1572 1284 1573
rect 1766 1576 1772 1577
rect 1766 1572 1767 1576
rect 1771 1572 1772 1576
rect 2062 1573 2068 1574
rect 110 1571 116 1572
rect 1766 1571 1772 1572
rect 1806 1572 1812 1573
rect 1806 1568 1807 1572
rect 1811 1568 1812 1572
rect 2062 1569 2063 1573
rect 2067 1569 2068 1573
rect 2062 1568 2068 1569
rect 2158 1573 2164 1574
rect 2158 1569 2159 1573
rect 2163 1569 2164 1573
rect 2158 1568 2164 1569
rect 2254 1573 2260 1574
rect 2254 1569 2255 1573
rect 2259 1569 2260 1573
rect 2254 1568 2260 1569
rect 2358 1573 2364 1574
rect 2358 1569 2359 1573
rect 2363 1569 2364 1573
rect 2358 1568 2364 1569
rect 2462 1573 2468 1574
rect 2462 1569 2463 1573
rect 2467 1569 2468 1573
rect 2462 1568 2468 1569
rect 2566 1573 2572 1574
rect 2566 1569 2567 1573
rect 2571 1569 2572 1573
rect 2566 1568 2572 1569
rect 2670 1573 2676 1574
rect 2670 1569 2671 1573
rect 2675 1569 2676 1573
rect 2670 1568 2676 1569
rect 2774 1573 2780 1574
rect 2774 1569 2775 1573
rect 2779 1569 2780 1573
rect 2774 1568 2780 1569
rect 2886 1573 2892 1574
rect 2886 1569 2887 1573
rect 2891 1569 2892 1573
rect 2886 1568 2892 1569
rect 3462 1572 3468 1573
rect 3462 1568 3463 1572
rect 3467 1568 3468 1572
rect 1806 1567 1812 1568
rect 3462 1567 3468 1568
rect 1806 1528 1812 1529
rect 3462 1528 3468 1529
rect 110 1524 116 1525
rect 1766 1524 1772 1525
rect 110 1520 111 1524
rect 115 1520 116 1524
rect 110 1519 116 1520
rect 182 1523 188 1524
rect 182 1519 183 1523
rect 187 1519 188 1523
rect 182 1518 188 1519
rect 326 1523 332 1524
rect 326 1519 327 1523
rect 331 1519 332 1523
rect 326 1518 332 1519
rect 470 1523 476 1524
rect 470 1519 471 1523
rect 475 1519 476 1523
rect 470 1518 476 1519
rect 622 1523 628 1524
rect 622 1519 623 1523
rect 627 1519 628 1523
rect 622 1518 628 1519
rect 766 1523 772 1524
rect 766 1519 767 1523
rect 771 1519 772 1523
rect 766 1518 772 1519
rect 910 1523 916 1524
rect 910 1519 911 1523
rect 915 1519 916 1523
rect 910 1518 916 1519
rect 1046 1523 1052 1524
rect 1046 1519 1047 1523
rect 1051 1519 1052 1523
rect 1046 1518 1052 1519
rect 1174 1523 1180 1524
rect 1174 1519 1175 1523
rect 1179 1519 1180 1523
rect 1174 1518 1180 1519
rect 1310 1523 1316 1524
rect 1310 1519 1311 1523
rect 1315 1519 1316 1523
rect 1310 1518 1316 1519
rect 1446 1523 1452 1524
rect 1446 1519 1447 1523
rect 1451 1519 1452 1523
rect 1766 1520 1767 1524
rect 1771 1520 1772 1524
rect 1806 1524 1807 1528
rect 1811 1524 1812 1528
rect 1806 1523 1812 1524
rect 1918 1527 1924 1528
rect 1918 1523 1919 1527
rect 1923 1523 1924 1527
rect 1918 1522 1924 1523
rect 2038 1527 2044 1528
rect 2038 1523 2039 1527
rect 2043 1523 2044 1527
rect 2038 1522 2044 1523
rect 2166 1527 2172 1528
rect 2166 1523 2167 1527
rect 2171 1523 2172 1527
rect 2166 1522 2172 1523
rect 2294 1527 2300 1528
rect 2294 1523 2295 1527
rect 2299 1523 2300 1527
rect 2294 1522 2300 1523
rect 2422 1527 2428 1528
rect 2422 1523 2423 1527
rect 2427 1523 2428 1527
rect 2422 1522 2428 1523
rect 2550 1527 2556 1528
rect 2550 1523 2551 1527
rect 2555 1523 2556 1527
rect 2550 1522 2556 1523
rect 2678 1527 2684 1528
rect 2678 1523 2679 1527
rect 2683 1523 2684 1527
rect 2678 1522 2684 1523
rect 2798 1527 2804 1528
rect 2798 1523 2799 1527
rect 2803 1523 2804 1527
rect 2798 1522 2804 1523
rect 2926 1527 2932 1528
rect 2926 1523 2927 1527
rect 2931 1523 2932 1527
rect 2926 1522 2932 1523
rect 3054 1527 3060 1528
rect 3054 1523 3055 1527
rect 3059 1523 3060 1527
rect 3462 1524 3463 1528
rect 3467 1524 3468 1528
rect 3462 1523 3468 1524
rect 3054 1522 3060 1523
rect 1766 1519 1772 1520
rect 1446 1518 1452 1519
rect 1806 1511 1812 1512
rect 110 1507 116 1508
rect 110 1503 111 1507
rect 115 1503 116 1507
rect 1766 1507 1772 1508
rect 110 1502 116 1503
rect 182 1504 188 1505
rect 182 1500 183 1504
rect 187 1500 188 1504
rect 182 1499 188 1500
rect 326 1504 332 1505
rect 326 1500 327 1504
rect 331 1500 332 1504
rect 326 1499 332 1500
rect 470 1504 476 1505
rect 470 1500 471 1504
rect 475 1500 476 1504
rect 470 1499 476 1500
rect 622 1504 628 1505
rect 622 1500 623 1504
rect 627 1500 628 1504
rect 622 1499 628 1500
rect 766 1504 772 1505
rect 766 1500 767 1504
rect 771 1500 772 1504
rect 766 1499 772 1500
rect 910 1504 916 1505
rect 910 1500 911 1504
rect 915 1500 916 1504
rect 910 1499 916 1500
rect 1046 1504 1052 1505
rect 1046 1500 1047 1504
rect 1051 1500 1052 1504
rect 1046 1499 1052 1500
rect 1174 1504 1180 1505
rect 1174 1500 1175 1504
rect 1179 1500 1180 1504
rect 1174 1499 1180 1500
rect 1310 1504 1316 1505
rect 1310 1500 1311 1504
rect 1315 1500 1316 1504
rect 1310 1499 1316 1500
rect 1446 1504 1452 1505
rect 1446 1500 1447 1504
rect 1451 1500 1452 1504
rect 1766 1503 1767 1507
rect 1771 1503 1772 1507
rect 1806 1507 1807 1511
rect 1811 1507 1812 1511
rect 3462 1511 3468 1512
rect 1806 1506 1812 1507
rect 1918 1508 1924 1509
rect 1918 1504 1919 1508
rect 1923 1504 1924 1508
rect 1918 1503 1924 1504
rect 2038 1508 2044 1509
rect 2038 1504 2039 1508
rect 2043 1504 2044 1508
rect 2038 1503 2044 1504
rect 2166 1508 2172 1509
rect 2166 1504 2167 1508
rect 2171 1504 2172 1508
rect 2166 1503 2172 1504
rect 2294 1508 2300 1509
rect 2294 1504 2295 1508
rect 2299 1504 2300 1508
rect 2294 1503 2300 1504
rect 2422 1508 2428 1509
rect 2422 1504 2423 1508
rect 2427 1504 2428 1508
rect 2422 1503 2428 1504
rect 2550 1508 2556 1509
rect 2550 1504 2551 1508
rect 2555 1504 2556 1508
rect 2550 1503 2556 1504
rect 2678 1508 2684 1509
rect 2678 1504 2679 1508
rect 2683 1504 2684 1508
rect 2678 1503 2684 1504
rect 2798 1508 2804 1509
rect 2798 1504 2799 1508
rect 2803 1504 2804 1508
rect 2798 1503 2804 1504
rect 2926 1508 2932 1509
rect 2926 1504 2927 1508
rect 2931 1504 2932 1508
rect 2926 1503 2932 1504
rect 3054 1508 3060 1509
rect 3054 1504 3055 1508
rect 3059 1504 3060 1508
rect 3462 1507 3463 1511
rect 3467 1507 3468 1511
rect 3462 1506 3468 1507
rect 3054 1503 3060 1504
rect 1766 1502 1772 1503
rect 1446 1499 1452 1500
rect 158 1456 164 1457
rect 110 1453 116 1454
rect 110 1449 111 1453
rect 115 1449 116 1453
rect 158 1452 159 1456
rect 163 1452 164 1456
rect 158 1451 164 1452
rect 374 1456 380 1457
rect 374 1452 375 1456
rect 379 1452 380 1456
rect 374 1451 380 1452
rect 582 1456 588 1457
rect 582 1452 583 1456
rect 587 1452 588 1456
rect 582 1451 588 1452
rect 782 1456 788 1457
rect 782 1452 783 1456
rect 787 1452 788 1456
rect 782 1451 788 1452
rect 958 1456 964 1457
rect 958 1452 959 1456
rect 963 1452 964 1456
rect 958 1451 964 1452
rect 1126 1456 1132 1457
rect 1126 1452 1127 1456
rect 1131 1452 1132 1456
rect 1126 1451 1132 1452
rect 1278 1456 1284 1457
rect 1278 1452 1279 1456
rect 1283 1452 1284 1456
rect 1278 1451 1284 1452
rect 1430 1456 1436 1457
rect 1430 1452 1431 1456
rect 1435 1452 1436 1456
rect 1430 1451 1436 1452
rect 1590 1456 1596 1457
rect 1590 1452 1591 1456
rect 1595 1452 1596 1456
rect 1830 1456 1836 1457
rect 1590 1451 1596 1452
rect 1766 1453 1772 1454
rect 110 1448 116 1449
rect 1766 1449 1767 1453
rect 1771 1449 1772 1453
rect 1766 1448 1772 1449
rect 1806 1453 1812 1454
rect 1806 1449 1807 1453
rect 1811 1449 1812 1453
rect 1830 1452 1831 1456
rect 1835 1452 1836 1456
rect 1830 1451 1836 1452
rect 1950 1456 1956 1457
rect 1950 1452 1951 1456
rect 1955 1452 1956 1456
rect 1950 1451 1956 1452
rect 2110 1456 2116 1457
rect 2110 1452 2111 1456
rect 2115 1452 2116 1456
rect 2110 1451 2116 1452
rect 2270 1456 2276 1457
rect 2270 1452 2271 1456
rect 2275 1452 2276 1456
rect 2270 1451 2276 1452
rect 2430 1456 2436 1457
rect 2430 1452 2431 1456
rect 2435 1452 2436 1456
rect 2430 1451 2436 1452
rect 2590 1456 2596 1457
rect 2590 1452 2591 1456
rect 2595 1452 2596 1456
rect 2590 1451 2596 1452
rect 2734 1456 2740 1457
rect 2734 1452 2735 1456
rect 2739 1452 2740 1456
rect 2734 1451 2740 1452
rect 2870 1456 2876 1457
rect 2870 1452 2871 1456
rect 2875 1452 2876 1456
rect 2870 1451 2876 1452
rect 3006 1456 3012 1457
rect 3006 1452 3007 1456
rect 3011 1452 3012 1456
rect 3006 1451 3012 1452
rect 3134 1456 3140 1457
rect 3134 1452 3135 1456
rect 3139 1452 3140 1456
rect 3134 1451 3140 1452
rect 3262 1456 3268 1457
rect 3262 1452 3263 1456
rect 3267 1452 3268 1456
rect 3262 1451 3268 1452
rect 3366 1456 3372 1457
rect 3366 1452 3367 1456
rect 3371 1452 3372 1456
rect 3366 1451 3372 1452
rect 3462 1453 3468 1454
rect 1806 1448 1812 1449
rect 3462 1449 3463 1453
rect 3467 1449 3468 1453
rect 3462 1448 3468 1449
rect 158 1437 164 1438
rect 110 1436 116 1437
rect 110 1432 111 1436
rect 115 1432 116 1436
rect 158 1433 159 1437
rect 163 1433 164 1437
rect 158 1432 164 1433
rect 374 1437 380 1438
rect 374 1433 375 1437
rect 379 1433 380 1437
rect 374 1432 380 1433
rect 582 1437 588 1438
rect 582 1433 583 1437
rect 587 1433 588 1437
rect 582 1432 588 1433
rect 782 1437 788 1438
rect 782 1433 783 1437
rect 787 1433 788 1437
rect 782 1432 788 1433
rect 958 1437 964 1438
rect 958 1433 959 1437
rect 963 1433 964 1437
rect 958 1432 964 1433
rect 1126 1437 1132 1438
rect 1126 1433 1127 1437
rect 1131 1433 1132 1437
rect 1126 1432 1132 1433
rect 1278 1437 1284 1438
rect 1278 1433 1279 1437
rect 1283 1433 1284 1437
rect 1278 1432 1284 1433
rect 1430 1437 1436 1438
rect 1430 1433 1431 1437
rect 1435 1433 1436 1437
rect 1430 1432 1436 1433
rect 1590 1437 1596 1438
rect 1830 1437 1836 1438
rect 1590 1433 1591 1437
rect 1595 1433 1596 1437
rect 1590 1432 1596 1433
rect 1766 1436 1772 1437
rect 1766 1432 1767 1436
rect 1771 1432 1772 1436
rect 110 1431 116 1432
rect 1766 1431 1772 1432
rect 1806 1436 1812 1437
rect 1806 1432 1807 1436
rect 1811 1432 1812 1436
rect 1830 1433 1831 1437
rect 1835 1433 1836 1437
rect 1830 1432 1836 1433
rect 1950 1437 1956 1438
rect 1950 1433 1951 1437
rect 1955 1433 1956 1437
rect 1950 1432 1956 1433
rect 2110 1437 2116 1438
rect 2110 1433 2111 1437
rect 2115 1433 2116 1437
rect 2110 1432 2116 1433
rect 2270 1437 2276 1438
rect 2270 1433 2271 1437
rect 2275 1433 2276 1437
rect 2270 1432 2276 1433
rect 2430 1437 2436 1438
rect 2430 1433 2431 1437
rect 2435 1433 2436 1437
rect 2430 1432 2436 1433
rect 2590 1437 2596 1438
rect 2590 1433 2591 1437
rect 2595 1433 2596 1437
rect 2590 1432 2596 1433
rect 2734 1437 2740 1438
rect 2734 1433 2735 1437
rect 2739 1433 2740 1437
rect 2734 1432 2740 1433
rect 2870 1437 2876 1438
rect 2870 1433 2871 1437
rect 2875 1433 2876 1437
rect 2870 1432 2876 1433
rect 3006 1437 3012 1438
rect 3006 1433 3007 1437
rect 3011 1433 3012 1437
rect 3006 1432 3012 1433
rect 3134 1437 3140 1438
rect 3134 1433 3135 1437
rect 3139 1433 3140 1437
rect 3134 1432 3140 1433
rect 3262 1437 3268 1438
rect 3262 1433 3263 1437
rect 3267 1433 3268 1437
rect 3262 1432 3268 1433
rect 3366 1437 3372 1438
rect 3366 1433 3367 1437
rect 3371 1433 3372 1437
rect 3366 1432 3372 1433
rect 3462 1436 3468 1437
rect 3462 1432 3463 1436
rect 3467 1432 3468 1436
rect 1806 1431 1812 1432
rect 3462 1431 3468 1432
rect 110 1388 116 1389
rect 1766 1388 1772 1389
rect 110 1384 111 1388
rect 115 1384 116 1388
rect 110 1383 116 1384
rect 134 1387 140 1388
rect 134 1383 135 1387
rect 139 1383 140 1387
rect 134 1382 140 1383
rect 302 1387 308 1388
rect 302 1383 303 1387
rect 307 1383 308 1387
rect 302 1382 308 1383
rect 494 1387 500 1388
rect 494 1383 495 1387
rect 499 1383 500 1387
rect 494 1382 500 1383
rect 678 1387 684 1388
rect 678 1383 679 1387
rect 683 1383 684 1387
rect 678 1382 684 1383
rect 854 1387 860 1388
rect 854 1383 855 1387
rect 859 1383 860 1387
rect 854 1382 860 1383
rect 1014 1387 1020 1388
rect 1014 1383 1015 1387
rect 1019 1383 1020 1387
rect 1014 1382 1020 1383
rect 1166 1387 1172 1388
rect 1166 1383 1167 1387
rect 1171 1383 1172 1387
rect 1166 1382 1172 1383
rect 1302 1387 1308 1388
rect 1302 1383 1303 1387
rect 1307 1383 1308 1387
rect 1302 1382 1308 1383
rect 1430 1387 1436 1388
rect 1430 1383 1431 1387
rect 1435 1383 1436 1387
rect 1430 1382 1436 1383
rect 1558 1387 1564 1388
rect 1558 1383 1559 1387
rect 1563 1383 1564 1387
rect 1558 1382 1564 1383
rect 1670 1387 1676 1388
rect 1670 1383 1671 1387
rect 1675 1383 1676 1387
rect 1766 1384 1767 1388
rect 1771 1384 1772 1388
rect 1766 1383 1772 1384
rect 1806 1388 1812 1389
rect 3462 1388 3468 1389
rect 1806 1384 1807 1388
rect 1811 1384 1812 1388
rect 1806 1383 1812 1384
rect 1830 1387 1836 1388
rect 1830 1383 1831 1387
rect 1835 1383 1836 1387
rect 1670 1382 1676 1383
rect 1830 1382 1836 1383
rect 2006 1387 2012 1388
rect 2006 1383 2007 1387
rect 2011 1383 2012 1387
rect 2006 1382 2012 1383
rect 2198 1387 2204 1388
rect 2198 1383 2199 1387
rect 2203 1383 2204 1387
rect 2198 1382 2204 1383
rect 2382 1387 2388 1388
rect 2382 1383 2383 1387
rect 2387 1383 2388 1387
rect 2382 1382 2388 1383
rect 2558 1387 2564 1388
rect 2558 1383 2559 1387
rect 2563 1383 2564 1387
rect 2558 1382 2564 1383
rect 2718 1387 2724 1388
rect 2718 1383 2719 1387
rect 2723 1383 2724 1387
rect 2718 1382 2724 1383
rect 2862 1387 2868 1388
rect 2862 1383 2863 1387
rect 2867 1383 2868 1387
rect 2862 1382 2868 1383
rect 2998 1387 3004 1388
rect 2998 1383 2999 1387
rect 3003 1383 3004 1387
rect 2998 1382 3004 1383
rect 3126 1387 3132 1388
rect 3126 1383 3127 1387
rect 3131 1383 3132 1387
rect 3126 1382 3132 1383
rect 3254 1387 3260 1388
rect 3254 1383 3255 1387
rect 3259 1383 3260 1387
rect 3254 1382 3260 1383
rect 3366 1387 3372 1388
rect 3366 1383 3367 1387
rect 3371 1383 3372 1387
rect 3462 1384 3463 1388
rect 3467 1384 3468 1388
rect 3462 1383 3468 1384
rect 3366 1382 3372 1383
rect 110 1371 116 1372
rect 110 1367 111 1371
rect 115 1367 116 1371
rect 1766 1371 1772 1372
rect 110 1366 116 1367
rect 134 1368 140 1369
rect 134 1364 135 1368
rect 139 1364 140 1368
rect 134 1363 140 1364
rect 302 1368 308 1369
rect 302 1364 303 1368
rect 307 1364 308 1368
rect 302 1363 308 1364
rect 494 1368 500 1369
rect 494 1364 495 1368
rect 499 1364 500 1368
rect 494 1363 500 1364
rect 678 1368 684 1369
rect 678 1364 679 1368
rect 683 1364 684 1368
rect 678 1363 684 1364
rect 854 1368 860 1369
rect 854 1364 855 1368
rect 859 1364 860 1368
rect 854 1363 860 1364
rect 1014 1368 1020 1369
rect 1014 1364 1015 1368
rect 1019 1364 1020 1368
rect 1014 1363 1020 1364
rect 1166 1368 1172 1369
rect 1166 1364 1167 1368
rect 1171 1364 1172 1368
rect 1166 1363 1172 1364
rect 1302 1368 1308 1369
rect 1302 1364 1303 1368
rect 1307 1364 1308 1368
rect 1302 1363 1308 1364
rect 1430 1368 1436 1369
rect 1430 1364 1431 1368
rect 1435 1364 1436 1368
rect 1430 1363 1436 1364
rect 1558 1368 1564 1369
rect 1558 1364 1559 1368
rect 1563 1364 1564 1368
rect 1558 1363 1564 1364
rect 1670 1368 1676 1369
rect 1670 1364 1671 1368
rect 1675 1364 1676 1368
rect 1766 1367 1767 1371
rect 1771 1367 1772 1371
rect 1766 1366 1772 1367
rect 1806 1371 1812 1372
rect 1806 1367 1807 1371
rect 1811 1367 1812 1371
rect 3462 1371 3468 1372
rect 1806 1366 1812 1367
rect 1830 1368 1836 1369
rect 1670 1363 1676 1364
rect 1830 1364 1831 1368
rect 1835 1364 1836 1368
rect 1830 1363 1836 1364
rect 2006 1368 2012 1369
rect 2006 1364 2007 1368
rect 2011 1364 2012 1368
rect 2006 1363 2012 1364
rect 2198 1368 2204 1369
rect 2198 1364 2199 1368
rect 2203 1364 2204 1368
rect 2198 1363 2204 1364
rect 2382 1368 2388 1369
rect 2382 1364 2383 1368
rect 2387 1364 2388 1368
rect 2382 1363 2388 1364
rect 2558 1368 2564 1369
rect 2558 1364 2559 1368
rect 2563 1364 2564 1368
rect 2558 1363 2564 1364
rect 2718 1368 2724 1369
rect 2718 1364 2719 1368
rect 2723 1364 2724 1368
rect 2718 1363 2724 1364
rect 2862 1368 2868 1369
rect 2862 1364 2863 1368
rect 2867 1364 2868 1368
rect 2862 1363 2868 1364
rect 2998 1368 3004 1369
rect 2998 1364 2999 1368
rect 3003 1364 3004 1368
rect 2998 1363 3004 1364
rect 3126 1368 3132 1369
rect 3126 1364 3127 1368
rect 3131 1364 3132 1368
rect 3126 1363 3132 1364
rect 3254 1368 3260 1369
rect 3254 1364 3255 1368
rect 3259 1364 3260 1368
rect 3254 1363 3260 1364
rect 3366 1368 3372 1369
rect 3366 1364 3367 1368
rect 3371 1364 3372 1368
rect 3462 1367 3463 1371
rect 3467 1367 3468 1371
rect 3462 1366 3468 1367
rect 3366 1363 3372 1364
rect 134 1320 140 1321
rect 110 1317 116 1318
rect 110 1313 111 1317
rect 115 1313 116 1317
rect 134 1316 135 1320
rect 139 1316 140 1320
rect 134 1315 140 1316
rect 246 1320 252 1321
rect 246 1316 247 1320
rect 251 1316 252 1320
rect 246 1315 252 1316
rect 398 1320 404 1321
rect 398 1316 399 1320
rect 403 1316 404 1320
rect 398 1315 404 1316
rect 558 1320 564 1321
rect 558 1316 559 1320
rect 563 1316 564 1320
rect 558 1315 564 1316
rect 726 1320 732 1321
rect 726 1316 727 1320
rect 731 1316 732 1320
rect 726 1315 732 1316
rect 894 1320 900 1321
rect 894 1316 895 1320
rect 899 1316 900 1320
rect 894 1315 900 1316
rect 1062 1320 1068 1321
rect 1062 1316 1063 1320
rect 1067 1316 1068 1320
rect 1062 1315 1068 1316
rect 1222 1320 1228 1321
rect 1222 1316 1223 1320
rect 1227 1316 1228 1320
rect 1222 1315 1228 1316
rect 1374 1320 1380 1321
rect 1374 1316 1375 1320
rect 1379 1316 1380 1320
rect 1374 1315 1380 1316
rect 1534 1320 1540 1321
rect 1534 1316 1535 1320
rect 1539 1316 1540 1320
rect 1534 1315 1540 1316
rect 1670 1320 1676 1321
rect 1670 1316 1671 1320
rect 1675 1316 1676 1320
rect 1670 1315 1676 1316
rect 1766 1317 1772 1318
rect 110 1312 116 1313
rect 1766 1313 1767 1317
rect 1771 1313 1772 1317
rect 1830 1316 1836 1317
rect 1766 1312 1772 1313
rect 1806 1313 1812 1314
rect 1806 1309 1807 1313
rect 1811 1309 1812 1313
rect 1830 1312 1831 1316
rect 1835 1312 1836 1316
rect 1830 1311 1836 1312
rect 1966 1316 1972 1317
rect 1966 1312 1967 1316
rect 1971 1312 1972 1316
rect 1966 1311 1972 1312
rect 2142 1316 2148 1317
rect 2142 1312 2143 1316
rect 2147 1312 2148 1316
rect 2142 1311 2148 1312
rect 2326 1316 2332 1317
rect 2326 1312 2327 1316
rect 2331 1312 2332 1316
rect 2326 1311 2332 1312
rect 2510 1316 2516 1317
rect 2510 1312 2511 1316
rect 2515 1312 2516 1316
rect 2510 1311 2516 1312
rect 2686 1316 2692 1317
rect 2686 1312 2687 1316
rect 2691 1312 2692 1316
rect 2686 1311 2692 1312
rect 2862 1316 2868 1317
rect 2862 1312 2863 1316
rect 2867 1312 2868 1316
rect 2862 1311 2868 1312
rect 3038 1316 3044 1317
rect 3038 1312 3039 1316
rect 3043 1312 3044 1316
rect 3038 1311 3044 1312
rect 3214 1316 3220 1317
rect 3214 1312 3215 1316
rect 3219 1312 3220 1316
rect 3214 1311 3220 1312
rect 3366 1316 3372 1317
rect 3366 1312 3367 1316
rect 3371 1312 3372 1316
rect 3366 1311 3372 1312
rect 3462 1313 3468 1314
rect 1806 1308 1812 1309
rect 3462 1309 3463 1313
rect 3467 1309 3468 1313
rect 3462 1308 3468 1309
rect 134 1301 140 1302
rect 110 1300 116 1301
rect 110 1296 111 1300
rect 115 1296 116 1300
rect 134 1297 135 1301
rect 139 1297 140 1301
rect 134 1296 140 1297
rect 246 1301 252 1302
rect 246 1297 247 1301
rect 251 1297 252 1301
rect 246 1296 252 1297
rect 398 1301 404 1302
rect 398 1297 399 1301
rect 403 1297 404 1301
rect 398 1296 404 1297
rect 558 1301 564 1302
rect 558 1297 559 1301
rect 563 1297 564 1301
rect 558 1296 564 1297
rect 726 1301 732 1302
rect 726 1297 727 1301
rect 731 1297 732 1301
rect 726 1296 732 1297
rect 894 1301 900 1302
rect 894 1297 895 1301
rect 899 1297 900 1301
rect 894 1296 900 1297
rect 1062 1301 1068 1302
rect 1062 1297 1063 1301
rect 1067 1297 1068 1301
rect 1062 1296 1068 1297
rect 1222 1301 1228 1302
rect 1222 1297 1223 1301
rect 1227 1297 1228 1301
rect 1222 1296 1228 1297
rect 1374 1301 1380 1302
rect 1374 1297 1375 1301
rect 1379 1297 1380 1301
rect 1374 1296 1380 1297
rect 1534 1301 1540 1302
rect 1534 1297 1535 1301
rect 1539 1297 1540 1301
rect 1534 1296 1540 1297
rect 1670 1301 1676 1302
rect 1670 1297 1671 1301
rect 1675 1297 1676 1301
rect 1670 1296 1676 1297
rect 1766 1300 1772 1301
rect 1766 1296 1767 1300
rect 1771 1296 1772 1300
rect 1830 1297 1836 1298
rect 110 1295 116 1296
rect 1766 1295 1772 1296
rect 1806 1296 1812 1297
rect 1806 1292 1807 1296
rect 1811 1292 1812 1296
rect 1830 1293 1831 1297
rect 1835 1293 1836 1297
rect 1830 1292 1836 1293
rect 1966 1297 1972 1298
rect 1966 1293 1967 1297
rect 1971 1293 1972 1297
rect 1966 1292 1972 1293
rect 2142 1297 2148 1298
rect 2142 1293 2143 1297
rect 2147 1293 2148 1297
rect 2142 1292 2148 1293
rect 2326 1297 2332 1298
rect 2326 1293 2327 1297
rect 2331 1293 2332 1297
rect 2326 1292 2332 1293
rect 2510 1297 2516 1298
rect 2510 1293 2511 1297
rect 2515 1293 2516 1297
rect 2510 1292 2516 1293
rect 2686 1297 2692 1298
rect 2686 1293 2687 1297
rect 2691 1293 2692 1297
rect 2686 1292 2692 1293
rect 2862 1297 2868 1298
rect 2862 1293 2863 1297
rect 2867 1293 2868 1297
rect 2862 1292 2868 1293
rect 3038 1297 3044 1298
rect 3038 1293 3039 1297
rect 3043 1293 3044 1297
rect 3038 1292 3044 1293
rect 3214 1297 3220 1298
rect 3214 1293 3215 1297
rect 3219 1293 3220 1297
rect 3214 1292 3220 1293
rect 3366 1297 3372 1298
rect 3366 1293 3367 1297
rect 3371 1293 3372 1297
rect 3366 1292 3372 1293
rect 3462 1296 3468 1297
rect 3462 1292 3463 1296
rect 3467 1292 3468 1296
rect 1806 1291 1812 1292
rect 3462 1291 3468 1292
rect 110 1252 116 1253
rect 1766 1252 1772 1253
rect 110 1248 111 1252
rect 115 1248 116 1252
rect 110 1247 116 1248
rect 134 1251 140 1252
rect 134 1247 135 1251
rect 139 1247 140 1251
rect 134 1246 140 1247
rect 222 1251 228 1252
rect 222 1247 223 1251
rect 227 1247 228 1251
rect 222 1246 228 1247
rect 318 1251 324 1252
rect 318 1247 319 1251
rect 323 1247 324 1251
rect 318 1246 324 1247
rect 430 1251 436 1252
rect 430 1247 431 1251
rect 435 1247 436 1251
rect 430 1246 436 1247
rect 550 1251 556 1252
rect 550 1247 551 1251
rect 555 1247 556 1251
rect 550 1246 556 1247
rect 678 1251 684 1252
rect 678 1247 679 1251
rect 683 1247 684 1251
rect 678 1246 684 1247
rect 822 1251 828 1252
rect 822 1247 823 1251
rect 827 1247 828 1251
rect 822 1246 828 1247
rect 974 1251 980 1252
rect 974 1247 975 1251
rect 979 1247 980 1251
rect 974 1246 980 1247
rect 1142 1251 1148 1252
rect 1142 1247 1143 1251
rect 1147 1247 1148 1251
rect 1142 1246 1148 1247
rect 1318 1251 1324 1252
rect 1318 1247 1319 1251
rect 1323 1247 1324 1251
rect 1318 1246 1324 1247
rect 1502 1251 1508 1252
rect 1502 1247 1503 1251
rect 1507 1247 1508 1251
rect 1502 1246 1508 1247
rect 1670 1251 1676 1252
rect 1670 1247 1671 1251
rect 1675 1247 1676 1251
rect 1766 1248 1767 1252
rect 1771 1248 1772 1252
rect 1766 1247 1772 1248
rect 1806 1252 1812 1253
rect 3462 1252 3468 1253
rect 1806 1248 1807 1252
rect 1811 1248 1812 1252
rect 1806 1247 1812 1248
rect 1830 1251 1836 1252
rect 1830 1247 1831 1251
rect 1835 1247 1836 1251
rect 1670 1246 1676 1247
rect 1830 1246 1836 1247
rect 2094 1251 2100 1252
rect 2094 1247 2095 1251
rect 2099 1247 2100 1251
rect 2094 1246 2100 1247
rect 2358 1251 2364 1252
rect 2358 1247 2359 1251
rect 2363 1247 2364 1251
rect 2358 1246 2364 1247
rect 2598 1251 2604 1252
rect 2598 1247 2599 1251
rect 2603 1247 2604 1251
rect 2598 1246 2604 1247
rect 2806 1251 2812 1252
rect 2806 1247 2807 1251
rect 2811 1247 2812 1251
rect 2806 1246 2812 1247
rect 3006 1251 3012 1252
rect 3006 1247 3007 1251
rect 3011 1247 3012 1251
rect 3006 1246 3012 1247
rect 3198 1251 3204 1252
rect 3198 1247 3199 1251
rect 3203 1247 3204 1251
rect 3198 1246 3204 1247
rect 3366 1251 3372 1252
rect 3366 1247 3367 1251
rect 3371 1247 3372 1251
rect 3462 1248 3463 1252
rect 3467 1248 3468 1252
rect 3462 1247 3468 1248
rect 3366 1246 3372 1247
rect 110 1235 116 1236
rect 110 1231 111 1235
rect 115 1231 116 1235
rect 1766 1235 1772 1236
rect 110 1230 116 1231
rect 134 1232 140 1233
rect 134 1228 135 1232
rect 139 1228 140 1232
rect 134 1227 140 1228
rect 222 1232 228 1233
rect 222 1228 223 1232
rect 227 1228 228 1232
rect 222 1227 228 1228
rect 318 1232 324 1233
rect 318 1228 319 1232
rect 323 1228 324 1232
rect 318 1227 324 1228
rect 430 1232 436 1233
rect 430 1228 431 1232
rect 435 1228 436 1232
rect 430 1227 436 1228
rect 550 1232 556 1233
rect 550 1228 551 1232
rect 555 1228 556 1232
rect 550 1227 556 1228
rect 678 1232 684 1233
rect 678 1228 679 1232
rect 683 1228 684 1232
rect 678 1227 684 1228
rect 822 1232 828 1233
rect 822 1228 823 1232
rect 827 1228 828 1232
rect 822 1227 828 1228
rect 974 1232 980 1233
rect 974 1228 975 1232
rect 979 1228 980 1232
rect 974 1227 980 1228
rect 1142 1232 1148 1233
rect 1142 1228 1143 1232
rect 1147 1228 1148 1232
rect 1142 1227 1148 1228
rect 1318 1232 1324 1233
rect 1318 1228 1319 1232
rect 1323 1228 1324 1232
rect 1318 1227 1324 1228
rect 1502 1232 1508 1233
rect 1502 1228 1503 1232
rect 1507 1228 1508 1232
rect 1502 1227 1508 1228
rect 1670 1232 1676 1233
rect 1670 1228 1671 1232
rect 1675 1228 1676 1232
rect 1766 1231 1767 1235
rect 1771 1231 1772 1235
rect 1766 1230 1772 1231
rect 1806 1235 1812 1236
rect 1806 1231 1807 1235
rect 1811 1231 1812 1235
rect 3462 1235 3468 1236
rect 1806 1230 1812 1231
rect 1830 1232 1836 1233
rect 1670 1227 1676 1228
rect 1830 1228 1831 1232
rect 1835 1228 1836 1232
rect 1830 1227 1836 1228
rect 2094 1232 2100 1233
rect 2094 1228 2095 1232
rect 2099 1228 2100 1232
rect 2094 1227 2100 1228
rect 2358 1232 2364 1233
rect 2358 1228 2359 1232
rect 2363 1228 2364 1232
rect 2358 1227 2364 1228
rect 2598 1232 2604 1233
rect 2598 1228 2599 1232
rect 2603 1228 2604 1232
rect 2598 1227 2604 1228
rect 2806 1232 2812 1233
rect 2806 1228 2807 1232
rect 2811 1228 2812 1232
rect 2806 1227 2812 1228
rect 3006 1232 3012 1233
rect 3006 1228 3007 1232
rect 3011 1228 3012 1232
rect 3006 1227 3012 1228
rect 3198 1232 3204 1233
rect 3198 1228 3199 1232
rect 3203 1228 3204 1232
rect 3198 1227 3204 1228
rect 3366 1232 3372 1233
rect 3366 1228 3367 1232
rect 3371 1228 3372 1232
rect 3462 1231 3463 1235
rect 3467 1231 3468 1235
rect 3462 1230 3468 1231
rect 3366 1227 3372 1228
rect 134 1180 140 1181
rect 110 1177 116 1178
rect 110 1173 111 1177
rect 115 1173 116 1177
rect 134 1176 135 1180
rect 139 1176 140 1180
rect 134 1175 140 1176
rect 230 1180 236 1181
rect 230 1176 231 1180
rect 235 1176 236 1180
rect 230 1175 236 1176
rect 358 1180 364 1181
rect 358 1176 359 1180
rect 363 1176 364 1180
rect 358 1175 364 1176
rect 486 1180 492 1181
rect 486 1176 487 1180
rect 491 1176 492 1180
rect 486 1175 492 1176
rect 614 1180 620 1181
rect 614 1176 615 1180
rect 619 1176 620 1180
rect 614 1175 620 1176
rect 742 1180 748 1181
rect 742 1176 743 1180
rect 747 1176 748 1180
rect 742 1175 748 1176
rect 870 1180 876 1181
rect 870 1176 871 1180
rect 875 1176 876 1180
rect 870 1175 876 1176
rect 990 1180 996 1181
rect 990 1176 991 1180
rect 995 1176 996 1180
rect 990 1175 996 1176
rect 1118 1180 1124 1181
rect 1118 1176 1119 1180
rect 1123 1176 1124 1180
rect 1118 1175 1124 1176
rect 1246 1180 1252 1181
rect 1246 1176 1247 1180
rect 1251 1176 1252 1180
rect 1934 1180 1940 1181
rect 1246 1175 1252 1176
rect 1766 1177 1772 1178
rect 110 1172 116 1173
rect 1766 1173 1767 1177
rect 1771 1173 1772 1177
rect 1766 1172 1772 1173
rect 1806 1177 1812 1178
rect 1806 1173 1807 1177
rect 1811 1173 1812 1177
rect 1934 1176 1935 1180
rect 1939 1176 1940 1180
rect 1934 1175 1940 1176
rect 2038 1180 2044 1181
rect 2038 1176 2039 1180
rect 2043 1176 2044 1180
rect 2038 1175 2044 1176
rect 2158 1180 2164 1181
rect 2158 1176 2159 1180
rect 2163 1176 2164 1180
rect 2158 1175 2164 1176
rect 2286 1180 2292 1181
rect 2286 1176 2287 1180
rect 2291 1176 2292 1180
rect 2286 1175 2292 1176
rect 2422 1180 2428 1181
rect 2422 1176 2423 1180
rect 2427 1176 2428 1180
rect 2422 1175 2428 1176
rect 2566 1180 2572 1181
rect 2566 1176 2567 1180
rect 2571 1176 2572 1180
rect 2566 1175 2572 1176
rect 2702 1180 2708 1181
rect 2702 1176 2703 1180
rect 2707 1176 2708 1180
rect 2702 1175 2708 1176
rect 2838 1180 2844 1181
rect 2838 1176 2839 1180
rect 2843 1176 2844 1180
rect 2838 1175 2844 1176
rect 2974 1180 2980 1181
rect 2974 1176 2975 1180
rect 2979 1176 2980 1180
rect 2974 1175 2980 1176
rect 3110 1180 3116 1181
rect 3110 1176 3111 1180
rect 3115 1176 3116 1180
rect 3110 1175 3116 1176
rect 3246 1180 3252 1181
rect 3246 1176 3247 1180
rect 3251 1176 3252 1180
rect 3246 1175 3252 1176
rect 3366 1180 3372 1181
rect 3366 1176 3367 1180
rect 3371 1176 3372 1180
rect 3366 1175 3372 1176
rect 3462 1177 3468 1178
rect 1806 1172 1812 1173
rect 3462 1173 3463 1177
rect 3467 1173 3468 1177
rect 3462 1172 3468 1173
rect 134 1161 140 1162
rect 110 1160 116 1161
rect 110 1156 111 1160
rect 115 1156 116 1160
rect 134 1157 135 1161
rect 139 1157 140 1161
rect 134 1156 140 1157
rect 230 1161 236 1162
rect 230 1157 231 1161
rect 235 1157 236 1161
rect 230 1156 236 1157
rect 358 1161 364 1162
rect 358 1157 359 1161
rect 363 1157 364 1161
rect 358 1156 364 1157
rect 486 1161 492 1162
rect 486 1157 487 1161
rect 491 1157 492 1161
rect 486 1156 492 1157
rect 614 1161 620 1162
rect 614 1157 615 1161
rect 619 1157 620 1161
rect 614 1156 620 1157
rect 742 1161 748 1162
rect 742 1157 743 1161
rect 747 1157 748 1161
rect 742 1156 748 1157
rect 870 1161 876 1162
rect 870 1157 871 1161
rect 875 1157 876 1161
rect 870 1156 876 1157
rect 990 1161 996 1162
rect 990 1157 991 1161
rect 995 1157 996 1161
rect 990 1156 996 1157
rect 1118 1161 1124 1162
rect 1118 1157 1119 1161
rect 1123 1157 1124 1161
rect 1118 1156 1124 1157
rect 1246 1161 1252 1162
rect 1934 1161 1940 1162
rect 1246 1157 1247 1161
rect 1251 1157 1252 1161
rect 1246 1156 1252 1157
rect 1766 1160 1772 1161
rect 1766 1156 1767 1160
rect 1771 1156 1772 1160
rect 110 1155 116 1156
rect 1766 1155 1772 1156
rect 1806 1160 1812 1161
rect 1806 1156 1807 1160
rect 1811 1156 1812 1160
rect 1934 1157 1935 1161
rect 1939 1157 1940 1161
rect 1934 1156 1940 1157
rect 2038 1161 2044 1162
rect 2038 1157 2039 1161
rect 2043 1157 2044 1161
rect 2038 1156 2044 1157
rect 2158 1161 2164 1162
rect 2158 1157 2159 1161
rect 2163 1157 2164 1161
rect 2158 1156 2164 1157
rect 2286 1161 2292 1162
rect 2286 1157 2287 1161
rect 2291 1157 2292 1161
rect 2286 1156 2292 1157
rect 2422 1161 2428 1162
rect 2422 1157 2423 1161
rect 2427 1157 2428 1161
rect 2422 1156 2428 1157
rect 2566 1161 2572 1162
rect 2566 1157 2567 1161
rect 2571 1157 2572 1161
rect 2566 1156 2572 1157
rect 2702 1161 2708 1162
rect 2702 1157 2703 1161
rect 2707 1157 2708 1161
rect 2702 1156 2708 1157
rect 2838 1161 2844 1162
rect 2838 1157 2839 1161
rect 2843 1157 2844 1161
rect 2838 1156 2844 1157
rect 2974 1161 2980 1162
rect 2974 1157 2975 1161
rect 2979 1157 2980 1161
rect 2974 1156 2980 1157
rect 3110 1161 3116 1162
rect 3110 1157 3111 1161
rect 3115 1157 3116 1161
rect 3110 1156 3116 1157
rect 3246 1161 3252 1162
rect 3246 1157 3247 1161
rect 3251 1157 3252 1161
rect 3246 1156 3252 1157
rect 3366 1161 3372 1162
rect 3366 1157 3367 1161
rect 3371 1157 3372 1161
rect 3366 1156 3372 1157
rect 3462 1160 3468 1161
rect 3462 1156 3463 1160
rect 3467 1156 3468 1160
rect 1806 1155 1812 1156
rect 3462 1155 3468 1156
rect 110 1112 116 1113
rect 1766 1112 1772 1113
rect 110 1108 111 1112
rect 115 1108 116 1112
rect 110 1107 116 1108
rect 246 1111 252 1112
rect 246 1107 247 1111
rect 251 1107 252 1111
rect 246 1106 252 1107
rect 366 1111 372 1112
rect 366 1107 367 1111
rect 371 1107 372 1111
rect 366 1106 372 1107
rect 494 1111 500 1112
rect 494 1107 495 1111
rect 499 1107 500 1111
rect 494 1106 500 1107
rect 622 1111 628 1112
rect 622 1107 623 1111
rect 627 1107 628 1111
rect 622 1106 628 1107
rect 758 1111 764 1112
rect 758 1107 759 1111
rect 763 1107 764 1111
rect 758 1106 764 1107
rect 886 1111 892 1112
rect 886 1107 887 1111
rect 891 1107 892 1111
rect 886 1106 892 1107
rect 1014 1111 1020 1112
rect 1014 1107 1015 1111
rect 1019 1107 1020 1111
rect 1014 1106 1020 1107
rect 1142 1111 1148 1112
rect 1142 1107 1143 1111
rect 1147 1107 1148 1111
rect 1142 1106 1148 1107
rect 1270 1111 1276 1112
rect 1270 1107 1271 1111
rect 1275 1107 1276 1111
rect 1270 1106 1276 1107
rect 1398 1111 1404 1112
rect 1398 1107 1399 1111
rect 1403 1107 1404 1111
rect 1766 1108 1767 1112
rect 1771 1108 1772 1112
rect 1766 1107 1772 1108
rect 1806 1108 1812 1109
rect 3462 1108 3468 1109
rect 1398 1106 1404 1107
rect 1806 1104 1807 1108
rect 1811 1104 1812 1108
rect 1806 1103 1812 1104
rect 1942 1107 1948 1108
rect 1942 1103 1943 1107
rect 1947 1103 1948 1107
rect 1942 1102 1948 1103
rect 2062 1107 2068 1108
rect 2062 1103 2063 1107
rect 2067 1103 2068 1107
rect 2062 1102 2068 1103
rect 2190 1107 2196 1108
rect 2190 1103 2191 1107
rect 2195 1103 2196 1107
rect 2190 1102 2196 1103
rect 2318 1107 2324 1108
rect 2318 1103 2319 1107
rect 2323 1103 2324 1107
rect 2318 1102 2324 1103
rect 2454 1107 2460 1108
rect 2454 1103 2455 1107
rect 2459 1103 2460 1107
rect 2454 1102 2460 1103
rect 2598 1107 2604 1108
rect 2598 1103 2599 1107
rect 2603 1103 2604 1107
rect 2598 1102 2604 1103
rect 2750 1107 2756 1108
rect 2750 1103 2751 1107
rect 2755 1103 2756 1107
rect 2750 1102 2756 1103
rect 2902 1107 2908 1108
rect 2902 1103 2903 1107
rect 2907 1103 2908 1107
rect 2902 1102 2908 1103
rect 3062 1107 3068 1108
rect 3062 1103 3063 1107
rect 3067 1103 3068 1107
rect 3062 1102 3068 1103
rect 3222 1107 3228 1108
rect 3222 1103 3223 1107
rect 3227 1103 3228 1107
rect 3222 1102 3228 1103
rect 3366 1107 3372 1108
rect 3366 1103 3367 1107
rect 3371 1103 3372 1107
rect 3462 1104 3463 1108
rect 3467 1104 3468 1108
rect 3462 1103 3468 1104
rect 3366 1102 3372 1103
rect 110 1095 116 1096
rect 110 1091 111 1095
rect 115 1091 116 1095
rect 1766 1095 1772 1096
rect 110 1090 116 1091
rect 246 1092 252 1093
rect 246 1088 247 1092
rect 251 1088 252 1092
rect 246 1087 252 1088
rect 366 1092 372 1093
rect 366 1088 367 1092
rect 371 1088 372 1092
rect 366 1087 372 1088
rect 494 1092 500 1093
rect 494 1088 495 1092
rect 499 1088 500 1092
rect 494 1087 500 1088
rect 622 1092 628 1093
rect 622 1088 623 1092
rect 627 1088 628 1092
rect 622 1087 628 1088
rect 758 1092 764 1093
rect 758 1088 759 1092
rect 763 1088 764 1092
rect 758 1087 764 1088
rect 886 1092 892 1093
rect 886 1088 887 1092
rect 891 1088 892 1092
rect 886 1087 892 1088
rect 1014 1092 1020 1093
rect 1014 1088 1015 1092
rect 1019 1088 1020 1092
rect 1014 1087 1020 1088
rect 1142 1092 1148 1093
rect 1142 1088 1143 1092
rect 1147 1088 1148 1092
rect 1142 1087 1148 1088
rect 1270 1092 1276 1093
rect 1270 1088 1271 1092
rect 1275 1088 1276 1092
rect 1270 1087 1276 1088
rect 1398 1092 1404 1093
rect 1398 1088 1399 1092
rect 1403 1088 1404 1092
rect 1766 1091 1767 1095
rect 1771 1091 1772 1095
rect 1766 1090 1772 1091
rect 1806 1091 1812 1092
rect 1398 1087 1404 1088
rect 1806 1087 1807 1091
rect 1811 1087 1812 1091
rect 3462 1091 3468 1092
rect 1806 1086 1812 1087
rect 1942 1088 1948 1089
rect 1942 1084 1943 1088
rect 1947 1084 1948 1088
rect 1942 1083 1948 1084
rect 2062 1088 2068 1089
rect 2062 1084 2063 1088
rect 2067 1084 2068 1088
rect 2062 1083 2068 1084
rect 2190 1088 2196 1089
rect 2190 1084 2191 1088
rect 2195 1084 2196 1088
rect 2190 1083 2196 1084
rect 2318 1088 2324 1089
rect 2318 1084 2319 1088
rect 2323 1084 2324 1088
rect 2318 1083 2324 1084
rect 2454 1088 2460 1089
rect 2454 1084 2455 1088
rect 2459 1084 2460 1088
rect 2454 1083 2460 1084
rect 2598 1088 2604 1089
rect 2598 1084 2599 1088
rect 2603 1084 2604 1088
rect 2598 1083 2604 1084
rect 2750 1088 2756 1089
rect 2750 1084 2751 1088
rect 2755 1084 2756 1088
rect 2750 1083 2756 1084
rect 2902 1088 2908 1089
rect 2902 1084 2903 1088
rect 2907 1084 2908 1088
rect 2902 1083 2908 1084
rect 3062 1088 3068 1089
rect 3062 1084 3063 1088
rect 3067 1084 3068 1088
rect 3062 1083 3068 1084
rect 3222 1088 3228 1089
rect 3222 1084 3223 1088
rect 3227 1084 3228 1088
rect 3222 1083 3228 1084
rect 3366 1088 3372 1089
rect 3366 1084 3367 1088
rect 3371 1084 3372 1088
rect 3462 1087 3463 1091
rect 3467 1087 3468 1091
rect 3462 1086 3468 1087
rect 3366 1083 3372 1084
rect 430 1044 436 1045
rect 110 1041 116 1042
rect 110 1037 111 1041
rect 115 1037 116 1041
rect 430 1040 431 1044
rect 435 1040 436 1044
rect 430 1039 436 1040
rect 542 1044 548 1045
rect 542 1040 543 1044
rect 547 1040 548 1044
rect 542 1039 548 1040
rect 662 1044 668 1045
rect 662 1040 663 1044
rect 667 1040 668 1044
rect 662 1039 668 1040
rect 790 1044 796 1045
rect 790 1040 791 1044
rect 795 1040 796 1044
rect 790 1039 796 1040
rect 918 1044 924 1045
rect 918 1040 919 1044
rect 923 1040 924 1044
rect 918 1039 924 1040
rect 1038 1044 1044 1045
rect 1038 1040 1039 1044
rect 1043 1040 1044 1044
rect 1038 1039 1044 1040
rect 1158 1044 1164 1045
rect 1158 1040 1159 1044
rect 1163 1040 1164 1044
rect 1158 1039 1164 1040
rect 1278 1044 1284 1045
rect 1278 1040 1279 1044
rect 1283 1040 1284 1044
rect 1278 1039 1284 1040
rect 1406 1044 1412 1045
rect 1406 1040 1407 1044
rect 1411 1040 1412 1044
rect 1406 1039 1412 1040
rect 1534 1044 1540 1045
rect 1534 1040 1535 1044
rect 1539 1040 1540 1044
rect 1534 1039 1540 1040
rect 1766 1041 1772 1042
rect 110 1036 116 1037
rect 1766 1037 1767 1041
rect 1771 1037 1772 1041
rect 1846 1040 1852 1041
rect 1766 1036 1772 1037
rect 1806 1037 1812 1038
rect 1806 1033 1807 1037
rect 1811 1033 1812 1037
rect 1846 1036 1847 1040
rect 1851 1036 1852 1040
rect 1846 1035 1852 1036
rect 1982 1040 1988 1041
rect 1982 1036 1983 1040
rect 1987 1036 1988 1040
rect 1982 1035 1988 1036
rect 2118 1040 2124 1041
rect 2118 1036 2119 1040
rect 2123 1036 2124 1040
rect 2118 1035 2124 1036
rect 2254 1040 2260 1041
rect 2254 1036 2255 1040
rect 2259 1036 2260 1040
rect 2254 1035 2260 1036
rect 2390 1040 2396 1041
rect 2390 1036 2391 1040
rect 2395 1036 2396 1040
rect 2390 1035 2396 1036
rect 2542 1040 2548 1041
rect 2542 1036 2543 1040
rect 2547 1036 2548 1040
rect 2542 1035 2548 1036
rect 2702 1040 2708 1041
rect 2702 1036 2703 1040
rect 2707 1036 2708 1040
rect 2702 1035 2708 1036
rect 2862 1040 2868 1041
rect 2862 1036 2863 1040
rect 2867 1036 2868 1040
rect 2862 1035 2868 1036
rect 3030 1040 3036 1041
rect 3030 1036 3031 1040
rect 3035 1036 3036 1040
rect 3030 1035 3036 1036
rect 3206 1040 3212 1041
rect 3206 1036 3207 1040
rect 3211 1036 3212 1040
rect 3206 1035 3212 1036
rect 3366 1040 3372 1041
rect 3366 1036 3367 1040
rect 3371 1036 3372 1040
rect 3366 1035 3372 1036
rect 3462 1037 3468 1038
rect 1806 1032 1812 1033
rect 3462 1033 3463 1037
rect 3467 1033 3468 1037
rect 3462 1032 3468 1033
rect 430 1025 436 1026
rect 110 1024 116 1025
rect 110 1020 111 1024
rect 115 1020 116 1024
rect 430 1021 431 1025
rect 435 1021 436 1025
rect 430 1020 436 1021
rect 542 1025 548 1026
rect 542 1021 543 1025
rect 547 1021 548 1025
rect 542 1020 548 1021
rect 662 1025 668 1026
rect 662 1021 663 1025
rect 667 1021 668 1025
rect 662 1020 668 1021
rect 790 1025 796 1026
rect 790 1021 791 1025
rect 795 1021 796 1025
rect 790 1020 796 1021
rect 918 1025 924 1026
rect 918 1021 919 1025
rect 923 1021 924 1025
rect 918 1020 924 1021
rect 1038 1025 1044 1026
rect 1038 1021 1039 1025
rect 1043 1021 1044 1025
rect 1038 1020 1044 1021
rect 1158 1025 1164 1026
rect 1158 1021 1159 1025
rect 1163 1021 1164 1025
rect 1158 1020 1164 1021
rect 1278 1025 1284 1026
rect 1278 1021 1279 1025
rect 1283 1021 1284 1025
rect 1278 1020 1284 1021
rect 1406 1025 1412 1026
rect 1406 1021 1407 1025
rect 1411 1021 1412 1025
rect 1406 1020 1412 1021
rect 1534 1025 1540 1026
rect 1534 1021 1535 1025
rect 1539 1021 1540 1025
rect 1534 1020 1540 1021
rect 1766 1024 1772 1025
rect 1766 1020 1767 1024
rect 1771 1020 1772 1024
rect 1846 1021 1852 1022
rect 110 1019 116 1020
rect 1766 1019 1772 1020
rect 1806 1020 1812 1021
rect 1806 1016 1807 1020
rect 1811 1016 1812 1020
rect 1846 1017 1847 1021
rect 1851 1017 1852 1021
rect 1846 1016 1852 1017
rect 1982 1021 1988 1022
rect 1982 1017 1983 1021
rect 1987 1017 1988 1021
rect 1982 1016 1988 1017
rect 2118 1021 2124 1022
rect 2118 1017 2119 1021
rect 2123 1017 2124 1021
rect 2118 1016 2124 1017
rect 2254 1021 2260 1022
rect 2254 1017 2255 1021
rect 2259 1017 2260 1021
rect 2254 1016 2260 1017
rect 2390 1021 2396 1022
rect 2390 1017 2391 1021
rect 2395 1017 2396 1021
rect 2390 1016 2396 1017
rect 2542 1021 2548 1022
rect 2542 1017 2543 1021
rect 2547 1017 2548 1021
rect 2542 1016 2548 1017
rect 2702 1021 2708 1022
rect 2702 1017 2703 1021
rect 2707 1017 2708 1021
rect 2702 1016 2708 1017
rect 2862 1021 2868 1022
rect 2862 1017 2863 1021
rect 2867 1017 2868 1021
rect 2862 1016 2868 1017
rect 3030 1021 3036 1022
rect 3030 1017 3031 1021
rect 3035 1017 3036 1021
rect 3030 1016 3036 1017
rect 3206 1021 3212 1022
rect 3206 1017 3207 1021
rect 3211 1017 3212 1021
rect 3206 1016 3212 1017
rect 3366 1021 3372 1022
rect 3366 1017 3367 1021
rect 3371 1017 3372 1021
rect 3366 1016 3372 1017
rect 3462 1020 3468 1021
rect 3462 1016 3463 1020
rect 3467 1016 3468 1020
rect 1806 1015 1812 1016
rect 3462 1015 3468 1016
rect 110 972 116 973
rect 1766 972 1772 973
rect 110 968 111 972
rect 115 968 116 972
rect 110 967 116 968
rect 566 971 572 972
rect 566 967 567 971
rect 571 967 572 971
rect 566 966 572 967
rect 678 971 684 972
rect 678 967 679 971
rect 683 967 684 971
rect 678 966 684 967
rect 790 971 796 972
rect 790 967 791 971
rect 795 967 796 971
rect 790 966 796 967
rect 910 971 916 972
rect 910 967 911 971
rect 915 967 916 971
rect 910 966 916 967
rect 1030 971 1036 972
rect 1030 967 1031 971
rect 1035 967 1036 971
rect 1030 966 1036 967
rect 1142 971 1148 972
rect 1142 967 1143 971
rect 1147 967 1148 971
rect 1142 966 1148 967
rect 1254 971 1260 972
rect 1254 967 1255 971
rect 1259 967 1260 971
rect 1254 966 1260 967
rect 1358 971 1364 972
rect 1358 967 1359 971
rect 1363 967 1364 971
rect 1358 966 1364 967
rect 1470 971 1476 972
rect 1470 967 1471 971
rect 1475 967 1476 971
rect 1470 966 1476 967
rect 1582 971 1588 972
rect 1582 967 1583 971
rect 1587 967 1588 971
rect 1582 966 1588 967
rect 1670 971 1676 972
rect 1670 967 1671 971
rect 1675 967 1676 971
rect 1766 968 1767 972
rect 1771 968 1772 972
rect 1766 967 1772 968
rect 1806 972 1812 973
rect 3462 972 3468 973
rect 1806 968 1807 972
rect 1811 968 1812 972
rect 1806 967 1812 968
rect 1830 971 1836 972
rect 1830 967 1831 971
rect 1835 967 1836 971
rect 1670 966 1676 967
rect 1830 966 1836 967
rect 1974 971 1980 972
rect 1974 967 1975 971
rect 1979 967 1980 971
rect 1974 966 1980 967
rect 2134 971 2140 972
rect 2134 967 2135 971
rect 2139 967 2140 971
rect 2134 966 2140 967
rect 2294 971 2300 972
rect 2294 967 2295 971
rect 2299 967 2300 971
rect 2294 966 2300 967
rect 2462 971 2468 972
rect 2462 967 2463 971
rect 2467 967 2468 971
rect 2462 966 2468 967
rect 2630 971 2636 972
rect 2630 967 2631 971
rect 2635 967 2636 971
rect 2630 966 2636 967
rect 2806 971 2812 972
rect 2806 967 2807 971
rect 2811 967 2812 971
rect 2806 966 2812 967
rect 2990 971 2996 972
rect 2990 967 2991 971
rect 2995 967 2996 971
rect 2990 966 2996 967
rect 3182 971 3188 972
rect 3182 967 3183 971
rect 3187 967 3188 971
rect 3182 966 3188 967
rect 3366 971 3372 972
rect 3366 967 3367 971
rect 3371 967 3372 971
rect 3462 968 3463 972
rect 3467 968 3468 972
rect 3462 967 3468 968
rect 3366 966 3372 967
rect 110 955 116 956
rect 110 951 111 955
rect 115 951 116 955
rect 1766 955 1772 956
rect 110 950 116 951
rect 566 952 572 953
rect 566 948 567 952
rect 571 948 572 952
rect 566 947 572 948
rect 678 952 684 953
rect 678 948 679 952
rect 683 948 684 952
rect 678 947 684 948
rect 790 952 796 953
rect 790 948 791 952
rect 795 948 796 952
rect 790 947 796 948
rect 910 952 916 953
rect 910 948 911 952
rect 915 948 916 952
rect 910 947 916 948
rect 1030 952 1036 953
rect 1030 948 1031 952
rect 1035 948 1036 952
rect 1030 947 1036 948
rect 1142 952 1148 953
rect 1142 948 1143 952
rect 1147 948 1148 952
rect 1142 947 1148 948
rect 1254 952 1260 953
rect 1254 948 1255 952
rect 1259 948 1260 952
rect 1254 947 1260 948
rect 1358 952 1364 953
rect 1358 948 1359 952
rect 1363 948 1364 952
rect 1358 947 1364 948
rect 1470 952 1476 953
rect 1470 948 1471 952
rect 1475 948 1476 952
rect 1470 947 1476 948
rect 1582 952 1588 953
rect 1582 948 1583 952
rect 1587 948 1588 952
rect 1582 947 1588 948
rect 1670 952 1676 953
rect 1670 948 1671 952
rect 1675 948 1676 952
rect 1766 951 1767 955
rect 1771 951 1772 955
rect 1766 950 1772 951
rect 1806 955 1812 956
rect 1806 951 1807 955
rect 1811 951 1812 955
rect 3462 955 3468 956
rect 1806 950 1812 951
rect 1830 952 1836 953
rect 1670 947 1676 948
rect 1830 948 1831 952
rect 1835 948 1836 952
rect 1830 947 1836 948
rect 1974 952 1980 953
rect 1974 948 1975 952
rect 1979 948 1980 952
rect 1974 947 1980 948
rect 2134 952 2140 953
rect 2134 948 2135 952
rect 2139 948 2140 952
rect 2134 947 2140 948
rect 2294 952 2300 953
rect 2294 948 2295 952
rect 2299 948 2300 952
rect 2294 947 2300 948
rect 2462 952 2468 953
rect 2462 948 2463 952
rect 2467 948 2468 952
rect 2462 947 2468 948
rect 2630 952 2636 953
rect 2630 948 2631 952
rect 2635 948 2636 952
rect 2630 947 2636 948
rect 2806 952 2812 953
rect 2806 948 2807 952
rect 2811 948 2812 952
rect 2806 947 2812 948
rect 2990 952 2996 953
rect 2990 948 2991 952
rect 2995 948 2996 952
rect 2990 947 2996 948
rect 3182 952 3188 953
rect 3182 948 3183 952
rect 3187 948 3188 952
rect 3182 947 3188 948
rect 3366 952 3372 953
rect 3366 948 3367 952
rect 3371 948 3372 952
rect 3462 951 3463 955
rect 3467 951 3468 955
rect 3462 950 3468 951
rect 3366 947 3372 948
rect 2126 908 2132 909
rect 1806 905 1812 906
rect 414 904 420 905
rect 110 901 116 902
rect 110 897 111 901
rect 115 897 116 901
rect 414 900 415 904
rect 419 900 420 904
rect 414 899 420 900
rect 558 904 564 905
rect 558 900 559 904
rect 563 900 564 904
rect 558 899 564 900
rect 726 904 732 905
rect 726 900 727 904
rect 731 900 732 904
rect 726 899 732 900
rect 910 904 916 905
rect 910 900 911 904
rect 915 900 916 904
rect 910 899 916 900
rect 1118 904 1124 905
rect 1118 900 1119 904
rect 1123 900 1124 904
rect 1118 899 1124 900
rect 1334 904 1340 905
rect 1334 900 1335 904
rect 1339 900 1340 904
rect 1334 899 1340 900
rect 1558 904 1564 905
rect 1558 900 1559 904
rect 1563 900 1564 904
rect 1558 899 1564 900
rect 1766 901 1772 902
rect 110 896 116 897
rect 1766 897 1767 901
rect 1771 897 1772 901
rect 1806 901 1807 905
rect 1811 901 1812 905
rect 2126 904 2127 908
rect 2131 904 2132 908
rect 2126 903 2132 904
rect 2214 908 2220 909
rect 2214 904 2215 908
rect 2219 904 2220 908
rect 2214 903 2220 904
rect 2302 908 2308 909
rect 2302 904 2303 908
rect 2307 904 2308 908
rect 2302 903 2308 904
rect 2390 908 2396 909
rect 2390 904 2391 908
rect 2395 904 2396 908
rect 2390 903 2396 904
rect 2478 908 2484 909
rect 2478 904 2479 908
rect 2483 904 2484 908
rect 2478 903 2484 904
rect 2566 908 2572 909
rect 2566 904 2567 908
rect 2571 904 2572 908
rect 2566 903 2572 904
rect 2654 908 2660 909
rect 2654 904 2655 908
rect 2659 904 2660 908
rect 2654 903 2660 904
rect 2742 908 2748 909
rect 2742 904 2743 908
rect 2747 904 2748 908
rect 2742 903 2748 904
rect 2830 908 2836 909
rect 2830 904 2831 908
rect 2835 904 2836 908
rect 2830 903 2836 904
rect 3462 905 3468 906
rect 1806 900 1812 901
rect 3462 901 3463 905
rect 3467 901 3468 905
rect 3462 900 3468 901
rect 1766 896 1772 897
rect 2126 889 2132 890
rect 1806 888 1812 889
rect 414 885 420 886
rect 110 884 116 885
rect 110 880 111 884
rect 115 880 116 884
rect 414 881 415 885
rect 419 881 420 885
rect 414 880 420 881
rect 558 885 564 886
rect 558 881 559 885
rect 563 881 564 885
rect 558 880 564 881
rect 726 885 732 886
rect 726 881 727 885
rect 731 881 732 885
rect 726 880 732 881
rect 910 885 916 886
rect 910 881 911 885
rect 915 881 916 885
rect 910 880 916 881
rect 1118 885 1124 886
rect 1118 881 1119 885
rect 1123 881 1124 885
rect 1118 880 1124 881
rect 1334 885 1340 886
rect 1334 881 1335 885
rect 1339 881 1340 885
rect 1334 880 1340 881
rect 1558 885 1564 886
rect 1558 881 1559 885
rect 1563 881 1564 885
rect 1558 880 1564 881
rect 1766 884 1772 885
rect 1766 880 1767 884
rect 1771 880 1772 884
rect 1806 884 1807 888
rect 1811 884 1812 888
rect 2126 885 2127 889
rect 2131 885 2132 889
rect 2126 884 2132 885
rect 2214 889 2220 890
rect 2214 885 2215 889
rect 2219 885 2220 889
rect 2214 884 2220 885
rect 2302 889 2308 890
rect 2302 885 2303 889
rect 2307 885 2308 889
rect 2302 884 2308 885
rect 2390 889 2396 890
rect 2390 885 2391 889
rect 2395 885 2396 889
rect 2390 884 2396 885
rect 2478 889 2484 890
rect 2478 885 2479 889
rect 2483 885 2484 889
rect 2478 884 2484 885
rect 2566 889 2572 890
rect 2566 885 2567 889
rect 2571 885 2572 889
rect 2566 884 2572 885
rect 2654 889 2660 890
rect 2654 885 2655 889
rect 2659 885 2660 889
rect 2654 884 2660 885
rect 2742 889 2748 890
rect 2742 885 2743 889
rect 2747 885 2748 889
rect 2742 884 2748 885
rect 2830 889 2836 890
rect 2830 885 2831 889
rect 2835 885 2836 889
rect 2830 884 2836 885
rect 3462 888 3468 889
rect 3462 884 3463 888
rect 3467 884 3468 888
rect 1806 883 1812 884
rect 3462 883 3468 884
rect 110 879 116 880
rect 1766 879 1772 880
rect 110 836 116 837
rect 1766 836 1772 837
rect 110 832 111 836
rect 115 832 116 836
rect 110 831 116 832
rect 134 835 140 836
rect 134 831 135 835
rect 139 831 140 835
rect 134 830 140 831
rect 230 835 236 836
rect 230 831 231 835
rect 235 831 236 835
rect 230 830 236 831
rect 358 835 364 836
rect 358 831 359 835
rect 363 831 364 835
rect 358 830 364 831
rect 486 835 492 836
rect 486 831 487 835
rect 491 831 492 835
rect 486 830 492 831
rect 622 835 628 836
rect 622 831 623 835
rect 627 831 628 835
rect 622 830 628 831
rect 750 835 756 836
rect 750 831 751 835
rect 755 831 756 835
rect 750 830 756 831
rect 878 835 884 836
rect 878 831 879 835
rect 883 831 884 835
rect 878 830 884 831
rect 1006 835 1012 836
rect 1006 831 1007 835
rect 1011 831 1012 835
rect 1006 830 1012 831
rect 1134 835 1140 836
rect 1134 831 1135 835
rect 1139 831 1140 835
rect 1134 830 1140 831
rect 1270 835 1276 836
rect 1270 831 1271 835
rect 1275 831 1276 835
rect 1766 832 1767 836
rect 1771 832 1772 836
rect 1766 831 1772 832
rect 1806 836 1812 837
rect 3462 836 3468 837
rect 1806 832 1807 836
rect 1811 832 1812 836
rect 1806 831 1812 832
rect 2158 835 2164 836
rect 2158 831 2159 835
rect 2163 831 2164 835
rect 1270 830 1276 831
rect 2158 830 2164 831
rect 2246 835 2252 836
rect 2246 831 2247 835
rect 2251 831 2252 835
rect 2246 830 2252 831
rect 2334 835 2340 836
rect 2334 831 2335 835
rect 2339 831 2340 835
rect 2334 830 2340 831
rect 2422 835 2428 836
rect 2422 831 2423 835
rect 2427 831 2428 835
rect 2422 830 2428 831
rect 2526 835 2532 836
rect 2526 831 2527 835
rect 2531 831 2532 835
rect 2526 830 2532 831
rect 2638 835 2644 836
rect 2638 831 2639 835
rect 2643 831 2644 835
rect 2638 830 2644 831
rect 2766 835 2772 836
rect 2766 831 2767 835
rect 2771 831 2772 835
rect 2766 830 2772 831
rect 2910 835 2916 836
rect 2910 831 2911 835
rect 2915 831 2916 835
rect 2910 830 2916 831
rect 3062 835 3068 836
rect 3062 831 3063 835
rect 3067 831 3068 835
rect 3062 830 3068 831
rect 3222 835 3228 836
rect 3222 831 3223 835
rect 3227 831 3228 835
rect 3222 830 3228 831
rect 3366 835 3372 836
rect 3366 831 3367 835
rect 3371 831 3372 835
rect 3462 832 3463 836
rect 3467 832 3468 836
rect 3462 831 3468 832
rect 3366 830 3372 831
rect 110 819 116 820
rect 110 815 111 819
rect 115 815 116 819
rect 1766 819 1772 820
rect 110 814 116 815
rect 134 816 140 817
rect 134 812 135 816
rect 139 812 140 816
rect 134 811 140 812
rect 230 816 236 817
rect 230 812 231 816
rect 235 812 236 816
rect 230 811 236 812
rect 358 816 364 817
rect 358 812 359 816
rect 363 812 364 816
rect 358 811 364 812
rect 486 816 492 817
rect 486 812 487 816
rect 491 812 492 816
rect 486 811 492 812
rect 622 816 628 817
rect 622 812 623 816
rect 627 812 628 816
rect 622 811 628 812
rect 750 816 756 817
rect 750 812 751 816
rect 755 812 756 816
rect 750 811 756 812
rect 878 816 884 817
rect 878 812 879 816
rect 883 812 884 816
rect 878 811 884 812
rect 1006 816 1012 817
rect 1006 812 1007 816
rect 1011 812 1012 816
rect 1006 811 1012 812
rect 1134 816 1140 817
rect 1134 812 1135 816
rect 1139 812 1140 816
rect 1134 811 1140 812
rect 1270 816 1276 817
rect 1270 812 1271 816
rect 1275 812 1276 816
rect 1766 815 1767 819
rect 1771 815 1772 819
rect 1766 814 1772 815
rect 1806 819 1812 820
rect 1806 815 1807 819
rect 1811 815 1812 819
rect 3462 819 3468 820
rect 1806 814 1812 815
rect 2158 816 2164 817
rect 1270 811 1276 812
rect 2158 812 2159 816
rect 2163 812 2164 816
rect 2158 811 2164 812
rect 2246 816 2252 817
rect 2246 812 2247 816
rect 2251 812 2252 816
rect 2246 811 2252 812
rect 2334 816 2340 817
rect 2334 812 2335 816
rect 2339 812 2340 816
rect 2334 811 2340 812
rect 2422 816 2428 817
rect 2422 812 2423 816
rect 2427 812 2428 816
rect 2422 811 2428 812
rect 2526 816 2532 817
rect 2526 812 2527 816
rect 2531 812 2532 816
rect 2526 811 2532 812
rect 2638 816 2644 817
rect 2638 812 2639 816
rect 2643 812 2644 816
rect 2638 811 2644 812
rect 2766 816 2772 817
rect 2766 812 2767 816
rect 2771 812 2772 816
rect 2766 811 2772 812
rect 2910 816 2916 817
rect 2910 812 2911 816
rect 2915 812 2916 816
rect 2910 811 2916 812
rect 3062 816 3068 817
rect 3062 812 3063 816
rect 3067 812 3068 816
rect 3062 811 3068 812
rect 3222 816 3228 817
rect 3222 812 3223 816
rect 3227 812 3228 816
rect 3222 811 3228 812
rect 3366 816 3372 817
rect 3366 812 3367 816
rect 3371 812 3372 816
rect 3462 815 3463 819
rect 3467 815 3468 819
rect 3462 814 3468 815
rect 3366 811 3372 812
rect 134 768 140 769
rect 110 765 116 766
rect 110 761 111 765
rect 115 761 116 765
rect 134 764 135 768
rect 139 764 140 768
rect 134 763 140 764
rect 222 768 228 769
rect 222 764 223 768
rect 227 764 228 768
rect 222 763 228 764
rect 342 768 348 769
rect 342 764 343 768
rect 347 764 348 768
rect 342 763 348 764
rect 470 768 476 769
rect 470 764 471 768
rect 475 764 476 768
rect 470 763 476 764
rect 606 768 612 769
rect 606 764 607 768
rect 611 764 612 768
rect 606 763 612 764
rect 742 768 748 769
rect 742 764 743 768
rect 747 764 748 768
rect 742 763 748 764
rect 886 768 892 769
rect 886 764 887 768
rect 891 764 892 768
rect 886 763 892 764
rect 1038 768 1044 769
rect 1038 764 1039 768
rect 1043 764 1044 768
rect 1038 763 1044 764
rect 1190 768 1196 769
rect 1190 764 1191 768
rect 1195 764 1196 768
rect 1190 763 1196 764
rect 1350 768 1356 769
rect 1350 764 1351 768
rect 1355 764 1356 768
rect 2062 768 2068 769
rect 1350 763 1356 764
rect 1766 765 1772 766
rect 110 760 116 761
rect 1766 761 1767 765
rect 1771 761 1772 765
rect 1766 760 1772 761
rect 1806 765 1812 766
rect 1806 761 1807 765
rect 1811 761 1812 765
rect 2062 764 2063 768
rect 2067 764 2068 768
rect 2062 763 2068 764
rect 2174 768 2180 769
rect 2174 764 2175 768
rect 2179 764 2180 768
rect 2174 763 2180 764
rect 2294 768 2300 769
rect 2294 764 2295 768
rect 2299 764 2300 768
rect 2294 763 2300 764
rect 2422 768 2428 769
rect 2422 764 2423 768
rect 2427 764 2428 768
rect 2422 763 2428 764
rect 2558 768 2564 769
rect 2558 764 2559 768
rect 2563 764 2564 768
rect 2558 763 2564 764
rect 2710 768 2716 769
rect 2710 764 2711 768
rect 2715 764 2716 768
rect 2710 763 2716 764
rect 2870 768 2876 769
rect 2870 764 2871 768
rect 2875 764 2876 768
rect 2870 763 2876 764
rect 3038 768 3044 769
rect 3038 764 3039 768
rect 3043 764 3044 768
rect 3038 763 3044 764
rect 3214 768 3220 769
rect 3214 764 3215 768
rect 3219 764 3220 768
rect 3214 763 3220 764
rect 3366 768 3372 769
rect 3366 764 3367 768
rect 3371 764 3372 768
rect 3366 763 3372 764
rect 3462 765 3468 766
rect 1806 760 1812 761
rect 3462 761 3463 765
rect 3467 761 3468 765
rect 3462 760 3468 761
rect 134 749 140 750
rect 110 748 116 749
rect 110 744 111 748
rect 115 744 116 748
rect 134 745 135 749
rect 139 745 140 749
rect 134 744 140 745
rect 222 749 228 750
rect 222 745 223 749
rect 227 745 228 749
rect 222 744 228 745
rect 342 749 348 750
rect 342 745 343 749
rect 347 745 348 749
rect 342 744 348 745
rect 470 749 476 750
rect 470 745 471 749
rect 475 745 476 749
rect 470 744 476 745
rect 606 749 612 750
rect 606 745 607 749
rect 611 745 612 749
rect 606 744 612 745
rect 742 749 748 750
rect 742 745 743 749
rect 747 745 748 749
rect 742 744 748 745
rect 886 749 892 750
rect 886 745 887 749
rect 891 745 892 749
rect 886 744 892 745
rect 1038 749 1044 750
rect 1038 745 1039 749
rect 1043 745 1044 749
rect 1038 744 1044 745
rect 1190 749 1196 750
rect 1190 745 1191 749
rect 1195 745 1196 749
rect 1190 744 1196 745
rect 1350 749 1356 750
rect 2062 749 2068 750
rect 1350 745 1351 749
rect 1355 745 1356 749
rect 1350 744 1356 745
rect 1766 748 1772 749
rect 1766 744 1767 748
rect 1771 744 1772 748
rect 110 743 116 744
rect 1766 743 1772 744
rect 1806 748 1812 749
rect 1806 744 1807 748
rect 1811 744 1812 748
rect 2062 745 2063 749
rect 2067 745 2068 749
rect 2062 744 2068 745
rect 2174 749 2180 750
rect 2174 745 2175 749
rect 2179 745 2180 749
rect 2174 744 2180 745
rect 2294 749 2300 750
rect 2294 745 2295 749
rect 2299 745 2300 749
rect 2294 744 2300 745
rect 2422 749 2428 750
rect 2422 745 2423 749
rect 2427 745 2428 749
rect 2422 744 2428 745
rect 2558 749 2564 750
rect 2558 745 2559 749
rect 2563 745 2564 749
rect 2558 744 2564 745
rect 2710 749 2716 750
rect 2710 745 2711 749
rect 2715 745 2716 749
rect 2710 744 2716 745
rect 2870 749 2876 750
rect 2870 745 2871 749
rect 2875 745 2876 749
rect 2870 744 2876 745
rect 3038 749 3044 750
rect 3038 745 3039 749
rect 3043 745 3044 749
rect 3038 744 3044 745
rect 3214 749 3220 750
rect 3214 745 3215 749
rect 3219 745 3220 749
rect 3214 744 3220 745
rect 3366 749 3372 750
rect 3366 745 3367 749
rect 3371 745 3372 749
rect 3366 744 3372 745
rect 3462 748 3468 749
rect 3462 744 3463 748
rect 3467 744 3468 748
rect 1806 743 1812 744
rect 3462 743 3468 744
rect 1806 704 1812 705
rect 3462 704 3468 705
rect 110 700 116 701
rect 1766 700 1772 701
rect 110 696 111 700
rect 115 696 116 700
rect 110 695 116 696
rect 166 699 172 700
rect 166 695 167 699
rect 171 695 172 699
rect 166 694 172 695
rect 294 699 300 700
rect 294 695 295 699
rect 299 695 300 699
rect 294 694 300 695
rect 430 699 436 700
rect 430 695 431 699
rect 435 695 436 699
rect 430 694 436 695
rect 574 699 580 700
rect 574 695 575 699
rect 579 695 580 699
rect 574 694 580 695
rect 726 699 732 700
rect 726 695 727 699
rect 731 695 732 699
rect 726 694 732 695
rect 878 699 884 700
rect 878 695 879 699
rect 883 695 884 699
rect 878 694 884 695
rect 1030 699 1036 700
rect 1030 695 1031 699
rect 1035 695 1036 699
rect 1030 694 1036 695
rect 1182 699 1188 700
rect 1182 695 1183 699
rect 1187 695 1188 699
rect 1182 694 1188 695
rect 1342 699 1348 700
rect 1342 695 1343 699
rect 1347 695 1348 699
rect 1342 694 1348 695
rect 1502 699 1508 700
rect 1502 695 1503 699
rect 1507 695 1508 699
rect 1766 696 1767 700
rect 1771 696 1772 700
rect 1806 700 1807 704
rect 1811 700 1812 704
rect 1806 699 1812 700
rect 1926 703 1932 704
rect 1926 699 1927 703
rect 1931 699 1932 703
rect 1926 698 1932 699
rect 2070 703 2076 704
rect 2070 699 2071 703
rect 2075 699 2076 703
rect 2070 698 2076 699
rect 2230 703 2236 704
rect 2230 699 2231 703
rect 2235 699 2236 703
rect 2230 698 2236 699
rect 2390 703 2396 704
rect 2390 699 2391 703
rect 2395 699 2396 703
rect 2390 698 2396 699
rect 2550 703 2556 704
rect 2550 699 2551 703
rect 2555 699 2556 703
rect 2550 698 2556 699
rect 2702 703 2708 704
rect 2702 699 2703 703
rect 2707 699 2708 703
rect 2702 698 2708 699
rect 2846 703 2852 704
rect 2846 699 2847 703
rect 2851 699 2852 703
rect 2846 698 2852 699
rect 2982 703 2988 704
rect 2982 699 2983 703
rect 2987 699 2988 703
rect 2982 698 2988 699
rect 3118 703 3124 704
rect 3118 699 3119 703
rect 3123 699 3124 703
rect 3118 698 3124 699
rect 3254 703 3260 704
rect 3254 699 3255 703
rect 3259 699 3260 703
rect 3254 698 3260 699
rect 3366 703 3372 704
rect 3366 699 3367 703
rect 3371 699 3372 703
rect 3462 700 3463 704
rect 3467 700 3468 704
rect 3462 699 3468 700
rect 3366 698 3372 699
rect 1766 695 1772 696
rect 1502 694 1508 695
rect 1806 687 1812 688
rect 110 683 116 684
rect 110 679 111 683
rect 115 679 116 683
rect 1766 683 1772 684
rect 110 678 116 679
rect 166 680 172 681
rect 166 676 167 680
rect 171 676 172 680
rect 166 675 172 676
rect 294 680 300 681
rect 294 676 295 680
rect 299 676 300 680
rect 294 675 300 676
rect 430 680 436 681
rect 430 676 431 680
rect 435 676 436 680
rect 430 675 436 676
rect 574 680 580 681
rect 574 676 575 680
rect 579 676 580 680
rect 574 675 580 676
rect 726 680 732 681
rect 726 676 727 680
rect 731 676 732 680
rect 726 675 732 676
rect 878 680 884 681
rect 878 676 879 680
rect 883 676 884 680
rect 878 675 884 676
rect 1030 680 1036 681
rect 1030 676 1031 680
rect 1035 676 1036 680
rect 1030 675 1036 676
rect 1182 680 1188 681
rect 1182 676 1183 680
rect 1187 676 1188 680
rect 1182 675 1188 676
rect 1342 680 1348 681
rect 1342 676 1343 680
rect 1347 676 1348 680
rect 1342 675 1348 676
rect 1502 680 1508 681
rect 1502 676 1503 680
rect 1507 676 1508 680
rect 1766 679 1767 683
rect 1771 679 1772 683
rect 1806 683 1807 687
rect 1811 683 1812 687
rect 3462 687 3468 688
rect 1806 682 1812 683
rect 1926 684 1932 685
rect 1926 680 1927 684
rect 1931 680 1932 684
rect 1926 679 1932 680
rect 2070 684 2076 685
rect 2070 680 2071 684
rect 2075 680 2076 684
rect 2070 679 2076 680
rect 2230 684 2236 685
rect 2230 680 2231 684
rect 2235 680 2236 684
rect 2230 679 2236 680
rect 2390 684 2396 685
rect 2390 680 2391 684
rect 2395 680 2396 684
rect 2390 679 2396 680
rect 2550 684 2556 685
rect 2550 680 2551 684
rect 2555 680 2556 684
rect 2550 679 2556 680
rect 2702 684 2708 685
rect 2702 680 2703 684
rect 2707 680 2708 684
rect 2702 679 2708 680
rect 2846 684 2852 685
rect 2846 680 2847 684
rect 2851 680 2852 684
rect 2846 679 2852 680
rect 2982 684 2988 685
rect 2982 680 2983 684
rect 2987 680 2988 684
rect 2982 679 2988 680
rect 3118 684 3124 685
rect 3118 680 3119 684
rect 3123 680 3124 684
rect 3118 679 3124 680
rect 3254 684 3260 685
rect 3254 680 3255 684
rect 3259 680 3260 684
rect 3254 679 3260 680
rect 3366 684 3372 685
rect 3366 680 3367 684
rect 3371 680 3372 684
rect 3462 683 3463 687
rect 3467 683 3468 687
rect 3462 682 3468 683
rect 3366 679 3372 680
rect 1766 678 1772 679
rect 1502 675 1508 676
rect 454 632 460 633
rect 110 629 116 630
rect 110 625 111 629
rect 115 625 116 629
rect 454 628 455 632
rect 459 628 460 632
rect 454 627 460 628
rect 558 632 564 633
rect 558 628 559 632
rect 563 628 564 632
rect 558 627 564 628
rect 678 632 684 633
rect 678 628 679 632
rect 683 628 684 632
rect 678 627 684 628
rect 798 632 804 633
rect 798 628 799 632
rect 803 628 804 632
rect 798 627 804 628
rect 926 632 932 633
rect 926 628 927 632
rect 931 628 932 632
rect 926 627 932 628
rect 1054 632 1060 633
rect 1054 628 1055 632
rect 1059 628 1060 632
rect 1054 627 1060 628
rect 1182 632 1188 633
rect 1182 628 1183 632
rect 1187 628 1188 632
rect 1182 627 1188 628
rect 1310 632 1316 633
rect 1310 628 1311 632
rect 1315 628 1316 632
rect 1310 627 1316 628
rect 1446 632 1452 633
rect 1446 628 1447 632
rect 1451 628 1452 632
rect 1446 627 1452 628
rect 1582 632 1588 633
rect 1582 628 1583 632
rect 1587 628 1588 632
rect 1830 632 1836 633
rect 1582 627 1588 628
rect 1766 629 1772 630
rect 110 624 116 625
rect 1766 625 1767 629
rect 1771 625 1772 629
rect 1766 624 1772 625
rect 1806 629 1812 630
rect 1806 625 1807 629
rect 1811 625 1812 629
rect 1830 628 1831 632
rect 1835 628 1836 632
rect 1830 627 1836 628
rect 1966 632 1972 633
rect 1966 628 1967 632
rect 1971 628 1972 632
rect 1966 627 1972 628
rect 2134 632 2140 633
rect 2134 628 2135 632
rect 2139 628 2140 632
rect 2134 627 2140 628
rect 2310 632 2316 633
rect 2310 628 2311 632
rect 2315 628 2316 632
rect 2310 627 2316 628
rect 2486 632 2492 633
rect 2486 628 2487 632
rect 2491 628 2492 632
rect 2486 627 2492 628
rect 2654 632 2660 633
rect 2654 628 2655 632
rect 2659 628 2660 632
rect 2654 627 2660 628
rect 2814 632 2820 633
rect 2814 628 2815 632
rect 2819 628 2820 632
rect 2814 627 2820 628
rect 2958 632 2964 633
rect 2958 628 2959 632
rect 2963 628 2964 632
rect 2958 627 2964 628
rect 3102 632 3108 633
rect 3102 628 3103 632
rect 3107 628 3108 632
rect 3102 627 3108 628
rect 3246 632 3252 633
rect 3246 628 3247 632
rect 3251 628 3252 632
rect 3246 627 3252 628
rect 3366 632 3372 633
rect 3366 628 3367 632
rect 3371 628 3372 632
rect 3366 627 3372 628
rect 3462 629 3468 630
rect 1806 624 1812 625
rect 3462 625 3463 629
rect 3467 625 3468 629
rect 3462 624 3468 625
rect 454 613 460 614
rect 110 612 116 613
rect 110 608 111 612
rect 115 608 116 612
rect 454 609 455 613
rect 459 609 460 613
rect 454 608 460 609
rect 558 613 564 614
rect 558 609 559 613
rect 563 609 564 613
rect 558 608 564 609
rect 678 613 684 614
rect 678 609 679 613
rect 683 609 684 613
rect 678 608 684 609
rect 798 613 804 614
rect 798 609 799 613
rect 803 609 804 613
rect 798 608 804 609
rect 926 613 932 614
rect 926 609 927 613
rect 931 609 932 613
rect 926 608 932 609
rect 1054 613 1060 614
rect 1054 609 1055 613
rect 1059 609 1060 613
rect 1054 608 1060 609
rect 1182 613 1188 614
rect 1182 609 1183 613
rect 1187 609 1188 613
rect 1182 608 1188 609
rect 1310 613 1316 614
rect 1310 609 1311 613
rect 1315 609 1316 613
rect 1310 608 1316 609
rect 1446 613 1452 614
rect 1446 609 1447 613
rect 1451 609 1452 613
rect 1446 608 1452 609
rect 1582 613 1588 614
rect 1830 613 1836 614
rect 1582 609 1583 613
rect 1587 609 1588 613
rect 1582 608 1588 609
rect 1766 612 1772 613
rect 1766 608 1767 612
rect 1771 608 1772 612
rect 110 607 116 608
rect 1766 607 1772 608
rect 1806 612 1812 613
rect 1806 608 1807 612
rect 1811 608 1812 612
rect 1830 609 1831 613
rect 1835 609 1836 613
rect 1830 608 1836 609
rect 1966 613 1972 614
rect 1966 609 1967 613
rect 1971 609 1972 613
rect 1966 608 1972 609
rect 2134 613 2140 614
rect 2134 609 2135 613
rect 2139 609 2140 613
rect 2134 608 2140 609
rect 2310 613 2316 614
rect 2310 609 2311 613
rect 2315 609 2316 613
rect 2310 608 2316 609
rect 2486 613 2492 614
rect 2486 609 2487 613
rect 2491 609 2492 613
rect 2486 608 2492 609
rect 2654 613 2660 614
rect 2654 609 2655 613
rect 2659 609 2660 613
rect 2654 608 2660 609
rect 2814 613 2820 614
rect 2814 609 2815 613
rect 2819 609 2820 613
rect 2814 608 2820 609
rect 2958 613 2964 614
rect 2958 609 2959 613
rect 2963 609 2964 613
rect 2958 608 2964 609
rect 3102 613 3108 614
rect 3102 609 3103 613
rect 3107 609 3108 613
rect 3102 608 3108 609
rect 3246 613 3252 614
rect 3246 609 3247 613
rect 3251 609 3252 613
rect 3246 608 3252 609
rect 3366 613 3372 614
rect 3366 609 3367 613
rect 3371 609 3372 613
rect 3366 608 3372 609
rect 3462 612 3468 613
rect 3462 608 3463 612
rect 3467 608 3468 612
rect 1806 607 1812 608
rect 3462 607 3468 608
rect 1806 568 1812 569
rect 3462 568 3468 569
rect 1806 564 1807 568
rect 1811 564 1812 568
rect 1806 563 1812 564
rect 1830 567 1836 568
rect 1830 563 1831 567
rect 1835 563 1836 567
rect 1830 562 1836 563
rect 1966 567 1972 568
rect 1966 563 1967 567
rect 1971 563 1972 567
rect 1966 562 1972 563
rect 2126 567 2132 568
rect 2126 563 2127 567
rect 2131 563 2132 567
rect 2126 562 2132 563
rect 2286 567 2292 568
rect 2286 563 2287 567
rect 2291 563 2292 567
rect 2286 562 2292 563
rect 2454 567 2460 568
rect 2454 563 2455 567
rect 2459 563 2460 567
rect 2454 562 2460 563
rect 2622 567 2628 568
rect 2622 563 2623 567
rect 2627 563 2628 567
rect 2622 562 2628 563
rect 2798 567 2804 568
rect 2798 563 2799 567
rect 2803 563 2804 567
rect 2798 562 2804 563
rect 2982 567 2988 568
rect 2982 563 2983 567
rect 2987 563 2988 567
rect 2982 562 2988 563
rect 3166 567 3172 568
rect 3166 563 3167 567
rect 3171 563 3172 567
rect 3166 562 3172 563
rect 3358 567 3364 568
rect 3358 563 3359 567
rect 3363 563 3364 567
rect 3462 564 3463 568
rect 3467 564 3468 568
rect 3462 563 3468 564
rect 3358 562 3364 563
rect 110 560 116 561
rect 1766 560 1772 561
rect 110 556 111 560
rect 115 556 116 560
rect 110 555 116 556
rect 598 559 604 560
rect 598 555 599 559
rect 603 555 604 559
rect 598 554 604 555
rect 702 559 708 560
rect 702 555 703 559
rect 707 555 708 559
rect 702 554 708 555
rect 814 559 820 560
rect 814 555 815 559
rect 819 555 820 559
rect 814 554 820 555
rect 926 559 932 560
rect 926 555 927 559
rect 931 555 932 559
rect 926 554 932 555
rect 1038 559 1044 560
rect 1038 555 1039 559
rect 1043 555 1044 559
rect 1038 554 1044 555
rect 1150 559 1156 560
rect 1150 555 1151 559
rect 1155 555 1156 559
rect 1150 554 1156 555
rect 1254 559 1260 560
rect 1254 555 1255 559
rect 1259 555 1260 559
rect 1254 554 1260 555
rect 1358 559 1364 560
rect 1358 555 1359 559
rect 1363 555 1364 559
rect 1358 554 1364 555
rect 1470 559 1476 560
rect 1470 555 1471 559
rect 1475 555 1476 559
rect 1470 554 1476 555
rect 1582 559 1588 560
rect 1582 555 1583 559
rect 1587 555 1588 559
rect 1582 554 1588 555
rect 1670 559 1676 560
rect 1670 555 1671 559
rect 1675 555 1676 559
rect 1766 556 1767 560
rect 1771 556 1772 560
rect 1766 555 1772 556
rect 1670 554 1676 555
rect 1806 551 1812 552
rect 1806 547 1807 551
rect 1811 547 1812 551
rect 3462 551 3468 552
rect 1806 546 1812 547
rect 1830 548 1836 549
rect 1830 544 1831 548
rect 1835 544 1836 548
rect 110 543 116 544
rect 110 539 111 543
rect 115 539 116 543
rect 1766 543 1772 544
rect 1830 543 1836 544
rect 1966 548 1972 549
rect 1966 544 1967 548
rect 1971 544 1972 548
rect 1966 543 1972 544
rect 2126 548 2132 549
rect 2126 544 2127 548
rect 2131 544 2132 548
rect 2126 543 2132 544
rect 2286 548 2292 549
rect 2286 544 2287 548
rect 2291 544 2292 548
rect 2286 543 2292 544
rect 2454 548 2460 549
rect 2454 544 2455 548
rect 2459 544 2460 548
rect 2454 543 2460 544
rect 2622 548 2628 549
rect 2622 544 2623 548
rect 2627 544 2628 548
rect 2622 543 2628 544
rect 2798 548 2804 549
rect 2798 544 2799 548
rect 2803 544 2804 548
rect 2798 543 2804 544
rect 2982 548 2988 549
rect 2982 544 2983 548
rect 2987 544 2988 548
rect 2982 543 2988 544
rect 3166 548 3172 549
rect 3166 544 3167 548
rect 3171 544 3172 548
rect 3166 543 3172 544
rect 3358 548 3364 549
rect 3358 544 3359 548
rect 3363 544 3364 548
rect 3462 547 3463 551
rect 3467 547 3468 551
rect 3462 546 3468 547
rect 3358 543 3364 544
rect 110 538 116 539
rect 598 540 604 541
rect 598 536 599 540
rect 603 536 604 540
rect 598 535 604 536
rect 702 540 708 541
rect 702 536 703 540
rect 707 536 708 540
rect 702 535 708 536
rect 814 540 820 541
rect 814 536 815 540
rect 819 536 820 540
rect 814 535 820 536
rect 926 540 932 541
rect 926 536 927 540
rect 931 536 932 540
rect 926 535 932 536
rect 1038 540 1044 541
rect 1038 536 1039 540
rect 1043 536 1044 540
rect 1038 535 1044 536
rect 1150 540 1156 541
rect 1150 536 1151 540
rect 1155 536 1156 540
rect 1150 535 1156 536
rect 1254 540 1260 541
rect 1254 536 1255 540
rect 1259 536 1260 540
rect 1254 535 1260 536
rect 1358 540 1364 541
rect 1358 536 1359 540
rect 1363 536 1364 540
rect 1358 535 1364 536
rect 1470 540 1476 541
rect 1470 536 1471 540
rect 1475 536 1476 540
rect 1470 535 1476 536
rect 1582 540 1588 541
rect 1582 536 1583 540
rect 1587 536 1588 540
rect 1582 535 1588 536
rect 1670 540 1676 541
rect 1670 536 1671 540
rect 1675 536 1676 540
rect 1766 539 1767 543
rect 1771 539 1772 543
rect 1766 538 1772 539
rect 1670 535 1676 536
rect 302 496 308 497
rect 110 493 116 494
rect 110 489 111 493
rect 115 489 116 493
rect 302 492 303 496
rect 307 492 308 496
rect 302 491 308 492
rect 430 496 436 497
rect 430 492 431 496
rect 435 492 436 496
rect 430 491 436 492
rect 566 496 572 497
rect 566 492 567 496
rect 571 492 572 496
rect 566 491 572 492
rect 702 496 708 497
rect 702 492 703 496
rect 707 492 708 496
rect 702 491 708 492
rect 846 496 852 497
rect 846 492 847 496
rect 851 492 852 496
rect 846 491 852 492
rect 982 496 988 497
rect 982 492 983 496
rect 987 492 988 496
rect 982 491 988 492
rect 1110 496 1116 497
rect 1110 492 1111 496
rect 1115 492 1116 496
rect 1110 491 1116 492
rect 1230 496 1236 497
rect 1230 492 1231 496
rect 1235 492 1236 496
rect 1230 491 1236 492
rect 1350 496 1356 497
rect 1350 492 1351 496
rect 1355 492 1356 496
rect 1350 491 1356 492
rect 1462 496 1468 497
rect 1462 492 1463 496
rect 1467 492 1468 496
rect 1462 491 1468 492
rect 1574 496 1580 497
rect 1574 492 1575 496
rect 1579 492 1580 496
rect 1574 491 1580 492
rect 1670 496 1676 497
rect 1670 492 1671 496
rect 1675 492 1676 496
rect 1670 491 1676 492
rect 1766 493 1772 494
rect 110 488 116 489
rect 1766 489 1767 493
rect 1771 489 1772 493
rect 1766 488 1772 489
rect 1830 488 1836 489
rect 1806 485 1812 486
rect 1806 481 1807 485
rect 1811 481 1812 485
rect 1830 484 1831 488
rect 1835 484 1836 488
rect 1830 483 1836 484
rect 1966 488 1972 489
rect 1966 484 1967 488
rect 1971 484 1972 488
rect 1966 483 1972 484
rect 2126 488 2132 489
rect 2126 484 2127 488
rect 2131 484 2132 488
rect 2126 483 2132 484
rect 2294 488 2300 489
rect 2294 484 2295 488
rect 2299 484 2300 488
rect 2294 483 2300 484
rect 2478 488 2484 489
rect 2478 484 2479 488
rect 2483 484 2484 488
rect 2478 483 2484 484
rect 2678 488 2684 489
rect 2678 484 2679 488
rect 2683 484 2684 488
rect 2678 483 2684 484
rect 2886 488 2892 489
rect 2886 484 2887 488
rect 2891 484 2892 488
rect 2886 483 2892 484
rect 3110 488 3116 489
rect 3110 484 3111 488
rect 3115 484 3116 488
rect 3110 483 3116 484
rect 3334 488 3340 489
rect 3334 484 3335 488
rect 3339 484 3340 488
rect 3334 483 3340 484
rect 3462 485 3468 486
rect 1806 480 1812 481
rect 3462 481 3463 485
rect 3467 481 3468 485
rect 3462 480 3468 481
rect 302 477 308 478
rect 110 476 116 477
rect 110 472 111 476
rect 115 472 116 476
rect 302 473 303 477
rect 307 473 308 477
rect 302 472 308 473
rect 430 477 436 478
rect 430 473 431 477
rect 435 473 436 477
rect 430 472 436 473
rect 566 477 572 478
rect 566 473 567 477
rect 571 473 572 477
rect 566 472 572 473
rect 702 477 708 478
rect 702 473 703 477
rect 707 473 708 477
rect 702 472 708 473
rect 846 477 852 478
rect 846 473 847 477
rect 851 473 852 477
rect 846 472 852 473
rect 982 477 988 478
rect 982 473 983 477
rect 987 473 988 477
rect 982 472 988 473
rect 1110 477 1116 478
rect 1110 473 1111 477
rect 1115 473 1116 477
rect 1110 472 1116 473
rect 1230 477 1236 478
rect 1230 473 1231 477
rect 1235 473 1236 477
rect 1230 472 1236 473
rect 1350 477 1356 478
rect 1350 473 1351 477
rect 1355 473 1356 477
rect 1350 472 1356 473
rect 1462 477 1468 478
rect 1462 473 1463 477
rect 1467 473 1468 477
rect 1462 472 1468 473
rect 1574 477 1580 478
rect 1574 473 1575 477
rect 1579 473 1580 477
rect 1574 472 1580 473
rect 1670 477 1676 478
rect 1670 473 1671 477
rect 1675 473 1676 477
rect 1670 472 1676 473
rect 1766 476 1772 477
rect 1766 472 1767 476
rect 1771 472 1772 476
rect 110 471 116 472
rect 1766 471 1772 472
rect 1830 469 1836 470
rect 1806 468 1812 469
rect 1806 464 1807 468
rect 1811 464 1812 468
rect 1830 465 1831 469
rect 1835 465 1836 469
rect 1830 464 1836 465
rect 1966 469 1972 470
rect 1966 465 1967 469
rect 1971 465 1972 469
rect 1966 464 1972 465
rect 2126 469 2132 470
rect 2126 465 2127 469
rect 2131 465 2132 469
rect 2126 464 2132 465
rect 2294 469 2300 470
rect 2294 465 2295 469
rect 2299 465 2300 469
rect 2294 464 2300 465
rect 2478 469 2484 470
rect 2478 465 2479 469
rect 2483 465 2484 469
rect 2478 464 2484 465
rect 2678 469 2684 470
rect 2678 465 2679 469
rect 2683 465 2684 469
rect 2678 464 2684 465
rect 2886 469 2892 470
rect 2886 465 2887 469
rect 2891 465 2892 469
rect 2886 464 2892 465
rect 3110 469 3116 470
rect 3110 465 3111 469
rect 3115 465 3116 469
rect 3110 464 3116 465
rect 3334 469 3340 470
rect 3334 465 3335 469
rect 3339 465 3340 469
rect 3334 464 3340 465
rect 3462 468 3468 469
rect 3462 464 3463 468
rect 3467 464 3468 468
rect 1806 463 1812 464
rect 3462 463 3468 464
rect 110 424 116 425
rect 1766 424 1772 425
rect 110 420 111 424
rect 115 420 116 424
rect 110 419 116 420
rect 134 423 140 424
rect 134 419 135 423
rect 139 419 140 423
rect 134 418 140 419
rect 254 423 260 424
rect 254 419 255 423
rect 259 419 260 423
rect 254 418 260 419
rect 414 423 420 424
rect 414 419 415 423
rect 419 419 420 423
rect 414 418 420 419
rect 582 423 588 424
rect 582 419 583 423
rect 587 419 588 423
rect 582 418 588 419
rect 742 423 748 424
rect 742 419 743 423
rect 747 419 748 423
rect 742 418 748 419
rect 902 423 908 424
rect 902 419 903 423
rect 907 419 908 423
rect 902 418 908 419
rect 1046 423 1052 424
rect 1046 419 1047 423
rect 1051 419 1052 423
rect 1046 418 1052 419
rect 1182 423 1188 424
rect 1182 419 1183 423
rect 1187 419 1188 423
rect 1182 418 1188 419
rect 1310 423 1316 424
rect 1310 419 1311 423
rect 1315 419 1316 423
rect 1310 418 1316 419
rect 1438 423 1444 424
rect 1438 419 1439 423
rect 1443 419 1444 423
rect 1438 418 1444 419
rect 1566 423 1572 424
rect 1566 419 1567 423
rect 1571 419 1572 423
rect 1566 418 1572 419
rect 1670 423 1676 424
rect 1670 419 1671 423
rect 1675 419 1676 423
rect 1766 420 1767 424
rect 1771 420 1772 424
rect 1766 419 1772 420
rect 1806 424 1812 425
rect 3462 424 3468 425
rect 1806 420 1807 424
rect 1811 420 1812 424
rect 1806 419 1812 420
rect 1830 423 1836 424
rect 1830 419 1831 423
rect 1835 419 1836 423
rect 1670 418 1676 419
rect 1830 418 1836 419
rect 1958 423 1964 424
rect 1958 419 1959 423
rect 1963 419 1964 423
rect 1958 418 1964 419
rect 2110 423 2116 424
rect 2110 419 2111 423
rect 2115 419 2116 423
rect 2110 418 2116 419
rect 2270 423 2276 424
rect 2270 419 2271 423
rect 2275 419 2276 423
rect 2270 418 2276 419
rect 2454 423 2460 424
rect 2454 419 2455 423
rect 2459 419 2460 423
rect 2454 418 2460 419
rect 2654 423 2660 424
rect 2654 419 2655 423
rect 2659 419 2660 423
rect 2654 418 2660 419
rect 2870 423 2876 424
rect 2870 419 2871 423
rect 2875 419 2876 423
rect 2870 418 2876 419
rect 3102 423 3108 424
rect 3102 419 3103 423
rect 3107 419 3108 423
rect 3102 418 3108 419
rect 3334 423 3340 424
rect 3334 419 3335 423
rect 3339 419 3340 423
rect 3462 420 3463 424
rect 3467 420 3468 424
rect 3462 419 3468 420
rect 3334 418 3340 419
rect 110 407 116 408
rect 110 403 111 407
rect 115 403 116 407
rect 1766 407 1772 408
rect 110 402 116 403
rect 134 404 140 405
rect 134 400 135 404
rect 139 400 140 404
rect 134 399 140 400
rect 254 404 260 405
rect 254 400 255 404
rect 259 400 260 404
rect 254 399 260 400
rect 414 404 420 405
rect 414 400 415 404
rect 419 400 420 404
rect 414 399 420 400
rect 582 404 588 405
rect 582 400 583 404
rect 587 400 588 404
rect 582 399 588 400
rect 742 404 748 405
rect 742 400 743 404
rect 747 400 748 404
rect 742 399 748 400
rect 902 404 908 405
rect 902 400 903 404
rect 907 400 908 404
rect 902 399 908 400
rect 1046 404 1052 405
rect 1046 400 1047 404
rect 1051 400 1052 404
rect 1046 399 1052 400
rect 1182 404 1188 405
rect 1182 400 1183 404
rect 1187 400 1188 404
rect 1182 399 1188 400
rect 1310 404 1316 405
rect 1310 400 1311 404
rect 1315 400 1316 404
rect 1310 399 1316 400
rect 1438 404 1444 405
rect 1438 400 1439 404
rect 1443 400 1444 404
rect 1438 399 1444 400
rect 1566 404 1572 405
rect 1566 400 1567 404
rect 1571 400 1572 404
rect 1566 399 1572 400
rect 1670 404 1676 405
rect 1670 400 1671 404
rect 1675 400 1676 404
rect 1766 403 1767 407
rect 1771 403 1772 407
rect 1766 402 1772 403
rect 1806 407 1812 408
rect 1806 403 1807 407
rect 1811 403 1812 407
rect 3462 407 3468 408
rect 1806 402 1812 403
rect 1830 404 1836 405
rect 1670 399 1676 400
rect 1830 400 1831 404
rect 1835 400 1836 404
rect 1830 399 1836 400
rect 1958 404 1964 405
rect 1958 400 1959 404
rect 1963 400 1964 404
rect 1958 399 1964 400
rect 2110 404 2116 405
rect 2110 400 2111 404
rect 2115 400 2116 404
rect 2110 399 2116 400
rect 2270 404 2276 405
rect 2270 400 2271 404
rect 2275 400 2276 404
rect 2270 399 2276 400
rect 2454 404 2460 405
rect 2454 400 2455 404
rect 2459 400 2460 404
rect 2454 399 2460 400
rect 2654 404 2660 405
rect 2654 400 2655 404
rect 2659 400 2660 404
rect 2654 399 2660 400
rect 2870 404 2876 405
rect 2870 400 2871 404
rect 2875 400 2876 404
rect 2870 399 2876 400
rect 3102 404 3108 405
rect 3102 400 3103 404
rect 3107 400 3108 404
rect 3102 399 3108 400
rect 3334 404 3340 405
rect 3334 400 3335 404
rect 3339 400 3340 404
rect 3462 403 3463 407
rect 3467 403 3468 407
rect 3462 402 3468 403
rect 3334 399 3340 400
rect 134 356 140 357
rect 110 353 116 354
rect 110 349 111 353
rect 115 349 116 353
rect 134 352 135 356
rect 139 352 140 356
rect 134 351 140 352
rect 222 356 228 357
rect 222 352 223 356
rect 227 352 228 356
rect 222 351 228 352
rect 342 356 348 357
rect 342 352 343 356
rect 347 352 348 356
rect 342 351 348 352
rect 470 356 476 357
rect 470 352 471 356
rect 475 352 476 356
rect 470 351 476 352
rect 598 356 604 357
rect 598 352 599 356
rect 603 352 604 356
rect 598 351 604 352
rect 718 356 724 357
rect 718 352 719 356
rect 723 352 724 356
rect 718 351 724 352
rect 838 356 844 357
rect 838 352 839 356
rect 843 352 844 356
rect 838 351 844 352
rect 958 356 964 357
rect 958 352 959 356
rect 963 352 964 356
rect 958 351 964 352
rect 1078 356 1084 357
rect 1078 352 1079 356
rect 1083 352 1084 356
rect 1078 351 1084 352
rect 1206 356 1212 357
rect 1206 352 1207 356
rect 1211 352 1212 356
rect 1926 356 1932 357
rect 1206 351 1212 352
rect 1766 353 1772 354
rect 110 348 116 349
rect 1766 349 1767 353
rect 1771 349 1772 353
rect 1766 348 1772 349
rect 1806 353 1812 354
rect 1806 349 1807 353
rect 1811 349 1812 353
rect 1926 352 1927 356
rect 1931 352 1932 356
rect 1926 351 1932 352
rect 2038 356 2044 357
rect 2038 352 2039 356
rect 2043 352 2044 356
rect 2038 351 2044 352
rect 2158 356 2164 357
rect 2158 352 2159 356
rect 2163 352 2164 356
rect 2158 351 2164 352
rect 2286 356 2292 357
rect 2286 352 2287 356
rect 2291 352 2292 356
rect 2286 351 2292 352
rect 2422 356 2428 357
rect 2422 352 2423 356
rect 2427 352 2428 356
rect 2422 351 2428 352
rect 2582 356 2588 357
rect 2582 352 2583 356
rect 2587 352 2588 356
rect 2582 351 2588 352
rect 2758 356 2764 357
rect 2758 352 2759 356
rect 2763 352 2764 356
rect 2758 351 2764 352
rect 2950 356 2956 357
rect 2950 352 2951 356
rect 2955 352 2956 356
rect 2950 351 2956 352
rect 3150 356 3156 357
rect 3150 352 3151 356
rect 3155 352 3156 356
rect 3150 351 3156 352
rect 3358 356 3364 357
rect 3358 352 3359 356
rect 3363 352 3364 356
rect 3358 351 3364 352
rect 3462 353 3468 354
rect 1806 348 1812 349
rect 3462 349 3463 353
rect 3467 349 3468 353
rect 3462 348 3468 349
rect 134 337 140 338
rect 110 336 116 337
rect 110 332 111 336
rect 115 332 116 336
rect 134 333 135 337
rect 139 333 140 337
rect 134 332 140 333
rect 222 337 228 338
rect 222 333 223 337
rect 227 333 228 337
rect 222 332 228 333
rect 342 337 348 338
rect 342 333 343 337
rect 347 333 348 337
rect 342 332 348 333
rect 470 337 476 338
rect 470 333 471 337
rect 475 333 476 337
rect 470 332 476 333
rect 598 337 604 338
rect 598 333 599 337
rect 603 333 604 337
rect 598 332 604 333
rect 718 337 724 338
rect 718 333 719 337
rect 723 333 724 337
rect 718 332 724 333
rect 838 337 844 338
rect 838 333 839 337
rect 843 333 844 337
rect 838 332 844 333
rect 958 337 964 338
rect 958 333 959 337
rect 963 333 964 337
rect 958 332 964 333
rect 1078 337 1084 338
rect 1078 333 1079 337
rect 1083 333 1084 337
rect 1078 332 1084 333
rect 1206 337 1212 338
rect 1926 337 1932 338
rect 1206 333 1207 337
rect 1211 333 1212 337
rect 1206 332 1212 333
rect 1766 336 1772 337
rect 1766 332 1767 336
rect 1771 332 1772 336
rect 110 331 116 332
rect 1766 331 1772 332
rect 1806 336 1812 337
rect 1806 332 1807 336
rect 1811 332 1812 336
rect 1926 333 1927 337
rect 1931 333 1932 337
rect 1926 332 1932 333
rect 2038 337 2044 338
rect 2038 333 2039 337
rect 2043 333 2044 337
rect 2038 332 2044 333
rect 2158 337 2164 338
rect 2158 333 2159 337
rect 2163 333 2164 337
rect 2158 332 2164 333
rect 2286 337 2292 338
rect 2286 333 2287 337
rect 2291 333 2292 337
rect 2286 332 2292 333
rect 2422 337 2428 338
rect 2422 333 2423 337
rect 2427 333 2428 337
rect 2422 332 2428 333
rect 2582 337 2588 338
rect 2582 333 2583 337
rect 2587 333 2588 337
rect 2582 332 2588 333
rect 2758 337 2764 338
rect 2758 333 2759 337
rect 2763 333 2764 337
rect 2758 332 2764 333
rect 2950 337 2956 338
rect 2950 333 2951 337
rect 2955 333 2956 337
rect 2950 332 2956 333
rect 3150 337 3156 338
rect 3150 333 3151 337
rect 3155 333 3156 337
rect 3150 332 3156 333
rect 3358 337 3364 338
rect 3358 333 3359 337
rect 3363 333 3364 337
rect 3358 332 3364 333
rect 3462 336 3468 337
rect 3462 332 3463 336
rect 3467 332 3468 336
rect 1806 331 1812 332
rect 3462 331 3468 332
rect 1806 292 1812 293
rect 3462 292 3468 293
rect 110 288 116 289
rect 1766 288 1772 289
rect 110 284 111 288
rect 115 284 116 288
rect 110 283 116 284
rect 262 287 268 288
rect 262 283 263 287
rect 267 283 268 287
rect 262 282 268 283
rect 374 287 380 288
rect 374 283 375 287
rect 379 283 380 287
rect 374 282 380 283
rect 486 287 492 288
rect 486 283 487 287
rect 491 283 492 287
rect 486 282 492 283
rect 598 287 604 288
rect 598 283 599 287
rect 603 283 604 287
rect 598 282 604 283
rect 710 287 716 288
rect 710 283 711 287
rect 715 283 716 287
rect 710 282 716 283
rect 814 287 820 288
rect 814 283 815 287
rect 819 283 820 287
rect 814 282 820 283
rect 918 287 924 288
rect 918 283 919 287
rect 923 283 924 287
rect 918 282 924 283
rect 1022 287 1028 288
rect 1022 283 1023 287
rect 1027 283 1028 287
rect 1022 282 1028 283
rect 1126 287 1132 288
rect 1126 283 1127 287
rect 1131 283 1132 287
rect 1126 282 1132 283
rect 1238 287 1244 288
rect 1238 283 1239 287
rect 1243 283 1244 287
rect 1766 284 1767 288
rect 1771 284 1772 288
rect 1806 288 1807 292
rect 1811 288 1812 292
rect 1806 287 1812 288
rect 2222 291 2228 292
rect 2222 287 2223 291
rect 2227 287 2228 291
rect 2222 286 2228 287
rect 2310 291 2316 292
rect 2310 287 2311 291
rect 2315 287 2316 291
rect 2310 286 2316 287
rect 2398 291 2404 292
rect 2398 287 2399 291
rect 2403 287 2404 291
rect 2398 286 2404 287
rect 2486 291 2492 292
rect 2486 287 2487 291
rect 2491 287 2492 291
rect 2486 286 2492 287
rect 2574 291 2580 292
rect 2574 287 2575 291
rect 2579 287 2580 291
rect 2574 286 2580 287
rect 2678 291 2684 292
rect 2678 287 2679 291
rect 2683 287 2684 291
rect 2678 286 2684 287
rect 2798 291 2804 292
rect 2798 287 2799 291
rect 2803 287 2804 291
rect 2798 286 2804 287
rect 2926 291 2932 292
rect 2926 287 2927 291
rect 2931 287 2932 291
rect 2926 286 2932 287
rect 3070 291 3076 292
rect 3070 287 3071 291
rect 3075 287 3076 291
rect 3070 286 3076 287
rect 3222 291 3228 292
rect 3222 287 3223 291
rect 3227 287 3228 291
rect 3222 286 3228 287
rect 3366 291 3372 292
rect 3366 287 3367 291
rect 3371 287 3372 291
rect 3462 288 3463 292
rect 3467 288 3468 292
rect 3462 287 3468 288
rect 3366 286 3372 287
rect 1766 283 1772 284
rect 1238 282 1244 283
rect 1806 275 1812 276
rect 110 271 116 272
rect 110 267 111 271
rect 115 267 116 271
rect 1766 271 1772 272
rect 110 266 116 267
rect 262 268 268 269
rect 262 264 263 268
rect 267 264 268 268
rect 262 263 268 264
rect 374 268 380 269
rect 374 264 375 268
rect 379 264 380 268
rect 374 263 380 264
rect 486 268 492 269
rect 486 264 487 268
rect 491 264 492 268
rect 486 263 492 264
rect 598 268 604 269
rect 598 264 599 268
rect 603 264 604 268
rect 598 263 604 264
rect 710 268 716 269
rect 710 264 711 268
rect 715 264 716 268
rect 710 263 716 264
rect 814 268 820 269
rect 814 264 815 268
rect 819 264 820 268
rect 814 263 820 264
rect 918 268 924 269
rect 918 264 919 268
rect 923 264 924 268
rect 918 263 924 264
rect 1022 268 1028 269
rect 1022 264 1023 268
rect 1027 264 1028 268
rect 1022 263 1028 264
rect 1126 268 1132 269
rect 1126 264 1127 268
rect 1131 264 1132 268
rect 1126 263 1132 264
rect 1238 268 1244 269
rect 1238 264 1239 268
rect 1243 264 1244 268
rect 1766 267 1767 271
rect 1771 267 1772 271
rect 1806 271 1807 275
rect 1811 271 1812 275
rect 3462 275 3468 276
rect 1806 270 1812 271
rect 2222 272 2228 273
rect 2222 268 2223 272
rect 2227 268 2228 272
rect 2222 267 2228 268
rect 2310 272 2316 273
rect 2310 268 2311 272
rect 2315 268 2316 272
rect 2310 267 2316 268
rect 2398 272 2404 273
rect 2398 268 2399 272
rect 2403 268 2404 272
rect 2398 267 2404 268
rect 2486 272 2492 273
rect 2486 268 2487 272
rect 2491 268 2492 272
rect 2486 267 2492 268
rect 2574 272 2580 273
rect 2574 268 2575 272
rect 2579 268 2580 272
rect 2574 267 2580 268
rect 2678 272 2684 273
rect 2678 268 2679 272
rect 2683 268 2684 272
rect 2678 267 2684 268
rect 2798 272 2804 273
rect 2798 268 2799 272
rect 2803 268 2804 272
rect 2798 267 2804 268
rect 2926 272 2932 273
rect 2926 268 2927 272
rect 2931 268 2932 272
rect 2926 267 2932 268
rect 3070 272 3076 273
rect 3070 268 3071 272
rect 3075 268 3076 272
rect 3070 267 3076 268
rect 3222 272 3228 273
rect 3222 268 3223 272
rect 3227 268 3228 272
rect 3222 267 3228 268
rect 3366 272 3372 273
rect 3366 268 3367 272
rect 3371 268 3372 272
rect 3462 271 3463 275
rect 3467 271 3468 275
rect 3462 270 3468 271
rect 3366 267 3372 268
rect 1766 266 1772 267
rect 1238 263 1244 264
rect 446 220 452 221
rect 110 217 116 218
rect 110 213 111 217
rect 115 213 116 217
rect 446 216 447 220
rect 451 216 452 220
rect 446 215 452 216
rect 534 220 540 221
rect 534 216 535 220
rect 539 216 540 220
rect 534 215 540 216
rect 622 220 628 221
rect 622 216 623 220
rect 627 216 628 220
rect 622 215 628 216
rect 710 220 716 221
rect 710 216 711 220
rect 715 216 716 220
rect 710 215 716 216
rect 806 220 812 221
rect 806 216 807 220
rect 811 216 812 220
rect 806 215 812 216
rect 902 220 908 221
rect 902 216 903 220
rect 907 216 908 220
rect 902 215 908 216
rect 998 220 1004 221
rect 998 216 999 220
rect 1003 216 1004 220
rect 998 215 1004 216
rect 1102 220 1108 221
rect 1102 216 1103 220
rect 1107 216 1108 220
rect 1102 215 1108 216
rect 1206 220 1212 221
rect 1206 216 1207 220
rect 1211 216 1212 220
rect 1206 215 1212 216
rect 1310 220 1316 221
rect 1310 216 1311 220
rect 1315 216 1316 220
rect 2142 220 2148 221
rect 1310 215 1316 216
rect 1766 217 1772 218
rect 110 212 116 213
rect 1766 213 1767 217
rect 1771 213 1772 217
rect 1766 212 1772 213
rect 1806 217 1812 218
rect 1806 213 1807 217
rect 1811 213 1812 217
rect 2142 216 2143 220
rect 2147 216 2148 220
rect 2142 215 2148 216
rect 2262 220 2268 221
rect 2262 216 2263 220
rect 2267 216 2268 220
rect 2262 215 2268 216
rect 2382 220 2388 221
rect 2382 216 2383 220
rect 2387 216 2388 220
rect 2382 215 2388 216
rect 2510 220 2516 221
rect 2510 216 2511 220
rect 2515 216 2516 220
rect 2510 215 2516 216
rect 2638 220 2644 221
rect 2638 216 2639 220
rect 2643 216 2644 220
rect 2638 215 2644 216
rect 2766 220 2772 221
rect 2766 216 2767 220
rect 2771 216 2772 220
rect 2766 215 2772 216
rect 2894 220 2900 221
rect 2894 216 2895 220
rect 2899 216 2900 220
rect 2894 215 2900 216
rect 3014 220 3020 221
rect 3014 216 3015 220
rect 3019 216 3020 220
rect 3014 215 3020 216
rect 3134 220 3140 221
rect 3134 216 3135 220
rect 3139 216 3140 220
rect 3134 215 3140 216
rect 3262 220 3268 221
rect 3262 216 3263 220
rect 3267 216 3268 220
rect 3262 215 3268 216
rect 3366 220 3372 221
rect 3366 216 3367 220
rect 3371 216 3372 220
rect 3366 215 3372 216
rect 3462 217 3468 218
rect 1806 212 1812 213
rect 3462 213 3463 217
rect 3467 213 3468 217
rect 3462 212 3468 213
rect 446 201 452 202
rect 110 200 116 201
rect 110 196 111 200
rect 115 196 116 200
rect 446 197 447 201
rect 451 197 452 201
rect 446 196 452 197
rect 534 201 540 202
rect 534 197 535 201
rect 539 197 540 201
rect 534 196 540 197
rect 622 201 628 202
rect 622 197 623 201
rect 627 197 628 201
rect 622 196 628 197
rect 710 201 716 202
rect 710 197 711 201
rect 715 197 716 201
rect 710 196 716 197
rect 806 201 812 202
rect 806 197 807 201
rect 811 197 812 201
rect 806 196 812 197
rect 902 201 908 202
rect 902 197 903 201
rect 907 197 908 201
rect 902 196 908 197
rect 998 201 1004 202
rect 998 197 999 201
rect 1003 197 1004 201
rect 998 196 1004 197
rect 1102 201 1108 202
rect 1102 197 1103 201
rect 1107 197 1108 201
rect 1102 196 1108 197
rect 1206 201 1212 202
rect 1206 197 1207 201
rect 1211 197 1212 201
rect 1206 196 1212 197
rect 1310 201 1316 202
rect 2142 201 2148 202
rect 1310 197 1311 201
rect 1315 197 1316 201
rect 1310 196 1316 197
rect 1766 200 1772 201
rect 1766 196 1767 200
rect 1771 196 1772 200
rect 110 195 116 196
rect 1766 195 1772 196
rect 1806 200 1812 201
rect 1806 196 1807 200
rect 1811 196 1812 200
rect 2142 197 2143 201
rect 2147 197 2148 201
rect 2142 196 2148 197
rect 2262 201 2268 202
rect 2262 197 2263 201
rect 2267 197 2268 201
rect 2262 196 2268 197
rect 2382 201 2388 202
rect 2382 197 2383 201
rect 2387 197 2388 201
rect 2382 196 2388 197
rect 2510 201 2516 202
rect 2510 197 2511 201
rect 2515 197 2516 201
rect 2510 196 2516 197
rect 2638 201 2644 202
rect 2638 197 2639 201
rect 2643 197 2644 201
rect 2638 196 2644 197
rect 2766 201 2772 202
rect 2766 197 2767 201
rect 2771 197 2772 201
rect 2766 196 2772 197
rect 2894 201 2900 202
rect 2894 197 2895 201
rect 2899 197 2900 201
rect 2894 196 2900 197
rect 3014 201 3020 202
rect 3014 197 3015 201
rect 3019 197 3020 201
rect 3014 196 3020 197
rect 3134 201 3140 202
rect 3134 197 3135 201
rect 3139 197 3140 201
rect 3134 196 3140 197
rect 3262 201 3268 202
rect 3262 197 3263 201
rect 3267 197 3268 201
rect 3262 196 3268 197
rect 3366 201 3372 202
rect 3366 197 3367 201
rect 3371 197 3372 201
rect 3366 196 3372 197
rect 3462 200 3468 201
rect 3462 196 3463 200
rect 3467 196 3468 200
rect 1806 195 1812 196
rect 3462 195 3468 196
rect 1806 132 1812 133
rect 3462 132 3468 133
rect 110 128 116 129
rect 1766 128 1772 129
rect 110 124 111 128
rect 115 124 116 128
rect 110 123 116 124
rect 262 127 268 128
rect 262 123 263 127
rect 267 123 268 127
rect 262 122 268 123
rect 350 127 356 128
rect 350 123 351 127
rect 355 123 356 127
rect 350 122 356 123
rect 438 127 444 128
rect 438 123 439 127
rect 443 123 444 127
rect 438 122 444 123
rect 526 127 532 128
rect 526 123 527 127
rect 531 123 532 127
rect 526 122 532 123
rect 614 127 620 128
rect 614 123 615 127
rect 619 123 620 127
rect 614 122 620 123
rect 702 127 708 128
rect 702 123 703 127
rect 707 123 708 127
rect 702 122 708 123
rect 790 127 796 128
rect 790 123 791 127
rect 795 123 796 127
rect 790 122 796 123
rect 878 127 884 128
rect 878 123 879 127
rect 883 123 884 127
rect 878 122 884 123
rect 966 127 972 128
rect 966 123 967 127
rect 971 123 972 127
rect 966 122 972 123
rect 1054 127 1060 128
rect 1054 123 1055 127
rect 1059 123 1060 127
rect 1054 122 1060 123
rect 1142 127 1148 128
rect 1142 123 1143 127
rect 1147 123 1148 127
rect 1142 122 1148 123
rect 1230 127 1236 128
rect 1230 123 1231 127
rect 1235 123 1236 127
rect 1230 122 1236 123
rect 1318 127 1324 128
rect 1318 123 1319 127
rect 1323 123 1324 127
rect 1318 122 1324 123
rect 1406 127 1412 128
rect 1406 123 1407 127
rect 1411 123 1412 127
rect 1406 122 1412 123
rect 1494 127 1500 128
rect 1494 123 1495 127
rect 1499 123 1500 127
rect 1494 122 1500 123
rect 1582 127 1588 128
rect 1582 123 1583 127
rect 1587 123 1588 127
rect 1582 122 1588 123
rect 1670 127 1676 128
rect 1670 123 1671 127
rect 1675 123 1676 127
rect 1766 124 1767 128
rect 1771 124 1772 128
rect 1806 128 1807 132
rect 1811 128 1812 132
rect 1806 127 1812 128
rect 1830 131 1836 132
rect 1830 127 1831 131
rect 1835 127 1836 131
rect 1830 126 1836 127
rect 1918 131 1924 132
rect 1918 127 1919 131
rect 1923 127 1924 131
rect 1918 126 1924 127
rect 2006 131 2012 132
rect 2006 127 2007 131
rect 2011 127 2012 131
rect 2006 126 2012 127
rect 2094 131 2100 132
rect 2094 127 2095 131
rect 2099 127 2100 131
rect 2094 126 2100 127
rect 2182 131 2188 132
rect 2182 127 2183 131
rect 2187 127 2188 131
rect 2182 126 2188 127
rect 2294 131 2300 132
rect 2294 127 2295 131
rect 2299 127 2300 131
rect 2294 126 2300 127
rect 2406 131 2412 132
rect 2406 127 2407 131
rect 2411 127 2412 131
rect 2406 126 2412 127
rect 2510 131 2516 132
rect 2510 127 2511 131
rect 2515 127 2516 131
rect 2510 126 2516 127
rect 2614 131 2620 132
rect 2614 127 2615 131
rect 2619 127 2620 131
rect 2614 126 2620 127
rect 2718 131 2724 132
rect 2718 127 2719 131
rect 2723 127 2724 131
rect 2718 126 2724 127
rect 2814 131 2820 132
rect 2814 127 2815 131
rect 2819 127 2820 131
rect 2814 126 2820 127
rect 2910 131 2916 132
rect 2910 127 2911 131
rect 2915 127 2916 131
rect 2910 126 2916 127
rect 3006 131 3012 132
rect 3006 127 3007 131
rect 3011 127 3012 131
rect 3006 126 3012 127
rect 3102 131 3108 132
rect 3102 127 3103 131
rect 3107 127 3108 131
rect 3102 126 3108 127
rect 3190 131 3196 132
rect 3190 127 3191 131
rect 3195 127 3196 131
rect 3190 126 3196 127
rect 3278 131 3284 132
rect 3278 127 3279 131
rect 3283 127 3284 131
rect 3278 126 3284 127
rect 3366 131 3372 132
rect 3366 127 3367 131
rect 3371 127 3372 131
rect 3462 128 3463 132
rect 3467 128 3468 132
rect 3462 127 3468 128
rect 3366 126 3372 127
rect 1766 123 1772 124
rect 1670 122 1676 123
rect 1806 115 1812 116
rect 110 111 116 112
rect 110 107 111 111
rect 115 107 116 111
rect 1766 111 1772 112
rect 110 106 116 107
rect 262 108 268 109
rect 262 104 263 108
rect 267 104 268 108
rect 262 103 268 104
rect 350 108 356 109
rect 350 104 351 108
rect 355 104 356 108
rect 350 103 356 104
rect 438 108 444 109
rect 438 104 439 108
rect 443 104 444 108
rect 438 103 444 104
rect 526 108 532 109
rect 526 104 527 108
rect 531 104 532 108
rect 526 103 532 104
rect 614 108 620 109
rect 614 104 615 108
rect 619 104 620 108
rect 614 103 620 104
rect 702 108 708 109
rect 702 104 703 108
rect 707 104 708 108
rect 702 103 708 104
rect 790 108 796 109
rect 790 104 791 108
rect 795 104 796 108
rect 790 103 796 104
rect 878 108 884 109
rect 878 104 879 108
rect 883 104 884 108
rect 878 103 884 104
rect 966 108 972 109
rect 966 104 967 108
rect 971 104 972 108
rect 966 103 972 104
rect 1054 108 1060 109
rect 1054 104 1055 108
rect 1059 104 1060 108
rect 1054 103 1060 104
rect 1142 108 1148 109
rect 1142 104 1143 108
rect 1147 104 1148 108
rect 1142 103 1148 104
rect 1230 108 1236 109
rect 1230 104 1231 108
rect 1235 104 1236 108
rect 1230 103 1236 104
rect 1318 108 1324 109
rect 1318 104 1319 108
rect 1323 104 1324 108
rect 1318 103 1324 104
rect 1406 108 1412 109
rect 1406 104 1407 108
rect 1411 104 1412 108
rect 1406 103 1412 104
rect 1494 108 1500 109
rect 1494 104 1495 108
rect 1499 104 1500 108
rect 1494 103 1500 104
rect 1582 108 1588 109
rect 1582 104 1583 108
rect 1587 104 1588 108
rect 1582 103 1588 104
rect 1670 108 1676 109
rect 1670 104 1671 108
rect 1675 104 1676 108
rect 1766 107 1767 111
rect 1771 107 1772 111
rect 1806 111 1807 115
rect 1811 111 1812 115
rect 3462 115 3468 116
rect 1806 110 1812 111
rect 1830 112 1836 113
rect 1830 108 1831 112
rect 1835 108 1836 112
rect 1830 107 1836 108
rect 1918 112 1924 113
rect 1918 108 1919 112
rect 1923 108 1924 112
rect 1918 107 1924 108
rect 2006 112 2012 113
rect 2006 108 2007 112
rect 2011 108 2012 112
rect 2006 107 2012 108
rect 2094 112 2100 113
rect 2094 108 2095 112
rect 2099 108 2100 112
rect 2094 107 2100 108
rect 2182 112 2188 113
rect 2182 108 2183 112
rect 2187 108 2188 112
rect 2182 107 2188 108
rect 2294 112 2300 113
rect 2294 108 2295 112
rect 2299 108 2300 112
rect 2294 107 2300 108
rect 2406 112 2412 113
rect 2406 108 2407 112
rect 2411 108 2412 112
rect 2406 107 2412 108
rect 2510 112 2516 113
rect 2510 108 2511 112
rect 2515 108 2516 112
rect 2510 107 2516 108
rect 2614 112 2620 113
rect 2614 108 2615 112
rect 2619 108 2620 112
rect 2614 107 2620 108
rect 2718 112 2724 113
rect 2718 108 2719 112
rect 2723 108 2724 112
rect 2718 107 2724 108
rect 2814 112 2820 113
rect 2814 108 2815 112
rect 2819 108 2820 112
rect 2814 107 2820 108
rect 2910 112 2916 113
rect 2910 108 2911 112
rect 2915 108 2916 112
rect 2910 107 2916 108
rect 3006 112 3012 113
rect 3006 108 3007 112
rect 3011 108 3012 112
rect 3006 107 3012 108
rect 3102 112 3108 113
rect 3102 108 3103 112
rect 3107 108 3108 112
rect 3102 107 3108 108
rect 3190 112 3196 113
rect 3190 108 3191 112
rect 3195 108 3196 112
rect 3190 107 3196 108
rect 3278 112 3284 113
rect 3278 108 3279 112
rect 3283 108 3284 112
rect 3278 107 3284 108
rect 3366 112 3372 113
rect 3366 108 3367 112
rect 3371 108 3372 112
rect 3462 111 3463 115
rect 3467 111 3468 115
rect 3462 110 3468 111
rect 3366 107 3372 108
rect 1766 106 1772 107
rect 1670 103 1676 104
<< m3c >>
rect 111 3480 115 3484
rect 135 3479 139 3483
rect 271 3479 275 3483
rect 439 3479 443 3483
rect 615 3479 619 3483
rect 791 3479 795 3483
rect 959 3479 963 3483
rect 1119 3479 1123 3483
rect 1263 3479 1267 3483
rect 1407 3479 1411 3483
rect 1551 3479 1555 3483
rect 1671 3479 1675 3483
rect 1767 3480 1771 3484
rect 1807 3468 1811 3472
rect 111 3463 115 3467
rect 1831 3467 1835 3471
rect 135 3460 139 3464
rect 271 3460 275 3464
rect 439 3460 443 3464
rect 615 3460 619 3464
rect 791 3460 795 3464
rect 959 3460 963 3464
rect 1119 3460 1123 3464
rect 1263 3460 1267 3464
rect 1407 3460 1411 3464
rect 1551 3460 1555 3464
rect 1671 3460 1675 3464
rect 1767 3463 1771 3467
rect 1975 3467 1979 3471
rect 2143 3467 2147 3471
rect 2311 3467 2315 3471
rect 2479 3467 2483 3471
rect 2639 3467 2643 3471
rect 2799 3467 2803 3471
rect 2967 3467 2971 3471
rect 3463 3468 3467 3472
rect 1807 3451 1811 3455
rect 1831 3448 1835 3452
rect 1975 3448 1979 3452
rect 2143 3448 2147 3452
rect 2311 3448 2315 3452
rect 2479 3448 2483 3452
rect 2639 3448 2643 3452
rect 2799 3448 2803 3452
rect 2967 3448 2971 3452
rect 3463 3451 3467 3455
rect 111 3409 115 3413
rect 135 3412 139 3416
rect 255 3412 259 3416
rect 415 3412 419 3416
rect 575 3412 579 3416
rect 735 3412 739 3416
rect 895 3412 899 3416
rect 1063 3412 1067 3416
rect 1231 3412 1235 3416
rect 1399 3412 1403 3416
rect 1767 3409 1771 3413
rect 1807 3401 1811 3405
rect 2031 3404 2035 3408
rect 2151 3404 2155 3408
rect 2271 3404 2275 3408
rect 2391 3404 2395 3408
rect 2511 3404 2515 3408
rect 2623 3404 2627 3408
rect 2727 3404 2731 3408
rect 2831 3404 2835 3408
rect 2935 3404 2939 3408
rect 3039 3404 3043 3408
rect 3151 3404 3155 3408
rect 3463 3401 3467 3405
rect 111 3392 115 3396
rect 135 3393 139 3397
rect 255 3393 259 3397
rect 415 3393 419 3397
rect 575 3393 579 3397
rect 735 3393 739 3397
rect 895 3393 899 3397
rect 1063 3393 1067 3397
rect 1231 3393 1235 3397
rect 1399 3393 1403 3397
rect 1767 3392 1771 3396
rect 1807 3384 1811 3388
rect 2031 3385 2035 3389
rect 2151 3385 2155 3389
rect 2271 3385 2275 3389
rect 2391 3385 2395 3389
rect 2511 3385 2515 3389
rect 2623 3385 2627 3389
rect 2727 3385 2731 3389
rect 2831 3385 2835 3389
rect 2935 3385 2939 3389
rect 3039 3385 3043 3389
rect 3151 3385 3155 3389
rect 3463 3384 3467 3388
rect 111 3340 115 3344
rect 135 3339 139 3343
rect 327 3339 331 3343
rect 535 3339 539 3343
rect 743 3339 747 3343
rect 935 3339 939 3343
rect 1119 3339 1123 3343
rect 1295 3339 1299 3343
rect 1463 3339 1467 3343
rect 1639 3339 1643 3343
rect 1767 3340 1771 3344
rect 1807 3336 1811 3340
rect 2159 3335 2163 3339
rect 2295 3335 2299 3339
rect 2431 3335 2435 3339
rect 2567 3335 2571 3339
rect 2703 3335 2707 3339
rect 2839 3335 2843 3339
rect 2975 3335 2979 3339
rect 3119 3335 3123 3339
rect 3463 3336 3467 3340
rect 111 3323 115 3327
rect 135 3320 139 3324
rect 327 3320 331 3324
rect 535 3320 539 3324
rect 743 3320 747 3324
rect 935 3320 939 3324
rect 1119 3320 1123 3324
rect 1295 3320 1299 3324
rect 1463 3320 1467 3324
rect 1639 3320 1643 3324
rect 1767 3323 1771 3327
rect 1807 3319 1811 3323
rect 2159 3316 2163 3320
rect 2295 3316 2299 3320
rect 2431 3316 2435 3320
rect 2567 3316 2571 3320
rect 2703 3316 2707 3320
rect 2839 3316 2843 3320
rect 2975 3316 2979 3320
rect 3119 3316 3123 3320
rect 3463 3319 3467 3323
rect 111 3265 115 3269
rect 135 3268 139 3272
rect 279 3268 283 3272
rect 463 3268 467 3272
rect 647 3268 651 3272
rect 831 3268 835 3272
rect 1007 3268 1011 3272
rect 1175 3268 1179 3272
rect 1343 3268 1347 3272
rect 1503 3268 1507 3272
rect 1671 3268 1675 3272
rect 1767 3265 1771 3269
rect 1807 3269 1811 3273
rect 2087 3272 2091 3276
rect 2239 3272 2243 3276
rect 2399 3272 2403 3276
rect 2559 3272 2563 3276
rect 2719 3272 2723 3276
rect 2879 3272 2883 3276
rect 3039 3272 3043 3276
rect 3199 3272 3203 3276
rect 3463 3269 3467 3273
rect 111 3248 115 3252
rect 135 3249 139 3253
rect 279 3249 283 3253
rect 463 3249 467 3253
rect 647 3249 651 3253
rect 831 3249 835 3253
rect 1007 3249 1011 3253
rect 1175 3249 1179 3253
rect 1343 3249 1347 3253
rect 1503 3249 1507 3253
rect 1671 3249 1675 3253
rect 1767 3248 1771 3252
rect 1807 3252 1811 3256
rect 2087 3253 2091 3257
rect 2239 3253 2243 3257
rect 2399 3253 2403 3257
rect 2559 3253 2563 3257
rect 2719 3253 2723 3257
rect 2879 3253 2883 3257
rect 3039 3253 3043 3257
rect 3199 3253 3203 3257
rect 3463 3252 3467 3256
rect 1807 3204 1811 3208
rect 1911 3203 1915 3207
rect 2047 3203 2051 3207
rect 2199 3203 2203 3207
rect 2359 3203 2363 3207
rect 2527 3203 2531 3207
rect 2687 3203 2691 3207
rect 2847 3203 2851 3207
rect 3007 3203 3011 3207
rect 3167 3203 3171 3207
rect 3335 3203 3339 3207
rect 3463 3204 3467 3208
rect 111 3196 115 3200
rect 183 3195 187 3199
rect 327 3195 331 3199
rect 487 3195 491 3199
rect 647 3195 651 3199
rect 807 3195 811 3199
rect 967 3195 971 3199
rect 1135 3195 1139 3199
rect 1303 3195 1307 3199
rect 1471 3195 1475 3199
rect 1767 3196 1771 3200
rect 1807 3187 1811 3191
rect 1911 3184 1915 3188
rect 111 3179 115 3183
rect 2047 3184 2051 3188
rect 2199 3184 2203 3188
rect 2359 3184 2363 3188
rect 2527 3184 2531 3188
rect 2687 3184 2691 3188
rect 2847 3184 2851 3188
rect 3007 3184 3011 3188
rect 3167 3184 3171 3188
rect 3335 3184 3339 3188
rect 3463 3187 3467 3191
rect 183 3176 187 3180
rect 327 3176 331 3180
rect 487 3176 491 3180
rect 647 3176 651 3180
rect 807 3176 811 3180
rect 967 3176 971 3180
rect 1135 3176 1139 3180
rect 1303 3176 1307 3180
rect 1471 3176 1475 3180
rect 1767 3179 1771 3183
rect 1807 3137 1811 3141
rect 1831 3140 1835 3144
rect 2007 3140 2011 3144
rect 2207 3140 2211 3144
rect 2399 3140 2403 3144
rect 2583 3140 2587 3144
rect 2759 3140 2763 3144
rect 2919 3140 2923 3144
rect 3079 3140 3083 3144
rect 3231 3140 3235 3144
rect 3367 3140 3371 3144
rect 111 3129 115 3133
rect 367 3132 371 3136
rect 487 3132 491 3136
rect 607 3132 611 3136
rect 727 3132 731 3136
rect 847 3132 851 3136
rect 967 3132 971 3136
rect 1079 3132 1083 3136
rect 1199 3132 1203 3136
rect 3463 3137 3467 3141
rect 1319 3132 1323 3136
rect 1767 3129 1771 3133
rect 1807 3120 1811 3124
rect 1831 3121 1835 3125
rect 2007 3121 2011 3125
rect 2207 3121 2211 3125
rect 2399 3121 2403 3125
rect 2583 3121 2587 3125
rect 2759 3121 2763 3125
rect 2919 3121 2923 3125
rect 3079 3121 3083 3125
rect 3231 3121 3235 3125
rect 3367 3121 3371 3125
rect 3463 3120 3467 3124
rect 111 3112 115 3116
rect 367 3113 371 3117
rect 487 3113 491 3117
rect 607 3113 611 3117
rect 727 3113 731 3117
rect 847 3113 851 3117
rect 967 3113 971 3117
rect 1079 3113 1083 3117
rect 1199 3113 1203 3117
rect 1319 3113 1323 3117
rect 1767 3112 1771 3116
rect 111 3064 115 3068
rect 439 3063 443 3067
rect 527 3063 531 3067
rect 615 3063 619 3067
rect 703 3063 707 3067
rect 791 3063 795 3067
rect 879 3063 883 3067
rect 967 3063 971 3067
rect 1055 3063 1059 3067
rect 1143 3063 1147 3067
rect 1767 3064 1771 3068
rect 1807 3068 1811 3072
rect 1831 3067 1835 3071
rect 1959 3067 1963 3071
rect 2119 3067 2123 3071
rect 2295 3067 2299 3071
rect 2487 3067 2491 3071
rect 2695 3067 2699 3071
rect 2919 3067 2923 3071
rect 3151 3067 3155 3071
rect 3367 3067 3371 3071
rect 3463 3068 3467 3072
rect 111 3047 115 3051
rect 439 3044 443 3048
rect 527 3044 531 3048
rect 615 3044 619 3048
rect 703 3044 707 3048
rect 791 3044 795 3048
rect 879 3044 883 3048
rect 967 3044 971 3048
rect 1055 3044 1059 3048
rect 1143 3044 1147 3048
rect 1767 3047 1771 3051
rect 1807 3051 1811 3055
rect 1831 3048 1835 3052
rect 1959 3048 1963 3052
rect 2119 3048 2123 3052
rect 2295 3048 2299 3052
rect 2487 3048 2491 3052
rect 2695 3048 2699 3052
rect 2919 3048 2923 3052
rect 3151 3048 3155 3052
rect 3367 3048 3371 3052
rect 3463 3051 3467 3055
rect 111 2989 115 2993
rect 503 2992 507 2996
rect 591 2992 595 2996
rect 679 2992 683 2996
rect 767 2992 771 2996
rect 855 2992 859 2996
rect 943 2992 947 2996
rect 1031 2992 1035 2996
rect 1119 2992 1123 2996
rect 1207 2992 1211 2996
rect 1295 2992 1299 2996
rect 1767 2989 1771 2993
rect 1807 2985 1811 2989
rect 1831 2988 1835 2992
rect 1919 2988 1923 2992
rect 2031 2988 2035 2992
rect 2143 2988 2147 2992
rect 2247 2988 2251 2992
rect 2359 2988 2363 2992
rect 2479 2988 2483 2992
rect 2623 2988 2627 2992
rect 2791 2988 2795 2992
rect 2983 2988 2987 2992
rect 3183 2988 3187 2992
rect 3367 2988 3371 2992
rect 3463 2985 3467 2989
rect 111 2972 115 2976
rect 503 2973 507 2977
rect 591 2973 595 2977
rect 679 2973 683 2977
rect 767 2973 771 2977
rect 855 2973 859 2977
rect 943 2973 947 2977
rect 1031 2973 1035 2977
rect 1119 2973 1123 2977
rect 1207 2973 1211 2977
rect 1295 2973 1299 2977
rect 1767 2972 1771 2976
rect 1807 2968 1811 2972
rect 1831 2969 1835 2973
rect 1919 2969 1923 2973
rect 2031 2969 2035 2973
rect 2143 2969 2147 2973
rect 2247 2969 2251 2973
rect 2359 2969 2363 2973
rect 2479 2969 2483 2973
rect 2623 2969 2627 2973
rect 2791 2969 2795 2973
rect 2983 2969 2987 2973
rect 3183 2969 3187 2973
rect 3367 2969 3371 2973
rect 3463 2968 3467 2972
rect 111 2916 115 2920
rect 327 2915 331 2919
rect 447 2915 451 2919
rect 575 2915 579 2919
rect 711 2915 715 2919
rect 847 2915 851 2919
rect 975 2915 979 2919
rect 1103 2915 1107 2919
rect 1231 2915 1235 2919
rect 1359 2915 1363 2919
rect 1495 2915 1499 2919
rect 1767 2916 1771 2920
rect 1807 2912 1811 2916
rect 1831 2911 1835 2915
rect 2015 2911 2019 2915
rect 2215 2911 2219 2915
rect 2407 2911 2411 2915
rect 2591 2911 2595 2915
rect 2759 2911 2763 2915
rect 2911 2911 2915 2915
rect 3063 2911 3067 2915
rect 3207 2911 3211 2915
rect 3359 2911 3363 2915
rect 3463 2912 3467 2916
rect 111 2899 115 2903
rect 327 2896 331 2900
rect 447 2896 451 2900
rect 575 2896 579 2900
rect 711 2896 715 2900
rect 847 2896 851 2900
rect 975 2896 979 2900
rect 1103 2896 1107 2900
rect 1231 2896 1235 2900
rect 1359 2896 1363 2900
rect 1495 2896 1499 2900
rect 1767 2899 1771 2903
rect 1807 2895 1811 2899
rect 1831 2892 1835 2896
rect 2015 2892 2019 2896
rect 2215 2892 2219 2896
rect 2407 2892 2411 2896
rect 2591 2892 2595 2896
rect 2759 2892 2763 2896
rect 2911 2892 2915 2896
rect 3063 2892 3067 2896
rect 3207 2892 3211 2896
rect 3359 2892 3363 2896
rect 3463 2895 3467 2899
rect 111 2841 115 2845
rect 135 2844 139 2848
rect 255 2844 259 2848
rect 415 2844 419 2848
rect 575 2844 579 2848
rect 735 2844 739 2848
rect 895 2844 899 2848
rect 1047 2844 1051 2848
rect 1191 2844 1195 2848
rect 1343 2844 1347 2848
rect 1495 2844 1499 2848
rect 1767 2841 1771 2845
rect 1807 2845 1811 2849
rect 1831 2848 1835 2852
rect 1999 2848 2003 2852
rect 2191 2848 2195 2852
rect 2383 2848 2387 2852
rect 2567 2848 2571 2852
rect 2735 2848 2739 2852
rect 2903 2848 2907 2852
rect 3063 2848 3067 2852
rect 3223 2848 3227 2852
rect 3367 2848 3371 2852
rect 3463 2845 3467 2849
rect 111 2824 115 2828
rect 135 2825 139 2829
rect 255 2825 259 2829
rect 415 2825 419 2829
rect 575 2825 579 2829
rect 735 2825 739 2829
rect 895 2825 899 2829
rect 1047 2825 1051 2829
rect 1191 2825 1195 2829
rect 1343 2825 1347 2829
rect 1495 2825 1499 2829
rect 1767 2824 1771 2828
rect 1807 2828 1811 2832
rect 1831 2829 1835 2833
rect 1999 2829 2003 2833
rect 2191 2829 2195 2833
rect 2383 2829 2387 2833
rect 2567 2829 2571 2833
rect 2735 2829 2739 2833
rect 2903 2829 2907 2833
rect 3063 2829 3067 2833
rect 3223 2829 3227 2833
rect 3367 2829 3371 2833
rect 3463 2828 3467 2832
rect 1807 2780 1811 2784
rect 1831 2779 1835 2783
rect 2015 2779 2019 2783
rect 2215 2779 2219 2783
rect 2407 2779 2411 2783
rect 2583 2779 2587 2783
rect 2751 2779 2755 2783
rect 2911 2779 2915 2783
rect 3071 2779 3075 2783
rect 3231 2779 3235 2783
rect 3367 2779 3371 2783
rect 3463 2780 3467 2784
rect 111 2768 115 2772
rect 135 2767 139 2771
rect 247 2767 251 2771
rect 391 2767 395 2771
rect 543 2767 547 2771
rect 695 2767 699 2771
rect 855 2767 859 2771
rect 1023 2767 1027 2771
rect 1191 2767 1195 2771
rect 1359 2767 1363 2771
rect 1527 2767 1531 2771
rect 1671 2767 1675 2771
rect 1767 2768 1771 2772
rect 1807 2763 1811 2767
rect 1831 2760 1835 2764
rect 2015 2760 2019 2764
rect 2215 2760 2219 2764
rect 2407 2760 2411 2764
rect 2583 2760 2587 2764
rect 2751 2760 2755 2764
rect 2911 2760 2915 2764
rect 3071 2760 3075 2764
rect 3231 2760 3235 2764
rect 3367 2760 3371 2764
rect 3463 2763 3467 2767
rect 111 2751 115 2755
rect 135 2748 139 2752
rect 247 2748 251 2752
rect 391 2748 395 2752
rect 543 2748 547 2752
rect 695 2748 699 2752
rect 855 2748 859 2752
rect 1023 2748 1027 2752
rect 1191 2748 1195 2752
rect 1359 2748 1363 2752
rect 1527 2748 1531 2752
rect 1671 2748 1675 2752
rect 1767 2751 1771 2755
rect 111 2693 115 2697
rect 247 2696 251 2700
rect 359 2696 363 2700
rect 479 2696 483 2700
rect 615 2696 619 2700
rect 759 2696 763 2700
rect 911 2696 915 2700
rect 1063 2696 1067 2700
rect 1215 2696 1219 2700
rect 1375 2696 1379 2700
rect 1535 2696 1539 2700
rect 1671 2696 1675 2700
rect 1767 2693 1771 2697
rect 1807 2697 1811 2701
rect 2039 2700 2043 2704
rect 2159 2700 2163 2704
rect 2279 2700 2283 2704
rect 2407 2700 2411 2704
rect 2543 2700 2547 2704
rect 2687 2700 2691 2704
rect 2847 2700 2851 2704
rect 3023 2700 3027 2704
rect 3207 2700 3211 2704
rect 3367 2700 3371 2704
rect 3463 2697 3467 2701
rect 111 2676 115 2680
rect 247 2677 251 2681
rect 359 2677 363 2681
rect 479 2677 483 2681
rect 615 2677 619 2681
rect 759 2677 763 2681
rect 911 2677 915 2681
rect 1063 2677 1067 2681
rect 1215 2677 1219 2681
rect 1375 2677 1379 2681
rect 1535 2677 1539 2681
rect 1671 2677 1675 2681
rect 1767 2676 1771 2680
rect 1807 2680 1811 2684
rect 2039 2681 2043 2685
rect 2159 2681 2163 2685
rect 2279 2681 2283 2685
rect 2407 2681 2411 2685
rect 2543 2681 2547 2685
rect 2687 2681 2691 2685
rect 2847 2681 2851 2685
rect 3023 2681 3027 2685
rect 3207 2681 3211 2685
rect 3367 2681 3371 2685
rect 3463 2680 3467 2684
rect 111 2624 115 2628
rect 463 2623 467 2627
rect 551 2623 555 2627
rect 639 2623 643 2627
rect 743 2623 747 2627
rect 855 2623 859 2627
rect 983 2623 987 2627
rect 1127 2623 1131 2627
rect 1279 2623 1283 2627
rect 1439 2623 1443 2627
rect 1607 2623 1611 2627
rect 1767 2624 1771 2628
rect 1807 2624 1811 2628
rect 1871 2623 1875 2627
rect 1967 2623 1971 2627
rect 2071 2623 2075 2627
rect 2183 2623 2187 2627
rect 2295 2623 2299 2627
rect 2431 2623 2435 2627
rect 2583 2623 2587 2627
rect 2759 2623 2763 2627
rect 2959 2623 2963 2627
rect 3167 2623 3171 2627
rect 3367 2623 3371 2627
rect 3463 2624 3467 2628
rect 111 2607 115 2611
rect 463 2604 467 2608
rect 551 2604 555 2608
rect 639 2604 643 2608
rect 743 2604 747 2608
rect 855 2604 859 2608
rect 983 2604 987 2608
rect 1127 2604 1131 2608
rect 1279 2604 1283 2608
rect 1439 2604 1443 2608
rect 1607 2604 1611 2608
rect 1767 2607 1771 2611
rect 1807 2607 1811 2611
rect 1871 2604 1875 2608
rect 1967 2604 1971 2608
rect 2071 2604 2075 2608
rect 2183 2604 2187 2608
rect 2295 2604 2299 2608
rect 2431 2604 2435 2608
rect 2583 2604 2587 2608
rect 2759 2604 2763 2608
rect 2959 2604 2963 2608
rect 3167 2604 3171 2608
rect 3367 2604 3371 2608
rect 3463 2607 3467 2611
rect 111 2549 115 2553
rect 503 2552 507 2556
rect 591 2552 595 2556
rect 679 2552 683 2556
rect 775 2552 779 2556
rect 879 2552 883 2556
rect 991 2552 995 2556
rect 1103 2552 1107 2556
rect 1223 2552 1227 2556
rect 1351 2552 1355 2556
rect 1479 2552 1483 2556
rect 1607 2552 1611 2556
rect 1767 2549 1771 2553
rect 1807 2545 1811 2549
rect 1831 2548 1835 2552
rect 1919 2548 1923 2552
rect 2007 2548 2011 2552
rect 2111 2548 2115 2552
rect 2223 2548 2227 2552
rect 2343 2548 2347 2552
rect 2487 2548 2491 2552
rect 2647 2548 2651 2552
rect 2815 2548 2819 2552
rect 2999 2548 3003 2552
rect 3191 2548 3195 2552
rect 3367 2548 3371 2552
rect 3463 2545 3467 2549
rect 111 2532 115 2536
rect 503 2533 507 2537
rect 591 2533 595 2537
rect 679 2533 683 2537
rect 775 2533 779 2537
rect 879 2533 883 2537
rect 991 2533 995 2537
rect 1103 2533 1107 2537
rect 1223 2533 1227 2537
rect 1351 2533 1355 2537
rect 1479 2533 1483 2537
rect 1607 2533 1611 2537
rect 1767 2532 1771 2536
rect 1807 2528 1811 2532
rect 1831 2529 1835 2533
rect 1919 2529 1923 2533
rect 2007 2529 2011 2533
rect 2111 2529 2115 2533
rect 2223 2529 2227 2533
rect 2343 2529 2347 2533
rect 2487 2529 2491 2533
rect 2647 2529 2651 2533
rect 2815 2529 2819 2533
rect 2999 2529 3003 2533
rect 3191 2529 3195 2533
rect 3367 2529 3371 2533
rect 3463 2528 3467 2532
rect 111 2480 115 2484
rect 551 2479 555 2483
rect 735 2479 739 2483
rect 911 2479 915 2483
rect 1079 2479 1083 2483
rect 1239 2479 1243 2483
rect 1399 2479 1403 2483
rect 1567 2479 1571 2483
rect 1767 2480 1771 2484
rect 1807 2484 1811 2488
rect 1951 2483 1955 2487
rect 2039 2483 2043 2487
rect 2135 2483 2139 2487
rect 2239 2483 2243 2487
rect 2367 2483 2371 2487
rect 2527 2483 2531 2487
rect 2711 2483 2715 2487
rect 2919 2483 2923 2487
rect 3143 2483 3147 2487
rect 3367 2483 3371 2487
rect 3463 2484 3467 2488
rect 111 2463 115 2467
rect 551 2460 555 2464
rect 735 2460 739 2464
rect 911 2460 915 2464
rect 1079 2460 1083 2464
rect 1239 2460 1243 2464
rect 1399 2460 1403 2464
rect 1567 2460 1571 2464
rect 1767 2463 1771 2467
rect 1807 2467 1811 2471
rect 1951 2464 1955 2468
rect 2039 2464 2043 2468
rect 2135 2464 2139 2468
rect 2239 2464 2243 2468
rect 2367 2464 2371 2468
rect 2527 2464 2531 2468
rect 2711 2464 2715 2468
rect 2919 2464 2923 2468
rect 3143 2464 3147 2468
rect 3367 2464 3371 2468
rect 3463 2467 3467 2471
rect 111 2413 115 2417
rect 415 2416 419 2420
rect 503 2416 507 2420
rect 599 2416 603 2420
rect 703 2416 707 2420
rect 807 2416 811 2420
rect 919 2416 923 2420
rect 1039 2416 1043 2420
rect 1167 2416 1171 2420
rect 1295 2416 1299 2420
rect 1423 2416 1427 2420
rect 1767 2413 1771 2417
rect 1807 2409 1811 2413
rect 2215 2412 2219 2416
rect 2303 2412 2307 2416
rect 2391 2412 2395 2416
rect 2479 2412 2483 2416
rect 2567 2412 2571 2416
rect 2655 2412 2659 2416
rect 2743 2412 2747 2416
rect 2839 2412 2843 2416
rect 2935 2412 2939 2416
rect 3463 2409 3467 2413
rect 111 2396 115 2400
rect 415 2397 419 2401
rect 503 2397 507 2401
rect 599 2397 603 2401
rect 703 2397 707 2401
rect 807 2397 811 2401
rect 919 2397 923 2401
rect 1039 2397 1043 2401
rect 1167 2397 1171 2401
rect 1295 2397 1299 2401
rect 1423 2397 1427 2401
rect 1767 2396 1771 2400
rect 1807 2392 1811 2396
rect 2215 2393 2219 2397
rect 2303 2393 2307 2397
rect 2391 2393 2395 2397
rect 2479 2393 2483 2397
rect 2567 2393 2571 2397
rect 2655 2393 2659 2397
rect 2743 2393 2747 2397
rect 2839 2393 2843 2397
rect 2935 2393 2939 2397
rect 3463 2392 3467 2396
rect 111 2348 115 2352
rect 319 2347 323 2351
rect 431 2347 435 2351
rect 543 2347 547 2351
rect 655 2347 659 2351
rect 767 2347 771 2351
rect 879 2347 883 2351
rect 991 2347 995 2351
rect 1103 2347 1107 2351
rect 1215 2347 1219 2351
rect 1335 2347 1339 2351
rect 1767 2348 1771 2352
rect 1807 2348 1811 2352
rect 2167 2347 2171 2351
rect 2263 2347 2267 2351
rect 2367 2347 2371 2351
rect 2471 2347 2475 2351
rect 2575 2347 2579 2351
rect 2687 2347 2691 2351
rect 2799 2347 2803 2351
rect 2911 2347 2915 2351
rect 3023 2347 3027 2351
rect 3463 2348 3467 2352
rect 111 2331 115 2335
rect 319 2328 323 2332
rect 431 2328 435 2332
rect 543 2328 547 2332
rect 655 2328 659 2332
rect 767 2328 771 2332
rect 879 2328 883 2332
rect 991 2328 995 2332
rect 1103 2328 1107 2332
rect 1215 2328 1219 2332
rect 1335 2328 1339 2332
rect 1767 2331 1771 2335
rect 1807 2331 1811 2335
rect 2167 2328 2171 2332
rect 2263 2328 2267 2332
rect 2367 2328 2371 2332
rect 2471 2328 2475 2332
rect 2575 2328 2579 2332
rect 2687 2328 2691 2332
rect 2799 2328 2803 2332
rect 2911 2328 2915 2332
rect 3023 2328 3027 2332
rect 3463 2331 3467 2335
rect 111 2273 115 2277
rect 151 2276 155 2280
rect 271 2276 275 2280
rect 391 2276 395 2280
rect 519 2276 523 2280
rect 647 2276 651 2280
rect 775 2276 779 2280
rect 895 2276 899 2280
rect 1015 2276 1019 2280
rect 1143 2276 1147 2280
rect 1271 2276 1275 2280
rect 1767 2273 1771 2277
rect 1807 2273 1811 2277
rect 1887 2276 1891 2280
rect 2039 2276 2043 2280
rect 2199 2276 2203 2280
rect 2375 2276 2379 2280
rect 2551 2276 2555 2280
rect 2719 2276 2723 2280
rect 2887 2276 2891 2280
rect 3055 2276 3059 2280
rect 3223 2276 3227 2280
rect 3367 2276 3371 2280
rect 3463 2273 3467 2277
rect 111 2256 115 2260
rect 151 2257 155 2261
rect 271 2257 275 2261
rect 391 2257 395 2261
rect 519 2257 523 2261
rect 647 2257 651 2261
rect 775 2257 779 2261
rect 895 2257 899 2261
rect 1015 2257 1019 2261
rect 1143 2257 1147 2261
rect 1271 2257 1275 2261
rect 1767 2256 1771 2260
rect 1807 2256 1811 2260
rect 1887 2257 1891 2261
rect 2039 2257 2043 2261
rect 2199 2257 2203 2261
rect 2375 2257 2379 2261
rect 2551 2257 2555 2261
rect 2719 2257 2723 2261
rect 2887 2257 2891 2261
rect 3055 2257 3059 2261
rect 3223 2257 3227 2261
rect 3367 2257 3371 2261
rect 3463 2256 3467 2260
rect 111 2208 115 2212
rect 135 2207 139 2211
rect 247 2207 251 2211
rect 407 2207 411 2211
rect 583 2207 587 2211
rect 767 2207 771 2211
rect 951 2207 955 2211
rect 1135 2207 1139 2211
rect 1319 2207 1323 2211
rect 1503 2207 1507 2211
rect 1671 2207 1675 2211
rect 1767 2208 1771 2212
rect 1807 2212 1811 2216
rect 1831 2211 1835 2215
rect 1967 2211 1971 2215
rect 2135 2211 2139 2215
rect 2311 2211 2315 2215
rect 2487 2211 2491 2215
rect 2655 2211 2659 2215
rect 2815 2211 2819 2215
rect 2959 2211 2963 2215
rect 3103 2211 3107 2215
rect 3247 2211 3251 2215
rect 3367 2211 3371 2215
rect 3463 2212 3467 2216
rect 111 2191 115 2195
rect 135 2188 139 2192
rect 247 2188 251 2192
rect 407 2188 411 2192
rect 583 2188 587 2192
rect 767 2188 771 2192
rect 951 2188 955 2192
rect 1135 2188 1139 2192
rect 1319 2188 1323 2192
rect 1503 2188 1507 2192
rect 1671 2188 1675 2192
rect 1767 2191 1771 2195
rect 1807 2195 1811 2199
rect 1831 2192 1835 2196
rect 1967 2192 1971 2196
rect 2135 2192 2139 2196
rect 2311 2192 2315 2196
rect 2487 2192 2491 2196
rect 2655 2192 2659 2196
rect 2815 2192 2819 2196
rect 2959 2192 2963 2196
rect 3103 2192 3107 2196
rect 3247 2192 3251 2196
rect 3367 2192 3371 2196
rect 3463 2195 3467 2199
rect 1807 2145 1811 2149
rect 2927 2148 2931 2152
rect 3015 2148 3019 2152
rect 3103 2148 3107 2152
rect 3191 2148 3195 2152
rect 3279 2148 3283 2152
rect 3367 2148 3371 2152
rect 3463 2145 3467 2149
rect 111 2133 115 2137
rect 135 2136 139 2140
rect 247 2136 251 2140
rect 391 2136 395 2140
rect 543 2136 547 2140
rect 695 2136 699 2140
rect 839 2136 843 2140
rect 975 2136 979 2140
rect 1103 2136 1107 2140
rect 1231 2136 1235 2140
rect 1351 2136 1355 2140
rect 1463 2136 1467 2140
rect 1575 2136 1579 2140
rect 1671 2136 1675 2140
rect 1767 2133 1771 2137
rect 1807 2128 1811 2132
rect 2927 2129 2931 2133
rect 3015 2129 3019 2133
rect 3103 2129 3107 2133
rect 3191 2129 3195 2133
rect 3279 2129 3283 2133
rect 3367 2129 3371 2133
rect 3463 2128 3467 2132
rect 111 2116 115 2120
rect 135 2117 139 2121
rect 247 2117 251 2121
rect 391 2117 395 2121
rect 543 2117 547 2121
rect 695 2117 699 2121
rect 839 2117 843 2121
rect 975 2117 979 2121
rect 1103 2117 1107 2121
rect 1231 2117 1235 2121
rect 1351 2117 1355 2121
rect 1463 2117 1467 2121
rect 1575 2117 1579 2121
rect 1671 2117 1675 2121
rect 1767 2116 1771 2120
rect 1807 2076 1811 2080
rect 1831 2075 1835 2079
rect 1991 2075 1995 2079
rect 2167 2075 2171 2079
rect 2343 2075 2347 2079
rect 2503 2075 2507 2079
rect 2655 2075 2659 2079
rect 2791 2075 2795 2079
rect 2919 2075 2923 2079
rect 3039 2075 3043 2079
rect 3159 2075 3163 2079
rect 3271 2075 3275 2079
rect 3367 2075 3371 2079
rect 3463 2076 3467 2080
rect 111 2068 115 2072
rect 135 2067 139 2071
rect 223 2067 227 2071
rect 343 2067 347 2071
rect 463 2067 467 2071
rect 583 2067 587 2071
rect 703 2067 707 2071
rect 823 2067 827 2071
rect 935 2067 939 2071
rect 1047 2067 1051 2071
rect 1159 2067 1163 2071
rect 1279 2067 1283 2071
rect 1767 2068 1771 2072
rect 1807 2059 1811 2063
rect 1831 2056 1835 2060
rect 111 2051 115 2055
rect 1991 2056 1995 2060
rect 2167 2056 2171 2060
rect 2343 2056 2347 2060
rect 2503 2056 2507 2060
rect 2655 2056 2659 2060
rect 2791 2056 2795 2060
rect 2919 2056 2923 2060
rect 3039 2056 3043 2060
rect 3159 2056 3163 2060
rect 3271 2056 3275 2060
rect 3367 2056 3371 2060
rect 3463 2059 3467 2063
rect 135 2048 139 2052
rect 223 2048 227 2052
rect 343 2048 347 2052
rect 463 2048 467 2052
rect 583 2048 587 2052
rect 703 2048 707 2052
rect 823 2048 827 2052
rect 935 2048 939 2052
rect 1047 2048 1051 2052
rect 1159 2048 1163 2052
rect 1279 2048 1283 2052
rect 1767 2051 1771 2055
rect 1807 2005 1811 2009
rect 1831 2008 1835 2012
rect 2015 2008 2019 2012
rect 2223 2008 2227 2012
rect 2431 2008 2435 2012
rect 2631 2008 2635 2012
rect 2823 2008 2827 2012
rect 3007 2008 3011 2012
rect 3199 2008 3203 2012
rect 3367 2008 3371 2012
rect 3463 2005 3467 2009
rect 111 1993 115 1997
rect 135 1996 139 2000
rect 239 1996 243 2000
rect 367 1996 371 2000
rect 503 1996 507 2000
rect 639 1996 643 2000
rect 775 1996 779 2000
rect 911 1996 915 2000
rect 1047 1996 1051 2000
rect 1183 1996 1187 2000
rect 1327 1996 1331 2000
rect 1767 1993 1771 1997
rect 1807 1988 1811 1992
rect 1831 1989 1835 1993
rect 2015 1989 2019 1993
rect 2223 1989 2227 1993
rect 2431 1989 2435 1993
rect 2631 1989 2635 1993
rect 2823 1989 2827 1993
rect 3007 1989 3011 1993
rect 3199 1989 3203 1993
rect 3367 1989 3371 1993
rect 3463 1988 3467 1992
rect 111 1976 115 1980
rect 135 1977 139 1981
rect 239 1977 243 1981
rect 367 1977 371 1981
rect 503 1977 507 1981
rect 639 1977 643 1981
rect 775 1977 779 1981
rect 911 1977 915 1981
rect 1047 1977 1051 1981
rect 1183 1977 1187 1981
rect 1327 1977 1331 1981
rect 1767 1976 1771 1980
rect 1807 1940 1811 1944
rect 1863 1939 1867 1943
rect 1999 1939 2003 1943
rect 2143 1939 2147 1943
rect 2287 1939 2291 1943
rect 2431 1939 2435 1943
rect 2575 1939 2579 1943
rect 2711 1939 2715 1943
rect 2831 1939 2835 1943
rect 2951 1939 2955 1943
rect 3063 1939 3067 1943
rect 3167 1939 3171 1943
rect 3279 1939 3283 1943
rect 3367 1939 3371 1943
rect 3463 1940 3467 1944
rect 111 1928 115 1932
rect 295 1927 299 1931
rect 423 1927 427 1931
rect 559 1927 563 1931
rect 703 1927 707 1931
rect 855 1927 859 1931
rect 1007 1927 1011 1931
rect 1159 1927 1163 1931
rect 1311 1927 1315 1931
rect 1471 1927 1475 1931
rect 1767 1928 1771 1932
rect 1807 1923 1811 1927
rect 1863 1920 1867 1924
rect 1999 1920 2003 1924
rect 2143 1920 2147 1924
rect 2287 1920 2291 1924
rect 2431 1920 2435 1924
rect 2575 1920 2579 1924
rect 2711 1920 2715 1924
rect 2831 1920 2835 1924
rect 2951 1920 2955 1924
rect 3063 1920 3067 1924
rect 3167 1920 3171 1924
rect 3279 1920 3283 1924
rect 3367 1920 3371 1924
rect 3463 1923 3467 1927
rect 111 1911 115 1915
rect 295 1908 299 1912
rect 423 1908 427 1912
rect 559 1908 563 1912
rect 703 1908 707 1912
rect 855 1908 859 1912
rect 1007 1908 1011 1912
rect 1159 1908 1163 1912
rect 1311 1908 1315 1912
rect 1471 1908 1475 1912
rect 1767 1911 1771 1915
rect 1807 1869 1811 1873
rect 2015 1872 2019 1876
rect 2111 1872 2115 1876
rect 2215 1872 2219 1876
rect 2327 1872 2331 1876
rect 2439 1872 2443 1876
rect 2543 1872 2547 1876
rect 2647 1872 2651 1876
rect 2759 1872 2763 1876
rect 2871 1872 2875 1876
rect 2983 1872 2987 1876
rect 111 1861 115 1865
rect 431 1864 435 1868
rect 575 1864 579 1868
rect 727 1864 731 1868
rect 887 1864 891 1868
rect 1047 1864 1051 1868
rect 1199 1864 1203 1868
rect 1351 1864 1355 1868
rect 1511 1864 1515 1868
rect 3463 1869 3467 1873
rect 1671 1864 1675 1868
rect 1767 1861 1771 1865
rect 1807 1852 1811 1856
rect 2015 1853 2019 1857
rect 2111 1853 2115 1857
rect 2215 1853 2219 1857
rect 2327 1853 2331 1857
rect 2439 1853 2443 1857
rect 2543 1853 2547 1857
rect 2647 1853 2651 1857
rect 2759 1853 2763 1857
rect 2871 1853 2875 1857
rect 2983 1853 2987 1857
rect 3463 1852 3467 1856
rect 111 1844 115 1848
rect 431 1845 435 1849
rect 575 1845 579 1849
rect 727 1845 731 1849
rect 887 1845 891 1849
rect 1047 1845 1051 1849
rect 1199 1845 1203 1849
rect 1351 1845 1355 1849
rect 1511 1845 1515 1849
rect 1671 1845 1675 1849
rect 1767 1844 1771 1848
rect 111 1796 115 1800
rect 511 1795 515 1799
rect 631 1795 635 1799
rect 759 1795 763 1799
rect 887 1795 891 1799
rect 1023 1795 1027 1799
rect 1151 1795 1155 1799
rect 1279 1795 1283 1799
rect 1407 1795 1411 1799
rect 1535 1795 1539 1799
rect 1671 1795 1675 1799
rect 1767 1796 1771 1800
rect 1807 1800 1811 1804
rect 2103 1799 2107 1803
rect 2191 1799 2195 1803
rect 2279 1799 2283 1803
rect 2367 1799 2371 1803
rect 2455 1799 2459 1803
rect 2543 1799 2547 1803
rect 2631 1799 2635 1803
rect 2719 1799 2723 1803
rect 2807 1799 2811 1803
rect 2895 1799 2899 1803
rect 3463 1800 3467 1804
rect 111 1779 115 1783
rect 511 1776 515 1780
rect 631 1776 635 1780
rect 759 1776 763 1780
rect 887 1776 891 1780
rect 1023 1776 1027 1780
rect 1151 1776 1155 1780
rect 1279 1776 1283 1780
rect 1407 1776 1411 1780
rect 1535 1776 1539 1780
rect 1671 1776 1675 1780
rect 1767 1779 1771 1783
rect 1807 1783 1811 1787
rect 2103 1780 2107 1784
rect 2191 1780 2195 1784
rect 2279 1780 2283 1784
rect 2367 1780 2371 1784
rect 2455 1780 2459 1784
rect 2543 1780 2547 1784
rect 2631 1780 2635 1784
rect 2719 1780 2723 1784
rect 2807 1780 2811 1784
rect 2895 1780 2899 1784
rect 3463 1783 3467 1787
rect 111 1725 115 1729
rect 439 1728 443 1732
rect 535 1728 539 1732
rect 639 1728 643 1732
rect 743 1728 747 1732
rect 847 1728 851 1732
rect 951 1728 955 1732
rect 1055 1728 1059 1732
rect 1159 1728 1163 1732
rect 1271 1728 1275 1732
rect 1383 1728 1387 1732
rect 1767 1725 1771 1729
rect 1807 1721 1811 1725
rect 2143 1724 2147 1728
rect 2231 1724 2235 1728
rect 2319 1724 2323 1728
rect 2407 1724 2411 1728
rect 2495 1724 2499 1728
rect 2583 1724 2587 1728
rect 2671 1724 2675 1728
rect 2759 1724 2763 1728
rect 2847 1724 2851 1728
rect 3463 1721 3467 1725
rect 111 1708 115 1712
rect 439 1709 443 1713
rect 535 1709 539 1713
rect 639 1709 643 1713
rect 743 1709 747 1713
rect 847 1709 851 1713
rect 951 1709 955 1713
rect 1055 1709 1059 1713
rect 1159 1709 1163 1713
rect 1271 1709 1275 1713
rect 1383 1709 1387 1713
rect 1767 1708 1771 1712
rect 1807 1704 1811 1708
rect 2143 1705 2147 1709
rect 2231 1705 2235 1709
rect 2319 1705 2323 1709
rect 2407 1705 2411 1709
rect 2495 1705 2499 1709
rect 2583 1705 2587 1709
rect 2671 1705 2675 1709
rect 2759 1705 2763 1709
rect 2847 1705 2851 1709
rect 3463 1704 3467 1708
rect 111 1660 115 1664
rect 399 1659 403 1663
rect 487 1659 491 1663
rect 575 1659 579 1663
rect 663 1659 667 1663
rect 759 1659 763 1663
rect 855 1659 859 1663
rect 951 1659 955 1663
rect 1047 1659 1051 1663
rect 1143 1659 1147 1663
rect 1767 1660 1771 1664
rect 1807 1656 1811 1660
rect 2103 1655 2107 1659
rect 2191 1655 2195 1659
rect 2279 1655 2283 1659
rect 2367 1655 2371 1659
rect 2455 1655 2459 1659
rect 2543 1655 2547 1659
rect 2631 1655 2635 1659
rect 2719 1655 2723 1659
rect 2807 1655 2811 1659
rect 2895 1655 2899 1659
rect 3463 1656 3467 1660
rect 111 1643 115 1647
rect 399 1640 403 1644
rect 487 1640 491 1644
rect 575 1640 579 1644
rect 663 1640 667 1644
rect 759 1640 763 1644
rect 855 1640 859 1644
rect 951 1640 955 1644
rect 1047 1640 1051 1644
rect 1143 1640 1147 1644
rect 1767 1643 1771 1647
rect 1807 1639 1811 1643
rect 2103 1636 2107 1640
rect 2191 1636 2195 1640
rect 2279 1636 2283 1640
rect 2367 1636 2371 1640
rect 2455 1636 2459 1640
rect 2543 1636 2547 1640
rect 2631 1636 2635 1640
rect 2719 1636 2723 1640
rect 2807 1636 2811 1640
rect 2895 1636 2899 1640
rect 3463 1639 3467 1643
rect 111 1589 115 1593
rect 279 1592 283 1596
rect 383 1592 387 1596
rect 495 1592 499 1596
rect 607 1592 611 1596
rect 719 1592 723 1596
rect 831 1592 835 1596
rect 943 1592 947 1596
rect 1055 1592 1059 1596
rect 1167 1592 1171 1596
rect 1279 1592 1283 1596
rect 1767 1589 1771 1593
rect 1807 1585 1811 1589
rect 2063 1588 2067 1592
rect 2159 1588 2163 1592
rect 2255 1588 2259 1592
rect 2359 1588 2363 1592
rect 2463 1588 2467 1592
rect 2567 1588 2571 1592
rect 2671 1588 2675 1592
rect 2775 1588 2779 1592
rect 2887 1588 2891 1592
rect 3463 1585 3467 1589
rect 111 1572 115 1576
rect 279 1573 283 1577
rect 383 1573 387 1577
rect 495 1573 499 1577
rect 607 1573 611 1577
rect 719 1573 723 1577
rect 831 1573 835 1577
rect 943 1573 947 1577
rect 1055 1573 1059 1577
rect 1167 1573 1171 1577
rect 1279 1573 1283 1577
rect 1767 1572 1771 1576
rect 1807 1568 1811 1572
rect 2063 1569 2067 1573
rect 2159 1569 2163 1573
rect 2255 1569 2259 1573
rect 2359 1569 2363 1573
rect 2463 1569 2467 1573
rect 2567 1569 2571 1573
rect 2671 1569 2675 1573
rect 2775 1569 2779 1573
rect 2887 1569 2891 1573
rect 3463 1568 3467 1572
rect 111 1520 115 1524
rect 183 1519 187 1523
rect 327 1519 331 1523
rect 471 1519 475 1523
rect 623 1519 627 1523
rect 767 1519 771 1523
rect 911 1519 915 1523
rect 1047 1519 1051 1523
rect 1175 1519 1179 1523
rect 1311 1519 1315 1523
rect 1447 1519 1451 1523
rect 1767 1520 1771 1524
rect 1807 1524 1811 1528
rect 1919 1523 1923 1527
rect 2039 1523 2043 1527
rect 2167 1523 2171 1527
rect 2295 1523 2299 1527
rect 2423 1523 2427 1527
rect 2551 1523 2555 1527
rect 2679 1523 2683 1527
rect 2799 1523 2803 1527
rect 2927 1523 2931 1527
rect 3055 1523 3059 1527
rect 3463 1524 3467 1528
rect 111 1503 115 1507
rect 183 1500 187 1504
rect 327 1500 331 1504
rect 471 1500 475 1504
rect 623 1500 627 1504
rect 767 1500 771 1504
rect 911 1500 915 1504
rect 1047 1500 1051 1504
rect 1175 1500 1179 1504
rect 1311 1500 1315 1504
rect 1447 1500 1451 1504
rect 1767 1503 1771 1507
rect 1807 1507 1811 1511
rect 1919 1504 1923 1508
rect 2039 1504 2043 1508
rect 2167 1504 2171 1508
rect 2295 1504 2299 1508
rect 2423 1504 2427 1508
rect 2551 1504 2555 1508
rect 2679 1504 2683 1508
rect 2799 1504 2803 1508
rect 2927 1504 2931 1508
rect 3055 1504 3059 1508
rect 3463 1507 3467 1511
rect 111 1449 115 1453
rect 159 1452 163 1456
rect 375 1452 379 1456
rect 583 1452 587 1456
rect 783 1452 787 1456
rect 959 1452 963 1456
rect 1127 1452 1131 1456
rect 1279 1452 1283 1456
rect 1431 1452 1435 1456
rect 1591 1452 1595 1456
rect 1767 1449 1771 1453
rect 1807 1449 1811 1453
rect 1831 1452 1835 1456
rect 1951 1452 1955 1456
rect 2111 1452 2115 1456
rect 2271 1452 2275 1456
rect 2431 1452 2435 1456
rect 2591 1452 2595 1456
rect 2735 1452 2739 1456
rect 2871 1452 2875 1456
rect 3007 1452 3011 1456
rect 3135 1452 3139 1456
rect 3263 1452 3267 1456
rect 3367 1452 3371 1456
rect 3463 1449 3467 1453
rect 111 1432 115 1436
rect 159 1433 163 1437
rect 375 1433 379 1437
rect 583 1433 587 1437
rect 783 1433 787 1437
rect 959 1433 963 1437
rect 1127 1433 1131 1437
rect 1279 1433 1283 1437
rect 1431 1433 1435 1437
rect 1591 1433 1595 1437
rect 1767 1432 1771 1436
rect 1807 1432 1811 1436
rect 1831 1433 1835 1437
rect 1951 1433 1955 1437
rect 2111 1433 2115 1437
rect 2271 1433 2275 1437
rect 2431 1433 2435 1437
rect 2591 1433 2595 1437
rect 2735 1433 2739 1437
rect 2871 1433 2875 1437
rect 3007 1433 3011 1437
rect 3135 1433 3139 1437
rect 3263 1433 3267 1437
rect 3367 1433 3371 1437
rect 3463 1432 3467 1436
rect 111 1384 115 1388
rect 135 1383 139 1387
rect 303 1383 307 1387
rect 495 1383 499 1387
rect 679 1383 683 1387
rect 855 1383 859 1387
rect 1015 1383 1019 1387
rect 1167 1383 1171 1387
rect 1303 1383 1307 1387
rect 1431 1383 1435 1387
rect 1559 1383 1563 1387
rect 1671 1383 1675 1387
rect 1767 1384 1771 1388
rect 1807 1384 1811 1388
rect 1831 1383 1835 1387
rect 2007 1383 2011 1387
rect 2199 1383 2203 1387
rect 2383 1383 2387 1387
rect 2559 1383 2563 1387
rect 2719 1383 2723 1387
rect 2863 1383 2867 1387
rect 2999 1383 3003 1387
rect 3127 1383 3131 1387
rect 3255 1383 3259 1387
rect 3367 1383 3371 1387
rect 3463 1384 3467 1388
rect 111 1367 115 1371
rect 135 1364 139 1368
rect 303 1364 307 1368
rect 495 1364 499 1368
rect 679 1364 683 1368
rect 855 1364 859 1368
rect 1015 1364 1019 1368
rect 1167 1364 1171 1368
rect 1303 1364 1307 1368
rect 1431 1364 1435 1368
rect 1559 1364 1563 1368
rect 1671 1364 1675 1368
rect 1767 1367 1771 1371
rect 1807 1367 1811 1371
rect 1831 1364 1835 1368
rect 2007 1364 2011 1368
rect 2199 1364 2203 1368
rect 2383 1364 2387 1368
rect 2559 1364 2563 1368
rect 2719 1364 2723 1368
rect 2863 1364 2867 1368
rect 2999 1364 3003 1368
rect 3127 1364 3131 1368
rect 3255 1364 3259 1368
rect 3367 1364 3371 1368
rect 3463 1367 3467 1371
rect 111 1313 115 1317
rect 135 1316 139 1320
rect 247 1316 251 1320
rect 399 1316 403 1320
rect 559 1316 563 1320
rect 727 1316 731 1320
rect 895 1316 899 1320
rect 1063 1316 1067 1320
rect 1223 1316 1227 1320
rect 1375 1316 1379 1320
rect 1535 1316 1539 1320
rect 1671 1316 1675 1320
rect 1767 1313 1771 1317
rect 1807 1309 1811 1313
rect 1831 1312 1835 1316
rect 1967 1312 1971 1316
rect 2143 1312 2147 1316
rect 2327 1312 2331 1316
rect 2511 1312 2515 1316
rect 2687 1312 2691 1316
rect 2863 1312 2867 1316
rect 3039 1312 3043 1316
rect 3215 1312 3219 1316
rect 3367 1312 3371 1316
rect 3463 1309 3467 1313
rect 111 1296 115 1300
rect 135 1297 139 1301
rect 247 1297 251 1301
rect 399 1297 403 1301
rect 559 1297 563 1301
rect 727 1297 731 1301
rect 895 1297 899 1301
rect 1063 1297 1067 1301
rect 1223 1297 1227 1301
rect 1375 1297 1379 1301
rect 1535 1297 1539 1301
rect 1671 1297 1675 1301
rect 1767 1296 1771 1300
rect 1807 1292 1811 1296
rect 1831 1293 1835 1297
rect 1967 1293 1971 1297
rect 2143 1293 2147 1297
rect 2327 1293 2331 1297
rect 2511 1293 2515 1297
rect 2687 1293 2691 1297
rect 2863 1293 2867 1297
rect 3039 1293 3043 1297
rect 3215 1293 3219 1297
rect 3367 1293 3371 1297
rect 3463 1292 3467 1296
rect 111 1248 115 1252
rect 135 1247 139 1251
rect 223 1247 227 1251
rect 319 1247 323 1251
rect 431 1247 435 1251
rect 551 1247 555 1251
rect 679 1247 683 1251
rect 823 1247 827 1251
rect 975 1247 979 1251
rect 1143 1247 1147 1251
rect 1319 1247 1323 1251
rect 1503 1247 1507 1251
rect 1671 1247 1675 1251
rect 1767 1248 1771 1252
rect 1807 1248 1811 1252
rect 1831 1247 1835 1251
rect 2095 1247 2099 1251
rect 2359 1247 2363 1251
rect 2599 1247 2603 1251
rect 2807 1247 2811 1251
rect 3007 1247 3011 1251
rect 3199 1247 3203 1251
rect 3367 1247 3371 1251
rect 3463 1248 3467 1252
rect 111 1231 115 1235
rect 135 1228 139 1232
rect 223 1228 227 1232
rect 319 1228 323 1232
rect 431 1228 435 1232
rect 551 1228 555 1232
rect 679 1228 683 1232
rect 823 1228 827 1232
rect 975 1228 979 1232
rect 1143 1228 1147 1232
rect 1319 1228 1323 1232
rect 1503 1228 1507 1232
rect 1671 1228 1675 1232
rect 1767 1231 1771 1235
rect 1807 1231 1811 1235
rect 1831 1228 1835 1232
rect 2095 1228 2099 1232
rect 2359 1228 2363 1232
rect 2599 1228 2603 1232
rect 2807 1228 2811 1232
rect 3007 1228 3011 1232
rect 3199 1228 3203 1232
rect 3367 1228 3371 1232
rect 3463 1231 3467 1235
rect 111 1173 115 1177
rect 135 1176 139 1180
rect 231 1176 235 1180
rect 359 1176 363 1180
rect 487 1176 491 1180
rect 615 1176 619 1180
rect 743 1176 747 1180
rect 871 1176 875 1180
rect 991 1176 995 1180
rect 1119 1176 1123 1180
rect 1247 1176 1251 1180
rect 1767 1173 1771 1177
rect 1807 1173 1811 1177
rect 1935 1176 1939 1180
rect 2039 1176 2043 1180
rect 2159 1176 2163 1180
rect 2287 1176 2291 1180
rect 2423 1176 2427 1180
rect 2567 1176 2571 1180
rect 2703 1176 2707 1180
rect 2839 1176 2843 1180
rect 2975 1176 2979 1180
rect 3111 1176 3115 1180
rect 3247 1176 3251 1180
rect 3367 1176 3371 1180
rect 3463 1173 3467 1177
rect 111 1156 115 1160
rect 135 1157 139 1161
rect 231 1157 235 1161
rect 359 1157 363 1161
rect 487 1157 491 1161
rect 615 1157 619 1161
rect 743 1157 747 1161
rect 871 1157 875 1161
rect 991 1157 995 1161
rect 1119 1157 1123 1161
rect 1247 1157 1251 1161
rect 1767 1156 1771 1160
rect 1807 1156 1811 1160
rect 1935 1157 1939 1161
rect 2039 1157 2043 1161
rect 2159 1157 2163 1161
rect 2287 1157 2291 1161
rect 2423 1157 2427 1161
rect 2567 1157 2571 1161
rect 2703 1157 2707 1161
rect 2839 1157 2843 1161
rect 2975 1157 2979 1161
rect 3111 1157 3115 1161
rect 3247 1157 3251 1161
rect 3367 1157 3371 1161
rect 3463 1156 3467 1160
rect 111 1108 115 1112
rect 247 1107 251 1111
rect 367 1107 371 1111
rect 495 1107 499 1111
rect 623 1107 627 1111
rect 759 1107 763 1111
rect 887 1107 891 1111
rect 1015 1107 1019 1111
rect 1143 1107 1147 1111
rect 1271 1107 1275 1111
rect 1399 1107 1403 1111
rect 1767 1108 1771 1112
rect 1807 1104 1811 1108
rect 1943 1103 1947 1107
rect 2063 1103 2067 1107
rect 2191 1103 2195 1107
rect 2319 1103 2323 1107
rect 2455 1103 2459 1107
rect 2599 1103 2603 1107
rect 2751 1103 2755 1107
rect 2903 1103 2907 1107
rect 3063 1103 3067 1107
rect 3223 1103 3227 1107
rect 3367 1103 3371 1107
rect 3463 1104 3467 1108
rect 111 1091 115 1095
rect 247 1088 251 1092
rect 367 1088 371 1092
rect 495 1088 499 1092
rect 623 1088 627 1092
rect 759 1088 763 1092
rect 887 1088 891 1092
rect 1015 1088 1019 1092
rect 1143 1088 1147 1092
rect 1271 1088 1275 1092
rect 1399 1088 1403 1092
rect 1767 1091 1771 1095
rect 1807 1087 1811 1091
rect 1943 1084 1947 1088
rect 2063 1084 2067 1088
rect 2191 1084 2195 1088
rect 2319 1084 2323 1088
rect 2455 1084 2459 1088
rect 2599 1084 2603 1088
rect 2751 1084 2755 1088
rect 2903 1084 2907 1088
rect 3063 1084 3067 1088
rect 3223 1084 3227 1088
rect 3367 1084 3371 1088
rect 3463 1087 3467 1091
rect 111 1037 115 1041
rect 431 1040 435 1044
rect 543 1040 547 1044
rect 663 1040 667 1044
rect 791 1040 795 1044
rect 919 1040 923 1044
rect 1039 1040 1043 1044
rect 1159 1040 1163 1044
rect 1279 1040 1283 1044
rect 1407 1040 1411 1044
rect 1535 1040 1539 1044
rect 1767 1037 1771 1041
rect 1807 1033 1811 1037
rect 1847 1036 1851 1040
rect 1983 1036 1987 1040
rect 2119 1036 2123 1040
rect 2255 1036 2259 1040
rect 2391 1036 2395 1040
rect 2543 1036 2547 1040
rect 2703 1036 2707 1040
rect 2863 1036 2867 1040
rect 3031 1036 3035 1040
rect 3207 1036 3211 1040
rect 3367 1036 3371 1040
rect 3463 1033 3467 1037
rect 111 1020 115 1024
rect 431 1021 435 1025
rect 543 1021 547 1025
rect 663 1021 667 1025
rect 791 1021 795 1025
rect 919 1021 923 1025
rect 1039 1021 1043 1025
rect 1159 1021 1163 1025
rect 1279 1021 1283 1025
rect 1407 1021 1411 1025
rect 1535 1021 1539 1025
rect 1767 1020 1771 1024
rect 1807 1016 1811 1020
rect 1847 1017 1851 1021
rect 1983 1017 1987 1021
rect 2119 1017 2123 1021
rect 2255 1017 2259 1021
rect 2391 1017 2395 1021
rect 2543 1017 2547 1021
rect 2703 1017 2707 1021
rect 2863 1017 2867 1021
rect 3031 1017 3035 1021
rect 3207 1017 3211 1021
rect 3367 1017 3371 1021
rect 3463 1016 3467 1020
rect 111 968 115 972
rect 567 967 571 971
rect 679 967 683 971
rect 791 967 795 971
rect 911 967 915 971
rect 1031 967 1035 971
rect 1143 967 1147 971
rect 1255 967 1259 971
rect 1359 967 1363 971
rect 1471 967 1475 971
rect 1583 967 1587 971
rect 1671 967 1675 971
rect 1767 968 1771 972
rect 1807 968 1811 972
rect 1831 967 1835 971
rect 1975 967 1979 971
rect 2135 967 2139 971
rect 2295 967 2299 971
rect 2463 967 2467 971
rect 2631 967 2635 971
rect 2807 967 2811 971
rect 2991 967 2995 971
rect 3183 967 3187 971
rect 3367 967 3371 971
rect 3463 968 3467 972
rect 111 951 115 955
rect 567 948 571 952
rect 679 948 683 952
rect 791 948 795 952
rect 911 948 915 952
rect 1031 948 1035 952
rect 1143 948 1147 952
rect 1255 948 1259 952
rect 1359 948 1363 952
rect 1471 948 1475 952
rect 1583 948 1587 952
rect 1671 948 1675 952
rect 1767 951 1771 955
rect 1807 951 1811 955
rect 1831 948 1835 952
rect 1975 948 1979 952
rect 2135 948 2139 952
rect 2295 948 2299 952
rect 2463 948 2467 952
rect 2631 948 2635 952
rect 2807 948 2811 952
rect 2991 948 2995 952
rect 3183 948 3187 952
rect 3367 948 3371 952
rect 3463 951 3467 955
rect 111 897 115 901
rect 415 900 419 904
rect 559 900 563 904
rect 727 900 731 904
rect 911 900 915 904
rect 1119 900 1123 904
rect 1335 900 1339 904
rect 1559 900 1563 904
rect 1767 897 1771 901
rect 1807 901 1811 905
rect 2127 904 2131 908
rect 2215 904 2219 908
rect 2303 904 2307 908
rect 2391 904 2395 908
rect 2479 904 2483 908
rect 2567 904 2571 908
rect 2655 904 2659 908
rect 2743 904 2747 908
rect 2831 904 2835 908
rect 3463 901 3467 905
rect 111 880 115 884
rect 415 881 419 885
rect 559 881 563 885
rect 727 881 731 885
rect 911 881 915 885
rect 1119 881 1123 885
rect 1335 881 1339 885
rect 1559 881 1563 885
rect 1767 880 1771 884
rect 1807 884 1811 888
rect 2127 885 2131 889
rect 2215 885 2219 889
rect 2303 885 2307 889
rect 2391 885 2395 889
rect 2479 885 2483 889
rect 2567 885 2571 889
rect 2655 885 2659 889
rect 2743 885 2747 889
rect 2831 885 2835 889
rect 3463 884 3467 888
rect 111 832 115 836
rect 135 831 139 835
rect 231 831 235 835
rect 359 831 363 835
rect 487 831 491 835
rect 623 831 627 835
rect 751 831 755 835
rect 879 831 883 835
rect 1007 831 1011 835
rect 1135 831 1139 835
rect 1271 831 1275 835
rect 1767 832 1771 836
rect 1807 832 1811 836
rect 2159 831 2163 835
rect 2247 831 2251 835
rect 2335 831 2339 835
rect 2423 831 2427 835
rect 2527 831 2531 835
rect 2639 831 2643 835
rect 2767 831 2771 835
rect 2911 831 2915 835
rect 3063 831 3067 835
rect 3223 831 3227 835
rect 3367 831 3371 835
rect 3463 832 3467 836
rect 111 815 115 819
rect 135 812 139 816
rect 231 812 235 816
rect 359 812 363 816
rect 487 812 491 816
rect 623 812 627 816
rect 751 812 755 816
rect 879 812 883 816
rect 1007 812 1011 816
rect 1135 812 1139 816
rect 1271 812 1275 816
rect 1767 815 1771 819
rect 1807 815 1811 819
rect 2159 812 2163 816
rect 2247 812 2251 816
rect 2335 812 2339 816
rect 2423 812 2427 816
rect 2527 812 2531 816
rect 2639 812 2643 816
rect 2767 812 2771 816
rect 2911 812 2915 816
rect 3063 812 3067 816
rect 3223 812 3227 816
rect 3367 812 3371 816
rect 3463 815 3467 819
rect 111 761 115 765
rect 135 764 139 768
rect 223 764 227 768
rect 343 764 347 768
rect 471 764 475 768
rect 607 764 611 768
rect 743 764 747 768
rect 887 764 891 768
rect 1039 764 1043 768
rect 1191 764 1195 768
rect 1351 764 1355 768
rect 1767 761 1771 765
rect 1807 761 1811 765
rect 2063 764 2067 768
rect 2175 764 2179 768
rect 2295 764 2299 768
rect 2423 764 2427 768
rect 2559 764 2563 768
rect 2711 764 2715 768
rect 2871 764 2875 768
rect 3039 764 3043 768
rect 3215 764 3219 768
rect 3367 764 3371 768
rect 3463 761 3467 765
rect 111 744 115 748
rect 135 745 139 749
rect 223 745 227 749
rect 343 745 347 749
rect 471 745 475 749
rect 607 745 611 749
rect 743 745 747 749
rect 887 745 891 749
rect 1039 745 1043 749
rect 1191 745 1195 749
rect 1351 745 1355 749
rect 1767 744 1771 748
rect 1807 744 1811 748
rect 2063 745 2067 749
rect 2175 745 2179 749
rect 2295 745 2299 749
rect 2423 745 2427 749
rect 2559 745 2563 749
rect 2711 745 2715 749
rect 2871 745 2875 749
rect 3039 745 3043 749
rect 3215 745 3219 749
rect 3367 745 3371 749
rect 3463 744 3467 748
rect 111 696 115 700
rect 167 695 171 699
rect 295 695 299 699
rect 431 695 435 699
rect 575 695 579 699
rect 727 695 731 699
rect 879 695 883 699
rect 1031 695 1035 699
rect 1183 695 1187 699
rect 1343 695 1347 699
rect 1503 695 1507 699
rect 1767 696 1771 700
rect 1807 700 1811 704
rect 1927 699 1931 703
rect 2071 699 2075 703
rect 2231 699 2235 703
rect 2391 699 2395 703
rect 2551 699 2555 703
rect 2703 699 2707 703
rect 2847 699 2851 703
rect 2983 699 2987 703
rect 3119 699 3123 703
rect 3255 699 3259 703
rect 3367 699 3371 703
rect 3463 700 3467 704
rect 111 679 115 683
rect 167 676 171 680
rect 295 676 299 680
rect 431 676 435 680
rect 575 676 579 680
rect 727 676 731 680
rect 879 676 883 680
rect 1031 676 1035 680
rect 1183 676 1187 680
rect 1343 676 1347 680
rect 1503 676 1507 680
rect 1767 679 1771 683
rect 1807 683 1811 687
rect 1927 680 1931 684
rect 2071 680 2075 684
rect 2231 680 2235 684
rect 2391 680 2395 684
rect 2551 680 2555 684
rect 2703 680 2707 684
rect 2847 680 2851 684
rect 2983 680 2987 684
rect 3119 680 3123 684
rect 3255 680 3259 684
rect 3367 680 3371 684
rect 3463 683 3467 687
rect 111 625 115 629
rect 455 628 459 632
rect 559 628 563 632
rect 679 628 683 632
rect 799 628 803 632
rect 927 628 931 632
rect 1055 628 1059 632
rect 1183 628 1187 632
rect 1311 628 1315 632
rect 1447 628 1451 632
rect 1583 628 1587 632
rect 1767 625 1771 629
rect 1807 625 1811 629
rect 1831 628 1835 632
rect 1967 628 1971 632
rect 2135 628 2139 632
rect 2311 628 2315 632
rect 2487 628 2491 632
rect 2655 628 2659 632
rect 2815 628 2819 632
rect 2959 628 2963 632
rect 3103 628 3107 632
rect 3247 628 3251 632
rect 3367 628 3371 632
rect 3463 625 3467 629
rect 111 608 115 612
rect 455 609 459 613
rect 559 609 563 613
rect 679 609 683 613
rect 799 609 803 613
rect 927 609 931 613
rect 1055 609 1059 613
rect 1183 609 1187 613
rect 1311 609 1315 613
rect 1447 609 1451 613
rect 1583 609 1587 613
rect 1767 608 1771 612
rect 1807 608 1811 612
rect 1831 609 1835 613
rect 1967 609 1971 613
rect 2135 609 2139 613
rect 2311 609 2315 613
rect 2487 609 2491 613
rect 2655 609 2659 613
rect 2815 609 2819 613
rect 2959 609 2963 613
rect 3103 609 3107 613
rect 3247 609 3251 613
rect 3367 609 3371 613
rect 3463 608 3467 612
rect 1807 564 1811 568
rect 1831 563 1835 567
rect 1967 563 1971 567
rect 2127 563 2131 567
rect 2287 563 2291 567
rect 2455 563 2459 567
rect 2623 563 2627 567
rect 2799 563 2803 567
rect 2983 563 2987 567
rect 3167 563 3171 567
rect 3359 563 3363 567
rect 3463 564 3467 568
rect 111 556 115 560
rect 599 555 603 559
rect 703 555 707 559
rect 815 555 819 559
rect 927 555 931 559
rect 1039 555 1043 559
rect 1151 555 1155 559
rect 1255 555 1259 559
rect 1359 555 1363 559
rect 1471 555 1475 559
rect 1583 555 1587 559
rect 1671 555 1675 559
rect 1767 556 1771 560
rect 1807 547 1811 551
rect 1831 544 1835 548
rect 111 539 115 543
rect 1967 544 1971 548
rect 2127 544 2131 548
rect 2287 544 2291 548
rect 2455 544 2459 548
rect 2623 544 2627 548
rect 2799 544 2803 548
rect 2983 544 2987 548
rect 3167 544 3171 548
rect 3359 544 3363 548
rect 3463 547 3467 551
rect 599 536 603 540
rect 703 536 707 540
rect 815 536 819 540
rect 927 536 931 540
rect 1039 536 1043 540
rect 1151 536 1155 540
rect 1255 536 1259 540
rect 1359 536 1363 540
rect 1471 536 1475 540
rect 1583 536 1587 540
rect 1671 536 1675 540
rect 1767 539 1771 543
rect 111 489 115 493
rect 303 492 307 496
rect 431 492 435 496
rect 567 492 571 496
rect 703 492 707 496
rect 847 492 851 496
rect 983 492 987 496
rect 1111 492 1115 496
rect 1231 492 1235 496
rect 1351 492 1355 496
rect 1463 492 1467 496
rect 1575 492 1579 496
rect 1671 492 1675 496
rect 1767 489 1771 493
rect 1807 481 1811 485
rect 1831 484 1835 488
rect 1967 484 1971 488
rect 2127 484 2131 488
rect 2295 484 2299 488
rect 2479 484 2483 488
rect 2679 484 2683 488
rect 2887 484 2891 488
rect 3111 484 3115 488
rect 3335 484 3339 488
rect 3463 481 3467 485
rect 111 472 115 476
rect 303 473 307 477
rect 431 473 435 477
rect 567 473 571 477
rect 703 473 707 477
rect 847 473 851 477
rect 983 473 987 477
rect 1111 473 1115 477
rect 1231 473 1235 477
rect 1351 473 1355 477
rect 1463 473 1467 477
rect 1575 473 1579 477
rect 1671 473 1675 477
rect 1767 472 1771 476
rect 1807 464 1811 468
rect 1831 465 1835 469
rect 1967 465 1971 469
rect 2127 465 2131 469
rect 2295 465 2299 469
rect 2479 465 2483 469
rect 2679 465 2683 469
rect 2887 465 2891 469
rect 3111 465 3115 469
rect 3335 465 3339 469
rect 3463 464 3467 468
rect 111 420 115 424
rect 135 419 139 423
rect 255 419 259 423
rect 415 419 419 423
rect 583 419 587 423
rect 743 419 747 423
rect 903 419 907 423
rect 1047 419 1051 423
rect 1183 419 1187 423
rect 1311 419 1315 423
rect 1439 419 1443 423
rect 1567 419 1571 423
rect 1671 419 1675 423
rect 1767 420 1771 424
rect 1807 420 1811 424
rect 1831 419 1835 423
rect 1959 419 1963 423
rect 2111 419 2115 423
rect 2271 419 2275 423
rect 2455 419 2459 423
rect 2655 419 2659 423
rect 2871 419 2875 423
rect 3103 419 3107 423
rect 3335 419 3339 423
rect 3463 420 3467 424
rect 111 403 115 407
rect 135 400 139 404
rect 255 400 259 404
rect 415 400 419 404
rect 583 400 587 404
rect 743 400 747 404
rect 903 400 907 404
rect 1047 400 1051 404
rect 1183 400 1187 404
rect 1311 400 1315 404
rect 1439 400 1443 404
rect 1567 400 1571 404
rect 1671 400 1675 404
rect 1767 403 1771 407
rect 1807 403 1811 407
rect 1831 400 1835 404
rect 1959 400 1963 404
rect 2111 400 2115 404
rect 2271 400 2275 404
rect 2455 400 2459 404
rect 2655 400 2659 404
rect 2871 400 2875 404
rect 3103 400 3107 404
rect 3335 400 3339 404
rect 3463 403 3467 407
rect 111 349 115 353
rect 135 352 139 356
rect 223 352 227 356
rect 343 352 347 356
rect 471 352 475 356
rect 599 352 603 356
rect 719 352 723 356
rect 839 352 843 356
rect 959 352 963 356
rect 1079 352 1083 356
rect 1207 352 1211 356
rect 1767 349 1771 353
rect 1807 349 1811 353
rect 1927 352 1931 356
rect 2039 352 2043 356
rect 2159 352 2163 356
rect 2287 352 2291 356
rect 2423 352 2427 356
rect 2583 352 2587 356
rect 2759 352 2763 356
rect 2951 352 2955 356
rect 3151 352 3155 356
rect 3359 352 3363 356
rect 3463 349 3467 353
rect 111 332 115 336
rect 135 333 139 337
rect 223 333 227 337
rect 343 333 347 337
rect 471 333 475 337
rect 599 333 603 337
rect 719 333 723 337
rect 839 333 843 337
rect 959 333 963 337
rect 1079 333 1083 337
rect 1207 333 1211 337
rect 1767 332 1771 336
rect 1807 332 1811 336
rect 1927 333 1931 337
rect 2039 333 2043 337
rect 2159 333 2163 337
rect 2287 333 2291 337
rect 2423 333 2427 337
rect 2583 333 2587 337
rect 2759 333 2763 337
rect 2951 333 2955 337
rect 3151 333 3155 337
rect 3359 333 3363 337
rect 3463 332 3467 336
rect 111 284 115 288
rect 263 283 267 287
rect 375 283 379 287
rect 487 283 491 287
rect 599 283 603 287
rect 711 283 715 287
rect 815 283 819 287
rect 919 283 923 287
rect 1023 283 1027 287
rect 1127 283 1131 287
rect 1239 283 1243 287
rect 1767 284 1771 288
rect 1807 288 1811 292
rect 2223 287 2227 291
rect 2311 287 2315 291
rect 2399 287 2403 291
rect 2487 287 2491 291
rect 2575 287 2579 291
rect 2679 287 2683 291
rect 2799 287 2803 291
rect 2927 287 2931 291
rect 3071 287 3075 291
rect 3223 287 3227 291
rect 3367 287 3371 291
rect 3463 288 3467 292
rect 111 267 115 271
rect 263 264 267 268
rect 375 264 379 268
rect 487 264 491 268
rect 599 264 603 268
rect 711 264 715 268
rect 815 264 819 268
rect 919 264 923 268
rect 1023 264 1027 268
rect 1127 264 1131 268
rect 1239 264 1243 268
rect 1767 267 1771 271
rect 1807 271 1811 275
rect 2223 268 2227 272
rect 2311 268 2315 272
rect 2399 268 2403 272
rect 2487 268 2491 272
rect 2575 268 2579 272
rect 2679 268 2683 272
rect 2799 268 2803 272
rect 2927 268 2931 272
rect 3071 268 3075 272
rect 3223 268 3227 272
rect 3367 268 3371 272
rect 3463 271 3467 275
rect 111 213 115 217
rect 447 216 451 220
rect 535 216 539 220
rect 623 216 627 220
rect 711 216 715 220
rect 807 216 811 220
rect 903 216 907 220
rect 999 216 1003 220
rect 1103 216 1107 220
rect 1207 216 1211 220
rect 1311 216 1315 220
rect 1767 213 1771 217
rect 1807 213 1811 217
rect 2143 216 2147 220
rect 2263 216 2267 220
rect 2383 216 2387 220
rect 2511 216 2515 220
rect 2639 216 2643 220
rect 2767 216 2771 220
rect 2895 216 2899 220
rect 3015 216 3019 220
rect 3135 216 3139 220
rect 3263 216 3267 220
rect 3367 216 3371 220
rect 3463 213 3467 217
rect 111 196 115 200
rect 447 197 451 201
rect 535 197 539 201
rect 623 197 627 201
rect 711 197 715 201
rect 807 197 811 201
rect 903 197 907 201
rect 999 197 1003 201
rect 1103 197 1107 201
rect 1207 197 1211 201
rect 1311 197 1315 201
rect 1767 196 1771 200
rect 1807 196 1811 200
rect 2143 197 2147 201
rect 2263 197 2267 201
rect 2383 197 2387 201
rect 2511 197 2515 201
rect 2639 197 2643 201
rect 2767 197 2771 201
rect 2895 197 2899 201
rect 3015 197 3019 201
rect 3135 197 3139 201
rect 3263 197 3267 201
rect 3367 197 3371 201
rect 3463 196 3467 200
rect 111 124 115 128
rect 263 123 267 127
rect 351 123 355 127
rect 439 123 443 127
rect 527 123 531 127
rect 615 123 619 127
rect 703 123 707 127
rect 791 123 795 127
rect 879 123 883 127
rect 967 123 971 127
rect 1055 123 1059 127
rect 1143 123 1147 127
rect 1231 123 1235 127
rect 1319 123 1323 127
rect 1407 123 1411 127
rect 1495 123 1499 127
rect 1583 123 1587 127
rect 1671 123 1675 127
rect 1767 124 1771 128
rect 1807 128 1811 132
rect 1831 127 1835 131
rect 1919 127 1923 131
rect 2007 127 2011 131
rect 2095 127 2099 131
rect 2183 127 2187 131
rect 2295 127 2299 131
rect 2407 127 2411 131
rect 2511 127 2515 131
rect 2615 127 2619 131
rect 2719 127 2723 131
rect 2815 127 2819 131
rect 2911 127 2915 131
rect 3007 127 3011 131
rect 3103 127 3107 131
rect 3191 127 3195 131
rect 3279 127 3283 131
rect 3367 127 3371 131
rect 3463 128 3467 132
rect 111 107 115 111
rect 263 104 267 108
rect 351 104 355 108
rect 439 104 443 108
rect 527 104 531 108
rect 615 104 619 108
rect 703 104 707 108
rect 791 104 795 108
rect 879 104 883 108
rect 967 104 971 108
rect 1055 104 1059 108
rect 1143 104 1147 108
rect 1231 104 1235 108
rect 1319 104 1323 108
rect 1407 104 1411 108
rect 1495 104 1499 108
rect 1583 104 1587 108
rect 1671 104 1675 108
rect 1767 107 1771 111
rect 1807 111 1811 115
rect 1831 108 1835 112
rect 1919 108 1923 112
rect 2007 108 2011 112
rect 2095 108 2099 112
rect 2183 108 2187 112
rect 2295 108 2299 112
rect 2407 108 2411 112
rect 2511 108 2515 112
rect 2615 108 2619 112
rect 2719 108 2723 112
rect 2815 108 2819 112
rect 2911 108 2915 112
rect 3007 108 3011 112
rect 3103 108 3107 112
rect 3191 108 3195 112
rect 3279 108 3283 112
rect 3367 108 3371 112
rect 3463 111 3467 115
<< m3 >>
rect 111 3506 115 3507
rect 111 3501 115 3502
rect 135 3506 139 3507
rect 135 3501 139 3502
rect 271 3506 275 3507
rect 271 3501 275 3502
rect 439 3506 443 3507
rect 439 3501 443 3502
rect 615 3506 619 3507
rect 615 3501 619 3502
rect 791 3506 795 3507
rect 791 3501 795 3502
rect 959 3506 963 3507
rect 959 3501 963 3502
rect 1119 3506 1123 3507
rect 1119 3501 1123 3502
rect 1263 3506 1267 3507
rect 1263 3501 1267 3502
rect 1407 3506 1411 3507
rect 1407 3501 1411 3502
rect 1551 3506 1555 3507
rect 1551 3501 1555 3502
rect 1671 3506 1675 3507
rect 1671 3501 1675 3502
rect 1767 3506 1771 3507
rect 1767 3501 1771 3502
rect 112 3485 114 3501
rect 110 3484 116 3485
rect 136 3484 138 3501
rect 272 3484 274 3501
rect 440 3484 442 3501
rect 616 3484 618 3501
rect 792 3484 794 3501
rect 960 3484 962 3501
rect 1120 3484 1122 3501
rect 1264 3484 1266 3501
rect 1408 3484 1410 3501
rect 1552 3484 1554 3501
rect 1672 3484 1674 3501
rect 1768 3485 1770 3501
rect 1807 3494 1811 3495
rect 1807 3489 1811 3490
rect 1831 3494 1835 3495
rect 1831 3489 1835 3490
rect 1975 3494 1979 3495
rect 1975 3489 1979 3490
rect 2143 3494 2147 3495
rect 2143 3489 2147 3490
rect 2311 3494 2315 3495
rect 2311 3489 2315 3490
rect 2479 3494 2483 3495
rect 2479 3489 2483 3490
rect 2639 3494 2643 3495
rect 2639 3489 2643 3490
rect 2799 3494 2803 3495
rect 2799 3489 2803 3490
rect 2967 3494 2971 3495
rect 2967 3489 2971 3490
rect 3463 3494 3467 3495
rect 3463 3489 3467 3490
rect 1766 3484 1772 3485
rect 110 3480 111 3484
rect 115 3480 116 3484
rect 110 3479 116 3480
rect 134 3483 140 3484
rect 134 3479 135 3483
rect 139 3479 140 3483
rect 134 3478 140 3479
rect 270 3483 276 3484
rect 270 3479 271 3483
rect 275 3479 276 3483
rect 270 3478 276 3479
rect 438 3483 444 3484
rect 438 3479 439 3483
rect 443 3479 444 3483
rect 438 3478 444 3479
rect 614 3483 620 3484
rect 614 3479 615 3483
rect 619 3479 620 3483
rect 614 3478 620 3479
rect 790 3483 796 3484
rect 790 3479 791 3483
rect 795 3479 796 3483
rect 790 3478 796 3479
rect 958 3483 964 3484
rect 958 3479 959 3483
rect 963 3479 964 3483
rect 958 3478 964 3479
rect 1118 3483 1124 3484
rect 1118 3479 1119 3483
rect 1123 3479 1124 3483
rect 1118 3478 1124 3479
rect 1262 3483 1268 3484
rect 1262 3479 1263 3483
rect 1267 3479 1268 3483
rect 1262 3478 1268 3479
rect 1406 3483 1412 3484
rect 1406 3479 1407 3483
rect 1411 3479 1412 3483
rect 1406 3478 1412 3479
rect 1550 3483 1556 3484
rect 1550 3479 1551 3483
rect 1555 3479 1556 3483
rect 1550 3478 1556 3479
rect 1670 3483 1676 3484
rect 1670 3479 1671 3483
rect 1675 3479 1676 3483
rect 1766 3480 1767 3484
rect 1771 3480 1772 3484
rect 1766 3479 1772 3480
rect 1670 3478 1676 3479
rect 1808 3473 1810 3489
rect 1806 3472 1812 3473
rect 1832 3472 1834 3489
rect 1976 3472 1978 3489
rect 2144 3472 2146 3489
rect 2312 3472 2314 3489
rect 2480 3472 2482 3489
rect 2640 3472 2642 3489
rect 2800 3472 2802 3489
rect 2968 3472 2970 3489
rect 3464 3473 3466 3489
rect 3462 3472 3468 3473
rect 1806 3468 1807 3472
rect 1811 3468 1812 3472
rect 110 3467 116 3468
rect 110 3463 111 3467
rect 115 3463 116 3467
rect 1766 3467 1772 3468
rect 1806 3467 1812 3468
rect 1830 3471 1836 3472
rect 1830 3467 1831 3471
rect 1835 3467 1836 3471
rect 110 3462 116 3463
rect 134 3464 140 3465
rect 112 3439 114 3462
rect 134 3460 135 3464
rect 139 3460 140 3464
rect 134 3459 140 3460
rect 270 3464 276 3465
rect 270 3460 271 3464
rect 275 3460 276 3464
rect 270 3459 276 3460
rect 438 3464 444 3465
rect 438 3460 439 3464
rect 443 3460 444 3464
rect 438 3459 444 3460
rect 614 3464 620 3465
rect 614 3460 615 3464
rect 619 3460 620 3464
rect 614 3459 620 3460
rect 790 3464 796 3465
rect 790 3460 791 3464
rect 795 3460 796 3464
rect 790 3459 796 3460
rect 958 3464 964 3465
rect 958 3460 959 3464
rect 963 3460 964 3464
rect 958 3459 964 3460
rect 1118 3464 1124 3465
rect 1118 3460 1119 3464
rect 1123 3460 1124 3464
rect 1118 3459 1124 3460
rect 1262 3464 1268 3465
rect 1262 3460 1263 3464
rect 1267 3460 1268 3464
rect 1262 3459 1268 3460
rect 1406 3464 1412 3465
rect 1406 3460 1407 3464
rect 1411 3460 1412 3464
rect 1406 3459 1412 3460
rect 1550 3464 1556 3465
rect 1550 3460 1551 3464
rect 1555 3460 1556 3464
rect 1550 3459 1556 3460
rect 1670 3464 1676 3465
rect 1670 3460 1671 3464
rect 1675 3460 1676 3464
rect 1766 3463 1767 3467
rect 1771 3463 1772 3467
rect 1830 3466 1836 3467
rect 1974 3471 1980 3472
rect 1974 3467 1975 3471
rect 1979 3467 1980 3471
rect 1974 3466 1980 3467
rect 2142 3471 2148 3472
rect 2142 3467 2143 3471
rect 2147 3467 2148 3471
rect 2142 3466 2148 3467
rect 2310 3471 2316 3472
rect 2310 3467 2311 3471
rect 2315 3467 2316 3471
rect 2310 3466 2316 3467
rect 2478 3471 2484 3472
rect 2478 3467 2479 3471
rect 2483 3467 2484 3471
rect 2478 3466 2484 3467
rect 2638 3471 2644 3472
rect 2638 3467 2639 3471
rect 2643 3467 2644 3471
rect 2638 3466 2644 3467
rect 2798 3471 2804 3472
rect 2798 3467 2799 3471
rect 2803 3467 2804 3471
rect 2798 3466 2804 3467
rect 2966 3471 2972 3472
rect 2966 3467 2967 3471
rect 2971 3467 2972 3471
rect 3462 3468 3463 3472
rect 3467 3468 3468 3472
rect 3462 3467 3468 3468
rect 2966 3466 2972 3467
rect 1766 3462 1772 3463
rect 1670 3459 1676 3460
rect 136 3439 138 3459
rect 272 3439 274 3459
rect 440 3439 442 3459
rect 616 3439 618 3459
rect 792 3439 794 3459
rect 960 3439 962 3459
rect 1120 3439 1122 3459
rect 1264 3439 1266 3459
rect 1408 3439 1410 3459
rect 1552 3439 1554 3459
rect 1672 3439 1674 3459
rect 1768 3439 1770 3462
rect 1806 3455 1812 3456
rect 1806 3451 1807 3455
rect 1811 3451 1812 3455
rect 3462 3455 3468 3456
rect 1806 3450 1812 3451
rect 1830 3452 1836 3453
rect 111 3438 115 3439
rect 111 3433 115 3434
rect 135 3438 139 3439
rect 135 3433 139 3434
rect 255 3438 259 3439
rect 255 3433 259 3434
rect 271 3438 275 3439
rect 271 3433 275 3434
rect 415 3438 419 3439
rect 415 3433 419 3434
rect 439 3438 443 3439
rect 439 3433 443 3434
rect 575 3438 579 3439
rect 575 3433 579 3434
rect 615 3438 619 3439
rect 615 3433 619 3434
rect 735 3438 739 3439
rect 735 3433 739 3434
rect 791 3438 795 3439
rect 791 3433 795 3434
rect 895 3438 899 3439
rect 895 3433 899 3434
rect 959 3438 963 3439
rect 959 3433 963 3434
rect 1063 3438 1067 3439
rect 1063 3433 1067 3434
rect 1119 3438 1123 3439
rect 1119 3433 1123 3434
rect 1231 3438 1235 3439
rect 1231 3433 1235 3434
rect 1263 3438 1267 3439
rect 1263 3433 1267 3434
rect 1399 3438 1403 3439
rect 1399 3433 1403 3434
rect 1407 3438 1411 3439
rect 1407 3433 1411 3434
rect 1551 3438 1555 3439
rect 1551 3433 1555 3434
rect 1671 3438 1675 3439
rect 1671 3433 1675 3434
rect 1767 3438 1771 3439
rect 1767 3433 1771 3434
rect 112 3414 114 3433
rect 136 3417 138 3433
rect 256 3417 258 3433
rect 416 3417 418 3433
rect 576 3417 578 3433
rect 736 3417 738 3433
rect 896 3417 898 3433
rect 1064 3417 1066 3433
rect 1232 3417 1234 3433
rect 1400 3417 1402 3433
rect 134 3416 140 3417
rect 110 3413 116 3414
rect 110 3409 111 3413
rect 115 3409 116 3413
rect 134 3412 135 3416
rect 139 3412 140 3416
rect 134 3411 140 3412
rect 254 3416 260 3417
rect 254 3412 255 3416
rect 259 3412 260 3416
rect 254 3411 260 3412
rect 414 3416 420 3417
rect 414 3412 415 3416
rect 419 3412 420 3416
rect 414 3411 420 3412
rect 574 3416 580 3417
rect 574 3412 575 3416
rect 579 3412 580 3416
rect 574 3411 580 3412
rect 734 3416 740 3417
rect 734 3412 735 3416
rect 739 3412 740 3416
rect 734 3411 740 3412
rect 894 3416 900 3417
rect 894 3412 895 3416
rect 899 3412 900 3416
rect 894 3411 900 3412
rect 1062 3416 1068 3417
rect 1062 3412 1063 3416
rect 1067 3412 1068 3416
rect 1062 3411 1068 3412
rect 1230 3416 1236 3417
rect 1230 3412 1231 3416
rect 1235 3412 1236 3416
rect 1230 3411 1236 3412
rect 1398 3416 1404 3417
rect 1398 3412 1399 3416
rect 1403 3412 1404 3416
rect 1768 3414 1770 3433
rect 1808 3431 1810 3450
rect 1830 3448 1831 3452
rect 1835 3448 1836 3452
rect 1830 3447 1836 3448
rect 1974 3452 1980 3453
rect 1974 3448 1975 3452
rect 1979 3448 1980 3452
rect 1974 3447 1980 3448
rect 2142 3452 2148 3453
rect 2142 3448 2143 3452
rect 2147 3448 2148 3452
rect 2142 3447 2148 3448
rect 2310 3452 2316 3453
rect 2310 3448 2311 3452
rect 2315 3448 2316 3452
rect 2310 3447 2316 3448
rect 2478 3452 2484 3453
rect 2478 3448 2479 3452
rect 2483 3448 2484 3452
rect 2478 3447 2484 3448
rect 2638 3452 2644 3453
rect 2638 3448 2639 3452
rect 2643 3448 2644 3452
rect 2638 3447 2644 3448
rect 2798 3452 2804 3453
rect 2798 3448 2799 3452
rect 2803 3448 2804 3452
rect 2798 3447 2804 3448
rect 2966 3452 2972 3453
rect 2966 3448 2967 3452
rect 2971 3448 2972 3452
rect 3462 3451 3463 3455
rect 3467 3451 3468 3455
rect 3462 3450 3468 3451
rect 2966 3447 2972 3448
rect 1832 3431 1834 3447
rect 1976 3431 1978 3447
rect 2144 3431 2146 3447
rect 2312 3431 2314 3447
rect 2480 3431 2482 3447
rect 2640 3431 2642 3447
rect 2800 3431 2802 3447
rect 2968 3431 2970 3447
rect 3464 3431 3466 3450
rect 1807 3430 1811 3431
rect 1807 3425 1811 3426
rect 1831 3430 1835 3431
rect 1831 3425 1835 3426
rect 1975 3430 1979 3431
rect 1975 3425 1979 3426
rect 2031 3430 2035 3431
rect 2031 3425 2035 3426
rect 2143 3430 2147 3431
rect 2143 3425 2147 3426
rect 2151 3430 2155 3431
rect 2151 3425 2155 3426
rect 2271 3430 2275 3431
rect 2271 3425 2275 3426
rect 2311 3430 2315 3431
rect 2311 3425 2315 3426
rect 2391 3430 2395 3431
rect 2391 3425 2395 3426
rect 2479 3430 2483 3431
rect 2479 3425 2483 3426
rect 2511 3430 2515 3431
rect 2511 3425 2515 3426
rect 2623 3430 2627 3431
rect 2623 3425 2627 3426
rect 2639 3430 2643 3431
rect 2639 3425 2643 3426
rect 2727 3430 2731 3431
rect 2727 3425 2731 3426
rect 2799 3430 2803 3431
rect 2799 3425 2803 3426
rect 2831 3430 2835 3431
rect 2831 3425 2835 3426
rect 2935 3430 2939 3431
rect 2935 3425 2939 3426
rect 2967 3430 2971 3431
rect 2967 3425 2971 3426
rect 3039 3430 3043 3431
rect 3039 3425 3043 3426
rect 3151 3430 3155 3431
rect 3151 3425 3155 3426
rect 3463 3430 3467 3431
rect 3463 3425 3467 3426
rect 1398 3411 1404 3412
rect 1766 3413 1772 3414
rect 110 3408 116 3409
rect 1766 3409 1767 3413
rect 1771 3409 1772 3413
rect 1766 3408 1772 3409
rect 1808 3406 1810 3425
rect 2032 3409 2034 3425
rect 2152 3409 2154 3425
rect 2272 3409 2274 3425
rect 2392 3409 2394 3425
rect 2512 3409 2514 3425
rect 2624 3409 2626 3425
rect 2728 3409 2730 3425
rect 2832 3409 2834 3425
rect 2936 3409 2938 3425
rect 3040 3409 3042 3425
rect 3152 3409 3154 3425
rect 2030 3408 2036 3409
rect 1806 3405 1812 3406
rect 1806 3401 1807 3405
rect 1811 3401 1812 3405
rect 2030 3404 2031 3408
rect 2035 3404 2036 3408
rect 2030 3403 2036 3404
rect 2150 3408 2156 3409
rect 2150 3404 2151 3408
rect 2155 3404 2156 3408
rect 2150 3403 2156 3404
rect 2270 3408 2276 3409
rect 2270 3404 2271 3408
rect 2275 3404 2276 3408
rect 2270 3403 2276 3404
rect 2390 3408 2396 3409
rect 2390 3404 2391 3408
rect 2395 3404 2396 3408
rect 2390 3403 2396 3404
rect 2510 3408 2516 3409
rect 2510 3404 2511 3408
rect 2515 3404 2516 3408
rect 2510 3403 2516 3404
rect 2622 3408 2628 3409
rect 2622 3404 2623 3408
rect 2627 3404 2628 3408
rect 2622 3403 2628 3404
rect 2726 3408 2732 3409
rect 2726 3404 2727 3408
rect 2731 3404 2732 3408
rect 2726 3403 2732 3404
rect 2830 3408 2836 3409
rect 2830 3404 2831 3408
rect 2835 3404 2836 3408
rect 2830 3403 2836 3404
rect 2934 3408 2940 3409
rect 2934 3404 2935 3408
rect 2939 3404 2940 3408
rect 2934 3403 2940 3404
rect 3038 3408 3044 3409
rect 3038 3404 3039 3408
rect 3043 3404 3044 3408
rect 3038 3403 3044 3404
rect 3150 3408 3156 3409
rect 3150 3404 3151 3408
rect 3155 3404 3156 3408
rect 3464 3406 3466 3425
rect 3150 3403 3156 3404
rect 3462 3405 3468 3406
rect 1806 3400 1812 3401
rect 3462 3401 3463 3405
rect 3467 3401 3468 3405
rect 3462 3400 3468 3401
rect 134 3397 140 3398
rect 110 3396 116 3397
rect 110 3392 111 3396
rect 115 3392 116 3396
rect 134 3393 135 3397
rect 139 3393 140 3397
rect 134 3392 140 3393
rect 254 3397 260 3398
rect 254 3393 255 3397
rect 259 3393 260 3397
rect 254 3392 260 3393
rect 414 3397 420 3398
rect 414 3393 415 3397
rect 419 3393 420 3397
rect 414 3392 420 3393
rect 574 3397 580 3398
rect 574 3393 575 3397
rect 579 3393 580 3397
rect 574 3392 580 3393
rect 734 3397 740 3398
rect 734 3393 735 3397
rect 739 3393 740 3397
rect 734 3392 740 3393
rect 894 3397 900 3398
rect 894 3393 895 3397
rect 899 3393 900 3397
rect 894 3392 900 3393
rect 1062 3397 1068 3398
rect 1062 3393 1063 3397
rect 1067 3393 1068 3397
rect 1062 3392 1068 3393
rect 1230 3397 1236 3398
rect 1230 3393 1231 3397
rect 1235 3393 1236 3397
rect 1230 3392 1236 3393
rect 1398 3397 1404 3398
rect 1398 3393 1399 3397
rect 1403 3393 1404 3397
rect 1398 3392 1404 3393
rect 1766 3396 1772 3397
rect 1766 3392 1767 3396
rect 1771 3392 1772 3396
rect 110 3391 116 3392
rect 112 3367 114 3391
rect 136 3367 138 3392
rect 256 3367 258 3392
rect 416 3367 418 3392
rect 576 3367 578 3392
rect 736 3367 738 3392
rect 896 3367 898 3392
rect 1064 3367 1066 3392
rect 1232 3367 1234 3392
rect 1400 3367 1402 3392
rect 1766 3391 1772 3392
rect 1768 3367 1770 3391
rect 2030 3389 2036 3390
rect 1806 3388 1812 3389
rect 1806 3384 1807 3388
rect 1811 3384 1812 3388
rect 2030 3385 2031 3389
rect 2035 3385 2036 3389
rect 2030 3384 2036 3385
rect 2150 3389 2156 3390
rect 2150 3385 2151 3389
rect 2155 3385 2156 3389
rect 2150 3384 2156 3385
rect 2270 3389 2276 3390
rect 2270 3385 2271 3389
rect 2275 3385 2276 3389
rect 2270 3384 2276 3385
rect 2390 3389 2396 3390
rect 2390 3385 2391 3389
rect 2395 3385 2396 3389
rect 2390 3384 2396 3385
rect 2510 3389 2516 3390
rect 2510 3385 2511 3389
rect 2515 3385 2516 3389
rect 2510 3384 2516 3385
rect 2622 3389 2628 3390
rect 2622 3385 2623 3389
rect 2627 3385 2628 3389
rect 2622 3384 2628 3385
rect 2726 3389 2732 3390
rect 2726 3385 2727 3389
rect 2731 3385 2732 3389
rect 2726 3384 2732 3385
rect 2830 3389 2836 3390
rect 2830 3385 2831 3389
rect 2835 3385 2836 3389
rect 2830 3384 2836 3385
rect 2934 3389 2940 3390
rect 2934 3385 2935 3389
rect 2939 3385 2940 3389
rect 2934 3384 2940 3385
rect 3038 3389 3044 3390
rect 3038 3385 3039 3389
rect 3043 3385 3044 3389
rect 3038 3384 3044 3385
rect 3150 3389 3156 3390
rect 3150 3385 3151 3389
rect 3155 3385 3156 3389
rect 3150 3384 3156 3385
rect 3462 3388 3468 3389
rect 3462 3384 3463 3388
rect 3467 3384 3468 3388
rect 1806 3383 1812 3384
rect 111 3366 115 3367
rect 111 3361 115 3362
rect 135 3366 139 3367
rect 135 3361 139 3362
rect 255 3366 259 3367
rect 255 3361 259 3362
rect 327 3366 331 3367
rect 327 3361 331 3362
rect 415 3366 419 3367
rect 415 3361 419 3362
rect 535 3366 539 3367
rect 535 3361 539 3362
rect 575 3366 579 3367
rect 575 3361 579 3362
rect 735 3366 739 3367
rect 735 3361 739 3362
rect 743 3366 747 3367
rect 743 3361 747 3362
rect 895 3366 899 3367
rect 895 3361 899 3362
rect 935 3366 939 3367
rect 935 3361 939 3362
rect 1063 3366 1067 3367
rect 1063 3361 1067 3362
rect 1119 3366 1123 3367
rect 1119 3361 1123 3362
rect 1231 3366 1235 3367
rect 1231 3361 1235 3362
rect 1295 3366 1299 3367
rect 1295 3361 1299 3362
rect 1399 3366 1403 3367
rect 1399 3361 1403 3362
rect 1463 3366 1467 3367
rect 1463 3361 1467 3362
rect 1639 3366 1643 3367
rect 1639 3361 1643 3362
rect 1767 3366 1771 3367
rect 1808 3363 1810 3383
rect 2032 3363 2034 3384
rect 2152 3363 2154 3384
rect 2272 3363 2274 3384
rect 2392 3363 2394 3384
rect 2512 3363 2514 3384
rect 2624 3363 2626 3384
rect 2728 3363 2730 3384
rect 2832 3363 2834 3384
rect 2936 3363 2938 3384
rect 3040 3363 3042 3384
rect 3152 3363 3154 3384
rect 3462 3383 3468 3384
rect 3464 3363 3466 3383
rect 1767 3361 1771 3362
rect 1807 3362 1811 3363
rect 112 3345 114 3361
rect 110 3344 116 3345
rect 136 3344 138 3361
rect 328 3344 330 3361
rect 536 3344 538 3361
rect 744 3344 746 3361
rect 936 3344 938 3361
rect 1120 3344 1122 3361
rect 1296 3344 1298 3361
rect 1464 3344 1466 3361
rect 1640 3344 1642 3361
rect 1768 3345 1770 3361
rect 1807 3357 1811 3358
rect 2031 3362 2035 3363
rect 2031 3357 2035 3358
rect 2151 3362 2155 3363
rect 2151 3357 2155 3358
rect 2159 3362 2163 3363
rect 2159 3357 2163 3358
rect 2271 3362 2275 3363
rect 2271 3357 2275 3358
rect 2295 3362 2299 3363
rect 2295 3357 2299 3358
rect 2391 3362 2395 3363
rect 2391 3357 2395 3358
rect 2431 3362 2435 3363
rect 2431 3357 2435 3358
rect 2511 3362 2515 3363
rect 2511 3357 2515 3358
rect 2567 3362 2571 3363
rect 2567 3357 2571 3358
rect 2623 3362 2627 3363
rect 2623 3357 2627 3358
rect 2703 3362 2707 3363
rect 2703 3357 2707 3358
rect 2727 3362 2731 3363
rect 2727 3357 2731 3358
rect 2831 3362 2835 3363
rect 2831 3357 2835 3358
rect 2839 3362 2843 3363
rect 2839 3357 2843 3358
rect 2935 3362 2939 3363
rect 2935 3357 2939 3358
rect 2975 3362 2979 3363
rect 2975 3357 2979 3358
rect 3039 3362 3043 3363
rect 3039 3357 3043 3358
rect 3119 3362 3123 3363
rect 3119 3357 3123 3358
rect 3151 3362 3155 3363
rect 3151 3357 3155 3358
rect 3463 3362 3467 3363
rect 3463 3357 3467 3358
rect 1766 3344 1772 3345
rect 110 3340 111 3344
rect 115 3340 116 3344
rect 110 3339 116 3340
rect 134 3343 140 3344
rect 134 3339 135 3343
rect 139 3339 140 3343
rect 134 3338 140 3339
rect 326 3343 332 3344
rect 326 3339 327 3343
rect 331 3339 332 3343
rect 326 3338 332 3339
rect 534 3343 540 3344
rect 534 3339 535 3343
rect 539 3339 540 3343
rect 534 3338 540 3339
rect 742 3343 748 3344
rect 742 3339 743 3343
rect 747 3339 748 3343
rect 742 3338 748 3339
rect 934 3343 940 3344
rect 934 3339 935 3343
rect 939 3339 940 3343
rect 934 3338 940 3339
rect 1118 3343 1124 3344
rect 1118 3339 1119 3343
rect 1123 3339 1124 3343
rect 1118 3338 1124 3339
rect 1294 3343 1300 3344
rect 1294 3339 1295 3343
rect 1299 3339 1300 3343
rect 1294 3338 1300 3339
rect 1462 3343 1468 3344
rect 1462 3339 1463 3343
rect 1467 3339 1468 3343
rect 1462 3338 1468 3339
rect 1638 3343 1644 3344
rect 1638 3339 1639 3343
rect 1643 3339 1644 3343
rect 1766 3340 1767 3344
rect 1771 3340 1772 3344
rect 1808 3341 1810 3357
rect 1766 3339 1772 3340
rect 1806 3340 1812 3341
rect 2160 3340 2162 3357
rect 2296 3340 2298 3357
rect 2432 3340 2434 3357
rect 2568 3340 2570 3357
rect 2704 3340 2706 3357
rect 2840 3340 2842 3357
rect 2976 3340 2978 3357
rect 3120 3340 3122 3357
rect 3464 3341 3466 3357
rect 3462 3340 3468 3341
rect 1638 3338 1644 3339
rect 1806 3336 1807 3340
rect 1811 3336 1812 3340
rect 1806 3335 1812 3336
rect 2158 3339 2164 3340
rect 2158 3335 2159 3339
rect 2163 3335 2164 3339
rect 2158 3334 2164 3335
rect 2294 3339 2300 3340
rect 2294 3335 2295 3339
rect 2299 3335 2300 3339
rect 2294 3334 2300 3335
rect 2430 3339 2436 3340
rect 2430 3335 2431 3339
rect 2435 3335 2436 3339
rect 2430 3334 2436 3335
rect 2566 3339 2572 3340
rect 2566 3335 2567 3339
rect 2571 3335 2572 3339
rect 2566 3334 2572 3335
rect 2702 3339 2708 3340
rect 2702 3335 2703 3339
rect 2707 3335 2708 3339
rect 2702 3334 2708 3335
rect 2838 3339 2844 3340
rect 2838 3335 2839 3339
rect 2843 3335 2844 3339
rect 2838 3334 2844 3335
rect 2974 3339 2980 3340
rect 2974 3335 2975 3339
rect 2979 3335 2980 3339
rect 2974 3334 2980 3335
rect 3118 3339 3124 3340
rect 3118 3335 3119 3339
rect 3123 3335 3124 3339
rect 3462 3336 3463 3340
rect 3467 3336 3468 3340
rect 3462 3335 3468 3336
rect 3118 3334 3124 3335
rect 110 3327 116 3328
rect 110 3323 111 3327
rect 115 3323 116 3327
rect 1766 3327 1772 3328
rect 110 3322 116 3323
rect 134 3324 140 3325
rect 112 3295 114 3322
rect 134 3320 135 3324
rect 139 3320 140 3324
rect 134 3319 140 3320
rect 326 3324 332 3325
rect 326 3320 327 3324
rect 331 3320 332 3324
rect 326 3319 332 3320
rect 534 3324 540 3325
rect 534 3320 535 3324
rect 539 3320 540 3324
rect 534 3319 540 3320
rect 742 3324 748 3325
rect 742 3320 743 3324
rect 747 3320 748 3324
rect 742 3319 748 3320
rect 934 3324 940 3325
rect 934 3320 935 3324
rect 939 3320 940 3324
rect 934 3319 940 3320
rect 1118 3324 1124 3325
rect 1118 3320 1119 3324
rect 1123 3320 1124 3324
rect 1118 3319 1124 3320
rect 1294 3324 1300 3325
rect 1294 3320 1295 3324
rect 1299 3320 1300 3324
rect 1294 3319 1300 3320
rect 1462 3324 1468 3325
rect 1462 3320 1463 3324
rect 1467 3320 1468 3324
rect 1462 3319 1468 3320
rect 1638 3324 1644 3325
rect 1638 3320 1639 3324
rect 1643 3320 1644 3324
rect 1766 3323 1767 3327
rect 1771 3323 1772 3327
rect 1766 3322 1772 3323
rect 1806 3323 1812 3324
rect 1638 3319 1644 3320
rect 136 3295 138 3319
rect 328 3295 330 3319
rect 536 3295 538 3319
rect 744 3295 746 3319
rect 936 3295 938 3319
rect 1120 3295 1122 3319
rect 1296 3295 1298 3319
rect 1464 3295 1466 3319
rect 1640 3295 1642 3319
rect 1768 3295 1770 3322
rect 1806 3319 1807 3323
rect 1811 3319 1812 3323
rect 3462 3323 3468 3324
rect 1806 3318 1812 3319
rect 2158 3320 2164 3321
rect 1808 3299 1810 3318
rect 2158 3316 2159 3320
rect 2163 3316 2164 3320
rect 2158 3315 2164 3316
rect 2294 3320 2300 3321
rect 2294 3316 2295 3320
rect 2299 3316 2300 3320
rect 2294 3315 2300 3316
rect 2430 3320 2436 3321
rect 2430 3316 2431 3320
rect 2435 3316 2436 3320
rect 2430 3315 2436 3316
rect 2566 3320 2572 3321
rect 2566 3316 2567 3320
rect 2571 3316 2572 3320
rect 2566 3315 2572 3316
rect 2702 3320 2708 3321
rect 2702 3316 2703 3320
rect 2707 3316 2708 3320
rect 2702 3315 2708 3316
rect 2838 3320 2844 3321
rect 2838 3316 2839 3320
rect 2843 3316 2844 3320
rect 2838 3315 2844 3316
rect 2974 3320 2980 3321
rect 2974 3316 2975 3320
rect 2979 3316 2980 3320
rect 2974 3315 2980 3316
rect 3118 3320 3124 3321
rect 3118 3316 3119 3320
rect 3123 3316 3124 3320
rect 3462 3319 3463 3323
rect 3467 3319 3468 3323
rect 3462 3318 3468 3319
rect 3118 3315 3124 3316
rect 2160 3299 2162 3315
rect 2296 3299 2298 3315
rect 2432 3299 2434 3315
rect 2568 3299 2570 3315
rect 2704 3299 2706 3315
rect 2840 3299 2842 3315
rect 2976 3299 2978 3315
rect 3120 3299 3122 3315
rect 3464 3299 3466 3318
rect 1807 3298 1811 3299
rect 111 3294 115 3295
rect 111 3289 115 3290
rect 135 3294 139 3295
rect 135 3289 139 3290
rect 279 3294 283 3295
rect 279 3289 283 3290
rect 327 3294 331 3295
rect 327 3289 331 3290
rect 463 3294 467 3295
rect 463 3289 467 3290
rect 535 3294 539 3295
rect 535 3289 539 3290
rect 647 3294 651 3295
rect 647 3289 651 3290
rect 743 3294 747 3295
rect 743 3289 747 3290
rect 831 3294 835 3295
rect 831 3289 835 3290
rect 935 3294 939 3295
rect 935 3289 939 3290
rect 1007 3294 1011 3295
rect 1007 3289 1011 3290
rect 1119 3294 1123 3295
rect 1119 3289 1123 3290
rect 1175 3294 1179 3295
rect 1175 3289 1179 3290
rect 1295 3294 1299 3295
rect 1295 3289 1299 3290
rect 1343 3294 1347 3295
rect 1343 3289 1347 3290
rect 1463 3294 1467 3295
rect 1463 3289 1467 3290
rect 1503 3294 1507 3295
rect 1503 3289 1507 3290
rect 1639 3294 1643 3295
rect 1639 3289 1643 3290
rect 1671 3294 1675 3295
rect 1671 3289 1675 3290
rect 1767 3294 1771 3295
rect 1807 3293 1811 3294
rect 2087 3298 2091 3299
rect 2087 3293 2091 3294
rect 2159 3298 2163 3299
rect 2159 3293 2163 3294
rect 2239 3298 2243 3299
rect 2239 3293 2243 3294
rect 2295 3298 2299 3299
rect 2295 3293 2299 3294
rect 2399 3298 2403 3299
rect 2399 3293 2403 3294
rect 2431 3298 2435 3299
rect 2431 3293 2435 3294
rect 2559 3298 2563 3299
rect 2559 3293 2563 3294
rect 2567 3298 2571 3299
rect 2567 3293 2571 3294
rect 2703 3298 2707 3299
rect 2703 3293 2707 3294
rect 2719 3298 2723 3299
rect 2719 3293 2723 3294
rect 2839 3298 2843 3299
rect 2839 3293 2843 3294
rect 2879 3298 2883 3299
rect 2879 3293 2883 3294
rect 2975 3298 2979 3299
rect 2975 3293 2979 3294
rect 3039 3298 3043 3299
rect 3039 3293 3043 3294
rect 3119 3298 3123 3299
rect 3119 3293 3123 3294
rect 3199 3298 3203 3299
rect 3199 3293 3203 3294
rect 3463 3298 3467 3299
rect 3463 3293 3467 3294
rect 1767 3289 1771 3290
rect 112 3270 114 3289
rect 136 3273 138 3289
rect 280 3273 282 3289
rect 464 3273 466 3289
rect 648 3273 650 3289
rect 832 3273 834 3289
rect 1008 3273 1010 3289
rect 1176 3273 1178 3289
rect 1344 3273 1346 3289
rect 1504 3273 1506 3289
rect 1672 3273 1674 3289
rect 134 3272 140 3273
rect 110 3269 116 3270
rect 110 3265 111 3269
rect 115 3265 116 3269
rect 134 3268 135 3272
rect 139 3268 140 3272
rect 134 3267 140 3268
rect 278 3272 284 3273
rect 278 3268 279 3272
rect 283 3268 284 3272
rect 278 3267 284 3268
rect 462 3272 468 3273
rect 462 3268 463 3272
rect 467 3268 468 3272
rect 462 3267 468 3268
rect 646 3272 652 3273
rect 646 3268 647 3272
rect 651 3268 652 3272
rect 646 3267 652 3268
rect 830 3272 836 3273
rect 830 3268 831 3272
rect 835 3268 836 3272
rect 830 3267 836 3268
rect 1006 3272 1012 3273
rect 1006 3268 1007 3272
rect 1011 3268 1012 3272
rect 1006 3267 1012 3268
rect 1174 3272 1180 3273
rect 1174 3268 1175 3272
rect 1179 3268 1180 3272
rect 1174 3267 1180 3268
rect 1342 3272 1348 3273
rect 1342 3268 1343 3272
rect 1347 3268 1348 3272
rect 1342 3267 1348 3268
rect 1502 3272 1508 3273
rect 1502 3268 1503 3272
rect 1507 3268 1508 3272
rect 1502 3267 1508 3268
rect 1670 3272 1676 3273
rect 1670 3268 1671 3272
rect 1675 3268 1676 3272
rect 1768 3270 1770 3289
rect 1808 3274 1810 3293
rect 2088 3277 2090 3293
rect 2240 3277 2242 3293
rect 2400 3277 2402 3293
rect 2560 3277 2562 3293
rect 2720 3277 2722 3293
rect 2880 3277 2882 3293
rect 3040 3277 3042 3293
rect 3200 3277 3202 3293
rect 2086 3276 2092 3277
rect 1806 3273 1812 3274
rect 1670 3267 1676 3268
rect 1766 3269 1772 3270
rect 110 3264 116 3265
rect 1766 3265 1767 3269
rect 1771 3265 1772 3269
rect 1806 3269 1807 3273
rect 1811 3269 1812 3273
rect 2086 3272 2087 3276
rect 2091 3272 2092 3276
rect 2086 3271 2092 3272
rect 2238 3276 2244 3277
rect 2238 3272 2239 3276
rect 2243 3272 2244 3276
rect 2238 3271 2244 3272
rect 2398 3276 2404 3277
rect 2398 3272 2399 3276
rect 2403 3272 2404 3276
rect 2398 3271 2404 3272
rect 2558 3276 2564 3277
rect 2558 3272 2559 3276
rect 2563 3272 2564 3276
rect 2558 3271 2564 3272
rect 2718 3276 2724 3277
rect 2718 3272 2719 3276
rect 2723 3272 2724 3276
rect 2718 3271 2724 3272
rect 2878 3276 2884 3277
rect 2878 3272 2879 3276
rect 2883 3272 2884 3276
rect 2878 3271 2884 3272
rect 3038 3276 3044 3277
rect 3038 3272 3039 3276
rect 3043 3272 3044 3276
rect 3038 3271 3044 3272
rect 3198 3276 3204 3277
rect 3198 3272 3199 3276
rect 3203 3272 3204 3276
rect 3464 3274 3466 3293
rect 3198 3271 3204 3272
rect 3462 3273 3468 3274
rect 1806 3268 1812 3269
rect 3462 3269 3463 3273
rect 3467 3269 3468 3273
rect 3462 3268 3468 3269
rect 1766 3264 1772 3265
rect 2086 3257 2092 3258
rect 1806 3256 1812 3257
rect 134 3253 140 3254
rect 110 3252 116 3253
rect 110 3248 111 3252
rect 115 3248 116 3252
rect 134 3249 135 3253
rect 139 3249 140 3253
rect 134 3248 140 3249
rect 278 3253 284 3254
rect 278 3249 279 3253
rect 283 3249 284 3253
rect 278 3248 284 3249
rect 462 3253 468 3254
rect 462 3249 463 3253
rect 467 3249 468 3253
rect 462 3248 468 3249
rect 646 3253 652 3254
rect 646 3249 647 3253
rect 651 3249 652 3253
rect 646 3248 652 3249
rect 830 3253 836 3254
rect 830 3249 831 3253
rect 835 3249 836 3253
rect 830 3248 836 3249
rect 1006 3253 1012 3254
rect 1006 3249 1007 3253
rect 1011 3249 1012 3253
rect 1006 3248 1012 3249
rect 1174 3253 1180 3254
rect 1174 3249 1175 3253
rect 1179 3249 1180 3253
rect 1174 3248 1180 3249
rect 1342 3253 1348 3254
rect 1342 3249 1343 3253
rect 1347 3249 1348 3253
rect 1342 3248 1348 3249
rect 1502 3253 1508 3254
rect 1502 3249 1503 3253
rect 1507 3249 1508 3253
rect 1502 3248 1508 3249
rect 1670 3253 1676 3254
rect 1670 3249 1671 3253
rect 1675 3249 1676 3253
rect 1670 3248 1676 3249
rect 1766 3252 1772 3253
rect 1766 3248 1767 3252
rect 1771 3248 1772 3252
rect 1806 3252 1807 3256
rect 1811 3252 1812 3256
rect 2086 3253 2087 3257
rect 2091 3253 2092 3257
rect 2086 3252 2092 3253
rect 2238 3257 2244 3258
rect 2238 3253 2239 3257
rect 2243 3253 2244 3257
rect 2238 3252 2244 3253
rect 2398 3257 2404 3258
rect 2398 3253 2399 3257
rect 2403 3253 2404 3257
rect 2398 3252 2404 3253
rect 2558 3257 2564 3258
rect 2558 3253 2559 3257
rect 2563 3253 2564 3257
rect 2558 3252 2564 3253
rect 2718 3257 2724 3258
rect 2718 3253 2719 3257
rect 2723 3253 2724 3257
rect 2718 3252 2724 3253
rect 2878 3257 2884 3258
rect 2878 3253 2879 3257
rect 2883 3253 2884 3257
rect 2878 3252 2884 3253
rect 3038 3257 3044 3258
rect 3038 3253 3039 3257
rect 3043 3253 3044 3257
rect 3038 3252 3044 3253
rect 3198 3257 3204 3258
rect 3198 3253 3199 3257
rect 3203 3253 3204 3257
rect 3198 3252 3204 3253
rect 3462 3256 3468 3257
rect 3462 3252 3463 3256
rect 3467 3252 3468 3256
rect 1806 3251 1812 3252
rect 110 3247 116 3248
rect 112 3223 114 3247
rect 136 3223 138 3248
rect 280 3223 282 3248
rect 464 3223 466 3248
rect 648 3223 650 3248
rect 832 3223 834 3248
rect 1008 3223 1010 3248
rect 1176 3223 1178 3248
rect 1344 3223 1346 3248
rect 1504 3223 1506 3248
rect 1672 3223 1674 3248
rect 1766 3247 1772 3248
rect 1768 3223 1770 3247
rect 1808 3231 1810 3251
rect 2088 3231 2090 3252
rect 2240 3231 2242 3252
rect 2400 3231 2402 3252
rect 2560 3231 2562 3252
rect 2720 3231 2722 3252
rect 2880 3231 2882 3252
rect 3040 3231 3042 3252
rect 3200 3231 3202 3252
rect 3462 3251 3468 3252
rect 3464 3231 3466 3251
rect 1807 3230 1811 3231
rect 1807 3225 1811 3226
rect 1911 3230 1915 3231
rect 1911 3225 1915 3226
rect 2047 3230 2051 3231
rect 2047 3225 2051 3226
rect 2087 3230 2091 3231
rect 2087 3225 2091 3226
rect 2199 3230 2203 3231
rect 2199 3225 2203 3226
rect 2239 3230 2243 3231
rect 2239 3225 2243 3226
rect 2359 3230 2363 3231
rect 2359 3225 2363 3226
rect 2399 3230 2403 3231
rect 2399 3225 2403 3226
rect 2527 3230 2531 3231
rect 2527 3225 2531 3226
rect 2559 3230 2563 3231
rect 2559 3225 2563 3226
rect 2687 3230 2691 3231
rect 2687 3225 2691 3226
rect 2719 3230 2723 3231
rect 2719 3225 2723 3226
rect 2847 3230 2851 3231
rect 2847 3225 2851 3226
rect 2879 3230 2883 3231
rect 2879 3225 2883 3226
rect 3007 3230 3011 3231
rect 3007 3225 3011 3226
rect 3039 3230 3043 3231
rect 3039 3225 3043 3226
rect 3167 3230 3171 3231
rect 3167 3225 3171 3226
rect 3199 3230 3203 3231
rect 3199 3225 3203 3226
rect 3335 3230 3339 3231
rect 3335 3225 3339 3226
rect 3463 3230 3467 3231
rect 3463 3225 3467 3226
rect 111 3222 115 3223
rect 111 3217 115 3218
rect 135 3222 139 3223
rect 135 3217 139 3218
rect 183 3222 187 3223
rect 183 3217 187 3218
rect 279 3222 283 3223
rect 279 3217 283 3218
rect 327 3222 331 3223
rect 327 3217 331 3218
rect 463 3222 467 3223
rect 463 3217 467 3218
rect 487 3222 491 3223
rect 487 3217 491 3218
rect 647 3222 651 3223
rect 647 3217 651 3218
rect 807 3222 811 3223
rect 807 3217 811 3218
rect 831 3222 835 3223
rect 831 3217 835 3218
rect 967 3222 971 3223
rect 967 3217 971 3218
rect 1007 3222 1011 3223
rect 1007 3217 1011 3218
rect 1135 3222 1139 3223
rect 1135 3217 1139 3218
rect 1175 3222 1179 3223
rect 1175 3217 1179 3218
rect 1303 3222 1307 3223
rect 1303 3217 1307 3218
rect 1343 3222 1347 3223
rect 1343 3217 1347 3218
rect 1471 3222 1475 3223
rect 1471 3217 1475 3218
rect 1503 3222 1507 3223
rect 1503 3217 1507 3218
rect 1671 3222 1675 3223
rect 1671 3217 1675 3218
rect 1767 3222 1771 3223
rect 1767 3217 1771 3218
rect 112 3201 114 3217
rect 110 3200 116 3201
rect 184 3200 186 3217
rect 328 3200 330 3217
rect 488 3200 490 3217
rect 648 3200 650 3217
rect 808 3200 810 3217
rect 968 3200 970 3217
rect 1136 3200 1138 3217
rect 1304 3200 1306 3217
rect 1472 3200 1474 3217
rect 1768 3201 1770 3217
rect 1808 3209 1810 3225
rect 1806 3208 1812 3209
rect 1912 3208 1914 3225
rect 2048 3208 2050 3225
rect 2200 3208 2202 3225
rect 2360 3208 2362 3225
rect 2528 3208 2530 3225
rect 2688 3208 2690 3225
rect 2848 3208 2850 3225
rect 3008 3208 3010 3225
rect 3168 3208 3170 3225
rect 3336 3208 3338 3225
rect 3464 3209 3466 3225
rect 3462 3208 3468 3209
rect 1806 3204 1807 3208
rect 1811 3204 1812 3208
rect 1806 3203 1812 3204
rect 1910 3207 1916 3208
rect 1910 3203 1911 3207
rect 1915 3203 1916 3207
rect 1910 3202 1916 3203
rect 2046 3207 2052 3208
rect 2046 3203 2047 3207
rect 2051 3203 2052 3207
rect 2046 3202 2052 3203
rect 2198 3207 2204 3208
rect 2198 3203 2199 3207
rect 2203 3203 2204 3207
rect 2198 3202 2204 3203
rect 2358 3207 2364 3208
rect 2358 3203 2359 3207
rect 2363 3203 2364 3207
rect 2358 3202 2364 3203
rect 2526 3207 2532 3208
rect 2526 3203 2527 3207
rect 2531 3203 2532 3207
rect 2526 3202 2532 3203
rect 2686 3207 2692 3208
rect 2686 3203 2687 3207
rect 2691 3203 2692 3207
rect 2686 3202 2692 3203
rect 2846 3207 2852 3208
rect 2846 3203 2847 3207
rect 2851 3203 2852 3207
rect 2846 3202 2852 3203
rect 3006 3207 3012 3208
rect 3006 3203 3007 3207
rect 3011 3203 3012 3207
rect 3006 3202 3012 3203
rect 3166 3207 3172 3208
rect 3166 3203 3167 3207
rect 3171 3203 3172 3207
rect 3166 3202 3172 3203
rect 3334 3207 3340 3208
rect 3334 3203 3335 3207
rect 3339 3203 3340 3207
rect 3462 3204 3463 3208
rect 3467 3204 3468 3208
rect 3462 3203 3468 3204
rect 3334 3202 3340 3203
rect 1766 3200 1772 3201
rect 110 3196 111 3200
rect 115 3196 116 3200
rect 110 3195 116 3196
rect 182 3199 188 3200
rect 182 3195 183 3199
rect 187 3195 188 3199
rect 182 3194 188 3195
rect 326 3199 332 3200
rect 326 3195 327 3199
rect 331 3195 332 3199
rect 326 3194 332 3195
rect 486 3199 492 3200
rect 486 3195 487 3199
rect 491 3195 492 3199
rect 486 3194 492 3195
rect 646 3199 652 3200
rect 646 3195 647 3199
rect 651 3195 652 3199
rect 646 3194 652 3195
rect 806 3199 812 3200
rect 806 3195 807 3199
rect 811 3195 812 3199
rect 806 3194 812 3195
rect 966 3199 972 3200
rect 966 3195 967 3199
rect 971 3195 972 3199
rect 966 3194 972 3195
rect 1134 3199 1140 3200
rect 1134 3195 1135 3199
rect 1139 3195 1140 3199
rect 1134 3194 1140 3195
rect 1302 3199 1308 3200
rect 1302 3195 1303 3199
rect 1307 3195 1308 3199
rect 1302 3194 1308 3195
rect 1470 3199 1476 3200
rect 1470 3195 1471 3199
rect 1475 3195 1476 3199
rect 1766 3196 1767 3200
rect 1771 3196 1772 3200
rect 1766 3195 1772 3196
rect 1470 3194 1476 3195
rect 1806 3191 1812 3192
rect 1806 3187 1807 3191
rect 1811 3187 1812 3191
rect 3462 3191 3468 3192
rect 1806 3186 1812 3187
rect 1910 3188 1916 3189
rect 110 3183 116 3184
rect 110 3179 111 3183
rect 115 3179 116 3183
rect 1766 3183 1772 3184
rect 110 3178 116 3179
rect 182 3180 188 3181
rect 112 3159 114 3178
rect 182 3176 183 3180
rect 187 3176 188 3180
rect 182 3175 188 3176
rect 326 3180 332 3181
rect 326 3176 327 3180
rect 331 3176 332 3180
rect 326 3175 332 3176
rect 486 3180 492 3181
rect 486 3176 487 3180
rect 491 3176 492 3180
rect 486 3175 492 3176
rect 646 3180 652 3181
rect 646 3176 647 3180
rect 651 3176 652 3180
rect 646 3175 652 3176
rect 806 3180 812 3181
rect 806 3176 807 3180
rect 811 3176 812 3180
rect 806 3175 812 3176
rect 966 3180 972 3181
rect 966 3176 967 3180
rect 971 3176 972 3180
rect 966 3175 972 3176
rect 1134 3180 1140 3181
rect 1134 3176 1135 3180
rect 1139 3176 1140 3180
rect 1134 3175 1140 3176
rect 1302 3180 1308 3181
rect 1302 3176 1303 3180
rect 1307 3176 1308 3180
rect 1302 3175 1308 3176
rect 1470 3180 1476 3181
rect 1470 3176 1471 3180
rect 1475 3176 1476 3180
rect 1766 3179 1767 3183
rect 1771 3179 1772 3183
rect 1766 3178 1772 3179
rect 1470 3175 1476 3176
rect 184 3159 186 3175
rect 328 3159 330 3175
rect 488 3159 490 3175
rect 648 3159 650 3175
rect 808 3159 810 3175
rect 968 3159 970 3175
rect 1136 3159 1138 3175
rect 1304 3159 1306 3175
rect 1472 3159 1474 3175
rect 1768 3159 1770 3178
rect 1808 3167 1810 3186
rect 1910 3184 1911 3188
rect 1915 3184 1916 3188
rect 1910 3183 1916 3184
rect 2046 3188 2052 3189
rect 2046 3184 2047 3188
rect 2051 3184 2052 3188
rect 2046 3183 2052 3184
rect 2198 3188 2204 3189
rect 2198 3184 2199 3188
rect 2203 3184 2204 3188
rect 2198 3183 2204 3184
rect 2358 3188 2364 3189
rect 2358 3184 2359 3188
rect 2363 3184 2364 3188
rect 2358 3183 2364 3184
rect 2526 3188 2532 3189
rect 2526 3184 2527 3188
rect 2531 3184 2532 3188
rect 2526 3183 2532 3184
rect 2686 3188 2692 3189
rect 2686 3184 2687 3188
rect 2691 3184 2692 3188
rect 2686 3183 2692 3184
rect 2846 3188 2852 3189
rect 2846 3184 2847 3188
rect 2851 3184 2852 3188
rect 2846 3183 2852 3184
rect 3006 3188 3012 3189
rect 3006 3184 3007 3188
rect 3011 3184 3012 3188
rect 3006 3183 3012 3184
rect 3166 3188 3172 3189
rect 3166 3184 3167 3188
rect 3171 3184 3172 3188
rect 3166 3183 3172 3184
rect 3334 3188 3340 3189
rect 3334 3184 3335 3188
rect 3339 3184 3340 3188
rect 3462 3187 3463 3191
rect 3467 3187 3468 3191
rect 3462 3186 3468 3187
rect 3334 3183 3340 3184
rect 1912 3167 1914 3183
rect 2048 3167 2050 3183
rect 2200 3167 2202 3183
rect 2360 3167 2362 3183
rect 2528 3167 2530 3183
rect 2688 3167 2690 3183
rect 2848 3167 2850 3183
rect 3008 3167 3010 3183
rect 3168 3167 3170 3183
rect 3336 3167 3338 3183
rect 3464 3167 3466 3186
rect 1807 3166 1811 3167
rect 1807 3161 1811 3162
rect 1831 3166 1835 3167
rect 1831 3161 1835 3162
rect 1911 3166 1915 3167
rect 1911 3161 1915 3162
rect 2007 3166 2011 3167
rect 2007 3161 2011 3162
rect 2047 3166 2051 3167
rect 2047 3161 2051 3162
rect 2199 3166 2203 3167
rect 2199 3161 2203 3162
rect 2207 3166 2211 3167
rect 2207 3161 2211 3162
rect 2359 3166 2363 3167
rect 2359 3161 2363 3162
rect 2399 3166 2403 3167
rect 2399 3161 2403 3162
rect 2527 3166 2531 3167
rect 2527 3161 2531 3162
rect 2583 3166 2587 3167
rect 2583 3161 2587 3162
rect 2687 3166 2691 3167
rect 2687 3161 2691 3162
rect 2759 3166 2763 3167
rect 2759 3161 2763 3162
rect 2847 3166 2851 3167
rect 2847 3161 2851 3162
rect 2919 3166 2923 3167
rect 2919 3161 2923 3162
rect 3007 3166 3011 3167
rect 3007 3161 3011 3162
rect 3079 3166 3083 3167
rect 3079 3161 3083 3162
rect 3167 3166 3171 3167
rect 3167 3161 3171 3162
rect 3231 3166 3235 3167
rect 3231 3161 3235 3162
rect 3335 3166 3339 3167
rect 3335 3161 3339 3162
rect 3367 3166 3371 3167
rect 3367 3161 3371 3162
rect 3463 3166 3467 3167
rect 3463 3161 3467 3162
rect 111 3158 115 3159
rect 111 3153 115 3154
rect 183 3158 187 3159
rect 183 3153 187 3154
rect 327 3158 331 3159
rect 327 3153 331 3154
rect 367 3158 371 3159
rect 367 3153 371 3154
rect 487 3158 491 3159
rect 487 3153 491 3154
rect 607 3158 611 3159
rect 607 3153 611 3154
rect 647 3158 651 3159
rect 647 3153 651 3154
rect 727 3158 731 3159
rect 727 3153 731 3154
rect 807 3158 811 3159
rect 807 3153 811 3154
rect 847 3158 851 3159
rect 847 3153 851 3154
rect 967 3158 971 3159
rect 967 3153 971 3154
rect 1079 3158 1083 3159
rect 1079 3153 1083 3154
rect 1135 3158 1139 3159
rect 1135 3153 1139 3154
rect 1199 3158 1203 3159
rect 1199 3153 1203 3154
rect 1303 3158 1307 3159
rect 1303 3153 1307 3154
rect 1319 3158 1323 3159
rect 1319 3153 1323 3154
rect 1471 3158 1475 3159
rect 1471 3153 1475 3154
rect 1767 3158 1771 3159
rect 1767 3153 1771 3154
rect 112 3134 114 3153
rect 368 3137 370 3153
rect 488 3137 490 3153
rect 608 3137 610 3153
rect 728 3137 730 3153
rect 848 3137 850 3153
rect 968 3137 970 3153
rect 1080 3137 1082 3153
rect 1200 3137 1202 3153
rect 1320 3137 1322 3153
rect 366 3136 372 3137
rect 110 3133 116 3134
rect 110 3129 111 3133
rect 115 3129 116 3133
rect 366 3132 367 3136
rect 371 3132 372 3136
rect 366 3131 372 3132
rect 486 3136 492 3137
rect 486 3132 487 3136
rect 491 3132 492 3136
rect 486 3131 492 3132
rect 606 3136 612 3137
rect 606 3132 607 3136
rect 611 3132 612 3136
rect 606 3131 612 3132
rect 726 3136 732 3137
rect 726 3132 727 3136
rect 731 3132 732 3136
rect 726 3131 732 3132
rect 846 3136 852 3137
rect 846 3132 847 3136
rect 851 3132 852 3136
rect 846 3131 852 3132
rect 966 3136 972 3137
rect 966 3132 967 3136
rect 971 3132 972 3136
rect 966 3131 972 3132
rect 1078 3136 1084 3137
rect 1078 3132 1079 3136
rect 1083 3132 1084 3136
rect 1078 3131 1084 3132
rect 1198 3136 1204 3137
rect 1198 3132 1199 3136
rect 1203 3132 1204 3136
rect 1198 3131 1204 3132
rect 1318 3136 1324 3137
rect 1318 3132 1319 3136
rect 1323 3132 1324 3136
rect 1768 3134 1770 3153
rect 1808 3142 1810 3161
rect 1832 3145 1834 3161
rect 2008 3145 2010 3161
rect 2208 3145 2210 3161
rect 2400 3145 2402 3161
rect 2584 3145 2586 3161
rect 2760 3145 2762 3161
rect 2920 3145 2922 3161
rect 3080 3145 3082 3161
rect 3232 3145 3234 3161
rect 3368 3145 3370 3161
rect 1830 3144 1836 3145
rect 1806 3141 1812 3142
rect 1806 3137 1807 3141
rect 1811 3137 1812 3141
rect 1830 3140 1831 3144
rect 1835 3140 1836 3144
rect 1830 3139 1836 3140
rect 2006 3144 2012 3145
rect 2006 3140 2007 3144
rect 2011 3140 2012 3144
rect 2006 3139 2012 3140
rect 2206 3144 2212 3145
rect 2206 3140 2207 3144
rect 2211 3140 2212 3144
rect 2206 3139 2212 3140
rect 2398 3144 2404 3145
rect 2398 3140 2399 3144
rect 2403 3140 2404 3144
rect 2398 3139 2404 3140
rect 2582 3144 2588 3145
rect 2582 3140 2583 3144
rect 2587 3140 2588 3144
rect 2582 3139 2588 3140
rect 2758 3144 2764 3145
rect 2758 3140 2759 3144
rect 2763 3140 2764 3144
rect 2758 3139 2764 3140
rect 2918 3144 2924 3145
rect 2918 3140 2919 3144
rect 2923 3140 2924 3144
rect 2918 3139 2924 3140
rect 3078 3144 3084 3145
rect 3078 3140 3079 3144
rect 3083 3140 3084 3144
rect 3078 3139 3084 3140
rect 3230 3144 3236 3145
rect 3230 3140 3231 3144
rect 3235 3140 3236 3144
rect 3230 3139 3236 3140
rect 3366 3144 3372 3145
rect 3366 3140 3367 3144
rect 3371 3140 3372 3144
rect 3464 3142 3466 3161
rect 3366 3139 3372 3140
rect 3462 3141 3468 3142
rect 1806 3136 1812 3137
rect 3462 3137 3463 3141
rect 3467 3137 3468 3141
rect 3462 3136 3468 3137
rect 1318 3131 1324 3132
rect 1766 3133 1772 3134
rect 110 3128 116 3129
rect 1766 3129 1767 3133
rect 1771 3129 1772 3133
rect 1766 3128 1772 3129
rect 1830 3125 1836 3126
rect 1806 3124 1812 3125
rect 1806 3120 1807 3124
rect 1811 3120 1812 3124
rect 1830 3121 1831 3125
rect 1835 3121 1836 3125
rect 1830 3120 1836 3121
rect 2006 3125 2012 3126
rect 2006 3121 2007 3125
rect 2011 3121 2012 3125
rect 2006 3120 2012 3121
rect 2206 3125 2212 3126
rect 2206 3121 2207 3125
rect 2211 3121 2212 3125
rect 2206 3120 2212 3121
rect 2398 3125 2404 3126
rect 2398 3121 2399 3125
rect 2403 3121 2404 3125
rect 2398 3120 2404 3121
rect 2582 3125 2588 3126
rect 2582 3121 2583 3125
rect 2587 3121 2588 3125
rect 2582 3120 2588 3121
rect 2758 3125 2764 3126
rect 2758 3121 2759 3125
rect 2763 3121 2764 3125
rect 2758 3120 2764 3121
rect 2918 3125 2924 3126
rect 2918 3121 2919 3125
rect 2923 3121 2924 3125
rect 2918 3120 2924 3121
rect 3078 3125 3084 3126
rect 3078 3121 3079 3125
rect 3083 3121 3084 3125
rect 3078 3120 3084 3121
rect 3230 3125 3236 3126
rect 3230 3121 3231 3125
rect 3235 3121 3236 3125
rect 3230 3120 3236 3121
rect 3366 3125 3372 3126
rect 3366 3121 3367 3125
rect 3371 3121 3372 3125
rect 3366 3120 3372 3121
rect 3462 3124 3468 3125
rect 3462 3120 3463 3124
rect 3467 3120 3468 3124
rect 1806 3119 1812 3120
rect 366 3117 372 3118
rect 110 3116 116 3117
rect 110 3112 111 3116
rect 115 3112 116 3116
rect 366 3113 367 3117
rect 371 3113 372 3117
rect 366 3112 372 3113
rect 486 3117 492 3118
rect 486 3113 487 3117
rect 491 3113 492 3117
rect 486 3112 492 3113
rect 606 3117 612 3118
rect 606 3113 607 3117
rect 611 3113 612 3117
rect 606 3112 612 3113
rect 726 3117 732 3118
rect 726 3113 727 3117
rect 731 3113 732 3117
rect 726 3112 732 3113
rect 846 3117 852 3118
rect 846 3113 847 3117
rect 851 3113 852 3117
rect 846 3112 852 3113
rect 966 3117 972 3118
rect 966 3113 967 3117
rect 971 3113 972 3117
rect 966 3112 972 3113
rect 1078 3117 1084 3118
rect 1078 3113 1079 3117
rect 1083 3113 1084 3117
rect 1078 3112 1084 3113
rect 1198 3117 1204 3118
rect 1198 3113 1199 3117
rect 1203 3113 1204 3117
rect 1198 3112 1204 3113
rect 1318 3117 1324 3118
rect 1318 3113 1319 3117
rect 1323 3113 1324 3117
rect 1318 3112 1324 3113
rect 1766 3116 1772 3117
rect 1766 3112 1767 3116
rect 1771 3112 1772 3116
rect 110 3111 116 3112
rect 112 3091 114 3111
rect 368 3091 370 3112
rect 488 3091 490 3112
rect 608 3091 610 3112
rect 728 3091 730 3112
rect 848 3091 850 3112
rect 968 3091 970 3112
rect 1080 3091 1082 3112
rect 1200 3091 1202 3112
rect 1320 3091 1322 3112
rect 1766 3111 1772 3112
rect 1768 3091 1770 3111
rect 1808 3095 1810 3119
rect 1832 3095 1834 3120
rect 2008 3095 2010 3120
rect 2208 3095 2210 3120
rect 2400 3095 2402 3120
rect 2584 3095 2586 3120
rect 2760 3095 2762 3120
rect 2920 3095 2922 3120
rect 3080 3095 3082 3120
rect 3232 3095 3234 3120
rect 3368 3095 3370 3120
rect 3462 3119 3468 3120
rect 3464 3095 3466 3119
rect 1807 3094 1811 3095
rect 111 3090 115 3091
rect 111 3085 115 3086
rect 367 3090 371 3091
rect 367 3085 371 3086
rect 439 3090 443 3091
rect 439 3085 443 3086
rect 487 3090 491 3091
rect 487 3085 491 3086
rect 527 3090 531 3091
rect 527 3085 531 3086
rect 607 3090 611 3091
rect 607 3085 611 3086
rect 615 3090 619 3091
rect 615 3085 619 3086
rect 703 3090 707 3091
rect 703 3085 707 3086
rect 727 3090 731 3091
rect 727 3085 731 3086
rect 791 3090 795 3091
rect 791 3085 795 3086
rect 847 3090 851 3091
rect 847 3085 851 3086
rect 879 3090 883 3091
rect 879 3085 883 3086
rect 967 3090 971 3091
rect 967 3085 971 3086
rect 1055 3090 1059 3091
rect 1055 3085 1059 3086
rect 1079 3090 1083 3091
rect 1079 3085 1083 3086
rect 1143 3090 1147 3091
rect 1143 3085 1147 3086
rect 1199 3090 1203 3091
rect 1199 3085 1203 3086
rect 1319 3090 1323 3091
rect 1319 3085 1323 3086
rect 1767 3090 1771 3091
rect 1807 3089 1811 3090
rect 1831 3094 1835 3095
rect 1831 3089 1835 3090
rect 1959 3094 1963 3095
rect 1959 3089 1963 3090
rect 2007 3094 2011 3095
rect 2007 3089 2011 3090
rect 2119 3094 2123 3095
rect 2119 3089 2123 3090
rect 2207 3094 2211 3095
rect 2207 3089 2211 3090
rect 2295 3094 2299 3095
rect 2295 3089 2299 3090
rect 2399 3094 2403 3095
rect 2399 3089 2403 3090
rect 2487 3094 2491 3095
rect 2487 3089 2491 3090
rect 2583 3094 2587 3095
rect 2583 3089 2587 3090
rect 2695 3094 2699 3095
rect 2695 3089 2699 3090
rect 2759 3094 2763 3095
rect 2759 3089 2763 3090
rect 2919 3094 2923 3095
rect 2919 3089 2923 3090
rect 3079 3094 3083 3095
rect 3079 3089 3083 3090
rect 3151 3094 3155 3095
rect 3151 3089 3155 3090
rect 3231 3094 3235 3095
rect 3231 3089 3235 3090
rect 3367 3094 3371 3095
rect 3367 3089 3371 3090
rect 3463 3094 3467 3095
rect 3463 3089 3467 3090
rect 1767 3085 1771 3086
rect 112 3069 114 3085
rect 110 3068 116 3069
rect 440 3068 442 3085
rect 528 3068 530 3085
rect 616 3068 618 3085
rect 704 3068 706 3085
rect 792 3068 794 3085
rect 880 3068 882 3085
rect 968 3068 970 3085
rect 1056 3068 1058 3085
rect 1144 3068 1146 3085
rect 1768 3069 1770 3085
rect 1808 3073 1810 3089
rect 1806 3072 1812 3073
rect 1832 3072 1834 3089
rect 1960 3072 1962 3089
rect 2120 3072 2122 3089
rect 2296 3072 2298 3089
rect 2488 3072 2490 3089
rect 2696 3072 2698 3089
rect 2920 3072 2922 3089
rect 3152 3072 3154 3089
rect 3368 3072 3370 3089
rect 3464 3073 3466 3089
rect 3462 3072 3468 3073
rect 1766 3068 1772 3069
rect 110 3064 111 3068
rect 115 3064 116 3068
rect 110 3063 116 3064
rect 438 3067 444 3068
rect 438 3063 439 3067
rect 443 3063 444 3067
rect 438 3062 444 3063
rect 526 3067 532 3068
rect 526 3063 527 3067
rect 531 3063 532 3067
rect 526 3062 532 3063
rect 614 3067 620 3068
rect 614 3063 615 3067
rect 619 3063 620 3067
rect 614 3062 620 3063
rect 702 3067 708 3068
rect 702 3063 703 3067
rect 707 3063 708 3067
rect 702 3062 708 3063
rect 790 3067 796 3068
rect 790 3063 791 3067
rect 795 3063 796 3067
rect 790 3062 796 3063
rect 878 3067 884 3068
rect 878 3063 879 3067
rect 883 3063 884 3067
rect 878 3062 884 3063
rect 966 3067 972 3068
rect 966 3063 967 3067
rect 971 3063 972 3067
rect 966 3062 972 3063
rect 1054 3067 1060 3068
rect 1054 3063 1055 3067
rect 1059 3063 1060 3067
rect 1054 3062 1060 3063
rect 1142 3067 1148 3068
rect 1142 3063 1143 3067
rect 1147 3063 1148 3067
rect 1766 3064 1767 3068
rect 1771 3064 1772 3068
rect 1806 3068 1807 3072
rect 1811 3068 1812 3072
rect 1806 3067 1812 3068
rect 1830 3071 1836 3072
rect 1830 3067 1831 3071
rect 1835 3067 1836 3071
rect 1830 3066 1836 3067
rect 1958 3071 1964 3072
rect 1958 3067 1959 3071
rect 1963 3067 1964 3071
rect 1958 3066 1964 3067
rect 2118 3071 2124 3072
rect 2118 3067 2119 3071
rect 2123 3067 2124 3071
rect 2118 3066 2124 3067
rect 2294 3071 2300 3072
rect 2294 3067 2295 3071
rect 2299 3067 2300 3071
rect 2294 3066 2300 3067
rect 2486 3071 2492 3072
rect 2486 3067 2487 3071
rect 2491 3067 2492 3071
rect 2486 3066 2492 3067
rect 2694 3071 2700 3072
rect 2694 3067 2695 3071
rect 2699 3067 2700 3071
rect 2694 3066 2700 3067
rect 2918 3071 2924 3072
rect 2918 3067 2919 3071
rect 2923 3067 2924 3071
rect 2918 3066 2924 3067
rect 3150 3071 3156 3072
rect 3150 3067 3151 3071
rect 3155 3067 3156 3071
rect 3150 3066 3156 3067
rect 3366 3071 3372 3072
rect 3366 3067 3367 3071
rect 3371 3067 3372 3071
rect 3462 3068 3463 3072
rect 3467 3068 3468 3072
rect 3462 3067 3468 3068
rect 3366 3066 3372 3067
rect 1766 3063 1772 3064
rect 1142 3062 1148 3063
rect 1806 3055 1812 3056
rect 110 3051 116 3052
rect 110 3047 111 3051
rect 115 3047 116 3051
rect 1766 3051 1772 3052
rect 110 3046 116 3047
rect 438 3048 444 3049
rect 112 3019 114 3046
rect 438 3044 439 3048
rect 443 3044 444 3048
rect 438 3043 444 3044
rect 526 3048 532 3049
rect 526 3044 527 3048
rect 531 3044 532 3048
rect 526 3043 532 3044
rect 614 3048 620 3049
rect 614 3044 615 3048
rect 619 3044 620 3048
rect 614 3043 620 3044
rect 702 3048 708 3049
rect 702 3044 703 3048
rect 707 3044 708 3048
rect 702 3043 708 3044
rect 790 3048 796 3049
rect 790 3044 791 3048
rect 795 3044 796 3048
rect 790 3043 796 3044
rect 878 3048 884 3049
rect 878 3044 879 3048
rect 883 3044 884 3048
rect 878 3043 884 3044
rect 966 3048 972 3049
rect 966 3044 967 3048
rect 971 3044 972 3048
rect 966 3043 972 3044
rect 1054 3048 1060 3049
rect 1054 3044 1055 3048
rect 1059 3044 1060 3048
rect 1054 3043 1060 3044
rect 1142 3048 1148 3049
rect 1142 3044 1143 3048
rect 1147 3044 1148 3048
rect 1766 3047 1767 3051
rect 1771 3047 1772 3051
rect 1806 3051 1807 3055
rect 1811 3051 1812 3055
rect 3462 3055 3468 3056
rect 1806 3050 1812 3051
rect 1830 3052 1836 3053
rect 1766 3046 1772 3047
rect 1142 3043 1148 3044
rect 440 3019 442 3043
rect 528 3019 530 3043
rect 616 3019 618 3043
rect 704 3019 706 3043
rect 792 3019 794 3043
rect 880 3019 882 3043
rect 968 3019 970 3043
rect 1056 3019 1058 3043
rect 1144 3019 1146 3043
rect 1768 3019 1770 3046
rect 111 3018 115 3019
rect 111 3013 115 3014
rect 439 3018 443 3019
rect 439 3013 443 3014
rect 503 3018 507 3019
rect 503 3013 507 3014
rect 527 3018 531 3019
rect 527 3013 531 3014
rect 591 3018 595 3019
rect 591 3013 595 3014
rect 615 3018 619 3019
rect 615 3013 619 3014
rect 679 3018 683 3019
rect 679 3013 683 3014
rect 703 3018 707 3019
rect 703 3013 707 3014
rect 767 3018 771 3019
rect 767 3013 771 3014
rect 791 3018 795 3019
rect 791 3013 795 3014
rect 855 3018 859 3019
rect 855 3013 859 3014
rect 879 3018 883 3019
rect 879 3013 883 3014
rect 943 3018 947 3019
rect 943 3013 947 3014
rect 967 3018 971 3019
rect 967 3013 971 3014
rect 1031 3018 1035 3019
rect 1031 3013 1035 3014
rect 1055 3018 1059 3019
rect 1055 3013 1059 3014
rect 1119 3018 1123 3019
rect 1119 3013 1123 3014
rect 1143 3018 1147 3019
rect 1143 3013 1147 3014
rect 1207 3018 1211 3019
rect 1207 3013 1211 3014
rect 1295 3018 1299 3019
rect 1295 3013 1299 3014
rect 1767 3018 1771 3019
rect 1808 3015 1810 3050
rect 1830 3048 1831 3052
rect 1835 3048 1836 3052
rect 1830 3047 1836 3048
rect 1958 3052 1964 3053
rect 1958 3048 1959 3052
rect 1963 3048 1964 3052
rect 1958 3047 1964 3048
rect 2118 3052 2124 3053
rect 2118 3048 2119 3052
rect 2123 3048 2124 3052
rect 2118 3047 2124 3048
rect 2294 3052 2300 3053
rect 2294 3048 2295 3052
rect 2299 3048 2300 3052
rect 2294 3047 2300 3048
rect 2486 3052 2492 3053
rect 2486 3048 2487 3052
rect 2491 3048 2492 3052
rect 2486 3047 2492 3048
rect 2694 3052 2700 3053
rect 2694 3048 2695 3052
rect 2699 3048 2700 3052
rect 2694 3047 2700 3048
rect 2918 3052 2924 3053
rect 2918 3048 2919 3052
rect 2923 3048 2924 3052
rect 2918 3047 2924 3048
rect 3150 3052 3156 3053
rect 3150 3048 3151 3052
rect 3155 3048 3156 3052
rect 3150 3047 3156 3048
rect 3366 3052 3372 3053
rect 3366 3048 3367 3052
rect 3371 3048 3372 3052
rect 3462 3051 3463 3055
rect 3467 3051 3468 3055
rect 3462 3050 3468 3051
rect 3366 3047 3372 3048
rect 1832 3015 1834 3047
rect 1960 3015 1962 3047
rect 2120 3015 2122 3047
rect 2296 3015 2298 3047
rect 2488 3015 2490 3047
rect 2696 3015 2698 3047
rect 2920 3015 2922 3047
rect 3152 3015 3154 3047
rect 3368 3015 3370 3047
rect 3464 3015 3466 3050
rect 1767 3013 1771 3014
rect 1807 3014 1811 3015
rect 112 2994 114 3013
rect 504 2997 506 3013
rect 592 2997 594 3013
rect 680 2997 682 3013
rect 768 2997 770 3013
rect 856 2997 858 3013
rect 944 2997 946 3013
rect 1032 2997 1034 3013
rect 1120 2997 1122 3013
rect 1208 2997 1210 3013
rect 1296 2997 1298 3013
rect 502 2996 508 2997
rect 110 2993 116 2994
rect 110 2989 111 2993
rect 115 2989 116 2993
rect 502 2992 503 2996
rect 507 2992 508 2996
rect 502 2991 508 2992
rect 590 2996 596 2997
rect 590 2992 591 2996
rect 595 2992 596 2996
rect 590 2991 596 2992
rect 678 2996 684 2997
rect 678 2992 679 2996
rect 683 2992 684 2996
rect 678 2991 684 2992
rect 766 2996 772 2997
rect 766 2992 767 2996
rect 771 2992 772 2996
rect 766 2991 772 2992
rect 854 2996 860 2997
rect 854 2992 855 2996
rect 859 2992 860 2996
rect 854 2991 860 2992
rect 942 2996 948 2997
rect 942 2992 943 2996
rect 947 2992 948 2996
rect 942 2991 948 2992
rect 1030 2996 1036 2997
rect 1030 2992 1031 2996
rect 1035 2992 1036 2996
rect 1030 2991 1036 2992
rect 1118 2996 1124 2997
rect 1118 2992 1119 2996
rect 1123 2992 1124 2996
rect 1118 2991 1124 2992
rect 1206 2996 1212 2997
rect 1206 2992 1207 2996
rect 1211 2992 1212 2996
rect 1206 2991 1212 2992
rect 1294 2996 1300 2997
rect 1294 2992 1295 2996
rect 1299 2992 1300 2996
rect 1768 2994 1770 3013
rect 1807 3009 1811 3010
rect 1831 3014 1835 3015
rect 1831 3009 1835 3010
rect 1919 3014 1923 3015
rect 1919 3009 1923 3010
rect 1959 3014 1963 3015
rect 1959 3009 1963 3010
rect 2031 3014 2035 3015
rect 2031 3009 2035 3010
rect 2119 3014 2123 3015
rect 2119 3009 2123 3010
rect 2143 3014 2147 3015
rect 2143 3009 2147 3010
rect 2247 3014 2251 3015
rect 2247 3009 2251 3010
rect 2295 3014 2299 3015
rect 2295 3009 2299 3010
rect 2359 3014 2363 3015
rect 2359 3009 2363 3010
rect 2479 3014 2483 3015
rect 2479 3009 2483 3010
rect 2487 3014 2491 3015
rect 2487 3009 2491 3010
rect 2623 3014 2627 3015
rect 2623 3009 2627 3010
rect 2695 3014 2699 3015
rect 2695 3009 2699 3010
rect 2791 3014 2795 3015
rect 2791 3009 2795 3010
rect 2919 3014 2923 3015
rect 2919 3009 2923 3010
rect 2983 3014 2987 3015
rect 2983 3009 2987 3010
rect 3151 3014 3155 3015
rect 3151 3009 3155 3010
rect 3183 3014 3187 3015
rect 3183 3009 3187 3010
rect 3367 3014 3371 3015
rect 3367 3009 3371 3010
rect 3463 3014 3467 3015
rect 3463 3009 3467 3010
rect 1294 2991 1300 2992
rect 1766 2993 1772 2994
rect 110 2988 116 2989
rect 1766 2989 1767 2993
rect 1771 2989 1772 2993
rect 1808 2990 1810 3009
rect 1832 2993 1834 3009
rect 1920 2993 1922 3009
rect 2032 2993 2034 3009
rect 2144 2993 2146 3009
rect 2248 2993 2250 3009
rect 2360 2993 2362 3009
rect 2480 2993 2482 3009
rect 2624 2993 2626 3009
rect 2792 2993 2794 3009
rect 2984 2993 2986 3009
rect 3184 2993 3186 3009
rect 3368 2993 3370 3009
rect 1830 2992 1836 2993
rect 1766 2988 1772 2989
rect 1806 2989 1812 2990
rect 1806 2985 1807 2989
rect 1811 2985 1812 2989
rect 1830 2988 1831 2992
rect 1835 2988 1836 2992
rect 1830 2987 1836 2988
rect 1918 2992 1924 2993
rect 1918 2988 1919 2992
rect 1923 2988 1924 2992
rect 1918 2987 1924 2988
rect 2030 2992 2036 2993
rect 2030 2988 2031 2992
rect 2035 2988 2036 2992
rect 2030 2987 2036 2988
rect 2142 2992 2148 2993
rect 2142 2988 2143 2992
rect 2147 2988 2148 2992
rect 2142 2987 2148 2988
rect 2246 2992 2252 2993
rect 2246 2988 2247 2992
rect 2251 2988 2252 2992
rect 2246 2987 2252 2988
rect 2358 2992 2364 2993
rect 2358 2988 2359 2992
rect 2363 2988 2364 2992
rect 2358 2987 2364 2988
rect 2478 2992 2484 2993
rect 2478 2988 2479 2992
rect 2483 2988 2484 2992
rect 2478 2987 2484 2988
rect 2622 2992 2628 2993
rect 2622 2988 2623 2992
rect 2627 2988 2628 2992
rect 2622 2987 2628 2988
rect 2790 2992 2796 2993
rect 2790 2988 2791 2992
rect 2795 2988 2796 2992
rect 2790 2987 2796 2988
rect 2982 2992 2988 2993
rect 2982 2988 2983 2992
rect 2987 2988 2988 2992
rect 2982 2987 2988 2988
rect 3182 2992 3188 2993
rect 3182 2988 3183 2992
rect 3187 2988 3188 2992
rect 3182 2987 3188 2988
rect 3366 2992 3372 2993
rect 3366 2988 3367 2992
rect 3371 2988 3372 2992
rect 3464 2990 3466 3009
rect 3366 2987 3372 2988
rect 3462 2989 3468 2990
rect 1806 2984 1812 2985
rect 3462 2985 3463 2989
rect 3467 2985 3468 2989
rect 3462 2984 3468 2985
rect 502 2977 508 2978
rect 110 2976 116 2977
rect 110 2972 111 2976
rect 115 2972 116 2976
rect 502 2973 503 2977
rect 507 2973 508 2977
rect 502 2972 508 2973
rect 590 2977 596 2978
rect 590 2973 591 2977
rect 595 2973 596 2977
rect 590 2972 596 2973
rect 678 2977 684 2978
rect 678 2973 679 2977
rect 683 2973 684 2977
rect 678 2972 684 2973
rect 766 2977 772 2978
rect 766 2973 767 2977
rect 771 2973 772 2977
rect 766 2972 772 2973
rect 854 2977 860 2978
rect 854 2973 855 2977
rect 859 2973 860 2977
rect 854 2972 860 2973
rect 942 2977 948 2978
rect 942 2973 943 2977
rect 947 2973 948 2977
rect 942 2972 948 2973
rect 1030 2977 1036 2978
rect 1030 2973 1031 2977
rect 1035 2973 1036 2977
rect 1030 2972 1036 2973
rect 1118 2977 1124 2978
rect 1118 2973 1119 2977
rect 1123 2973 1124 2977
rect 1118 2972 1124 2973
rect 1206 2977 1212 2978
rect 1206 2973 1207 2977
rect 1211 2973 1212 2977
rect 1206 2972 1212 2973
rect 1294 2977 1300 2978
rect 1294 2973 1295 2977
rect 1299 2973 1300 2977
rect 1294 2972 1300 2973
rect 1766 2976 1772 2977
rect 1766 2972 1767 2976
rect 1771 2972 1772 2976
rect 1830 2973 1836 2974
rect 110 2971 116 2972
rect 112 2943 114 2971
rect 504 2943 506 2972
rect 592 2943 594 2972
rect 680 2943 682 2972
rect 768 2943 770 2972
rect 856 2943 858 2972
rect 944 2943 946 2972
rect 1032 2943 1034 2972
rect 1120 2943 1122 2972
rect 1208 2943 1210 2972
rect 1296 2943 1298 2972
rect 1766 2971 1772 2972
rect 1806 2972 1812 2973
rect 1768 2943 1770 2971
rect 1806 2968 1807 2972
rect 1811 2968 1812 2972
rect 1830 2969 1831 2973
rect 1835 2969 1836 2973
rect 1830 2968 1836 2969
rect 1918 2973 1924 2974
rect 1918 2969 1919 2973
rect 1923 2969 1924 2973
rect 1918 2968 1924 2969
rect 2030 2973 2036 2974
rect 2030 2969 2031 2973
rect 2035 2969 2036 2973
rect 2030 2968 2036 2969
rect 2142 2973 2148 2974
rect 2142 2969 2143 2973
rect 2147 2969 2148 2973
rect 2142 2968 2148 2969
rect 2246 2973 2252 2974
rect 2246 2969 2247 2973
rect 2251 2969 2252 2973
rect 2246 2968 2252 2969
rect 2358 2973 2364 2974
rect 2358 2969 2359 2973
rect 2363 2969 2364 2973
rect 2358 2968 2364 2969
rect 2478 2973 2484 2974
rect 2478 2969 2479 2973
rect 2483 2969 2484 2973
rect 2478 2968 2484 2969
rect 2622 2973 2628 2974
rect 2622 2969 2623 2973
rect 2627 2969 2628 2973
rect 2622 2968 2628 2969
rect 2790 2973 2796 2974
rect 2790 2969 2791 2973
rect 2795 2969 2796 2973
rect 2790 2968 2796 2969
rect 2982 2973 2988 2974
rect 2982 2969 2983 2973
rect 2987 2969 2988 2973
rect 2982 2968 2988 2969
rect 3182 2973 3188 2974
rect 3182 2969 3183 2973
rect 3187 2969 3188 2973
rect 3182 2968 3188 2969
rect 3366 2973 3372 2974
rect 3366 2969 3367 2973
rect 3371 2969 3372 2973
rect 3366 2968 3372 2969
rect 3462 2972 3468 2973
rect 3462 2968 3463 2972
rect 3467 2968 3468 2972
rect 1806 2967 1812 2968
rect 111 2942 115 2943
rect 111 2937 115 2938
rect 327 2942 331 2943
rect 327 2937 331 2938
rect 447 2942 451 2943
rect 447 2937 451 2938
rect 503 2942 507 2943
rect 503 2937 507 2938
rect 575 2942 579 2943
rect 575 2937 579 2938
rect 591 2942 595 2943
rect 591 2937 595 2938
rect 679 2942 683 2943
rect 679 2937 683 2938
rect 711 2942 715 2943
rect 711 2937 715 2938
rect 767 2942 771 2943
rect 767 2937 771 2938
rect 847 2942 851 2943
rect 847 2937 851 2938
rect 855 2942 859 2943
rect 855 2937 859 2938
rect 943 2942 947 2943
rect 943 2937 947 2938
rect 975 2942 979 2943
rect 975 2937 979 2938
rect 1031 2942 1035 2943
rect 1031 2937 1035 2938
rect 1103 2942 1107 2943
rect 1103 2937 1107 2938
rect 1119 2942 1123 2943
rect 1119 2937 1123 2938
rect 1207 2942 1211 2943
rect 1207 2937 1211 2938
rect 1231 2942 1235 2943
rect 1231 2937 1235 2938
rect 1295 2942 1299 2943
rect 1295 2937 1299 2938
rect 1359 2942 1363 2943
rect 1359 2937 1363 2938
rect 1495 2942 1499 2943
rect 1495 2937 1499 2938
rect 1767 2942 1771 2943
rect 1808 2939 1810 2967
rect 1832 2939 1834 2968
rect 1920 2939 1922 2968
rect 2032 2939 2034 2968
rect 2144 2939 2146 2968
rect 2248 2939 2250 2968
rect 2360 2939 2362 2968
rect 2480 2939 2482 2968
rect 2624 2939 2626 2968
rect 2792 2939 2794 2968
rect 2984 2939 2986 2968
rect 3184 2939 3186 2968
rect 3368 2939 3370 2968
rect 3462 2967 3468 2968
rect 3464 2939 3466 2967
rect 1767 2937 1771 2938
rect 1807 2938 1811 2939
rect 112 2921 114 2937
rect 110 2920 116 2921
rect 328 2920 330 2937
rect 448 2920 450 2937
rect 576 2920 578 2937
rect 712 2920 714 2937
rect 848 2920 850 2937
rect 976 2920 978 2937
rect 1104 2920 1106 2937
rect 1232 2920 1234 2937
rect 1360 2920 1362 2937
rect 1496 2920 1498 2937
rect 1768 2921 1770 2937
rect 1807 2933 1811 2934
rect 1831 2938 1835 2939
rect 1831 2933 1835 2934
rect 1919 2938 1923 2939
rect 1919 2933 1923 2934
rect 2015 2938 2019 2939
rect 2015 2933 2019 2934
rect 2031 2938 2035 2939
rect 2031 2933 2035 2934
rect 2143 2938 2147 2939
rect 2143 2933 2147 2934
rect 2215 2938 2219 2939
rect 2215 2933 2219 2934
rect 2247 2938 2251 2939
rect 2247 2933 2251 2934
rect 2359 2938 2363 2939
rect 2359 2933 2363 2934
rect 2407 2938 2411 2939
rect 2407 2933 2411 2934
rect 2479 2938 2483 2939
rect 2479 2933 2483 2934
rect 2591 2938 2595 2939
rect 2591 2933 2595 2934
rect 2623 2938 2627 2939
rect 2623 2933 2627 2934
rect 2759 2938 2763 2939
rect 2759 2933 2763 2934
rect 2791 2938 2795 2939
rect 2791 2933 2795 2934
rect 2911 2938 2915 2939
rect 2911 2933 2915 2934
rect 2983 2938 2987 2939
rect 2983 2933 2987 2934
rect 3063 2938 3067 2939
rect 3063 2933 3067 2934
rect 3183 2938 3187 2939
rect 3183 2933 3187 2934
rect 3207 2938 3211 2939
rect 3207 2933 3211 2934
rect 3359 2938 3363 2939
rect 3359 2933 3363 2934
rect 3367 2938 3371 2939
rect 3367 2933 3371 2934
rect 3463 2938 3467 2939
rect 3463 2933 3467 2934
rect 1766 2920 1772 2921
rect 110 2916 111 2920
rect 115 2916 116 2920
rect 110 2915 116 2916
rect 326 2919 332 2920
rect 326 2915 327 2919
rect 331 2915 332 2919
rect 326 2914 332 2915
rect 446 2919 452 2920
rect 446 2915 447 2919
rect 451 2915 452 2919
rect 446 2914 452 2915
rect 574 2919 580 2920
rect 574 2915 575 2919
rect 579 2915 580 2919
rect 574 2914 580 2915
rect 710 2919 716 2920
rect 710 2915 711 2919
rect 715 2915 716 2919
rect 710 2914 716 2915
rect 846 2919 852 2920
rect 846 2915 847 2919
rect 851 2915 852 2919
rect 846 2914 852 2915
rect 974 2919 980 2920
rect 974 2915 975 2919
rect 979 2915 980 2919
rect 974 2914 980 2915
rect 1102 2919 1108 2920
rect 1102 2915 1103 2919
rect 1107 2915 1108 2919
rect 1102 2914 1108 2915
rect 1230 2919 1236 2920
rect 1230 2915 1231 2919
rect 1235 2915 1236 2919
rect 1230 2914 1236 2915
rect 1358 2919 1364 2920
rect 1358 2915 1359 2919
rect 1363 2915 1364 2919
rect 1358 2914 1364 2915
rect 1494 2919 1500 2920
rect 1494 2915 1495 2919
rect 1499 2915 1500 2919
rect 1766 2916 1767 2920
rect 1771 2916 1772 2920
rect 1808 2917 1810 2933
rect 1766 2915 1772 2916
rect 1806 2916 1812 2917
rect 1832 2916 1834 2933
rect 2016 2916 2018 2933
rect 2216 2916 2218 2933
rect 2408 2916 2410 2933
rect 2592 2916 2594 2933
rect 2760 2916 2762 2933
rect 2912 2916 2914 2933
rect 3064 2916 3066 2933
rect 3208 2916 3210 2933
rect 3360 2916 3362 2933
rect 3464 2917 3466 2933
rect 3462 2916 3468 2917
rect 1494 2914 1500 2915
rect 1806 2912 1807 2916
rect 1811 2912 1812 2916
rect 1806 2911 1812 2912
rect 1830 2915 1836 2916
rect 1830 2911 1831 2915
rect 1835 2911 1836 2915
rect 1830 2910 1836 2911
rect 2014 2915 2020 2916
rect 2014 2911 2015 2915
rect 2019 2911 2020 2915
rect 2014 2910 2020 2911
rect 2214 2915 2220 2916
rect 2214 2911 2215 2915
rect 2219 2911 2220 2915
rect 2214 2910 2220 2911
rect 2406 2915 2412 2916
rect 2406 2911 2407 2915
rect 2411 2911 2412 2915
rect 2406 2910 2412 2911
rect 2590 2915 2596 2916
rect 2590 2911 2591 2915
rect 2595 2911 2596 2915
rect 2590 2910 2596 2911
rect 2758 2915 2764 2916
rect 2758 2911 2759 2915
rect 2763 2911 2764 2915
rect 2758 2910 2764 2911
rect 2910 2915 2916 2916
rect 2910 2911 2911 2915
rect 2915 2911 2916 2915
rect 2910 2910 2916 2911
rect 3062 2915 3068 2916
rect 3062 2911 3063 2915
rect 3067 2911 3068 2915
rect 3062 2910 3068 2911
rect 3206 2915 3212 2916
rect 3206 2911 3207 2915
rect 3211 2911 3212 2915
rect 3206 2910 3212 2911
rect 3358 2915 3364 2916
rect 3358 2911 3359 2915
rect 3363 2911 3364 2915
rect 3462 2912 3463 2916
rect 3467 2912 3468 2916
rect 3462 2911 3468 2912
rect 3358 2910 3364 2911
rect 110 2903 116 2904
rect 110 2899 111 2903
rect 115 2899 116 2903
rect 1766 2903 1772 2904
rect 110 2898 116 2899
rect 326 2900 332 2901
rect 112 2871 114 2898
rect 326 2896 327 2900
rect 331 2896 332 2900
rect 326 2895 332 2896
rect 446 2900 452 2901
rect 446 2896 447 2900
rect 451 2896 452 2900
rect 446 2895 452 2896
rect 574 2900 580 2901
rect 574 2896 575 2900
rect 579 2896 580 2900
rect 574 2895 580 2896
rect 710 2900 716 2901
rect 710 2896 711 2900
rect 715 2896 716 2900
rect 710 2895 716 2896
rect 846 2900 852 2901
rect 846 2896 847 2900
rect 851 2896 852 2900
rect 846 2895 852 2896
rect 974 2900 980 2901
rect 974 2896 975 2900
rect 979 2896 980 2900
rect 974 2895 980 2896
rect 1102 2900 1108 2901
rect 1102 2896 1103 2900
rect 1107 2896 1108 2900
rect 1102 2895 1108 2896
rect 1230 2900 1236 2901
rect 1230 2896 1231 2900
rect 1235 2896 1236 2900
rect 1230 2895 1236 2896
rect 1358 2900 1364 2901
rect 1358 2896 1359 2900
rect 1363 2896 1364 2900
rect 1358 2895 1364 2896
rect 1494 2900 1500 2901
rect 1494 2896 1495 2900
rect 1499 2896 1500 2900
rect 1766 2899 1767 2903
rect 1771 2899 1772 2903
rect 1766 2898 1772 2899
rect 1806 2899 1812 2900
rect 1494 2895 1500 2896
rect 328 2871 330 2895
rect 448 2871 450 2895
rect 576 2871 578 2895
rect 712 2871 714 2895
rect 848 2871 850 2895
rect 976 2871 978 2895
rect 1104 2871 1106 2895
rect 1232 2871 1234 2895
rect 1360 2871 1362 2895
rect 1496 2871 1498 2895
rect 1768 2871 1770 2898
rect 1806 2895 1807 2899
rect 1811 2895 1812 2899
rect 3462 2899 3468 2900
rect 1806 2894 1812 2895
rect 1830 2896 1836 2897
rect 1808 2875 1810 2894
rect 1830 2892 1831 2896
rect 1835 2892 1836 2896
rect 1830 2891 1836 2892
rect 2014 2896 2020 2897
rect 2014 2892 2015 2896
rect 2019 2892 2020 2896
rect 2014 2891 2020 2892
rect 2214 2896 2220 2897
rect 2214 2892 2215 2896
rect 2219 2892 2220 2896
rect 2214 2891 2220 2892
rect 2406 2896 2412 2897
rect 2406 2892 2407 2896
rect 2411 2892 2412 2896
rect 2406 2891 2412 2892
rect 2590 2896 2596 2897
rect 2590 2892 2591 2896
rect 2595 2892 2596 2896
rect 2590 2891 2596 2892
rect 2758 2896 2764 2897
rect 2758 2892 2759 2896
rect 2763 2892 2764 2896
rect 2758 2891 2764 2892
rect 2910 2896 2916 2897
rect 2910 2892 2911 2896
rect 2915 2892 2916 2896
rect 2910 2891 2916 2892
rect 3062 2896 3068 2897
rect 3062 2892 3063 2896
rect 3067 2892 3068 2896
rect 3062 2891 3068 2892
rect 3206 2896 3212 2897
rect 3206 2892 3207 2896
rect 3211 2892 3212 2896
rect 3206 2891 3212 2892
rect 3358 2896 3364 2897
rect 3358 2892 3359 2896
rect 3363 2892 3364 2896
rect 3462 2895 3463 2899
rect 3467 2895 3468 2899
rect 3462 2894 3468 2895
rect 3358 2891 3364 2892
rect 1832 2875 1834 2891
rect 2016 2875 2018 2891
rect 2216 2875 2218 2891
rect 2408 2875 2410 2891
rect 2592 2875 2594 2891
rect 2760 2875 2762 2891
rect 2912 2875 2914 2891
rect 3064 2875 3066 2891
rect 3208 2875 3210 2891
rect 3360 2875 3362 2891
rect 3464 2875 3466 2894
rect 1807 2874 1811 2875
rect 111 2870 115 2871
rect 111 2865 115 2866
rect 135 2870 139 2871
rect 135 2865 139 2866
rect 255 2870 259 2871
rect 255 2865 259 2866
rect 327 2870 331 2871
rect 327 2865 331 2866
rect 415 2870 419 2871
rect 415 2865 419 2866
rect 447 2870 451 2871
rect 447 2865 451 2866
rect 575 2870 579 2871
rect 575 2865 579 2866
rect 711 2870 715 2871
rect 711 2865 715 2866
rect 735 2870 739 2871
rect 735 2865 739 2866
rect 847 2870 851 2871
rect 847 2865 851 2866
rect 895 2870 899 2871
rect 895 2865 899 2866
rect 975 2870 979 2871
rect 975 2865 979 2866
rect 1047 2870 1051 2871
rect 1047 2865 1051 2866
rect 1103 2870 1107 2871
rect 1103 2865 1107 2866
rect 1191 2870 1195 2871
rect 1191 2865 1195 2866
rect 1231 2870 1235 2871
rect 1231 2865 1235 2866
rect 1343 2870 1347 2871
rect 1343 2865 1347 2866
rect 1359 2870 1363 2871
rect 1359 2865 1363 2866
rect 1495 2870 1499 2871
rect 1495 2865 1499 2866
rect 1767 2870 1771 2871
rect 1807 2869 1811 2870
rect 1831 2874 1835 2875
rect 1831 2869 1835 2870
rect 1999 2874 2003 2875
rect 1999 2869 2003 2870
rect 2015 2874 2019 2875
rect 2015 2869 2019 2870
rect 2191 2874 2195 2875
rect 2191 2869 2195 2870
rect 2215 2874 2219 2875
rect 2215 2869 2219 2870
rect 2383 2874 2387 2875
rect 2383 2869 2387 2870
rect 2407 2874 2411 2875
rect 2407 2869 2411 2870
rect 2567 2874 2571 2875
rect 2567 2869 2571 2870
rect 2591 2874 2595 2875
rect 2591 2869 2595 2870
rect 2735 2874 2739 2875
rect 2735 2869 2739 2870
rect 2759 2874 2763 2875
rect 2759 2869 2763 2870
rect 2903 2874 2907 2875
rect 2903 2869 2907 2870
rect 2911 2874 2915 2875
rect 2911 2869 2915 2870
rect 3063 2874 3067 2875
rect 3063 2869 3067 2870
rect 3207 2874 3211 2875
rect 3207 2869 3211 2870
rect 3223 2874 3227 2875
rect 3223 2869 3227 2870
rect 3359 2874 3363 2875
rect 3359 2869 3363 2870
rect 3367 2874 3371 2875
rect 3367 2869 3371 2870
rect 3463 2874 3467 2875
rect 3463 2869 3467 2870
rect 1767 2865 1771 2866
rect 112 2846 114 2865
rect 136 2849 138 2865
rect 256 2849 258 2865
rect 416 2849 418 2865
rect 576 2849 578 2865
rect 736 2849 738 2865
rect 896 2849 898 2865
rect 1048 2849 1050 2865
rect 1192 2849 1194 2865
rect 1344 2849 1346 2865
rect 1496 2849 1498 2865
rect 134 2848 140 2849
rect 110 2845 116 2846
rect 110 2841 111 2845
rect 115 2841 116 2845
rect 134 2844 135 2848
rect 139 2844 140 2848
rect 134 2843 140 2844
rect 254 2848 260 2849
rect 254 2844 255 2848
rect 259 2844 260 2848
rect 254 2843 260 2844
rect 414 2848 420 2849
rect 414 2844 415 2848
rect 419 2844 420 2848
rect 414 2843 420 2844
rect 574 2848 580 2849
rect 574 2844 575 2848
rect 579 2844 580 2848
rect 574 2843 580 2844
rect 734 2848 740 2849
rect 734 2844 735 2848
rect 739 2844 740 2848
rect 734 2843 740 2844
rect 894 2848 900 2849
rect 894 2844 895 2848
rect 899 2844 900 2848
rect 894 2843 900 2844
rect 1046 2848 1052 2849
rect 1046 2844 1047 2848
rect 1051 2844 1052 2848
rect 1046 2843 1052 2844
rect 1190 2848 1196 2849
rect 1190 2844 1191 2848
rect 1195 2844 1196 2848
rect 1190 2843 1196 2844
rect 1342 2848 1348 2849
rect 1342 2844 1343 2848
rect 1347 2844 1348 2848
rect 1342 2843 1348 2844
rect 1494 2848 1500 2849
rect 1494 2844 1495 2848
rect 1499 2844 1500 2848
rect 1768 2846 1770 2865
rect 1808 2850 1810 2869
rect 1832 2853 1834 2869
rect 2000 2853 2002 2869
rect 2192 2853 2194 2869
rect 2384 2853 2386 2869
rect 2568 2853 2570 2869
rect 2736 2853 2738 2869
rect 2904 2853 2906 2869
rect 3064 2853 3066 2869
rect 3224 2853 3226 2869
rect 3368 2853 3370 2869
rect 1830 2852 1836 2853
rect 1806 2849 1812 2850
rect 1494 2843 1500 2844
rect 1766 2845 1772 2846
rect 110 2840 116 2841
rect 1766 2841 1767 2845
rect 1771 2841 1772 2845
rect 1806 2845 1807 2849
rect 1811 2845 1812 2849
rect 1830 2848 1831 2852
rect 1835 2848 1836 2852
rect 1830 2847 1836 2848
rect 1998 2852 2004 2853
rect 1998 2848 1999 2852
rect 2003 2848 2004 2852
rect 1998 2847 2004 2848
rect 2190 2852 2196 2853
rect 2190 2848 2191 2852
rect 2195 2848 2196 2852
rect 2190 2847 2196 2848
rect 2382 2852 2388 2853
rect 2382 2848 2383 2852
rect 2387 2848 2388 2852
rect 2382 2847 2388 2848
rect 2566 2852 2572 2853
rect 2566 2848 2567 2852
rect 2571 2848 2572 2852
rect 2566 2847 2572 2848
rect 2734 2852 2740 2853
rect 2734 2848 2735 2852
rect 2739 2848 2740 2852
rect 2734 2847 2740 2848
rect 2902 2852 2908 2853
rect 2902 2848 2903 2852
rect 2907 2848 2908 2852
rect 2902 2847 2908 2848
rect 3062 2852 3068 2853
rect 3062 2848 3063 2852
rect 3067 2848 3068 2852
rect 3062 2847 3068 2848
rect 3222 2852 3228 2853
rect 3222 2848 3223 2852
rect 3227 2848 3228 2852
rect 3222 2847 3228 2848
rect 3366 2852 3372 2853
rect 3366 2848 3367 2852
rect 3371 2848 3372 2852
rect 3464 2850 3466 2869
rect 3366 2847 3372 2848
rect 3462 2849 3468 2850
rect 1806 2844 1812 2845
rect 3462 2845 3463 2849
rect 3467 2845 3468 2849
rect 3462 2844 3468 2845
rect 1766 2840 1772 2841
rect 1830 2833 1836 2834
rect 1806 2832 1812 2833
rect 134 2829 140 2830
rect 110 2828 116 2829
rect 110 2824 111 2828
rect 115 2824 116 2828
rect 134 2825 135 2829
rect 139 2825 140 2829
rect 134 2824 140 2825
rect 254 2829 260 2830
rect 254 2825 255 2829
rect 259 2825 260 2829
rect 254 2824 260 2825
rect 414 2829 420 2830
rect 414 2825 415 2829
rect 419 2825 420 2829
rect 414 2824 420 2825
rect 574 2829 580 2830
rect 574 2825 575 2829
rect 579 2825 580 2829
rect 574 2824 580 2825
rect 734 2829 740 2830
rect 734 2825 735 2829
rect 739 2825 740 2829
rect 734 2824 740 2825
rect 894 2829 900 2830
rect 894 2825 895 2829
rect 899 2825 900 2829
rect 894 2824 900 2825
rect 1046 2829 1052 2830
rect 1046 2825 1047 2829
rect 1051 2825 1052 2829
rect 1046 2824 1052 2825
rect 1190 2829 1196 2830
rect 1190 2825 1191 2829
rect 1195 2825 1196 2829
rect 1190 2824 1196 2825
rect 1342 2829 1348 2830
rect 1342 2825 1343 2829
rect 1347 2825 1348 2829
rect 1342 2824 1348 2825
rect 1494 2829 1500 2830
rect 1494 2825 1495 2829
rect 1499 2825 1500 2829
rect 1494 2824 1500 2825
rect 1766 2828 1772 2829
rect 1766 2824 1767 2828
rect 1771 2824 1772 2828
rect 1806 2828 1807 2832
rect 1811 2828 1812 2832
rect 1830 2829 1831 2833
rect 1835 2829 1836 2833
rect 1830 2828 1836 2829
rect 1998 2833 2004 2834
rect 1998 2829 1999 2833
rect 2003 2829 2004 2833
rect 1998 2828 2004 2829
rect 2190 2833 2196 2834
rect 2190 2829 2191 2833
rect 2195 2829 2196 2833
rect 2190 2828 2196 2829
rect 2382 2833 2388 2834
rect 2382 2829 2383 2833
rect 2387 2829 2388 2833
rect 2382 2828 2388 2829
rect 2566 2833 2572 2834
rect 2566 2829 2567 2833
rect 2571 2829 2572 2833
rect 2566 2828 2572 2829
rect 2734 2833 2740 2834
rect 2734 2829 2735 2833
rect 2739 2829 2740 2833
rect 2734 2828 2740 2829
rect 2902 2833 2908 2834
rect 2902 2829 2903 2833
rect 2907 2829 2908 2833
rect 2902 2828 2908 2829
rect 3062 2833 3068 2834
rect 3062 2829 3063 2833
rect 3067 2829 3068 2833
rect 3062 2828 3068 2829
rect 3222 2833 3228 2834
rect 3222 2829 3223 2833
rect 3227 2829 3228 2833
rect 3222 2828 3228 2829
rect 3366 2833 3372 2834
rect 3366 2829 3367 2833
rect 3371 2829 3372 2833
rect 3366 2828 3372 2829
rect 3462 2832 3468 2833
rect 3462 2828 3463 2832
rect 3467 2828 3468 2832
rect 1806 2827 1812 2828
rect 110 2823 116 2824
rect 112 2795 114 2823
rect 136 2795 138 2824
rect 256 2795 258 2824
rect 416 2795 418 2824
rect 576 2795 578 2824
rect 736 2795 738 2824
rect 896 2795 898 2824
rect 1048 2795 1050 2824
rect 1192 2795 1194 2824
rect 1344 2795 1346 2824
rect 1496 2795 1498 2824
rect 1766 2823 1772 2824
rect 1768 2795 1770 2823
rect 1808 2807 1810 2827
rect 1832 2807 1834 2828
rect 2000 2807 2002 2828
rect 2192 2807 2194 2828
rect 2384 2807 2386 2828
rect 2568 2807 2570 2828
rect 2736 2807 2738 2828
rect 2904 2807 2906 2828
rect 3064 2807 3066 2828
rect 3224 2807 3226 2828
rect 3368 2807 3370 2828
rect 3462 2827 3468 2828
rect 3464 2807 3466 2827
rect 1807 2806 1811 2807
rect 1807 2801 1811 2802
rect 1831 2806 1835 2807
rect 1831 2801 1835 2802
rect 1999 2806 2003 2807
rect 1999 2801 2003 2802
rect 2015 2806 2019 2807
rect 2015 2801 2019 2802
rect 2191 2806 2195 2807
rect 2191 2801 2195 2802
rect 2215 2806 2219 2807
rect 2215 2801 2219 2802
rect 2383 2806 2387 2807
rect 2383 2801 2387 2802
rect 2407 2806 2411 2807
rect 2407 2801 2411 2802
rect 2567 2806 2571 2807
rect 2567 2801 2571 2802
rect 2583 2806 2587 2807
rect 2583 2801 2587 2802
rect 2735 2806 2739 2807
rect 2735 2801 2739 2802
rect 2751 2806 2755 2807
rect 2751 2801 2755 2802
rect 2903 2806 2907 2807
rect 2903 2801 2907 2802
rect 2911 2806 2915 2807
rect 2911 2801 2915 2802
rect 3063 2806 3067 2807
rect 3063 2801 3067 2802
rect 3071 2806 3075 2807
rect 3071 2801 3075 2802
rect 3223 2806 3227 2807
rect 3223 2801 3227 2802
rect 3231 2806 3235 2807
rect 3231 2801 3235 2802
rect 3367 2806 3371 2807
rect 3367 2801 3371 2802
rect 3463 2806 3467 2807
rect 3463 2801 3467 2802
rect 111 2794 115 2795
rect 111 2789 115 2790
rect 135 2794 139 2795
rect 135 2789 139 2790
rect 247 2794 251 2795
rect 247 2789 251 2790
rect 255 2794 259 2795
rect 255 2789 259 2790
rect 391 2794 395 2795
rect 391 2789 395 2790
rect 415 2794 419 2795
rect 415 2789 419 2790
rect 543 2794 547 2795
rect 543 2789 547 2790
rect 575 2794 579 2795
rect 575 2789 579 2790
rect 695 2794 699 2795
rect 695 2789 699 2790
rect 735 2794 739 2795
rect 735 2789 739 2790
rect 855 2794 859 2795
rect 855 2789 859 2790
rect 895 2794 899 2795
rect 895 2789 899 2790
rect 1023 2794 1027 2795
rect 1023 2789 1027 2790
rect 1047 2794 1051 2795
rect 1047 2789 1051 2790
rect 1191 2794 1195 2795
rect 1191 2789 1195 2790
rect 1343 2794 1347 2795
rect 1343 2789 1347 2790
rect 1359 2794 1363 2795
rect 1359 2789 1363 2790
rect 1495 2794 1499 2795
rect 1495 2789 1499 2790
rect 1527 2794 1531 2795
rect 1527 2789 1531 2790
rect 1671 2794 1675 2795
rect 1671 2789 1675 2790
rect 1767 2794 1771 2795
rect 1767 2789 1771 2790
rect 112 2773 114 2789
rect 110 2772 116 2773
rect 136 2772 138 2789
rect 248 2772 250 2789
rect 392 2772 394 2789
rect 544 2772 546 2789
rect 696 2772 698 2789
rect 856 2772 858 2789
rect 1024 2772 1026 2789
rect 1192 2772 1194 2789
rect 1360 2772 1362 2789
rect 1528 2772 1530 2789
rect 1672 2772 1674 2789
rect 1768 2773 1770 2789
rect 1808 2785 1810 2801
rect 1806 2784 1812 2785
rect 1832 2784 1834 2801
rect 2016 2784 2018 2801
rect 2216 2784 2218 2801
rect 2408 2784 2410 2801
rect 2584 2784 2586 2801
rect 2752 2784 2754 2801
rect 2912 2784 2914 2801
rect 3072 2784 3074 2801
rect 3232 2784 3234 2801
rect 3368 2784 3370 2801
rect 3464 2785 3466 2801
rect 3462 2784 3468 2785
rect 1806 2780 1807 2784
rect 1811 2780 1812 2784
rect 1806 2779 1812 2780
rect 1830 2783 1836 2784
rect 1830 2779 1831 2783
rect 1835 2779 1836 2783
rect 1830 2778 1836 2779
rect 2014 2783 2020 2784
rect 2014 2779 2015 2783
rect 2019 2779 2020 2783
rect 2014 2778 2020 2779
rect 2214 2783 2220 2784
rect 2214 2779 2215 2783
rect 2219 2779 2220 2783
rect 2214 2778 2220 2779
rect 2406 2783 2412 2784
rect 2406 2779 2407 2783
rect 2411 2779 2412 2783
rect 2406 2778 2412 2779
rect 2582 2783 2588 2784
rect 2582 2779 2583 2783
rect 2587 2779 2588 2783
rect 2582 2778 2588 2779
rect 2750 2783 2756 2784
rect 2750 2779 2751 2783
rect 2755 2779 2756 2783
rect 2750 2778 2756 2779
rect 2910 2783 2916 2784
rect 2910 2779 2911 2783
rect 2915 2779 2916 2783
rect 2910 2778 2916 2779
rect 3070 2783 3076 2784
rect 3070 2779 3071 2783
rect 3075 2779 3076 2783
rect 3070 2778 3076 2779
rect 3230 2783 3236 2784
rect 3230 2779 3231 2783
rect 3235 2779 3236 2783
rect 3230 2778 3236 2779
rect 3366 2783 3372 2784
rect 3366 2779 3367 2783
rect 3371 2779 3372 2783
rect 3462 2780 3463 2784
rect 3467 2780 3468 2784
rect 3462 2779 3468 2780
rect 3366 2778 3372 2779
rect 1766 2772 1772 2773
rect 110 2768 111 2772
rect 115 2768 116 2772
rect 110 2767 116 2768
rect 134 2771 140 2772
rect 134 2767 135 2771
rect 139 2767 140 2771
rect 134 2766 140 2767
rect 246 2771 252 2772
rect 246 2767 247 2771
rect 251 2767 252 2771
rect 246 2766 252 2767
rect 390 2771 396 2772
rect 390 2767 391 2771
rect 395 2767 396 2771
rect 390 2766 396 2767
rect 542 2771 548 2772
rect 542 2767 543 2771
rect 547 2767 548 2771
rect 542 2766 548 2767
rect 694 2771 700 2772
rect 694 2767 695 2771
rect 699 2767 700 2771
rect 694 2766 700 2767
rect 854 2771 860 2772
rect 854 2767 855 2771
rect 859 2767 860 2771
rect 854 2766 860 2767
rect 1022 2771 1028 2772
rect 1022 2767 1023 2771
rect 1027 2767 1028 2771
rect 1022 2766 1028 2767
rect 1190 2771 1196 2772
rect 1190 2767 1191 2771
rect 1195 2767 1196 2771
rect 1190 2766 1196 2767
rect 1358 2771 1364 2772
rect 1358 2767 1359 2771
rect 1363 2767 1364 2771
rect 1358 2766 1364 2767
rect 1526 2771 1532 2772
rect 1526 2767 1527 2771
rect 1531 2767 1532 2771
rect 1526 2766 1532 2767
rect 1670 2771 1676 2772
rect 1670 2767 1671 2771
rect 1675 2767 1676 2771
rect 1766 2768 1767 2772
rect 1771 2768 1772 2772
rect 1766 2767 1772 2768
rect 1806 2767 1812 2768
rect 1670 2766 1676 2767
rect 1806 2763 1807 2767
rect 1811 2763 1812 2767
rect 3462 2767 3468 2768
rect 1806 2762 1812 2763
rect 1830 2764 1836 2765
rect 110 2755 116 2756
rect 110 2751 111 2755
rect 115 2751 116 2755
rect 1766 2755 1772 2756
rect 110 2750 116 2751
rect 134 2752 140 2753
rect 112 2723 114 2750
rect 134 2748 135 2752
rect 139 2748 140 2752
rect 134 2747 140 2748
rect 246 2752 252 2753
rect 246 2748 247 2752
rect 251 2748 252 2752
rect 246 2747 252 2748
rect 390 2752 396 2753
rect 390 2748 391 2752
rect 395 2748 396 2752
rect 390 2747 396 2748
rect 542 2752 548 2753
rect 542 2748 543 2752
rect 547 2748 548 2752
rect 542 2747 548 2748
rect 694 2752 700 2753
rect 694 2748 695 2752
rect 699 2748 700 2752
rect 694 2747 700 2748
rect 854 2752 860 2753
rect 854 2748 855 2752
rect 859 2748 860 2752
rect 854 2747 860 2748
rect 1022 2752 1028 2753
rect 1022 2748 1023 2752
rect 1027 2748 1028 2752
rect 1022 2747 1028 2748
rect 1190 2752 1196 2753
rect 1190 2748 1191 2752
rect 1195 2748 1196 2752
rect 1190 2747 1196 2748
rect 1358 2752 1364 2753
rect 1358 2748 1359 2752
rect 1363 2748 1364 2752
rect 1358 2747 1364 2748
rect 1526 2752 1532 2753
rect 1526 2748 1527 2752
rect 1531 2748 1532 2752
rect 1526 2747 1532 2748
rect 1670 2752 1676 2753
rect 1670 2748 1671 2752
rect 1675 2748 1676 2752
rect 1766 2751 1767 2755
rect 1771 2751 1772 2755
rect 1766 2750 1772 2751
rect 1670 2747 1676 2748
rect 136 2723 138 2747
rect 248 2723 250 2747
rect 392 2723 394 2747
rect 544 2723 546 2747
rect 696 2723 698 2747
rect 856 2723 858 2747
rect 1024 2723 1026 2747
rect 1192 2723 1194 2747
rect 1360 2723 1362 2747
rect 1528 2723 1530 2747
rect 1672 2723 1674 2747
rect 1768 2723 1770 2750
rect 1808 2727 1810 2762
rect 1830 2760 1831 2764
rect 1835 2760 1836 2764
rect 1830 2759 1836 2760
rect 2014 2764 2020 2765
rect 2014 2760 2015 2764
rect 2019 2760 2020 2764
rect 2014 2759 2020 2760
rect 2214 2764 2220 2765
rect 2214 2760 2215 2764
rect 2219 2760 2220 2764
rect 2214 2759 2220 2760
rect 2406 2764 2412 2765
rect 2406 2760 2407 2764
rect 2411 2760 2412 2764
rect 2406 2759 2412 2760
rect 2582 2764 2588 2765
rect 2582 2760 2583 2764
rect 2587 2760 2588 2764
rect 2582 2759 2588 2760
rect 2750 2764 2756 2765
rect 2750 2760 2751 2764
rect 2755 2760 2756 2764
rect 2750 2759 2756 2760
rect 2910 2764 2916 2765
rect 2910 2760 2911 2764
rect 2915 2760 2916 2764
rect 2910 2759 2916 2760
rect 3070 2764 3076 2765
rect 3070 2760 3071 2764
rect 3075 2760 3076 2764
rect 3070 2759 3076 2760
rect 3230 2764 3236 2765
rect 3230 2760 3231 2764
rect 3235 2760 3236 2764
rect 3230 2759 3236 2760
rect 3366 2764 3372 2765
rect 3366 2760 3367 2764
rect 3371 2760 3372 2764
rect 3462 2763 3463 2767
rect 3467 2763 3468 2767
rect 3462 2762 3468 2763
rect 3366 2759 3372 2760
rect 1832 2727 1834 2759
rect 2016 2727 2018 2759
rect 2216 2727 2218 2759
rect 2408 2727 2410 2759
rect 2584 2727 2586 2759
rect 2752 2727 2754 2759
rect 2912 2727 2914 2759
rect 3072 2727 3074 2759
rect 3232 2727 3234 2759
rect 3368 2727 3370 2759
rect 3464 2727 3466 2762
rect 1807 2726 1811 2727
rect 111 2722 115 2723
rect 111 2717 115 2718
rect 135 2722 139 2723
rect 135 2717 139 2718
rect 247 2722 251 2723
rect 247 2717 251 2718
rect 359 2722 363 2723
rect 359 2717 363 2718
rect 391 2722 395 2723
rect 391 2717 395 2718
rect 479 2722 483 2723
rect 479 2717 483 2718
rect 543 2722 547 2723
rect 543 2717 547 2718
rect 615 2722 619 2723
rect 615 2717 619 2718
rect 695 2722 699 2723
rect 695 2717 699 2718
rect 759 2722 763 2723
rect 759 2717 763 2718
rect 855 2722 859 2723
rect 855 2717 859 2718
rect 911 2722 915 2723
rect 911 2717 915 2718
rect 1023 2722 1027 2723
rect 1023 2717 1027 2718
rect 1063 2722 1067 2723
rect 1063 2717 1067 2718
rect 1191 2722 1195 2723
rect 1191 2717 1195 2718
rect 1215 2722 1219 2723
rect 1215 2717 1219 2718
rect 1359 2722 1363 2723
rect 1359 2717 1363 2718
rect 1375 2722 1379 2723
rect 1375 2717 1379 2718
rect 1527 2722 1531 2723
rect 1527 2717 1531 2718
rect 1535 2722 1539 2723
rect 1535 2717 1539 2718
rect 1671 2722 1675 2723
rect 1671 2717 1675 2718
rect 1767 2722 1771 2723
rect 1807 2721 1811 2722
rect 1831 2726 1835 2727
rect 1831 2721 1835 2722
rect 2015 2726 2019 2727
rect 2015 2721 2019 2722
rect 2039 2726 2043 2727
rect 2039 2721 2043 2722
rect 2159 2726 2163 2727
rect 2159 2721 2163 2722
rect 2215 2726 2219 2727
rect 2215 2721 2219 2722
rect 2279 2726 2283 2727
rect 2279 2721 2283 2722
rect 2407 2726 2411 2727
rect 2407 2721 2411 2722
rect 2543 2726 2547 2727
rect 2543 2721 2547 2722
rect 2583 2726 2587 2727
rect 2583 2721 2587 2722
rect 2687 2726 2691 2727
rect 2687 2721 2691 2722
rect 2751 2726 2755 2727
rect 2751 2721 2755 2722
rect 2847 2726 2851 2727
rect 2847 2721 2851 2722
rect 2911 2726 2915 2727
rect 2911 2721 2915 2722
rect 3023 2726 3027 2727
rect 3023 2721 3027 2722
rect 3071 2726 3075 2727
rect 3071 2721 3075 2722
rect 3207 2726 3211 2727
rect 3207 2721 3211 2722
rect 3231 2726 3235 2727
rect 3231 2721 3235 2722
rect 3367 2726 3371 2727
rect 3367 2721 3371 2722
rect 3463 2726 3467 2727
rect 3463 2721 3467 2722
rect 1767 2717 1771 2718
rect 112 2698 114 2717
rect 248 2701 250 2717
rect 360 2701 362 2717
rect 480 2701 482 2717
rect 616 2701 618 2717
rect 760 2701 762 2717
rect 912 2701 914 2717
rect 1064 2701 1066 2717
rect 1216 2701 1218 2717
rect 1376 2701 1378 2717
rect 1536 2701 1538 2717
rect 1672 2701 1674 2717
rect 246 2700 252 2701
rect 110 2697 116 2698
rect 110 2693 111 2697
rect 115 2693 116 2697
rect 246 2696 247 2700
rect 251 2696 252 2700
rect 246 2695 252 2696
rect 358 2700 364 2701
rect 358 2696 359 2700
rect 363 2696 364 2700
rect 358 2695 364 2696
rect 478 2700 484 2701
rect 478 2696 479 2700
rect 483 2696 484 2700
rect 478 2695 484 2696
rect 614 2700 620 2701
rect 614 2696 615 2700
rect 619 2696 620 2700
rect 614 2695 620 2696
rect 758 2700 764 2701
rect 758 2696 759 2700
rect 763 2696 764 2700
rect 758 2695 764 2696
rect 910 2700 916 2701
rect 910 2696 911 2700
rect 915 2696 916 2700
rect 910 2695 916 2696
rect 1062 2700 1068 2701
rect 1062 2696 1063 2700
rect 1067 2696 1068 2700
rect 1062 2695 1068 2696
rect 1214 2700 1220 2701
rect 1214 2696 1215 2700
rect 1219 2696 1220 2700
rect 1214 2695 1220 2696
rect 1374 2700 1380 2701
rect 1374 2696 1375 2700
rect 1379 2696 1380 2700
rect 1374 2695 1380 2696
rect 1534 2700 1540 2701
rect 1534 2696 1535 2700
rect 1539 2696 1540 2700
rect 1534 2695 1540 2696
rect 1670 2700 1676 2701
rect 1670 2696 1671 2700
rect 1675 2696 1676 2700
rect 1768 2698 1770 2717
rect 1808 2702 1810 2721
rect 2040 2705 2042 2721
rect 2160 2705 2162 2721
rect 2280 2705 2282 2721
rect 2408 2705 2410 2721
rect 2544 2705 2546 2721
rect 2688 2705 2690 2721
rect 2848 2705 2850 2721
rect 3024 2705 3026 2721
rect 3208 2705 3210 2721
rect 3368 2705 3370 2721
rect 2038 2704 2044 2705
rect 1806 2701 1812 2702
rect 1670 2695 1676 2696
rect 1766 2697 1772 2698
rect 110 2692 116 2693
rect 1766 2693 1767 2697
rect 1771 2693 1772 2697
rect 1806 2697 1807 2701
rect 1811 2697 1812 2701
rect 2038 2700 2039 2704
rect 2043 2700 2044 2704
rect 2038 2699 2044 2700
rect 2158 2704 2164 2705
rect 2158 2700 2159 2704
rect 2163 2700 2164 2704
rect 2158 2699 2164 2700
rect 2278 2704 2284 2705
rect 2278 2700 2279 2704
rect 2283 2700 2284 2704
rect 2278 2699 2284 2700
rect 2406 2704 2412 2705
rect 2406 2700 2407 2704
rect 2411 2700 2412 2704
rect 2406 2699 2412 2700
rect 2542 2704 2548 2705
rect 2542 2700 2543 2704
rect 2547 2700 2548 2704
rect 2542 2699 2548 2700
rect 2686 2704 2692 2705
rect 2686 2700 2687 2704
rect 2691 2700 2692 2704
rect 2686 2699 2692 2700
rect 2846 2704 2852 2705
rect 2846 2700 2847 2704
rect 2851 2700 2852 2704
rect 2846 2699 2852 2700
rect 3022 2704 3028 2705
rect 3022 2700 3023 2704
rect 3027 2700 3028 2704
rect 3022 2699 3028 2700
rect 3206 2704 3212 2705
rect 3206 2700 3207 2704
rect 3211 2700 3212 2704
rect 3206 2699 3212 2700
rect 3366 2704 3372 2705
rect 3366 2700 3367 2704
rect 3371 2700 3372 2704
rect 3464 2702 3466 2721
rect 3366 2699 3372 2700
rect 3462 2701 3468 2702
rect 1806 2696 1812 2697
rect 3462 2697 3463 2701
rect 3467 2697 3468 2701
rect 3462 2696 3468 2697
rect 1766 2692 1772 2693
rect 2038 2685 2044 2686
rect 1806 2684 1812 2685
rect 246 2681 252 2682
rect 110 2680 116 2681
rect 110 2676 111 2680
rect 115 2676 116 2680
rect 246 2677 247 2681
rect 251 2677 252 2681
rect 246 2676 252 2677
rect 358 2681 364 2682
rect 358 2677 359 2681
rect 363 2677 364 2681
rect 358 2676 364 2677
rect 478 2681 484 2682
rect 478 2677 479 2681
rect 483 2677 484 2681
rect 478 2676 484 2677
rect 614 2681 620 2682
rect 614 2677 615 2681
rect 619 2677 620 2681
rect 614 2676 620 2677
rect 758 2681 764 2682
rect 758 2677 759 2681
rect 763 2677 764 2681
rect 758 2676 764 2677
rect 910 2681 916 2682
rect 910 2677 911 2681
rect 915 2677 916 2681
rect 910 2676 916 2677
rect 1062 2681 1068 2682
rect 1062 2677 1063 2681
rect 1067 2677 1068 2681
rect 1062 2676 1068 2677
rect 1214 2681 1220 2682
rect 1214 2677 1215 2681
rect 1219 2677 1220 2681
rect 1214 2676 1220 2677
rect 1374 2681 1380 2682
rect 1374 2677 1375 2681
rect 1379 2677 1380 2681
rect 1374 2676 1380 2677
rect 1534 2681 1540 2682
rect 1534 2677 1535 2681
rect 1539 2677 1540 2681
rect 1534 2676 1540 2677
rect 1670 2681 1676 2682
rect 1670 2677 1671 2681
rect 1675 2677 1676 2681
rect 1670 2676 1676 2677
rect 1766 2680 1772 2681
rect 1766 2676 1767 2680
rect 1771 2676 1772 2680
rect 1806 2680 1807 2684
rect 1811 2680 1812 2684
rect 2038 2681 2039 2685
rect 2043 2681 2044 2685
rect 2038 2680 2044 2681
rect 2158 2685 2164 2686
rect 2158 2681 2159 2685
rect 2163 2681 2164 2685
rect 2158 2680 2164 2681
rect 2278 2685 2284 2686
rect 2278 2681 2279 2685
rect 2283 2681 2284 2685
rect 2278 2680 2284 2681
rect 2406 2685 2412 2686
rect 2406 2681 2407 2685
rect 2411 2681 2412 2685
rect 2406 2680 2412 2681
rect 2542 2685 2548 2686
rect 2542 2681 2543 2685
rect 2547 2681 2548 2685
rect 2542 2680 2548 2681
rect 2686 2685 2692 2686
rect 2686 2681 2687 2685
rect 2691 2681 2692 2685
rect 2686 2680 2692 2681
rect 2846 2685 2852 2686
rect 2846 2681 2847 2685
rect 2851 2681 2852 2685
rect 2846 2680 2852 2681
rect 3022 2685 3028 2686
rect 3022 2681 3023 2685
rect 3027 2681 3028 2685
rect 3022 2680 3028 2681
rect 3206 2685 3212 2686
rect 3206 2681 3207 2685
rect 3211 2681 3212 2685
rect 3206 2680 3212 2681
rect 3366 2685 3372 2686
rect 3366 2681 3367 2685
rect 3371 2681 3372 2685
rect 3366 2680 3372 2681
rect 3462 2684 3468 2685
rect 3462 2680 3463 2684
rect 3467 2680 3468 2684
rect 1806 2679 1812 2680
rect 110 2675 116 2676
rect 112 2651 114 2675
rect 248 2651 250 2676
rect 360 2651 362 2676
rect 480 2651 482 2676
rect 616 2651 618 2676
rect 760 2651 762 2676
rect 912 2651 914 2676
rect 1064 2651 1066 2676
rect 1216 2651 1218 2676
rect 1376 2651 1378 2676
rect 1536 2651 1538 2676
rect 1672 2651 1674 2676
rect 1766 2675 1772 2676
rect 1768 2651 1770 2675
rect 1808 2651 1810 2679
rect 2040 2651 2042 2680
rect 2160 2651 2162 2680
rect 2280 2651 2282 2680
rect 2408 2651 2410 2680
rect 2544 2651 2546 2680
rect 2688 2651 2690 2680
rect 2848 2651 2850 2680
rect 3024 2651 3026 2680
rect 3208 2651 3210 2680
rect 3368 2651 3370 2680
rect 3462 2679 3468 2680
rect 3464 2651 3466 2679
rect 111 2650 115 2651
rect 111 2645 115 2646
rect 247 2650 251 2651
rect 247 2645 251 2646
rect 359 2650 363 2651
rect 359 2645 363 2646
rect 463 2650 467 2651
rect 463 2645 467 2646
rect 479 2650 483 2651
rect 479 2645 483 2646
rect 551 2650 555 2651
rect 551 2645 555 2646
rect 615 2650 619 2651
rect 615 2645 619 2646
rect 639 2650 643 2651
rect 639 2645 643 2646
rect 743 2650 747 2651
rect 743 2645 747 2646
rect 759 2650 763 2651
rect 759 2645 763 2646
rect 855 2650 859 2651
rect 855 2645 859 2646
rect 911 2650 915 2651
rect 911 2645 915 2646
rect 983 2650 987 2651
rect 983 2645 987 2646
rect 1063 2650 1067 2651
rect 1063 2645 1067 2646
rect 1127 2650 1131 2651
rect 1127 2645 1131 2646
rect 1215 2650 1219 2651
rect 1215 2645 1219 2646
rect 1279 2650 1283 2651
rect 1279 2645 1283 2646
rect 1375 2650 1379 2651
rect 1375 2645 1379 2646
rect 1439 2650 1443 2651
rect 1439 2645 1443 2646
rect 1535 2650 1539 2651
rect 1535 2645 1539 2646
rect 1607 2650 1611 2651
rect 1607 2645 1611 2646
rect 1671 2650 1675 2651
rect 1671 2645 1675 2646
rect 1767 2650 1771 2651
rect 1767 2645 1771 2646
rect 1807 2650 1811 2651
rect 1807 2645 1811 2646
rect 1871 2650 1875 2651
rect 1871 2645 1875 2646
rect 1967 2650 1971 2651
rect 1967 2645 1971 2646
rect 2039 2650 2043 2651
rect 2039 2645 2043 2646
rect 2071 2650 2075 2651
rect 2071 2645 2075 2646
rect 2159 2650 2163 2651
rect 2159 2645 2163 2646
rect 2183 2650 2187 2651
rect 2183 2645 2187 2646
rect 2279 2650 2283 2651
rect 2279 2645 2283 2646
rect 2295 2650 2299 2651
rect 2295 2645 2299 2646
rect 2407 2650 2411 2651
rect 2407 2645 2411 2646
rect 2431 2650 2435 2651
rect 2431 2645 2435 2646
rect 2543 2650 2547 2651
rect 2543 2645 2547 2646
rect 2583 2650 2587 2651
rect 2583 2645 2587 2646
rect 2687 2650 2691 2651
rect 2687 2645 2691 2646
rect 2759 2650 2763 2651
rect 2759 2645 2763 2646
rect 2847 2650 2851 2651
rect 2847 2645 2851 2646
rect 2959 2650 2963 2651
rect 2959 2645 2963 2646
rect 3023 2650 3027 2651
rect 3023 2645 3027 2646
rect 3167 2650 3171 2651
rect 3167 2645 3171 2646
rect 3207 2650 3211 2651
rect 3207 2645 3211 2646
rect 3367 2650 3371 2651
rect 3367 2645 3371 2646
rect 3463 2650 3467 2651
rect 3463 2645 3467 2646
rect 112 2629 114 2645
rect 110 2628 116 2629
rect 464 2628 466 2645
rect 552 2628 554 2645
rect 640 2628 642 2645
rect 744 2628 746 2645
rect 856 2628 858 2645
rect 984 2628 986 2645
rect 1128 2628 1130 2645
rect 1280 2628 1282 2645
rect 1440 2628 1442 2645
rect 1608 2628 1610 2645
rect 1768 2629 1770 2645
rect 1808 2629 1810 2645
rect 1766 2628 1772 2629
rect 110 2624 111 2628
rect 115 2624 116 2628
rect 110 2623 116 2624
rect 462 2627 468 2628
rect 462 2623 463 2627
rect 467 2623 468 2627
rect 462 2622 468 2623
rect 550 2627 556 2628
rect 550 2623 551 2627
rect 555 2623 556 2627
rect 550 2622 556 2623
rect 638 2627 644 2628
rect 638 2623 639 2627
rect 643 2623 644 2627
rect 638 2622 644 2623
rect 742 2627 748 2628
rect 742 2623 743 2627
rect 747 2623 748 2627
rect 742 2622 748 2623
rect 854 2627 860 2628
rect 854 2623 855 2627
rect 859 2623 860 2627
rect 854 2622 860 2623
rect 982 2627 988 2628
rect 982 2623 983 2627
rect 987 2623 988 2627
rect 982 2622 988 2623
rect 1126 2627 1132 2628
rect 1126 2623 1127 2627
rect 1131 2623 1132 2627
rect 1126 2622 1132 2623
rect 1278 2627 1284 2628
rect 1278 2623 1279 2627
rect 1283 2623 1284 2627
rect 1278 2622 1284 2623
rect 1438 2627 1444 2628
rect 1438 2623 1439 2627
rect 1443 2623 1444 2627
rect 1438 2622 1444 2623
rect 1606 2627 1612 2628
rect 1606 2623 1607 2627
rect 1611 2623 1612 2627
rect 1766 2624 1767 2628
rect 1771 2624 1772 2628
rect 1766 2623 1772 2624
rect 1806 2628 1812 2629
rect 1872 2628 1874 2645
rect 1968 2628 1970 2645
rect 2072 2628 2074 2645
rect 2184 2628 2186 2645
rect 2296 2628 2298 2645
rect 2432 2628 2434 2645
rect 2584 2628 2586 2645
rect 2760 2628 2762 2645
rect 2960 2628 2962 2645
rect 3168 2628 3170 2645
rect 3368 2628 3370 2645
rect 3464 2629 3466 2645
rect 3462 2628 3468 2629
rect 1806 2624 1807 2628
rect 1811 2624 1812 2628
rect 1806 2623 1812 2624
rect 1870 2627 1876 2628
rect 1870 2623 1871 2627
rect 1875 2623 1876 2627
rect 1606 2622 1612 2623
rect 1870 2622 1876 2623
rect 1966 2627 1972 2628
rect 1966 2623 1967 2627
rect 1971 2623 1972 2627
rect 1966 2622 1972 2623
rect 2070 2627 2076 2628
rect 2070 2623 2071 2627
rect 2075 2623 2076 2627
rect 2070 2622 2076 2623
rect 2182 2627 2188 2628
rect 2182 2623 2183 2627
rect 2187 2623 2188 2627
rect 2182 2622 2188 2623
rect 2294 2627 2300 2628
rect 2294 2623 2295 2627
rect 2299 2623 2300 2627
rect 2294 2622 2300 2623
rect 2430 2627 2436 2628
rect 2430 2623 2431 2627
rect 2435 2623 2436 2627
rect 2430 2622 2436 2623
rect 2582 2627 2588 2628
rect 2582 2623 2583 2627
rect 2587 2623 2588 2627
rect 2582 2622 2588 2623
rect 2758 2627 2764 2628
rect 2758 2623 2759 2627
rect 2763 2623 2764 2627
rect 2758 2622 2764 2623
rect 2958 2627 2964 2628
rect 2958 2623 2959 2627
rect 2963 2623 2964 2627
rect 2958 2622 2964 2623
rect 3166 2627 3172 2628
rect 3166 2623 3167 2627
rect 3171 2623 3172 2627
rect 3166 2622 3172 2623
rect 3366 2627 3372 2628
rect 3366 2623 3367 2627
rect 3371 2623 3372 2627
rect 3462 2624 3463 2628
rect 3467 2624 3468 2628
rect 3462 2623 3468 2624
rect 3366 2622 3372 2623
rect 110 2611 116 2612
rect 110 2607 111 2611
rect 115 2607 116 2611
rect 1766 2611 1772 2612
rect 110 2606 116 2607
rect 462 2608 468 2609
rect 112 2579 114 2606
rect 462 2604 463 2608
rect 467 2604 468 2608
rect 462 2603 468 2604
rect 550 2608 556 2609
rect 550 2604 551 2608
rect 555 2604 556 2608
rect 550 2603 556 2604
rect 638 2608 644 2609
rect 638 2604 639 2608
rect 643 2604 644 2608
rect 638 2603 644 2604
rect 742 2608 748 2609
rect 742 2604 743 2608
rect 747 2604 748 2608
rect 742 2603 748 2604
rect 854 2608 860 2609
rect 854 2604 855 2608
rect 859 2604 860 2608
rect 854 2603 860 2604
rect 982 2608 988 2609
rect 982 2604 983 2608
rect 987 2604 988 2608
rect 982 2603 988 2604
rect 1126 2608 1132 2609
rect 1126 2604 1127 2608
rect 1131 2604 1132 2608
rect 1126 2603 1132 2604
rect 1278 2608 1284 2609
rect 1278 2604 1279 2608
rect 1283 2604 1284 2608
rect 1278 2603 1284 2604
rect 1438 2608 1444 2609
rect 1438 2604 1439 2608
rect 1443 2604 1444 2608
rect 1438 2603 1444 2604
rect 1606 2608 1612 2609
rect 1606 2604 1607 2608
rect 1611 2604 1612 2608
rect 1766 2607 1767 2611
rect 1771 2607 1772 2611
rect 1766 2606 1772 2607
rect 1806 2611 1812 2612
rect 1806 2607 1807 2611
rect 1811 2607 1812 2611
rect 3462 2611 3468 2612
rect 1806 2606 1812 2607
rect 1870 2608 1876 2609
rect 1606 2603 1612 2604
rect 464 2579 466 2603
rect 552 2579 554 2603
rect 640 2579 642 2603
rect 744 2579 746 2603
rect 856 2579 858 2603
rect 984 2579 986 2603
rect 1128 2579 1130 2603
rect 1280 2579 1282 2603
rect 1440 2579 1442 2603
rect 1608 2579 1610 2603
rect 1768 2579 1770 2606
rect 111 2578 115 2579
rect 111 2573 115 2574
rect 463 2578 467 2579
rect 463 2573 467 2574
rect 503 2578 507 2579
rect 503 2573 507 2574
rect 551 2578 555 2579
rect 551 2573 555 2574
rect 591 2578 595 2579
rect 591 2573 595 2574
rect 639 2578 643 2579
rect 639 2573 643 2574
rect 679 2578 683 2579
rect 679 2573 683 2574
rect 743 2578 747 2579
rect 743 2573 747 2574
rect 775 2578 779 2579
rect 775 2573 779 2574
rect 855 2578 859 2579
rect 855 2573 859 2574
rect 879 2578 883 2579
rect 879 2573 883 2574
rect 983 2578 987 2579
rect 983 2573 987 2574
rect 991 2578 995 2579
rect 991 2573 995 2574
rect 1103 2578 1107 2579
rect 1103 2573 1107 2574
rect 1127 2578 1131 2579
rect 1127 2573 1131 2574
rect 1223 2578 1227 2579
rect 1223 2573 1227 2574
rect 1279 2578 1283 2579
rect 1279 2573 1283 2574
rect 1351 2578 1355 2579
rect 1351 2573 1355 2574
rect 1439 2578 1443 2579
rect 1439 2573 1443 2574
rect 1479 2578 1483 2579
rect 1479 2573 1483 2574
rect 1607 2578 1611 2579
rect 1607 2573 1611 2574
rect 1767 2578 1771 2579
rect 1808 2575 1810 2606
rect 1870 2604 1871 2608
rect 1875 2604 1876 2608
rect 1870 2603 1876 2604
rect 1966 2608 1972 2609
rect 1966 2604 1967 2608
rect 1971 2604 1972 2608
rect 1966 2603 1972 2604
rect 2070 2608 2076 2609
rect 2070 2604 2071 2608
rect 2075 2604 2076 2608
rect 2070 2603 2076 2604
rect 2182 2608 2188 2609
rect 2182 2604 2183 2608
rect 2187 2604 2188 2608
rect 2182 2603 2188 2604
rect 2294 2608 2300 2609
rect 2294 2604 2295 2608
rect 2299 2604 2300 2608
rect 2294 2603 2300 2604
rect 2430 2608 2436 2609
rect 2430 2604 2431 2608
rect 2435 2604 2436 2608
rect 2430 2603 2436 2604
rect 2582 2608 2588 2609
rect 2582 2604 2583 2608
rect 2587 2604 2588 2608
rect 2582 2603 2588 2604
rect 2758 2608 2764 2609
rect 2758 2604 2759 2608
rect 2763 2604 2764 2608
rect 2758 2603 2764 2604
rect 2958 2608 2964 2609
rect 2958 2604 2959 2608
rect 2963 2604 2964 2608
rect 2958 2603 2964 2604
rect 3166 2608 3172 2609
rect 3166 2604 3167 2608
rect 3171 2604 3172 2608
rect 3166 2603 3172 2604
rect 3366 2608 3372 2609
rect 3366 2604 3367 2608
rect 3371 2604 3372 2608
rect 3462 2607 3463 2611
rect 3467 2607 3468 2611
rect 3462 2606 3468 2607
rect 3366 2603 3372 2604
rect 1872 2575 1874 2603
rect 1968 2575 1970 2603
rect 2072 2575 2074 2603
rect 2184 2575 2186 2603
rect 2296 2575 2298 2603
rect 2432 2575 2434 2603
rect 2584 2575 2586 2603
rect 2760 2575 2762 2603
rect 2960 2575 2962 2603
rect 3168 2575 3170 2603
rect 3368 2575 3370 2603
rect 3464 2575 3466 2606
rect 1767 2573 1771 2574
rect 1807 2574 1811 2575
rect 112 2554 114 2573
rect 504 2557 506 2573
rect 592 2557 594 2573
rect 680 2557 682 2573
rect 776 2557 778 2573
rect 880 2557 882 2573
rect 992 2557 994 2573
rect 1104 2557 1106 2573
rect 1224 2557 1226 2573
rect 1352 2557 1354 2573
rect 1480 2557 1482 2573
rect 1608 2557 1610 2573
rect 502 2556 508 2557
rect 110 2553 116 2554
rect 110 2549 111 2553
rect 115 2549 116 2553
rect 502 2552 503 2556
rect 507 2552 508 2556
rect 502 2551 508 2552
rect 590 2556 596 2557
rect 590 2552 591 2556
rect 595 2552 596 2556
rect 590 2551 596 2552
rect 678 2556 684 2557
rect 678 2552 679 2556
rect 683 2552 684 2556
rect 678 2551 684 2552
rect 774 2556 780 2557
rect 774 2552 775 2556
rect 779 2552 780 2556
rect 774 2551 780 2552
rect 878 2556 884 2557
rect 878 2552 879 2556
rect 883 2552 884 2556
rect 878 2551 884 2552
rect 990 2556 996 2557
rect 990 2552 991 2556
rect 995 2552 996 2556
rect 990 2551 996 2552
rect 1102 2556 1108 2557
rect 1102 2552 1103 2556
rect 1107 2552 1108 2556
rect 1102 2551 1108 2552
rect 1222 2556 1228 2557
rect 1222 2552 1223 2556
rect 1227 2552 1228 2556
rect 1222 2551 1228 2552
rect 1350 2556 1356 2557
rect 1350 2552 1351 2556
rect 1355 2552 1356 2556
rect 1350 2551 1356 2552
rect 1478 2556 1484 2557
rect 1478 2552 1479 2556
rect 1483 2552 1484 2556
rect 1478 2551 1484 2552
rect 1606 2556 1612 2557
rect 1606 2552 1607 2556
rect 1611 2552 1612 2556
rect 1768 2554 1770 2573
rect 1807 2569 1811 2570
rect 1831 2574 1835 2575
rect 1831 2569 1835 2570
rect 1871 2574 1875 2575
rect 1871 2569 1875 2570
rect 1919 2574 1923 2575
rect 1919 2569 1923 2570
rect 1967 2574 1971 2575
rect 1967 2569 1971 2570
rect 2007 2574 2011 2575
rect 2007 2569 2011 2570
rect 2071 2574 2075 2575
rect 2071 2569 2075 2570
rect 2111 2574 2115 2575
rect 2111 2569 2115 2570
rect 2183 2574 2187 2575
rect 2183 2569 2187 2570
rect 2223 2574 2227 2575
rect 2223 2569 2227 2570
rect 2295 2574 2299 2575
rect 2295 2569 2299 2570
rect 2343 2574 2347 2575
rect 2343 2569 2347 2570
rect 2431 2574 2435 2575
rect 2431 2569 2435 2570
rect 2487 2574 2491 2575
rect 2487 2569 2491 2570
rect 2583 2574 2587 2575
rect 2583 2569 2587 2570
rect 2647 2574 2651 2575
rect 2647 2569 2651 2570
rect 2759 2574 2763 2575
rect 2759 2569 2763 2570
rect 2815 2574 2819 2575
rect 2815 2569 2819 2570
rect 2959 2574 2963 2575
rect 2959 2569 2963 2570
rect 2999 2574 3003 2575
rect 2999 2569 3003 2570
rect 3167 2574 3171 2575
rect 3167 2569 3171 2570
rect 3191 2574 3195 2575
rect 3191 2569 3195 2570
rect 3367 2574 3371 2575
rect 3367 2569 3371 2570
rect 3463 2574 3467 2575
rect 3463 2569 3467 2570
rect 1606 2551 1612 2552
rect 1766 2553 1772 2554
rect 110 2548 116 2549
rect 1766 2549 1767 2553
rect 1771 2549 1772 2553
rect 1808 2550 1810 2569
rect 1832 2553 1834 2569
rect 1920 2553 1922 2569
rect 2008 2553 2010 2569
rect 2112 2553 2114 2569
rect 2224 2553 2226 2569
rect 2344 2553 2346 2569
rect 2488 2553 2490 2569
rect 2648 2553 2650 2569
rect 2816 2553 2818 2569
rect 3000 2553 3002 2569
rect 3192 2553 3194 2569
rect 3368 2553 3370 2569
rect 1830 2552 1836 2553
rect 1766 2548 1772 2549
rect 1806 2549 1812 2550
rect 1806 2545 1807 2549
rect 1811 2545 1812 2549
rect 1830 2548 1831 2552
rect 1835 2548 1836 2552
rect 1830 2547 1836 2548
rect 1918 2552 1924 2553
rect 1918 2548 1919 2552
rect 1923 2548 1924 2552
rect 1918 2547 1924 2548
rect 2006 2552 2012 2553
rect 2006 2548 2007 2552
rect 2011 2548 2012 2552
rect 2006 2547 2012 2548
rect 2110 2552 2116 2553
rect 2110 2548 2111 2552
rect 2115 2548 2116 2552
rect 2110 2547 2116 2548
rect 2222 2552 2228 2553
rect 2222 2548 2223 2552
rect 2227 2548 2228 2552
rect 2222 2547 2228 2548
rect 2342 2552 2348 2553
rect 2342 2548 2343 2552
rect 2347 2548 2348 2552
rect 2342 2547 2348 2548
rect 2486 2552 2492 2553
rect 2486 2548 2487 2552
rect 2491 2548 2492 2552
rect 2486 2547 2492 2548
rect 2646 2552 2652 2553
rect 2646 2548 2647 2552
rect 2651 2548 2652 2552
rect 2646 2547 2652 2548
rect 2814 2552 2820 2553
rect 2814 2548 2815 2552
rect 2819 2548 2820 2552
rect 2814 2547 2820 2548
rect 2998 2552 3004 2553
rect 2998 2548 2999 2552
rect 3003 2548 3004 2552
rect 2998 2547 3004 2548
rect 3190 2552 3196 2553
rect 3190 2548 3191 2552
rect 3195 2548 3196 2552
rect 3190 2547 3196 2548
rect 3366 2552 3372 2553
rect 3366 2548 3367 2552
rect 3371 2548 3372 2552
rect 3464 2550 3466 2569
rect 3366 2547 3372 2548
rect 3462 2549 3468 2550
rect 1806 2544 1812 2545
rect 3462 2545 3463 2549
rect 3467 2545 3468 2549
rect 3462 2544 3468 2545
rect 502 2537 508 2538
rect 110 2536 116 2537
rect 110 2532 111 2536
rect 115 2532 116 2536
rect 502 2533 503 2537
rect 507 2533 508 2537
rect 502 2532 508 2533
rect 590 2537 596 2538
rect 590 2533 591 2537
rect 595 2533 596 2537
rect 590 2532 596 2533
rect 678 2537 684 2538
rect 678 2533 679 2537
rect 683 2533 684 2537
rect 678 2532 684 2533
rect 774 2537 780 2538
rect 774 2533 775 2537
rect 779 2533 780 2537
rect 774 2532 780 2533
rect 878 2537 884 2538
rect 878 2533 879 2537
rect 883 2533 884 2537
rect 878 2532 884 2533
rect 990 2537 996 2538
rect 990 2533 991 2537
rect 995 2533 996 2537
rect 990 2532 996 2533
rect 1102 2537 1108 2538
rect 1102 2533 1103 2537
rect 1107 2533 1108 2537
rect 1102 2532 1108 2533
rect 1222 2537 1228 2538
rect 1222 2533 1223 2537
rect 1227 2533 1228 2537
rect 1222 2532 1228 2533
rect 1350 2537 1356 2538
rect 1350 2533 1351 2537
rect 1355 2533 1356 2537
rect 1350 2532 1356 2533
rect 1478 2537 1484 2538
rect 1478 2533 1479 2537
rect 1483 2533 1484 2537
rect 1478 2532 1484 2533
rect 1606 2537 1612 2538
rect 1606 2533 1607 2537
rect 1611 2533 1612 2537
rect 1606 2532 1612 2533
rect 1766 2536 1772 2537
rect 1766 2532 1767 2536
rect 1771 2532 1772 2536
rect 1830 2533 1836 2534
rect 110 2531 116 2532
rect 112 2507 114 2531
rect 504 2507 506 2532
rect 592 2507 594 2532
rect 680 2507 682 2532
rect 776 2507 778 2532
rect 880 2507 882 2532
rect 992 2507 994 2532
rect 1104 2507 1106 2532
rect 1224 2507 1226 2532
rect 1352 2507 1354 2532
rect 1480 2507 1482 2532
rect 1608 2507 1610 2532
rect 1766 2531 1772 2532
rect 1806 2532 1812 2533
rect 1768 2507 1770 2531
rect 1806 2528 1807 2532
rect 1811 2528 1812 2532
rect 1830 2529 1831 2533
rect 1835 2529 1836 2533
rect 1830 2528 1836 2529
rect 1918 2533 1924 2534
rect 1918 2529 1919 2533
rect 1923 2529 1924 2533
rect 1918 2528 1924 2529
rect 2006 2533 2012 2534
rect 2006 2529 2007 2533
rect 2011 2529 2012 2533
rect 2006 2528 2012 2529
rect 2110 2533 2116 2534
rect 2110 2529 2111 2533
rect 2115 2529 2116 2533
rect 2110 2528 2116 2529
rect 2222 2533 2228 2534
rect 2222 2529 2223 2533
rect 2227 2529 2228 2533
rect 2222 2528 2228 2529
rect 2342 2533 2348 2534
rect 2342 2529 2343 2533
rect 2347 2529 2348 2533
rect 2342 2528 2348 2529
rect 2486 2533 2492 2534
rect 2486 2529 2487 2533
rect 2491 2529 2492 2533
rect 2486 2528 2492 2529
rect 2646 2533 2652 2534
rect 2646 2529 2647 2533
rect 2651 2529 2652 2533
rect 2646 2528 2652 2529
rect 2814 2533 2820 2534
rect 2814 2529 2815 2533
rect 2819 2529 2820 2533
rect 2814 2528 2820 2529
rect 2998 2533 3004 2534
rect 2998 2529 2999 2533
rect 3003 2529 3004 2533
rect 2998 2528 3004 2529
rect 3190 2533 3196 2534
rect 3190 2529 3191 2533
rect 3195 2529 3196 2533
rect 3190 2528 3196 2529
rect 3366 2533 3372 2534
rect 3366 2529 3367 2533
rect 3371 2529 3372 2533
rect 3366 2528 3372 2529
rect 3462 2532 3468 2533
rect 3462 2528 3463 2532
rect 3467 2528 3468 2532
rect 1806 2527 1812 2528
rect 1808 2511 1810 2527
rect 1832 2511 1834 2528
rect 1920 2511 1922 2528
rect 2008 2511 2010 2528
rect 2112 2511 2114 2528
rect 2224 2511 2226 2528
rect 2344 2511 2346 2528
rect 2488 2511 2490 2528
rect 2648 2511 2650 2528
rect 2816 2511 2818 2528
rect 3000 2511 3002 2528
rect 3192 2511 3194 2528
rect 3368 2511 3370 2528
rect 3462 2527 3468 2528
rect 3464 2511 3466 2527
rect 1807 2510 1811 2511
rect 111 2506 115 2507
rect 111 2501 115 2502
rect 503 2506 507 2507
rect 503 2501 507 2502
rect 551 2506 555 2507
rect 551 2501 555 2502
rect 591 2506 595 2507
rect 591 2501 595 2502
rect 679 2506 683 2507
rect 679 2501 683 2502
rect 735 2506 739 2507
rect 735 2501 739 2502
rect 775 2506 779 2507
rect 775 2501 779 2502
rect 879 2506 883 2507
rect 879 2501 883 2502
rect 911 2506 915 2507
rect 911 2501 915 2502
rect 991 2506 995 2507
rect 991 2501 995 2502
rect 1079 2506 1083 2507
rect 1079 2501 1083 2502
rect 1103 2506 1107 2507
rect 1103 2501 1107 2502
rect 1223 2506 1227 2507
rect 1223 2501 1227 2502
rect 1239 2506 1243 2507
rect 1239 2501 1243 2502
rect 1351 2506 1355 2507
rect 1351 2501 1355 2502
rect 1399 2506 1403 2507
rect 1399 2501 1403 2502
rect 1479 2506 1483 2507
rect 1479 2501 1483 2502
rect 1567 2506 1571 2507
rect 1567 2501 1571 2502
rect 1607 2506 1611 2507
rect 1607 2501 1611 2502
rect 1767 2506 1771 2507
rect 1807 2505 1811 2506
rect 1831 2510 1835 2511
rect 1831 2505 1835 2506
rect 1919 2510 1923 2511
rect 1919 2505 1923 2506
rect 1951 2510 1955 2511
rect 1951 2505 1955 2506
rect 2007 2510 2011 2511
rect 2007 2505 2011 2506
rect 2039 2510 2043 2511
rect 2039 2505 2043 2506
rect 2111 2510 2115 2511
rect 2111 2505 2115 2506
rect 2135 2510 2139 2511
rect 2135 2505 2139 2506
rect 2223 2510 2227 2511
rect 2223 2505 2227 2506
rect 2239 2510 2243 2511
rect 2239 2505 2243 2506
rect 2343 2510 2347 2511
rect 2343 2505 2347 2506
rect 2367 2510 2371 2511
rect 2367 2505 2371 2506
rect 2487 2510 2491 2511
rect 2487 2505 2491 2506
rect 2527 2510 2531 2511
rect 2527 2505 2531 2506
rect 2647 2510 2651 2511
rect 2647 2505 2651 2506
rect 2711 2510 2715 2511
rect 2711 2505 2715 2506
rect 2815 2510 2819 2511
rect 2815 2505 2819 2506
rect 2919 2510 2923 2511
rect 2919 2505 2923 2506
rect 2999 2510 3003 2511
rect 2999 2505 3003 2506
rect 3143 2510 3147 2511
rect 3143 2505 3147 2506
rect 3191 2510 3195 2511
rect 3191 2505 3195 2506
rect 3367 2510 3371 2511
rect 3367 2505 3371 2506
rect 3463 2510 3467 2511
rect 3463 2505 3467 2506
rect 1767 2501 1771 2502
rect 112 2485 114 2501
rect 110 2484 116 2485
rect 552 2484 554 2501
rect 736 2484 738 2501
rect 912 2484 914 2501
rect 1080 2484 1082 2501
rect 1240 2484 1242 2501
rect 1400 2484 1402 2501
rect 1568 2484 1570 2501
rect 1768 2485 1770 2501
rect 1808 2489 1810 2505
rect 1806 2488 1812 2489
rect 1952 2488 1954 2505
rect 2040 2488 2042 2505
rect 2136 2488 2138 2505
rect 2240 2488 2242 2505
rect 2368 2488 2370 2505
rect 2528 2488 2530 2505
rect 2712 2488 2714 2505
rect 2920 2488 2922 2505
rect 3144 2488 3146 2505
rect 3368 2488 3370 2505
rect 3464 2489 3466 2505
rect 3462 2488 3468 2489
rect 1766 2484 1772 2485
rect 110 2480 111 2484
rect 115 2480 116 2484
rect 110 2479 116 2480
rect 550 2483 556 2484
rect 550 2479 551 2483
rect 555 2479 556 2483
rect 550 2478 556 2479
rect 734 2483 740 2484
rect 734 2479 735 2483
rect 739 2479 740 2483
rect 734 2478 740 2479
rect 910 2483 916 2484
rect 910 2479 911 2483
rect 915 2479 916 2483
rect 910 2478 916 2479
rect 1078 2483 1084 2484
rect 1078 2479 1079 2483
rect 1083 2479 1084 2483
rect 1078 2478 1084 2479
rect 1238 2483 1244 2484
rect 1238 2479 1239 2483
rect 1243 2479 1244 2483
rect 1238 2478 1244 2479
rect 1398 2483 1404 2484
rect 1398 2479 1399 2483
rect 1403 2479 1404 2483
rect 1398 2478 1404 2479
rect 1566 2483 1572 2484
rect 1566 2479 1567 2483
rect 1571 2479 1572 2483
rect 1766 2480 1767 2484
rect 1771 2480 1772 2484
rect 1806 2484 1807 2488
rect 1811 2484 1812 2488
rect 1806 2483 1812 2484
rect 1950 2487 1956 2488
rect 1950 2483 1951 2487
rect 1955 2483 1956 2487
rect 1950 2482 1956 2483
rect 2038 2487 2044 2488
rect 2038 2483 2039 2487
rect 2043 2483 2044 2487
rect 2038 2482 2044 2483
rect 2134 2487 2140 2488
rect 2134 2483 2135 2487
rect 2139 2483 2140 2487
rect 2134 2482 2140 2483
rect 2238 2487 2244 2488
rect 2238 2483 2239 2487
rect 2243 2483 2244 2487
rect 2238 2482 2244 2483
rect 2366 2487 2372 2488
rect 2366 2483 2367 2487
rect 2371 2483 2372 2487
rect 2366 2482 2372 2483
rect 2526 2487 2532 2488
rect 2526 2483 2527 2487
rect 2531 2483 2532 2487
rect 2526 2482 2532 2483
rect 2710 2487 2716 2488
rect 2710 2483 2711 2487
rect 2715 2483 2716 2487
rect 2710 2482 2716 2483
rect 2918 2487 2924 2488
rect 2918 2483 2919 2487
rect 2923 2483 2924 2487
rect 2918 2482 2924 2483
rect 3142 2487 3148 2488
rect 3142 2483 3143 2487
rect 3147 2483 3148 2487
rect 3142 2482 3148 2483
rect 3366 2487 3372 2488
rect 3366 2483 3367 2487
rect 3371 2483 3372 2487
rect 3462 2484 3463 2488
rect 3467 2484 3468 2488
rect 3462 2483 3468 2484
rect 3366 2482 3372 2483
rect 1766 2479 1772 2480
rect 1566 2478 1572 2479
rect 1806 2471 1812 2472
rect 110 2467 116 2468
rect 110 2463 111 2467
rect 115 2463 116 2467
rect 1766 2467 1772 2468
rect 110 2462 116 2463
rect 550 2464 556 2465
rect 112 2443 114 2462
rect 550 2460 551 2464
rect 555 2460 556 2464
rect 550 2459 556 2460
rect 734 2464 740 2465
rect 734 2460 735 2464
rect 739 2460 740 2464
rect 734 2459 740 2460
rect 910 2464 916 2465
rect 910 2460 911 2464
rect 915 2460 916 2464
rect 910 2459 916 2460
rect 1078 2464 1084 2465
rect 1078 2460 1079 2464
rect 1083 2460 1084 2464
rect 1078 2459 1084 2460
rect 1238 2464 1244 2465
rect 1238 2460 1239 2464
rect 1243 2460 1244 2464
rect 1238 2459 1244 2460
rect 1398 2464 1404 2465
rect 1398 2460 1399 2464
rect 1403 2460 1404 2464
rect 1398 2459 1404 2460
rect 1566 2464 1572 2465
rect 1566 2460 1567 2464
rect 1571 2460 1572 2464
rect 1766 2463 1767 2467
rect 1771 2463 1772 2467
rect 1806 2467 1807 2471
rect 1811 2467 1812 2471
rect 3462 2471 3468 2472
rect 1806 2466 1812 2467
rect 1950 2468 1956 2469
rect 1766 2462 1772 2463
rect 1566 2459 1572 2460
rect 552 2443 554 2459
rect 736 2443 738 2459
rect 912 2443 914 2459
rect 1080 2443 1082 2459
rect 1240 2443 1242 2459
rect 1400 2443 1402 2459
rect 1568 2443 1570 2459
rect 1768 2443 1770 2462
rect 111 2442 115 2443
rect 111 2437 115 2438
rect 415 2442 419 2443
rect 415 2437 419 2438
rect 503 2442 507 2443
rect 503 2437 507 2438
rect 551 2442 555 2443
rect 551 2437 555 2438
rect 599 2442 603 2443
rect 599 2437 603 2438
rect 703 2442 707 2443
rect 703 2437 707 2438
rect 735 2442 739 2443
rect 735 2437 739 2438
rect 807 2442 811 2443
rect 807 2437 811 2438
rect 911 2442 915 2443
rect 911 2437 915 2438
rect 919 2442 923 2443
rect 919 2437 923 2438
rect 1039 2442 1043 2443
rect 1039 2437 1043 2438
rect 1079 2442 1083 2443
rect 1079 2437 1083 2438
rect 1167 2442 1171 2443
rect 1167 2437 1171 2438
rect 1239 2442 1243 2443
rect 1239 2437 1243 2438
rect 1295 2442 1299 2443
rect 1295 2437 1299 2438
rect 1399 2442 1403 2443
rect 1399 2437 1403 2438
rect 1423 2442 1427 2443
rect 1423 2437 1427 2438
rect 1567 2442 1571 2443
rect 1567 2437 1571 2438
rect 1767 2442 1771 2443
rect 1808 2439 1810 2466
rect 1950 2464 1951 2468
rect 1955 2464 1956 2468
rect 1950 2463 1956 2464
rect 2038 2468 2044 2469
rect 2038 2464 2039 2468
rect 2043 2464 2044 2468
rect 2038 2463 2044 2464
rect 2134 2468 2140 2469
rect 2134 2464 2135 2468
rect 2139 2464 2140 2468
rect 2134 2463 2140 2464
rect 2238 2468 2244 2469
rect 2238 2464 2239 2468
rect 2243 2464 2244 2468
rect 2238 2463 2244 2464
rect 2366 2468 2372 2469
rect 2366 2464 2367 2468
rect 2371 2464 2372 2468
rect 2366 2463 2372 2464
rect 2526 2468 2532 2469
rect 2526 2464 2527 2468
rect 2531 2464 2532 2468
rect 2526 2463 2532 2464
rect 2710 2468 2716 2469
rect 2710 2464 2711 2468
rect 2715 2464 2716 2468
rect 2710 2463 2716 2464
rect 2918 2468 2924 2469
rect 2918 2464 2919 2468
rect 2923 2464 2924 2468
rect 2918 2463 2924 2464
rect 3142 2468 3148 2469
rect 3142 2464 3143 2468
rect 3147 2464 3148 2468
rect 3142 2463 3148 2464
rect 3366 2468 3372 2469
rect 3366 2464 3367 2468
rect 3371 2464 3372 2468
rect 3462 2467 3463 2471
rect 3467 2467 3468 2471
rect 3462 2466 3468 2467
rect 3366 2463 3372 2464
rect 1952 2439 1954 2463
rect 2040 2439 2042 2463
rect 2136 2439 2138 2463
rect 2240 2439 2242 2463
rect 2368 2439 2370 2463
rect 2528 2439 2530 2463
rect 2712 2439 2714 2463
rect 2920 2439 2922 2463
rect 3144 2439 3146 2463
rect 3368 2439 3370 2463
rect 3464 2439 3466 2466
rect 1767 2437 1771 2438
rect 1807 2438 1811 2439
rect 112 2418 114 2437
rect 416 2421 418 2437
rect 504 2421 506 2437
rect 600 2421 602 2437
rect 704 2421 706 2437
rect 808 2421 810 2437
rect 920 2421 922 2437
rect 1040 2421 1042 2437
rect 1168 2421 1170 2437
rect 1296 2421 1298 2437
rect 1424 2421 1426 2437
rect 414 2420 420 2421
rect 110 2417 116 2418
rect 110 2413 111 2417
rect 115 2413 116 2417
rect 414 2416 415 2420
rect 419 2416 420 2420
rect 414 2415 420 2416
rect 502 2420 508 2421
rect 502 2416 503 2420
rect 507 2416 508 2420
rect 502 2415 508 2416
rect 598 2420 604 2421
rect 598 2416 599 2420
rect 603 2416 604 2420
rect 598 2415 604 2416
rect 702 2420 708 2421
rect 702 2416 703 2420
rect 707 2416 708 2420
rect 702 2415 708 2416
rect 806 2420 812 2421
rect 806 2416 807 2420
rect 811 2416 812 2420
rect 806 2415 812 2416
rect 918 2420 924 2421
rect 918 2416 919 2420
rect 923 2416 924 2420
rect 918 2415 924 2416
rect 1038 2420 1044 2421
rect 1038 2416 1039 2420
rect 1043 2416 1044 2420
rect 1038 2415 1044 2416
rect 1166 2420 1172 2421
rect 1166 2416 1167 2420
rect 1171 2416 1172 2420
rect 1166 2415 1172 2416
rect 1294 2420 1300 2421
rect 1294 2416 1295 2420
rect 1299 2416 1300 2420
rect 1294 2415 1300 2416
rect 1422 2420 1428 2421
rect 1422 2416 1423 2420
rect 1427 2416 1428 2420
rect 1768 2418 1770 2437
rect 1807 2433 1811 2434
rect 1951 2438 1955 2439
rect 1951 2433 1955 2434
rect 2039 2438 2043 2439
rect 2039 2433 2043 2434
rect 2135 2438 2139 2439
rect 2135 2433 2139 2434
rect 2215 2438 2219 2439
rect 2215 2433 2219 2434
rect 2239 2438 2243 2439
rect 2239 2433 2243 2434
rect 2303 2438 2307 2439
rect 2303 2433 2307 2434
rect 2367 2438 2371 2439
rect 2367 2433 2371 2434
rect 2391 2438 2395 2439
rect 2391 2433 2395 2434
rect 2479 2438 2483 2439
rect 2479 2433 2483 2434
rect 2527 2438 2531 2439
rect 2527 2433 2531 2434
rect 2567 2438 2571 2439
rect 2567 2433 2571 2434
rect 2655 2438 2659 2439
rect 2655 2433 2659 2434
rect 2711 2438 2715 2439
rect 2711 2433 2715 2434
rect 2743 2438 2747 2439
rect 2743 2433 2747 2434
rect 2839 2438 2843 2439
rect 2839 2433 2843 2434
rect 2919 2438 2923 2439
rect 2919 2433 2923 2434
rect 2935 2438 2939 2439
rect 2935 2433 2939 2434
rect 3143 2438 3147 2439
rect 3143 2433 3147 2434
rect 3367 2438 3371 2439
rect 3367 2433 3371 2434
rect 3463 2438 3467 2439
rect 3463 2433 3467 2434
rect 1422 2415 1428 2416
rect 1766 2417 1772 2418
rect 110 2412 116 2413
rect 1766 2413 1767 2417
rect 1771 2413 1772 2417
rect 1808 2414 1810 2433
rect 2216 2417 2218 2433
rect 2304 2417 2306 2433
rect 2392 2417 2394 2433
rect 2480 2417 2482 2433
rect 2568 2417 2570 2433
rect 2656 2417 2658 2433
rect 2744 2417 2746 2433
rect 2840 2417 2842 2433
rect 2936 2417 2938 2433
rect 2214 2416 2220 2417
rect 1766 2412 1772 2413
rect 1806 2413 1812 2414
rect 1806 2409 1807 2413
rect 1811 2409 1812 2413
rect 2214 2412 2215 2416
rect 2219 2412 2220 2416
rect 2214 2411 2220 2412
rect 2302 2416 2308 2417
rect 2302 2412 2303 2416
rect 2307 2412 2308 2416
rect 2302 2411 2308 2412
rect 2390 2416 2396 2417
rect 2390 2412 2391 2416
rect 2395 2412 2396 2416
rect 2390 2411 2396 2412
rect 2478 2416 2484 2417
rect 2478 2412 2479 2416
rect 2483 2412 2484 2416
rect 2478 2411 2484 2412
rect 2566 2416 2572 2417
rect 2566 2412 2567 2416
rect 2571 2412 2572 2416
rect 2566 2411 2572 2412
rect 2654 2416 2660 2417
rect 2654 2412 2655 2416
rect 2659 2412 2660 2416
rect 2654 2411 2660 2412
rect 2742 2416 2748 2417
rect 2742 2412 2743 2416
rect 2747 2412 2748 2416
rect 2742 2411 2748 2412
rect 2838 2416 2844 2417
rect 2838 2412 2839 2416
rect 2843 2412 2844 2416
rect 2838 2411 2844 2412
rect 2934 2416 2940 2417
rect 2934 2412 2935 2416
rect 2939 2412 2940 2416
rect 3464 2414 3466 2433
rect 2934 2411 2940 2412
rect 3462 2413 3468 2414
rect 1806 2408 1812 2409
rect 3462 2409 3463 2413
rect 3467 2409 3468 2413
rect 3462 2408 3468 2409
rect 414 2401 420 2402
rect 110 2400 116 2401
rect 110 2396 111 2400
rect 115 2396 116 2400
rect 414 2397 415 2401
rect 419 2397 420 2401
rect 414 2396 420 2397
rect 502 2401 508 2402
rect 502 2397 503 2401
rect 507 2397 508 2401
rect 502 2396 508 2397
rect 598 2401 604 2402
rect 598 2397 599 2401
rect 603 2397 604 2401
rect 598 2396 604 2397
rect 702 2401 708 2402
rect 702 2397 703 2401
rect 707 2397 708 2401
rect 702 2396 708 2397
rect 806 2401 812 2402
rect 806 2397 807 2401
rect 811 2397 812 2401
rect 806 2396 812 2397
rect 918 2401 924 2402
rect 918 2397 919 2401
rect 923 2397 924 2401
rect 918 2396 924 2397
rect 1038 2401 1044 2402
rect 1038 2397 1039 2401
rect 1043 2397 1044 2401
rect 1038 2396 1044 2397
rect 1166 2401 1172 2402
rect 1166 2397 1167 2401
rect 1171 2397 1172 2401
rect 1166 2396 1172 2397
rect 1294 2401 1300 2402
rect 1294 2397 1295 2401
rect 1299 2397 1300 2401
rect 1294 2396 1300 2397
rect 1422 2401 1428 2402
rect 1422 2397 1423 2401
rect 1427 2397 1428 2401
rect 1422 2396 1428 2397
rect 1766 2400 1772 2401
rect 1766 2396 1767 2400
rect 1771 2396 1772 2400
rect 2214 2397 2220 2398
rect 110 2395 116 2396
rect 112 2375 114 2395
rect 416 2375 418 2396
rect 504 2375 506 2396
rect 600 2375 602 2396
rect 704 2375 706 2396
rect 808 2375 810 2396
rect 920 2375 922 2396
rect 1040 2375 1042 2396
rect 1168 2375 1170 2396
rect 1296 2375 1298 2396
rect 1424 2375 1426 2396
rect 1766 2395 1772 2396
rect 1806 2396 1812 2397
rect 1768 2375 1770 2395
rect 1806 2392 1807 2396
rect 1811 2392 1812 2396
rect 2214 2393 2215 2397
rect 2219 2393 2220 2397
rect 2214 2392 2220 2393
rect 2302 2397 2308 2398
rect 2302 2393 2303 2397
rect 2307 2393 2308 2397
rect 2302 2392 2308 2393
rect 2390 2397 2396 2398
rect 2390 2393 2391 2397
rect 2395 2393 2396 2397
rect 2390 2392 2396 2393
rect 2478 2397 2484 2398
rect 2478 2393 2479 2397
rect 2483 2393 2484 2397
rect 2478 2392 2484 2393
rect 2566 2397 2572 2398
rect 2566 2393 2567 2397
rect 2571 2393 2572 2397
rect 2566 2392 2572 2393
rect 2654 2397 2660 2398
rect 2654 2393 2655 2397
rect 2659 2393 2660 2397
rect 2654 2392 2660 2393
rect 2742 2397 2748 2398
rect 2742 2393 2743 2397
rect 2747 2393 2748 2397
rect 2742 2392 2748 2393
rect 2838 2397 2844 2398
rect 2838 2393 2839 2397
rect 2843 2393 2844 2397
rect 2838 2392 2844 2393
rect 2934 2397 2940 2398
rect 2934 2393 2935 2397
rect 2939 2393 2940 2397
rect 2934 2392 2940 2393
rect 3462 2396 3468 2397
rect 3462 2392 3463 2396
rect 3467 2392 3468 2396
rect 1806 2391 1812 2392
rect 1808 2375 1810 2391
rect 2216 2375 2218 2392
rect 2304 2375 2306 2392
rect 2392 2375 2394 2392
rect 2480 2375 2482 2392
rect 2568 2375 2570 2392
rect 2656 2375 2658 2392
rect 2744 2375 2746 2392
rect 2840 2375 2842 2392
rect 2936 2375 2938 2392
rect 3462 2391 3468 2392
rect 3464 2375 3466 2391
rect 111 2374 115 2375
rect 111 2369 115 2370
rect 319 2374 323 2375
rect 319 2369 323 2370
rect 415 2374 419 2375
rect 415 2369 419 2370
rect 431 2374 435 2375
rect 431 2369 435 2370
rect 503 2374 507 2375
rect 503 2369 507 2370
rect 543 2374 547 2375
rect 543 2369 547 2370
rect 599 2374 603 2375
rect 599 2369 603 2370
rect 655 2374 659 2375
rect 655 2369 659 2370
rect 703 2374 707 2375
rect 703 2369 707 2370
rect 767 2374 771 2375
rect 767 2369 771 2370
rect 807 2374 811 2375
rect 807 2369 811 2370
rect 879 2374 883 2375
rect 879 2369 883 2370
rect 919 2374 923 2375
rect 919 2369 923 2370
rect 991 2374 995 2375
rect 991 2369 995 2370
rect 1039 2374 1043 2375
rect 1039 2369 1043 2370
rect 1103 2374 1107 2375
rect 1103 2369 1107 2370
rect 1167 2374 1171 2375
rect 1167 2369 1171 2370
rect 1215 2374 1219 2375
rect 1215 2369 1219 2370
rect 1295 2374 1299 2375
rect 1295 2369 1299 2370
rect 1335 2374 1339 2375
rect 1335 2369 1339 2370
rect 1423 2374 1427 2375
rect 1423 2369 1427 2370
rect 1767 2374 1771 2375
rect 1767 2369 1771 2370
rect 1807 2374 1811 2375
rect 1807 2369 1811 2370
rect 2167 2374 2171 2375
rect 2167 2369 2171 2370
rect 2215 2374 2219 2375
rect 2215 2369 2219 2370
rect 2263 2374 2267 2375
rect 2263 2369 2267 2370
rect 2303 2374 2307 2375
rect 2303 2369 2307 2370
rect 2367 2374 2371 2375
rect 2367 2369 2371 2370
rect 2391 2374 2395 2375
rect 2391 2369 2395 2370
rect 2471 2374 2475 2375
rect 2471 2369 2475 2370
rect 2479 2374 2483 2375
rect 2479 2369 2483 2370
rect 2567 2374 2571 2375
rect 2567 2369 2571 2370
rect 2575 2374 2579 2375
rect 2575 2369 2579 2370
rect 2655 2374 2659 2375
rect 2655 2369 2659 2370
rect 2687 2374 2691 2375
rect 2687 2369 2691 2370
rect 2743 2374 2747 2375
rect 2743 2369 2747 2370
rect 2799 2374 2803 2375
rect 2799 2369 2803 2370
rect 2839 2374 2843 2375
rect 2839 2369 2843 2370
rect 2911 2374 2915 2375
rect 2911 2369 2915 2370
rect 2935 2374 2939 2375
rect 2935 2369 2939 2370
rect 3023 2374 3027 2375
rect 3023 2369 3027 2370
rect 3463 2374 3467 2375
rect 3463 2369 3467 2370
rect 112 2353 114 2369
rect 110 2352 116 2353
rect 320 2352 322 2369
rect 432 2352 434 2369
rect 544 2352 546 2369
rect 656 2352 658 2369
rect 768 2352 770 2369
rect 880 2352 882 2369
rect 992 2352 994 2369
rect 1104 2352 1106 2369
rect 1216 2352 1218 2369
rect 1336 2352 1338 2369
rect 1768 2353 1770 2369
rect 1808 2353 1810 2369
rect 1766 2352 1772 2353
rect 110 2348 111 2352
rect 115 2348 116 2352
rect 110 2347 116 2348
rect 318 2351 324 2352
rect 318 2347 319 2351
rect 323 2347 324 2351
rect 318 2346 324 2347
rect 430 2351 436 2352
rect 430 2347 431 2351
rect 435 2347 436 2351
rect 430 2346 436 2347
rect 542 2351 548 2352
rect 542 2347 543 2351
rect 547 2347 548 2351
rect 542 2346 548 2347
rect 654 2351 660 2352
rect 654 2347 655 2351
rect 659 2347 660 2351
rect 654 2346 660 2347
rect 766 2351 772 2352
rect 766 2347 767 2351
rect 771 2347 772 2351
rect 766 2346 772 2347
rect 878 2351 884 2352
rect 878 2347 879 2351
rect 883 2347 884 2351
rect 878 2346 884 2347
rect 990 2351 996 2352
rect 990 2347 991 2351
rect 995 2347 996 2351
rect 990 2346 996 2347
rect 1102 2351 1108 2352
rect 1102 2347 1103 2351
rect 1107 2347 1108 2351
rect 1102 2346 1108 2347
rect 1214 2351 1220 2352
rect 1214 2347 1215 2351
rect 1219 2347 1220 2351
rect 1214 2346 1220 2347
rect 1334 2351 1340 2352
rect 1334 2347 1335 2351
rect 1339 2347 1340 2351
rect 1766 2348 1767 2352
rect 1771 2348 1772 2352
rect 1766 2347 1772 2348
rect 1806 2352 1812 2353
rect 2168 2352 2170 2369
rect 2264 2352 2266 2369
rect 2368 2352 2370 2369
rect 2472 2352 2474 2369
rect 2576 2352 2578 2369
rect 2688 2352 2690 2369
rect 2800 2352 2802 2369
rect 2912 2352 2914 2369
rect 3024 2352 3026 2369
rect 3464 2353 3466 2369
rect 3462 2352 3468 2353
rect 1806 2348 1807 2352
rect 1811 2348 1812 2352
rect 1806 2347 1812 2348
rect 2166 2351 2172 2352
rect 2166 2347 2167 2351
rect 2171 2347 2172 2351
rect 1334 2346 1340 2347
rect 2166 2346 2172 2347
rect 2262 2351 2268 2352
rect 2262 2347 2263 2351
rect 2267 2347 2268 2351
rect 2262 2346 2268 2347
rect 2366 2351 2372 2352
rect 2366 2347 2367 2351
rect 2371 2347 2372 2351
rect 2366 2346 2372 2347
rect 2470 2351 2476 2352
rect 2470 2347 2471 2351
rect 2475 2347 2476 2351
rect 2470 2346 2476 2347
rect 2574 2351 2580 2352
rect 2574 2347 2575 2351
rect 2579 2347 2580 2351
rect 2574 2346 2580 2347
rect 2686 2351 2692 2352
rect 2686 2347 2687 2351
rect 2691 2347 2692 2351
rect 2686 2346 2692 2347
rect 2798 2351 2804 2352
rect 2798 2347 2799 2351
rect 2803 2347 2804 2351
rect 2798 2346 2804 2347
rect 2910 2351 2916 2352
rect 2910 2347 2911 2351
rect 2915 2347 2916 2351
rect 2910 2346 2916 2347
rect 3022 2351 3028 2352
rect 3022 2347 3023 2351
rect 3027 2347 3028 2351
rect 3462 2348 3463 2352
rect 3467 2348 3468 2352
rect 3462 2347 3468 2348
rect 3022 2346 3028 2347
rect 110 2335 116 2336
rect 110 2331 111 2335
rect 115 2331 116 2335
rect 1766 2335 1772 2336
rect 110 2330 116 2331
rect 318 2332 324 2333
rect 112 2303 114 2330
rect 318 2328 319 2332
rect 323 2328 324 2332
rect 318 2327 324 2328
rect 430 2332 436 2333
rect 430 2328 431 2332
rect 435 2328 436 2332
rect 430 2327 436 2328
rect 542 2332 548 2333
rect 542 2328 543 2332
rect 547 2328 548 2332
rect 542 2327 548 2328
rect 654 2332 660 2333
rect 654 2328 655 2332
rect 659 2328 660 2332
rect 654 2327 660 2328
rect 766 2332 772 2333
rect 766 2328 767 2332
rect 771 2328 772 2332
rect 766 2327 772 2328
rect 878 2332 884 2333
rect 878 2328 879 2332
rect 883 2328 884 2332
rect 878 2327 884 2328
rect 990 2332 996 2333
rect 990 2328 991 2332
rect 995 2328 996 2332
rect 990 2327 996 2328
rect 1102 2332 1108 2333
rect 1102 2328 1103 2332
rect 1107 2328 1108 2332
rect 1102 2327 1108 2328
rect 1214 2332 1220 2333
rect 1214 2328 1215 2332
rect 1219 2328 1220 2332
rect 1214 2327 1220 2328
rect 1334 2332 1340 2333
rect 1334 2328 1335 2332
rect 1339 2328 1340 2332
rect 1766 2331 1767 2335
rect 1771 2331 1772 2335
rect 1766 2330 1772 2331
rect 1806 2335 1812 2336
rect 1806 2331 1807 2335
rect 1811 2331 1812 2335
rect 3462 2335 3468 2336
rect 1806 2330 1812 2331
rect 2166 2332 2172 2333
rect 1334 2327 1340 2328
rect 320 2303 322 2327
rect 432 2303 434 2327
rect 544 2303 546 2327
rect 656 2303 658 2327
rect 768 2303 770 2327
rect 880 2303 882 2327
rect 992 2303 994 2327
rect 1104 2303 1106 2327
rect 1216 2303 1218 2327
rect 1336 2303 1338 2327
rect 1768 2303 1770 2330
rect 1808 2303 1810 2330
rect 2166 2328 2167 2332
rect 2171 2328 2172 2332
rect 2166 2327 2172 2328
rect 2262 2332 2268 2333
rect 2262 2328 2263 2332
rect 2267 2328 2268 2332
rect 2262 2327 2268 2328
rect 2366 2332 2372 2333
rect 2366 2328 2367 2332
rect 2371 2328 2372 2332
rect 2366 2327 2372 2328
rect 2470 2332 2476 2333
rect 2470 2328 2471 2332
rect 2475 2328 2476 2332
rect 2470 2327 2476 2328
rect 2574 2332 2580 2333
rect 2574 2328 2575 2332
rect 2579 2328 2580 2332
rect 2574 2327 2580 2328
rect 2686 2332 2692 2333
rect 2686 2328 2687 2332
rect 2691 2328 2692 2332
rect 2686 2327 2692 2328
rect 2798 2332 2804 2333
rect 2798 2328 2799 2332
rect 2803 2328 2804 2332
rect 2798 2327 2804 2328
rect 2910 2332 2916 2333
rect 2910 2328 2911 2332
rect 2915 2328 2916 2332
rect 2910 2327 2916 2328
rect 3022 2332 3028 2333
rect 3022 2328 3023 2332
rect 3027 2328 3028 2332
rect 3462 2331 3463 2335
rect 3467 2331 3468 2335
rect 3462 2330 3468 2331
rect 3022 2327 3028 2328
rect 2168 2303 2170 2327
rect 2264 2303 2266 2327
rect 2368 2303 2370 2327
rect 2472 2303 2474 2327
rect 2576 2303 2578 2327
rect 2688 2303 2690 2327
rect 2800 2303 2802 2327
rect 2912 2303 2914 2327
rect 3024 2303 3026 2327
rect 3464 2303 3466 2330
rect 111 2302 115 2303
rect 111 2297 115 2298
rect 151 2302 155 2303
rect 151 2297 155 2298
rect 271 2302 275 2303
rect 271 2297 275 2298
rect 319 2302 323 2303
rect 319 2297 323 2298
rect 391 2302 395 2303
rect 391 2297 395 2298
rect 431 2302 435 2303
rect 431 2297 435 2298
rect 519 2302 523 2303
rect 519 2297 523 2298
rect 543 2302 547 2303
rect 543 2297 547 2298
rect 647 2302 651 2303
rect 647 2297 651 2298
rect 655 2302 659 2303
rect 655 2297 659 2298
rect 767 2302 771 2303
rect 767 2297 771 2298
rect 775 2302 779 2303
rect 775 2297 779 2298
rect 879 2302 883 2303
rect 879 2297 883 2298
rect 895 2302 899 2303
rect 895 2297 899 2298
rect 991 2302 995 2303
rect 991 2297 995 2298
rect 1015 2302 1019 2303
rect 1015 2297 1019 2298
rect 1103 2302 1107 2303
rect 1103 2297 1107 2298
rect 1143 2302 1147 2303
rect 1143 2297 1147 2298
rect 1215 2302 1219 2303
rect 1215 2297 1219 2298
rect 1271 2302 1275 2303
rect 1271 2297 1275 2298
rect 1335 2302 1339 2303
rect 1335 2297 1339 2298
rect 1767 2302 1771 2303
rect 1767 2297 1771 2298
rect 1807 2302 1811 2303
rect 1807 2297 1811 2298
rect 1887 2302 1891 2303
rect 1887 2297 1891 2298
rect 2039 2302 2043 2303
rect 2039 2297 2043 2298
rect 2167 2302 2171 2303
rect 2167 2297 2171 2298
rect 2199 2302 2203 2303
rect 2199 2297 2203 2298
rect 2263 2302 2267 2303
rect 2263 2297 2267 2298
rect 2367 2302 2371 2303
rect 2367 2297 2371 2298
rect 2375 2302 2379 2303
rect 2375 2297 2379 2298
rect 2471 2302 2475 2303
rect 2471 2297 2475 2298
rect 2551 2302 2555 2303
rect 2551 2297 2555 2298
rect 2575 2302 2579 2303
rect 2575 2297 2579 2298
rect 2687 2302 2691 2303
rect 2687 2297 2691 2298
rect 2719 2302 2723 2303
rect 2719 2297 2723 2298
rect 2799 2302 2803 2303
rect 2799 2297 2803 2298
rect 2887 2302 2891 2303
rect 2887 2297 2891 2298
rect 2911 2302 2915 2303
rect 2911 2297 2915 2298
rect 3023 2302 3027 2303
rect 3023 2297 3027 2298
rect 3055 2302 3059 2303
rect 3055 2297 3059 2298
rect 3223 2302 3227 2303
rect 3223 2297 3227 2298
rect 3367 2302 3371 2303
rect 3367 2297 3371 2298
rect 3463 2302 3467 2303
rect 3463 2297 3467 2298
rect 112 2278 114 2297
rect 152 2281 154 2297
rect 272 2281 274 2297
rect 392 2281 394 2297
rect 520 2281 522 2297
rect 648 2281 650 2297
rect 776 2281 778 2297
rect 896 2281 898 2297
rect 1016 2281 1018 2297
rect 1144 2281 1146 2297
rect 1272 2281 1274 2297
rect 150 2280 156 2281
rect 110 2277 116 2278
rect 110 2273 111 2277
rect 115 2273 116 2277
rect 150 2276 151 2280
rect 155 2276 156 2280
rect 150 2275 156 2276
rect 270 2280 276 2281
rect 270 2276 271 2280
rect 275 2276 276 2280
rect 270 2275 276 2276
rect 390 2280 396 2281
rect 390 2276 391 2280
rect 395 2276 396 2280
rect 390 2275 396 2276
rect 518 2280 524 2281
rect 518 2276 519 2280
rect 523 2276 524 2280
rect 518 2275 524 2276
rect 646 2280 652 2281
rect 646 2276 647 2280
rect 651 2276 652 2280
rect 646 2275 652 2276
rect 774 2280 780 2281
rect 774 2276 775 2280
rect 779 2276 780 2280
rect 774 2275 780 2276
rect 894 2280 900 2281
rect 894 2276 895 2280
rect 899 2276 900 2280
rect 894 2275 900 2276
rect 1014 2280 1020 2281
rect 1014 2276 1015 2280
rect 1019 2276 1020 2280
rect 1014 2275 1020 2276
rect 1142 2280 1148 2281
rect 1142 2276 1143 2280
rect 1147 2276 1148 2280
rect 1142 2275 1148 2276
rect 1270 2280 1276 2281
rect 1270 2276 1271 2280
rect 1275 2276 1276 2280
rect 1768 2278 1770 2297
rect 1808 2278 1810 2297
rect 1888 2281 1890 2297
rect 2040 2281 2042 2297
rect 2200 2281 2202 2297
rect 2376 2281 2378 2297
rect 2552 2281 2554 2297
rect 2720 2281 2722 2297
rect 2888 2281 2890 2297
rect 3056 2281 3058 2297
rect 3224 2281 3226 2297
rect 3368 2281 3370 2297
rect 1886 2280 1892 2281
rect 1270 2275 1276 2276
rect 1766 2277 1772 2278
rect 110 2272 116 2273
rect 1766 2273 1767 2277
rect 1771 2273 1772 2277
rect 1766 2272 1772 2273
rect 1806 2277 1812 2278
rect 1806 2273 1807 2277
rect 1811 2273 1812 2277
rect 1886 2276 1887 2280
rect 1891 2276 1892 2280
rect 1886 2275 1892 2276
rect 2038 2280 2044 2281
rect 2038 2276 2039 2280
rect 2043 2276 2044 2280
rect 2038 2275 2044 2276
rect 2198 2280 2204 2281
rect 2198 2276 2199 2280
rect 2203 2276 2204 2280
rect 2198 2275 2204 2276
rect 2374 2280 2380 2281
rect 2374 2276 2375 2280
rect 2379 2276 2380 2280
rect 2374 2275 2380 2276
rect 2550 2280 2556 2281
rect 2550 2276 2551 2280
rect 2555 2276 2556 2280
rect 2550 2275 2556 2276
rect 2718 2280 2724 2281
rect 2718 2276 2719 2280
rect 2723 2276 2724 2280
rect 2718 2275 2724 2276
rect 2886 2280 2892 2281
rect 2886 2276 2887 2280
rect 2891 2276 2892 2280
rect 2886 2275 2892 2276
rect 3054 2280 3060 2281
rect 3054 2276 3055 2280
rect 3059 2276 3060 2280
rect 3054 2275 3060 2276
rect 3222 2280 3228 2281
rect 3222 2276 3223 2280
rect 3227 2276 3228 2280
rect 3222 2275 3228 2276
rect 3366 2280 3372 2281
rect 3366 2276 3367 2280
rect 3371 2276 3372 2280
rect 3464 2278 3466 2297
rect 3366 2275 3372 2276
rect 3462 2277 3468 2278
rect 1806 2272 1812 2273
rect 3462 2273 3463 2277
rect 3467 2273 3468 2277
rect 3462 2272 3468 2273
rect 150 2261 156 2262
rect 110 2260 116 2261
rect 110 2256 111 2260
rect 115 2256 116 2260
rect 150 2257 151 2261
rect 155 2257 156 2261
rect 150 2256 156 2257
rect 270 2261 276 2262
rect 270 2257 271 2261
rect 275 2257 276 2261
rect 270 2256 276 2257
rect 390 2261 396 2262
rect 390 2257 391 2261
rect 395 2257 396 2261
rect 390 2256 396 2257
rect 518 2261 524 2262
rect 518 2257 519 2261
rect 523 2257 524 2261
rect 518 2256 524 2257
rect 646 2261 652 2262
rect 646 2257 647 2261
rect 651 2257 652 2261
rect 646 2256 652 2257
rect 774 2261 780 2262
rect 774 2257 775 2261
rect 779 2257 780 2261
rect 774 2256 780 2257
rect 894 2261 900 2262
rect 894 2257 895 2261
rect 899 2257 900 2261
rect 894 2256 900 2257
rect 1014 2261 1020 2262
rect 1014 2257 1015 2261
rect 1019 2257 1020 2261
rect 1014 2256 1020 2257
rect 1142 2261 1148 2262
rect 1142 2257 1143 2261
rect 1147 2257 1148 2261
rect 1142 2256 1148 2257
rect 1270 2261 1276 2262
rect 1886 2261 1892 2262
rect 1270 2257 1271 2261
rect 1275 2257 1276 2261
rect 1270 2256 1276 2257
rect 1766 2260 1772 2261
rect 1766 2256 1767 2260
rect 1771 2256 1772 2260
rect 110 2255 116 2256
rect 112 2235 114 2255
rect 152 2235 154 2256
rect 272 2235 274 2256
rect 392 2235 394 2256
rect 520 2235 522 2256
rect 648 2235 650 2256
rect 776 2235 778 2256
rect 896 2235 898 2256
rect 1016 2235 1018 2256
rect 1144 2235 1146 2256
rect 1272 2235 1274 2256
rect 1766 2255 1772 2256
rect 1806 2260 1812 2261
rect 1806 2256 1807 2260
rect 1811 2256 1812 2260
rect 1886 2257 1887 2261
rect 1891 2257 1892 2261
rect 1886 2256 1892 2257
rect 2038 2261 2044 2262
rect 2038 2257 2039 2261
rect 2043 2257 2044 2261
rect 2038 2256 2044 2257
rect 2198 2261 2204 2262
rect 2198 2257 2199 2261
rect 2203 2257 2204 2261
rect 2198 2256 2204 2257
rect 2374 2261 2380 2262
rect 2374 2257 2375 2261
rect 2379 2257 2380 2261
rect 2374 2256 2380 2257
rect 2550 2261 2556 2262
rect 2550 2257 2551 2261
rect 2555 2257 2556 2261
rect 2550 2256 2556 2257
rect 2718 2261 2724 2262
rect 2718 2257 2719 2261
rect 2723 2257 2724 2261
rect 2718 2256 2724 2257
rect 2886 2261 2892 2262
rect 2886 2257 2887 2261
rect 2891 2257 2892 2261
rect 2886 2256 2892 2257
rect 3054 2261 3060 2262
rect 3054 2257 3055 2261
rect 3059 2257 3060 2261
rect 3054 2256 3060 2257
rect 3222 2261 3228 2262
rect 3222 2257 3223 2261
rect 3227 2257 3228 2261
rect 3222 2256 3228 2257
rect 3366 2261 3372 2262
rect 3366 2257 3367 2261
rect 3371 2257 3372 2261
rect 3366 2256 3372 2257
rect 3462 2260 3468 2261
rect 3462 2256 3463 2260
rect 3467 2256 3468 2260
rect 1806 2255 1812 2256
rect 1768 2235 1770 2255
rect 1808 2239 1810 2255
rect 1888 2239 1890 2256
rect 2040 2239 2042 2256
rect 2200 2239 2202 2256
rect 2376 2239 2378 2256
rect 2552 2239 2554 2256
rect 2720 2239 2722 2256
rect 2888 2239 2890 2256
rect 3056 2239 3058 2256
rect 3224 2239 3226 2256
rect 3368 2239 3370 2256
rect 3462 2255 3468 2256
rect 3464 2239 3466 2255
rect 1807 2238 1811 2239
rect 111 2234 115 2235
rect 111 2229 115 2230
rect 135 2234 139 2235
rect 135 2229 139 2230
rect 151 2234 155 2235
rect 151 2229 155 2230
rect 247 2234 251 2235
rect 247 2229 251 2230
rect 271 2234 275 2235
rect 271 2229 275 2230
rect 391 2234 395 2235
rect 391 2229 395 2230
rect 407 2234 411 2235
rect 407 2229 411 2230
rect 519 2234 523 2235
rect 519 2229 523 2230
rect 583 2234 587 2235
rect 583 2229 587 2230
rect 647 2234 651 2235
rect 647 2229 651 2230
rect 767 2234 771 2235
rect 767 2229 771 2230
rect 775 2234 779 2235
rect 775 2229 779 2230
rect 895 2234 899 2235
rect 895 2229 899 2230
rect 951 2234 955 2235
rect 951 2229 955 2230
rect 1015 2234 1019 2235
rect 1015 2229 1019 2230
rect 1135 2234 1139 2235
rect 1135 2229 1139 2230
rect 1143 2234 1147 2235
rect 1143 2229 1147 2230
rect 1271 2234 1275 2235
rect 1271 2229 1275 2230
rect 1319 2234 1323 2235
rect 1319 2229 1323 2230
rect 1503 2234 1507 2235
rect 1503 2229 1507 2230
rect 1671 2234 1675 2235
rect 1671 2229 1675 2230
rect 1767 2234 1771 2235
rect 1807 2233 1811 2234
rect 1831 2238 1835 2239
rect 1831 2233 1835 2234
rect 1887 2238 1891 2239
rect 1887 2233 1891 2234
rect 1967 2238 1971 2239
rect 1967 2233 1971 2234
rect 2039 2238 2043 2239
rect 2039 2233 2043 2234
rect 2135 2238 2139 2239
rect 2135 2233 2139 2234
rect 2199 2238 2203 2239
rect 2199 2233 2203 2234
rect 2311 2238 2315 2239
rect 2311 2233 2315 2234
rect 2375 2238 2379 2239
rect 2375 2233 2379 2234
rect 2487 2238 2491 2239
rect 2487 2233 2491 2234
rect 2551 2238 2555 2239
rect 2551 2233 2555 2234
rect 2655 2238 2659 2239
rect 2655 2233 2659 2234
rect 2719 2238 2723 2239
rect 2719 2233 2723 2234
rect 2815 2238 2819 2239
rect 2815 2233 2819 2234
rect 2887 2238 2891 2239
rect 2887 2233 2891 2234
rect 2959 2238 2963 2239
rect 2959 2233 2963 2234
rect 3055 2238 3059 2239
rect 3055 2233 3059 2234
rect 3103 2238 3107 2239
rect 3103 2233 3107 2234
rect 3223 2238 3227 2239
rect 3223 2233 3227 2234
rect 3247 2238 3251 2239
rect 3247 2233 3251 2234
rect 3367 2238 3371 2239
rect 3367 2233 3371 2234
rect 3463 2238 3467 2239
rect 3463 2233 3467 2234
rect 1767 2229 1771 2230
rect 112 2213 114 2229
rect 110 2212 116 2213
rect 136 2212 138 2229
rect 248 2212 250 2229
rect 408 2212 410 2229
rect 584 2212 586 2229
rect 768 2212 770 2229
rect 952 2212 954 2229
rect 1136 2212 1138 2229
rect 1320 2212 1322 2229
rect 1504 2212 1506 2229
rect 1672 2212 1674 2229
rect 1768 2213 1770 2229
rect 1808 2217 1810 2233
rect 1806 2216 1812 2217
rect 1832 2216 1834 2233
rect 1968 2216 1970 2233
rect 2136 2216 2138 2233
rect 2312 2216 2314 2233
rect 2488 2216 2490 2233
rect 2656 2216 2658 2233
rect 2816 2216 2818 2233
rect 2960 2216 2962 2233
rect 3104 2216 3106 2233
rect 3248 2216 3250 2233
rect 3368 2216 3370 2233
rect 3464 2217 3466 2233
rect 3462 2216 3468 2217
rect 1766 2212 1772 2213
rect 110 2208 111 2212
rect 115 2208 116 2212
rect 110 2207 116 2208
rect 134 2211 140 2212
rect 134 2207 135 2211
rect 139 2207 140 2211
rect 134 2206 140 2207
rect 246 2211 252 2212
rect 246 2207 247 2211
rect 251 2207 252 2211
rect 246 2206 252 2207
rect 406 2211 412 2212
rect 406 2207 407 2211
rect 411 2207 412 2211
rect 406 2206 412 2207
rect 582 2211 588 2212
rect 582 2207 583 2211
rect 587 2207 588 2211
rect 582 2206 588 2207
rect 766 2211 772 2212
rect 766 2207 767 2211
rect 771 2207 772 2211
rect 766 2206 772 2207
rect 950 2211 956 2212
rect 950 2207 951 2211
rect 955 2207 956 2211
rect 950 2206 956 2207
rect 1134 2211 1140 2212
rect 1134 2207 1135 2211
rect 1139 2207 1140 2211
rect 1134 2206 1140 2207
rect 1318 2211 1324 2212
rect 1318 2207 1319 2211
rect 1323 2207 1324 2211
rect 1318 2206 1324 2207
rect 1502 2211 1508 2212
rect 1502 2207 1503 2211
rect 1507 2207 1508 2211
rect 1502 2206 1508 2207
rect 1670 2211 1676 2212
rect 1670 2207 1671 2211
rect 1675 2207 1676 2211
rect 1766 2208 1767 2212
rect 1771 2208 1772 2212
rect 1806 2212 1807 2216
rect 1811 2212 1812 2216
rect 1806 2211 1812 2212
rect 1830 2215 1836 2216
rect 1830 2211 1831 2215
rect 1835 2211 1836 2215
rect 1830 2210 1836 2211
rect 1966 2215 1972 2216
rect 1966 2211 1967 2215
rect 1971 2211 1972 2215
rect 1966 2210 1972 2211
rect 2134 2215 2140 2216
rect 2134 2211 2135 2215
rect 2139 2211 2140 2215
rect 2134 2210 2140 2211
rect 2310 2215 2316 2216
rect 2310 2211 2311 2215
rect 2315 2211 2316 2215
rect 2310 2210 2316 2211
rect 2486 2215 2492 2216
rect 2486 2211 2487 2215
rect 2491 2211 2492 2215
rect 2486 2210 2492 2211
rect 2654 2215 2660 2216
rect 2654 2211 2655 2215
rect 2659 2211 2660 2215
rect 2654 2210 2660 2211
rect 2814 2215 2820 2216
rect 2814 2211 2815 2215
rect 2819 2211 2820 2215
rect 2814 2210 2820 2211
rect 2958 2215 2964 2216
rect 2958 2211 2959 2215
rect 2963 2211 2964 2215
rect 2958 2210 2964 2211
rect 3102 2215 3108 2216
rect 3102 2211 3103 2215
rect 3107 2211 3108 2215
rect 3102 2210 3108 2211
rect 3246 2215 3252 2216
rect 3246 2211 3247 2215
rect 3251 2211 3252 2215
rect 3246 2210 3252 2211
rect 3366 2215 3372 2216
rect 3366 2211 3367 2215
rect 3371 2211 3372 2215
rect 3462 2212 3463 2216
rect 3467 2212 3468 2216
rect 3462 2211 3468 2212
rect 3366 2210 3372 2211
rect 1766 2207 1772 2208
rect 1670 2206 1676 2207
rect 1806 2199 1812 2200
rect 110 2195 116 2196
rect 110 2191 111 2195
rect 115 2191 116 2195
rect 1766 2195 1772 2196
rect 110 2190 116 2191
rect 134 2192 140 2193
rect 112 2163 114 2190
rect 134 2188 135 2192
rect 139 2188 140 2192
rect 134 2187 140 2188
rect 246 2192 252 2193
rect 246 2188 247 2192
rect 251 2188 252 2192
rect 246 2187 252 2188
rect 406 2192 412 2193
rect 406 2188 407 2192
rect 411 2188 412 2192
rect 406 2187 412 2188
rect 582 2192 588 2193
rect 582 2188 583 2192
rect 587 2188 588 2192
rect 582 2187 588 2188
rect 766 2192 772 2193
rect 766 2188 767 2192
rect 771 2188 772 2192
rect 766 2187 772 2188
rect 950 2192 956 2193
rect 950 2188 951 2192
rect 955 2188 956 2192
rect 950 2187 956 2188
rect 1134 2192 1140 2193
rect 1134 2188 1135 2192
rect 1139 2188 1140 2192
rect 1134 2187 1140 2188
rect 1318 2192 1324 2193
rect 1318 2188 1319 2192
rect 1323 2188 1324 2192
rect 1318 2187 1324 2188
rect 1502 2192 1508 2193
rect 1502 2188 1503 2192
rect 1507 2188 1508 2192
rect 1502 2187 1508 2188
rect 1670 2192 1676 2193
rect 1670 2188 1671 2192
rect 1675 2188 1676 2192
rect 1766 2191 1767 2195
rect 1771 2191 1772 2195
rect 1806 2195 1807 2199
rect 1811 2195 1812 2199
rect 3462 2199 3468 2200
rect 1806 2194 1812 2195
rect 1830 2196 1836 2197
rect 1766 2190 1772 2191
rect 1670 2187 1676 2188
rect 136 2163 138 2187
rect 248 2163 250 2187
rect 408 2163 410 2187
rect 584 2163 586 2187
rect 768 2163 770 2187
rect 952 2163 954 2187
rect 1136 2163 1138 2187
rect 1320 2163 1322 2187
rect 1504 2163 1506 2187
rect 1672 2163 1674 2187
rect 1768 2163 1770 2190
rect 1808 2175 1810 2194
rect 1830 2192 1831 2196
rect 1835 2192 1836 2196
rect 1830 2191 1836 2192
rect 1966 2196 1972 2197
rect 1966 2192 1967 2196
rect 1971 2192 1972 2196
rect 1966 2191 1972 2192
rect 2134 2196 2140 2197
rect 2134 2192 2135 2196
rect 2139 2192 2140 2196
rect 2134 2191 2140 2192
rect 2310 2196 2316 2197
rect 2310 2192 2311 2196
rect 2315 2192 2316 2196
rect 2310 2191 2316 2192
rect 2486 2196 2492 2197
rect 2486 2192 2487 2196
rect 2491 2192 2492 2196
rect 2486 2191 2492 2192
rect 2654 2196 2660 2197
rect 2654 2192 2655 2196
rect 2659 2192 2660 2196
rect 2654 2191 2660 2192
rect 2814 2196 2820 2197
rect 2814 2192 2815 2196
rect 2819 2192 2820 2196
rect 2814 2191 2820 2192
rect 2958 2196 2964 2197
rect 2958 2192 2959 2196
rect 2963 2192 2964 2196
rect 2958 2191 2964 2192
rect 3102 2196 3108 2197
rect 3102 2192 3103 2196
rect 3107 2192 3108 2196
rect 3102 2191 3108 2192
rect 3246 2196 3252 2197
rect 3246 2192 3247 2196
rect 3251 2192 3252 2196
rect 3246 2191 3252 2192
rect 3366 2196 3372 2197
rect 3366 2192 3367 2196
rect 3371 2192 3372 2196
rect 3462 2195 3463 2199
rect 3467 2195 3468 2199
rect 3462 2194 3468 2195
rect 3366 2191 3372 2192
rect 1832 2175 1834 2191
rect 1968 2175 1970 2191
rect 2136 2175 2138 2191
rect 2312 2175 2314 2191
rect 2488 2175 2490 2191
rect 2656 2175 2658 2191
rect 2816 2175 2818 2191
rect 2960 2175 2962 2191
rect 3104 2175 3106 2191
rect 3248 2175 3250 2191
rect 3368 2175 3370 2191
rect 3464 2175 3466 2194
rect 1807 2174 1811 2175
rect 1807 2169 1811 2170
rect 1831 2174 1835 2175
rect 1831 2169 1835 2170
rect 1967 2174 1971 2175
rect 1967 2169 1971 2170
rect 2135 2174 2139 2175
rect 2135 2169 2139 2170
rect 2311 2174 2315 2175
rect 2311 2169 2315 2170
rect 2487 2174 2491 2175
rect 2487 2169 2491 2170
rect 2655 2174 2659 2175
rect 2655 2169 2659 2170
rect 2815 2174 2819 2175
rect 2815 2169 2819 2170
rect 2927 2174 2931 2175
rect 2927 2169 2931 2170
rect 2959 2174 2963 2175
rect 2959 2169 2963 2170
rect 3015 2174 3019 2175
rect 3015 2169 3019 2170
rect 3103 2174 3107 2175
rect 3103 2169 3107 2170
rect 3191 2174 3195 2175
rect 3191 2169 3195 2170
rect 3247 2174 3251 2175
rect 3247 2169 3251 2170
rect 3279 2174 3283 2175
rect 3279 2169 3283 2170
rect 3367 2174 3371 2175
rect 3367 2169 3371 2170
rect 3463 2174 3467 2175
rect 3463 2169 3467 2170
rect 111 2162 115 2163
rect 111 2157 115 2158
rect 135 2162 139 2163
rect 135 2157 139 2158
rect 247 2162 251 2163
rect 247 2157 251 2158
rect 391 2162 395 2163
rect 391 2157 395 2158
rect 407 2162 411 2163
rect 407 2157 411 2158
rect 543 2162 547 2163
rect 543 2157 547 2158
rect 583 2162 587 2163
rect 583 2157 587 2158
rect 695 2162 699 2163
rect 695 2157 699 2158
rect 767 2162 771 2163
rect 767 2157 771 2158
rect 839 2162 843 2163
rect 839 2157 843 2158
rect 951 2162 955 2163
rect 951 2157 955 2158
rect 975 2162 979 2163
rect 975 2157 979 2158
rect 1103 2162 1107 2163
rect 1103 2157 1107 2158
rect 1135 2162 1139 2163
rect 1135 2157 1139 2158
rect 1231 2162 1235 2163
rect 1231 2157 1235 2158
rect 1319 2162 1323 2163
rect 1319 2157 1323 2158
rect 1351 2162 1355 2163
rect 1351 2157 1355 2158
rect 1463 2162 1467 2163
rect 1463 2157 1467 2158
rect 1503 2162 1507 2163
rect 1503 2157 1507 2158
rect 1575 2162 1579 2163
rect 1575 2157 1579 2158
rect 1671 2162 1675 2163
rect 1671 2157 1675 2158
rect 1767 2162 1771 2163
rect 1767 2157 1771 2158
rect 112 2138 114 2157
rect 136 2141 138 2157
rect 248 2141 250 2157
rect 392 2141 394 2157
rect 544 2141 546 2157
rect 696 2141 698 2157
rect 840 2141 842 2157
rect 976 2141 978 2157
rect 1104 2141 1106 2157
rect 1232 2141 1234 2157
rect 1352 2141 1354 2157
rect 1464 2141 1466 2157
rect 1576 2141 1578 2157
rect 1672 2141 1674 2157
rect 134 2140 140 2141
rect 110 2137 116 2138
rect 110 2133 111 2137
rect 115 2133 116 2137
rect 134 2136 135 2140
rect 139 2136 140 2140
rect 134 2135 140 2136
rect 246 2140 252 2141
rect 246 2136 247 2140
rect 251 2136 252 2140
rect 246 2135 252 2136
rect 390 2140 396 2141
rect 390 2136 391 2140
rect 395 2136 396 2140
rect 390 2135 396 2136
rect 542 2140 548 2141
rect 542 2136 543 2140
rect 547 2136 548 2140
rect 542 2135 548 2136
rect 694 2140 700 2141
rect 694 2136 695 2140
rect 699 2136 700 2140
rect 694 2135 700 2136
rect 838 2140 844 2141
rect 838 2136 839 2140
rect 843 2136 844 2140
rect 838 2135 844 2136
rect 974 2140 980 2141
rect 974 2136 975 2140
rect 979 2136 980 2140
rect 974 2135 980 2136
rect 1102 2140 1108 2141
rect 1102 2136 1103 2140
rect 1107 2136 1108 2140
rect 1102 2135 1108 2136
rect 1230 2140 1236 2141
rect 1230 2136 1231 2140
rect 1235 2136 1236 2140
rect 1230 2135 1236 2136
rect 1350 2140 1356 2141
rect 1350 2136 1351 2140
rect 1355 2136 1356 2140
rect 1350 2135 1356 2136
rect 1462 2140 1468 2141
rect 1462 2136 1463 2140
rect 1467 2136 1468 2140
rect 1462 2135 1468 2136
rect 1574 2140 1580 2141
rect 1574 2136 1575 2140
rect 1579 2136 1580 2140
rect 1574 2135 1580 2136
rect 1670 2140 1676 2141
rect 1670 2136 1671 2140
rect 1675 2136 1676 2140
rect 1768 2138 1770 2157
rect 1808 2150 1810 2169
rect 2928 2153 2930 2169
rect 3016 2153 3018 2169
rect 3104 2153 3106 2169
rect 3192 2153 3194 2169
rect 3280 2153 3282 2169
rect 3368 2153 3370 2169
rect 2926 2152 2932 2153
rect 1806 2149 1812 2150
rect 1806 2145 1807 2149
rect 1811 2145 1812 2149
rect 2926 2148 2927 2152
rect 2931 2148 2932 2152
rect 2926 2147 2932 2148
rect 3014 2152 3020 2153
rect 3014 2148 3015 2152
rect 3019 2148 3020 2152
rect 3014 2147 3020 2148
rect 3102 2152 3108 2153
rect 3102 2148 3103 2152
rect 3107 2148 3108 2152
rect 3102 2147 3108 2148
rect 3190 2152 3196 2153
rect 3190 2148 3191 2152
rect 3195 2148 3196 2152
rect 3190 2147 3196 2148
rect 3278 2152 3284 2153
rect 3278 2148 3279 2152
rect 3283 2148 3284 2152
rect 3278 2147 3284 2148
rect 3366 2152 3372 2153
rect 3366 2148 3367 2152
rect 3371 2148 3372 2152
rect 3464 2150 3466 2169
rect 3366 2147 3372 2148
rect 3462 2149 3468 2150
rect 1806 2144 1812 2145
rect 3462 2145 3463 2149
rect 3467 2145 3468 2149
rect 3462 2144 3468 2145
rect 1670 2135 1676 2136
rect 1766 2137 1772 2138
rect 110 2132 116 2133
rect 1766 2133 1767 2137
rect 1771 2133 1772 2137
rect 2926 2133 2932 2134
rect 1766 2132 1772 2133
rect 1806 2132 1812 2133
rect 1806 2128 1807 2132
rect 1811 2128 1812 2132
rect 2926 2129 2927 2133
rect 2931 2129 2932 2133
rect 2926 2128 2932 2129
rect 3014 2133 3020 2134
rect 3014 2129 3015 2133
rect 3019 2129 3020 2133
rect 3014 2128 3020 2129
rect 3102 2133 3108 2134
rect 3102 2129 3103 2133
rect 3107 2129 3108 2133
rect 3102 2128 3108 2129
rect 3190 2133 3196 2134
rect 3190 2129 3191 2133
rect 3195 2129 3196 2133
rect 3190 2128 3196 2129
rect 3278 2133 3284 2134
rect 3278 2129 3279 2133
rect 3283 2129 3284 2133
rect 3278 2128 3284 2129
rect 3366 2133 3372 2134
rect 3366 2129 3367 2133
rect 3371 2129 3372 2133
rect 3366 2128 3372 2129
rect 3462 2132 3468 2133
rect 3462 2128 3463 2132
rect 3467 2128 3468 2132
rect 1806 2127 1812 2128
rect 134 2121 140 2122
rect 110 2120 116 2121
rect 110 2116 111 2120
rect 115 2116 116 2120
rect 134 2117 135 2121
rect 139 2117 140 2121
rect 134 2116 140 2117
rect 246 2121 252 2122
rect 246 2117 247 2121
rect 251 2117 252 2121
rect 246 2116 252 2117
rect 390 2121 396 2122
rect 390 2117 391 2121
rect 395 2117 396 2121
rect 390 2116 396 2117
rect 542 2121 548 2122
rect 542 2117 543 2121
rect 547 2117 548 2121
rect 542 2116 548 2117
rect 694 2121 700 2122
rect 694 2117 695 2121
rect 699 2117 700 2121
rect 694 2116 700 2117
rect 838 2121 844 2122
rect 838 2117 839 2121
rect 843 2117 844 2121
rect 838 2116 844 2117
rect 974 2121 980 2122
rect 974 2117 975 2121
rect 979 2117 980 2121
rect 974 2116 980 2117
rect 1102 2121 1108 2122
rect 1102 2117 1103 2121
rect 1107 2117 1108 2121
rect 1102 2116 1108 2117
rect 1230 2121 1236 2122
rect 1230 2117 1231 2121
rect 1235 2117 1236 2121
rect 1230 2116 1236 2117
rect 1350 2121 1356 2122
rect 1350 2117 1351 2121
rect 1355 2117 1356 2121
rect 1350 2116 1356 2117
rect 1462 2121 1468 2122
rect 1462 2117 1463 2121
rect 1467 2117 1468 2121
rect 1462 2116 1468 2117
rect 1574 2121 1580 2122
rect 1574 2117 1575 2121
rect 1579 2117 1580 2121
rect 1574 2116 1580 2117
rect 1670 2121 1676 2122
rect 1670 2117 1671 2121
rect 1675 2117 1676 2121
rect 1670 2116 1676 2117
rect 1766 2120 1772 2121
rect 1766 2116 1767 2120
rect 1771 2116 1772 2120
rect 110 2115 116 2116
rect 112 2095 114 2115
rect 136 2095 138 2116
rect 248 2095 250 2116
rect 392 2095 394 2116
rect 544 2095 546 2116
rect 696 2095 698 2116
rect 840 2095 842 2116
rect 976 2095 978 2116
rect 1104 2095 1106 2116
rect 1232 2095 1234 2116
rect 1352 2095 1354 2116
rect 1464 2095 1466 2116
rect 1576 2095 1578 2116
rect 1672 2095 1674 2116
rect 1766 2115 1772 2116
rect 1768 2095 1770 2115
rect 1808 2103 1810 2127
rect 2928 2103 2930 2128
rect 3016 2103 3018 2128
rect 3104 2103 3106 2128
rect 3192 2103 3194 2128
rect 3280 2103 3282 2128
rect 3368 2103 3370 2128
rect 3462 2127 3468 2128
rect 3464 2103 3466 2127
rect 1807 2102 1811 2103
rect 1807 2097 1811 2098
rect 1831 2102 1835 2103
rect 1831 2097 1835 2098
rect 1991 2102 1995 2103
rect 1991 2097 1995 2098
rect 2167 2102 2171 2103
rect 2167 2097 2171 2098
rect 2343 2102 2347 2103
rect 2343 2097 2347 2098
rect 2503 2102 2507 2103
rect 2503 2097 2507 2098
rect 2655 2102 2659 2103
rect 2655 2097 2659 2098
rect 2791 2102 2795 2103
rect 2791 2097 2795 2098
rect 2919 2102 2923 2103
rect 2919 2097 2923 2098
rect 2927 2102 2931 2103
rect 2927 2097 2931 2098
rect 3015 2102 3019 2103
rect 3015 2097 3019 2098
rect 3039 2102 3043 2103
rect 3039 2097 3043 2098
rect 3103 2102 3107 2103
rect 3103 2097 3107 2098
rect 3159 2102 3163 2103
rect 3159 2097 3163 2098
rect 3191 2102 3195 2103
rect 3191 2097 3195 2098
rect 3271 2102 3275 2103
rect 3271 2097 3275 2098
rect 3279 2102 3283 2103
rect 3279 2097 3283 2098
rect 3367 2102 3371 2103
rect 3367 2097 3371 2098
rect 3463 2102 3467 2103
rect 3463 2097 3467 2098
rect 111 2094 115 2095
rect 111 2089 115 2090
rect 135 2094 139 2095
rect 135 2089 139 2090
rect 223 2094 227 2095
rect 223 2089 227 2090
rect 247 2094 251 2095
rect 247 2089 251 2090
rect 343 2094 347 2095
rect 343 2089 347 2090
rect 391 2094 395 2095
rect 391 2089 395 2090
rect 463 2094 467 2095
rect 463 2089 467 2090
rect 543 2094 547 2095
rect 543 2089 547 2090
rect 583 2094 587 2095
rect 583 2089 587 2090
rect 695 2094 699 2095
rect 695 2089 699 2090
rect 703 2094 707 2095
rect 703 2089 707 2090
rect 823 2094 827 2095
rect 823 2089 827 2090
rect 839 2094 843 2095
rect 839 2089 843 2090
rect 935 2094 939 2095
rect 935 2089 939 2090
rect 975 2094 979 2095
rect 975 2089 979 2090
rect 1047 2094 1051 2095
rect 1047 2089 1051 2090
rect 1103 2094 1107 2095
rect 1103 2089 1107 2090
rect 1159 2094 1163 2095
rect 1159 2089 1163 2090
rect 1231 2094 1235 2095
rect 1231 2089 1235 2090
rect 1279 2094 1283 2095
rect 1279 2089 1283 2090
rect 1351 2094 1355 2095
rect 1351 2089 1355 2090
rect 1463 2094 1467 2095
rect 1463 2089 1467 2090
rect 1575 2094 1579 2095
rect 1575 2089 1579 2090
rect 1671 2094 1675 2095
rect 1671 2089 1675 2090
rect 1767 2094 1771 2095
rect 1767 2089 1771 2090
rect 112 2073 114 2089
rect 110 2072 116 2073
rect 136 2072 138 2089
rect 224 2072 226 2089
rect 344 2072 346 2089
rect 464 2072 466 2089
rect 584 2072 586 2089
rect 704 2072 706 2089
rect 824 2072 826 2089
rect 936 2072 938 2089
rect 1048 2072 1050 2089
rect 1160 2072 1162 2089
rect 1280 2072 1282 2089
rect 1768 2073 1770 2089
rect 1808 2081 1810 2097
rect 1806 2080 1812 2081
rect 1832 2080 1834 2097
rect 1992 2080 1994 2097
rect 2168 2080 2170 2097
rect 2344 2080 2346 2097
rect 2504 2080 2506 2097
rect 2656 2080 2658 2097
rect 2792 2080 2794 2097
rect 2920 2080 2922 2097
rect 3040 2080 3042 2097
rect 3160 2080 3162 2097
rect 3272 2080 3274 2097
rect 3368 2080 3370 2097
rect 3464 2081 3466 2097
rect 3462 2080 3468 2081
rect 1806 2076 1807 2080
rect 1811 2076 1812 2080
rect 1806 2075 1812 2076
rect 1830 2079 1836 2080
rect 1830 2075 1831 2079
rect 1835 2075 1836 2079
rect 1830 2074 1836 2075
rect 1990 2079 1996 2080
rect 1990 2075 1991 2079
rect 1995 2075 1996 2079
rect 1990 2074 1996 2075
rect 2166 2079 2172 2080
rect 2166 2075 2167 2079
rect 2171 2075 2172 2079
rect 2166 2074 2172 2075
rect 2342 2079 2348 2080
rect 2342 2075 2343 2079
rect 2347 2075 2348 2079
rect 2342 2074 2348 2075
rect 2502 2079 2508 2080
rect 2502 2075 2503 2079
rect 2507 2075 2508 2079
rect 2502 2074 2508 2075
rect 2654 2079 2660 2080
rect 2654 2075 2655 2079
rect 2659 2075 2660 2079
rect 2654 2074 2660 2075
rect 2790 2079 2796 2080
rect 2790 2075 2791 2079
rect 2795 2075 2796 2079
rect 2790 2074 2796 2075
rect 2918 2079 2924 2080
rect 2918 2075 2919 2079
rect 2923 2075 2924 2079
rect 2918 2074 2924 2075
rect 3038 2079 3044 2080
rect 3038 2075 3039 2079
rect 3043 2075 3044 2079
rect 3038 2074 3044 2075
rect 3158 2079 3164 2080
rect 3158 2075 3159 2079
rect 3163 2075 3164 2079
rect 3158 2074 3164 2075
rect 3270 2079 3276 2080
rect 3270 2075 3271 2079
rect 3275 2075 3276 2079
rect 3270 2074 3276 2075
rect 3366 2079 3372 2080
rect 3366 2075 3367 2079
rect 3371 2075 3372 2079
rect 3462 2076 3463 2080
rect 3467 2076 3468 2080
rect 3462 2075 3468 2076
rect 3366 2074 3372 2075
rect 1766 2072 1772 2073
rect 110 2068 111 2072
rect 115 2068 116 2072
rect 110 2067 116 2068
rect 134 2071 140 2072
rect 134 2067 135 2071
rect 139 2067 140 2071
rect 134 2066 140 2067
rect 222 2071 228 2072
rect 222 2067 223 2071
rect 227 2067 228 2071
rect 222 2066 228 2067
rect 342 2071 348 2072
rect 342 2067 343 2071
rect 347 2067 348 2071
rect 342 2066 348 2067
rect 462 2071 468 2072
rect 462 2067 463 2071
rect 467 2067 468 2071
rect 462 2066 468 2067
rect 582 2071 588 2072
rect 582 2067 583 2071
rect 587 2067 588 2071
rect 582 2066 588 2067
rect 702 2071 708 2072
rect 702 2067 703 2071
rect 707 2067 708 2071
rect 702 2066 708 2067
rect 822 2071 828 2072
rect 822 2067 823 2071
rect 827 2067 828 2071
rect 822 2066 828 2067
rect 934 2071 940 2072
rect 934 2067 935 2071
rect 939 2067 940 2071
rect 934 2066 940 2067
rect 1046 2071 1052 2072
rect 1046 2067 1047 2071
rect 1051 2067 1052 2071
rect 1046 2066 1052 2067
rect 1158 2071 1164 2072
rect 1158 2067 1159 2071
rect 1163 2067 1164 2071
rect 1158 2066 1164 2067
rect 1278 2071 1284 2072
rect 1278 2067 1279 2071
rect 1283 2067 1284 2071
rect 1766 2068 1767 2072
rect 1771 2068 1772 2072
rect 1766 2067 1772 2068
rect 1278 2066 1284 2067
rect 1806 2063 1812 2064
rect 1806 2059 1807 2063
rect 1811 2059 1812 2063
rect 3462 2063 3468 2064
rect 1806 2058 1812 2059
rect 1830 2060 1836 2061
rect 110 2055 116 2056
rect 110 2051 111 2055
rect 115 2051 116 2055
rect 1766 2055 1772 2056
rect 110 2050 116 2051
rect 134 2052 140 2053
rect 112 2023 114 2050
rect 134 2048 135 2052
rect 139 2048 140 2052
rect 134 2047 140 2048
rect 222 2052 228 2053
rect 222 2048 223 2052
rect 227 2048 228 2052
rect 222 2047 228 2048
rect 342 2052 348 2053
rect 342 2048 343 2052
rect 347 2048 348 2052
rect 342 2047 348 2048
rect 462 2052 468 2053
rect 462 2048 463 2052
rect 467 2048 468 2052
rect 462 2047 468 2048
rect 582 2052 588 2053
rect 582 2048 583 2052
rect 587 2048 588 2052
rect 582 2047 588 2048
rect 702 2052 708 2053
rect 702 2048 703 2052
rect 707 2048 708 2052
rect 702 2047 708 2048
rect 822 2052 828 2053
rect 822 2048 823 2052
rect 827 2048 828 2052
rect 822 2047 828 2048
rect 934 2052 940 2053
rect 934 2048 935 2052
rect 939 2048 940 2052
rect 934 2047 940 2048
rect 1046 2052 1052 2053
rect 1046 2048 1047 2052
rect 1051 2048 1052 2052
rect 1046 2047 1052 2048
rect 1158 2052 1164 2053
rect 1158 2048 1159 2052
rect 1163 2048 1164 2052
rect 1158 2047 1164 2048
rect 1278 2052 1284 2053
rect 1278 2048 1279 2052
rect 1283 2048 1284 2052
rect 1766 2051 1767 2055
rect 1771 2051 1772 2055
rect 1766 2050 1772 2051
rect 1278 2047 1284 2048
rect 136 2023 138 2047
rect 224 2023 226 2047
rect 344 2023 346 2047
rect 464 2023 466 2047
rect 584 2023 586 2047
rect 704 2023 706 2047
rect 824 2023 826 2047
rect 936 2023 938 2047
rect 1048 2023 1050 2047
rect 1160 2023 1162 2047
rect 1280 2023 1282 2047
rect 1768 2023 1770 2050
rect 1808 2035 1810 2058
rect 1830 2056 1831 2060
rect 1835 2056 1836 2060
rect 1830 2055 1836 2056
rect 1990 2060 1996 2061
rect 1990 2056 1991 2060
rect 1995 2056 1996 2060
rect 1990 2055 1996 2056
rect 2166 2060 2172 2061
rect 2166 2056 2167 2060
rect 2171 2056 2172 2060
rect 2166 2055 2172 2056
rect 2342 2060 2348 2061
rect 2342 2056 2343 2060
rect 2347 2056 2348 2060
rect 2342 2055 2348 2056
rect 2502 2060 2508 2061
rect 2502 2056 2503 2060
rect 2507 2056 2508 2060
rect 2502 2055 2508 2056
rect 2654 2060 2660 2061
rect 2654 2056 2655 2060
rect 2659 2056 2660 2060
rect 2654 2055 2660 2056
rect 2790 2060 2796 2061
rect 2790 2056 2791 2060
rect 2795 2056 2796 2060
rect 2790 2055 2796 2056
rect 2918 2060 2924 2061
rect 2918 2056 2919 2060
rect 2923 2056 2924 2060
rect 2918 2055 2924 2056
rect 3038 2060 3044 2061
rect 3038 2056 3039 2060
rect 3043 2056 3044 2060
rect 3038 2055 3044 2056
rect 3158 2060 3164 2061
rect 3158 2056 3159 2060
rect 3163 2056 3164 2060
rect 3158 2055 3164 2056
rect 3270 2060 3276 2061
rect 3270 2056 3271 2060
rect 3275 2056 3276 2060
rect 3270 2055 3276 2056
rect 3366 2060 3372 2061
rect 3366 2056 3367 2060
rect 3371 2056 3372 2060
rect 3462 2059 3463 2063
rect 3467 2059 3468 2063
rect 3462 2058 3468 2059
rect 3366 2055 3372 2056
rect 1832 2035 1834 2055
rect 1992 2035 1994 2055
rect 2168 2035 2170 2055
rect 2344 2035 2346 2055
rect 2504 2035 2506 2055
rect 2656 2035 2658 2055
rect 2792 2035 2794 2055
rect 2920 2035 2922 2055
rect 3040 2035 3042 2055
rect 3160 2035 3162 2055
rect 3272 2035 3274 2055
rect 3368 2035 3370 2055
rect 3464 2035 3466 2058
rect 1807 2034 1811 2035
rect 1807 2029 1811 2030
rect 1831 2034 1835 2035
rect 1831 2029 1835 2030
rect 1991 2034 1995 2035
rect 1991 2029 1995 2030
rect 2015 2034 2019 2035
rect 2015 2029 2019 2030
rect 2167 2034 2171 2035
rect 2167 2029 2171 2030
rect 2223 2034 2227 2035
rect 2223 2029 2227 2030
rect 2343 2034 2347 2035
rect 2343 2029 2347 2030
rect 2431 2034 2435 2035
rect 2431 2029 2435 2030
rect 2503 2034 2507 2035
rect 2503 2029 2507 2030
rect 2631 2034 2635 2035
rect 2631 2029 2635 2030
rect 2655 2034 2659 2035
rect 2655 2029 2659 2030
rect 2791 2034 2795 2035
rect 2791 2029 2795 2030
rect 2823 2034 2827 2035
rect 2823 2029 2827 2030
rect 2919 2034 2923 2035
rect 2919 2029 2923 2030
rect 3007 2034 3011 2035
rect 3007 2029 3011 2030
rect 3039 2034 3043 2035
rect 3039 2029 3043 2030
rect 3159 2034 3163 2035
rect 3159 2029 3163 2030
rect 3199 2034 3203 2035
rect 3199 2029 3203 2030
rect 3271 2034 3275 2035
rect 3271 2029 3275 2030
rect 3367 2034 3371 2035
rect 3367 2029 3371 2030
rect 3463 2034 3467 2035
rect 3463 2029 3467 2030
rect 111 2022 115 2023
rect 111 2017 115 2018
rect 135 2022 139 2023
rect 135 2017 139 2018
rect 223 2022 227 2023
rect 223 2017 227 2018
rect 239 2022 243 2023
rect 239 2017 243 2018
rect 343 2022 347 2023
rect 343 2017 347 2018
rect 367 2022 371 2023
rect 367 2017 371 2018
rect 463 2022 467 2023
rect 463 2017 467 2018
rect 503 2022 507 2023
rect 503 2017 507 2018
rect 583 2022 587 2023
rect 583 2017 587 2018
rect 639 2022 643 2023
rect 639 2017 643 2018
rect 703 2022 707 2023
rect 703 2017 707 2018
rect 775 2022 779 2023
rect 775 2017 779 2018
rect 823 2022 827 2023
rect 823 2017 827 2018
rect 911 2022 915 2023
rect 911 2017 915 2018
rect 935 2022 939 2023
rect 935 2017 939 2018
rect 1047 2022 1051 2023
rect 1047 2017 1051 2018
rect 1159 2022 1163 2023
rect 1159 2017 1163 2018
rect 1183 2022 1187 2023
rect 1183 2017 1187 2018
rect 1279 2022 1283 2023
rect 1279 2017 1283 2018
rect 1327 2022 1331 2023
rect 1327 2017 1331 2018
rect 1767 2022 1771 2023
rect 1767 2017 1771 2018
rect 112 1998 114 2017
rect 136 2001 138 2017
rect 240 2001 242 2017
rect 368 2001 370 2017
rect 504 2001 506 2017
rect 640 2001 642 2017
rect 776 2001 778 2017
rect 912 2001 914 2017
rect 1048 2001 1050 2017
rect 1184 2001 1186 2017
rect 1328 2001 1330 2017
rect 134 2000 140 2001
rect 110 1997 116 1998
rect 110 1993 111 1997
rect 115 1993 116 1997
rect 134 1996 135 2000
rect 139 1996 140 2000
rect 134 1995 140 1996
rect 238 2000 244 2001
rect 238 1996 239 2000
rect 243 1996 244 2000
rect 238 1995 244 1996
rect 366 2000 372 2001
rect 366 1996 367 2000
rect 371 1996 372 2000
rect 366 1995 372 1996
rect 502 2000 508 2001
rect 502 1996 503 2000
rect 507 1996 508 2000
rect 502 1995 508 1996
rect 638 2000 644 2001
rect 638 1996 639 2000
rect 643 1996 644 2000
rect 638 1995 644 1996
rect 774 2000 780 2001
rect 774 1996 775 2000
rect 779 1996 780 2000
rect 774 1995 780 1996
rect 910 2000 916 2001
rect 910 1996 911 2000
rect 915 1996 916 2000
rect 910 1995 916 1996
rect 1046 2000 1052 2001
rect 1046 1996 1047 2000
rect 1051 1996 1052 2000
rect 1046 1995 1052 1996
rect 1182 2000 1188 2001
rect 1182 1996 1183 2000
rect 1187 1996 1188 2000
rect 1182 1995 1188 1996
rect 1326 2000 1332 2001
rect 1326 1996 1327 2000
rect 1331 1996 1332 2000
rect 1768 1998 1770 2017
rect 1808 2010 1810 2029
rect 1832 2013 1834 2029
rect 2016 2013 2018 2029
rect 2224 2013 2226 2029
rect 2432 2013 2434 2029
rect 2632 2013 2634 2029
rect 2824 2013 2826 2029
rect 3008 2013 3010 2029
rect 3200 2013 3202 2029
rect 3368 2013 3370 2029
rect 1830 2012 1836 2013
rect 1806 2009 1812 2010
rect 1806 2005 1807 2009
rect 1811 2005 1812 2009
rect 1830 2008 1831 2012
rect 1835 2008 1836 2012
rect 1830 2007 1836 2008
rect 2014 2012 2020 2013
rect 2014 2008 2015 2012
rect 2019 2008 2020 2012
rect 2014 2007 2020 2008
rect 2222 2012 2228 2013
rect 2222 2008 2223 2012
rect 2227 2008 2228 2012
rect 2222 2007 2228 2008
rect 2430 2012 2436 2013
rect 2430 2008 2431 2012
rect 2435 2008 2436 2012
rect 2430 2007 2436 2008
rect 2630 2012 2636 2013
rect 2630 2008 2631 2012
rect 2635 2008 2636 2012
rect 2630 2007 2636 2008
rect 2822 2012 2828 2013
rect 2822 2008 2823 2012
rect 2827 2008 2828 2012
rect 2822 2007 2828 2008
rect 3006 2012 3012 2013
rect 3006 2008 3007 2012
rect 3011 2008 3012 2012
rect 3006 2007 3012 2008
rect 3198 2012 3204 2013
rect 3198 2008 3199 2012
rect 3203 2008 3204 2012
rect 3198 2007 3204 2008
rect 3366 2012 3372 2013
rect 3366 2008 3367 2012
rect 3371 2008 3372 2012
rect 3464 2010 3466 2029
rect 3366 2007 3372 2008
rect 3462 2009 3468 2010
rect 1806 2004 1812 2005
rect 3462 2005 3463 2009
rect 3467 2005 3468 2009
rect 3462 2004 3468 2005
rect 1326 1995 1332 1996
rect 1766 1997 1772 1998
rect 110 1992 116 1993
rect 1766 1993 1767 1997
rect 1771 1993 1772 1997
rect 1830 1993 1836 1994
rect 1766 1992 1772 1993
rect 1806 1992 1812 1993
rect 1806 1988 1807 1992
rect 1811 1988 1812 1992
rect 1830 1989 1831 1993
rect 1835 1989 1836 1993
rect 1830 1988 1836 1989
rect 2014 1993 2020 1994
rect 2014 1989 2015 1993
rect 2019 1989 2020 1993
rect 2014 1988 2020 1989
rect 2222 1993 2228 1994
rect 2222 1989 2223 1993
rect 2227 1989 2228 1993
rect 2222 1988 2228 1989
rect 2430 1993 2436 1994
rect 2430 1989 2431 1993
rect 2435 1989 2436 1993
rect 2430 1988 2436 1989
rect 2630 1993 2636 1994
rect 2630 1989 2631 1993
rect 2635 1989 2636 1993
rect 2630 1988 2636 1989
rect 2822 1993 2828 1994
rect 2822 1989 2823 1993
rect 2827 1989 2828 1993
rect 2822 1988 2828 1989
rect 3006 1993 3012 1994
rect 3006 1989 3007 1993
rect 3011 1989 3012 1993
rect 3006 1988 3012 1989
rect 3198 1993 3204 1994
rect 3198 1989 3199 1993
rect 3203 1989 3204 1993
rect 3198 1988 3204 1989
rect 3366 1993 3372 1994
rect 3366 1989 3367 1993
rect 3371 1989 3372 1993
rect 3366 1988 3372 1989
rect 3462 1992 3468 1993
rect 3462 1988 3463 1992
rect 3467 1988 3468 1992
rect 1806 1987 1812 1988
rect 134 1981 140 1982
rect 110 1980 116 1981
rect 110 1976 111 1980
rect 115 1976 116 1980
rect 134 1977 135 1981
rect 139 1977 140 1981
rect 134 1976 140 1977
rect 238 1981 244 1982
rect 238 1977 239 1981
rect 243 1977 244 1981
rect 238 1976 244 1977
rect 366 1981 372 1982
rect 366 1977 367 1981
rect 371 1977 372 1981
rect 366 1976 372 1977
rect 502 1981 508 1982
rect 502 1977 503 1981
rect 507 1977 508 1981
rect 502 1976 508 1977
rect 638 1981 644 1982
rect 638 1977 639 1981
rect 643 1977 644 1981
rect 638 1976 644 1977
rect 774 1981 780 1982
rect 774 1977 775 1981
rect 779 1977 780 1981
rect 774 1976 780 1977
rect 910 1981 916 1982
rect 910 1977 911 1981
rect 915 1977 916 1981
rect 910 1976 916 1977
rect 1046 1981 1052 1982
rect 1046 1977 1047 1981
rect 1051 1977 1052 1981
rect 1046 1976 1052 1977
rect 1182 1981 1188 1982
rect 1182 1977 1183 1981
rect 1187 1977 1188 1981
rect 1182 1976 1188 1977
rect 1326 1981 1332 1982
rect 1326 1977 1327 1981
rect 1331 1977 1332 1981
rect 1326 1976 1332 1977
rect 1766 1980 1772 1981
rect 1766 1976 1767 1980
rect 1771 1976 1772 1980
rect 110 1975 116 1976
rect 112 1955 114 1975
rect 136 1955 138 1976
rect 240 1955 242 1976
rect 368 1955 370 1976
rect 504 1955 506 1976
rect 640 1955 642 1976
rect 776 1955 778 1976
rect 912 1955 914 1976
rect 1048 1955 1050 1976
rect 1184 1955 1186 1976
rect 1328 1955 1330 1976
rect 1766 1975 1772 1976
rect 1768 1955 1770 1975
rect 1808 1967 1810 1987
rect 1832 1967 1834 1988
rect 2016 1967 2018 1988
rect 2224 1967 2226 1988
rect 2432 1967 2434 1988
rect 2632 1967 2634 1988
rect 2824 1967 2826 1988
rect 3008 1967 3010 1988
rect 3200 1967 3202 1988
rect 3368 1967 3370 1988
rect 3462 1987 3468 1988
rect 3464 1967 3466 1987
rect 1807 1966 1811 1967
rect 1807 1961 1811 1962
rect 1831 1966 1835 1967
rect 1831 1961 1835 1962
rect 1863 1966 1867 1967
rect 1863 1961 1867 1962
rect 1999 1966 2003 1967
rect 1999 1961 2003 1962
rect 2015 1966 2019 1967
rect 2015 1961 2019 1962
rect 2143 1966 2147 1967
rect 2143 1961 2147 1962
rect 2223 1966 2227 1967
rect 2223 1961 2227 1962
rect 2287 1966 2291 1967
rect 2287 1961 2291 1962
rect 2431 1966 2435 1967
rect 2431 1961 2435 1962
rect 2575 1966 2579 1967
rect 2575 1961 2579 1962
rect 2631 1966 2635 1967
rect 2631 1961 2635 1962
rect 2711 1966 2715 1967
rect 2711 1961 2715 1962
rect 2823 1966 2827 1967
rect 2823 1961 2827 1962
rect 2831 1966 2835 1967
rect 2831 1961 2835 1962
rect 2951 1966 2955 1967
rect 2951 1961 2955 1962
rect 3007 1966 3011 1967
rect 3007 1961 3011 1962
rect 3063 1966 3067 1967
rect 3063 1961 3067 1962
rect 3167 1966 3171 1967
rect 3167 1961 3171 1962
rect 3199 1966 3203 1967
rect 3199 1961 3203 1962
rect 3279 1966 3283 1967
rect 3279 1961 3283 1962
rect 3367 1966 3371 1967
rect 3367 1961 3371 1962
rect 3463 1966 3467 1967
rect 3463 1961 3467 1962
rect 111 1954 115 1955
rect 111 1949 115 1950
rect 135 1954 139 1955
rect 135 1949 139 1950
rect 239 1954 243 1955
rect 239 1949 243 1950
rect 295 1954 299 1955
rect 295 1949 299 1950
rect 367 1954 371 1955
rect 367 1949 371 1950
rect 423 1954 427 1955
rect 423 1949 427 1950
rect 503 1954 507 1955
rect 503 1949 507 1950
rect 559 1954 563 1955
rect 559 1949 563 1950
rect 639 1954 643 1955
rect 639 1949 643 1950
rect 703 1954 707 1955
rect 703 1949 707 1950
rect 775 1954 779 1955
rect 775 1949 779 1950
rect 855 1954 859 1955
rect 855 1949 859 1950
rect 911 1954 915 1955
rect 911 1949 915 1950
rect 1007 1954 1011 1955
rect 1007 1949 1011 1950
rect 1047 1954 1051 1955
rect 1047 1949 1051 1950
rect 1159 1954 1163 1955
rect 1159 1949 1163 1950
rect 1183 1954 1187 1955
rect 1183 1949 1187 1950
rect 1311 1954 1315 1955
rect 1311 1949 1315 1950
rect 1327 1954 1331 1955
rect 1327 1949 1331 1950
rect 1471 1954 1475 1955
rect 1471 1949 1475 1950
rect 1767 1954 1771 1955
rect 1767 1949 1771 1950
rect 112 1933 114 1949
rect 110 1932 116 1933
rect 296 1932 298 1949
rect 424 1932 426 1949
rect 560 1932 562 1949
rect 704 1932 706 1949
rect 856 1932 858 1949
rect 1008 1932 1010 1949
rect 1160 1932 1162 1949
rect 1312 1932 1314 1949
rect 1472 1932 1474 1949
rect 1768 1933 1770 1949
rect 1808 1945 1810 1961
rect 1806 1944 1812 1945
rect 1864 1944 1866 1961
rect 2000 1944 2002 1961
rect 2144 1944 2146 1961
rect 2288 1944 2290 1961
rect 2432 1944 2434 1961
rect 2576 1944 2578 1961
rect 2712 1944 2714 1961
rect 2832 1944 2834 1961
rect 2952 1944 2954 1961
rect 3064 1944 3066 1961
rect 3168 1944 3170 1961
rect 3280 1944 3282 1961
rect 3368 1944 3370 1961
rect 3464 1945 3466 1961
rect 3462 1944 3468 1945
rect 1806 1940 1807 1944
rect 1811 1940 1812 1944
rect 1806 1939 1812 1940
rect 1862 1943 1868 1944
rect 1862 1939 1863 1943
rect 1867 1939 1868 1943
rect 1862 1938 1868 1939
rect 1998 1943 2004 1944
rect 1998 1939 1999 1943
rect 2003 1939 2004 1943
rect 1998 1938 2004 1939
rect 2142 1943 2148 1944
rect 2142 1939 2143 1943
rect 2147 1939 2148 1943
rect 2142 1938 2148 1939
rect 2286 1943 2292 1944
rect 2286 1939 2287 1943
rect 2291 1939 2292 1943
rect 2286 1938 2292 1939
rect 2430 1943 2436 1944
rect 2430 1939 2431 1943
rect 2435 1939 2436 1943
rect 2430 1938 2436 1939
rect 2574 1943 2580 1944
rect 2574 1939 2575 1943
rect 2579 1939 2580 1943
rect 2574 1938 2580 1939
rect 2710 1943 2716 1944
rect 2710 1939 2711 1943
rect 2715 1939 2716 1943
rect 2710 1938 2716 1939
rect 2830 1943 2836 1944
rect 2830 1939 2831 1943
rect 2835 1939 2836 1943
rect 2830 1938 2836 1939
rect 2950 1943 2956 1944
rect 2950 1939 2951 1943
rect 2955 1939 2956 1943
rect 2950 1938 2956 1939
rect 3062 1943 3068 1944
rect 3062 1939 3063 1943
rect 3067 1939 3068 1943
rect 3062 1938 3068 1939
rect 3166 1943 3172 1944
rect 3166 1939 3167 1943
rect 3171 1939 3172 1943
rect 3166 1938 3172 1939
rect 3278 1943 3284 1944
rect 3278 1939 3279 1943
rect 3283 1939 3284 1943
rect 3278 1938 3284 1939
rect 3366 1943 3372 1944
rect 3366 1939 3367 1943
rect 3371 1939 3372 1943
rect 3462 1940 3463 1944
rect 3467 1940 3468 1944
rect 3462 1939 3468 1940
rect 3366 1938 3372 1939
rect 1766 1932 1772 1933
rect 110 1928 111 1932
rect 115 1928 116 1932
rect 110 1927 116 1928
rect 294 1931 300 1932
rect 294 1927 295 1931
rect 299 1927 300 1931
rect 294 1926 300 1927
rect 422 1931 428 1932
rect 422 1927 423 1931
rect 427 1927 428 1931
rect 422 1926 428 1927
rect 558 1931 564 1932
rect 558 1927 559 1931
rect 563 1927 564 1931
rect 558 1926 564 1927
rect 702 1931 708 1932
rect 702 1927 703 1931
rect 707 1927 708 1931
rect 702 1926 708 1927
rect 854 1931 860 1932
rect 854 1927 855 1931
rect 859 1927 860 1931
rect 854 1926 860 1927
rect 1006 1931 1012 1932
rect 1006 1927 1007 1931
rect 1011 1927 1012 1931
rect 1006 1926 1012 1927
rect 1158 1931 1164 1932
rect 1158 1927 1159 1931
rect 1163 1927 1164 1931
rect 1158 1926 1164 1927
rect 1310 1931 1316 1932
rect 1310 1927 1311 1931
rect 1315 1927 1316 1931
rect 1310 1926 1316 1927
rect 1470 1931 1476 1932
rect 1470 1927 1471 1931
rect 1475 1927 1476 1931
rect 1766 1928 1767 1932
rect 1771 1928 1772 1932
rect 1766 1927 1772 1928
rect 1806 1927 1812 1928
rect 1470 1926 1476 1927
rect 1806 1923 1807 1927
rect 1811 1923 1812 1927
rect 3462 1927 3468 1928
rect 1806 1922 1812 1923
rect 1862 1924 1868 1925
rect 110 1915 116 1916
rect 110 1911 111 1915
rect 115 1911 116 1915
rect 1766 1915 1772 1916
rect 110 1910 116 1911
rect 294 1912 300 1913
rect 112 1891 114 1910
rect 294 1908 295 1912
rect 299 1908 300 1912
rect 294 1907 300 1908
rect 422 1912 428 1913
rect 422 1908 423 1912
rect 427 1908 428 1912
rect 422 1907 428 1908
rect 558 1912 564 1913
rect 558 1908 559 1912
rect 563 1908 564 1912
rect 558 1907 564 1908
rect 702 1912 708 1913
rect 702 1908 703 1912
rect 707 1908 708 1912
rect 702 1907 708 1908
rect 854 1912 860 1913
rect 854 1908 855 1912
rect 859 1908 860 1912
rect 854 1907 860 1908
rect 1006 1912 1012 1913
rect 1006 1908 1007 1912
rect 1011 1908 1012 1912
rect 1006 1907 1012 1908
rect 1158 1912 1164 1913
rect 1158 1908 1159 1912
rect 1163 1908 1164 1912
rect 1158 1907 1164 1908
rect 1310 1912 1316 1913
rect 1310 1908 1311 1912
rect 1315 1908 1316 1912
rect 1310 1907 1316 1908
rect 1470 1912 1476 1913
rect 1470 1908 1471 1912
rect 1475 1908 1476 1912
rect 1766 1911 1767 1915
rect 1771 1911 1772 1915
rect 1766 1910 1772 1911
rect 1470 1907 1476 1908
rect 296 1891 298 1907
rect 424 1891 426 1907
rect 560 1891 562 1907
rect 704 1891 706 1907
rect 856 1891 858 1907
rect 1008 1891 1010 1907
rect 1160 1891 1162 1907
rect 1312 1891 1314 1907
rect 1472 1891 1474 1907
rect 1768 1891 1770 1910
rect 1808 1899 1810 1922
rect 1862 1920 1863 1924
rect 1867 1920 1868 1924
rect 1862 1919 1868 1920
rect 1998 1924 2004 1925
rect 1998 1920 1999 1924
rect 2003 1920 2004 1924
rect 1998 1919 2004 1920
rect 2142 1924 2148 1925
rect 2142 1920 2143 1924
rect 2147 1920 2148 1924
rect 2142 1919 2148 1920
rect 2286 1924 2292 1925
rect 2286 1920 2287 1924
rect 2291 1920 2292 1924
rect 2286 1919 2292 1920
rect 2430 1924 2436 1925
rect 2430 1920 2431 1924
rect 2435 1920 2436 1924
rect 2430 1919 2436 1920
rect 2574 1924 2580 1925
rect 2574 1920 2575 1924
rect 2579 1920 2580 1924
rect 2574 1919 2580 1920
rect 2710 1924 2716 1925
rect 2710 1920 2711 1924
rect 2715 1920 2716 1924
rect 2710 1919 2716 1920
rect 2830 1924 2836 1925
rect 2830 1920 2831 1924
rect 2835 1920 2836 1924
rect 2830 1919 2836 1920
rect 2950 1924 2956 1925
rect 2950 1920 2951 1924
rect 2955 1920 2956 1924
rect 2950 1919 2956 1920
rect 3062 1924 3068 1925
rect 3062 1920 3063 1924
rect 3067 1920 3068 1924
rect 3062 1919 3068 1920
rect 3166 1924 3172 1925
rect 3166 1920 3167 1924
rect 3171 1920 3172 1924
rect 3166 1919 3172 1920
rect 3278 1924 3284 1925
rect 3278 1920 3279 1924
rect 3283 1920 3284 1924
rect 3278 1919 3284 1920
rect 3366 1924 3372 1925
rect 3366 1920 3367 1924
rect 3371 1920 3372 1924
rect 3462 1923 3463 1927
rect 3467 1923 3468 1927
rect 3462 1922 3468 1923
rect 3366 1919 3372 1920
rect 1864 1899 1866 1919
rect 2000 1899 2002 1919
rect 2144 1899 2146 1919
rect 2288 1899 2290 1919
rect 2432 1899 2434 1919
rect 2576 1899 2578 1919
rect 2712 1899 2714 1919
rect 2832 1899 2834 1919
rect 2952 1899 2954 1919
rect 3064 1899 3066 1919
rect 3168 1899 3170 1919
rect 3280 1899 3282 1919
rect 3368 1899 3370 1919
rect 3464 1899 3466 1922
rect 1807 1898 1811 1899
rect 1807 1893 1811 1894
rect 1863 1898 1867 1899
rect 1863 1893 1867 1894
rect 1999 1898 2003 1899
rect 1999 1893 2003 1894
rect 2015 1898 2019 1899
rect 2015 1893 2019 1894
rect 2111 1898 2115 1899
rect 2111 1893 2115 1894
rect 2143 1898 2147 1899
rect 2143 1893 2147 1894
rect 2215 1898 2219 1899
rect 2215 1893 2219 1894
rect 2287 1898 2291 1899
rect 2287 1893 2291 1894
rect 2327 1898 2331 1899
rect 2327 1893 2331 1894
rect 2431 1898 2435 1899
rect 2431 1893 2435 1894
rect 2439 1898 2443 1899
rect 2439 1893 2443 1894
rect 2543 1898 2547 1899
rect 2543 1893 2547 1894
rect 2575 1898 2579 1899
rect 2575 1893 2579 1894
rect 2647 1898 2651 1899
rect 2647 1893 2651 1894
rect 2711 1898 2715 1899
rect 2711 1893 2715 1894
rect 2759 1898 2763 1899
rect 2759 1893 2763 1894
rect 2831 1898 2835 1899
rect 2831 1893 2835 1894
rect 2871 1898 2875 1899
rect 2871 1893 2875 1894
rect 2951 1898 2955 1899
rect 2951 1893 2955 1894
rect 2983 1898 2987 1899
rect 2983 1893 2987 1894
rect 3063 1898 3067 1899
rect 3063 1893 3067 1894
rect 3167 1898 3171 1899
rect 3167 1893 3171 1894
rect 3279 1898 3283 1899
rect 3279 1893 3283 1894
rect 3367 1898 3371 1899
rect 3367 1893 3371 1894
rect 3463 1898 3467 1899
rect 3463 1893 3467 1894
rect 111 1890 115 1891
rect 111 1885 115 1886
rect 295 1890 299 1891
rect 295 1885 299 1886
rect 423 1890 427 1891
rect 423 1885 427 1886
rect 431 1890 435 1891
rect 431 1885 435 1886
rect 559 1890 563 1891
rect 559 1885 563 1886
rect 575 1890 579 1891
rect 575 1885 579 1886
rect 703 1890 707 1891
rect 703 1885 707 1886
rect 727 1890 731 1891
rect 727 1885 731 1886
rect 855 1890 859 1891
rect 855 1885 859 1886
rect 887 1890 891 1891
rect 887 1885 891 1886
rect 1007 1890 1011 1891
rect 1007 1885 1011 1886
rect 1047 1890 1051 1891
rect 1047 1885 1051 1886
rect 1159 1890 1163 1891
rect 1159 1885 1163 1886
rect 1199 1890 1203 1891
rect 1199 1885 1203 1886
rect 1311 1890 1315 1891
rect 1311 1885 1315 1886
rect 1351 1890 1355 1891
rect 1351 1885 1355 1886
rect 1471 1890 1475 1891
rect 1471 1885 1475 1886
rect 1511 1890 1515 1891
rect 1511 1885 1515 1886
rect 1671 1890 1675 1891
rect 1671 1885 1675 1886
rect 1767 1890 1771 1891
rect 1767 1885 1771 1886
rect 112 1866 114 1885
rect 432 1869 434 1885
rect 576 1869 578 1885
rect 728 1869 730 1885
rect 888 1869 890 1885
rect 1048 1869 1050 1885
rect 1200 1869 1202 1885
rect 1352 1869 1354 1885
rect 1512 1869 1514 1885
rect 1672 1869 1674 1885
rect 430 1868 436 1869
rect 110 1865 116 1866
rect 110 1861 111 1865
rect 115 1861 116 1865
rect 430 1864 431 1868
rect 435 1864 436 1868
rect 430 1863 436 1864
rect 574 1868 580 1869
rect 574 1864 575 1868
rect 579 1864 580 1868
rect 574 1863 580 1864
rect 726 1868 732 1869
rect 726 1864 727 1868
rect 731 1864 732 1868
rect 726 1863 732 1864
rect 886 1868 892 1869
rect 886 1864 887 1868
rect 891 1864 892 1868
rect 886 1863 892 1864
rect 1046 1868 1052 1869
rect 1046 1864 1047 1868
rect 1051 1864 1052 1868
rect 1046 1863 1052 1864
rect 1198 1868 1204 1869
rect 1198 1864 1199 1868
rect 1203 1864 1204 1868
rect 1198 1863 1204 1864
rect 1350 1868 1356 1869
rect 1350 1864 1351 1868
rect 1355 1864 1356 1868
rect 1350 1863 1356 1864
rect 1510 1868 1516 1869
rect 1510 1864 1511 1868
rect 1515 1864 1516 1868
rect 1510 1863 1516 1864
rect 1670 1868 1676 1869
rect 1670 1864 1671 1868
rect 1675 1864 1676 1868
rect 1768 1866 1770 1885
rect 1808 1874 1810 1893
rect 2016 1877 2018 1893
rect 2112 1877 2114 1893
rect 2216 1877 2218 1893
rect 2328 1877 2330 1893
rect 2440 1877 2442 1893
rect 2544 1877 2546 1893
rect 2648 1877 2650 1893
rect 2760 1877 2762 1893
rect 2872 1877 2874 1893
rect 2984 1877 2986 1893
rect 2014 1876 2020 1877
rect 1806 1873 1812 1874
rect 1806 1869 1807 1873
rect 1811 1869 1812 1873
rect 2014 1872 2015 1876
rect 2019 1872 2020 1876
rect 2014 1871 2020 1872
rect 2110 1876 2116 1877
rect 2110 1872 2111 1876
rect 2115 1872 2116 1876
rect 2110 1871 2116 1872
rect 2214 1876 2220 1877
rect 2214 1872 2215 1876
rect 2219 1872 2220 1876
rect 2214 1871 2220 1872
rect 2326 1876 2332 1877
rect 2326 1872 2327 1876
rect 2331 1872 2332 1876
rect 2326 1871 2332 1872
rect 2438 1876 2444 1877
rect 2438 1872 2439 1876
rect 2443 1872 2444 1876
rect 2438 1871 2444 1872
rect 2542 1876 2548 1877
rect 2542 1872 2543 1876
rect 2547 1872 2548 1876
rect 2542 1871 2548 1872
rect 2646 1876 2652 1877
rect 2646 1872 2647 1876
rect 2651 1872 2652 1876
rect 2646 1871 2652 1872
rect 2758 1876 2764 1877
rect 2758 1872 2759 1876
rect 2763 1872 2764 1876
rect 2758 1871 2764 1872
rect 2870 1876 2876 1877
rect 2870 1872 2871 1876
rect 2875 1872 2876 1876
rect 2870 1871 2876 1872
rect 2982 1876 2988 1877
rect 2982 1872 2983 1876
rect 2987 1872 2988 1876
rect 3464 1874 3466 1893
rect 2982 1871 2988 1872
rect 3462 1873 3468 1874
rect 1806 1868 1812 1869
rect 3462 1869 3463 1873
rect 3467 1869 3468 1873
rect 3462 1868 3468 1869
rect 1670 1863 1676 1864
rect 1766 1865 1772 1866
rect 110 1860 116 1861
rect 1766 1861 1767 1865
rect 1771 1861 1772 1865
rect 1766 1860 1772 1861
rect 2014 1857 2020 1858
rect 1806 1856 1812 1857
rect 1806 1852 1807 1856
rect 1811 1852 1812 1856
rect 2014 1853 2015 1857
rect 2019 1853 2020 1857
rect 2014 1852 2020 1853
rect 2110 1857 2116 1858
rect 2110 1853 2111 1857
rect 2115 1853 2116 1857
rect 2110 1852 2116 1853
rect 2214 1857 2220 1858
rect 2214 1853 2215 1857
rect 2219 1853 2220 1857
rect 2214 1852 2220 1853
rect 2326 1857 2332 1858
rect 2326 1853 2327 1857
rect 2331 1853 2332 1857
rect 2326 1852 2332 1853
rect 2438 1857 2444 1858
rect 2438 1853 2439 1857
rect 2443 1853 2444 1857
rect 2438 1852 2444 1853
rect 2542 1857 2548 1858
rect 2542 1853 2543 1857
rect 2547 1853 2548 1857
rect 2542 1852 2548 1853
rect 2646 1857 2652 1858
rect 2646 1853 2647 1857
rect 2651 1853 2652 1857
rect 2646 1852 2652 1853
rect 2758 1857 2764 1858
rect 2758 1853 2759 1857
rect 2763 1853 2764 1857
rect 2758 1852 2764 1853
rect 2870 1857 2876 1858
rect 2870 1853 2871 1857
rect 2875 1853 2876 1857
rect 2870 1852 2876 1853
rect 2982 1857 2988 1858
rect 2982 1853 2983 1857
rect 2987 1853 2988 1857
rect 2982 1852 2988 1853
rect 3462 1856 3468 1857
rect 3462 1852 3463 1856
rect 3467 1852 3468 1856
rect 1806 1851 1812 1852
rect 430 1849 436 1850
rect 110 1848 116 1849
rect 110 1844 111 1848
rect 115 1844 116 1848
rect 430 1845 431 1849
rect 435 1845 436 1849
rect 430 1844 436 1845
rect 574 1849 580 1850
rect 574 1845 575 1849
rect 579 1845 580 1849
rect 574 1844 580 1845
rect 726 1849 732 1850
rect 726 1845 727 1849
rect 731 1845 732 1849
rect 726 1844 732 1845
rect 886 1849 892 1850
rect 886 1845 887 1849
rect 891 1845 892 1849
rect 886 1844 892 1845
rect 1046 1849 1052 1850
rect 1046 1845 1047 1849
rect 1051 1845 1052 1849
rect 1046 1844 1052 1845
rect 1198 1849 1204 1850
rect 1198 1845 1199 1849
rect 1203 1845 1204 1849
rect 1198 1844 1204 1845
rect 1350 1849 1356 1850
rect 1350 1845 1351 1849
rect 1355 1845 1356 1849
rect 1350 1844 1356 1845
rect 1510 1849 1516 1850
rect 1510 1845 1511 1849
rect 1515 1845 1516 1849
rect 1510 1844 1516 1845
rect 1670 1849 1676 1850
rect 1670 1845 1671 1849
rect 1675 1845 1676 1849
rect 1670 1844 1676 1845
rect 1766 1848 1772 1849
rect 1766 1844 1767 1848
rect 1771 1844 1772 1848
rect 110 1843 116 1844
rect 112 1823 114 1843
rect 432 1823 434 1844
rect 576 1823 578 1844
rect 728 1823 730 1844
rect 888 1823 890 1844
rect 1048 1823 1050 1844
rect 1200 1823 1202 1844
rect 1352 1823 1354 1844
rect 1512 1823 1514 1844
rect 1672 1823 1674 1844
rect 1766 1843 1772 1844
rect 1768 1823 1770 1843
rect 1808 1827 1810 1851
rect 2016 1827 2018 1852
rect 2112 1827 2114 1852
rect 2216 1827 2218 1852
rect 2328 1827 2330 1852
rect 2440 1827 2442 1852
rect 2544 1827 2546 1852
rect 2648 1827 2650 1852
rect 2760 1827 2762 1852
rect 2872 1827 2874 1852
rect 2984 1827 2986 1852
rect 3462 1851 3468 1852
rect 3464 1827 3466 1851
rect 1807 1826 1811 1827
rect 111 1822 115 1823
rect 111 1817 115 1818
rect 431 1822 435 1823
rect 431 1817 435 1818
rect 511 1822 515 1823
rect 511 1817 515 1818
rect 575 1822 579 1823
rect 575 1817 579 1818
rect 631 1822 635 1823
rect 631 1817 635 1818
rect 727 1822 731 1823
rect 727 1817 731 1818
rect 759 1822 763 1823
rect 759 1817 763 1818
rect 887 1822 891 1823
rect 887 1817 891 1818
rect 1023 1822 1027 1823
rect 1023 1817 1027 1818
rect 1047 1822 1051 1823
rect 1047 1817 1051 1818
rect 1151 1822 1155 1823
rect 1151 1817 1155 1818
rect 1199 1822 1203 1823
rect 1199 1817 1203 1818
rect 1279 1822 1283 1823
rect 1279 1817 1283 1818
rect 1351 1822 1355 1823
rect 1351 1817 1355 1818
rect 1407 1822 1411 1823
rect 1407 1817 1411 1818
rect 1511 1822 1515 1823
rect 1511 1817 1515 1818
rect 1535 1822 1539 1823
rect 1535 1817 1539 1818
rect 1671 1822 1675 1823
rect 1671 1817 1675 1818
rect 1767 1822 1771 1823
rect 1807 1821 1811 1822
rect 2015 1826 2019 1827
rect 2015 1821 2019 1822
rect 2103 1826 2107 1827
rect 2103 1821 2107 1822
rect 2111 1826 2115 1827
rect 2111 1821 2115 1822
rect 2191 1826 2195 1827
rect 2191 1821 2195 1822
rect 2215 1826 2219 1827
rect 2215 1821 2219 1822
rect 2279 1826 2283 1827
rect 2279 1821 2283 1822
rect 2327 1826 2331 1827
rect 2327 1821 2331 1822
rect 2367 1826 2371 1827
rect 2367 1821 2371 1822
rect 2439 1826 2443 1827
rect 2439 1821 2443 1822
rect 2455 1826 2459 1827
rect 2455 1821 2459 1822
rect 2543 1826 2547 1827
rect 2543 1821 2547 1822
rect 2631 1826 2635 1827
rect 2631 1821 2635 1822
rect 2647 1826 2651 1827
rect 2647 1821 2651 1822
rect 2719 1826 2723 1827
rect 2719 1821 2723 1822
rect 2759 1826 2763 1827
rect 2759 1821 2763 1822
rect 2807 1826 2811 1827
rect 2807 1821 2811 1822
rect 2871 1826 2875 1827
rect 2871 1821 2875 1822
rect 2895 1826 2899 1827
rect 2895 1821 2899 1822
rect 2983 1826 2987 1827
rect 2983 1821 2987 1822
rect 3463 1826 3467 1827
rect 3463 1821 3467 1822
rect 1767 1817 1771 1818
rect 112 1801 114 1817
rect 110 1800 116 1801
rect 512 1800 514 1817
rect 632 1800 634 1817
rect 760 1800 762 1817
rect 888 1800 890 1817
rect 1024 1800 1026 1817
rect 1152 1800 1154 1817
rect 1280 1800 1282 1817
rect 1408 1800 1410 1817
rect 1536 1800 1538 1817
rect 1672 1800 1674 1817
rect 1768 1801 1770 1817
rect 1808 1805 1810 1821
rect 1806 1804 1812 1805
rect 2104 1804 2106 1821
rect 2192 1804 2194 1821
rect 2280 1804 2282 1821
rect 2368 1804 2370 1821
rect 2456 1804 2458 1821
rect 2544 1804 2546 1821
rect 2632 1804 2634 1821
rect 2720 1804 2722 1821
rect 2808 1804 2810 1821
rect 2896 1804 2898 1821
rect 3464 1805 3466 1821
rect 3462 1804 3468 1805
rect 1766 1800 1772 1801
rect 110 1796 111 1800
rect 115 1796 116 1800
rect 110 1795 116 1796
rect 510 1799 516 1800
rect 510 1795 511 1799
rect 515 1795 516 1799
rect 510 1794 516 1795
rect 630 1799 636 1800
rect 630 1795 631 1799
rect 635 1795 636 1799
rect 630 1794 636 1795
rect 758 1799 764 1800
rect 758 1795 759 1799
rect 763 1795 764 1799
rect 758 1794 764 1795
rect 886 1799 892 1800
rect 886 1795 887 1799
rect 891 1795 892 1799
rect 886 1794 892 1795
rect 1022 1799 1028 1800
rect 1022 1795 1023 1799
rect 1027 1795 1028 1799
rect 1022 1794 1028 1795
rect 1150 1799 1156 1800
rect 1150 1795 1151 1799
rect 1155 1795 1156 1799
rect 1150 1794 1156 1795
rect 1278 1799 1284 1800
rect 1278 1795 1279 1799
rect 1283 1795 1284 1799
rect 1278 1794 1284 1795
rect 1406 1799 1412 1800
rect 1406 1795 1407 1799
rect 1411 1795 1412 1799
rect 1406 1794 1412 1795
rect 1534 1799 1540 1800
rect 1534 1795 1535 1799
rect 1539 1795 1540 1799
rect 1534 1794 1540 1795
rect 1670 1799 1676 1800
rect 1670 1795 1671 1799
rect 1675 1795 1676 1799
rect 1766 1796 1767 1800
rect 1771 1796 1772 1800
rect 1806 1800 1807 1804
rect 1811 1800 1812 1804
rect 1806 1799 1812 1800
rect 2102 1803 2108 1804
rect 2102 1799 2103 1803
rect 2107 1799 2108 1803
rect 2102 1798 2108 1799
rect 2190 1803 2196 1804
rect 2190 1799 2191 1803
rect 2195 1799 2196 1803
rect 2190 1798 2196 1799
rect 2278 1803 2284 1804
rect 2278 1799 2279 1803
rect 2283 1799 2284 1803
rect 2278 1798 2284 1799
rect 2366 1803 2372 1804
rect 2366 1799 2367 1803
rect 2371 1799 2372 1803
rect 2366 1798 2372 1799
rect 2454 1803 2460 1804
rect 2454 1799 2455 1803
rect 2459 1799 2460 1803
rect 2454 1798 2460 1799
rect 2542 1803 2548 1804
rect 2542 1799 2543 1803
rect 2547 1799 2548 1803
rect 2542 1798 2548 1799
rect 2630 1803 2636 1804
rect 2630 1799 2631 1803
rect 2635 1799 2636 1803
rect 2630 1798 2636 1799
rect 2718 1803 2724 1804
rect 2718 1799 2719 1803
rect 2723 1799 2724 1803
rect 2718 1798 2724 1799
rect 2806 1803 2812 1804
rect 2806 1799 2807 1803
rect 2811 1799 2812 1803
rect 2806 1798 2812 1799
rect 2894 1803 2900 1804
rect 2894 1799 2895 1803
rect 2899 1799 2900 1803
rect 3462 1800 3463 1804
rect 3467 1800 3468 1804
rect 3462 1799 3468 1800
rect 2894 1798 2900 1799
rect 1766 1795 1772 1796
rect 1670 1794 1676 1795
rect 1806 1787 1812 1788
rect 110 1783 116 1784
rect 110 1779 111 1783
rect 115 1779 116 1783
rect 1766 1783 1772 1784
rect 110 1778 116 1779
rect 510 1780 516 1781
rect 112 1755 114 1778
rect 510 1776 511 1780
rect 515 1776 516 1780
rect 510 1775 516 1776
rect 630 1780 636 1781
rect 630 1776 631 1780
rect 635 1776 636 1780
rect 630 1775 636 1776
rect 758 1780 764 1781
rect 758 1776 759 1780
rect 763 1776 764 1780
rect 758 1775 764 1776
rect 886 1780 892 1781
rect 886 1776 887 1780
rect 891 1776 892 1780
rect 886 1775 892 1776
rect 1022 1780 1028 1781
rect 1022 1776 1023 1780
rect 1027 1776 1028 1780
rect 1022 1775 1028 1776
rect 1150 1780 1156 1781
rect 1150 1776 1151 1780
rect 1155 1776 1156 1780
rect 1150 1775 1156 1776
rect 1278 1780 1284 1781
rect 1278 1776 1279 1780
rect 1283 1776 1284 1780
rect 1278 1775 1284 1776
rect 1406 1780 1412 1781
rect 1406 1776 1407 1780
rect 1411 1776 1412 1780
rect 1406 1775 1412 1776
rect 1534 1780 1540 1781
rect 1534 1776 1535 1780
rect 1539 1776 1540 1780
rect 1534 1775 1540 1776
rect 1670 1780 1676 1781
rect 1670 1776 1671 1780
rect 1675 1776 1676 1780
rect 1766 1779 1767 1783
rect 1771 1779 1772 1783
rect 1806 1783 1807 1787
rect 1811 1783 1812 1787
rect 3462 1787 3468 1788
rect 1806 1782 1812 1783
rect 2102 1784 2108 1785
rect 1766 1778 1772 1779
rect 1670 1775 1676 1776
rect 512 1755 514 1775
rect 632 1755 634 1775
rect 760 1755 762 1775
rect 888 1755 890 1775
rect 1024 1755 1026 1775
rect 1152 1755 1154 1775
rect 1280 1755 1282 1775
rect 1408 1755 1410 1775
rect 1536 1755 1538 1775
rect 1672 1755 1674 1775
rect 1768 1755 1770 1778
rect 111 1754 115 1755
rect 111 1749 115 1750
rect 439 1754 443 1755
rect 439 1749 443 1750
rect 511 1754 515 1755
rect 511 1749 515 1750
rect 535 1754 539 1755
rect 535 1749 539 1750
rect 631 1754 635 1755
rect 631 1749 635 1750
rect 639 1754 643 1755
rect 639 1749 643 1750
rect 743 1754 747 1755
rect 743 1749 747 1750
rect 759 1754 763 1755
rect 759 1749 763 1750
rect 847 1754 851 1755
rect 847 1749 851 1750
rect 887 1754 891 1755
rect 887 1749 891 1750
rect 951 1754 955 1755
rect 951 1749 955 1750
rect 1023 1754 1027 1755
rect 1023 1749 1027 1750
rect 1055 1754 1059 1755
rect 1055 1749 1059 1750
rect 1151 1754 1155 1755
rect 1151 1749 1155 1750
rect 1159 1754 1163 1755
rect 1159 1749 1163 1750
rect 1271 1754 1275 1755
rect 1271 1749 1275 1750
rect 1279 1754 1283 1755
rect 1279 1749 1283 1750
rect 1383 1754 1387 1755
rect 1383 1749 1387 1750
rect 1407 1754 1411 1755
rect 1407 1749 1411 1750
rect 1535 1754 1539 1755
rect 1535 1749 1539 1750
rect 1671 1754 1675 1755
rect 1671 1749 1675 1750
rect 1767 1754 1771 1755
rect 1808 1751 1810 1782
rect 2102 1780 2103 1784
rect 2107 1780 2108 1784
rect 2102 1779 2108 1780
rect 2190 1784 2196 1785
rect 2190 1780 2191 1784
rect 2195 1780 2196 1784
rect 2190 1779 2196 1780
rect 2278 1784 2284 1785
rect 2278 1780 2279 1784
rect 2283 1780 2284 1784
rect 2278 1779 2284 1780
rect 2366 1784 2372 1785
rect 2366 1780 2367 1784
rect 2371 1780 2372 1784
rect 2366 1779 2372 1780
rect 2454 1784 2460 1785
rect 2454 1780 2455 1784
rect 2459 1780 2460 1784
rect 2454 1779 2460 1780
rect 2542 1784 2548 1785
rect 2542 1780 2543 1784
rect 2547 1780 2548 1784
rect 2542 1779 2548 1780
rect 2630 1784 2636 1785
rect 2630 1780 2631 1784
rect 2635 1780 2636 1784
rect 2630 1779 2636 1780
rect 2718 1784 2724 1785
rect 2718 1780 2719 1784
rect 2723 1780 2724 1784
rect 2718 1779 2724 1780
rect 2806 1784 2812 1785
rect 2806 1780 2807 1784
rect 2811 1780 2812 1784
rect 2806 1779 2812 1780
rect 2894 1784 2900 1785
rect 2894 1780 2895 1784
rect 2899 1780 2900 1784
rect 3462 1783 3463 1787
rect 3467 1783 3468 1787
rect 3462 1782 3468 1783
rect 2894 1779 2900 1780
rect 2104 1751 2106 1779
rect 2192 1751 2194 1779
rect 2280 1751 2282 1779
rect 2368 1751 2370 1779
rect 2456 1751 2458 1779
rect 2544 1751 2546 1779
rect 2632 1751 2634 1779
rect 2720 1751 2722 1779
rect 2808 1751 2810 1779
rect 2896 1751 2898 1779
rect 3464 1751 3466 1782
rect 1767 1749 1771 1750
rect 1807 1750 1811 1751
rect 112 1730 114 1749
rect 440 1733 442 1749
rect 536 1733 538 1749
rect 640 1733 642 1749
rect 744 1733 746 1749
rect 848 1733 850 1749
rect 952 1733 954 1749
rect 1056 1733 1058 1749
rect 1160 1733 1162 1749
rect 1272 1733 1274 1749
rect 1384 1733 1386 1749
rect 438 1732 444 1733
rect 110 1729 116 1730
rect 110 1725 111 1729
rect 115 1725 116 1729
rect 438 1728 439 1732
rect 443 1728 444 1732
rect 438 1727 444 1728
rect 534 1732 540 1733
rect 534 1728 535 1732
rect 539 1728 540 1732
rect 534 1727 540 1728
rect 638 1732 644 1733
rect 638 1728 639 1732
rect 643 1728 644 1732
rect 638 1727 644 1728
rect 742 1732 748 1733
rect 742 1728 743 1732
rect 747 1728 748 1732
rect 742 1727 748 1728
rect 846 1732 852 1733
rect 846 1728 847 1732
rect 851 1728 852 1732
rect 846 1727 852 1728
rect 950 1732 956 1733
rect 950 1728 951 1732
rect 955 1728 956 1732
rect 950 1727 956 1728
rect 1054 1732 1060 1733
rect 1054 1728 1055 1732
rect 1059 1728 1060 1732
rect 1054 1727 1060 1728
rect 1158 1732 1164 1733
rect 1158 1728 1159 1732
rect 1163 1728 1164 1732
rect 1158 1727 1164 1728
rect 1270 1732 1276 1733
rect 1270 1728 1271 1732
rect 1275 1728 1276 1732
rect 1270 1727 1276 1728
rect 1382 1732 1388 1733
rect 1382 1728 1383 1732
rect 1387 1728 1388 1732
rect 1768 1730 1770 1749
rect 1807 1745 1811 1746
rect 2103 1750 2107 1751
rect 2103 1745 2107 1746
rect 2143 1750 2147 1751
rect 2143 1745 2147 1746
rect 2191 1750 2195 1751
rect 2191 1745 2195 1746
rect 2231 1750 2235 1751
rect 2231 1745 2235 1746
rect 2279 1750 2283 1751
rect 2279 1745 2283 1746
rect 2319 1750 2323 1751
rect 2319 1745 2323 1746
rect 2367 1750 2371 1751
rect 2367 1745 2371 1746
rect 2407 1750 2411 1751
rect 2407 1745 2411 1746
rect 2455 1750 2459 1751
rect 2455 1745 2459 1746
rect 2495 1750 2499 1751
rect 2495 1745 2499 1746
rect 2543 1750 2547 1751
rect 2543 1745 2547 1746
rect 2583 1750 2587 1751
rect 2583 1745 2587 1746
rect 2631 1750 2635 1751
rect 2631 1745 2635 1746
rect 2671 1750 2675 1751
rect 2671 1745 2675 1746
rect 2719 1750 2723 1751
rect 2719 1745 2723 1746
rect 2759 1750 2763 1751
rect 2759 1745 2763 1746
rect 2807 1750 2811 1751
rect 2807 1745 2811 1746
rect 2847 1750 2851 1751
rect 2847 1745 2851 1746
rect 2895 1750 2899 1751
rect 2895 1745 2899 1746
rect 3463 1750 3467 1751
rect 3463 1745 3467 1746
rect 1382 1727 1388 1728
rect 1766 1729 1772 1730
rect 110 1724 116 1725
rect 1766 1725 1767 1729
rect 1771 1725 1772 1729
rect 1808 1726 1810 1745
rect 2144 1729 2146 1745
rect 2232 1729 2234 1745
rect 2320 1729 2322 1745
rect 2408 1729 2410 1745
rect 2496 1729 2498 1745
rect 2584 1729 2586 1745
rect 2672 1729 2674 1745
rect 2760 1729 2762 1745
rect 2848 1729 2850 1745
rect 2142 1728 2148 1729
rect 1766 1724 1772 1725
rect 1806 1725 1812 1726
rect 1806 1721 1807 1725
rect 1811 1721 1812 1725
rect 2142 1724 2143 1728
rect 2147 1724 2148 1728
rect 2142 1723 2148 1724
rect 2230 1728 2236 1729
rect 2230 1724 2231 1728
rect 2235 1724 2236 1728
rect 2230 1723 2236 1724
rect 2318 1728 2324 1729
rect 2318 1724 2319 1728
rect 2323 1724 2324 1728
rect 2318 1723 2324 1724
rect 2406 1728 2412 1729
rect 2406 1724 2407 1728
rect 2411 1724 2412 1728
rect 2406 1723 2412 1724
rect 2494 1728 2500 1729
rect 2494 1724 2495 1728
rect 2499 1724 2500 1728
rect 2494 1723 2500 1724
rect 2582 1728 2588 1729
rect 2582 1724 2583 1728
rect 2587 1724 2588 1728
rect 2582 1723 2588 1724
rect 2670 1728 2676 1729
rect 2670 1724 2671 1728
rect 2675 1724 2676 1728
rect 2670 1723 2676 1724
rect 2758 1728 2764 1729
rect 2758 1724 2759 1728
rect 2763 1724 2764 1728
rect 2758 1723 2764 1724
rect 2846 1728 2852 1729
rect 2846 1724 2847 1728
rect 2851 1724 2852 1728
rect 3464 1726 3466 1745
rect 2846 1723 2852 1724
rect 3462 1725 3468 1726
rect 1806 1720 1812 1721
rect 3462 1721 3463 1725
rect 3467 1721 3468 1725
rect 3462 1720 3468 1721
rect 438 1713 444 1714
rect 110 1712 116 1713
rect 110 1708 111 1712
rect 115 1708 116 1712
rect 438 1709 439 1713
rect 443 1709 444 1713
rect 438 1708 444 1709
rect 534 1713 540 1714
rect 534 1709 535 1713
rect 539 1709 540 1713
rect 534 1708 540 1709
rect 638 1713 644 1714
rect 638 1709 639 1713
rect 643 1709 644 1713
rect 638 1708 644 1709
rect 742 1713 748 1714
rect 742 1709 743 1713
rect 747 1709 748 1713
rect 742 1708 748 1709
rect 846 1713 852 1714
rect 846 1709 847 1713
rect 851 1709 852 1713
rect 846 1708 852 1709
rect 950 1713 956 1714
rect 950 1709 951 1713
rect 955 1709 956 1713
rect 950 1708 956 1709
rect 1054 1713 1060 1714
rect 1054 1709 1055 1713
rect 1059 1709 1060 1713
rect 1054 1708 1060 1709
rect 1158 1713 1164 1714
rect 1158 1709 1159 1713
rect 1163 1709 1164 1713
rect 1158 1708 1164 1709
rect 1270 1713 1276 1714
rect 1270 1709 1271 1713
rect 1275 1709 1276 1713
rect 1270 1708 1276 1709
rect 1382 1713 1388 1714
rect 1382 1709 1383 1713
rect 1387 1709 1388 1713
rect 1382 1708 1388 1709
rect 1766 1712 1772 1713
rect 1766 1708 1767 1712
rect 1771 1708 1772 1712
rect 2142 1709 2148 1710
rect 110 1707 116 1708
rect 112 1687 114 1707
rect 440 1687 442 1708
rect 536 1687 538 1708
rect 640 1687 642 1708
rect 744 1687 746 1708
rect 848 1687 850 1708
rect 952 1687 954 1708
rect 1056 1687 1058 1708
rect 1160 1687 1162 1708
rect 1272 1687 1274 1708
rect 1384 1687 1386 1708
rect 1766 1707 1772 1708
rect 1806 1708 1812 1709
rect 1768 1687 1770 1707
rect 1806 1704 1807 1708
rect 1811 1704 1812 1708
rect 2142 1705 2143 1709
rect 2147 1705 2148 1709
rect 2142 1704 2148 1705
rect 2230 1709 2236 1710
rect 2230 1705 2231 1709
rect 2235 1705 2236 1709
rect 2230 1704 2236 1705
rect 2318 1709 2324 1710
rect 2318 1705 2319 1709
rect 2323 1705 2324 1709
rect 2318 1704 2324 1705
rect 2406 1709 2412 1710
rect 2406 1705 2407 1709
rect 2411 1705 2412 1709
rect 2406 1704 2412 1705
rect 2494 1709 2500 1710
rect 2494 1705 2495 1709
rect 2499 1705 2500 1709
rect 2494 1704 2500 1705
rect 2582 1709 2588 1710
rect 2582 1705 2583 1709
rect 2587 1705 2588 1709
rect 2582 1704 2588 1705
rect 2670 1709 2676 1710
rect 2670 1705 2671 1709
rect 2675 1705 2676 1709
rect 2670 1704 2676 1705
rect 2758 1709 2764 1710
rect 2758 1705 2759 1709
rect 2763 1705 2764 1709
rect 2758 1704 2764 1705
rect 2846 1709 2852 1710
rect 2846 1705 2847 1709
rect 2851 1705 2852 1709
rect 2846 1704 2852 1705
rect 3462 1708 3468 1709
rect 3462 1704 3463 1708
rect 3467 1704 3468 1708
rect 1806 1703 1812 1704
rect 111 1686 115 1687
rect 111 1681 115 1682
rect 399 1686 403 1687
rect 399 1681 403 1682
rect 439 1686 443 1687
rect 439 1681 443 1682
rect 487 1686 491 1687
rect 487 1681 491 1682
rect 535 1686 539 1687
rect 535 1681 539 1682
rect 575 1686 579 1687
rect 575 1681 579 1682
rect 639 1686 643 1687
rect 639 1681 643 1682
rect 663 1686 667 1687
rect 663 1681 667 1682
rect 743 1686 747 1687
rect 743 1681 747 1682
rect 759 1686 763 1687
rect 759 1681 763 1682
rect 847 1686 851 1687
rect 847 1681 851 1682
rect 855 1686 859 1687
rect 855 1681 859 1682
rect 951 1686 955 1687
rect 951 1681 955 1682
rect 1047 1686 1051 1687
rect 1047 1681 1051 1682
rect 1055 1686 1059 1687
rect 1055 1681 1059 1682
rect 1143 1686 1147 1687
rect 1143 1681 1147 1682
rect 1159 1686 1163 1687
rect 1159 1681 1163 1682
rect 1271 1686 1275 1687
rect 1271 1681 1275 1682
rect 1383 1686 1387 1687
rect 1383 1681 1387 1682
rect 1767 1686 1771 1687
rect 1808 1683 1810 1703
rect 2144 1683 2146 1704
rect 2232 1683 2234 1704
rect 2320 1683 2322 1704
rect 2408 1683 2410 1704
rect 2496 1683 2498 1704
rect 2584 1683 2586 1704
rect 2672 1683 2674 1704
rect 2760 1683 2762 1704
rect 2848 1683 2850 1704
rect 3462 1703 3468 1704
rect 3464 1683 3466 1703
rect 1767 1681 1771 1682
rect 1807 1682 1811 1683
rect 112 1665 114 1681
rect 110 1664 116 1665
rect 400 1664 402 1681
rect 488 1664 490 1681
rect 576 1664 578 1681
rect 664 1664 666 1681
rect 760 1664 762 1681
rect 856 1664 858 1681
rect 952 1664 954 1681
rect 1048 1664 1050 1681
rect 1144 1664 1146 1681
rect 1768 1665 1770 1681
rect 1807 1677 1811 1678
rect 2103 1682 2107 1683
rect 2103 1677 2107 1678
rect 2143 1682 2147 1683
rect 2143 1677 2147 1678
rect 2191 1682 2195 1683
rect 2191 1677 2195 1678
rect 2231 1682 2235 1683
rect 2231 1677 2235 1678
rect 2279 1682 2283 1683
rect 2279 1677 2283 1678
rect 2319 1682 2323 1683
rect 2319 1677 2323 1678
rect 2367 1682 2371 1683
rect 2367 1677 2371 1678
rect 2407 1682 2411 1683
rect 2407 1677 2411 1678
rect 2455 1682 2459 1683
rect 2455 1677 2459 1678
rect 2495 1682 2499 1683
rect 2495 1677 2499 1678
rect 2543 1682 2547 1683
rect 2543 1677 2547 1678
rect 2583 1682 2587 1683
rect 2583 1677 2587 1678
rect 2631 1682 2635 1683
rect 2631 1677 2635 1678
rect 2671 1682 2675 1683
rect 2671 1677 2675 1678
rect 2719 1682 2723 1683
rect 2719 1677 2723 1678
rect 2759 1682 2763 1683
rect 2759 1677 2763 1678
rect 2807 1682 2811 1683
rect 2807 1677 2811 1678
rect 2847 1682 2851 1683
rect 2847 1677 2851 1678
rect 2895 1682 2899 1683
rect 2895 1677 2899 1678
rect 3463 1682 3467 1683
rect 3463 1677 3467 1678
rect 1766 1664 1772 1665
rect 110 1660 111 1664
rect 115 1660 116 1664
rect 110 1659 116 1660
rect 398 1663 404 1664
rect 398 1659 399 1663
rect 403 1659 404 1663
rect 398 1658 404 1659
rect 486 1663 492 1664
rect 486 1659 487 1663
rect 491 1659 492 1663
rect 486 1658 492 1659
rect 574 1663 580 1664
rect 574 1659 575 1663
rect 579 1659 580 1663
rect 574 1658 580 1659
rect 662 1663 668 1664
rect 662 1659 663 1663
rect 667 1659 668 1663
rect 662 1658 668 1659
rect 758 1663 764 1664
rect 758 1659 759 1663
rect 763 1659 764 1663
rect 758 1658 764 1659
rect 854 1663 860 1664
rect 854 1659 855 1663
rect 859 1659 860 1663
rect 854 1658 860 1659
rect 950 1663 956 1664
rect 950 1659 951 1663
rect 955 1659 956 1663
rect 950 1658 956 1659
rect 1046 1663 1052 1664
rect 1046 1659 1047 1663
rect 1051 1659 1052 1663
rect 1046 1658 1052 1659
rect 1142 1663 1148 1664
rect 1142 1659 1143 1663
rect 1147 1659 1148 1663
rect 1766 1660 1767 1664
rect 1771 1660 1772 1664
rect 1808 1661 1810 1677
rect 1766 1659 1772 1660
rect 1806 1660 1812 1661
rect 2104 1660 2106 1677
rect 2192 1660 2194 1677
rect 2280 1660 2282 1677
rect 2368 1660 2370 1677
rect 2456 1660 2458 1677
rect 2544 1660 2546 1677
rect 2632 1660 2634 1677
rect 2720 1660 2722 1677
rect 2808 1660 2810 1677
rect 2896 1660 2898 1677
rect 3464 1661 3466 1677
rect 3462 1660 3468 1661
rect 1142 1658 1148 1659
rect 1806 1656 1807 1660
rect 1811 1656 1812 1660
rect 1806 1655 1812 1656
rect 2102 1659 2108 1660
rect 2102 1655 2103 1659
rect 2107 1655 2108 1659
rect 2102 1654 2108 1655
rect 2190 1659 2196 1660
rect 2190 1655 2191 1659
rect 2195 1655 2196 1659
rect 2190 1654 2196 1655
rect 2278 1659 2284 1660
rect 2278 1655 2279 1659
rect 2283 1655 2284 1659
rect 2278 1654 2284 1655
rect 2366 1659 2372 1660
rect 2366 1655 2367 1659
rect 2371 1655 2372 1659
rect 2366 1654 2372 1655
rect 2454 1659 2460 1660
rect 2454 1655 2455 1659
rect 2459 1655 2460 1659
rect 2454 1654 2460 1655
rect 2542 1659 2548 1660
rect 2542 1655 2543 1659
rect 2547 1655 2548 1659
rect 2542 1654 2548 1655
rect 2630 1659 2636 1660
rect 2630 1655 2631 1659
rect 2635 1655 2636 1659
rect 2630 1654 2636 1655
rect 2718 1659 2724 1660
rect 2718 1655 2719 1659
rect 2723 1655 2724 1659
rect 2718 1654 2724 1655
rect 2806 1659 2812 1660
rect 2806 1655 2807 1659
rect 2811 1655 2812 1659
rect 2806 1654 2812 1655
rect 2894 1659 2900 1660
rect 2894 1655 2895 1659
rect 2899 1655 2900 1659
rect 3462 1656 3463 1660
rect 3467 1656 3468 1660
rect 3462 1655 3468 1656
rect 2894 1654 2900 1655
rect 110 1647 116 1648
rect 110 1643 111 1647
rect 115 1643 116 1647
rect 1766 1647 1772 1648
rect 110 1642 116 1643
rect 398 1644 404 1645
rect 112 1619 114 1642
rect 398 1640 399 1644
rect 403 1640 404 1644
rect 398 1639 404 1640
rect 486 1644 492 1645
rect 486 1640 487 1644
rect 491 1640 492 1644
rect 486 1639 492 1640
rect 574 1644 580 1645
rect 574 1640 575 1644
rect 579 1640 580 1644
rect 574 1639 580 1640
rect 662 1644 668 1645
rect 662 1640 663 1644
rect 667 1640 668 1644
rect 662 1639 668 1640
rect 758 1644 764 1645
rect 758 1640 759 1644
rect 763 1640 764 1644
rect 758 1639 764 1640
rect 854 1644 860 1645
rect 854 1640 855 1644
rect 859 1640 860 1644
rect 854 1639 860 1640
rect 950 1644 956 1645
rect 950 1640 951 1644
rect 955 1640 956 1644
rect 950 1639 956 1640
rect 1046 1644 1052 1645
rect 1046 1640 1047 1644
rect 1051 1640 1052 1644
rect 1046 1639 1052 1640
rect 1142 1644 1148 1645
rect 1142 1640 1143 1644
rect 1147 1640 1148 1644
rect 1766 1643 1767 1647
rect 1771 1643 1772 1647
rect 1766 1642 1772 1643
rect 1806 1643 1812 1644
rect 1142 1639 1148 1640
rect 400 1619 402 1639
rect 488 1619 490 1639
rect 576 1619 578 1639
rect 664 1619 666 1639
rect 760 1619 762 1639
rect 856 1619 858 1639
rect 952 1619 954 1639
rect 1048 1619 1050 1639
rect 1144 1619 1146 1639
rect 1768 1619 1770 1642
rect 1806 1639 1807 1643
rect 1811 1639 1812 1643
rect 3462 1643 3468 1644
rect 1806 1638 1812 1639
rect 2102 1640 2108 1641
rect 111 1618 115 1619
rect 111 1613 115 1614
rect 279 1618 283 1619
rect 279 1613 283 1614
rect 383 1618 387 1619
rect 383 1613 387 1614
rect 399 1618 403 1619
rect 399 1613 403 1614
rect 487 1618 491 1619
rect 487 1613 491 1614
rect 495 1618 499 1619
rect 495 1613 499 1614
rect 575 1618 579 1619
rect 575 1613 579 1614
rect 607 1618 611 1619
rect 607 1613 611 1614
rect 663 1618 667 1619
rect 663 1613 667 1614
rect 719 1618 723 1619
rect 719 1613 723 1614
rect 759 1618 763 1619
rect 759 1613 763 1614
rect 831 1618 835 1619
rect 831 1613 835 1614
rect 855 1618 859 1619
rect 855 1613 859 1614
rect 943 1618 947 1619
rect 943 1613 947 1614
rect 951 1618 955 1619
rect 951 1613 955 1614
rect 1047 1618 1051 1619
rect 1047 1613 1051 1614
rect 1055 1618 1059 1619
rect 1055 1613 1059 1614
rect 1143 1618 1147 1619
rect 1143 1613 1147 1614
rect 1167 1618 1171 1619
rect 1167 1613 1171 1614
rect 1279 1618 1283 1619
rect 1279 1613 1283 1614
rect 1767 1618 1771 1619
rect 1808 1615 1810 1638
rect 2102 1636 2103 1640
rect 2107 1636 2108 1640
rect 2102 1635 2108 1636
rect 2190 1640 2196 1641
rect 2190 1636 2191 1640
rect 2195 1636 2196 1640
rect 2190 1635 2196 1636
rect 2278 1640 2284 1641
rect 2278 1636 2279 1640
rect 2283 1636 2284 1640
rect 2278 1635 2284 1636
rect 2366 1640 2372 1641
rect 2366 1636 2367 1640
rect 2371 1636 2372 1640
rect 2366 1635 2372 1636
rect 2454 1640 2460 1641
rect 2454 1636 2455 1640
rect 2459 1636 2460 1640
rect 2454 1635 2460 1636
rect 2542 1640 2548 1641
rect 2542 1636 2543 1640
rect 2547 1636 2548 1640
rect 2542 1635 2548 1636
rect 2630 1640 2636 1641
rect 2630 1636 2631 1640
rect 2635 1636 2636 1640
rect 2630 1635 2636 1636
rect 2718 1640 2724 1641
rect 2718 1636 2719 1640
rect 2723 1636 2724 1640
rect 2718 1635 2724 1636
rect 2806 1640 2812 1641
rect 2806 1636 2807 1640
rect 2811 1636 2812 1640
rect 2806 1635 2812 1636
rect 2894 1640 2900 1641
rect 2894 1636 2895 1640
rect 2899 1636 2900 1640
rect 3462 1639 3463 1643
rect 3467 1639 3468 1643
rect 3462 1638 3468 1639
rect 2894 1635 2900 1636
rect 2104 1615 2106 1635
rect 2192 1615 2194 1635
rect 2280 1615 2282 1635
rect 2368 1615 2370 1635
rect 2456 1615 2458 1635
rect 2544 1615 2546 1635
rect 2632 1615 2634 1635
rect 2720 1615 2722 1635
rect 2808 1615 2810 1635
rect 2896 1615 2898 1635
rect 3464 1615 3466 1638
rect 1767 1613 1771 1614
rect 1807 1614 1811 1615
rect 112 1594 114 1613
rect 280 1597 282 1613
rect 384 1597 386 1613
rect 496 1597 498 1613
rect 608 1597 610 1613
rect 720 1597 722 1613
rect 832 1597 834 1613
rect 944 1597 946 1613
rect 1056 1597 1058 1613
rect 1168 1597 1170 1613
rect 1280 1597 1282 1613
rect 278 1596 284 1597
rect 110 1593 116 1594
rect 110 1589 111 1593
rect 115 1589 116 1593
rect 278 1592 279 1596
rect 283 1592 284 1596
rect 278 1591 284 1592
rect 382 1596 388 1597
rect 382 1592 383 1596
rect 387 1592 388 1596
rect 382 1591 388 1592
rect 494 1596 500 1597
rect 494 1592 495 1596
rect 499 1592 500 1596
rect 494 1591 500 1592
rect 606 1596 612 1597
rect 606 1592 607 1596
rect 611 1592 612 1596
rect 606 1591 612 1592
rect 718 1596 724 1597
rect 718 1592 719 1596
rect 723 1592 724 1596
rect 718 1591 724 1592
rect 830 1596 836 1597
rect 830 1592 831 1596
rect 835 1592 836 1596
rect 830 1591 836 1592
rect 942 1596 948 1597
rect 942 1592 943 1596
rect 947 1592 948 1596
rect 942 1591 948 1592
rect 1054 1596 1060 1597
rect 1054 1592 1055 1596
rect 1059 1592 1060 1596
rect 1054 1591 1060 1592
rect 1166 1596 1172 1597
rect 1166 1592 1167 1596
rect 1171 1592 1172 1596
rect 1166 1591 1172 1592
rect 1278 1596 1284 1597
rect 1278 1592 1279 1596
rect 1283 1592 1284 1596
rect 1768 1594 1770 1613
rect 1807 1609 1811 1610
rect 2063 1614 2067 1615
rect 2063 1609 2067 1610
rect 2103 1614 2107 1615
rect 2103 1609 2107 1610
rect 2159 1614 2163 1615
rect 2159 1609 2163 1610
rect 2191 1614 2195 1615
rect 2191 1609 2195 1610
rect 2255 1614 2259 1615
rect 2255 1609 2259 1610
rect 2279 1614 2283 1615
rect 2279 1609 2283 1610
rect 2359 1614 2363 1615
rect 2359 1609 2363 1610
rect 2367 1614 2371 1615
rect 2367 1609 2371 1610
rect 2455 1614 2459 1615
rect 2455 1609 2459 1610
rect 2463 1614 2467 1615
rect 2463 1609 2467 1610
rect 2543 1614 2547 1615
rect 2543 1609 2547 1610
rect 2567 1614 2571 1615
rect 2567 1609 2571 1610
rect 2631 1614 2635 1615
rect 2631 1609 2635 1610
rect 2671 1614 2675 1615
rect 2671 1609 2675 1610
rect 2719 1614 2723 1615
rect 2719 1609 2723 1610
rect 2775 1614 2779 1615
rect 2775 1609 2779 1610
rect 2807 1614 2811 1615
rect 2807 1609 2811 1610
rect 2887 1614 2891 1615
rect 2887 1609 2891 1610
rect 2895 1614 2899 1615
rect 2895 1609 2899 1610
rect 3463 1614 3467 1615
rect 3463 1609 3467 1610
rect 1278 1591 1284 1592
rect 1766 1593 1772 1594
rect 110 1588 116 1589
rect 1766 1589 1767 1593
rect 1771 1589 1772 1593
rect 1808 1590 1810 1609
rect 2064 1593 2066 1609
rect 2160 1593 2162 1609
rect 2256 1593 2258 1609
rect 2360 1593 2362 1609
rect 2464 1593 2466 1609
rect 2568 1593 2570 1609
rect 2672 1593 2674 1609
rect 2776 1593 2778 1609
rect 2888 1593 2890 1609
rect 2062 1592 2068 1593
rect 1766 1588 1772 1589
rect 1806 1589 1812 1590
rect 1806 1585 1807 1589
rect 1811 1585 1812 1589
rect 2062 1588 2063 1592
rect 2067 1588 2068 1592
rect 2062 1587 2068 1588
rect 2158 1592 2164 1593
rect 2158 1588 2159 1592
rect 2163 1588 2164 1592
rect 2158 1587 2164 1588
rect 2254 1592 2260 1593
rect 2254 1588 2255 1592
rect 2259 1588 2260 1592
rect 2254 1587 2260 1588
rect 2358 1592 2364 1593
rect 2358 1588 2359 1592
rect 2363 1588 2364 1592
rect 2358 1587 2364 1588
rect 2462 1592 2468 1593
rect 2462 1588 2463 1592
rect 2467 1588 2468 1592
rect 2462 1587 2468 1588
rect 2566 1592 2572 1593
rect 2566 1588 2567 1592
rect 2571 1588 2572 1592
rect 2566 1587 2572 1588
rect 2670 1592 2676 1593
rect 2670 1588 2671 1592
rect 2675 1588 2676 1592
rect 2670 1587 2676 1588
rect 2774 1592 2780 1593
rect 2774 1588 2775 1592
rect 2779 1588 2780 1592
rect 2774 1587 2780 1588
rect 2886 1592 2892 1593
rect 2886 1588 2887 1592
rect 2891 1588 2892 1592
rect 3464 1590 3466 1609
rect 2886 1587 2892 1588
rect 3462 1589 3468 1590
rect 1806 1584 1812 1585
rect 3462 1585 3463 1589
rect 3467 1585 3468 1589
rect 3462 1584 3468 1585
rect 278 1577 284 1578
rect 110 1576 116 1577
rect 110 1572 111 1576
rect 115 1572 116 1576
rect 278 1573 279 1577
rect 283 1573 284 1577
rect 278 1572 284 1573
rect 382 1577 388 1578
rect 382 1573 383 1577
rect 387 1573 388 1577
rect 382 1572 388 1573
rect 494 1577 500 1578
rect 494 1573 495 1577
rect 499 1573 500 1577
rect 494 1572 500 1573
rect 606 1577 612 1578
rect 606 1573 607 1577
rect 611 1573 612 1577
rect 606 1572 612 1573
rect 718 1577 724 1578
rect 718 1573 719 1577
rect 723 1573 724 1577
rect 718 1572 724 1573
rect 830 1577 836 1578
rect 830 1573 831 1577
rect 835 1573 836 1577
rect 830 1572 836 1573
rect 942 1577 948 1578
rect 942 1573 943 1577
rect 947 1573 948 1577
rect 942 1572 948 1573
rect 1054 1577 1060 1578
rect 1054 1573 1055 1577
rect 1059 1573 1060 1577
rect 1054 1572 1060 1573
rect 1166 1577 1172 1578
rect 1166 1573 1167 1577
rect 1171 1573 1172 1577
rect 1166 1572 1172 1573
rect 1278 1577 1284 1578
rect 1278 1573 1279 1577
rect 1283 1573 1284 1577
rect 1278 1572 1284 1573
rect 1766 1576 1772 1577
rect 1766 1572 1767 1576
rect 1771 1572 1772 1576
rect 2062 1573 2068 1574
rect 110 1571 116 1572
rect 112 1547 114 1571
rect 280 1547 282 1572
rect 384 1547 386 1572
rect 496 1547 498 1572
rect 608 1547 610 1572
rect 720 1547 722 1572
rect 832 1547 834 1572
rect 944 1547 946 1572
rect 1056 1547 1058 1572
rect 1168 1547 1170 1572
rect 1280 1547 1282 1572
rect 1766 1571 1772 1572
rect 1806 1572 1812 1573
rect 1768 1547 1770 1571
rect 1806 1568 1807 1572
rect 1811 1568 1812 1572
rect 2062 1569 2063 1573
rect 2067 1569 2068 1573
rect 2062 1568 2068 1569
rect 2158 1573 2164 1574
rect 2158 1569 2159 1573
rect 2163 1569 2164 1573
rect 2158 1568 2164 1569
rect 2254 1573 2260 1574
rect 2254 1569 2255 1573
rect 2259 1569 2260 1573
rect 2254 1568 2260 1569
rect 2358 1573 2364 1574
rect 2358 1569 2359 1573
rect 2363 1569 2364 1573
rect 2358 1568 2364 1569
rect 2462 1573 2468 1574
rect 2462 1569 2463 1573
rect 2467 1569 2468 1573
rect 2462 1568 2468 1569
rect 2566 1573 2572 1574
rect 2566 1569 2567 1573
rect 2571 1569 2572 1573
rect 2566 1568 2572 1569
rect 2670 1573 2676 1574
rect 2670 1569 2671 1573
rect 2675 1569 2676 1573
rect 2670 1568 2676 1569
rect 2774 1573 2780 1574
rect 2774 1569 2775 1573
rect 2779 1569 2780 1573
rect 2774 1568 2780 1569
rect 2886 1573 2892 1574
rect 2886 1569 2887 1573
rect 2891 1569 2892 1573
rect 2886 1568 2892 1569
rect 3462 1572 3468 1573
rect 3462 1568 3463 1572
rect 3467 1568 3468 1572
rect 1806 1567 1812 1568
rect 1808 1551 1810 1567
rect 2064 1551 2066 1568
rect 2160 1551 2162 1568
rect 2256 1551 2258 1568
rect 2360 1551 2362 1568
rect 2464 1551 2466 1568
rect 2568 1551 2570 1568
rect 2672 1551 2674 1568
rect 2776 1551 2778 1568
rect 2888 1551 2890 1568
rect 3462 1567 3468 1568
rect 3464 1551 3466 1567
rect 1807 1550 1811 1551
rect 111 1546 115 1547
rect 111 1541 115 1542
rect 183 1546 187 1547
rect 183 1541 187 1542
rect 279 1546 283 1547
rect 279 1541 283 1542
rect 327 1546 331 1547
rect 327 1541 331 1542
rect 383 1546 387 1547
rect 383 1541 387 1542
rect 471 1546 475 1547
rect 471 1541 475 1542
rect 495 1546 499 1547
rect 495 1541 499 1542
rect 607 1546 611 1547
rect 607 1541 611 1542
rect 623 1546 627 1547
rect 623 1541 627 1542
rect 719 1546 723 1547
rect 719 1541 723 1542
rect 767 1546 771 1547
rect 767 1541 771 1542
rect 831 1546 835 1547
rect 831 1541 835 1542
rect 911 1546 915 1547
rect 911 1541 915 1542
rect 943 1546 947 1547
rect 943 1541 947 1542
rect 1047 1546 1051 1547
rect 1047 1541 1051 1542
rect 1055 1546 1059 1547
rect 1055 1541 1059 1542
rect 1167 1546 1171 1547
rect 1167 1541 1171 1542
rect 1175 1546 1179 1547
rect 1175 1541 1179 1542
rect 1279 1546 1283 1547
rect 1279 1541 1283 1542
rect 1311 1546 1315 1547
rect 1311 1541 1315 1542
rect 1447 1546 1451 1547
rect 1447 1541 1451 1542
rect 1767 1546 1771 1547
rect 1807 1545 1811 1546
rect 1919 1550 1923 1551
rect 1919 1545 1923 1546
rect 2039 1550 2043 1551
rect 2039 1545 2043 1546
rect 2063 1550 2067 1551
rect 2063 1545 2067 1546
rect 2159 1550 2163 1551
rect 2159 1545 2163 1546
rect 2167 1550 2171 1551
rect 2167 1545 2171 1546
rect 2255 1550 2259 1551
rect 2255 1545 2259 1546
rect 2295 1550 2299 1551
rect 2295 1545 2299 1546
rect 2359 1550 2363 1551
rect 2359 1545 2363 1546
rect 2423 1550 2427 1551
rect 2423 1545 2427 1546
rect 2463 1550 2467 1551
rect 2463 1545 2467 1546
rect 2551 1550 2555 1551
rect 2551 1545 2555 1546
rect 2567 1550 2571 1551
rect 2567 1545 2571 1546
rect 2671 1550 2675 1551
rect 2671 1545 2675 1546
rect 2679 1550 2683 1551
rect 2679 1545 2683 1546
rect 2775 1550 2779 1551
rect 2775 1545 2779 1546
rect 2799 1550 2803 1551
rect 2799 1545 2803 1546
rect 2887 1550 2891 1551
rect 2887 1545 2891 1546
rect 2927 1550 2931 1551
rect 2927 1545 2931 1546
rect 3055 1550 3059 1551
rect 3055 1545 3059 1546
rect 3463 1550 3467 1551
rect 3463 1545 3467 1546
rect 1767 1541 1771 1542
rect 112 1525 114 1541
rect 110 1524 116 1525
rect 184 1524 186 1541
rect 328 1524 330 1541
rect 472 1524 474 1541
rect 624 1524 626 1541
rect 768 1524 770 1541
rect 912 1524 914 1541
rect 1048 1524 1050 1541
rect 1176 1524 1178 1541
rect 1312 1524 1314 1541
rect 1448 1524 1450 1541
rect 1768 1525 1770 1541
rect 1808 1529 1810 1545
rect 1806 1528 1812 1529
rect 1920 1528 1922 1545
rect 2040 1528 2042 1545
rect 2168 1528 2170 1545
rect 2296 1528 2298 1545
rect 2424 1528 2426 1545
rect 2552 1528 2554 1545
rect 2680 1528 2682 1545
rect 2800 1528 2802 1545
rect 2928 1528 2930 1545
rect 3056 1528 3058 1545
rect 3464 1529 3466 1545
rect 3462 1528 3468 1529
rect 1766 1524 1772 1525
rect 110 1520 111 1524
rect 115 1520 116 1524
rect 110 1519 116 1520
rect 182 1523 188 1524
rect 182 1519 183 1523
rect 187 1519 188 1523
rect 182 1518 188 1519
rect 326 1523 332 1524
rect 326 1519 327 1523
rect 331 1519 332 1523
rect 326 1518 332 1519
rect 470 1523 476 1524
rect 470 1519 471 1523
rect 475 1519 476 1523
rect 470 1518 476 1519
rect 622 1523 628 1524
rect 622 1519 623 1523
rect 627 1519 628 1523
rect 622 1518 628 1519
rect 766 1523 772 1524
rect 766 1519 767 1523
rect 771 1519 772 1523
rect 766 1518 772 1519
rect 910 1523 916 1524
rect 910 1519 911 1523
rect 915 1519 916 1523
rect 910 1518 916 1519
rect 1046 1523 1052 1524
rect 1046 1519 1047 1523
rect 1051 1519 1052 1523
rect 1046 1518 1052 1519
rect 1174 1523 1180 1524
rect 1174 1519 1175 1523
rect 1179 1519 1180 1523
rect 1174 1518 1180 1519
rect 1310 1523 1316 1524
rect 1310 1519 1311 1523
rect 1315 1519 1316 1523
rect 1310 1518 1316 1519
rect 1446 1523 1452 1524
rect 1446 1519 1447 1523
rect 1451 1519 1452 1523
rect 1766 1520 1767 1524
rect 1771 1520 1772 1524
rect 1806 1524 1807 1528
rect 1811 1524 1812 1528
rect 1806 1523 1812 1524
rect 1918 1527 1924 1528
rect 1918 1523 1919 1527
rect 1923 1523 1924 1527
rect 1918 1522 1924 1523
rect 2038 1527 2044 1528
rect 2038 1523 2039 1527
rect 2043 1523 2044 1527
rect 2038 1522 2044 1523
rect 2166 1527 2172 1528
rect 2166 1523 2167 1527
rect 2171 1523 2172 1527
rect 2166 1522 2172 1523
rect 2294 1527 2300 1528
rect 2294 1523 2295 1527
rect 2299 1523 2300 1527
rect 2294 1522 2300 1523
rect 2422 1527 2428 1528
rect 2422 1523 2423 1527
rect 2427 1523 2428 1527
rect 2422 1522 2428 1523
rect 2550 1527 2556 1528
rect 2550 1523 2551 1527
rect 2555 1523 2556 1527
rect 2550 1522 2556 1523
rect 2678 1527 2684 1528
rect 2678 1523 2679 1527
rect 2683 1523 2684 1527
rect 2678 1522 2684 1523
rect 2798 1527 2804 1528
rect 2798 1523 2799 1527
rect 2803 1523 2804 1527
rect 2798 1522 2804 1523
rect 2926 1527 2932 1528
rect 2926 1523 2927 1527
rect 2931 1523 2932 1527
rect 2926 1522 2932 1523
rect 3054 1527 3060 1528
rect 3054 1523 3055 1527
rect 3059 1523 3060 1527
rect 3462 1524 3463 1528
rect 3467 1524 3468 1528
rect 3462 1523 3468 1524
rect 3054 1522 3060 1523
rect 1766 1519 1772 1520
rect 1446 1518 1452 1519
rect 1806 1511 1812 1512
rect 110 1507 116 1508
rect 110 1503 111 1507
rect 115 1503 116 1507
rect 1766 1507 1772 1508
rect 110 1502 116 1503
rect 182 1504 188 1505
rect 112 1479 114 1502
rect 182 1500 183 1504
rect 187 1500 188 1504
rect 182 1499 188 1500
rect 326 1504 332 1505
rect 326 1500 327 1504
rect 331 1500 332 1504
rect 326 1499 332 1500
rect 470 1504 476 1505
rect 470 1500 471 1504
rect 475 1500 476 1504
rect 470 1499 476 1500
rect 622 1504 628 1505
rect 622 1500 623 1504
rect 627 1500 628 1504
rect 622 1499 628 1500
rect 766 1504 772 1505
rect 766 1500 767 1504
rect 771 1500 772 1504
rect 766 1499 772 1500
rect 910 1504 916 1505
rect 910 1500 911 1504
rect 915 1500 916 1504
rect 910 1499 916 1500
rect 1046 1504 1052 1505
rect 1046 1500 1047 1504
rect 1051 1500 1052 1504
rect 1046 1499 1052 1500
rect 1174 1504 1180 1505
rect 1174 1500 1175 1504
rect 1179 1500 1180 1504
rect 1174 1499 1180 1500
rect 1310 1504 1316 1505
rect 1310 1500 1311 1504
rect 1315 1500 1316 1504
rect 1310 1499 1316 1500
rect 1446 1504 1452 1505
rect 1446 1500 1447 1504
rect 1451 1500 1452 1504
rect 1766 1503 1767 1507
rect 1771 1503 1772 1507
rect 1806 1507 1807 1511
rect 1811 1507 1812 1511
rect 3462 1511 3468 1512
rect 1806 1506 1812 1507
rect 1918 1508 1924 1509
rect 1766 1502 1772 1503
rect 1446 1499 1452 1500
rect 184 1479 186 1499
rect 328 1479 330 1499
rect 472 1479 474 1499
rect 624 1479 626 1499
rect 768 1479 770 1499
rect 912 1479 914 1499
rect 1048 1479 1050 1499
rect 1176 1479 1178 1499
rect 1312 1479 1314 1499
rect 1448 1479 1450 1499
rect 1768 1479 1770 1502
rect 1808 1479 1810 1506
rect 1918 1504 1919 1508
rect 1923 1504 1924 1508
rect 1918 1503 1924 1504
rect 2038 1508 2044 1509
rect 2038 1504 2039 1508
rect 2043 1504 2044 1508
rect 2038 1503 2044 1504
rect 2166 1508 2172 1509
rect 2166 1504 2167 1508
rect 2171 1504 2172 1508
rect 2166 1503 2172 1504
rect 2294 1508 2300 1509
rect 2294 1504 2295 1508
rect 2299 1504 2300 1508
rect 2294 1503 2300 1504
rect 2422 1508 2428 1509
rect 2422 1504 2423 1508
rect 2427 1504 2428 1508
rect 2422 1503 2428 1504
rect 2550 1508 2556 1509
rect 2550 1504 2551 1508
rect 2555 1504 2556 1508
rect 2550 1503 2556 1504
rect 2678 1508 2684 1509
rect 2678 1504 2679 1508
rect 2683 1504 2684 1508
rect 2678 1503 2684 1504
rect 2798 1508 2804 1509
rect 2798 1504 2799 1508
rect 2803 1504 2804 1508
rect 2798 1503 2804 1504
rect 2926 1508 2932 1509
rect 2926 1504 2927 1508
rect 2931 1504 2932 1508
rect 2926 1503 2932 1504
rect 3054 1508 3060 1509
rect 3054 1504 3055 1508
rect 3059 1504 3060 1508
rect 3462 1507 3463 1511
rect 3467 1507 3468 1511
rect 3462 1506 3468 1507
rect 3054 1503 3060 1504
rect 1920 1479 1922 1503
rect 2040 1479 2042 1503
rect 2168 1479 2170 1503
rect 2296 1479 2298 1503
rect 2424 1479 2426 1503
rect 2552 1479 2554 1503
rect 2680 1479 2682 1503
rect 2800 1479 2802 1503
rect 2928 1479 2930 1503
rect 3056 1479 3058 1503
rect 3464 1479 3466 1506
rect 111 1478 115 1479
rect 111 1473 115 1474
rect 159 1478 163 1479
rect 159 1473 163 1474
rect 183 1478 187 1479
rect 183 1473 187 1474
rect 327 1478 331 1479
rect 327 1473 331 1474
rect 375 1478 379 1479
rect 375 1473 379 1474
rect 471 1478 475 1479
rect 471 1473 475 1474
rect 583 1478 587 1479
rect 583 1473 587 1474
rect 623 1478 627 1479
rect 623 1473 627 1474
rect 767 1478 771 1479
rect 767 1473 771 1474
rect 783 1478 787 1479
rect 783 1473 787 1474
rect 911 1478 915 1479
rect 911 1473 915 1474
rect 959 1478 963 1479
rect 959 1473 963 1474
rect 1047 1478 1051 1479
rect 1047 1473 1051 1474
rect 1127 1478 1131 1479
rect 1127 1473 1131 1474
rect 1175 1478 1179 1479
rect 1175 1473 1179 1474
rect 1279 1478 1283 1479
rect 1279 1473 1283 1474
rect 1311 1478 1315 1479
rect 1311 1473 1315 1474
rect 1431 1478 1435 1479
rect 1431 1473 1435 1474
rect 1447 1478 1451 1479
rect 1447 1473 1451 1474
rect 1591 1478 1595 1479
rect 1591 1473 1595 1474
rect 1767 1478 1771 1479
rect 1767 1473 1771 1474
rect 1807 1478 1811 1479
rect 1807 1473 1811 1474
rect 1831 1478 1835 1479
rect 1831 1473 1835 1474
rect 1919 1478 1923 1479
rect 1919 1473 1923 1474
rect 1951 1478 1955 1479
rect 1951 1473 1955 1474
rect 2039 1478 2043 1479
rect 2039 1473 2043 1474
rect 2111 1478 2115 1479
rect 2111 1473 2115 1474
rect 2167 1478 2171 1479
rect 2167 1473 2171 1474
rect 2271 1478 2275 1479
rect 2271 1473 2275 1474
rect 2295 1478 2299 1479
rect 2295 1473 2299 1474
rect 2423 1478 2427 1479
rect 2423 1473 2427 1474
rect 2431 1478 2435 1479
rect 2431 1473 2435 1474
rect 2551 1478 2555 1479
rect 2551 1473 2555 1474
rect 2591 1478 2595 1479
rect 2591 1473 2595 1474
rect 2679 1478 2683 1479
rect 2679 1473 2683 1474
rect 2735 1478 2739 1479
rect 2735 1473 2739 1474
rect 2799 1478 2803 1479
rect 2799 1473 2803 1474
rect 2871 1478 2875 1479
rect 2871 1473 2875 1474
rect 2927 1478 2931 1479
rect 2927 1473 2931 1474
rect 3007 1478 3011 1479
rect 3007 1473 3011 1474
rect 3055 1478 3059 1479
rect 3055 1473 3059 1474
rect 3135 1478 3139 1479
rect 3135 1473 3139 1474
rect 3263 1478 3267 1479
rect 3263 1473 3267 1474
rect 3367 1478 3371 1479
rect 3367 1473 3371 1474
rect 3463 1478 3467 1479
rect 3463 1473 3467 1474
rect 112 1454 114 1473
rect 160 1457 162 1473
rect 376 1457 378 1473
rect 584 1457 586 1473
rect 784 1457 786 1473
rect 960 1457 962 1473
rect 1128 1457 1130 1473
rect 1280 1457 1282 1473
rect 1432 1457 1434 1473
rect 1592 1457 1594 1473
rect 158 1456 164 1457
rect 110 1453 116 1454
rect 110 1449 111 1453
rect 115 1449 116 1453
rect 158 1452 159 1456
rect 163 1452 164 1456
rect 158 1451 164 1452
rect 374 1456 380 1457
rect 374 1452 375 1456
rect 379 1452 380 1456
rect 374 1451 380 1452
rect 582 1456 588 1457
rect 582 1452 583 1456
rect 587 1452 588 1456
rect 582 1451 588 1452
rect 782 1456 788 1457
rect 782 1452 783 1456
rect 787 1452 788 1456
rect 782 1451 788 1452
rect 958 1456 964 1457
rect 958 1452 959 1456
rect 963 1452 964 1456
rect 958 1451 964 1452
rect 1126 1456 1132 1457
rect 1126 1452 1127 1456
rect 1131 1452 1132 1456
rect 1126 1451 1132 1452
rect 1278 1456 1284 1457
rect 1278 1452 1279 1456
rect 1283 1452 1284 1456
rect 1278 1451 1284 1452
rect 1430 1456 1436 1457
rect 1430 1452 1431 1456
rect 1435 1452 1436 1456
rect 1430 1451 1436 1452
rect 1590 1456 1596 1457
rect 1590 1452 1591 1456
rect 1595 1452 1596 1456
rect 1768 1454 1770 1473
rect 1808 1454 1810 1473
rect 1832 1457 1834 1473
rect 1952 1457 1954 1473
rect 2112 1457 2114 1473
rect 2272 1457 2274 1473
rect 2432 1457 2434 1473
rect 2592 1457 2594 1473
rect 2736 1457 2738 1473
rect 2872 1457 2874 1473
rect 3008 1457 3010 1473
rect 3136 1457 3138 1473
rect 3264 1457 3266 1473
rect 3368 1457 3370 1473
rect 1830 1456 1836 1457
rect 1590 1451 1596 1452
rect 1766 1453 1772 1454
rect 110 1448 116 1449
rect 1766 1449 1767 1453
rect 1771 1449 1772 1453
rect 1766 1448 1772 1449
rect 1806 1453 1812 1454
rect 1806 1449 1807 1453
rect 1811 1449 1812 1453
rect 1830 1452 1831 1456
rect 1835 1452 1836 1456
rect 1830 1451 1836 1452
rect 1950 1456 1956 1457
rect 1950 1452 1951 1456
rect 1955 1452 1956 1456
rect 1950 1451 1956 1452
rect 2110 1456 2116 1457
rect 2110 1452 2111 1456
rect 2115 1452 2116 1456
rect 2110 1451 2116 1452
rect 2270 1456 2276 1457
rect 2270 1452 2271 1456
rect 2275 1452 2276 1456
rect 2270 1451 2276 1452
rect 2430 1456 2436 1457
rect 2430 1452 2431 1456
rect 2435 1452 2436 1456
rect 2430 1451 2436 1452
rect 2590 1456 2596 1457
rect 2590 1452 2591 1456
rect 2595 1452 2596 1456
rect 2590 1451 2596 1452
rect 2734 1456 2740 1457
rect 2734 1452 2735 1456
rect 2739 1452 2740 1456
rect 2734 1451 2740 1452
rect 2870 1456 2876 1457
rect 2870 1452 2871 1456
rect 2875 1452 2876 1456
rect 2870 1451 2876 1452
rect 3006 1456 3012 1457
rect 3006 1452 3007 1456
rect 3011 1452 3012 1456
rect 3006 1451 3012 1452
rect 3134 1456 3140 1457
rect 3134 1452 3135 1456
rect 3139 1452 3140 1456
rect 3134 1451 3140 1452
rect 3262 1456 3268 1457
rect 3262 1452 3263 1456
rect 3267 1452 3268 1456
rect 3262 1451 3268 1452
rect 3366 1456 3372 1457
rect 3366 1452 3367 1456
rect 3371 1452 3372 1456
rect 3464 1454 3466 1473
rect 3366 1451 3372 1452
rect 3462 1453 3468 1454
rect 1806 1448 1812 1449
rect 3462 1449 3463 1453
rect 3467 1449 3468 1453
rect 3462 1448 3468 1449
rect 158 1437 164 1438
rect 110 1436 116 1437
rect 110 1432 111 1436
rect 115 1432 116 1436
rect 158 1433 159 1437
rect 163 1433 164 1437
rect 158 1432 164 1433
rect 374 1437 380 1438
rect 374 1433 375 1437
rect 379 1433 380 1437
rect 374 1432 380 1433
rect 582 1437 588 1438
rect 582 1433 583 1437
rect 587 1433 588 1437
rect 582 1432 588 1433
rect 782 1437 788 1438
rect 782 1433 783 1437
rect 787 1433 788 1437
rect 782 1432 788 1433
rect 958 1437 964 1438
rect 958 1433 959 1437
rect 963 1433 964 1437
rect 958 1432 964 1433
rect 1126 1437 1132 1438
rect 1126 1433 1127 1437
rect 1131 1433 1132 1437
rect 1126 1432 1132 1433
rect 1278 1437 1284 1438
rect 1278 1433 1279 1437
rect 1283 1433 1284 1437
rect 1278 1432 1284 1433
rect 1430 1437 1436 1438
rect 1430 1433 1431 1437
rect 1435 1433 1436 1437
rect 1430 1432 1436 1433
rect 1590 1437 1596 1438
rect 1830 1437 1836 1438
rect 1590 1433 1591 1437
rect 1595 1433 1596 1437
rect 1590 1432 1596 1433
rect 1766 1436 1772 1437
rect 1766 1432 1767 1436
rect 1771 1432 1772 1436
rect 110 1431 116 1432
rect 112 1411 114 1431
rect 160 1411 162 1432
rect 376 1411 378 1432
rect 584 1411 586 1432
rect 784 1411 786 1432
rect 960 1411 962 1432
rect 1128 1411 1130 1432
rect 1280 1411 1282 1432
rect 1432 1411 1434 1432
rect 1592 1411 1594 1432
rect 1766 1431 1772 1432
rect 1806 1436 1812 1437
rect 1806 1432 1807 1436
rect 1811 1432 1812 1436
rect 1830 1433 1831 1437
rect 1835 1433 1836 1437
rect 1830 1432 1836 1433
rect 1950 1437 1956 1438
rect 1950 1433 1951 1437
rect 1955 1433 1956 1437
rect 1950 1432 1956 1433
rect 2110 1437 2116 1438
rect 2110 1433 2111 1437
rect 2115 1433 2116 1437
rect 2110 1432 2116 1433
rect 2270 1437 2276 1438
rect 2270 1433 2271 1437
rect 2275 1433 2276 1437
rect 2270 1432 2276 1433
rect 2430 1437 2436 1438
rect 2430 1433 2431 1437
rect 2435 1433 2436 1437
rect 2430 1432 2436 1433
rect 2590 1437 2596 1438
rect 2590 1433 2591 1437
rect 2595 1433 2596 1437
rect 2590 1432 2596 1433
rect 2734 1437 2740 1438
rect 2734 1433 2735 1437
rect 2739 1433 2740 1437
rect 2734 1432 2740 1433
rect 2870 1437 2876 1438
rect 2870 1433 2871 1437
rect 2875 1433 2876 1437
rect 2870 1432 2876 1433
rect 3006 1437 3012 1438
rect 3006 1433 3007 1437
rect 3011 1433 3012 1437
rect 3006 1432 3012 1433
rect 3134 1437 3140 1438
rect 3134 1433 3135 1437
rect 3139 1433 3140 1437
rect 3134 1432 3140 1433
rect 3262 1437 3268 1438
rect 3262 1433 3263 1437
rect 3267 1433 3268 1437
rect 3262 1432 3268 1433
rect 3366 1437 3372 1438
rect 3366 1433 3367 1437
rect 3371 1433 3372 1437
rect 3366 1432 3372 1433
rect 3462 1436 3468 1437
rect 3462 1432 3463 1436
rect 3467 1432 3468 1436
rect 1806 1431 1812 1432
rect 1768 1411 1770 1431
rect 1808 1411 1810 1431
rect 1832 1411 1834 1432
rect 1952 1411 1954 1432
rect 2112 1411 2114 1432
rect 2272 1411 2274 1432
rect 2432 1411 2434 1432
rect 2592 1411 2594 1432
rect 2736 1411 2738 1432
rect 2872 1411 2874 1432
rect 3008 1411 3010 1432
rect 3136 1411 3138 1432
rect 3264 1411 3266 1432
rect 3368 1411 3370 1432
rect 3462 1431 3468 1432
rect 3464 1411 3466 1431
rect 111 1410 115 1411
rect 111 1405 115 1406
rect 135 1410 139 1411
rect 135 1405 139 1406
rect 159 1410 163 1411
rect 159 1405 163 1406
rect 303 1410 307 1411
rect 303 1405 307 1406
rect 375 1410 379 1411
rect 375 1405 379 1406
rect 495 1410 499 1411
rect 495 1405 499 1406
rect 583 1410 587 1411
rect 583 1405 587 1406
rect 679 1410 683 1411
rect 679 1405 683 1406
rect 783 1410 787 1411
rect 783 1405 787 1406
rect 855 1410 859 1411
rect 855 1405 859 1406
rect 959 1410 963 1411
rect 959 1405 963 1406
rect 1015 1410 1019 1411
rect 1015 1405 1019 1406
rect 1127 1410 1131 1411
rect 1127 1405 1131 1406
rect 1167 1410 1171 1411
rect 1167 1405 1171 1406
rect 1279 1410 1283 1411
rect 1279 1405 1283 1406
rect 1303 1410 1307 1411
rect 1303 1405 1307 1406
rect 1431 1410 1435 1411
rect 1431 1405 1435 1406
rect 1559 1410 1563 1411
rect 1559 1405 1563 1406
rect 1591 1410 1595 1411
rect 1591 1405 1595 1406
rect 1671 1410 1675 1411
rect 1671 1405 1675 1406
rect 1767 1410 1771 1411
rect 1767 1405 1771 1406
rect 1807 1410 1811 1411
rect 1807 1405 1811 1406
rect 1831 1410 1835 1411
rect 1831 1405 1835 1406
rect 1951 1410 1955 1411
rect 1951 1405 1955 1406
rect 2007 1410 2011 1411
rect 2007 1405 2011 1406
rect 2111 1410 2115 1411
rect 2111 1405 2115 1406
rect 2199 1410 2203 1411
rect 2199 1405 2203 1406
rect 2271 1410 2275 1411
rect 2271 1405 2275 1406
rect 2383 1410 2387 1411
rect 2383 1405 2387 1406
rect 2431 1410 2435 1411
rect 2431 1405 2435 1406
rect 2559 1410 2563 1411
rect 2559 1405 2563 1406
rect 2591 1410 2595 1411
rect 2591 1405 2595 1406
rect 2719 1410 2723 1411
rect 2719 1405 2723 1406
rect 2735 1410 2739 1411
rect 2735 1405 2739 1406
rect 2863 1410 2867 1411
rect 2863 1405 2867 1406
rect 2871 1410 2875 1411
rect 2871 1405 2875 1406
rect 2999 1410 3003 1411
rect 2999 1405 3003 1406
rect 3007 1410 3011 1411
rect 3007 1405 3011 1406
rect 3127 1410 3131 1411
rect 3127 1405 3131 1406
rect 3135 1410 3139 1411
rect 3135 1405 3139 1406
rect 3255 1410 3259 1411
rect 3255 1405 3259 1406
rect 3263 1410 3267 1411
rect 3263 1405 3267 1406
rect 3367 1410 3371 1411
rect 3367 1405 3371 1406
rect 3463 1410 3467 1411
rect 3463 1405 3467 1406
rect 112 1389 114 1405
rect 110 1388 116 1389
rect 136 1388 138 1405
rect 304 1388 306 1405
rect 496 1388 498 1405
rect 680 1388 682 1405
rect 856 1388 858 1405
rect 1016 1388 1018 1405
rect 1168 1388 1170 1405
rect 1304 1388 1306 1405
rect 1432 1388 1434 1405
rect 1560 1388 1562 1405
rect 1672 1388 1674 1405
rect 1768 1389 1770 1405
rect 1808 1389 1810 1405
rect 1766 1388 1772 1389
rect 110 1384 111 1388
rect 115 1384 116 1388
rect 110 1383 116 1384
rect 134 1387 140 1388
rect 134 1383 135 1387
rect 139 1383 140 1387
rect 134 1382 140 1383
rect 302 1387 308 1388
rect 302 1383 303 1387
rect 307 1383 308 1387
rect 302 1382 308 1383
rect 494 1387 500 1388
rect 494 1383 495 1387
rect 499 1383 500 1387
rect 494 1382 500 1383
rect 678 1387 684 1388
rect 678 1383 679 1387
rect 683 1383 684 1387
rect 678 1382 684 1383
rect 854 1387 860 1388
rect 854 1383 855 1387
rect 859 1383 860 1387
rect 854 1382 860 1383
rect 1014 1387 1020 1388
rect 1014 1383 1015 1387
rect 1019 1383 1020 1387
rect 1014 1382 1020 1383
rect 1166 1387 1172 1388
rect 1166 1383 1167 1387
rect 1171 1383 1172 1387
rect 1166 1382 1172 1383
rect 1302 1387 1308 1388
rect 1302 1383 1303 1387
rect 1307 1383 1308 1387
rect 1302 1382 1308 1383
rect 1430 1387 1436 1388
rect 1430 1383 1431 1387
rect 1435 1383 1436 1387
rect 1430 1382 1436 1383
rect 1558 1387 1564 1388
rect 1558 1383 1559 1387
rect 1563 1383 1564 1387
rect 1558 1382 1564 1383
rect 1670 1387 1676 1388
rect 1670 1383 1671 1387
rect 1675 1383 1676 1387
rect 1766 1384 1767 1388
rect 1771 1384 1772 1388
rect 1766 1383 1772 1384
rect 1806 1388 1812 1389
rect 1832 1388 1834 1405
rect 2008 1388 2010 1405
rect 2200 1388 2202 1405
rect 2384 1388 2386 1405
rect 2560 1388 2562 1405
rect 2720 1388 2722 1405
rect 2864 1388 2866 1405
rect 3000 1388 3002 1405
rect 3128 1388 3130 1405
rect 3256 1388 3258 1405
rect 3368 1388 3370 1405
rect 3464 1389 3466 1405
rect 3462 1388 3468 1389
rect 1806 1384 1807 1388
rect 1811 1384 1812 1388
rect 1806 1383 1812 1384
rect 1830 1387 1836 1388
rect 1830 1383 1831 1387
rect 1835 1383 1836 1387
rect 1670 1382 1676 1383
rect 1830 1382 1836 1383
rect 2006 1387 2012 1388
rect 2006 1383 2007 1387
rect 2011 1383 2012 1387
rect 2006 1382 2012 1383
rect 2198 1387 2204 1388
rect 2198 1383 2199 1387
rect 2203 1383 2204 1387
rect 2198 1382 2204 1383
rect 2382 1387 2388 1388
rect 2382 1383 2383 1387
rect 2387 1383 2388 1387
rect 2382 1382 2388 1383
rect 2558 1387 2564 1388
rect 2558 1383 2559 1387
rect 2563 1383 2564 1387
rect 2558 1382 2564 1383
rect 2718 1387 2724 1388
rect 2718 1383 2719 1387
rect 2723 1383 2724 1387
rect 2718 1382 2724 1383
rect 2862 1387 2868 1388
rect 2862 1383 2863 1387
rect 2867 1383 2868 1387
rect 2862 1382 2868 1383
rect 2998 1387 3004 1388
rect 2998 1383 2999 1387
rect 3003 1383 3004 1387
rect 2998 1382 3004 1383
rect 3126 1387 3132 1388
rect 3126 1383 3127 1387
rect 3131 1383 3132 1387
rect 3126 1382 3132 1383
rect 3254 1387 3260 1388
rect 3254 1383 3255 1387
rect 3259 1383 3260 1387
rect 3254 1382 3260 1383
rect 3366 1387 3372 1388
rect 3366 1383 3367 1387
rect 3371 1383 3372 1387
rect 3462 1384 3463 1388
rect 3467 1384 3468 1388
rect 3462 1383 3468 1384
rect 3366 1382 3372 1383
rect 110 1371 116 1372
rect 110 1367 111 1371
rect 115 1367 116 1371
rect 1766 1371 1772 1372
rect 110 1366 116 1367
rect 134 1368 140 1369
rect 112 1343 114 1366
rect 134 1364 135 1368
rect 139 1364 140 1368
rect 134 1363 140 1364
rect 302 1368 308 1369
rect 302 1364 303 1368
rect 307 1364 308 1368
rect 302 1363 308 1364
rect 494 1368 500 1369
rect 494 1364 495 1368
rect 499 1364 500 1368
rect 494 1363 500 1364
rect 678 1368 684 1369
rect 678 1364 679 1368
rect 683 1364 684 1368
rect 678 1363 684 1364
rect 854 1368 860 1369
rect 854 1364 855 1368
rect 859 1364 860 1368
rect 854 1363 860 1364
rect 1014 1368 1020 1369
rect 1014 1364 1015 1368
rect 1019 1364 1020 1368
rect 1014 1363 1020 1364
rect 1166 1368 1172 1369
rect 1166 1364 1167 1368
rect 1171 1364 1172 1368
rect 1166 1363 1172 1364
rect 1302 1368 1308 1369
rect 1302 1364 1303 1368
rect 1307 1364 1308 1368
rect 1302 1363 1308 1364
rect 1430 1368 1436 1369
rect 1430 1364 1431 1368
rect 1435 1364 1436 1368
rect 1430 1363 1436 1364
rect 1558 1368 1564 1369
rect 1558 1364 1559 1368
rect 1563 1364 1564 1368
rect 1558 1363 1564 1364
rect 1670 1368 1676 1369
rect 1670 1364 1671 1368
rect 1675 1364 1676 1368
rect 1766 1367 1767 1371
rect 1771 1367 1772 1371
rect 1766 1366 1772 1367
rect 1806 1371 1812 1372
rect 1806 1367 1807 1371
rect 1811 1367 1812 1371
rect 3462 1371 3468 1372
rect 1806 1366 1812 1367
rect 1830 1368 1836 1369
rect 1670 1363 1676 1364
rect 136 1343 138 1363
rect 304 1343 306 1363
rect 496 1343 498 1363
rect 680 1343 682 1363
rect 856 1343 858 1363
rect 1016 1343 1018 1363
rect 1168 1343 1170 1363
rect 1304 1343 1306 1363
rect 1432 1343 1434 1363
rect 1560 1343 1562 1363
rect 1672 1343 1674 1363
rect 1768 1343 1770 1366
rect 111 1342 115 1343
rect 111 1337 115 1338
rect 135 1342 139 1343
rect 135 1337 139 1338
rect 247 1342 251 1343
rect 247 1337 251 1338
rect 303 1342 307 1343
rect 303 1337 307 1338
rect 399 1342 403 1343
rect 399 1337 403 1338
rect 495 1342 499 1343
rect 495 1337 499 1338
rect 559 1342 563 1343
rect 559 1337 563 1338
rect 679 1342 683 1343
rect 679 1337 683 1338
rect 727 1342 731 1343
rect 727 1337 731 1338
rect 855 1342 859 1343
rect 855 1337 859 1338
rect 895 1342 899 1343
rect 895 1337 899 1338
rect 1015 1342 1019 1343
rect 1015 1337 1019 1338
rect 1063 1342 1067 1343
rect 1063 1337 1067 1338
rect 1167 1342 1171 1343
rect 1167 1337 1171 1338
rect 1223 1342 1227 1343
rect 1223 1337 1227 1338
rect 1303 1342 1307 1343
rect 1303 1337 1307 1338
rect 1375 1342 1379 1343
rect 1375 1337 1379 1338
rect 1431 1342 1435 1343
rect 1431 1337 1435 1338
rect 1535 1342 1539 1343
rect 1535 1337 1539 1338
rect 1559 1342 1563 1343
rect 1559 1337 1563 1338
rect 1671 1342 1675 1343
rect 1671 1337 1675 1338
rect 1767 1342 1771 1343
rect 1808 1339 1810 1366
rect 1830 1364 1831 1368
rect 1835 1364 1836 1368
rect 1830 1363 1836 1364
rect 2006 1368 2012 1369
rect 2006 1364 2007 1368
rect 2011 1364 2012 1368
rect 2006 1363 2012 1364
rect 2198 1368 2204 1369
rect 2198 1364 2199 1368
rect 2203 1364 2204 1368
rect 2198 1363 2204 1364
rect 2382 1368 2388 1369
rect 2382 1364 2383 1368
rect 2387 1364 2388 1368
rect 2382 1363 2388 1364
rect 2558 1368 2564 1369
rect 2558 1364 2559 1368
rect 2563 1364 2564 1368
rect 2558 1363 2564 1364
rect 2718 1368 2724 1369
rect 2718 1364 2719 1368
rect 2723 1364 2724 1368
rect 2718 1363 2724 1364
rect 2862 1368 2868 1369
rect 2862 1364 2863 1368
rect 2867 1364 2868 1368
rect 2862 1363 2868 1364
rect 2998 1368 3004 1369
rect 2998 1364 2999 1368
rect 3003 1364 3004 1368
rect 2998 1363 3004 1364
rect 3126 1368 3132 1369
rect 3126 1364 3127 1368
rect 3131 1364 3132 1368
rect 3126 1363 3132 1364
rect 3254 1368 3260 1369
rect 3254 1364 3255 1368
rect 3259 1364 3260 1368
rect 3254 1363 3260 1364
rect 3366 1368 3372 1369
rect 3366 1364 3367 1368
rect 3371 1364 3372 1368
rect 3462 1367 3463 1371
rect 3467 1367 3468 1371
rect 3462 1366 3468 1367
rect 3366 1363 3372 1364
rect 1832 1339 1834 1363
rect 2008 1339 2010 1363
rect 2200 1339 2202 1363
rect 2384 1339 2386 1363
rect 2560 1339 2562 1363
rect 2720 1339 2722 1363
rect 2864 1339 2866 1363
rect 3000 1339 3002 1363
rect 3128 1339 3130 1363
rect 3256 1339 3258 1363
rect 3368 1339 3370 1363
rect 3464 1339 3466 1366
rect 1767 1337 1771 1338
rect 1807 1338 1811 1339
rect 112 1318 114 1337
rect 136 1321 138 1337
rect 248 1321 250 1337
rect 400 1321 402 1337
rect 560 1321 562 1337
rect 728 1321 730 1337
rect 896 1321 898 1337
rect 1064 1321 1066 1337
rect 1224 1321 1226 1337
rect 1376 1321 1378 1337
rect 1536 1321 1538 1337
rect 1672 1321 1674 1337
rect 134 1320 140 1321
rect 110 1317 116 1318
rect 110 1313 111 1317
rect 115 1313 116 1317
rect 134 1316 135 1320
rect 139 1316 140 1320
rect 134 1315 140 1316
rect 246 1320 252 1321
rect 246 1316 247 1320
rect 251 1316 252 1320
rect 246 1315 252 1316
rect 398 1320 404 1321
rect 398 1316 399 1320
rect 403 1316 404 1320
rect 398 1315 404 1316
rect 558 1320 564 1321
rect 558 1316 559 1320
rect 563 1316 564 1320
rect 558 1315 564 1316
rect 726 1320 732 1321
rect 726 1316 727 1320
rect 731 1316 732 1320
rect 726 1315 732 1316
rect 894 1320 900 1321
rect 894 1316 895 1320
rect 899 1316 900 1320
rect 894 1315 900 1316
rect 1062 1320 1068 1321
rect 1062 1316 1063 1320
rect 1067 1316 1068 1320
rect 1062 1315 1068 1316
rect 1222 1320 1228 1321
rect 1222 1316 1223 1320
rect 1227 1316 1228 1320
rect 1222 1315 1228 1316
rect 1374 1320 1380 1321
rect 1374 1316 1375 1320
rect 1379 1316 1380 1320
rect 1374 1315 1380 1316
rect 1534 1320 1540 1321
rect 1534 1316 1535 1320
rect 1539 1316 1540 1320
rect 1534 1315 1540 1316
rect 1670 1320 1676 1321
rect 1670 1316 1671 1320
rect 1675 1316 1676 1320
rect 1768 1318 1770 1337
rect 1807 1333 1811 1334
rect 1831 1338 1835 1339
rect 1831 1333 1835 1334
rect 1967 1338 1971 1339
rect 1967 1333 1971 1334
rect 2007 1338 2011 1339
rect 2007 1333 2011 1334
rect 2143 1338 2147 1339
rect 2143 1333 2147 1334
rect 2199 1338 2203 1339
rect 2199 1333 2203 1334
rect 2327 1338 2331 1339
rect 2327 1333 2331 1334
rect 2383 1338 2387 1339
rect 2383 1333 2387 1334
rect 2511 1338 2515 1339
rect 2511 1333 2515 1334
rect 2559 1338 2563 1339
rect 2559 1333 2563 1334
rect 2687 1338 2691 1339
rect 2687 1333 2691 1334
rect 2719 1338 2723 1339
rect 2719 1333 2723 1334
rect 2863 1338 2867 1339
rect 2863 1333 2867 1334
rect 2999 1338 3003 1339
rect 2999 1333 3003 1334
rect 3039 1338 3043 1339
rect 3039 1333 3043 1334
rect 3127 1338 3131 1339
rect 3127 1333 3131 1334
rect 3215 1338 3219 1339
rect 3215 1333 3219 1334
rect 3255 1338 3259 1339
rect 3255 1333 3259 1334
rect 3367 1338 3371 1339
rect 3367 1333 3371 1334
rect 3463 1338 3467 1339
rect 3463 1333 3467 1334
rect 1670 1315 1676 1316
rect 1766 1317 1772 1318
rect 110 1312 116 1313
rect 1766 1313 1767 1317
rect 1771 1313 1772 1317
rect 1808 1314 1810 1333
rect 1832 1317 1834 1333
rect 1968 1317 1970 1333
rect 2144 1317 2146 1333
rect 2328 1317 2330 1333
rect 2512 1317 2514 1333
rect 2688 1317 2690 1333
rect 2864 1317 2866 1333
rect 3040 1317 3042 1333
rect 3216 1317 3218 1333
rect 3368 1317 3370 1333
rect 1830 1316 1836 1317
rect 1766 1312 1772 1313
rect 1806 1313 1812 1314
rect 1806 1309 1807 1313
rect 1811 1309 1812 1313
rect 1830 1312 1831 1316
rect 1835 1312 1836 1316
rect 1830 1311 1836 1312
rect 1966 1316 1972 1317
rect 1966 1312 1967 1316
rect 1971 1312 1972 1316
rect 1966 1311 1972 1312
rect 2142 1316 2148 1317
rect 2142 1312 2143 1316
rect 2147 1312 2148 1316
rect 2142 1311 2148 1312
rect 2326 1316 2332 1317
rect 2326 1312 2327 1316
rect 2331 1312 2332 1316
rect 2326 1311 2332 1312
rect 2510 1316 2516 1317
rect 2510 1312 2511 1316
rect 2515 1312 2516 1316
rect 2510 1311 2516 1312
rect 2686 1316 2692 1317
rect 2686 1312 2687 1316
rect 2691 1312 2692 1316
rect 2686 1311 2692 1312
rect 2862 1316 2868 1317
rect 2862 1312 2863 1316
rect 2867 1312 2868 1316
rect 2862 1311 2868 1312
rect 3038 1316 3044 1317
rect 3038 1312 3039 1316
rect 3043 1312 3044 1316
rect 3038 1311 3044 1312
rect 3214 1316 3220 1317
rect 3214 1312 3215 1316
rect 3219 1312 3220 1316
rect 3214 1311 3220 1312
rect 3366 1316 3372 1317
rect 3366 1312 3367 1316
rect 3371 1312 3372 1316
rect 3464 1314 3466 1333
rect 3366 1311 3372 1312
rect 3462 1313 3468 1314
rect 1806 1308 1812 1309
rect 3462 1309 3463 1313
rect 3467 1309 3468 1313
rect 3462 1308 3468 1309
rect 134 1301 140 1302
rect 110 1300 116 1301
rect 110 1296 111 1300
rect 115 1296 116 1300
rect 134 1297 135 1301
rect 139 1297 140 1301
rect 134 1296 140 1297
rect 246 1301 252 1302
rect 246 1297 247 1301
rect 251 1297 252 1301
rect 246 1296 252 1297
rect 398 1301 404 1302
rect 398 1297 399 1301
rect 403 1297 404 1301
rect 398 1296 404 1297
rect 558 1301 564 1302
rect 558 1297 559 1301
rect 563 1297 564 1301
rect 558 1296 564 1297
rect 726 1301 732 1302
rect 726 1297 727 1301
rect 731 1297 732 1301
rect 726 1296 732 1297
rect 894 1301 900 1302
rect 894 1297 895 1301
rect 899 1297 900 1301
rect 894 1296 900 1297
rect 1062 1301 1068 1302
rect 1062 1297 1063 1301
rect 1067 1297 1068 1301
rect 1062 1296 1068 1297
rect 1222 1301 1228 1302
rect 1222 1297 1223 1301
rect 1227 1297 1228 1301
rect 1222 1296 1228 1297
rect 1374 1301 1380 1302
rect 1374 1297 1375 1301
rect 1379 1297 1380 1301
rect 1374 1296 1380 1297
rect 1534 1301 1540 1302
rect 1534 1297 1535 1301
rect 1539 1297 1540 1301
rect 1534 1296 1540 1297
rect 1670 1301 1676 1302
rect 1670 1297 1671 1301
rect 1675 1297 1676 1301
rect 1670 1296 1676 1297
rect 1766 1300 1772 1301
rect 1766 1296 1767 1300
rect 1771 1296 1772 1300
rect 1830 1297 1836 1298
rect 110 1295 116 1296
rect 112 1275 114 1295
rect 136 1275 138 1296
rect 248 1275 250 1296
rect 400 1275 402 1296
rect 560 1275 562 1296
rect 728 1275 730 1296
rect 896 1275 898 1296
rect 1064 1275 1066 1296
rect 1224 1275 1226 1296
rect 1376 1275 1378 1296
rect 1536 1275 1538 1296
rect 1672 1275 1674 1296
rect 1766 1295 1772 1296
rect 1806 1296 1812 1297
rect 1768 1275 1770 1295
rect 1806 1292 1807 1296
rect 1811 1292 1812 1296
rect 1830 1293 1831 1297
rect 1835 1293 1836 1297
rect 1830 1292 1836 1293
rect 1966 1297 1972 1298
rect 1966 1293 1967 1297
rect 1971 1293 1972 1297
rect 1966 1292 1972 1293
rect 2142 1297 2148 1298
rect 2142 1293 2143 1297
rect 2147 1293 2148 1297
rect 2142 1292 2148 1293
rect 2326 1297 2332 1298
rect 2326 1293 2327 1297
rect 2331 1293 2332 1297
rect 2326 1292 2332 1293
rect 2510 1297 2516 1298
rect 2510 1293 2511 1297
rect 2515 1293 2516 1297
rect 2510 1292 2516 1293
rect 2686 1297 2692 1298
rect 2686 1293 2687 1297
rect 2691 1293 2692 1297
rect 2686 1292 2692 1293
rect 2862 1297 2868 1298
rect 2862 1293 2863 1297
rect 2867 1293 2868 1297
rect 2862 1292 2868 1293
rect 3038 1297 3044 1298
rect 3038 1293 3039 1297
rect 3043 1293 3044 1297
rect 3038 1292 3044 1293
rect 3214 1297 3220 1298
rect 3214 1293 3215 1297
rect 3219 1293 3220 1297
rect 3214 1292 3220 1293
rect 3366 1297 3372 1298
rect 3366 1293 3367 1297
rect 3371 1293 3372 1297
rect 3366 1292 3372 1293
rect 3462 1296 3468 1297
rect 3462 1292 3463 1296
rect 3467 1292 3468 1296
rect 1806 1291 1812 1292
rect 1808 1275 1810 1291
rect 1832 1275 1834 1292
rect 1968 1275 1970 1292
rect 2144 1275 2146 1292
rect 2328 1275 2330 1292
rect 2512 1275 2514 1292
rect 2688 1275 2690 1292
rect 2864 1275 2866 1292
rect 3040 1275 3042 1292
rect 3216 1275 3218 1292
rect 3368 1275 3370 1292
rect 3462 1291 3468 1292
rect 3464 1275 3466 1291
rect 111 1274 115 1275
rect 111 1269 115 1270
rect 135 1274 139 1275
rect 135 1269 139 1270
rect 223 1274 227 1275
rect 223 1269 227 1270
rect 247 1274 251 1275
rect 247 1269 251 1270
rect 319 1274 323 1275
rect 319 1269 323 1270
rect 399 1274 403 1275
rect 399 1269 403 1270
rect 431 1274 435 1275
rect 431 1269 435 1270
rect 551 1274 555 1275
rect 551 1269 555 1270
rect 559 1274 563 1275
rect 559 1269 563 1270
rect 679 1274 683 1275
rect 679 1269 683 1270
rect 727 1274 731 1275
rect 727 1269 731 1270
rect 823 1274 827 1275
rect 823 1269 827 1270
rect 895 1274 899 1275
rect 895 1269 899 1270
rect 975 1274 979 1275
rect 975 1269 979 1270
rect 1063 1274 1067 1275
rect 1063 1269 1067 1270
rect 1143 1274 1147 1275
rect 1143 1269 1147 1270
rect 1223 1274 1227 1275
rect 1223 1269 1227 1270
rect 1319 1274 1323 1275
rect 1319 1269 1323 1270
rect 1375 1274 1379 1275
rect 1375 1269 1379 1270
rect 1503 1274 1507 1275
rect 1503 1269 1507 1270
rect 1535 1274 1539 1275
rect 1535 1269 1539 1270
rect 1671 1274 1675 1275
rect 1671 1269 1675 1270
rect 1767 1274 1771 1275
rect 1767 1269 1771 1270
rect 1807 1274 1811 1275
rect 1807 1269 1811 1270
rect 1831 1274 1835 1275
rect 1831 1269 1835 1270
rect 1967 1274 1971 1275
rect 1967 1269 1971 1270
rect 2095 1274 2099 1275
rect 2095 1269 2099 1270
rect 2143 1274 2147 1275
rect 2143 1269 2147 1270
rect 2327 1274 2331 1275
rect 2327 1269 2331 1270
rect 2359 1274 2363 1275
rect 2359 1269 2363 1270
rect 2511 1274 2515 1275
rect 2511 1269 2515 1270
rect 2599 1274 2603 1275
rect 2599 1269 2603 1270
rect 2687 1274 2691 1275
rect 2687 1269 2691 1270
rect 2807 1274 2811 1275
rect 2807 1269 2811 1270
rect 2863 1274 2867 1275
rect 2863 1269 2867 1270
rect 3007 1274 3011 1275
rect 3007 1269 3011 1270
rect 3039 1274 3043 1275
rect 3039 1269 3043 1270
rect 3199 1274 3203 1275
rect 3199 1269 3203 1270
rect 3215 1274 3219 1275
rect 3215 1269 3219 1270
rect 3367 1274 3371 1275
rect 3367 1269 3371 1270
rect 3463 1274 3467 1275
rect 3463 1269 3467 1270
rect 112 1253 114 1269
rect 110 1252 116 1253
rect 136 1252 138 1269
rect 224 1252 226 1269
rect 320 1252 322 1269
rect 432 1252 434 1269
rect 552 1252 554 1269
rect 680 1252 682 1269
rect 824 1252 826 1269
rect 976 1252 978 1269
rect 1144 1252 1146 1269
rect 1320 1252 1322 1269
rect 1504 1252 1506 1269
rect 1672 1252 1674 1269
rect 1768 1253 1770 1269
rect 1808 1253 1810 1269
rect 1766 1252 1772 1253
rect 110 1248 111 1252
rect 115 1248 116 1252
rect 110 1247 116 1248
rect 134 1251 140 1252
rect 134 1247 135 1251
rect 139 1247 140 1251
rect 134 1246 140 1247
rect 222 1251 228 1252
rect 222 1247 223 1251
rect 227 1247 228 1251
rect 222 1246 228 1247
rect 318 1251 324 1252
rect 318 1247 319 1251
rect 323 1247 324 1251
rect 318 1246 324 1247
rect 430 1251 436 1252
rect 430 1247 431 1251
rect 435 1247 436 1251
rect 430 1246 436 1247
rect 550 1251 556 1252
rect 550 1247 551 1251
rect 555 1247 556 1251
rect 550 1246 556 1247
rect 678 1251 684 1252
rect 678 1247 679 1251
rect 683 1247 684 1251
rect 678 1246 684 1247
rect 822 1251 828 1252
rect 822 1247 823 1251
rect 827 1247 828 1251
rect 822 1246 828 1247
rect 974 1251 980 1252
rect 974 1247 975 1251
rect 979 1247 980 1251
rect 974 1246 980 1247
rect 1142 1251 1148 1252
rect 1142 1247 1143 1251
rect 1147 1247 1148 1251
rect 1142 1246 1148 1247
rect 1318 1251 1324 1252
rect 1318 1247 1319 1251
rect 1323 1247 1324 1251
rect 1318 1246 1324 1247
rect 1502 1251 1508 1252
rect 1502 1247 1503 1251
rect 1507 1247 1508 1251
rect 1502 1246 1508 1247
rect 1670 1251 1676 1252
rect 1670 1247 1671 1251
rect 1675 1247 1676 1251
rect 1766 1248 1767 1252
rect 1771 1248 1772 1252
rect 1766 1247 1772 1248
rect 1806 1252 1812 1253
rect 1832 1252 1834 1269
rect 2096 1252 2098 1269
rect 2360 1252 2362 1269
rect 2600 1252 2602 1269
rect 2808 1252 2810 1269
rect 3008 1252 3010 1269
rect 3200 1252 3202 1269
rect 3368 1252 3370 1269
rect 3464 1253 3466 1269
rect 3462 1252 3468 1253
rect 1806 1248 1807 1252
rect 1811 1248 1812 1252
rect 1806 1247 1812 1248
rect 1830 1251 1836 1252
rect 1830 1247 1831 1251
rect 1835 1247 1836 1251
rect 1670 1246 1676 1247
rect 1830 1246 1836 1247
rect 2094 1251 2100 1252
rect 2094 1247 2095 1251
rect 2099 1247 2100 1251
rect 2094 1246 2100 1247
rect 2358 1251 2364 1252
rect 2358 1247 2359 1251
rect 2363 1247 2364 1251
rect 2358 1246 2364 1247
rect 2598 1251 2604 1252
rect 2598 1247 2599 1251
rect 2603 1247 2604 1251
rect 2598 1246 2604 1247
rect 2806 1251 2812 1252
rect 2806 1247 2807 1251
rect 2811 1247 2812 1251
rect 2806 1246 2812 1247
rect 3006 1251 3012 1252
rect 3006 1247 3007 1251
rect 3011 1247 3012 1251
rect 3006 1246 3012 1247
rect 3198 1251 3204 1252
rect 3198 1247 3199 1251
rect 3203 1247 3204 1251
rect 3198 1246 3204 1247
rect 3366 1251 3372 1252
rect 3366 1247 3367 1251
rect 3371 1247 3372 1251
rect 3462 1248 3463 1252
rect 3467 1248 3468 1252
rect 3462 1247 3468 1248
rect 3366 1246 3372 1247
rect 110 1235 116 1236
rect 110 1231 111 1235
rect 115 1231 116 1235
rect 1766 1235 1772 1236
rect 110 1230 116 1231
rect 134 1232 140 1233
rect 112 1203 114 1230
rect 134 1228 135 1232
rect 139 1228 140 1232
rect 134 1227 140 1228
rect 222 1232 228 1233
rect 222 1228 223 1232
rect 227 1228 228 1232
rect 222 1227 228 1228
rect 318 1232 324 1233
rect 318 1228 319 1232
rect 323 1228 324 1232
rect 318 1227 324 1228
rect 430 1232 436 1233
rect 430 1228 431 1232
rect 435 1228 436 1232
rect 430 1227 436 1228
rect 550 1232 556 1233
rect 550 1228 551 1232
rect 555 1228 556 1232
rect 550 1227 556 1228
rect 678 1232 684 1233
rect 678 1228 679 1232
rect 683 1228 684 1232
rect 678 1227 684 1228
rect 822 1232 828 1233
rect 822 1228 823 1232
rect 827 1228 828 1232
rect 822 1227 828 1228
rect 974 1232 980 1233
rect 974 1228 975 1232
rect 979 1228 980 1232
rect 974 1227 980 1228
rect 1142 1232 1148 1233
rect 1142 1228 1143 1232
rect 1147 1228 1148 1232
rect 1142 1227 1148 1228
rect 1318 1232 1324 1233
rect 1318 1228 1319 1232
rect 1323 1228 1324 1232
rect 1318 1227 1324 1228
rect 1502 1232 1508 1233
rect 1502 1228 1503 1232
rect 1507 1228 1508 1232
rect 1502 1227 1508 1228
rect 1670 1232 1676 1233
rect 1670 1228 1671 1232
rect 1675 1228 1676 1232
rect 1766 1231 1767 1235
rect 1771 1231 1772 1235
rect 1766 1230 1772 1231
rect 1806 1235 1812 1236
rect 1806 1231 1807 1235
rect 1811 1231 1812 1235
rect 3462 1235 3468 1236
rect 1806 1230 1812 1231
rect 1830 1232 1836 1233
rect 1670 1227 1676 1228
rect 136 1203 138 1227
rect 224 1203 226 1227
rect 320 1203 322 1227
rect 432 1203 434 1227
rect 552 1203 554 1227
rect 680 1203 682 1227
rect 824 1203 826 1227
rect 976 1203 978 1227
rect 1144 1203 1146 1227
rect 1320 1203 1322 1227
rect 1504 1203 1506 1227
rect 1672 1203 1674 1227
rect 1768 1203 1770 1230
rect 1808 1203 1810 1230
rect 1830 1228 1831 1232
rect 1835 1228 1836 1232
rect 1830 1227 1836 1228
rect 2094 1232 2100 1233
rect 2094 1228 2095 1232
rect 2099 1228 2100 1232
rect 2094 1227 2100 1228
rect 2358 1232 2364 1233
rect 2358 1228 2359 1232
rect 2363 1228 2364 1232
rect 2358 1227 2364 1228
rect 2598 1232 2604 1233
rect 2598 1228 2599 1232
rect 2603 1228 2604 1232
rect 2598 1227 2604 1228
rect 2806 1232 2812 1233
rect 2806 1228 2807 1232
rect 2811 1228 2812 1232
rect 2806 1227 2812 1228
rect 3006 1232 3012 1233
rect 3006 1228 3007 1232
rect 3011 1228 3012 1232
rect 3006 1227 3012 1228
rect 3198 1232 3204 1233
rect 3198 1228 3199 1232
rect 3203 1228 3204 1232
rect 3198 1227 3204 1228
rect 3366 1232 3372 1233
rect 3366 1228 3367 1232
rect 3371 1228 3372 1232
rect 3462 1231 3463 1235
rect 3467 1231 3468 1235
rect 3462 1230 3468 1231
rect 3366 1227 3372 1228
rect 1832 1203 1834 1227
rect 2096 1203 2098 1227
rect 2360 1203 2362 1227
rect 2600 1203 2602 1227
rect 2808 1203 2810 1227
rect 3008 1203 3010 1227
rect 3200 1203 3202 1227
rect 3368 1203 3370 1227
rect 3464 1203 3466 1230
rect 111 1202 115 1203
rect 111 1197 115 1198
rect 135 1202 139 1203
rect 135 1197 139 1198
rect 223 1202 227 1203
rect 223 1197 227 1198
rect 231 1202 235 1203
rect 231 1197 235 1198
rect 319 1202 323 1203
rect 319 1197 323 1198
rect 359 1202 363 1203
rect 359 1197 363 1198
rect 431 1202 435 1203
rect 431 1197 435 1198
rect 487 1202 491 1203
rect 487 1197 491 1198
rect 551 1202 555 1203
rect 551 1197 555 1198
rect 615 1202 619 1203
rect 615 1197 619 1198
rect 679 1202 683 1203
rect 679 1197 683 1198
rect 743 1202 747 1203
rect 743 1197 747 1198
rect 823 1202 827 1203
rect 823 1197 827 1198
rect 871 1202 875 1203
rect 871 1197 875 1198
rect 975 1202 979 1203
rect 975 1197 979 1198
rect 991 1202 995 1203
rect 991 1197 995 1198
rect 1119 1202 1123 1203
rect 1119 1197 1123 1198
rect 1143 1202 1147 1203
rect 1143 1197 1147 1198
rect 1247 1202 1251 1203
rect 1247 1197 1251 1198
rect 1319 1202 1323 1203
rect 1319 1197 1323 1198
rect 1503 1202 1507 1203
rect 1503 1197 1507 1198
rect 1671 1202 1675 1203
rect 1671 1197 1675 1198
rect 1767 1202 1771 1203
rect 1767 1197 1771 1198
rect 1807 1202 1811 1203
rect 1807 1197 1811 1198
rect 1831 1202 1835 1203
rect 1831 1197 1835 1198
rect 1935 1202 1939 1203
rect 1935 1197 1939 1198
rect 2039 1202 2043 1203
rect 2039 1197 2043 1198
rect 2095 1202 2099 1203
rect 2095 1197 2099 1198
rect 2159 1202 2163 1203
rect 2159 1197 2163 1198
rect 2287 1202 2291 1203
rect 2287 1197 2291 1198
rect 2359 1202 2363 1203
rect 2359 1197 2363 1198
rect 2423 1202 2427 1203
rect 2423 1197 2427 1198
rect 2567 1202 2571 1203
rect 2567 1197 2571 1198
rect 2599 1202 2603 1203
rect 2599 1197 2603 1198
rect 2703 1202 2707 1203
rect 2703 1197 2707 1198
rect 2807 1202 2811 1203
rect 2807 1197 2811 1198
rect 2839 1202 2843 1203
rect 2839 1197 2843 1198
rect 2975 1202 2979 1203
rect 2975 1197 2979 1198
rect 3007 1202 3011 1203
rect 3007 1197 3011 1198
rect 3111 1202 3115 1203
rect 3111 1197 3115 1198
rect 3199 1202 3203 1203
rect 3199 1197 3203 1198
rect 3247 1202 3251 1203
rect 3247 1197 3251 1198
rect 3367 1202 3371 1203
rect 3367 1197 3371 1198
rect 3463 1202 3467 1203
rect 3463 1197 3467 1198
rect 112 1178 114 1197
rect 136 1181 138 1197
rect 232 1181 234 1197
rect 360 1181 362 1197
rect 488 1181 490 1197
rect 616 1181 618 1197
rect 744 1181 746 1197
rect 872 1181 874 1197
rect 992 1181 994 1197
rect 1120 1181 1122 1197
rect 1248 1181 1250 1197
rect 134 1180 140 1181
rect 110 1177 116 1178
rect 110 1173 111 1177
rect 115 1173 116 1177
rect 134 1176 135 1180
rect 139 1176 140 1180
rect 134 1175 140 1176
rect 230 1180 236 1181
rect 230 1176 231 1180
rect 235 1176 236 1180
rect 230 1175 236 1176
rect 358 1180 364 1181
rect 358 1176 359 1180
rect 363 1176 364 1180
rect 358 1175 364 1176
rect 486 1180 492 1181
rect 486 1176 487 1180
rect 491 1176 492 1180
rect 486 1175 492 1176
rect 614 1180 620 1181
rect 614 1176 615 1180
rect 619 1176 620 1180
rect 614 1175 620 1176
rect 742 1180 748 1181
rect 742 1176 743 1180
rect 747 1176 748 1180
rect 742 1175 748 1176
rect 870 1180 876 1181
rect 870 1176 871 1180
rect 875 1176 876 1180
rect 870 1175 876 1176
rect 990 1180 996 1181
rect 990 1176 991 1180
rect 995 1176 996 1180
rect 990 1175 996 1176
rect 1118 1180 1124 1181
rect 1118 1176 1119 1180
rect 1123 1176 1124 1180
rect 1118 1175 1124 1176
rect 1246 1180 1252 1181
rect 1246 1176 1247 1180
rect 1251 1176 1252 1180
rect 1768 1178 1770 1197
rect 1808 1178 1810 1197
rect 1936 1181 1938 1197
rect 2040 1181 2042 1197
rect 2160 1181 2162 1197
rect 2288 1181 2290 1197
rect 2424 1181 2426 1197
rect 2568 1181 2570 1197
rect 2704 1181 2706 1197
rect 2840 1181 2842 1197
rect 2976 1181 2978 1197
rect 3112 1181 3114 1197
rect 3248 1181 3250 1197
rect 3368 1181 3370 1197
rect 1934 1180 1940 1181
rect 1246 1175 1252 1176
rect 1766 1177 1772 1178
rect 110 1172 116 1173
rect 1766 1173 1767 1177
rect 1771 1173 1772 1177
rect 1766 1172 1772 1173
rect 1806 1177 1812 1178
rect 1806 1173 1807 1177
rect 1811 1173 1812 1177
rect 1934 1176 1935 1180
rect 1939 1176 1940 1180
rect 1934 1175 1940 1176
rect 2038 1180 2044 1181
rect 2038 1176 2039 1180
rect 2043 1176 2044 1180
rect 2038 1175 2044 1176
rect 2158 1180 2164 1181
rect 2158 1176 2159 1180
rect 2163 1176 2164 1180
rect 2158 1175 2164 1176
rect 2286 1180 2292 1181
rect 2286 1176 2287 1180
rect 2291 1176 2292 1180
rect 2286 1175 2292 1176
rect 2422 1180 2428 1181
rect 2422 1176 2423 1180
rect 2427 1176 2428 1180
rect 2422 1175 2428 1176
rect 2566 1180 2572 1181
rect 2566 1176 2567 1180
rect 2571 1176 2572 1180
rect 2566 1175 2572 1176
rect 2702 1180 2708 1181
rect 2702 1176 2703 1180
rect 2707 1176 2708 1180
rect 2702 1175 2708 1176
rect 2838 1180 2844 1181
rect 2838 1176 2839 1180
rect 2843 1176 2844 1180
rect 2838 1175 2844 1176
rect 2974 1180 2980 1181
rect 2974 1176 2975 1180
rect 2979 1176 2980 1180
rect 2974 1175 2980 1176
rect 3110 1180 3116 1181
rect 3110 1176 3111 1180
rect 3115 1176 3116 1180
rect 3110 1175 3116 1176
rect 3246 1180 3252 1181
rect 3246 1176 3247 1180
rect 3251 1176 3252 1180
rect 3246 1175 3252 1176
rect 3366 1180 3372 1181
rect 3366 1176 3367 1180
rect 3371 1176 3372 1180
rect 3464 1178 3466 1197
rect 3366 1175 3372 1176
rect 3462 1177 3468 1178
rect 1806 1172 1812 1173
rect 3462 1173 3463 1177
rect 3467 1173 3468 1177
rect 3462 1172 3468 1173
rect 134 1161 140 1162
rect 110 1160 116 1161
rect 110 1156 111 1160
rect 115 1156 116 1160
rect 134 1157 135 1161
rect 139 1157 140 1161
rect 134 1156 140 1157
rect 230 1161 236 1162
rect 230 1157 231 1161
rect 235 1157 236 1161
rect 230 1156 236 1157
rect 358 1161 364 1162
rect 358 1157 359 1161
rect 363 1157 364 1161
rect 358 1156 364 1157
rect 486 1161 492 1162
rect 486 1157 487 1161
rect 491 1157 492 1161
rect 486 1156 492 1157
rect 614 1161 620 1162
rect 614 1157 615 1161
rect 619 1157 620 1161
rect 614 1156 620 1157
rect 742 1161 748 1162
rect 742 1157 743 1161
rect 747 1157 748 1161
rect 742 1156 748 1157
rect 870 1161 876 1162
rect 870 1157 871 1161
rect 875 1157 876 1161
rect 870 1156 876 1157
rect 990 1161 996 1162
rect 990 1157 991 1161
rect 995 1157 996 1161
rect 990 1156 996 1157
rect 1118 1161 1124 1162
rect 1118 1157 1119 1161
rect 1123 1157 1124 1161
rect 1118 1156 1124 1157
rect 1246 1161 1252 1162
rect 1934 1161 1940 1162
rect 1246 1157 1247 1161
rect 1251 1157 1252 1161
rect 1246 1156 1252 1157
rect 1766 1160 1772 1161
rect 1766 1156 1767 1160
rect 1771 1156 1772 1160
rect 110 1155 116 1156
rect 112 1135 114 1155
rect 136 1135 138 1156
rect 232 1135 234 1156
rect 360 1135 362 1156
rect 488 1135 490 1156
rect 616 1135 618 1156
rect 744 1135 746 1156
rect 872 1135 874 1156
rect 992 1135 994 1156
rect 1120 1135 1122 1156
rect 1248 1135 1250 1156
rect 1766 1155 1772 1156
rect 1806 1160 1812 1161
rect 1806 1156 1807 1160
rect 1811 1156 1812 1160
rect 1934 1157 1935 1161
rect 1939 1157 1940 1161
rect 1934 1156 1940 1157
rect 2038 1161 2044 1162
rect 2038 1157 2039 1161
rect 2043 1157 2044 1161
rect 2038 1156 2044 1157
rect 2158 1161 2164 1162
rect 2158 1157 2159 1161
rect 2163 1157 2164 1161
rect 2158 1156 2164 1157
rect 2286 1161 2292 1162
rect 2286 1157 2287 1161
rect 2291 1157 2292 1161
rect 2286 1156 2292 1157
rect 2422 1161 2428 1162
rect 2422 1157 2423 1161
rect 2427 1157 2428 1161
rect 2422 1156 2428 1157
rect 2566 1161 2572 1162
rect 2566 1157 2567 1161
rect 2571 1157 2572 1161
rect 2566 1156 2572 1157
rect 2702 1161 2708 1162
rect 2702 1157 2703 1161
rect 2707 1157 2708 1161
rect 2702 1156 2708 1157
rect 2838 1161 2844 1162
rect 2838 1157 2839 1161
rect 2843 1157 2844 1161
rect 2838 1156 2844 1157
rect 2974 1161 2980 1162
rect 2974 1157 2975 1161
rect 2979 1157 2980 1161
rect 2974 1156 2980 1157
rect 3110 1161 3116 1162
rect 3110 1157 3111 1161
rect 3115 1157 3116 1161
rect 3110 1156 3116 1157
rect 3246 1161 3252 1162
rect 3246 1157 3247 1161
rect 3251 1157 3252 1161
rect 3246 1156 3252 1157
rect 3366 1161 3372 1162
rect 3366 1157 3367 1161
rect 3371 1157 3372 1161
rect 3366 1156 3372 1157
rect 3462 1160 3468 1161
rect 3462 1156 3463 1160
rect 3467 1156 3468 1160
rect 1806 1155 1812 1156
rect 1768 1135 1770 1155
rect 111 1134 115 1135
rect 111 1129 115 1130
rect 135 1134 139 1135
rect 135 1129 139 1130
rect 231 1134 235 1135
rect 231 1129 235 1130
rect 247 1134 251 1135
rect 247 1129 251 1130
rect 359 1134 363 1135
rect 359 1129 363 1130
rect 367 1134 371 1135
rect 367 1129 371 1130
rect 487 1134 491 1135
rect 487 1129 491 1130
rect 495 1134 499 1135
rect 495 1129 499 1130
rect 615 1134 619 1135
rect 615 1129 619 1130
rect 623 1134 627 1135
rect 623 1129 627 1130
rect 743 1134 747 1135
rect 743 1129 747 1130
rect 759 1134 763 1135
rect 759 1129 763 1130
rect 871 1134 875 1135
rect 871 1129 875 1130
rect 887 1134 891 1135
rect 887 1129 891 1130
rect 991 1134 995 1135
rect 991 1129 995 1130
rect 1015 1134 1019 1135
rect 1015 1129 1019 1130
rect 1119 1134 1123 1135
rect 1119 1129 1123 1130
rect 1143 1134 1147 1135
rect 1143 1129 1147 1130
rect 1247 1134 1251 1135
rect 1247 1129 1251 1130
rect 1271 1134 1275 1135
rect 1271 1129 1275 1130
rect 1399 1134 1403 1135
rect 1399 1129 1403 1130
rect 1767 1134 1771 1135
rect 1808 1131 1810 1155
rect 1936 1131 1938 1156
rect 2040 1131 2042 1156
rect 2160 1131 2162 1156
rect 2288 1131 2290 1156
rect 2424 1131 2426 1156
rect 2568 1131 2570 1156
rect 2704 1131 2706 1156
rect 2840 1131 2842 1156
rect 2976 1131 2978 1156
rect 3112 1131 3114 1156
rect 3248 1131 3250 1156
rect 3368 1131 3370 1156
rect 3462 1155 3468 1156
rect 3464 1131 3466 1155
rect 1767 1129 1771 1130
rect 1807 1130 1811 1131
rect 112 1113 114 1129
rect 110 1112 116 1113
rect 248 1112 250 1129
rect 368 1112 370 1129
rect 496 1112 498 1129
rect 624 1112 626 1129
rect 760 1112 762 1129
rect 888 1112 890 1129
rect 1016 1112 1018 1129
rect 1144 1112 1146 1129
rect 1272 1112 1274 1129
rect 1400 1112 1402 1129
rect 1768 1113 1770 1129
rect 1807 1125 1811 1126
rect 1935 1130 1939 1131
rect 1935 1125 1939 1126
rect 1943 1130 1947 1131
rect 1943 1125 1947 1126
rect 2039 1130 2043 1131
rect 2039 1125 2043 1126
rect 2063 1130 2067 1131
rect 2063 1125 2067 1126
rect 2159 1130 2163 1131
rect 2159 1125 2163 1126
rect 2191 1130 2195 1131
rect 2191 1125 2195 1126
rect 2287 1130 2291 1131
rect 2287 1125 2291 1126
rect 2319 1130 2323 1131
rect 2319 1125 2323 1126
rect 2423 1130 2427 1131
rect 2423 1125 2427 1126
rect 2455 1130 2459 1131
rect 2455 1125 2459 1126
rect 2567 1130 2571 1131
rect 2567 1125 2571 1126
rect 2599 1130 2603 1131
rect 2599 1125 2603 1126
rect 2703 1130 2707 1131
rect 2703 1125 2707 1126
rect 2751 1130 2755 1131
rect 2751 1125 2755 1126
rect 2839 1130 2843 1131
rect 2839 1125 2843 1126
rect 2903 1130 2907 1131
rect 2903 1125 2907 1126
rect 2975 1130 2979 1131
rect 2975 1125 2979 1126
rect 3063 1130 3067 1131
rect 3063 1125 3067 1126
rect 3111 1130 3115 1131
rect 3111 1125 3115 1126
rect 3223 1130 3227 1131
rect 3223 1125 3227 1126
rect 3247 1130 3251 1131
rect 3247 1125 3251 1126
rect 3367 1130 3371 1131
rect 3367 1125 3371 1126
rect 3463 1130 3467 1131
rect 3463 1125 3467 1126
rect 1766 1112 1772 1113
rect 110 1108 111 1112
rect 115 1108 116 1112
rect 110 1107 116 1108
rect 246 1111 252 1112
rect 246 1107 247 1111
rect 251 1107 252 1111
rect 246 1106 252 1107
rect 366 1111 372 1112
rect 366 1107 367 1111
rect 371 1107 372 1111
rect 366 1106 372 1107
rect 494 1111 500 1112
rect 494 1107 495 1111
rect 499 1107 500 1111
rect 494 1106 500 1107
rect 622 1111 628 1112
rect 622 1107 623 1111
rect 627 1107 628 1111
rect 622 1106 628 1107
rect 758 1111 764 1112
rect 758 1107 759 1111
rect 763 1107 764 1111
rect 758 1106 764 1107
rect 886 1111 892 1112
rect 886 1107 887 1111
rect 891 1107 892 1111
rect 886 1106 892 1107
rect 1014 1111 1020 1112
rect 1014 1107 1015 1111
rect 1019 1107 1020 1111
rect 1014 1106 1020 1107
rect 1142 1111 1148 1112
rect 1142 1107 1143 1111
rect 1147 1107 1148 1111
rect 1142 1106 1148 1107
rect 1270 1111 1276 1112
rect 1270 1107 1271 1111
rect 1275 1107 1276 1111
rect 1270 1106 1276 1107
rect 1398 1111 1404 1112
rect 1398 1107 1399 1111
rect 1403 1107 1404 1111
rect 1766 1108 1767 1112
rect 1771 1108 1772 1112
rect 1808 1109 1810 1125
rect 1766 1107 1772 1108
rect 1806 1108 1812 1109
rect 1944 1108 1946 1125
rect 2064 1108 2066 1125
rect 2192 1108 2194 1125
rect 2320 1108 2322 1125
rect 2456 1108 2458 1125
rect 2600 1108 2602 1125
rect 2752 1108 2754 1125
rect 2904 1108 2906 1125
rect 3064 1108 3066 1125
rect 3224 1108 3226 1125
rect 3368 1108 3370 1125
rect 3464 1109 3466 1125
rect 3462 1108 3468 1109
rect 1398 1106 1404 1107
rect 1806 1104 1807 1108
rect 1811 1104 1812 1108
rect 1806 1103 1812 1104
rect 1942 1107 1948 1108
rect 1942 1103 1943 1107
rect 1947 1103 1948 1107
rect 1942 1102 1948 1103
rect 2062 1107 2068 1108
rect 2062 1103 2063 1107
rect 2067 1103 2068 1107
rect 2062 1102 2068 1103
rect 2190 1107 2196 1108
rect 2190 1103 2191 1107
rect 2195 1103 2196 1107
rect 2190 1102 2196 1103
rect 2318 1107 2324 1108
rect 2318 1103 2319 1107
rect 2323 1103 2324 1107
rect 2318 1102 2324 1103
rect 2454 1107 2460 1108
rect 2454 1103 2455 1107
rect 2459 1103 2460 1107
rect 2454 1102 2460 1103
rect 2598 1107 2604 1108
rect 2598 1103 2599 1107
rect 2603 1103 2604 1107
rect 2598 1102 2604 1103
rect 2750 1107 2756 1108
rect 2750 1103 2751 1107
rect 2755 1103 2756 1107
rect 2750 1102 2756 1103
rect 2902 1107 2908 1108
rect 2902 1103 2903 1107
rect 2907 1103 2908 1107
rect 2902 1102 2908 1103
rect 3062 1107 3068 1108
rect 3062 1103 3063 1107
rect 3067 1103 3068 1107
rect 3062 1102 3068 1103
rect 3222 1107 3228 1108
rect 3222 1103 3223 1107
rect 3227 1103 3228 1107
rect 3222 1102 3228 1103
rect 3366 1107 3372 1108
rect 3366 1103 3367 1107
rect 3371 1103 3372 1107
rect 3462 1104 3463 1108
rect 3467 1104 3468 1108
rect 3462 1103 3468 1104
rect 3366 1102 3372 1103
rect 110 1095 116 1096
rect 110 1091 111 1095
rect 115 1091 116 1095
rect 1766 1095 1772 1096
rect 110 1090 116 1091
rect 246 1092 252 1093
rect 112 1067 114 1090
rect 246 1088 247 1092
rect 251 1088 252 1092
rect 246 1087 252 1088
rect 366 1092 372 1093
rect 366 1088 367 1092
rect 371 1088 372 1092
rect 366 1087 372 1088
rect 494 1092 500 1093
rect 494 1088 495 1092
rect 499 1088 500 1092
rect 494 1087 500 1088
rect 622 1092 628 1093
rect 622 1088 623 1092
rect 627 1088 628 1092
rect 622 1087 628 1088
rect 758 1092 764 1093
rect 758 1088 759 1092
rect 763 1088 764 1092
rect 758 1087 764 1088
rect 886 1092 892 1093
rect 886 1088 887 1092
rect 891 1088 892 1092
rect 886 1087 892 1088
rect 1014 1092 1020 1093
rect 1014 1088 1015 1092
rect 1019 1088 1020 1092
rect 1014 1087 1020 1088
rect 1142 1092 1148 1093
rect 1142 1088 1143 1092
rect 1147 1088 1148 1092
rect 1142 1087 1148 1088
rect 1270 1092 1276 1093
rect 1270 1088 1271 1092
rect 1275 1088 1276 1092
rect 1270 1087 1276 1088
rect 1398 1092 1404 1093
rect 1398 1088 1399 1092
rect 1403 1088 1404 1092
rect 1766 1091 1767 1095
rect 1771 1091 1772 1095
rect 1766 1090 1772 1091
rect 1806 1091 1812 1092
rect 1398 1087 1404 1088
rect 248 1067 250 1087
rect 368 1067 370 1087
rect 496 1067 498 1087
rect 624 1067 626 1087
rect 760 1067 762 1087
rect 888 1067 890 1087
rect 1016 1067 1018 1087
rect 1144 1067 1146 1087
rect 1272 1067 1274 1087
rect 1400 1067 1402 1087
rect 1768 1067 1770 1090
rect 1806 1087 1807 1091
rect 1811 1087 1812 1091
rect 3462 1091 3468 1092
rect 1806 1086 1812 1087
rect 1942 1088 1948 1089
rect 111 1066 115 1067
rect 111 1061 115 1062
rect 247 1066 251 1067
rect 247 1061 251 1062
rect 367 1066 371 1067
rect 367 1061 371 1062
rect 431 1066 435 1067
rect 431 1061 435 1062
rect 495 1066 499 1067
rect 495 1061 499 1062
rect 543 1066 547 1067
rect 543 1061 547 1062
rect 623 1066 627 1067
rect 623 1061 627 1062
rect 663 1066 667 1067
rect 663 1061 667 1062
rect 759 1066 763 1067
rect 759 1061 763 1062
rect 791 1066 795 1067
rect 791 1061 795 1062
rect 887 1066 891 1067
rect 887 1061 891 1062
rect 919 1066 923 1067
rect 919 1061 923 1062
rect 1015 1066 1019 1067
rect 1015 1061 1019 1062
rect 1039 1066 1043 1067
rect 1039 1061 1043 1062
rect 1143 1066 1147 1067
rect 1143 1061 1147 1062
rect 1159 1066 1163 1067
rect 1159 1061 1163 1062
rect 1271 1066 1275 1067
rect 1271 1061 1275 1062
rect 1279 1066 1283 1067
rect 1279 1061 1283 1062
rect 1399 1066 1403 1067
rect 1399 1061 1403 1062
rect 1407 1066 1411 1067
rect 1407 1061 1411 1062
rect 1535 1066 1539 1067
rect 1535 1061 1539 1062
rect 1767 1066 1771 1067
rect 1808 1063 1810 1086
rect 1942 1084 1943 1088
rect 1947 1084 1948 1088
rect 1942 1083 1948 1084
rect 2062 1088 2068 1089
rect 2062 1084 2063 1088
rect 2067 1084 2068 1088
rect 2062 1083 2068 1084
rect 2190 1088 2196 1089
rect 2190 1084 2191 1088
rect 2195 1084 2196 1088
rect 2190 1083 2196 1084
rect 2318 1088 2324 1089
rect 2318 1084 2319 1088
rect 2323 1084 2324 1088
rect 2318 1083 2324 1084
rect 2454 1088 2460 1089
rect 2454 1084 2455 1088
rect 2459 1084 2460 1088
rect 2454 1083 2460 1084
rect 2598 1088 2604 1089
rect 2598 1084 2599 1088
rect 2603 1084 2604 1088
rect 2598 1083 2604 1084
rect 2750 1088 2756 1089
rect 2750 1084 2751 1088
rect 2755 1084 2756 1088
rect 2750 1083 2756 1084
rect 2902 1088 2908 1089
rect 2902 1084 2903 1088
rect 2907 1084 2908 1088
rect 2902 1083 2908 1084
rect 3062 1088 3068 1089
rect 3062 1084 3063 1088
rect 3067 1084 3068 1088
rect 3062 1083 3068 1084
rect 3222 1088 3228 1089
rect 3222 1084 3223 1088
rect 3227 1084 3228 1088
rect 3222 1083 3228 1084
rect 3366 1088 3372 1089
rect 3366 1084 3367 1088
rect 3371 1084 3372 1088
rect 3462 1087 3463 1091
rect 3467 1087 3468 1091
rect 3462 1086 3468 1087
rect 3366 1083 3372 1084
rect 1944 1063 1946 1083
rect 2064 1063 2066 1083
rect 2192 1063 2194 1083
rect 2320 1063 2322 1083
rect 2456 1063 2458 1083
rect 2600 1063 2602 1083
rect 2752 1063 2754 1083
rect 2904 1063 2906 1083
rect 3064 1063 3066 1083
rect 3224 1063 3226 1083
rect 3368 1063 3370 1083
rect 3464 1063 3466 1086
rect 1767 1061 1771 1062
rect 1807 1062 1811 1063
rect 112 1042 114 1061
rect 432 1045 434 1061
rect 544 1045 546 1061
rect 664 1045 666 1061
rect 792 1045 794 1061
rect 920 1045 922 1061
rect 1040 1045 1042 1061
rect 1160 1045 1162 1061
rect 1280 1045 1282 1061
rect 1408 1045 1410 1061
rect 1536 1045 1538 1061
rect 430 1044 436 1045
rect 110 1041 116 1042
rect 110 1037 111 1041
rect 115 1037 116 1041
rect 430 1040 431 1044
rect 435 1040 436 1044
rect 430 1039 436 1040
rect 542 1044 548 1045
rect 542 1040 543 1044
rect 547 1040 548 1044
rect 542 1039 548 1040
rect 662 1044 668 1045
rect 662 1040 663 1044
rect 667 1040 668 1044
rect 662 1039 668 1040
rect 790 1044 796 1045
rect 790 1040 791 1044
rect 795 1040 796 1044
rect 790 1039 796 1040
rect 918 1044 924 1045
rect 918 1040 919 1044
rect 923 1040 924 1044
rect 918 1039 924 1040
rect 1038 1044 1044 1045
rect 1038 1040 1039 1044
rect 1043 1040 1044 1044
rect 1038 1039 1044 1040
rect 1158 1044 1164 1045
rect 1158 1040 1159 1044
rect 1163 1040 1164 1044
rect 1158 1039 1164 1040
rect 1278 1044 1284 1045
rect 1278 1040 1279 1044
rect 1283 1040 1284 1044
rect 1278 1039 1284 1040
rect 1406 1044 1412 1045
rect 1406 1040 1407 1044
rect 1411 1040 1412 1044
rect 1406 1039 1412 1040
rect 1534 1044 1540 1045
rect 1534 1040 1535 1044
rect 1539 1040 1540 1044
rect 1768 1042 1770 1061
rect 1807 1057 1811 1058
rect 1847 1062 1851 1063
rect 1847 1057 1851 1058
rect 1943 1062 1947 1063
rect 1943 1057 1947 1058
rect 1983 1062 1987 1063
rect 1983 1057 1987 1058
rect 2063 1062 2067 1063
rect 2063 1057 2067 1058
rect 2119 1062 2123 1063
rect 2119 1057 2123 1058
rect 2191 1062 2195 1063
rect 2191 1057 2195 1058
rect 2255 1062 2259 1063
rect 2255 1057 2259 1058
rect 2319 1062 2323 1063
rect 2319 1057 2323 1058
rect 2391 1062 2395 1063
rect 2391 1057 2395 1058
rect 2455 1062 2459 1063
rect 2455 1057 2459 1058
rect 2543 1062 2547 1063
rect 2543 1057 2547 1058
rect 2599 1062 2603 1063
rect 2599 1057 2603 1058
rect 2703 1062 2707 1063
rect 2703 1057 2707 1058
rect 2751 1062 2755 1063
rect 2751 1057 2755 1058
rect 2863 1062 2867 1063
rect 2863 1057 2867 1058
rect 2903 1062 2907 1063
rect 2903 1057 2907 1058
rect 3031 1062 3035 1063
rect 3031 1057 3035 1058
rect 3063 1062 3067 1063
rect 3063 1057 3067 1058
rect 3207 1062 3211 1063
rect 3207 1057 3211 1058
rect 3223 1062 3227 1063
rect 3223 1057 3227 1058
rect 3367 1062 3371 1063
rect 3367 1057 3371 1058
rect 3463 1062 3467 1063
rect 3463 1057 3467 1058
rect 1534 1039 1540 1040
rect 1766 1041 1772 1042
rect 110 1036 116 1037
rect 1766 1037 1767 1041
rect 1771 1037 1772 1041
rect 1808 1038 1810 1057
rect 1848 1041 1850 1057
rect 1984 1041 1986 1057
rect 2120 1041 2122 1057
rect 2256 1041 2258 1057
rect 2392 1041 2394 1057
rect 2544 1041 2546 1057
rect 2704 1041 2706 1057
rect 2864 1041 2866 1057
rect 3032 1041 3034 1057
rect 3208 1041 3210 1057
rect 3368 1041 3370 1057
rect 1846 1040 1852 1041
rect 1766 1036 1772 1037
rect 1806 1037 1812 1038
rect 1806 1033 1807 1037
rect 1811 1033 1812 1037
rect 1846 1036 1847 1040
rect 1851 1036 1852 1040
rect 1846 1035 1852 1036
rect 1982 1040 1988 1041
rect 1982 1036 1983 1040
rect 1987 1036 1988 1040
rect 1982 1035 1988 1036
rect 2118 1040 2124 1041
rect 2118 1036 2119 1040
rect 2123 1036 2124 1040
rect 2118 1035 2124 1036
rect 2254 1040 2260 1041
rect 2254 1036 2255 1040
rect 2259 1036 2260 1040
rect 2254 1035 2260 1036
rect 2390 1040 2396 1041
rect 2390 1036 2391 1040
rect 2395 1036 2396 1040
rect 2390 1035 2396 1036
rect 2542 1040 2548 1041
rect 2542 1036 2543 1040
rect 2547 1036 2548 1040
rect 2542 1035 2548 1036
rect 2702 1040 2708 1041
rect 2702 1036 2703 1040
rect 2707 1036 2708 1040
rect 2702 1035 2708 1036
rect 2862 1040 2868 1041
rect 2862 1036 2863 1040
rect 2867 1036 2868 1040
rect 2862 1035 2868 1036
rect 3030 1040 3036 1041
rect 3030 1036 3031 1040
rect 3035 1036 3036 1040
rect 3030 1035 3036 1036
rect 3206 1040 3212 1041
rect 3206 1036 3207 1040
rect 3211 1036 3212 1040
rect 3206 1035 3212 1036
rect 3366 1040 3372 1041
rect 3366 1036 3367 1040
rect 3371 1036 3372 1040
rect 3464 1038 3466 1057
rect 3366 1035 3372 1036
rect 3462 1037 3468 1038
rect 1806 1032 1812 1033
rect 3462 1033 3463 1037
rect 3467 1033 3468 1037
rect 3462 1032 3468 1033
rect 430 1025 436 1026
rect 110 1024 116 1025
rect 110 1020 111 1024
rect 115 1020 116 1024
rect 430 1021 431 1025
rect 435 1021 436 1025
rect 430 1020 436 1021
rect 542 1025 548 1026
rect 542 1021 543 1025
rect 547 1021 548 1025
rect 542 1020 548 1021
rect 662 1025 668 1026
rect 662 1021 663 1025
rect 667 1021 668 1025
rect 662 1020 668 1021
rect 790 1025 796 1026
rect 790 1021 791 1025
rect 795 1021 796 1025
rect 790 1020 796 1021
rect 918 1025 924 1026
rect 918 1021 919 1025
rect 923 1021 924 1025
rect 918 1020 924 1021
rect 1038 1025 1044 1026
rect 1038 1021 1039 1025
rect 1043 1021 1044 1025
rect 1038 1020 1044 1021
rect 1158 1025 1164 1026
rect 1158 1021 1159 1025
rect 1163 1021 1164 1025
rect 1158 1020 1164 1021
rect 1278 1025 1284 1026
rect 1278 1021 1279 1025
rect 1283 1021 1284 1025
rect 1278 1020 1284 1021
rect 1406 1025 1412 1026
rect 1406 1021 1407 1025
rect 1411 1021 1412 1025
rect 1406 1020 1412 1021
rect 1534 1025 1540 1026
rect 1534 1021 1535 1025
rect 1539 1021 1540 1025
rect 1534 1020 1540 1021
rect 1766 1024 1772 1025
rect 1766 1020 1767 1024
rect 1771 1020 1772 1024
rect 1846 1021 1852 1022
rect 110 1019 116 1020
rect 112 995 114 1019
rect 432 995 434 1020
rect 544 995 546 1020
rect 664 995 666 1020
rect 792 995 794 1020
rect 920 995 922 1020
rect 1040 995 1042 1020
rect 1160 995 1162 1020
rect 1280 995 1282 1020
rect 1408 995 1410 1020
rect 1536 995 1538 1020
rect 1766 1019 1772 1020
rect 1806 1020 1812 1021
rect 1768 995 1770 1019
rect 1806 1016 1807 1020
rect 1811 1016 1812 1020
rect 1846 1017 1847 1021
rect 1851 1017 1852 1021
rect 1846 1016 1852 1017
rect 1982 1021 1988 1022
rect 1982 1017 1983 1021
rect 1987 1017 1988 1021
rect 1982 1016 1988 1017
rect 2118 1021 2124 1022
rect 2118 1017 2119 1021
rect 2123 1017 2124 1021
rect 2118 1016 2124 1017
rect 2254 1021 2260 1022
rect 2254 1017 2255 1021
rect 2259 1017 2260 1021
rect 2254 1016 2260 1017
rect 2390 1021 2396 1022
rect 2390 1017 2391 1021
rect 2395 1017 2396 1021
rect 2390 1016 2396 1017
rect 2542 1021 2548 1022
rect 2542 1017 2543 1021
rect 2547 1017 2548 1021
rect 2542 1016 2548 1017
rect 2702 1021 2708 1022
rect 2702 1017 2703 1021
rect 2707 1017 2708 1021
rect 2702 1016 2708 1017
rect 2862 1021 2868 1022
rect 2862 1017 2863 1021
rect 2867 1017 2868 1021
rect 2862 1016 2868 1017
rect 3030 1021 3036 1022
rect 3030 1017 3031 1021
rect 3035 1017 3036 1021
rect 3030 1016 3036 1017
rect 3206 1021 3212 1022
rect 3206 1017 3207 1021
rect 3211 1017 3212 1021
rect 3206 1016 3212 1017
rect 3366 1021 3372 1022
rect 3366 1017 3367 1021
rect 3371 1017 3372 1021
rect 3366 1016 3372 1017
rect 3462 1020 3468 1021
rect 3462 1016 3463 1020
rect 3467 1016 3468 1020
rect 1806 1015 1812 1016
rect 1808 995 1810 1015
rect 1848 995 1850 1016
rect 1984 995 1986 1016
rect 2120 995 2122 1016
rect 2256 995 2258 1016
rect 2392 995 2394 1016
rect 2544 995 2546 1016
rect 2704 995 2706 1016
rect 2864 995 2866 1016
rect 3032 995 3034 1016
rect 3208 995 3210 1016
rect 3368 995 3370 1016
rect 3462 1015 3468 1016
rect 3464 995 3466 1015
rect 111 994 115 995
rect 111 989 115 990
rect 431 994 435 995
rect 431 989 435 990
rect 543 994 547 995
rect 543 989 547 990
rect 567 994 571 995
rect 567 989 571 990
rect 663 994 667 995
rect 663 989 667 990
rect 679 994 683 995
rect 679 989 683 990
rect 791 994 795 995
rect 791 989 795 990
rect 911 994 915 995
rect 911 989 915 990
rect 919 994 923 995
rect 919 989 923 990
rect 1031 994 1035 995
rect 1031 989 1035 990
rect 1039 994 1043 995
rect 1039 989 1043 990
rect 1143 994 1147 995
rect 1143 989 1147 990
rect 1159 994 1163 995
rect 1159 989 1163 990
rect 1255 994 1259 995
rect 1255 989 1259 990
rect 1279 994 1283 995
rect 1279 989 1283 990
rect 1359 994 1363 995
rect 1359 989 1363 990
rect 1407 994 1411 995
rect 1407 989 1411 990
rect 1471 994 1475 995
rect 1471 989 1475 990
rect 1535 994 1539 995
rect 1535 989 1539 990
rect 1583 994 1587 995
rect 1583 989 1587 990
rect 1671 994 1675 995
rect 1671 989 1675 990
rect 1767 994 1771 995
rect 1767 989 1771 990
rect 1807 994 1811 995
rect 1807 989 1811 990
rect 1831 994 1835 995
rect 1831 989 1835 990
rect 1847 994 1851 995
rect 1847 989 1851 990
rect 1975 994 1979 995
rect 1975 989 1979 990
rect 1983 994 1987 995
rect 1983 989 1987 990
rect 2119 994 2123 995
rect 2119 989 2123 990
rect 2135 994 2139 995
rect 2135 989 2139 990
rect 2255 994 2259 995
rect 2255 989 2259 990
rect 2295 994 2299 995
rect 2295 989 2299 990
rect 2391 994 2395 995
rect 2391 989 2395 990
rect 2463 994 2467 995
rect 2463 989 2467 990
rect 2543 994 2547 995
rect 2543 989 2547 990
rect 2631 994 2635 995
rect 2631 989 2635 990
rect 2703 994 2707 995
rect 2703 989 2707 990
rect 2807 994 2811 995
rect 2807 989 2811 990
rect 2863 994 2867 995
rect 2863 989 2867 990
rect 2991 994 2995 995
rect 2991 989 2995 990
rect 3031 994 3035 995
rect 3031 989 3035 990
rect 3183 994 3187 995
rect 3183 989 3187 990
rect 3207 994 3211 995
rect 3207 989 3211 990
rect 3367 994 3371 995
rect 3367 989 3371 990
rect 3463 994 3467 995
rect 3463 989 3467 990
rect 112 973 114 989
rect 110 972 116 973
rect 568 972 570 989
rect 680 972 682 989
rect 792 972 794 989
rect 912 972 914 989
rect 1032 972 1034 989
rect 1144 972 1146 989
rect 1256 972 1258 989
rect 1360 972 1362 989
rect 1472 972 1474 989
rect 1584 972 1586 989
rect 1672 972 1674 989
rect 1768 973 1770 989
rect 1808 973 1810 989
rect 1766 972 1772 973
rect 110 968 111 972
rect 115 968 116 972
rect 110 967 116 968
rect 566 971 572 972
rect 566 967 567 971
rect 571 967 572 971
rect 566 966 572 967
rect 678 971 684 972
rect 678 967 679 971
rect 683 967 684 971
rect 678 966 684 967
rect 790 971 796 972
rect 790 967 791 971
rect 795 967 796 971
rect 790 966 796 967
rect 910 971 916 972
rect 910 967 911 971
rect 915 967 916 971
rect 910 966 916 967
rect 1030 971 1036 972
rect 1030 967 1031 971
rect 1035 967 1036 971
rect 1030 966 1036 967
rect 1142 971 1148 972
rect 1142 967 1143 971
rect 1147 967 1148 971
rect 1142 966 1148 967
rect 1254 971 1260 972
rect 1254 967 1255 971
rect 1259 967 1260 971
rect 1254 966 1260 967
rect 1358 971 1364 972
rect 1358 967 1359 971
rect 1363 967 1364 971
rect 1358 966 1364 967
rect 1470 971 1476 972
rect 1470 967 1471 971
rect 1475 967 1476 971
rect 1470 966 1476 967
rect 1582 971 1588 972
rect 1582 967 1583 971
rect 1587 967 1588 971
rect 1582 966 1588 967
rect 1670 971 1676 972
rect 1670 967 1671 971
rect 1675 967 1676 971
rect 1766 968 1767 972
rect 1771 968 1772 972
rect 1766 967 1772 968
rect 1806 972 1812 973
rect 1832 972 1834 989
rect 1976 972 1978 989
rect 2136 972 2138 989
rect 2296 972 2298 989
rect 2464 972 2466 989
rect 2632 972 2634 989
rect 2808 972 2810 989
rect 2992 972 2994 989
rect 3184 972 3186 989
rect 3368 972 3370 989
rect 3464 973 3466 989
rect 3462 972 3468 973
rect 1806 968 1807 972
rect 1811 968 1812 972
rect 1806 967 1812 968
rect 1830 971 1836 972
rect 1830 967 1831 971
rect 1835 967 1836 971
rect 1670 966 1676 967
rect 1830 966 1836 967
rect 1974 971 1980 972
rect 1974 967 1975 971
rect 1979 967 1980 971
rect 1974 966 1980 967
rect 2134 971 2140 972
rect 2134 967 2135 971
rect 2139 967 2140 971
rect 2134 966 2140 967
rect 2294 971 2300 972
rect 2294 967 2295 971
rect 2299 967 2300 971
rect 2294 966 2300 967
rect 2462 971 2468 972
rect 2462 967 2463 971
rect 2467 967 2468 971
rect 2462 966 2468 967
rect 2630 971 2636 972
rect 2630 967 2631 971
rect 2635 967 2636 971
rect 2630 966 2636 967
rect 2806 971 2812 972
rect 2806 967 2807 971
rect 2811 967 2812 971
rect 2806 966 2812 967
rect 2990 971 2996 972
rect 2990 967 2991 971
rect 2995 967 2996 971
rect 2990 966 2996 967
rect 3182 971 3188 972
rect 3182 967 3183 971
rect 3187 967 3188 971
rect 3182 966 3188 967
rect 3366 971 3372 972
rect 3366 967 3367 971
rect 3371 967 3372 971
rect 3462 968 3463 972
rect 3467 968 3468 972
rect 3462 967 3468 968
rect 3366 966 3372 967
rect 110 955 116 956
rect 110 951 111 955
rect 115 951 116 955
rect 1766 955 1772 956
rect 110 950 116 951
rect 566 952 572 953
rect 112 927 114 950
rect 566 948 567 952
rect 571 948 572 952
rect 566 947 572 948
rect 678 952 684 953
rect 678 948 679 952
rect 683 948 684 952
rect 678 947 684 948
rect 790 952 796 953
rect 790 948 791 952
rect 795 948 796 952
rect 790 947 796 948
rect 910 952 916 953
rect 910 948 911 952
rect 915 948 916 952
rect 910 947 916 948
rect 1030 952 1036 953
rect 1030 948 1031 952
rect 1035 948 1036 952
rect 1030 947 1036 948
rect 1142 952 1148 953
rect 1142 948 1143 952
rect 1147 948 1148 952
rect 1142 947 1148 948
rect 1254 952 1260 953
rect 1254 948 1255 952
rect 1259 948 1260 952
rect 1254 947 1260 948
rect 1358 952 1364 953
rect 1358 948 1359 952
rect 1363 948 1364 952
rect 1358 947 1364 948
rect 1470 952 1476 953
rect 1470 948 1471 952
rect 1475 948 1476 952
rect 1470 947 1476 948
rect 1582 952 1588 953
rect 1582 948 1583 952
rect 1587 948 1588 952
rect 1582 947 1588 948
rect 1670 952 1676 953
rect 1670 948 1671 952
rect 1675 948 1676 952
rect 1766 951 1767 955
rect 1771 951 1772 955
rect 1766 950 1772 951
rect 1806 955 1812 956
rect 1806 951 1807 955
rect 1811 951 1812 955
rect 3462 955 3468 956
rect 1806 950 1812 951
rect 1830 952 1836 953
rect 1670 947 1676 948
rect 568 927 570 947
rect 680 927 682 947
rect 792 927 794 947
rect 912 927 914 947
rect 1032 927 1034 947
rect 1144 927 1146 947
rect 1256 927 1258 947
rect 1360 927 1362 947
rect 1472 927 1474 947
rect 1584 927 1586 947
rect 1672 927 1674 947
rect 1768 927 1770 950
rect 1808 931 1810 950
rect 1830 948 1831 952
rect 1835 948 1836 952
rect 1830 947 1836 948
rect 1974 952 1980 953
rect 1974 948 1975 952
rect 1979 948 1980 952
rect 1974 947 1980 948
rect 2134 952 2140 953
rect 2134 948 2135 952
rect 2139 948 2140 952
rect 2134 947 2140 948
rect 2294 952 2300 953
rect 2294 948 2295 952
rect 2299 948 2300 952
rect 2294 947 2300 948
rect 2462 952 2468 953
rect 2462 948 2463 952
rect 2467 948 2468 952
rect 2462 947 2468 948
rect 2630 952 2636 953
rect 2630 948 2631 952
rect 2635 948 2636 952
rect 2630 947 2636 948
rect 2806 952 2812 953
rect 2806 948 2807 952
rect 2811 948 2812 952
rect 2806 947 2812 948
rect 2990 952 2996 953
rect 2990 948 2991 952
rect 2995 948 2996 952
rect 2990 947 2996 948
rect 3182 952 3188 953
rect 3182 948 3183 952
rect 3187 948 3188 952
rect 3182 947 3188 948
rect 3366 952 3372 953
rect 3366 948 3367 952
rect 3371 948 3372 952
rect 3462 951 3463 955
rect 3467 951 3468 955
rect 3462 950 3468 951
rect 3366 947 3372 948
rect 1832 931 1834 947
rect 1976 931 1978 947
rect 2136 931 2138 947
rect 2296 931 2298 947
rect 2464 931 2466 947
rect 2632 931 2634 947
rect 2808 931 2810 947
rect 2992 931 2994 947
rect 3184 931 3186 947
rect 3368 931 3370 947
rect 3464 931 3466 950
rect 1807 930 1811 931
rect 111 926 115 927
rect 111 921 115 922
rect 415 926 419 927
rect 415 921 419 922
rect 559 926 563 927
rect 559 921 563 922
rect 567 926 571 927
rect 567 921 571 922
rect 679 926 683 927
rect 679 921 683 922
rect 727 926 731 927
rect 727 921 731 922
rect 791 926 795 927
rect 791 921 795 922
rect 911 926 915 927
rect 911 921 915 922
rect 1031 926 1035 927
rect 1031 921 1035 922
rect 1119 926 1123 927
rect 1119 921 1123 922
rect 1143 926 1147 927
rect 1143 921 1147 922
rect 1255 926 1259 927
rect 1255 921 1259 922
rect 1335 926 1339 927
rect 1335 921 1339 922
rect 1359 926 1363 927
rect 1359 921 1363 922
rect 1471 926 1475 927
rect 1471 921 1475 922
rect 1559 926 1563 927
rect 1559 921 1563 922
rect 1583 926 1587 927
rect 1583 921 1587 922
rect 1671 926 1675 927
rect 1671 921 1675 922
rect 1767 926 1771 927
rect 1807 925 1811 926
rect 1831 930 1835 931
rect 1831 925 1835 926
rect 1975 930 1979 931
rect 1975 925 1979 926
rect 2127 930 2131 931
rect 2127 925 2131 926
rect 2135 930 2139 931
rect 2135 925 2139 926
rect 2215 930 2219 931
rect 2215 925 2219 926
rect 2295 930 2299 931
rect 2295 925 2299 926
rect 2303 930 2307 931
rect 2303 925 2307 926
rect 2391 930 2395 931
rect 2391 925 2395 926
rect 2463 930 2467 931
rect 2463 925 2467 926
rect 2479 930 2483 931
rect 2479 925 2483 926
rect 2567 930 2571 931
rect 2567 925 2571 926
rect 2631 930 2635 931
rect 2631 925 2635 926
rect 2655 930 2659 931
rect 2655 925 2659 926
rect 2743 930 2747 931
rect 2743 925 2747 926
rect 2807 930 2811 931
rect 2807 925 2811 926
rect 2831 930 2835 931
rect 2831 925 2835 926
rect 2991 930 2995 931
rect 2991 925 2995 926
rect 3183 930 3187 931
rect 3183 925 3187 926
rect 3367 930 3371 931
rect 3367 925 3371 926
rect 3463 930 3467 931
rect 3463 925 3467 926
rect 1767 921 1771 922
rect 112 902 114 921
rect 416 905 418 921
rect 560 905 562 921
rect 728 905 730 921
rect 912 905 914 921
rect 1120 905 1122 921
rect 1336 905 1338 921
rect 1560 905 1562 921
rect 414 904 420 905
rect 110 901 116 902
rect 110 897 111 901
rect 115 897 116 901
rect 414 900 415 904
rect 419 900 420 904
rect 414 899 420 900
rect 558 904 564 905
rect 558 900 559 904
rect 563 900 564 904
rect 558 899 564 900
rect 726 904 732 905
rect 726 900 727 904
rect 731 900 732 904
rect 726 899 732 900
rect 910 904 916 905
rect 910 900 911 904
rect 915 900 916 904
rect 910 899 916 900
rect 1118 904 1124 905
rect 1118 900 1119 904
rect 1123 900 1124 904
rect 1118 899 1124 900
rect 1334 904 1340 905
rect 1334 900 1335 904
rect 1339 900 1340 904
rect 1334 899 1340 900
rect 1558 904 1564 905
rect 1558 900 1559 904
rect 1563 900 1564 904
rect 1768 902 1770 921
rect 1808 906 1810 925
rect 2128 909 2130 925
rect 2216 909 2218 925
rect 2304 909 2306 925
rect 2392 909 2394 925
rect 2480 909 2482 925
rect 2568 909 2570 925
rect 2656 909 2658 925
rect 2744 909 2746 925
rect 2832 909 2834 925
rect 2126 908 2132 909
rect 1806 905 1812 906
rect 1558 899 1564 900
rect 1766 901 1772 902
rect 110 896 116 897
rect 1766 897 1767 901
rect 1771 897 1772 901
rect 1806 901 1807 905
rect 1811 901 1812 905
rect 2126 904 2127 908
rect 2131 904 2132 908
rect 2126 903 2132 904
rect 2214 908 2220 909
rect 2214 904 2215 908
rect 2219 904 2220 908
rect 2214 903 2220 904
rect 2302 908 2308 909
rect 2302 904 2303 908
rect 2307 904 2308 908
rect 2302 903 2308 904
rect 2390 908 2396 909
rect 2390 904 2391 908
rect 2395 904 2396 908
rect 2390 903 2396 904
rect 2478 908 2484 909
rect 2478 904 2479 908
rect 2483 904 2484 908
rect 2478 903 2484 904
rect 2566 908 2572 909
rect 2566 904 2567 908
rect 2571 904 2572 908
rect 2566 903 2572 904
rect 2654 908 2660 909
rect 2654 904 2655 908
rect 2659 904 2660 908
rect 2654 903 2660 904
rect 2742 908 2748 909
rect 2742 904 2743 908
rect 2747 904 2748 908
rect 2742 903 2748 904
rect 2830 908 2836 909
rect 2830 904 2831 908
rect 2835 904 2836 908
rect 3464 906 3466 925
rect 2830 903 2836 904
rect 3462 905 3468 906
rect 1806 900 1812 901
rect 3462 901 3463 905
rect 3467 901 3468 905
rect 3462 900 3468 901
rect 1766 896 1772 897
rect 2126 889 2132 890
rect 1806 888 1812 889
rect 414 885 420 886
rect 110 884 116 885
rect 110 880 111 884
rect 115 880 116 884
rect 414 881 415 885
rect 419 881 420 885
rect 414 880 420 881
rect 558 885 564 886
rect 558 881 559 885
rect 563 881 564 885
rect 558 880 564 881
rect 726 885 732 886
rect 726 881 727 885
rect 731 881 732 885
rect 726 880 732 881
rect 910 885 916 886
rect 910 881 911 885
rect 915 881 916 885
rect 910 880 916 881
rect 1118 885 1124 886
rect 1118 881 1119 885
rect 1123 881 1124 885
rect 1118 880 1124 881
rect 1334 885 1340 886
rect 1334 881 1335 885
rect 1339 881 1340 885
rect 1334 880 1340 881
rect 1558 885 1564 886
rect 1558 881 1559 885
rect 1563 881 1564 885
rect 1558 880 1564 881
rect 1766 884 1772 885
rect 1766 880 1767 884
rect 1771 880 1772 884
rect 1806 884 1807 888
rect 1811 884 1812 888
rect 2126 885 2127 889
rect 2131 885 2132 889
rect 2126 884 2132 885
rect 2214 889 2220 890
rect 2214 885 2215 889
rect 2219 885 2220 889
rect 2214 884 2220 885
rect 2302 889 2308 890
rect 2302 885 2303 889
rect 2307 885 2308 889
rect 2302 884 2308 885
rect 2390 889 2396 890
rect 2390 885 2391 889
rect 2395 885 2396 889
rect 2390 884 2396 885
rect 2478 889 2484 890
rect 2478 885 2479 889
rect 2483 885 2484 889
rect 2478 884 2484 885
rect 2566 889 2572 890
rect 2566 885 2567 889
rect 2571 885 2572 889
rect 2566 884 2572 885
rect 2654 889 2660 890
rect 2654 885 2655 889
rect 2659 885 2660 889
rect 2654 884 2660 885
rect 2742 889 2748 890
rect 2742 885 2743 889
rect 2747 885 2748 889
rect 2742 884 2748 885
rect 2830 889 2836 890
rect 2830 885 2831 889
rect 2835 885 2836 889
rect 2830 884 2836 885
rect 3462 888 3468 889
rect 3462 884 3463 888
rect 3467 884 3468 888
rect 1806 883 1812 884
rect 110 879 116 880
rect 112 859 114 879
rect 416 859 418 880
rect 560 859 562 880
rect 728 859 730 880
rect 912 859 914 880
rect 1120 859 1122 880
rect 1336 859 1338 880
rect 1560 859 1562 880
rect 1766 879 1772 880
rect 1768 859 1770 879
rect 1808 859 1810 883
rect 2128 859 2130 884
rect 2216 859 2218 884
rect 2304 859 2306 884
rect 2392 859 2394 884
rect 2480 859 2482 884
rect 2568 859 2570 884
rect 2656 859 2658 884
rect 2744 859 2746 884
rect 2832 859 2834 884
rect 3462 883 3468 884
rect 3464 859 3466 883
rect 111 858 115 859
rect 111 853 115 854
rect 135 858 139 859
rect 135 853 139 854
rect 231 858 235 859
rect 231 853 235 854
rect 359 858 363 859
rect 359 853 363 854
rect 415 858 419 859
rect 415 853 419 854
rect 487 858 491 859
rect 487 853 491 854
rect 559 858 563 859
rect 559 853 563 854
rect 623 858 627 859
rect 623 853 627 854
rect 727 858 731 859
rect 727 853 731 854
rect 751 858 755 859
rect 751 853 755 854
rect 879 858 883 859
rect 879 853 883 854
rect 911 858 915 859
rect 911 853 915 854
rect 1007 858 1011 859
rect 1007 853 1011 854
rect 1119 858 1123 859
rect 1119 853 1123 854
rect 1135 858 1139 859
rect 1135 853 1139 854
rect 1271 858 1275 859
rect 1271 853 1275 854
rect 1335 858 1339 859
rect 1335 853 1339 854
rect 1559 858 1563 859
rect 1559 853 1563 854
rect 1767 858 1771 859
rect 1767 853 1771 854
rect 1807 858 1811 859
rect 1807 853 1811 854
rect 2127 858 2131 859
rect 2127 853 2131 854
rect 2159 858 2163 859
rect 2159 853 2163 854
rect 2215 858 2219 859
rect 2215 853 2219 854
rect 2247 858 2251 859
rect 2247 853 2251 854
rect 2303 858 2307 859
rect 2303 853 2307 854
rect 2335 858 2339 859
rect 2335 853 2339 854
rect 2391 858 2395 859
rect 2391 853 2395 854
rect 2423 858 2427 859
rect 2423 853 2427 854
rect 2479 858 2483 859
rect 2479 853 2483 854
rect 2527 858 2531 859
rect 2527 853 2531 854
rect 2567 858 2571 859
rect 2567 853 2571 854
rect 2639 858 2643 859
rect 2639 853 2643 854
rect 2655 858 2659 859
rect 2655 853 2659 854
rect 2743 858 2747 859
rect 2743 853 2747 854
rect 2767 858 2771 859
rect 2767 853 2771 854
rect 2831 858 2835 859
rect 2831 853 2835 854
rect 2911 858 2915 859
rect 2911 853 2915 854
rect 3063 858 3067 859
rect 3063 853 3067 854
rect 3223 858 3227 859
rect 3223 853 3227 854
rect 3367 858 3371 859
rect 3367 853 3371 854
rect 3463 858 3467 859
rect 3463 853 3467 854
rect 112 837 114 853
rect 110 836 116 837
rect 136 836 138 853
rect 232 836 234 853
rect 360 836 362 853
rect 488 836 490 853
rect 624 836 626 853
rect 752 836 754 853
rect 880 836 882 853
rect 1008 836 1010 853
rect 1136 836 1138 853
rect 1272 836 1274 853
rect 1768 837 1770 853
rect 1808 837 1810 853
rect 1766 836 1772 837
rect 110 832 111 836
rect 115 832 116 836
rect 110 831 116 832
rect 134 835 140 836
rect 134 831 135 835
rect 139 831 140 835
rect 134 830 140 831
rect 230 835 236 836
rect 230 831 231 835
rect 235 831 236 835
rect 230 830 236 831
rect 358 835 364 836
rect 358 831 359 835
rect 363 831 364 835
rect 358 830 364 831
rect 486 835 492 836
rect 486 831 487 835
rect 491 831 492 835
rect 486 830 492 831
rect 622 835 628 836
rect 622 831 623 835
rect 627 831 628 835
rect 622 830 628 831
rect 750 835 756 836
rect 750 831 751 835
rect 755 831 756 835
rect 750 830 756 831
rect 878 835 884 836
rect 878 831 879 835
rect 883 831 884 835
rect 878 830 884 831
rect 1006 835 1012 836
rect 1006 831 1007 835
rect 1011 831 1012 835
rect 1006 830 1012 831
rect 1134 835 1140 836
rect 1134 831 1135 835
rect 1139 831 1140 835
rect 1134 830 1140 831
rect 1270 835 1276 836
rect 1270 831 1271 835
rect 1275 831 1276 835
rect 1766 832 1767 836
rect 1771 832 1772 836
rect 1766 831 1772 832
rect 1806 836 1812 837
rect 2160 836 2162 853
rect 2248 836 2250 853
rect 2336 836 2338 853
rect 2424 836 2426 853
rect 2528 836 2530 853
rect 2640 836 2642 853
rect 2768 836 2770 853
rect 2912 836 2914 853
rect 3064 836 3066 853
rect 3224 836 3226 853
rect 3368 836 3370 853
rect 3464 837 3466 853
rect 3462 836 3468 837
rect 1806 832 1807 836
rect 1811 832 1812 836
rect 1806 831 1812 832
rect 2158 835 2164 836
rect 2158 831 2159 835
rect 2163 831 2164 835
rect 1270 830 1276 831
rect 2158 830 2164 831
rect 2246 835 2252 836
rect 2246 831 2247 835
rect 2251 831 2252 835
rect 2246 830 2252 831
rect 2334 835 2340 836
rect 2334 831 2335 835
rect 2339 831 2340 835
rect 2334 830 2340 831
rect 2422 835 2428 836
rect 2422 831 2423 835
rect 2427 831 2428 835
rect 2422 830 2428 831
rect 2526 835 2532 836
rect 2526 831 2527 835
rect 2531 831 2532 835
rect 2526 830 2532 831
rect 2638 835 2644 836
rect 2638 831 2639 835
rect 2643 831 2644 835
rect 2638 830 2644 831
rect 2766 835 2772 836
rect 2766 831 2767 835
rect 2771 831 2772 835
rect 2766 830 2772 831
rect 2910 835 2916 836
rect 2910 831 2911 835
rect 2915 831 2916 835
rect 2910 830 2916 831
rect 3062 835 3068 836
rect 3062 831 3063 835
rect 3067 831 3068 835
rect 3062 830 3068 831
rect 3222 835 3228 836
rect 3222 831 3223 835
rect 3227 831 3228 835
rect 3222 830 3228 831
rect 3366 835 3372 836
rect 3366 831 3367 835
rect 3371 831 3372 835
rect 3462 832 3463 836
rect 3467 832 3468 836
rect 3462 831 3468 832
rect 3366 830 3372 831
rect 110 819 116 820
rect 110 815 111 819
rect 115 815 116 819
rect 1766 819 1772 820
rect 110 814 116 815
rect 134 816 140 817
rect 112 791 114 814
rect 134 812 135 816
rect 139 812 140 816
rect 134 811 140 812
rect 230 816 236 817
rect 230 812 231 816
rect 235 812 236 816
rect 230 811 236 812
rect 358 816 364 817
rect 358 812 359 816
rect 363 812 364 816
rect 358 811 364 812
rect 486 816 492 817
rect 486 812 487 816
rect 491 812 492 816
rect 486 811 492 812
rect 622 816 628 817
rect 622 812 623 816
rect 627 812 628 816
rect 622 811 628 812
rect 750 816 756 817
rect 750 812 751 816
rect 755 812 756 816
rect 750 811 756 812
rect 878 816 884 817
rect 878 812 879 816
rect 883 812 884 816
rect 878 811 884 812
rect 1006 816 1012 817
rect 1006 812 1007 816
rect 1011 812 1012 816
rect 1006 811 1012 812
rect 1134 816 1140 817
rect 1134 812 1135 816
rect 1139 812 1140 816
rect 1134 811 1140 812
rect 1270 816 1276 817
rect 1270 812 1271 816
rect 1275 812 1276 816
rect 1766 815 1767 819
rect 1771 815 1772 819
rect 1766 814 1772 815
rect 1806 819 1812 820
rect 1806 815 1807 819
rect 1811 815 1812 819
rect 3462 819 3468 820
rect 1806 814 1812 815
rect 2158 816 2164 817
rect 1270 811 1276 812
rect 136 791 138 811
rect 232 791 234 811
rect 360 791 362 811
rect 488 791 490 811
rect 624 791 626 811
rect 752 791 754 811
rect 880 791 882 811
rect 1008 791 1010 811
rect 1136 791 1138 811
rect 1272 791 1274 811
rect 1768 791 1770 814
rect 1808 791 1810 814
rect 2158 812 2159 816
rect 2163 812 2164 816
rect 2158 811 2164 812
rect 2246 816 2252 817
rect 2246 812 2247 816
rect 2251 812 2252 816
rect 2246 811 2252 812
rect 2334 816 2340 817
rect 2334 812 2335 816
rect 2339 812 2340 816
rect 2334 811 2340 812
rect 2422 816 2428 817
rect 2422 812 2423 816
rect 2427 812 2428 816
rect 2422 811 2428 812
rect 2526 816 2532 817
rect 2526 812 2527 816
rect 2531 812 2532 816
rect 2526 811 2532 812
rect 2638 816 2644 817
rect 2638 812 2639 816
rect 2643 812 2644 816
rect 2638 811 2644 812
rect 2766 816 2772 817
rect 2766 812 2767 816
rect 2771 812 2772 816
rect 2766 811 2772 812
rect 2910 816 2916 817
rect 2910 812 2911 816
rect 2915 812 2916 816
rect 2910 811 2916 812
rect 3062 816 3068 817
rect 3062 812 3063 816
rect 3067 812 3068 816
rect 3062 811 3068 812
rect 3222 816 3228 817
rect 3222 812 3223 816
rect 3227 812 3228 816
rect 3222 811 3228 812
rect 3366 816 3372 817
rect 3366 812 3367 816
rect 3371 812 3372 816
rect 3462 815 3463 819
rect 3467 815 3468 819
rect 3462 814 3468 815
rect 3366 811 3372 812
rect 2160 791 2162 811
rect 2248 791 2250 811
rect 2336 791 2338 811
rect 2424 791 2426 811
rect 2528 791 2530 811
rect 2640 791 2642 811
rect 2768 791 2770 811
rect 2912 791 2914 811
rect 3064 791 3066 811
rect 3224 791 3226 811
rect 3368 791 3370 811
rect 3464 791 3466 814
rect 111 790 115 791
rect 111 785 115 786
rect 135 790 139 791
rect 135 785 139 786
rect 223 790 227 791
rect 223 785 227 786
rect 231 790 235 791
rect 231 785 235 786
rect 343 790 347 791
rect 343 785 347 786
rect 359 790 363 791
rect 359 785 363 786
rect 471 790 475 791
rect 471 785 475 786
rect 487 790 491 791
rect 487 785 491 786
rect 607 790 611 791
rect 607 785 611 786
rect 623 790 627 791
rect 623 785 627 786
rect 743 790 747 791
rect 743 785 747 786
rect 751 790 755 791
rect 751 785 755 786
rect 879 790 883 791
rect 879 785 883 786
rect 887 790 891 791
rect 887 785 891 786
rect 1007 790 1011 791
rect 1007 785 1011 786
rect 1039 790 1043 791
rect 1039 785 1043 786
rect 1135 790 1139 791
rect 1135 785 1139 786
rect 1191 790 1195 791
rect 1191 785 1195 786
rect 1271 790 1275 791
rect 1271 785 1275 786
rect 1351 790 1355 791
rect 1351 785 1355 786
rect 1767 790 1771 791
rect 1767 785 1771 786
rect 1807 790 1811 791
rect 1807 785 1811 786
rect 2063 790 2067 791
rect 2063 785 2067 786
rect 2159 790 2163 791
rect 2159 785 2163 786
rect 2175 790 2179 791
rect 2175 785 2179 786
rect 2247 790 2251 791
rect 2247 785 2251 786
rect 2295 790 2299 791
rect 2295 785 2299 786
rect 2335 790 2339 791
rect 2335 785 2339 786
rect 2423 790 2427 791
rect 2423 785 2427 786
rect 2527 790 2531 791
rect 2527 785 2531 786
rect 2559 790 2563 791
rect 2559 785 2563 786
rect 2639 790 2643 791
rect 2639 785 2643 786
rect 2711 790 2715 791
rect 2711 785 2715 786
rect 2767 790 2771 791
rect 2767 785 2771 786
rect 2871 790 2875 791
rect 2871 785 2875 786
rect 2911 790 2915 791
rect 2911 785 2915 786
rect 3039 790 3043 791
rect 3039 785 3043 786
rect 3063 790 3067 791
rect 3063 785 3067 786
rect 3215 790 3219 791
rect 3215 785 3219 786
rect 3223 790 3227 791
rect 3223 785 3227 786
rect 3367 790 3371 791
rect 3367 785 3371 786
rect 3463 790 3467 791
rect 3463 785 3467 786
rect 112 766 114 785
rect 136 769 138 785
rect 224 769 226 785
rect 344 769 346 785
rect 472 769 474 785
rect 608 769 610 785
rect 744 769 746 785
rect 888 769 890 785
rect 1040 769 1042 785
rect 1192 769 1194 785
rect 1352 769 1354 785
rect 134 768 140 769
rect 110 765 116 766
rect 110 761 111 765
rect 115 761 116 765
rect 134 764 135 768
rect 139 764 140 768
rect 134 763 140 764
rect 222 768 228 769
rect 222 764 223 768
rect 227 764 228 768
rect 222 763 228 764
rect 342 768 348 769
rect 342 764 343 768
rect 347 764 348 768
rect 342 763 348 764
rect 470 768 476 769
rect 470 764 471 768
rect 475 764 476 768
rect 470 763 476 764
rect 606 768 612 769
rect 606 764 607 768
rect 611 764 612 768
rect 606 763 612 764
rect 742 768 748 769
rect 742 764 743 768
rect 747 764 748 768
rect 742 763 748 764
rect 886 768 892 769
rect 886 764 887 768
rect 891 764 892 768
rect 886 763 892 764
rect 1038 768 1044 769
rect 1038 764 1039 768
rect 1043 764 1044 768
rect 1038 763 1044 764
rect 1190 768 1196 769
rect 1190 764 1191 768
rect 1195 764 1196 768
rect 1190 763 1196 764
rect 1350 768 1356 769
rect 1350 764 1351 768
rect 1355 764 1356 768
rect 1768 766 1770 785
rect 1808 766 1810 785
rect 2064 769 2066 785
rect 2176 769 2178 785
rect 2296 769 2298 785
rect 2424 769 2426 785
rect 2560 769 2562 785
rect 2712 769 2714 785
rect 2872 769 2874 785
rect 3040 769 3042 785
rect 3216 769 3218 785
rect 3368 769 3370 785
rect 2062 768 2068 769
rect 1350 763 1356 764
rect 1766 765 1772 766
rect 110 760 116 761
rect 1766 761 1767 765
rect 1771 761 1772 765
rect 1766 760 1772 761
rect 1806 765 1812 766
rect 1806 761 1807 765
rect 1811 761 1812 765
rect 2062 764 2063 768
rect 2067 764 2068 768
rect 2062 763 2068 764
rect 2174 768 2180 769
rect 2174 764 2175 768
rect 2179 764 2180 768
rect 2174 763 2180 764
rect 2294 768 2300 769
rect 2294 764 2295 768
rect 2299 764 2300 768
rect 2294 763 2300 764
rect 2422 768 2428 769
rect 2422 764 2423 768
rect 2427 764 2428 768
rect 2422 763 2428 764
rect 2558 768 2564 769
rect 2558 764 2559 768
rect 2563 764 2564 768
rect 2558 763 2564 764
rect 2710 768 2716 769
rect 2710 764 2711 768
rect 2715 764 2716 768
rect 2710 763 2716 764
rect 2870 768 2876 769
rect 2870 764 2871 768
rect 2875 764 2876 768
rect 2870 763 2876 764
rect 3038 768 3044 769
rect 3038 764 3039 768
rect 3043 764 3044 768
rect 3038 763 3044 764
rect 3214 768 3220 769
rect 3214 764 3215 768
rect 3219 764 3220 768
rect 3214 763 3220 764
rect 3366 768 3372 769
rect 3366 764 3367 768
rect 3371 764 3372 768
rect 3464 766 3466 785
rect 3366 763 3372 764
rect 3462 765 3468 766
rect 1806 760 1812 761
rect 3462 761 3463 765
rect 3467 761 3468 765
rect 3462 760 3468 761
rect 134 749 140 750
rect 110 748 116 749
rect 110 744 111 748
rect 115 744 116 748
rect 134 745 135 749
rect 139 745 140 749
rect 134 744 140 745
rect 222 749 228 750
rect 222 745 223 749
rect 227 745 228 749
rect 222 744 228 745
rect 342 749 348 750
rect 342 745 343 749
rect 347 745 348 749
rect 342 744 348 745
rect 470 749 476 750
rect 470 745 471 749
rect 475 745 476 749
rect 470 744 476 745
rect 606 749 612 750
rect 606 745 607 749
rect 611 745 612 749
rect 606 744 612 745
rect 742 749 748 750
rect 742 745 743 749
rect 747 745 748 749
rect 742 744 748 745
rect 886 749 892 750
rect 886 745 887 749
rect 891 745 892 749
rect 886 744 892 745
rect 1038 749 1044 750
rect 1038 745 1039 749
rect 1043 745 1044 749
rect 1038 744 1044 745
rect 1190 749 1196 750
rect 1190 745 1191 749
rect 1195 745 1196 749
rect 1190 744 1196 745
rect 1350 749 1356 750
rect 2062 749 2068 750
rect 1350 745 1351 749
rect 1355 745 1356 749
rect 1350 744 1356 745
rect 1766 748 1772 749
rect 1766 744 1767 748
rect 1771 744 1772 748
rect 110 743 116 744
rect 112 723 114 743
rect 136 723 138 744
rect 224 723 226 744
rect 344 723 346 744
rect 472 723 474 744
rect 608 723 610 744
rect 744 723 746 744
rect 888 723 890 744
rect 1040 723 1042 744
rect 1192 723 1194 744
rect 1352 723 1354 744
rect 1766 743 1772 744
rect 1806 748 1812 749
rect 1806 744 1807 748
rect 1811 744 1812 748
rect 2062 745 2063 749
rect 2067 745 2068 749
rect 2062 744 2068 745
rect 2174 749 2180 750
rect 2174 745 2175 749
rect 2179 745 2180 749
rect 2174 744 2180 745
rect 2294 749 2300 750
rect 2294 745 2295 749
rect 2299 745 2300 749
rect 2294 744 2300 745
rect 2422 749 2428 750
rect 2422 745 2423 749
rect 2427 745 2428 749
rect 2422 744 2428 745
rect 2558 749 2564 750
rect 2558 745 2559 749
rect 2563 745 2564 749
rect 2558 744 2564 745
rect 2710 749 2716 750
rect 2710 745 2711 749
rect 2715 745 2716 749
rect 2710 744 2716 745
rect 2870 749 2876 750
rect 2870 745 2871 749
rect 2875 745 2876 749
rect 2870 744 2876 745
rect 3038 749 3044 750
rect 3038 745 3039 749
rect 3043 745 3044 749
rect 3038 744 3044 745
rect 3214 749 3220 750
rect 3214 745 3215 749
rect 3219 745 3220 749
rect 3214 744 3220 745
rect 3366 749 3372 750
rect 3366 745 3367 749
rect 3371 745 3372 749
rect 3366 744 3372 745
rect 3462 748 3468 749
rect 3462 744 3463 748
rect 3467 744 3468 748
rect 1806 743 1812 744
rect 1768 723 1770 743
rect 1808 727 1810 743
rect 2064 727 2066 744
rect 2176 727 2178 744
rect 2296 727 2298 744
rect 2424 727 2426 744
rect 2560 727 2562 744
rect 2712 727 2714 744
rect 2872 727 2874 744
rect 3040 727 3042 744
rect 3216 727 3218 744
rect 3368 727 3370 744
rect 3462 743 3468 744
rect 3464 727 3466 743
rect 1807 726 1811 727
rect 111 722 115 723
rect 111 717 115 718
rect 135 722 139 723
rect 135 717 139 718
rect 167 722 171 723
rect 167 717 171 718
rect 223 722 227 723
rect 223 717 227 718
rect 295 722 299 723
rect 295 717 299 718
rect 343 722 347 723
rect 343 717 347 718
rect 431 722 435 723
rect 431 717 435 718
rect 471 722 475 723
rect 471 717 475 718
rect 575 722 579 723
rect 575 717 579 718
rect 607 722 611 723
rect 607 717 611 718
rect 727 722 731 723
rect 727 717 731 718
rect 743 722 747 723
rect 743 717 747 718
rect 879 722 883 723
rect 879 717 883 718
rect 887 722 891 723
rect 887 717 891 718
rect 1031 722 1035 723
rect 1031 717 1035 718
rect 1039 722 1043 723
rect 1039 717 1043 718
rect 1183 722 1187 723
rect 1183 717 1187 718
rect 1191 722 1195 723
rect 1191 717 1195 718
rect 1343 722 1347 723
rect 1343 717 1347 718
rect 1351 722 1355 723
rect 1351 717 1355 718
rect 1503 722 1507 723
rect 1503 717 1507 718
rect 1767 722 1771 723
rect 1807 721 1811 722
rect 1927 726 1931 727
rect 1927 721 1931 722
rect 2063 726 2067 727
rect 2063 721 2067 722
rect 2071 726 2075 727
rect 2071 721 2075 722
rect 2175 726 2179 727
rect 2175 721 2179 722
rect 2231 726 2235 727
rect 2231 721 2235 722
rect 2295 726 2299 727
rect 2295 721 2299 722
rect 2391 726 2395 727
rect 2391 721 2395 722
rect 2423 726 2427 727
rect 2423 721 2427 722
rect 2551 726 2555 727
rect 2551 721 2555 722
rect 2559 726 2563 727
rect 2559 721 2563 722
rect 2703 726 2707 727
rect 2703 721 2707 722
rect 2711 726 2715 727
rect 2711 721 2715 722
rect 2847 726 2851 727
rect 2847 721 2851 722
rect 2871 726 2875 727
rect 2871 721 2875 722
rect 2983 726 2987 727
rect 2983 721 2987 722
rect 3039 726 3043 727
rect 3039 721 3043 722
rect 3119 726 3123 727
rect 3119 721 3123 722
rect 3215 726 3219 727
rect 3215 721 3219 722
rect 3255 726 3259 727
rect 3255 721 3259 722
rect 3367 726 3371 727
rect 3367 721 3371 722
rect 3463 726 3467 727
rect 3463 721 3467 722
rect 1767 717 1771 718
rect 112 701 114 717
rect 110 700 116 701
rect 168 700 170 717
rect 296 700 298 717
rect 432 700 434 717
rect 576 700 578 717
rect 728 700 730 717
rect 880 700 882 717
rect 1032 700 1034 717
rect 1184 700 1186 717
rect 1344 700 1346 717
rect 1504 700 1506 717
rect 1768 701 1770 717
rect 1808 705 1810 721
rect 1806 704 1812 705
rect 1928 704 1930 721
rect 2072 704 2074 721
rect 2232 704 2234 721
rect 2392 704 2394 721
rect 2552 704 2554 721
rect 2704 704 2706 721
rect 2848 704 2850 721
rect 2984 704 2986 721
rect 3120 704 3122 721
rect 3256 704 3258 721
rect 3368 704 3370 721
rect 3464 705 3466 721
rect 3462 704 3468 705
rect 1766 700 1772 701
rect 110 696 111 700
rect 115 696 116 700
rect 110 695 116 696
rect 166 699 172 700
rect 166 695 167 699
rect 171 695 172 699
rect 166 694 172 695
rect 294 699 300 700
rect 294 695 295 699
rect 299 695 300 699
rect 294 694 300 695
rect 430 699 436 700
rect 430 695 431 699
rect 435 695 436 699
rect 430 694 436 695
rect 574 699 580 700
rect 574 695 575 699
rect 579 695 580 699
rect 574 694 580 695
rect 726 699 732 700
rect 726 695 727 699
rect 731 695 732 699
rect 726 694 732 695
rect 878 699 884 700
rect 878 695 879 699
rect 883 695 884 699
rect 878 694 884 695
rect 1030 699 1036 700
rect 1030 695 1031 699
rect 1035 695 1036 699
rect 1030 694 1036 695
rect 1182 699 1188 700
rect 1182 695 1183 699
rect 1187 695 1188 699
rect 1182 694 1188 695
rect 1342 699 1348 700
rect 1342 695 1343 699
rect 1347 695 1348 699
rect 1342 694 1348 695
rect 1502 699 1508 700
rect 1502 695 1503 699
rect 1507 695 1508 699
rect 1766 696 1767 700
rect 1771 696 1772 700
rect 1806 700 1807 704
rect 1811 700 1812 704
rect 1806 699 1812 700
rect 1926 703 1932 704
rect 1926 699 1927 703
rect 1931 699 1932 703
rect 1926 698 1932 699
rect 2070 703 2076 704
rect 2070 699 2071 703
rect 2075 699 2076 703
rect 2070 698 2076 699
rect 2230 703 2236 704
rect 2230 699 2231 703
rect 2235 699 2236 703
rect 2230 698 2236 699
rect 2390 703 2396 704
rect 2390 699 2391 703
rect 2395 699 2396 703
rect 2390 698 2396 699
rect 2550 703 2556 704
rect 2550 699 2551 703
rect 2555 699 2556 703
rect 2550 698 2556 699
rect 2702 703 2708 704
rect 2702 699 2703 703
rect 2707 699 2708 703
rect 2702 698 2708 699
rect 2846 703 2852 704
rect 2846 699 2847 703
rect 2851 699 2852 703
rect 2846 698 2852 699
rect 2982 703 2988 704
rect 2982 699 2983 703
rect 2987 699 2988 703
rect 2982 698 2988 699
rect 3118 703 3124 704
rect 3118 699 3119 703
rect 3123 699 3124 703
rect 3118 698 3124 699
rect 3254 703 3260 704
rect 3254 699 3255 703
rect 3259 699 3260 703
rect 3254 698 3260 699
rect 3366 703 3372 704
rect 3366 699 3367 703
rect 3371 699 3372 703
rect 3462 700 3463 704
rect 3467 700 3468 704
rect 3462 699 3468 700
rect 3366 698 3372 699
rect 1766 695 1772 696
rect 1502 694 1508 695
rect 1806 687 1812 688
rect 110 683 116 684
rect 110 679 111 683
rect 115 679 116 683
rect 1766 683 1772 684
rect 110 678 116 679
rect 166 680 172 681
rect 112 655 114 678
rect 166 676 167 680
rect 171 676 172 680
rect 166 675 172 676
rect 294 680 300 681
rect 294 676 295 680
rect 299 676 300 680
rect 294 675 300 676
rect 430 680 436 681
rect 430 676 431 680
rect 435 676 436 680
rect 430 675 436 676
rect 574 680 580 681
rect 574 676 575 680
rect 579 676 580 680
rect 574 675 580 676
rect 726 680 732 681
rect 726 676 727 680
rect 731 676 732 680
rect 726 675 732 676
rect 878 680 884 681
rect 878 676 879 680
rect 883 676 884 680
rect 878 675 884 676
rect 1030 680 1036 681
rect 1030 676 1031 680
rect 1035 676 1036 680
rect 1030 675 1036 676
rect 1182 680 1188 681
rect 1182 676 1183 680
rect 1187 676 1188 680
rect 1182 675 1188 676
rect 1342 680 1348 681
rect 1342 676 1343 680
rect 1347 676 1348 680
rect 1342 675 1348 676
rect 1502 680 1508 681
rect 1502 676 1503 680
rect 1507 676 1508 680
rect 1766 679 1767 683
rect 1771 679 1772 683
rect 1806 683 1807 687
rect 1811 683 1812 687
rect 3462 687 3468 688
rect 1806 682 1812 683
rect 1926 684 1932 685
rect 1766 678 1772 679
rect 1502 675 1508 676
rect 168 655 170 675
rect 296 655 298 675
rect 432 655 434 675
rect 576 655 578 675
rect 728 655 730 675
rect 880 655 882 675
rect 1032 655 1034 675
rect 1184 655 1186 675
rect 1344 655 1346 675
rect 1504 655 1506 675
rect 1768 655 1770 678
rect 1808 655 1810 682
rect 1926 680 1927 684
rect 1931 680 1932 684
rect 1926 679 1932 680
rect 2070 684 2076 685
rect 2070 680 2071 684
rect 2075 680 2076 684
rect 2070 679 2076 680
rect 2230 684 2236 685
rect 2230 680 2231 684
rect 2235 680 2236 684
rect 2230 679 2236 680
rect 2390 684 2396 685
rect 2390 680 2391 684
rect 2395 680 2396 684
rect 2390 679 2396 680
rect 2550 684 2556 685
rect 2550 680 2551 684
rect 2555 680 2556 684
rect 2550 679 2556 680
rect 2702 684 2708 685
rect 2702 680 2703 684
rect 2707 680 2708 684
rect 2702 679 2708 680
rect 2846 684 2852 685
rect 2846 680 2847 684
rect 2851 680 2852 684
rect 2846 679 2852 680
rect 2982 684 2988 685
rect 2982 680 2983 684
rect 2987 680 2988 684
rect 2982 679 2988 680
rect 3118 684 3124 685
rect 3118 680 3119 684
rect 3123 680 3124 684
rect 3118 679 3124 680
rect 3254 684 3260 685
rect 3254 680 3255 684
rect 3259 680 3260 684
rect 3254 679 3260 680
rect 3366 684 3372 685
rect 3366 680 3367 684
rect 3371 680 3372 684
rect 3462 683 3463 687
rect 3467 683 3468 687
rect 3462 682 3468 683
rect 3366 679 3372 680
rect 1928 655 1930 679
rect 2072 655 2074 679
rect 2232 655 2234 679
rect 2392 655 2394 679
rect 2552 655 2554 679
rect 2704 655 2706 679
rect 2848 655 2850 679
rect 2984 655 2986 679
rect 3120 655 3122 679
rect 3256 655 3258 679
rect 3368 655 3370 679
rect 3464 655 3466 682
rect 111 654 115 655
rect 111 649 115 650
rect 167 654 171 655
rect 167 649 171 650
rect 295 654 299 655
rect 295 649 299 650
rect 431 654 435 655
rect 431 649 435 650
rect 455 654 459 655
rect 455 649 459 650
rect 559 654 563 655
rect 559 649 563 650
rect 575 654 579 655
rect 575 649 579 650
rect 679 654 683 655
rect 679 649 683 650
rect 727 654 731 655
rect 727 649 731 650
rect 799 654 803 655
rect 799 649 803 650
rect 879 654 883 655
rect 879 649 883 650
rect 927 654 931 655
rect 927 649 931 650
rect 1031 654 1035 655
rect 1031 649 1035 650
rect 1055 654 1059 655
rect 1055 649 1059 650
rect 1183 654 1187 655
rect 1183 649 1187 650
rect 1311 654 1315 655
rect 1311 649 1315 650
rect 1343 654 1347 655
rect 1343 649 1347 650
rect 1447 654 1451 655
rect 1447 649 1451 650
rect 1503 654 1507 655
rect 1503 649 1507 650
rect 1583 654 1587 655
rect 1583 649 1587 650
rect 1767 654 1771 655
rect 1767 649 1771 650
rect 1807 654 1811 655
rect 1807 649 1811 650
rect 1831 654 1835 655
rect 1831 649 1835 650
rect 1927 654 1931 655
rect 1927 649 1931 650
rect 1967 654 1971 655
rect 1967 649 1971 650
rect 2071 654 2075 655
rect 2071 649 2075 650
rect 2135 654 2139 655
rect 2135 649 2139 650
rect 2231 654 2235 655
rect 2231 649 2235 650
rect 2311 654 2315 655
rect 2311 649 2315 650
rect 2391 654 2395 655
rect 2391 649 2395 650
rect 2487 654 2491 655
rect 2487 649 2491 650
rect 2551 654 2555 655
rect 2551 649 2555 650
rect 2655 654 2659 655
rect 2655 649 2659 650
rect 2703 654 2707 655
rect 2703 649 2707 650
rect 2815 654 2819 655
rect 2815 649 2819 650
rect 2847 654 2851 655
rect 2847 649 2851 650
rect 2959 654 2963 655
rect 2959 649 2963 650
rect 2983 654 2987 655
rect 2983 649 2987 650
rect 3103 654 3107 655
rect 3103 649 3107 650
rect 3119 654 3123 655
rect 3119 649 3123 650
rect 3247 654 3251 655
rect 3247 649 3251 650
rect 3255 654 3259 655
rect 3255 649 3259 650
rect 3367 654 3371 655
rect 3367 649 3371 650
rect 3463 654 3467 655
rect 3463 649 3467 650
rect 112 630 114 649
rect 456 633 458 649
rect 560 633 562 649
rect 680 633 682 649
rect 800 633 802 649
rect 928 633 930 649
rect 1056 633 1058 649
rect 1184 633 1186 649
rect 1312 633 1314 649
rect 1448 633 1450 649
rect 1584 633 1586 649
rect 454 632 460 633
rect 110 629 116 630
rect 110 625 111 629
rect 115 625 116 629
rect 454 628 455 632
rect 459 628 460 632
rect 454 627 460 628
rect 558 632 564 633
rect 558 628 559 632
rect 563 628 564 632
rect 558 627 564 628
rect 678 632 684 633
rect 678 628 679 632
rect 683 628 684 632
rect 678 627 684 628
rect 798 632 804 633
rect 798 628 799 632
rect 803 628 804 632
rect 798 627 804 628
rect 926 632 932 633
rect 926 628 927 632
rect 931 628 932 632
rect 926 627 932 628
rect 1054 632 1060 633
rect 1054 628 1055 632
rect 1059 628 1060 632
rect 1054 627 1060 628
rect 1182 632 1188 633
rect 1182 628 1183 632
rect 1187 628 1188 632
rect 1182 627 1188 628
rect 1310 632 1316 633
rect 1310 628 1311 632
rect 1315 628 1316 632
rect 1310 627 1316 628
rect 1446 632 1452 633
rect 1446 628 1447 632
rect 1451 628 1452 632
rect 1446 627 1452 628
rect 1582 632 1588 633
rect 1582 628 1583 632
rect 1587 628 1588 632
rect 1768 630 1770 649
rect 1808 630 1810 649
rect 1832 633 1834 649
rect 1968 633 1970 649
rect 2136 633 2138 649
rect 2312 633 2314 649
rect 2488 633 2490 649
rect 2656 633 2658 649
rect 2816 633 2818 649
rect 2960 633 2962 649
rect 3104 633 3106 649
rect 3248 633 3250 649
rect 3368 633 3370 649
rect 1830 632 1836 633
rect 1582 627 1588 628
rect 1766 629 1772 630
rect 110 624 116 625
rect 1766 625 1767 629
rect 1771 625 1772 629
rect 1766 624 1772 625
rect 1806 629 1812 630
rect 1806 625 1807 629
rect 1811 625 1812 629
rect 1830 628 1831 632
rect 1835 628 1836 632
rect 1830 627 1836 628
rect 1966 632 1972 633
rect 1966 628 1967 632
rect 1971 628 1972 632
rect 1966 627 1972 628
rect 2134 632 2140 633
rect 2134 628 2135 632
rect 2139 628 2140 632
rect 2134 627 2140 628
rect 2310 632 2316 633
rect 2310 628 2311 632
rect 2315 628 2316 632
rect 2310 627 2316 628
rect 2486 632 2492 633
rect 2486 628 2487 632
rect 2491 628 2492 632
rect 2486 627 2492 628
rect 2654 632 2660 633
rect 2654 628 2655 632
rect 2659 628 2660 632
rect 2654 627 2660 628
rect 2814 632 2820 633
rect 2814 628 2815 632
rect 2819 628 2820 632
rect 2814 627 2820 628
rect 2958 632 2964 633
rect 2958 628 2959 632
rect 2963 628 2964 632
rect 2958 627 2964 628
rect 3102 632 3108 633
rect 3102 628 3103 632
rect 3107 628 3108 632
rect 3102 627 3108 628
rect 3246 632 3252 633
rect 3246 628 3247 632
rect 3251 628 3252 632
rect 3246 627 3252 628
rect 3366 632 3372 633
rect 3366 628 3367 632
rect 3371 628 3372 632
rect 3464 630 3466 649
rect 3366 627 3372 628
rect 3462 629 3468 630
rect 1806 624 1812 625
rect 3462 625 3463 629
rect 3467 625 3468 629
rect 3462 624 3468 625
rect 454 613 460 614
rect 110 612 116 613
rect 110 608 111 612
rect 115 608 116 612
rect 454 609 455 613
rect 459 609 460 613
rect 454 608 460 609
rect 558 613 564 614
rect 558 609 559 613
rect 563 609 564 613
rect 558 608 564 609
rect 678 613 684 614
rect 678 609 679 613
rect 683 609 684 613
rect 678 608 684 609
rect 798 613 804 614
rect 798 609 799 613
rect 803 609 804 613
rect 798 608 804 609
rect 926 613 932 614
rect 926 609 927 613
rect 931 609 932 613
rect 926 608 932 609
rect 1054 613 1060 614
rect 1054 609 1055 613
rect 1059 609 1060 613
rect 1054 608 1060 609
rect 1182 613 1188 614
rect 1182 609 1183 613
rect 1187 609 1188 613
rect 1182 608 1188 609
rect 1310 613 1316 614
rect 1310 609 1311 613
rect 1315 609 1316 613
rect 1310 608 1316 609
rect 1446 613 1452 614
rect 1446 609 1447 613
rect 1451 609 1452 613
rect 1446 608 1452 609
rect 1582 613 1588 614
rect 1830 613 1836 614
rect 1582 609 1583 613
rect 1587 609 1588 613
rect 1582 608 1588 609
rect 1766 612 1772 613
rect 1766 608 1767 612
rect 1771 608 1772 612
rect 110 607 116 608
rect 112 583 114 607
rect 456 583 458 608
rect 560 583 562 608
rect 680 583 682 608
rect 800 583 802 608
rect 928 583 930 608
rect 1056 583 1058 608
rect 1184 583 1186 608
rect 1312 583 1314 608
rect 1448 583 1450 608
rect 1584 583 1586 608
rect 1766 607 1772 608
rect 1806 612 1812 613
rect 1806 608 1807 612
rect 1811 608 1812 612
rect 1830 609 1831 613
rect 1835 609 1836 613
rect 1830 608 1836 609
rect 1966 613 1972 614
rect 1966 609 1967 613
rect 1971 609 1972 613
rect 1966 608 1972 609
rect 2134 613 2140 614
rect 2134 609 2135 613
rect 2139 609 2140 613
rect 2134 608 2140 609
rect 2310 613 2316 614
rect 2310 609 2311 613
rect 2315 609 2316 613
rect 2310 608 2316 609
rect 2486 613 2492 614
rect 2486 609 2487 613
rect 2491 609 2492 613
rect 2486 608 2492 609
rect 2654 613 2660 614
rect 2654 609 2655 613
rect 2659 609 2660 613
rect 2654 608 2660 609
rect 2814 613 2820 614
rect 2814 609 2815 613
rect 2819 609 2820 613
rect 2814 608 2820 609
rect 2958 613 2964 614
rect 2958 609 2959 613
rect 2963 609 2964 613
rect 2958 608 2964 609
rect 3102 613 3108 614
rect 3102 609 3103 613
rect 3107 609 3108 613
rect 3102 608 3108 609
rect 3246 613 3252 614
rect 3246 609 3247 613
rect 3251 609 3252 613
rect 3246 608 3252 609
rect 3366 613 3372 614
rect 3366 609 3367 613
rect 3371 609 3372 613
rect 3366 608 3372 609
rect 3462 612 3468 613
rect 3462 608 3463 612
rect 3467 608 3468 612
rect 1806 607 1812 608
rect 1768 583 1770 607
rect 1808 591 1810 607
rect 1832 591 1834 608
rect 1968 591 1970 608
rect 2136 591 2138 608
rect 2312 591 2314 608
rect 2488 591 2490 608
rect 2656 591 2658 608
rect 2816 591 2818 608
rect 2960 591 2962 608
rect 3104 591 3106 608
rect 3248 591 3250 608
rect 3368 591 3370 608
rect 3462 607 3468 608
rect 3464 591 3466 607
rect 1807 590 1811 591
rect 1807 585 1811 586
rect 1831 590 1835 591
rect 1831 585 1835 586
rect 1967 590 1971 591
rect 1967 585 1971 586
rect 2127 590 2131 591
rect 2127 585 2131 586
rect 2135 590 2139 591
rect 2135 585 2139 586
rect 2287 590 2291 591
rect 2287 585 2291 586
rect 2311 590 2315 591
rect 2311 585 2315 586
rect 2455 590 2459 591
rect 2455 585 2459 586
rect 2487 590 2491 591
rect 2487 585 2491 586
rect 2623 590 2627 591
rect 2623 585 2627 586
rect 2655 590 2659 591
rect 2655 585 2659 586
rect 2799 590 2803 591
rect 2799 585 2803 586
rect 2815 590 2819 591
rect 2815 585 2819 586
rect 2959 590 2963 591
rect 2959 585 2963 586
rect 2983 590 2987 591
rect 2983 585 2987 586
rect 3103 590 3107 591
rect 3103 585 3107 586
rect 3167 590 3171 591
rect 3167 585 3171 586
rect 3247 590 3251 591
rect 3247 585 3251 586
rect 3359 590 3363 591
rect 3359 585 3363 586
rect 3367 590 3371 591
rect 3367 585 3371 586
rect 3463 590 3467 591
rect 3463 585 3467 586
rect 111 582 115 583
rect 111 577 115 578
rect 455 582 459 583
rect 455 577 459 578
rect 559 582 563 583
rect 559 577 563 578
rect 599 582 603 583
rect 599 577 603 578
rect 679 582 683 583
rect 679 577 683 578
rect 703 582 707 583
rect 703 577 707 578
rect 799 582 803 583
rect 799 577 803 578
rect 815 582 819 583
rect 815 577 819 578
rect 927 582 931 583
rect 927 577 931 578
rect 1039 582 1043 583
rect 1039 577 1043 578
rect 1055 582 1059 583
rect 1055 577 1059 578
rect 1151 582 1155 583
rect 1151 577 1155 578
rect 1183 582 1187 583
rect 1183 577 1187 578
rect 1255 582 1259 583
rect 1255 577 1259 578
rect 1311 582 1315 583
rect 1311 577 1315 578
rect 1359 582 1363 583
rect 1359 577 1363 578
rect 1447 582 1451 583
rect 1447 577 1451 578
rect 1471 582 1475 583
rect 1471 577 1475 578
rect 1583 582 1587 583
rect 1583 577 1587 578
rect 1671 582 1675 583
rect 1671 577 1675 578
rect 1767 582 1771 583
rect 1767 577 1771 578
rect 112 561 114 577
rect 110 560 116 561
rect 600 560 602 577
rect 704 560 706 577
rect 816 560 818 577
rect 928 560 930 577
rect 1040 560 1042 577
rect 1152 560 1154 577
rect 1256 560 1258 577
rect 1360 560 1362 577
rect 1472 560 1474 577
rect 1584 560 1586 577
rect 1672 560 1674 577
rect 1768 561 1770 577
rect 1808 569 1810 585
rect 1806 568 1812 569
rect 1832 568 1834 585
rect 1968 568 1970 585
rect 2128 568 2130 585
rect 2288 568 2290 585
rect 2456 568 2458 585
rect 2624 568 2626 585
rect 2800 568 2802 585
rect 2984 568 2986 585
rect 3168 568 3170 585
rect 3360 568 3362 585
rect 3464 569 3466 585
rect 3462 568 3468 569
rect 1806 564 1807 568
rect 1811 564 1812 568
rect 1806 563 1812 564
rect 1830 567 1836 568
rect 1830 563 1831 567
rect 1835 563 1836 567
rect 1830 562 1836 563
rect 1966 567 1972 568
rect 1966 563 1967 567
rect 1971 563 1972 567
rect 1966 562 1972 563
rect 2126 567 2132 568
rect 2126 563 2127 567
rect 2131 563 2132 567
rect 2126 562 2132 563
rect 2286 567 2292 568
rect 2286 563 2287 567
rect 2291 563 2292 567
rect 2286 562 2292 563
rect 2454 567 2460 568
rect 2454 563 2455 567
rect 2459 563 2460 567
rect 2454 562 2460 563
rect 2622 567 2628 568
rect 2622 563 2623 567
rect 2627 563 2628 567
rect 2622 562 2628 563
rect 2798 567 2804 568
rect 2798 563 2799 567
rect 2803 563 2804 567
rect 2798 562 2804 563
rect 2982 567 2988 568
rect 2982 563 2983 567
rect 2987 563 2988 567
rect 2982 562 2988 563
rect 3166 567 3172 568
rect 3166 563 3167 567
rect 3171 563 3172 567
rect 3166 562 3172 563
rect 3358 567 3364 568
rect 3358 563 3359 567
rect 3363 563 3364 567
rect 3462 564 3463 568
rect 3467 564 3468 568
rect 3462 563 3468 564
rect 3358 562 3364 563
rect 1766 560 1772 561
rect 110 556 111 560
rect 115 556 116 560
rect 110 555 116 556
rect 598 559 604 560
rect 598 555 599 559
rect 603 555 604 559
rect 598 554 604 555
rect 702 559 708 560
rect 702 555 703 559
rect 707 555 708 559
rect 702 554 708 555
rect 814 559 820 560
rect 814 555 815 559
rect 819 555 820 559
rect 814 554 820 555
rect 926 559 932 560
rect 926 555 927 559
rect 931 555 932 559
rect 926 554 932 555
rect 1038 559 1044 560
rect 1038 555 1039 559
rect 1043 555 1044 559
rect 1038 554 1044 555
rect 1150 559 1156 560
rect 1150 555 1151 559
rect 1155 555 1156 559
rect 1150 554 1156 555
rect 1254 559 1260 560
rect 1254 555 1255 559
rect 1259 555 1260 559
rect 1254 554 1260 555
rect 1358 559 1364 560
rect 1358 555 1359 559
rect 1363 555 1364 559
rect 1358 554 1364 555
rect 1470 559 1476 560
rect 1470 555 1471 559
rect 1475 555 1476 559
rect 1470 554 1476 555
rect 1582 559 1588 560
rect 1582 555 1583 559
rect 1587 555 1588 559
rect 1582 554 1588 555
rect 1670 559 1676 560
rect 1670 555 1671 559
rect 1675 555 1676 559
rect 1766 556 1767 560
rect 1771 556 1772 560
rect 1766 555 1772 556
rect 1670 554 1676 555
rect 1806 551 1812 552
rect 1806 547 1807 551
rect 1811 547 1812 551
rect 3462 551 3468 552
rect 1806 546 1812 547
rect 1830 548 1836 549
rect 110 543 116 544
rect 110 539 111 543
rect 115 539 116 543
rect 1766 543 1772 544
rect 110 538 116 539
rect 598 540 604 541
rect 112 519 114 538
rect 598 536 599 540
rect 603 536 604 540
rect 598 535 604 536
rect 702 540 708 541
rect 702 536 703 540
rect 707 536 708 540
rect 702 535 708 536
rect 814 540 820 541
rect 814 536 815 540
rect 819 536 820 540
rect 814 535 820 536
rect 926 540 932 541
rect 926 536 927 540
rect 931 536 932 540
rect 926 535 932 536
rect 1038 540 1044 541
rect 1038 536 1039 540
rect 1043 536 1044 540
rect 1038 535 1044 536
rect 1150 540 1156 541
rect 1150 536 1151 540
rect 1155 536 1156 540
rect 1150 535 1156 536
rect 1254 540 1260 541
rect 1254 536 1255 540
rect 1259 536 1260 540
rect 1254 535 1260 536
rect 1358 540 1364 541
rect 1358 536 1359 540
rect 1363 536 1364 540
rect 1358 535 1364 536
rect 1470 540 1476 541
rect 1470 536 1471 540
rect 1475 536 1476 540
rect 1470 535 1476 536
rect 1582 540 1588 541
rect 1582 536 1583 540
rect 1587 536 1588 540
rect 1582 535 1588 536
rect 1670 540 1676 541
rect 1670 536 1671 540
rect 1675 536 1676 540
rect 1766 539 1767 543
rect 1771 539 1772 543
rect 1766 538 1772 539
rect 1670 535 1676 536
rect 600 519 602 535
rect 704 519 706 535
rect 816 519 818 535
rect 928 519 930 535
rect 1040 519 1042 535
rect 1152 519 1154 535
rect 1256 519 1258 535
rect 1360 519 1362 535
rect 1472 519 1474 535
rect 1584 519 1586 535
rect 1672 519 1674 535
rect 1768 519 1770 538
rect 111 518 115 519
rect 111 513 115 514
rect 303 518 307 519
rect 303 513 307 514
rect 431 518 435 519
rect 431 513 435 514
rect 567 518 571 519
rect 567 513 571 514
rect 599 518 603 519
rect 599 513 603 514
rect 703 518 707 519
rect 703 513 707 514
rect 815 518 819 519
rect 815 513 819 514
rect 847 518 851 519
rect 847 513 851 514
rect 927 518 931 519
rect 927 513 931 514
rect 983 518 987 519
rect 983 513 987 514
rect 1039 518 1043 519
rect 1039 513 1043 514
rect 1111 518 1115 519
rect 1111 513 1115 514
rect 1151 518 1155 519
rect 1151 513 1155 514
rect 1231 518 1235 519
rect 1231 513 1235 514
rect 1255 518 1259 519
rect 1255 513 1259 514
rect 1351 518 1355 519
rect 1351 513 1355 514
rect 1359 518 1363 519
rect 1359 513 1363 514
rect 1463 518 1467 519
rect 1463 513 1467 514
rect 1471 518 1475 519
rect 1471 513 1475 514
rect 1575 518 1579 519
rect 1575 513 1579 514
rect 1583 518 1587 519
rect 1583 513 1587 514
rect 1671 518 1675 519
rect 1671 513 1675 514
rect 1767 518 1771 519
rect 1767 513 1771 514
rect 112 494 114 513
rect 304 497 306 513
rect 432 497 434 513
rect 568 497 570 513
rect 704 497 706 513
rect 848 497 850 513
rect 984 497 986 513
rect 1112 497 1114 513
rect 1232 497 1234 513
rect 1352 497 1354 513
rect 1464 497 1466 513
rect 1576 497 1578 513
rect 1672 497 1674 513
rect 302 496 308 497
rect 110 493 116 494
rect 110 489 111 493
rect 115 489 116 493
rect 302 492 303 496
rect 307 492 308 496
rect 302 491 308 492
rect 430 496 436 497
rect 430 492 431 496
rect 435 492 436 496
rect 430 491 436 492
rect 566 496 572 497
rect 566 492 567 496
rect 571 492 572 496
rect 566 491 572 492
rect 702 496 708 497
rect 702 492 703 496
rect 707 492 708 496
rect 702 491 708 492
rect 846 496 852 497
rect 846 492 847 496
rect 851 492 852 496
rect 846 491 852 492
rect 982 496 988 497
rect 982 492 983 496
rect 987 492 988 496
rect 982 491 988 492
rect 1110 496 1116 497
rect 1110 492 1111 496
rect 1115 492 1116 496
rect 1110 491 1116 492
rect 1230 496 1236 497
rect 1230 492 1231 496
rect 1235 492 1236 496
rect 1230 491 1236 492
rect 1350 496 1356 497
rect 1350 492 1351 496
rect 1355 492 1356 496
rect 1350 491 1356 492
rect 1462 496 1468 497
rect 1462 492 1463 496
rect 1467 492 1468 496
rect 1462 491 1468 492
rect 1574 496 1580 497
rect 1574 492 1575 496
rect 1579 492 1580 496
rect 1574 491 1580 492
rect 1670 496 1676 497
rect 1670 492 1671 496
rect 1675 492 1676 496
rect 1768 494 1770 513
rect 1808 511 1810 546
rect 1830 544 1831 548
rect 1835 544 1836 548
rect 1830 543 1836 544
rect 1966 548 1972 549
rect 1966 544 1967 548
rect 1971 544 1972 548
rect 1966 543 1972 544
rect 2126 548 2132 549
rect 2126 544 2127 548
rect 2131 544 2132 548
rect 2126 543 2132 544
rect 2286 548 2292 549
rect 2286 544 2287 548
rect 2291 544 2292 548
rect 2286 543 2292 544
rect 2454 548 2460 549
rect 2454 544 2455 548
rect 2459 544 2460 548
rect 2454 543 2460 544
rect 2622 548 2628 549
rect 2622 544 2623 548
rect 2627 544 2628 548
rect 2622 543 2628 544
rect 2798 548 2804 549
rect 2798 544 2799 548
rect 2803 544 2804 548
rect 2798 543 2804 544
rect 2982 548 2988 549
rect 2982 544 2983 548
rect 2987 544 2988 548
rect 2982 543 2988 544
rect 3166 548 3172 549
rect 3166 544 3167 548
rect 3171 544 3172 548
rect 3166 543 3172 544
rect 3358 548 3364 549
rect 3358 544 3359 548
rect 3363 544 3364 548
rect 3462 547 3463 551
rect 3467 547 3468 551
rect 3462 546 3468 547
rect 3358 543 3364 544
rect 1832 511 1834 543
rect 1968 511 1970 543
rect 2128 511 2130 543
rect 2288 511 2290 543
rect 2456 511 2458 543
rect 2624 511 2626 543
rect 2800 511 2802 543
rect 2984 511 2986 543
rect 3168 511 3170 543
rect 3360 511 3362 543
rect 3464 511 3466 546
rect 1807 510 1811 511
rect 1807 505 1811 506
rect 1831 510 1835 511
rect 1831 505 1835 506
rect 1967 510 1971 511
rect 1967 505 1971 506
rect 2127 510 2131 511
rect 2127 505 2131 506
rect 2287 510 2291 511
rect 2287 505 2291 506
rect 2295 510 2299 511
rect 2295 505 2299 506
rect 2455 510 2459 511
rect 2455 505 2459 506
rect 2479 510 2483 511
rect 2479 505 2483 506
rect 2623 510 2627 511
rect 2623 505 2627 506
rect 2679 510 2683 511
rect 2679 505 2683 506
rect 2799 510 2803 511
rect 2799 505 2803 506
rect 2887 510 2891 511
rect 2887 505 2891 506
rect 2983 510 2987 511
rect 2983 505 2987 506
rect 3111 510 3115 511
rect 3111 505 3115 506
rect 3167 510 3171 511
rect 3167 505 3171 506
rect 3335 510 3339 511
rect 3335 505 3339 506
rect 3359 510 3363 511
rect 3359 505 3363 506
rect 3463 510 3467 511
rect 3463 505 3467 506
rect 1670 491 1676 492
rect 1766 493 1772 494
rect 110 488 116 489
rect 1766 489 1767 493
rect 1771 489 1772 493
rect 1766 488 1772 489
rect 1808 486 1810 505
rect 1832 489 1834 505
rect 1968 489 1970 505
rect 2128 489 2130 505
rect 2296 489 2298 505
rect 2480 489 2482 505
rect 2680 489 2682 505
rect 2888 489 2890 505
rect 3112 489 3114 505
rect 3336 489 3338 505
rect 1830 488 1836 489
rect 1806 485 1812 486
rect 1806 481 1807 485
rect 1811 481 1812 485
rect 1830 484 1831 488
rect 1835 484 1836 488
rect 1830 483 1836 484
rect 1966 488 1972 489
rect 1966 484 1967 488
rect 1971 484 1972 488
rect 1966 483 1972 484
rect 2126 488 2132 489
rect 2126 484 2127 488
rect 2131 484 2132 488
rect 2126 483 2132 484
rect 2294 488 2300 489
rect 2294 484 2295 488
rect 2299 484 2300 488
rect 2294 483 2300 484
rect 2478 488 2484 489
rect 2478 484 2479 488
rect 2483 484 2484 488
rect 2478 483 2484 484
rect 2678 488 2684 489
rect 2678 484 2679 488
rect 2683 484 2684 488
rect 2678 483 2684 484
rect 2886 488 2892 489
rect 2886 484 2887 488
rect 2891 484 2892 488
rect 2886 483 2892 484
rect 3110 488 3116 489
rect 3110 484 3111 488
rect 3115 484 3116 488
rect 3110 483 3116 484
rect 3334 488 3340 489
rect 3334 484 3335 488
rect 3339 484 3340 488
rect 3464 486 3466 505
rect 3334 483 3340 484
rect 3462 485 3468 486
rect 1806 480 1812 481
rect 3462 481 3463 485
rect 3467 481 3468 485
rect 3462 480 3468 481
rect 302 477 308 478
rect 110 476 116 477
rect 110 472 111 476
rect 115 472 116 476
rect 302 473 303 477
rect 307 473 308 477
rect 302 472 308 473
rect 430 477 436 478
rect 430 473 431 477
rect 435 473 436 477
rect 430 472 436 473
rect 566 477 572 478
rect 566 473 567 477
rect 571 473 572 477
rect 566 472 572 473
rect 702 477 708 478
rect 702 473 703 477
rect 707 473 708 477
rect 702 472 708 473
rect 846 477 852 478
rect 846 473 847 477
rect 851 473 852 477
rect 846 472 852 473
rect 982 477 988 478
rect 982 473 983 477
rect 987 473 988 477
rect 982 472 988 473
rect 1110 477 1116 478
rect 1110 473 1111 477
rect 1115 473 1116 477
rect 1110 472 1116 473
rect 1230 477 1236 478
rect 1230 473 1231 477
rect 1235 473 1236 477
rect 1230 472 1236 473
rect 1350 477 1356 478
rect 1350 473 1351 477
rect 1355 473 1356 477
rect 1350 472 1356 473
rect 1462 477 1468 478
rect 1462 473 1463 477
rect 1467 473 1468 477
rect 1462 472 1468 473
rect 1574 477 1580 478
rect 1574 473 1575 477
rect 1579 473 1580 477
rect 1574 472 1580 473
rect 1670 477 1676 478
rect 1670 473 1671 477
rect 1675 473 1676 477
rect 1670 472 1676 473
rect 1766 476 1772 477
rect 1766 472 1767 476
rect 1771 472 1772 476
rect 110 471 116 472
rect 112 447 114 471
rect 304 447 306 472
rect 432 447 434 472
rect 568 447 570 472
rect 704 447 706 472
rect 848 447 850 472
rect 984 447 986 472
rect 1112 447 1114 472
rect 1232 447 1234 472
rect 1352 447 1354 472
rect 1464 447 1466 472
rect 1576 447 1578 472
rect 1672 447 1674 472
rect 1766 471 1772 472
rect 1768 447 1770 471
rect 1830 469 1836 470
rect 1806 468 1812 469
rect 1806 464 1807 468
rect 1811 464 1812 468
rect 1830 465 1831 469
rect 1835 465 1836 469
rect 1830 464 1836 465
rect 1966 469 1972 470
rect 1966 465 1967 469
rect 1971 465 1972 469
rect 1966 464 1972 465
rect 2126 469 2132 470
rect 2126 465 2127 469
rect 2131 465 2132 469
rect 2126 464 2132 465
rect 2294 469 2300 470
rect 2294 465 2295 469
rect 2299 465 2300 469
rect 2294 464 2300 465
rect 2478 469 2484 470
rect 2478 465 2479 469
rect 2483 465 2484 469
rect 2478 464 2484 465
rect 2678 469 2684 470
rect 2678 465 2679 469
rect 2683 465 2684 469
rect 2678 464 2684 465
rect 2886 469 2892 470
rect 2886 465 2887 469
rect 2891 465 2892 469
rect 2886 464 2892 465
rect 3110 469 3116 470
rect 3110 465 3111 469
rect 3115 465 3116 469
rect 3110 464 3116 465
rect 3334 469 3340 470
rect 3334 465 3335 469
rect 3339 465 3340 469
rect 3334 464 3340 465
rect 3462 468 3468 469
rect 3462 464 3463 468
rect 3467 464 3468 468
rect 1806 463 1812 464
rect 1808 447 1810 463
rect 1832 447 1834 464
rect 1968 447 1970 464
rect 2128 447 2130 464
rect 2296 447 2298 464
rect 2480 447 2482 464
rect 2680 447 2682 464
rect 2888 447 2890 464
rect 3112 447 3114 464
rect 3336 447 3338 464
rect 3462 463 3468 464
rect 3464 447 3466 463
rect 111 446 115 447
rect 111 441 115 442
rect 135 446 139 447
rect 135 441 139 442
rect 255 446 259 447
rect 255 441 259 442
rect 303 446 307 447
rect 303 441 307 442
rect 415 446 419 447
rect 415 441 419 442
rect 431 446 435 447
rect 431 441 435 442
rect 567 446 571 447
rect 567 441 571 442
rect 583 446 587 447
rect 583 441 587 442
rect 703 446 707 447
rect 703 441 707 442
rect 743 446 747 447
rect 743 441 747 442
rect 847 446 851 447
rect 847 441 851 442
rect 903 446 907 447
rect 903 441 907 442
rect 983 446 987 447
rect 983 441 987 442
rect 1047 446 1051 447
rect 1047 441 1051 442
rect 1111 446 1115 447
rect 1111 441 1115 442
rect 1183 446 1187 447
rect 1183 441 1187 442
rect 1231 446 1235 447
rect 1231 441 1235 442
rect 1311 446 1315 447
rect 1311 441 1315 442
rect 1351 446 1355 447
rect 1351 441 1355 442
rect 1439 446 1443 447
rect 1439 441 1443 442
rect 1463 446 1467 447
rect 1463 441 1467 442
rect 1567 446 1571 447
rect 1567 441 1571 442
rect 1575 446 1579 447
rect 1575 441 1579 442
rect 1671 446 1675 447
rect 1671 441 1675 442
rect 1767 446 1771 447
rect 1767 441 1771 442
rect 1807 446 1811 447
rect 1807 441 1811 442
rect 1831 446 1835 447
rect 1831 441 1835 442
rect 1959 446 1963 447
rect 1959 441 1963 442
rect 1967 446 1971 447
rect 1967 441 1971 442
rect 2111 446 2115 447
rect 2111 441 2115 442
rect 2127 446 2131 447
rect 2127 441 2131 442
rect 2271 446 2275 447
rect 2271 441 2275 442
rect 2295 446 2299 447
rect 2295 441 2299 442
rect 2455 446 2459 447
rect 2455 441 2459 442
rect 2479 446 2483 447
rect 2479 441 2483 442
rect 2655 446 2659 447
rect 2655 441 2659 442
rect 2679 446 2683 447
rect 2679 441 2683 442
rect 2871 446 2875 447
rect 2871 441 2875 442
rect 2887 446 2891 447
rect 2887 441 2891 442
rect 3103 446 3107 447
rect 3103 441 3107 442
rect 3111 446 3115 447
rect 3111 441 3115 442
rect 3335 446 3339 447
rect 3335 441 3339 442
rect 3463 446 3467 447
rect 3463 441 3467 442
rect 112 425 114 441
rect 110 424 116 425
rect 136 424 138 441
rect 256 424 258 441
rect 416 424 418 441
rect 584 424 586 441
rect 744 424 746 441
rect 904 424 906 441
rect 1048 424 1050 441
rect 1184 424 1186 441
rect 1312 424 1314 441
rect 1440 424 1442 441
rect 1568 424 1570 441
rect 1672 424 1674 441
rect 1768 425 1770 441
rect 1808 425 1810 441
rect 1766 424 1772 425
rect 110 420 111 424
rect 115 420 116 424
rect 110 419 116 420
rect 134 423 140 424
rect 134 419 135 423
rect 139 419 140 423
rect 134 418 140 419
rect 254 423 260 424
rect 254 419 255 423
rect 259 419 260 423
rect 254 418 260 419
rect 414 423 420 424
rect 414 419 415 423
rect 419 419 420 423
rect 414 418 420 419
rect 582 423 588 424
rect 582 419 583 423
rect 587 419 588 423
rect 582 418 588 419
rect 742 423 748 424
rect 742 419 743 423
rect 747 419 748 423
rect 742 418 748 419
rect 902 423 908 424
rect 902 419 903 423
rect 907 419 908 423
rect 902 418 908 419
rect 1046 423 1052 424
rect 1046 419 1047 423
rect 1051 419 1052 423
rect 1046 418 1052 419
rect 1182 423 1188 424
rect 1182 419 1183 423
rect 1187 419 1188 423
rect 1182 418 1188 419
rect 1310 423 1316 424
rect 1310 419 1311 423
rect 1315 419 1316 423
rect 1310 418 1316 419
rect 1438 423 1444 424
rect 1438 419 1439 423
rect 1443 419 1444 423
rect 1438 418 1444 419
rect 1566 423 1572 424
rect 1566 419 1567 423
rect 1571 419 1572 423
rect 1566 418 1572 419
rect 1670 423 1676 424
rect 1670 419 1671 423
rect 1675 419 1676 423
rect 1766 420 1767 424
rect 1771 420 1772 424
rect 1766 419 1772 420
rect 1806 424 1812 425
rect 1832 424 1834 441
rect 1960 424 1962 441
rect 2112 424 2114 441
rect 2272 424 2274 441
rect 2456 424 2458 441
rect 2656 424 2658 441
rect 2872 424 2874 441
rect 3104 424 3106 441
rect 3336 424 3338 441
rect 3464 425 3466 441
rect 3462 424 3468 425
rect 1806 420 1807 424
rect 1811 420 1812 424
rect 1806 419 1812 420
rect 1830 423 1836 424
rect 1830 419 1831 423
rect 1835 419 1836 423
rect 1670 418 1676 419
rect 1830 418 1836 419
rect 1958 423 1964 424
rect 1958 419 1959 423
rect 1963 419 1964 423
rect 1958 418 1964 419
rect 2110 423 2116 424
rect 2110 419 2111 423
rect 2115 419 2116 423
rect 2110 418 2116 419
rect 2270 423 2276 424
rect 2270 419 2271 423
rect 2275 419 2276 423
rect 2270 418 2276 419
rect 2454 423 2460 424
rect 2454 419 2455 423
rect 2459 419 2460 423
rect 2454 418 2460 419
rect 2654 423 2660 424
rect 2654 419 2655 423
rect 2659 419 2660 423
rect 2654 418 2660 419
rect 2870 423 2876 424
rect 2870 419 2871 423
rect 2875 419 2876 423
rect 2870 418 2876 419
rect 3102 423 3108 424
rect 3102 419 3103 423
rect 3107 419 3108 423
rect 3102 418 3108 419
rect 3334 423 3340 424
rect 3334 419 3335 423
rect 3339 419 3340 423
rect 3462 420 3463 424
rect 3467 420 3468 424
rect 3462 419 3468 420
rect 3334 418 3340 419
rect 110 407 116 408
rect 110 403 111 407
rect 115 403 116 407
rect 1766 407 1772 408
rect 110 402 116 403
rect 134 404 140 405
rect 112 379 114 402
rect 134 400 135 404
rect 139 400 140 404
rect 134 399 140 400
rect 254 404 260 405
rect 254 400 255 404
rect 259 400 260 404
rect 254 399 260 400
rect 414 404 420 405
rect 414 400 415 404
rect 419 400 420 404
rect 414 399 420 400
rect 582 404 588 405
rect 582 400 583 404
rect 587 400 588 404
rect 582 399 588 400
rect 742 404 748 405
rect 742 400 743 404
rect 747 400 748 404
rect 742 399 748 400
rect 902 404 908 405
rect 902 400 903 404
rect 907 400 908 404
rect 902 399 908 400
rect 1046 404 1052 405
rect 1046 400 1047 404
rect 1051 400 1052 404
rect 1046 399 1052 400
rect 1182 404 1188 405
rect 1182 400 1183 404
rect 1187 400 1188 404
rect 1182 399 1188 400
rect 1310 404 1316 405
rect 1310 400 1311 404
rect 1315 400 1316 404
rect 1310 399 1316 400
rect 1438 404 1444 405
rect 1438 400 1439 404
rect 1443 400 1444 404
rect 1438 399 1444 400
rect 1566 404 1572 405
rect 1566 400 1567 404
rect 1571 400 1572 404
rect 1566 399 1572 400
rect 1670 404 1676 405
rect 1670 400 1671 404
rect 1675 400 1676 404
rect 1766 403 1767 407
rect 1771 403 1772 407
rect 1766 402 1772 403
rect 1806 407 1812 408
rect 1806 403 1807 407
rect 1811 403 1812 407
rect 3462 407 3468 408
rect 1806 402 1812 403
rect 1830 404 1836 405
rect 1670 399 1676 400
rect 136 379 138 399
rect 256 379 258 399
rect 416 379 418 399
rect 584 379 586 399
rect 744 379 746 399
rect 904 379 906 399
rect 1048 379 1050 399
rect 1184 379 1186 399
rect 1312 379 1314 399
rect 1440 379 1442 399
rect 1568 379 1570 399
rect 1672 379 1674 399
rect 1768 379 1770 402
rect 1808 379 1810 402
rect 1830 400 1831 404
rect 1835 400 1836 404
rect 1830 399 1836 400
rect 1958 404 1964 405
rect 1958 400 1959 404
rect 1963 400 1964 404
rect 1958 399 1964 400
rect 2110 404 2116 405
rect 2110 400 2111 404
rect 2115 400 2116 404
rect 2110 399 2116 400
rect 2270 404 2276 405
rect 2270 400 2271 404
rect 2275 400 2276 404
rect 2270 399 2276 400
rect 2454 404 2460 405
rect 2454 400 2455 404
rect 2459 400 2460 404
rect 2454 399 2460 400
rect 2654 404 2660 405
rect 2654 400 2655 404
rect 2659 400 2660 404
rect 2654 399 2660 400
rect 2870 404 2876 405
rect 2870 400 2871 404
rect 2875 400 2876 404
rect 2870 399 2876 400
rect 3102 404 3108 405
rect 3102 400 3103 404
rect 3107 400 3108 404
rect 3102 399 3108 400
rect 3334 404 3340 405
rect 3334 400 3335 404
rect 3339 400 3340 404
rect 3462 403 3463 407
rect 3467 403 3468 407
rect 3462 402 3468 403
rect 3334 399 3340 400
rect 1832 379 1834 399
rect 1960 379 1962 399
rect 2112 379 2114 399
rect 2272 379 2274 399
rect 2456 379 2458 399
rect 2656 379 2658 399
rect 2872 379 2874 399
rect 3104 379 3106 399
rect 3336 379 3338 399
rect 3464 379 3466 402
rect 111 378 115 379
rect 111 373 115 374
rect 135 378 139 379
rect 135 373 139 374
rect 223 378 227 379
rect 223 373 227 374
rect 255 378 259 379
rect 255 373 259 374
rect 343 378 347 379
rect 343 373 347 374
rect 415 378 419 379
rect 415 373 419 374
rect 471 378 475 379
rect 471 373 475 374
rect 583 378 587 379
rect 583 373 587 374
rect 599 378 603 379
rect 599 373 603 374
rect 719 378 723 379
rect 719 373 723 374
rect 743 378 747 379
rect 743 373 747 374
rect 839 378 843 379
rect 839 373 843 374
rect 903 378 907 379
rect 903 373 907 374
rect 959 378 963 379
rect 959 373 963 374
rect 1047 378 1051 379
rect 1047 373 1051 374
rect 1079 378 1083 379
rect 1079 373 1083 374
rect 1183 378 1187 379
rect 1183 373 1187 374
rect 1207 378 1211 379
rect 1207 373 1211 374
rect 1311 378 1315 379
rect 1311 373 1315 374
rect 1439 378 1443 379
rect 1439 373 1443 374
rect 1567 378 1571 379
rect 1567 373 1571 374
rect 1671 378 1675 379
rect 1671 373 1675 374
rect 1767 378 1771 379
rect 1767 373 1771 374
rect 1807 378 1811 379
rect 1807 373 1811 374
rect 1831 378 1835 379
rect 1831 373 1835 374
rect 1927 378 1931 379
rect 1927 373 1931 374
rect 1959 378 1963 379
rect 1959 373 1963 374
rect 2039 378 2043 379
rect 2039 373 2043 374
rect 2111 378 2115 379
rect 2111 373 2115 374
rect 2159 378 2163 379
rect 2159 373 2163 374
rect 2271 378 2275 379
rect 2271 373 2275 374
rect 2287 378 2291 379
rect 2287 373 2291 374
rect 2423 378 2427 379
rect 2423 373 2427 374
rect 2455 378 2459 379
rect 2455 373 2459 374
rect 2583 378 2587 379
rect 2583 373 2587 374
rect 2655 378 2659 379
rect 2655 373 2659 374
rect 2759 378 2763 379
rect 2759 373 2763 374
rect 2871 378 2875 379
rect 2871 373 2875 374
rect 2951 378 2955 379
rect 2951 373 2955 374
rect 3103 378 3107 379
rect 3103 373 3107 374
rect 3151 378 3155 379
rect 3151 373 3155 374
rect 3335 378 3339 379
rect 3335 373 3339 374
rect 3359 378 3363 379
rect 3359 373 3363 374
rect 3463 378 3467 379
rect 3463 373 3467 374
rect 112 354 114 373
rect 136 357 138 373
rect 224 357 226 373
rect 344 357 346 373
rect 472 357 474 373
rect 600 357 602 373
rect 720 357 722 373
rect 840 357 842 373
rect 960 357 962 373
rect 1080 357 1082 373
rect 1208 357 1210 373
rect 134 356 140 357
rect 110 353 116 354
rect 110 349 111 353
rect 115 349 116 353
rect 134 352 135 356
rect 139 352 140 356
rect 134 351 140 352
rect 222 356 228 357
rect 222 352 223 356
rect 227 352 228 356
rect 222 351 228 352
rect 342 356 348 357
rect 342 352 343 356
rect 347 352 348 356
rect 342 351 348 352
rect 470 356 476 357
rect 470 352 471 356
rect 475 352 476 356
rect 470 351 476 352
rect 598 356 604 357
rect 598 352 599 356
rect 603 352 604 356
rect 598 351 604 352
rect 718 356 724 357
rect 718 352 719 356
rect 723 352 724 356
rect 718 351 724 352
rect 838 356 844 357
rect 838 352 839 356
rect 843 352 844 356
rect 838 351 844 352
rect 958 356 964 357
rect 958 352 959 356
rect 963 352 964 356
rect 958 351 964 352
rect 1078 356 1084 357
rect 1078 352 1079 356
rect 1083 352 1084 356
rect 1078 351 1084 352
rect 1206 356 1212 357
rect 1206 352 1207 356
rect 1211 352 1212 356
rect 1768 354 1770 373
rect 1808 354 1810 373
rect 1928 357 1930 373
rect 2040 357 2042 373
rect 2160 357 2162 373
rect 2288 357 2290 373
rect 2424 357 2426 373
rect 2584 357 2586 373
rect 2760 357 2762 373
rect 2952 357 2954 373
rect 3152 357 3154 373
rect 3360 357 3362 373
rect 1926 356 1932 357
rect 1206 351 1212 352
rect 1766 353 1772 354
rect 110 348 116 349
rect 1766 349 1767 353
rect 1771 349 1772 353
rect 1766 348 1772 349
rect 1806 353 1812 354
rect 1806 349 1807 353
rect 1811 349 1812 353
rect 1926 352 1927 356
rect 1931 352 1932 356
rect 1926 351 1932 352
rect 2038 356 2044 357
rect 2038 352 2039 356
rect 2043 352 2044 356
rect 2038 351 2044 352
rect 2158 356 2164 357
rect 2158 352 2159 356
rect 2163 352 2164 356
rect 2158 351 2164 352
rect 2286 356 2292 357
rect 2286 352 2287 356
rect 2291 352 2292 356
rect 2286 351 2292 352
rect 2422 356 2428 357
rect 2422 352 2423 356
rect 2427 352 2428 356
rect 2422 351 2428 352
rect 2582 356 2588 357
rect 2582 352 2583 356
rect 2587 352 2588 356
rect 2582 351 2588 352
rect 2758 356 2764 357
rect 2758 352 2759 356
rect 2763 352 2764 356
rect 2758 351 2764 352
rect 2950 356 2956 357
rect 2950 352 2951 356
rect 2955 352 2956 356
rect 2950 351 2956 352
rect 3150 356 3156 357
rect 3150 352 3151 356
rect 3155 352 3156 356
rect 3150 351 3156 352
rect 3358 356 3364 357
rect 3358 352 3359 356
rect 3363 352 3364 356
rect 3464 354 3466 373
rect 3358 351 3364 352
rect 3462 353 3468 354
rect 1806 348 1812 349
rect 3462 349 3463 353
rect 3467 349 3468 353
rect 3462 348 3468 349
rect 134 337 140 338
rect 110 336 116 337
rect 110 332 111 336
rect 115 332 116 336
rect 134 333 135 337
rect 139 333 140 337
rect 134 332 140 333
rect 222 337 228 338
rect 222 333 223 337
rect 227 333 228 337
rect 222 332 228 333
rect 342 337 348 338
rect 342 333 343 337
rect 347 333 348 337
rect 342 332 348 333
rect 470 337 476 338
rect 470 333 471 337
rect 475 333 476 337
rect 470 332 476 333
rect 598 337 604 338
rect 598 333 599 337
rect 603 333 604 337
rect 598 332 604 333
rect 718 337 724 338
rect 718 333 719 337
rect 723 333 724 337
rect 718 332 724 333
rect 838 337 844 338
rect 838 333 839 337
rect 843 333 844 337
rect 838 332 844 333
rect 958 337 964 338
rect 958 333 959 337
rect 963 333 964 337
rect 958 332 964 333
rect 1078 337 1084 338
rect 1078 333 1079 337
rect 1083 333 1084 337
rect 1078 332 1084 333
rect 1206 337 1212 338
rect 1926 337 1932 338
rect 1206 333 1207 337
rect 1211 333 1212 337
rect 1206 332 1212 333
rect 1766 336 1772 337
rect 1766 332 1767 336
rect 1771 332 1772 336
rect 110 331 116 332
rect 112 311 114 331
rect 136 311 138 332
rect 224 311 226 332
rect 344 311 346 332
rect 472 311 474 332
rect 600 311 602 332
rect 720 311 722 332
rect 840 311 842 332
rect 960 311 962 332
rect 1080 311 1082 332
rect 1208 311 1210 332
rect 1766 331 1772 332
rect 1806 336 1812 337
rect 1806 332 1807 336
rect 1811 332 1812 336
rect 1926 333 1927 337
rect 1931 333 1932 337
rect 1926 332 1932 333
rect 2038 337 2044 338
rect 2038 333 2039 337
rect 2043 333 2044 337
rect 2038 332 2044 333
rect 2158 337 2164 338
rect 2158 333 2159 337
rect 2163 333 2164 337
rect 2158 332 2164 333
rect 2286 337 2292 338
rect 2286 333 2287 337
rect 2291 333 2292 337
rect 2286 332 2292 333
rect 2422 337 2428 338
rect 2422 333 2423 337
rect 2427 333 2428 337
rect 2422 332 2428 333
rect 2582 337 2588 338
rect 2582 333 2583 337
rect 2587 333 2588 337
rect 2582 332 2588 333
rect 2758 337 2764 338
rect 2758 333 2759 337
rect 2763 333 2764 337
rect 2758 332 2764 333
rect 2950 337 2956 338
rect 2950 333 2951 337
rect 2955 333 2956 337
rect 2950 332 2956 333
rect 3150 337 3156 338
rect 3150 333 3151 337
rect 3155 333 3156 337
rect 3150 332 3156 333
rect 3358 337 3364 338
rect 3358 333 3359 337
rect 3363 333 3364 337
rect 3358 332 3364 333
rect 3462 336 3468 337
rect 3462 332 3463 336
rect 3467 332 3468 336
rect 1806 331 1812 332
rect 1768 311 1770 331
rect 1808 315 1810 331
rect 1928 315 1930 332
rect 2040 315 2042 332
rect 2160 315 2162 332
rect 2288 315 2290 332
rect 2424 315 2426 332
rect 2584 315 2586 332
rect 2760 315 2762 332
rect 2952 315 2954 332
rect 3152 315 3154 332
rect 3360 315 3362 332
rect 3462 331 3468 332
rect 3464 315 3466 331
rect 1807 314 1811 315
rect 111 310 115 311
rect 111 305 115 306
rect 135 310 139 311
rect 135 305 139 306
rect 223 310 227 311
rect 223 305 227 306
rect 263 310 267 311
rect 263 305 267 306
rect 343 310 347 311
rect 343 305 347 306
rect 375 310 379 311
rect 375 305 379 306
rect 471 310 475 311
rect 471 305 475 306
rect 487 310 491 311
rect 487 305 491 306
rect 599 310 603 311
rect 599 305 603 306
rect 711 310 715 311
rect 711 305 715 306
rect 719 310 723 311
rect 719 305 723 306
rect 815 310 819 311
rect 815 305 819 306
rect 839 310 843 311
rect 839 305 843 306
rect 919 310 923 311
rect 919 305 923 306
rect 959 310 963 311
rect 959 305 963 306
rect 1023 310 1027 311
rect 1023 305 1027 306
rect 1079 310 1083 311
rect 1079 305 1083 306
rect 1127 310 1131 311
rect 1127 305 1131 306
rect 1207 310 1211 311
rect 1207 305 1211 306
rect 1239 310 1243 311
rect 1239 305 1243 306
rect 1767 310 1771 311
rect 1807 309 1811 310
rect 1927 314 1931 315
rect 1927 309 1931 310
rect 2039 314 2043 315
rect 2039 309 2043 310
rect 2159 314 2163 315
rect 2159 309 2163 310
rect 2223 314 2227 315
rect 2223 309 2227 310
rect 2287 314 2291 315
rect 2287 309 2291 310
rect 2311 314 2315 315
rect 2311 309 2315 310
rect 2399 314 2403 315
rect 2399 309 2403 310
rect 2423 314 2427 315
rect 2423 309 2427 310
rect 2487 314 2491 315
rect 2487 309 2491 310
rect 2575 314 2579 315
rect 2575 309 2579 310
rect 2583 314 2587 315
rect 2583 309 2587 310
rect 2679 314 2683 315
rect 2679 309 2683 310
rect 2759 314 2763 315
rect 2759 309 2763 310
rect 2799 314 2803 315
rect 2799 309 2803 310
rect 2927 314 2931 315
rect 2927 309 2931 310
rect 2951 314 2955 315
rect 2951 309 2955 310
rect 3071 314 3075 315
rect 3071 309 3075 310
rect 3151 314 3155 315
rect 3151 309 3155 310
rect 3223 314 3227 315
rect 3223 309 3227 310
rect 3359 314 3363 315
rect 3359 309 3363 310
rect 3367 314 3371 315
rect 3367 309 3371 310
rect 3463 314 3467 315
rect 3463 309 3467 310
rect 1767 305 1771 306
rect 112 289 114 305
rect 110 288 116 289
rect 264 288 266 305
rect 376 288 378 305
rect 488 288 490 305
rect 600 288 602 305
rect 712 288 714 305
rect 816 288 818 305
rect 920 288 922 305
rect 1024 288 1026 305
rect 1128 288 1130 305
rect 1240 288 1242 305
rect 1768 289 1770 305
rect 1808 293 1810 309
rect 1806 292 1812 293
rect 2224 292 2226 309
rect 2312 292 2314 309
rect 2400 292 2402 309
rect 2488 292 2490 309
rect 2576 292 2578 309
rect 2680 292 2682 309
rect 2800 292 2802 309
rect 2928 292 2930 309
rect 3072 292 3074 309
rect 3224 292 3226 309
rect 3368 292 3370 309
rect 3464 293 3466 309
rect 3462 292 3468 293
rect 1766 288 1772 289
rect 110 284 111 288
rect 115 284 116 288
rect 110 283 116 284
rect 262 287 268 288
rect 262 283 263 287
rect 267 283 268 287
rect 262 282 268 283
rect 374 287 380 288
rect 374 283 375 287
rect 379 283 380 287
rect 374 282 380 283
rect 486 287 492 288
rect 486 283 487 287
rect 491 283 492 287
rect 486 282 492 283
rect 598 287 604 288
rect 598 283 599 287
rect 603 283 604 287
rect 598 282 604 283
rect 710 287 716 288
rect 710 283 711 287
rect 715 283 716 287
rect 710 282 716 283
rect 814 287 820 288
rect 814 283 815 287
rect 819 283 820 287
rect 814 282 820 283
rect 918 287 924 288
rect 918 283 919 287
rect 923 283 924 287
rect 918 282 924 283
rect 1022 287 1028 288
rect 1022 283 1023 287
rect 1027 283 1028 287
rect 1022 282 1028 283
rect 1126 287 1132 288
rect 1126 283 1127 287
rect 1131 283 1132 287
rect 1126 282 1132 283
rect 1238 287 1244 288
rect 1238 283 1239 287
rect 1243 283 1244 287
rect 1766 284 1767 288
rect 1771 284 1772 288
rect 1806 288 1807 292
rect 1811 288 1812 292
rect 1806 287 1812 288
rect 2222 291 2228 292
rect 2222 287 2223 291
rect 2227 287 2228 291
rect 2222 286 2228 287
rect 2310 291 2316 292
rect 2310 287 2311 291
rect 2315 287 2316 291
rect 2310 286 2316 287
rect 2398 291 2404 292
rect 2398 287 2399 291
rect 2403 287 2404 291
rect 2398 286 2404 287
rect 2486 291 2492 292
rect 2486 287 2487 291
rect 2491 287 2492 291
rect 2486 286 2492 287
rect 2574 291 2580 292
rect 2574 287 2575 291
rect 2579 287 2580 291
rect 2574 286 2580 287
rect 2678 291 2684 292
rect 2678 287 2679 291
rect 2683 287 2684 291
rect 2678 286 2684 287
rect 2798 291 2804 292
rect 2798 287 2799 291
rect 2803 287 2804 291
rect 2798 286 2804 287
rect 2926 291 2932 292
rect 2926 287 2927 291
rect 2931 287 2932 291
rect 2926 286 2932 287
rect 3070 291 3076 292
rect 3070 287 3071 291
rect 3075 287 3076 291
rect 3070 286 3076 287
rect 3222 291 3228 292
rect 3222 287 3223 291
rect 3227 287 3228 291
rect 3222 286 3228 287
rect 3366 291 3372 292
rect 3366 287 3367 291
rect 3371 287 3372 291
rect 3462 288 3463 292
rect 3467 288 3468 292
rect 3462 287 3468 288
rect 3366 286 3372 287
rect 1766 283 1772 284
rect 1238 282 1244 283
rect 1806 275 1812 276
rect 110 271 116 272
rect 110 267 111 271
rect 115 267 116 271
rect 1766 271 1772 272
rect 110 266 116 267
rect 262 268 268 269
rect 112 243 114 266
rect 262 264 263 268
rect 267 264 268 268
rect 262 263 268 264
rect 374 268 380 269
rect 374 264 375 268
rect 379 264 380 268
rect 374 263 380 264
rect 486 268 492 269
rect 486 264 487 268
rect 491 264 492 268
rect 486 263 492 264
rect 598 268 604 269
rect 598 264 599 268
rect 603 264 604 268
rect 598 263 604 264
rect 710 268 716 269
rect 710 264 711 268
rect 715 264 716 268
rect 710 263 716 264
rect 814 268 820 269
rect 814 264 815 268
rect 819 264 820 268
rect 814 263 820 264
rect 918 268 924 269
rect 918 264 919 268
rect 923 264 924 268
rect 918 263 924 264
rect 1022 268 1028 269
rect 1022 264 1023 268
rect 1027 264 1028 268
rect 1022 263 1028 264
rect 1126 268 1132 269
rect 1126 264 1127 268
rect 1131 264 1132 268
rect 1126 263 1132 264
rect 1238 268 1244 269
rect 1238 264 1239 268
rect 1243 264 1244 268
rect 1766 267 1767 271
rect 1771 267 1772 271
rect 1806 271 1807 275
rect 1811 271 1812 275
rect 3462 275 3468 276
rect 1806 270 1812 271
rect 2222 272 2228 273
rect 1766 266 1772 267
rect 1238 263 1244 264
rect 264 243 266 263
rect 376 243 378 263
rect 488 243 490 263
rect 600 243 602 263
rect 712 243 714 263
rect 816 243 818 263
rect 920 243 922 263
rect 1024 243 1026 263
rect 1128 243 1130 263
rect 1240 243 1242 263
rect 1768 243 1770 266
rect 1808 243 1810 270
rect 2222 268 2223 272
rect 2227 268 2228 272
rect 2222 267 2228 268
rect 2310 272 2316 273
rect 2310 268 2311 272
rect 2315 268 2316 272
rect 2310 267 2316 268
rect 2398 272 2404 273
rect 2398 268 2399 272
rect 2403 268 2404 272
rect 2398 267 2404 268
rect 2486 272 2492 273
rect 2486 268 2487 272
rect 2491 268 2492 272
rect 2486 267 2492 268
rect 2574 272 2580 273
rect 2574 268 2575 272
rect 2579 268 2580 272
rect 2574 267 2580 268
rect 2678 272 2684 273
rect 2678 268 2679 272
rect 2683 268 2684 272
rect 2678 267 2684 268
rect 2798 272 2804 273
rect 2798 268 2799 272
rect 2803 268 2804 272
rect 2798 267 2804 268
rect 2926 272 2932 273
rect 2926 268 2927 272
rect 2931 268 2932 272
rect 2926 267 2932 268
rect 3070 272 3076 273
rect 3070 268 3071 272
rect 3075 268 3076 272
rect 3070 267 3076 268
rect 3222 272 3228 273
rect 3222 268 3223 272
rect 3227 268 3228 272
rect 3222 267 3228 268
rect 3366 272 3372 273
rect 3366 268 3367 272
rect 3371 268 3372 272
rect 3462 271 3463 275
rect 3467 271 3468 275
rect 3462 270 3468 271
rect 3366 267 3372 268
rect 2224 243 2226 267
rect 2312 243 2314 267
rect 2400 243 2402 267
rect 2488 243 2490 267
rect 2576 243 2578 267
rect 2680 243 2682 267
rect 2800 243 2802 267
rect 2928 243 2930 267
rect 3072 243 3074 267
rect 3224 243 3226 267
rect 3368 243 3370 267
rect 3464 243 3466 270
rect 111 242 115 243
rect 111 237 115 238
rect 263 242 267 243
rect 263 237 267 238
rect 375 242 379 243
rect 375 237 379 238
rect 447 242 451 243
rect 447 237 451 238
rect 487 242 491 243
rect 487 237 491 238
rect 535 242 539 243
rect 535 237 539 238
rect 599 242 603 243
rect 599 237 603 238
rect 623 242 627 243
rect 623 237 627 238
rect 711 242 715 243
rect 711 237 715 238
rect 807 242 811 243
rect 807 237 811 238
rect 815 242 819 243
rect 815 237 819 238
rect 903 242 907 243
rect 903 237 907 238
rect 919 242 923 243
rect 919 237 923 238
rect 999 242 1003 243
rect 999 237 1003 238
rect 1023 242 1027 243
rect 1023 237 1027 238
rect 1103 242 1107 243
rect 1103 237 1107 238
rect 1127 242 1131 243
rect 1127 237 1131 238
rect 1207 242 1211 243
rect 1207 237 1211 238
rect 1239 242 1243 243
rect 1239 237 1243 238
rect 1311 242 1315 243
rect 1311 237 1315 238
rect 1767 242 1771 243
rect 1767 237 1771 238
rect 1807 242 1811 243
rect 1807 237 1811 238
rect 2143 242 2147 243
rect 2143 237 2147 238
rect 2223 242 2227 243
rect 2223 237 2227 238
rect 2263 242 2267 243
rect 2263 237 2267 238
rect 2311 242 2315 243
rect 2311 237 2315 238
rect 2383 242 2387 243
rect 2383 237 2387 238
rect 2399 242 2403 243
rect 2399 237 2403 238
rect 2487 242 2491 243
rect 2487 237 2491 238
rect 2511 242 2515 243
rect 2511 237 2515 238
rect 2575 242 2579 243
rect 2575 237 2579 238
rect 2639 242 2643 243
rect 2639 237 2643 238
rect 2679 242 2683 243
rect 2679 237 2683 238
rect 2767 242 2771 243
rect 2767 237 2771 238
rect 2799 242 2803 243
rect 2799 237 2803 238
rect 2895 242 2899 243
rect 2895 237 2899 238
rect 2927 242 2931 243
rect 2927 237 2931 238
rect 3015 242 3019 243
rect 3015 237 3019 238
rect 3071 242 3075 243
rect 3071 237 3075 238
rect 3135 242 3139 243
rect 3135 237 3139 238
rect 3223 242 3227 243
rect 3223 237 3227 238
rect 3263 242 3267 243
rect 3263 237 3267 238
rect 3367 242 3371 243
rect 3367 237 3371 238
rect 3463 242 3467 243
rect 3463 237 3467 238
rect 112 218 114 237
rect 448 221 450 237
rect 536 221 538 237
rect 624 221 626 237
rect 712 221 714 237
rect 808 221 810 237
rect 904 221 906 237
rect 1000 221 1002 237
rect 1104 221 1106 237
rect 1208 221 1210 237
rect 1312 221 1314 237
rect 446 220 452 221
rect 110 217 116 218
rect 110 213 111 217
rect 115 213 116 217
rect 446 216 447 220
rect 451 216 452 220
rect 446 215 452 216
rect 534 220 540 221
rect 534 216 535 220
rect 539 216 540 220
rect 534 215 540 216
rect 622 220 628 221
rect 622 216 623 220
rect 627 216 628 220
rect 622 215 628 216
rect 710 220 716 221
rect 710 216 711 220
rect 715 216 716 220
rect 710 215 716 216
rect 806 220 812 221
rect 806 216 807 220
rect 811 216 812 220
rect 806 215 812 216
rect 902 220 908 221
rect 902 216 903 220
rect 907 216 908 220
rect 902 215 908 216
rect 998 220 1004 221
rect 998 216 999 220
rect 1003 216 1004 220
rect 998 215 1004 216
rect 1102 220 1108 221
rect 1102 216 1103 220
rect 1107 216 1108 220
rect 1102 215 1108 216
rect 1206 220 1212 221
rect 1206 216 1207 220
rect 1211 216 1212 220
rect 1206 215 1212 216
rect 1310 220 1316 221
rect 1310 216 1311 220
rect 1315 216 1316 220
rect 1768 218 1770 237
rect 1808 218 1810 237
rect 2144 221 2146 237
rect 2264 221 2266 237
rect 2384 221 2386 237
rect 2512 221 2514 237
rect 2640 221 2642 237
rect 2768 221 2770 237
rect 2896 221 2898 237
rect 3016 221 3018 237
rect 3136 221 3138 237
rect 3264 221 3266 237
rect 3368 221 3370 237
rect 2142 220 2148 221
rect 1310 215 1316 216
rect 1766 217 1772 218
rect 110 212 116 213
rect 1766 213 1767 217
rect 1771 213 1772 217
rect 1766 212 1772 213
rect 1806 217 1812 218
rect 1806 213 1807 217
rect 1811 213 1812 217
rect 2142 216 2143 220
rect 2147 216 2148 220
rect 2142 215 2148 216
rect 2262 220 2268 221
rect 2262 216 2263 220
rect 2267 216 2268 220
rect 2262 215 2268 216
rect 2382 220 2388 221
rect 2382 216 2383 220
rect 2387 216 2388 220
rect 2382 215 2388 216
rect 2510 220 2516 221
rect 2510 216 2511 220
rect 2515 216 2516 220
rect 2510 215 2516 216
rect 2638 220 2644 221
rect 2638 216 2639 220
rect 2643 216 2644 220
rect 2638 215 2644 216
rect 2766 220 2772 221
rect 2766 216 2767 220
rect 2771 216 2772 220
rect 2766 215 2772 216
rect 2894 220 2900 221
rect 2894 216 2895 220
rect 2899 216 2900 220
rect 2894 215 2900 216
rect 3014 220 3020 221
rect 3014 216 3015 220
rect 3019 216 3020 220
rect 3014 215 3020 216
rect 3134 220 3140 221
rect 3134 216 3135 220
rect 3139 216 3140 220
rect 3134 215 3140 216
rect 3262 220 3268 221
rect 3262 216 3263 220
rect 3267 216 3268 220
rect 3262 215 3268 216
rect 3366 220 3372 221
rect 3366 216 3367 220
rect 3371 216 3372 220
rect 3464 218 3466 237
rect 3366 215 3372 216
rect 3462 217 3468 218
rect 1806 212 1812 213
rect 3462 213 3463 217
rect 3467 213 3468 217
rect 3462 212 3468 213
rect 446 201 452 202
rect 110 200 116 201
rect 110 196 111 200
rect 115 196 116 200
rect 446 197 447 201
rect 451 197 452 201
rect 446 196 452 197
rect 534 201 540 202
rect 534 197 535 201
rect 539 197 540 201
rect 534 196 540 197
rect 622 201 628 202
rect 622 197 623 201
rect 627 197 628 201
rect 622 196 628 197
rect 710 201 716 202
rect 710 197 711 201
rect 715 197 716 201
rect 710 196 716 197
rect 806 201 812 202
rect 806 197 807 201
rect 811 197 812 201
rect 806 196 812 197
rect 902 201 908 202
rect 902 197 903 201
rect 907 197 908 201
rect 902 196 908 197
rect 998 201 1004 202
rect 998 197 999 201
rect 1003 197 1004 201
rect 998 196 1004 197
rect 1102 201 1108 202
rect 1102 197 1103 201
rect 1107 197 1108 201
rect 1102 196 1108 197
rect 1206 201 1212 202
rect 1206 197 1207 201
rect 1211 197 1212 201
rect 1206 196 1212 197
rect 1310 201 1316 202
rect 2142 201 2148 202
rect 1310 197 1311 201
rect 1315 197 1316 201
rect 1310 196 1316 197
rect 1766 200 1772 201
rect 1766 196 1767 200
rect 1771 196 1772 200
rect 110 195 116 196
rect 112 151 114 195
rect 448 151 450 196
rect 536 151 538 196
rect 624 151 626 196
rect 712 151 714 196
rect 808 151 810 196
rect 904 151 906 196
rect 1000 151 1002 196
rect 1104 151 1106 196
rect 1208 151 1210 196
rect 1312 151 1314 196
rect 1766 195 1772 196
rect 1806 200 1812 201
rect 1806 196 1807 200
rect 1811 196 1812 200
rect 2142 197 2143 201
rect 2147 197 2148 201
rect 2142 196 2148 197
rect 2262 201 2268 202
rect 2262 197 2263 201
rect 2267 197 2268 201
rect 2262 196 2268 197
rect 2382 201 2388 202
rect 2382 197 2383 201
rect 2387 197 2388 201
rect 2382 196 2388 197
rect 2510 201 2516 202
rect 2510 197 2511 201
rect 2515 197 2516 201
rect 2510 196 2516 197
rect 2638 201 2644 202
rect 2638 197 2639 201
rect 2643 197 2644 201
rect 2638 196 2644 197
rect 2766 201 2772 202
rect 2766 197 2767 201
rect 2771 197 2772 201
rect 2766 196 2772 197
rect 2894 201 2900 202
rect 2894 197 2895 201
rect 2899 197 2900 201
rect 2894 196 2900 197
rect 3014 201 3020 202
rect 3014 197 3015 201
rect 3019 197 3020 201
rect 3014 196 3020 197
rect 3134 201 3140 202
rect 3134 197 3135 201
rect 3139 197 3140 201
rect 3134 196 3140 197
rect 3262 201 3268 202
rect 3262 197 3263 201
rect 3267 197 3268 201
rect 3262 196 3268 197
rect 3366 201 3372 202
rect 3366 197 3367 201
rect 3371 197 3372 201
rect 3366 196 3372 197
rect 3462 200 3468 201
rect 3462 196 3463 200
rect 3467 196 3468 200
rect 1806 195 1812 196
rect 1768 151 1770 195
rect 1808 155 1810 195
rect 2144 155 2146 196
rect 2264 155 2266 196
rect 2384 155 2386 196
rect 2512 155 2514 196
rect 2640 155 2642 196
rect 2768 155 2770 196
rect 2896 155 2898 196
rect 3016 155 3018 196
rect 3136 155 3138 196
rect 3264 155 3266 196
rect 3368 155 3370 196
rect 3462 195 3468 196
rect 3464 155 3466 195
rect 1807 154 1811 155
rect 111 150 115 151
rect 111 145 115 146
rect 263 150 267 151
rect 263 145 267 146
rect 351 150 355 151
rect 351 145 355 146
rect 439 150 443 151
rect 439 145 443 146
rect 447 150 451 151
rect 447 145 451 146
rect 527 150 531 151
rect 527 145 531 146
rect 535 150 539 151
rect 535 145 539 146
rect 615 150 619 151
rect 615 145 619 146
rect 623 150 627 151
rect 623 145 627 146
rect 703 150 707 151
rect 703 145 707 146
rect 711 150 715 151
rect 711 145 715 146
rect 791 150 795 151
rect 791 145 795 146
rect 807 150 811 151
rect 807 145 811 146
rect 879 150 883 151
rect 879 145 883 146
rect 903 150 907 151
rect 903 145 907 146
rect 967 150 971 151
rect 967 145 971 146
rect 999 150 1003 151
rect 999 145 1003 146
rect 1055 150 1059 151
rect 1055 145 1059 146
rect 1103 150 1107 151
rect 1103 145 1107 146
rect 1143 150 1147 151
rect 1143 145 1147 146
rect 1207 150 1211 151
rect 1207 145 1211 146
rect 1231 150 1235 151
rect 1231 145 1235 146
rect 1311 150 1315 151
rect 1311 145 1315 146
rect 1319 150 1323 151
rect 1319 145 1323 146
rect 1407 150 1411 151
rect 1407 145 1411 146
rect 1495 150 1499 151
rect 1495 145 1499 146
rect 1583 150 1587 151
rect 1583 145 1587 146
rect 1671 150 1675 151
rect 1671 145 1675 146
rect 1767 150 1771 151
rect 1807 149 1811 150
rect 1831 154 1835 155
rect 1831 149 1835 150
rect 1919 154 1923 155
rect 1919 149 1923 150
rect 2007 154 2011 155
rect 2007 149 2011 150
rect 2095 154 2099 155
rect 2095 149 2099 150
rect 2143 154 2147 155
rect 2143 149 2147 150
rect 2183 154 2187 155
rect 2183 149 2187 150
rect 2263 154 2267 155
rect 2263 149 2267 150
rect 2295 154 2299 155
rect 2295 149 2299 150
rect 2383 154 2387 155
rect 2383 149 2387 150
rect 2407 154 2411 155
rect 2407 149 2411 150
rect 2511 154 2515 155
rect 2511 149 2515 150
rect 2615 154 2619 155
rect 2615 149 2619 150
rect 2639 154 2643 155
rect 2639 149 2643 150
rect 2719 154 2723 155
rect 2719 149 2723 150
rect 2767 154 2771 155
rect 2767 149 2771 150
rect 2815 154 2819 155
rect 2815 149 2819 150
rect 2895 154 2899 155
rect 2895 149 2899 150
rect 2911 154 2915 155
rect 2911 149 2915 150
rect 3007 154 3011 155
rect 3007 149 3011 150
rect 3015 154 3019 155
rect 3015 149 3019 150
rect 3103 154 3107 155
rect 3103 149 3107 150
rect 3135 154 3139 155
rect 3135 149 3139 150
rect 3191 154 3195 155
rect 3191 149 3195 150
rect 3263 154 3267 155
rect 3263 149 3267 150
rect 3279 154 3283 155
rect 3279 149 3283 150
rect 3367 154 3371 155
rect 3367 149 3371 150
rect 3463 154 3467 155
rect 3463 149 3467 150
rect 1767 145 1771 146
rect 112 129 114 145
rect 110 128 116 129
rect 264 128 266 145
rect 352 128 354 145
rect 440 128 442 145
rect 528 128 530 145
rect 616 128 618 145
rect 704 128 706 145
rect 792 128 794 145
rect 880 128 882 145
rect 968 128 970 145
rect 1056 128 1058 145
rect 1144 128 1146 145
rect 1232 128 1234 145
rect 1320 128 1322 145
rect 1408 128 1410 145
rect 1496 128 1498 145
rect 1584 128 1586 145
rect 1672 128 1674 145
rect 1768 129 1770 145
rect 1808 133 1810 149
rect 1806 132 1812 133
rect 1832 132 1834 149
rect 1920 132 1922 149
rect 2008 132 2010 149
rect 2096 132 2098 149
rect 2184 132 2186 149
rect 2296 132 2298 149
rect 2408 132 2410 149
rect 2512 132 2514 149
rect 2616 132 2618 149
rect 2720 132 2722 149
rect 2816 132 2818 149
rect 2912 132 2914 149
rect 3008 132 3010 149
rect 3104 132 3106 149
rect 3192 132 3194 149
rect 3280 132 3282 149
rect 3368 132 3370 149
rect 3464 133 3466 149
rect 3462 132 3468 133
rect 1766 128 1772 129
rect 110 124 111 128
rect 115 124 116 128
rect 110 123 116 124
rect 262 127 268 128
rect 262 123 263 127
rect 267 123 268 127
rect 262 122 268 123
rect 350 127 356 128
rect 350 123 351 127
rect 355 123 356 127
rect 350 122 356 123
rect 438 127 444 128
rect 438 123 439 127
rect 443 123 444 127
rect 438 122 444 123
rect 526 127 532 128
rect 526 123 527 127
rect 531 123 532 127
rect 526 122 532 123
rect 614 127 620 128
rect 614 123 615 127
rect 619 123 620 127
rect 614 122 620 123
rect 702 127 708 128
rect 702 123 703 127
rect 707 123 708 127
rect 702 122 708 123
rect 790 127 796 128
rect 790 123 791 127
rect 795 123 796 127
rect 790 122 796 123
rect 878 127 884 128
rect 878 123 879 127
rect 883 123 884 127
rect 878 122 884 123
rect 966 127 972 128
rect 966 123 967 127
rect 971 123 972 127
rect 966 122 972 123
rect 1054 127 1060 128
rect 1054 123 1055 127
rect 1059 123 1060 127
rect 1054 122 1060 123
rect 1142 127 1148 128
rect 1142 123 1143 127
rect 1147 123 1148 127
rect 1142 122 1148 123
rect 1230 127 1236 128
rect 1230 123 1231 127
rect 1235 123 1236 127
rect 1230 122 1236 123
rect 1318 127 1324 128
rect 1318 123 1319 127
rect 1323 123 1324 127
rect 1318 122 1324 123
rect 1406 127 1412 128
rect 1406 123 1407 127
rect 1411 123 1412 127
rect 1406 122 1412 123
rect 1494 127 1500 128
rect 1494 123 1495 127
rect 1499 123 1500 127
rect 1494 122 1500 123
rect 1582 127 1588 128
rect 1582 123 1583 127
rect 1587 123 1588 127
rect 1582 122 1588 123
rect 1670 127 1676 128
rect 1670 123 1671 127
rect 1675 123 1676 127
rect 1766 124 1767 128
rect 1771 124 1772 128
rect 1806 128 1807 132
rect 1811 128 1812 132
rect 1806 127 1812 128
rect 1830 131 1836 132
rect 1830 127 1831 131
rect 1835 127 1836 131
rect 1830 126 1836 127
rect 1918 131 1924 132
rect 1918 127 1919 131
rect 1923 127 1924 131
rect 1918 126 1924 127
rect 2006 131 2012 132
rect 2006 127 2007 131
rect 2011 127 2012 131
rect 2006 126 2012 127
rect 2094 131 2100 132
rect 2094 127 2095 131
rect 2099 127 2100 131
rect 2094 126 2100 127
rect 2182 131 2188 132
rect 2182 127 2183 131
rect 2187 127 2188 131
rect 2182 126 2188 127
rect 2294 131 2300 132
rect 2294 127 2295 131
rect 2299 127 2300 131
rect 2294 126 2300 127
rect 2406 131 2412 132
rect 2406 127 2407 131
rect 2411 127 2412 131
rect 2406 126 2412 127
rect 2510 131 2516 132
rect 2510 127 2511 131
rect 2515 127 2516 131
rect 2510 126 2516 127
rect 2614 131 2620 132
rect 2614 127 2615 131
rect 2619 127 2620 131
rect 2614 126 2620 127
rect 2718 131 2724 132
rect 2718 127 2719 131
rect 2723 127 2724 131
rect 2718 126 2724 127
rect 2814 131 2820 132
rect 2814 127 2815 131
rect 2819 127 2820 131
rect 2814 126 2820 127
rect 2910 131 2916 132
rect 2910 127 2911 131
rect 2915 127 2916 131
rect 2910 126 2916 127
rect 3006 131 3012 132
rect 3006 127 3007 131
rect 3011 127 3012 131
rect 3006 126 3012 127
rect 3102 131 3108 132
rect 3102 127 3103 131
rect 3107 127 3108 131
rect 3102 126 3108 127
rect 3190 131 3196 132
rect 3190 127 3191 131
rect 3195 127 3196 131
rect 3190 126 3196 127
rect 3278 131 3284 132
rect 3278 127 3279 131
rect 3283 127 3284 131
rect 3278 126 3284 127
rect 3366 131 3372 132
rect 3366 127 3367 131
rect 3371 127 3372 131
rect 3462 128 3463 132
rect 3467 128 3468 132
rect 3462 127 3468 128
rect 3366 126 3372 127
rect 1766 123 1772 124
rect 1670 122 1676 123
rect 1806 115 1812 116
rect 110 111 116 112
rect 110 107 111 111
rect 115 107 116 111
rect 1766 111 1772 112
rect 110 106 116 107
rect 262 108 268 109
rect 112 87 114 106
rect 262 104 263 108
rect 267 104 268 108
rect 262 103 268 104
rect 350 108 356 109
rect 350 104 351 108
rect 355 104 356 108
rect 350 103 356 104
rect 438 108 444 109
rect 438 104 439 108
rect 443 104 444 108
rect 438 103 444 104
rect 526 108 532 109
rect 526 104 527 108
rect 531 104 532 108
rect 526 103 532 104
rect 614 108 620 109
rect 614 104 615 108
rect 619 104 620 108
rect 614 103 620 104
rect 702 108 708 109
rect 702 104 703 108
rect 707 104 708 108
rect 702 103 708 104
rect 790 108 796 109
rect 790 104 791 108
rect 795 104 796 108
rect 790 103 796 104
rect 878 108 884 109
rect 878 104 879 108
rect 883 104 884 108
rect 878 103 884 104
rect 966 108 972 109
rect 966 104 967 108
rect 971 104 972 108
rect 966 103 972 104
rect 1054 108 1060 109
rect 1054 104 1055 108
rect 1059 104 1060 108
rect 1054 103 1060 104
rect 1142 108 1148 109
rect 1142 104 1143 108
rect 1147 104 1148 108
rect 1142 103 1148 104
rect 1230 108 1236 109
rect 1230 104 1231 108
rect 1235 104 1236 108
rect 1230 103 1236 104
rect 1318 108 1324 109
rect 1318 104 1319 108
rect 1323 104 1324 108
rect 1318 103 1324 104
rect 1406 108 1412 109
rect 1406 104 1407 108
rect 1411 104 1412 108
rect 1406 103 1412 104
rect 1494 108 1500 109
rect 1494 104 1495 108
rect 1499 104 1500 108
rect 1494 103 1500 104
rect 1582 108 1588 109
rect 1582 104 1583 108
rect 1587 104 1588 108
rect 1582 103 1588 104
rect 1670 108 1676 109
rect 1670 104 1671 108
rect 1675 104 1676 108
rect 1766 107 1767 111
rect 1771 107 1772 111
rect 1806 111 1807 115
rect 1811 111 1812 115
rect 3462 115 3468 116
rect 1806 110 1812 111
rect 1830 112 1836 113
rect 1766 106 1772 107
rect 1670 103 1676 104
rect 264 87 266 103
rect 352 87 354 103
rect 440 87 442 103
rect 528 87 530 103
rect 616 87 618 103
rect 704 87 706 103
rect 792 87 794 103
rect 880 87 882 103
rect 968 87 970 103
rect 1056 87 1058 103
rect 1144 87 1146 103
rect 1232 87 1234 103
rect 1320 87 1322 103
rect 1408 87 1410 103
rect 1496 87 1498 103
rect 1584 87 1586 103
rect 1672 87 1674 103
rect 1768 87 1770 106
rect 1808 91 1810 110
rect 1830 108 1831 112
rect 1835 108 1836 112
rect 1830 107 1836 108
rect 1918 112 1924 113
rect 1918 108 1919 112
rect 1923 108 1924 112
rect 1918 107 1924 108
rect 2006 112 2012 113
rect 2006 108 2007 112
rect 2011 108 2012 112
rect 2006 107 2012 108
rect 2094 112 2100 113
rect 2094 108 2095 112
rect 2099 108 2100 112
rect 2094 107 2100 108
rect 2182 112 2188 113
rect 2182 108 2183 112
rect 2187 108 2188 112
rect 2182 107 2188 108
rect 2294 112 2300 113
rect 2294 108 2295 112
rect 2299 108 2300 112
rect 2294 107 2300 108
rect 2406 112 2412 113
rect 2406 108 2407 112
rect 2411 108 2412 112
rect 2406 107 2412 108
rect 2510 112 2516 113
rect 2510 108 2511 112
rect 2515 108 2516 112
rect 2510 107 2516 108
rect 2614 112 2620 113
rect 2614 108 2615 112
rect 2619 108 2620 112
rect 2614 107 2620 108
rect 2718 112 2724 113
rect 2718 108 2719 112
rect 2723 108 2724 112
rect 2718 107 2724 108
rect 2814 112 2820 113
rect 2814 108 2815 112
rect 2819 108 2820 112
rect 2814 107 2820 108
rect 2910 112 2916 113
rect 2910 108 2911 112
rect 2915 108 2916 112
rect 2910 107 2916 108
rect 3006 112 3012 113
rect 3006 108 3007 112
rect 3011 108 3012 112
rect 3006 107 3012 108
rect 3102 112 3108 113
rect 3102 108 3103 112
rect 3107 108 3108 112
rect 3102 107 3108 108
rect 3190 112 3196 113
rect 3190 108 3191 112
rect 3195 108 3196 112
rect 3190 107 3196 108
rect 3278 112 3284 113
rect 3278 108 3279 112
rect 3283 108 3284 112
rect 3278 107 3284 108
rect 3366 112 3372 113
rect 3366 108 3367 112
rect 3371 108 3372 112
rect 3462 111 3463 115
rect 3467 111 3468 115
rect 3462 110 3468 111
rect 3366 107 3372 108
rect 1832 91 1834 107
rect 1920 91 1922 107
rect 2008 91 2010 107
rect 2096 91 2098 107
rect 2184 91 2186 107
rect 2296 91 2298 107
rect 2408 91 2410 107
rect 2512 91 2514 107
rect 2616 91 2618 107
rect 2720 91 2722 107
rect 2816 91 2818 107
rect 2912 91 2914 107
rect 3008 91 3010 107
rect 3104 91 3106 107
rect 3192 91 3194 107
rect 3280 91 3282 107
rect 3368 91 3370 107
rect 3464 91 3466 110
rect 1807 90 1811 91
rect 111 86 115 87
rect 111 81 115 82
rect 263 86 267 87
rect 263 81 267 82
rect 351 86 355 87
rect 351 81 355 82
rect 439 86 443 87
rect 439 81 443 82
rect 527 86 531 87
rect 527 81 531 82
rect 615 86 619 87
rect 615 81 619 82
rect 703 86 707 87
rect 703 81 707 82
rect 791 86 795 87
rect 791 81 795 82
rect 879 86 883 87
rect 879 81 883 82
rect 967 86 971 87
rect 967 81 971 82
rect 1055 86 1059 87
rect 1055 81 1059 82
rect 1143 86 1147 87
rect 1143 81 1147 82
rect 1231 86 1235 87
rect 1231 81 1235 82
rect 1319 86 1323 87
rect 1319 81 1323 82
rect 1407 86 1411 87
rect 1407 81 1411 82
rect 1495 86 1499 87
rect 1495 81 1499 82
rect 1583 86 1587 87
rect 1583 81 1587 82
rect 1671 86 1675 87
rect 1671 81 1675 82
rect 1767 86 1771 87
rect 1807 85 1811 86
rect 1831 90 1835 91
rect 1831 85 1835 86
rect 1919 90 1923 91
rect 1919 85 1923 86
rect 2007 90 2011 91
rect 2007 85 2011 86
rect 2095 90 2099 91
rect 2095 85 2099 86
rect 2183 90 2187 91
rect 2183 85 2187 86
rect 2295 90 2299 91
rect 2295 85 2299 86
rect 2407 90 2411 91
rect 2407 85 2411 86
rect 2511 90 2515 91
rect 2511 85 2515 86
rect 2615 90 2619 91
rect 2615 85 2619 86
rect 2719 90 2723 91
rect 2719 85 2723 86
rect 2815 90 2819 91
rect 2815 85 2819 86
rect 2911 90 2915 91
rect 2911 85 2915 86
rect 3007 90 3011 91
rect 3007 85 3011 86
rect 3103 90 3107 91
rect 3103 85 3107 86
rect 3191 90 3195 91
rect 3191 85 3195 86
rect 3279 90 3283 91
rect 3279 85 3283 86
rect 3367 90 3371 91
rect 3367 85 3371 86
rect 3463 90 3467 91
rect 3463 85 3467 86
rect 1767 81 1771 82
<< m4c >>
rect 111 3502 115 3506
rect 135 3502 139 3506
rect 271 3502 275 3506
rect 439 3502 443 3506
rect 615 3502 619 3506
rect 791 3502 795 3506
rect 959 3502 963 3506
rect 1119 3502 1123 3506
rect 1263 3502 1267 3506
rect 1407 3502 1411 3506
rect 1551 3502 1555 3506
rect 1671 3502 1675 3506
rect 1767 3502 1771 3506
rect 1807 3490 1811 3494
rect 1831 3490 1835 3494
rect 1975 3490 1979 3494
rect 2143 3490 2147 3494
rect 2311 3490 2315 3494
rect 2479 3490 2483 3494
rect 2639 3490 2643 3494
rect 2799 3490 2803 3494
rect 2967 3490 2971 3494
rect 3463 3490 3467 3494
rect 111 3434 115 3438
rect 135 3434 139 3438
rect 255 3434 259 3438
rect 271 3434 275 3438
rect 415 3434 419 3438
rect 439 3434 443 3438
rect 575 3434 579 3438
rect 615 3434 619 3438
rect 735 3434 739 3438
rect 791 3434 795 3438
rect 895 3434 899 3438
rect 959 3434 963 3438
rect 1063 3434 1067 3438
rect 1119 3434 1123 3438
rect 1231 3434 1235 3438
rect 1263 3434 1267 3438
rect 1399 3434 1403 3438
rect 1407 3434 1411 3438
rect 1551 3434 1555 3438
rect 1671 3434 1675 3438
rect 1767 3434 1771 3438
rect 1807 3426 1811 3430
rect 1831 3426 1835 3430
rect 1975 3426 1979 3430
rect 2031 3426 2035 3430
rect 2143 3426 2147 3430
rect 2151 3426 2155 3430
rect 2271 3426 2275 3430
rect 2311 3426 2315 3430
rect 2391 3426 2395 3430
rect 2479 3426 2483 3430
rect 2511 3426 2515 3430
rect 2623 3426 2627 3430
rect 2639 3426 2643 3430
rect 2727 3426 2731 3430
rect 2799 3426 2803 3430
rect 2831 3426 2835 3430
rect 2935 3426 2939 3430
rect 2967 3426 2971 3430
rect 3039 3426 3043 3430
rect 3151 3426 3155 3430
rect 3463 3426 3467 3430
rect 111 3362 115 3366
rect 135 3362 139 3366
rect 255 3362 259 3366
rect 327 3362 331 3366
rect 415 3362 419 3366
rect 535 3362 539 3366
rect 575 3362 579 3366
rect 735 3362 739 3366
rect 743 3362 747 3366
rect 895 3362 899 3366
rect 935 3362 939 3366
rect 1063 3362 1067 3366
rect 1119 3362 1123 3366
rect 1231 3362 1235 3366
rect 1295 3362 1299 3366
rect 1399 3362 1403 3366
rect 1463 3362 1467 3366
rect 1639 3362 1643 3366
rect 1767 3362 1771 3366
rect 1807 3358 1811 3362
rect 2031 3358 2035 3362
rect 2151 3358 2155 3362
rect 2159 3358 2163 3362
rect 2271 3358 2275 3362
rect 2295 3358 2299 3362
rect 2391 3358 2395 3362
rect 2431 3358 2435 3362
rect 2511 3358 2515 3362
rect 2567 3358 2571 3362
rect 2623 3358 2627 3362
rect 2703 3358 2707 3362
rect 2727 3358 2731 3362
rect 2831 3358 2835 3362
rect 2839 3358 2843 3362
rect 2935 3358 2939 3362
rect 2975 3358 2979 3362
rect 3039 3358 3043 3362
rect 3119 3358 3123 3362
rect 3151 3358 3155 3362
rect 3463 3358 3467 3362
rect 111 3290 115 3294
rect 135 3290 139 3294
rect 279 3290 283 3294
rect 327 3290 331 3294
rect 463 3290 467 3294
rect 535 3290 539 3294
rect 647 3290 651 3294
rect 743 3290 747 3294
rect 831 3290 835 3294
rect 935 3290 939 3294
rect 1007 3290 1011 3294
rect 1119 3290 1123 3294
rect 1175 3290 1179 3294
rect 1295 3290 1299 3294
rect 1343 3290 1347 3294
rect 1463 3290 1467 3294
rect 1503 3290 1507 3294
rect 1639 3290 1643 3294
rect 1671 3290 1675 3294
rect 1767 3290 1771 3294
rect 1807 3294 1811 3298
rect 2087 3294 2091 3298
rect 2159 3294 2163 3298
rect 2239 3294 2243 3298
rect 2295 3294 2299 3298
rect 2399 3294 2403 3298
rect 2431 3294 2435 3298
rect 2559 3294 2563 3298
rect 2567 3294 2571 3298
rect 2703 3294 2707 3298
rect 2719 3294 2723 3298
rect 2839 3294 2843 3298
rect 2879 3294 2883 3298
rect 2975 3294 2979 3298
rect 3039 3294 3043 3298
rect 3119 3294 3123 3298
rect 3199 3294 3203 3298
rect 3463 3294 3467 3298
rect 1807 3226 1811 3230
rect 1911 3226 1915 3230
rect 2047 3226 2051 3230
rect 2087 3226 2091 3230
rect 2199 3226 2203 3230
rect 2239 3226 2243 3230
rect 2359 3226 2363 3230
rect 2399 3226 2403 3230
rect 2527 3226 2531 3230
rect 2559 3226 2563 3230
rect 2687 3226 2691 3230
rect 2719 3226 2723 3230
rect 2847 3226 2851 3230
rect 2879 3226 2883 3230
rect 3007 3226 3011 3230
rect 3039 3226 3043 3230
rect 3167 3226 3171 3230
rect 3199 3226 3203 3230
rect 3335 3226 3339 3230
rect 3463 3226 3467 3230
rect 111 3218 115 3222
rect 135 3218 139 3222
rect 183 3218 187 3222
rect 279 3218 283 3222
rect 327 3218 331 3222
rect 463 3218 467 3222
rect 487 3218 491 3222
rect 647 3218 651 3222
rect 807 3218 811 3222
rect 831 3218 835 3222
rect 967 3218 971 3222
rect 1007 3218 1011 3222
rect 1135 3218 1139 3222
rect 1175 3218 1179 3222
rect 1303 3218 1307 3222
rect 1343 3218 1347 3222
rect 1471 3218 1475 3222
rect 1503 3218 1507 3222
rect 1671 3218 1675 3222
rect 1767 3218 1771 3222
rect 1807 3162 1811 3166
rect 1831 3162 1835 3166
rect 1911 3162 1915 3166
rect 2007 3162 2011 3166
rect 2047 3162 2051 3166
rect 2199 3162 2203 3166
rect 2207 3162 2211 3166
rect 2359 3162 2363 3166
rect 2399 3162 2403 3166
rect 2527 3162 2531 3166
rect 2583 3162 2587 3166
rect 2687 3162 2691 3166
rect 2759 3162 2763 3166
rect 2847 3162 2851 3166
rect 2919 3162 2923 3166
rect 3007 3162 3011 3166
rect 3079 3162 3083 3166
rect 3167 3162 3171 3166
rect 3231 3162 3235 3166
rect 3335 3162 3339 3166
rect 3367 3162 3371 3166
rect 3463 3162 3467 3166
rect 111 3154 115 3158
rect 183 3154 187 3158
rect 327 3154 331 3158
rect 367 3154 371 3158
rect 487 3154 491 3158
rect 607 3154 611 3158
rect 647 3154 651 3158
rect 727 3154 731 3158
rect 807 3154 811 3158
rect 847 3154 851 3158
rect 967 3154 971 3158
rect 1079 3154 1083 3158
rect 1135 3154 1139 3158
rect 1199 3154 1203 3158
rect 1303 3154 1307 3158
rect 1319 3154 1323 3158
rect 1471 3154 1475 3158
rect 1767 3154 1771 3158
rect 111 3086 115 3090
rect 367 3086 371 3090
rect 439 3086 443 3090
rect 487 3086 491 3090
rect 527 3086 531 3090
rect 607 3086 611 3090
rect 615 3086 619 3090
rect 703 3086 707 3090
rect 727 3086 731 3090
rect 791 3086 795 3090
rect 847 3086 851 3090
rect 879 3086 883 3090
rect 967 3086 971 3090
rect 1055 3086 1059 3090
rect 1079 3086 1083 3090
rect 1143 3086 1147 3090
rect 1199 3086 1203 3090
rect 1319 3086 1323 3090
rect 1767 3086 1771 3090
rect 1807 3090 1811 3094
rect 1831 3090 1835 3094
rect 1959 3090 1963 3094
rect 2007 3090 2011 3094
rect 2119 3090 2123 3094
rect 2207 3090 2211 3094
rect 2295 3090 2299 3094
rect 2399 3090 2403 3094
rect 2487 3090 2491 3094
rect 2583 3090 2587 3094
rect 2695 3090 2699 3094
rect 2759 3090 2763 3094
rect 2919 3090 2923 3094
rect 3079 3090 3083 3094
rect 3151 3090 3155 3094
rect 3231 3090 3235 3094
rect 3367 3090 3371 3094
rect 3463 3090 3467 3094
rect 111 3014 115 3018
rect 439 3014 443 3018
rect 503 3014 507 3018
rect 527 3014 531 3018
rect 591 3014 595 3018
rect 615 3014 619 3018
rect 679 3014 683 3018
rect 703 3014 707 3018
rect 767 3014 771 3018
rect 791 3014 795 3018
rect 855 3014 859 3018
rect 879 3014 883 3018
rect 943 3014 947 3018
rect 967 3014 971 3018
rect 1031 3014 1035 3018
rect 1055 3014 1059 3018
rect 1119 3014 1123 3018
rect 1143 3014 1147 3018
rect 1207 3014 1211 3018
rect 1295 3014 1299 3018
rect 1767 3014 1771 3018
rect 1807 3010 1811 3014
rect 1831 3010 1835 3014
rect 1919 3010 1923 3014
rect 1959 3010 1963 3014
rect 2031 3010 2035 3014
rect 2119 3010 2123 3014
rect 2143 3010 2147 3014
rect 2247 3010 2251 3014
rect 2295 3010 2299 3014
rect 2359 3010 2363 3014
rect 2479 3010 2483 3014
rect 2487 3010 2491 3014
rect 2623 3010 2627 3014
rect 2695 3010 2699 3014
rect 2791 3010 2795 3014
rect 2919 3010 2923 3014
rect 2983 3010 2987 3014
rect 3151 3010 3155 3014
rect 3183 3010 3187 3014
rect 3367 3010 3371 3014
rect 3463 3010 3467 3014
rect 111 2938 115 2942
rect 327 2938 331 2942
rect 447 2938 451 2942
rect 503 2938 507 2942
rect 575 2938 579 2942
rect 591 2938 595 2942
rect 679 2938 683 2942
rect 711 2938 715 2942
rect 767 2938 771 2942
rect 847 2938 851 2942
rect 855 2938 859 2942
rect 943 2938 947 2942
rect 975 2938 979 2942
rect 1031 2938 1035 2942
rect 1103 2938 1107 2942
rect 1119 2938 1123 2942
rect 1207 2938 1211 2942
rect 1231 2938 1235 2942
rect 1295 2938 1299 2942
rect 1359 2938 1363 2942
rect 1495 2938 1499 2942
rect 1767 2938 1771 2942
rect 1807 2934 1811 2938
rect 1831 2934 1835 2938
rect 1919 2934 1923 2938
rect 2015 2934 2019 2938
rect 2031 2934 2035 2938
rect 2143 2934 2147 2938
rect 2215 2934 2219 2938
rect 2247 2934 2251 2938
rect 2359 2934 2363 2938
rect 2407 2934 2411 2938
rect 2479 2934 2483 2938
rect 2591 2934 2595 2938
rect 2623 2934 2627 2938
rect 2759 2934 2763 2938
rect 2791 2934 2795 2938
rect 2911 2934 2915 2938
rect 2983 2934 2987 2938
rect 3063 2934 3067 2938
rect 3183 2934 3187 2938
rect 3207 2934 3211 2938
rect 3359 2934 3363 2938
rect 3367 2934 3371 2938
rect 3463 2934 3467 2938
rect 111 2866 115 2870
rect 135 2866 139 2870
rect 255 2866 259 2870
rect 327 2866 331 2870
rect 415 2866 419 2870
rect 447 2866 451 2870
rect 575 2866 579 2870
rect 711 2866 715 2870
rect 735 2866 739 2870
rect 847 2866 851 2870
rect 895 2866 899 2870
rect 975 2866 979 2870
rect 1047 2866 1051 2870
rect 1103 2866 1107 2870
rect 1191 2866 1195 2870
rect 1231 2866 1235 2870
rect 1343 2866 1347 2870
rect 1359 2866 1363 2870
rect 1495 2866 1499 2870
rect 1767 2866 1771 2870
rect 1807 2870 1811 2874
rect 1831 2870 1835 2874
rect 1999 2870 2003 2874
rect 2015 2870 2019 2874
rect 2191 2870 2195 2874
rect 2215 2870 2219 2874
rect 2383 2870 2387 2874
rect 2407 2870 2411 2874
rect 2567 2870 2571 2874
rect 2591 2870 2595 2874
rect 2735 2870 2739 2874
rect 2759 2870 2763 2874
rect 2903 2870 2907 2874
rect 2911 2870 2915 2874
rect 3063 2870 3067 2874
rect 3207 2870 3211 2874
rect 3223 2870 3227 2874
rect 3359 2870 3363 2874
rect 3367 2870 3371 2874
rect 3463 2870 3467 2874
rect 1807 2802 1811 2806
rect 1831 2802 1835 2806
rect 1999 2802 2003 2806
rect 2015 2802 2019 2806
rect 2191 2802 2195 2806
rect 2215 2802 2219 2806
rect 2383 2802 2387 2806
rect 2407 2802 2411 2806
rect 2567 2802 2571 2806
rect 2583 2802 2587 2806
rect 2735 2802 2739 2806
rect 2751 2802 2755 2806
rect 2903 2802 2907 2806
rect 2911 2802 2915 2806
rect 3063 2802 3067 2806
rect 3071 2802 3075 2806
rect 3223 2802 3227 2806
rect 3231 2802 3235 2806
rect 3367 2802 3371 2806
rect 3463 2802 3467 2806
rect 111 2790 115 2794
rect 135 2790 139 2794
rect 247 2790 251 2794
rect 255 2790 259 2794
rect 391 2790 395 2794
rect 415 2790 419 2794
rect 543 2790 547 2794
rect 575 2790 579 2794
rect 695 2790 699 2794
rect 735 2790 739 2794
rect 855 2790 859 2794
rect 895 2790 899 2794
rect 1023 2790 1027 2794
rect 1047 2790 1051 2794
rect 1191 2790 1195 2794
rect 1343 2790 1347 2794
rect 1359 2790 1363 2794
rect 1495 2790 1499 2794
rect 1527 2790 1531 2794
rect 1671 2790 1675 2794
rect 1767 2790 1771 2794
rect 111 2718 115 2722
rect 135 2718 139 2722
rect 247 2718 251 2722
rect 359 2718 363 2722
rect 391 2718 395 2722
rect 479 2718 483 2722
rect 543 2718 547 2722
rect 615 2718 619 2722
rect 695 2718 699 2722
rect 759 2718 763 2722
rect 855 2718 859 2722
rect 911 2718 915 2722
rect 1023 2718 1027 2722
rect 1063 2718 1067 2722
rect 1191 2718 1195 2722
rect 1215 2718 1219 2722
rect 1359 2718 1363 2722
rect 1375 2718 1379 2722
rect 1527 2718 1531 2722
rect 1535 2718 1539 2722
rect 1671 2718 1675 2722
rect 1767 2718 1771 2722
rect 1807 2722 1811 2726
rect 1831 2722 1835 2726
rect 2015 2722 2019 2726
rect 2039 2722 2043 2726
rect 2159 2722 2163 2726
rect 2215 2722 2219 2726
rect 2279 2722 2283 2726
rect 2407 2722 2411 2726
rect 2543 2722 2547 2726
rect 2583 2722 2587 2726
rect 2687 2722 2691 2726
rect 2751 2722 2755 2726
rect 2847 2722 2851 2726
rect 2911 2722 2915 2726
rect 3023 2722 3027 2726
rect 3071 2722 3075 2726
rect 3207 2722 3211 2726
rect 3231 2722 3235 2726
rect 3367 2722 3371 2726
rect 3463 2722 3467 2726
rect 111 2646 115 2650
rect 247 2646 251 2650
rect 359 2646 363 2650
rect 463 2646 467 2650
rect 479 2646 483 2650
rect 551 2646 555 2650
rect 615 2646 619 2650
rect 639 2646 643 2650
rect 743 2646 747 2650
rect 759 2646 763 2650
rect 855 2646 859 2650
rect 911 2646 915 2650
rect 983 2646 987 2650
rect 1063 2646 1067 2650
rect 1127 2646 1131 2650
rect 1215 2646 1219 2650
rect 1279 2646 1283 2650
rect 1375 2646 1379 2650
rect 1439 2646 1443 2650
rect 1535 2646 1539 2650
rect 1607 2646 1611 2650
rect 1671 2646 1675 2650
rect 1767 2646 1771 2650
rect 1807 2646 1811 2650
rect 1871 2646 1875 2650
rect 1967 2646 1971 2650
rect 2039 2646 2043 2650
rect 2071 2646 2075 2650
rect 2159 2646 2163 2650
rect 2183 2646 2187 2650
rect 2279 2646 2283 2650
rect 2295 2646 2299 2650
rect 2407 2646 2411 2650
rect 2431 2646 2435 2650
rect 2543 2646 2547 2650
rect 2583 2646 2587 2650
rect 2687 2646 2691 2650
rect 2759 2646 2763 2650
rect 2847 2646 2851 2650
rect 2959 2646 2963 2650
rect 3023 2646 3027 2650
rect 3167 2646 3171 2650
rect 3207 2646 3211 2650
rect 3367 2646 3371 2650
rect 3463 2646 3467 2650
rect 111 2574 115 2578
rect 463 2574 467 2578
rect 503 2574 507 2578
rect 551 2574 555 2578
rect 591 2574 595 2578
rect 639 2574 643 2578
rect 679 2574 683 2578
rect 743 2574 747 2578
rect 775 2574 779 2578
rect 855 2574 859 2578
rect 879 2574 883 2578
rect 983 2574 987 2578
rect 991 2574 995 2578
rect 1103 2574 1107 2578
rect 1127 2574 1131 2578
rect 1223 2574 1227 2578
rect 1279 2574 1283 2578
rect 1351 2574 1355 2578
rect 1439 2574 1443 2578
rect 1479 2574 1483 2578
rect 1607 2574 1611 2578
rect 1767 2574 1771 2578
rect 1807 2570 1811 2574
rect 1831 2570 1835 2574
rect 1871 2570 1875 2574
rect 1919 2570 1923 2574
rect 1967 2570 1971 2574
rect 2007 2570 2011 2574
rect 2071 2570 2075 2574
rect 2111 2570 2115 2574
rect 2183 2570 2187 2574
rect 2223 2570 2227 2574
rect 2295 2570 2299 2574
rect 2343 2570 2347 2574
rect 2431 2570 2435 2574
rect 2487 2570 2491 2574
rect 2583 2570 2587 2574
rect 2647 2570 2651 2574
rect 2759 2570 2763 2574
rect 2815 2570 2819 2574
rect 2959 2570 2963 2574
rect 2999 2570 3003 2574
rect 3167 2570 3171 2574
rect 3191 2570 3195 2574
rect 3367 2570 3371 2574
rect 3463 2570 3467 2574
rect 111 2502 115 2506
rect 503 2502 507 2506
rect 551 2502 555 2506
rect 591 2502 595 2506
rect 679 2502 683 2506
rect 735 2502 739 2506
rect 775 2502 779 2506
rect 879 2502 883 2506
rect 911 2502 915 2506
rect 991 2502 995 2506
rect 1079 2502 1083 2506
rect 1103 2502 1107 2506
rect 1223 2502 1227 2506
rect 1239 2502 1243 2506
rect 1351 2502 1355 2506
rect 1399 2502 1403 2506
rect 1479 2502 1483 2506
rect 1567 2502 1571 2506
rect 1607 2502 1611 2506
rect 1767 2502 1771 2506
rect 1807 2506 1811 2510
rect 1831 2506 1835 2510
rect 1919 2506 1923 2510
rect 1951 2506 1955 2510
rect 2007 2506 2011 2510
rect 2039 2506 2043 2510
rect 2111 2506 2115 2510
rect 2135 2506 2139 2510
rect 2223 2506 2227 2510
rect 2239 2506 2243 2510
rect 2343 2506 2347 2510
rect 2367 2506 2371 2510
rect 2487 2506 2491 2510
rect 2527 2506 2531 2510
rect 2647 2506 2651 2510
rect 2711 2506 2715 2510
rect 2815 2506 2819 2510
rect 2919 2506 2923 2510
rect 2999 2506 3003 2510
rect 3143 2506 3147 2510
rect 3191 2506 3195 2510
rect 3367 2506 3371 2510
rect 3463 2506 3467 2510
rect 111 2438 115 2442
rect 415 2438 419 2442
rect 503 2438 507 2442
rect 551 2438 555 2442
rect 599 2438 603 2442
rect 703 2438 707 2442
rect 735 2438 739 2442
rect 807 2438 811 2442
rect 911 2438 915 2442
rect 919 2438 923 2442
rect 1039 2438 1043 2442
rect 1079 2438 1083 2442
rect 1167 2438 1171 2442
rect 1239 2438 1243 2442
rect 1295 2438 1299 2442
rect 1399 2438 1403 2442
rect 1423 2438 1427 2442
rect 1567 2438 1571 2442
rect 1767 2438 1771 2442
rect 1807 2434 1811 2438
rect 1951 2434 1955 2438
rect 2039 2434 2043 2438
rect 2135 2434 2139 2438
rect 2215 2434 2219 2438
rect 2239 2434 2243 2438
rect 2303 2434 2307 2438
rect 2367 2434 2371 2438
rect 2391 2434 2395 2438
rect 2479 2434 2483 2438
rect 2527 2434 2531 2438
rect 2567 2434 2571 2438
rect 2655 2434 2659 2438
rect 2711 2434 2715 2438
rect 2743 2434 2747 2438
rect 2839 2434 2843 2438
rect 2919 2434 2923 2438
rect 2935 2434 2939 2438
rect 3143 2434 3147 2438
rect 3367 2434 3371 2438
rect 3463 2434 3467 2438
rect 111 2370 115 2374
rect 319 2370 323 2374
rect 415 2370 419 2374
rect 431 2370 435 2374
rect 503 2370 507 2374
rect 543 2370 547 2374
rect 599 2370 603 2374
rect 655 2370 659 2374
rect 703 2370 707 2374
rect 767 2370 771 2374
rect 807 2370 811 2374
rect 879 2370 883 2374
rect 919 2370 923 2374
rect 991 2370 995 2374
rect 1039 2370 1043 2374
rect 1103 2370 1107 2374
rect 1167 2370 1171 2374
rect 1215 2370 1219 2374
rect 1295 2370 1299 2374
rect 1335 2370 1339 2374
rect 1423 2370 1427 2374
rect 1767 2370 1771 2374
rect 1807 2370 1811 2374
rect 2167 2370 2171 2374
rect 2215 2370 2219 2374
rect 2263 2370 2267 2374
rect 2303 2370 2307 2374
rect 2367 2370 2371 2374
rect 2391 2370 2395 2374
rect 2471 2370 2475 2374
rect 2479 2370 2483 2374
rect 2567 2370 2571 2374
rect 2575 2370 2579 2374
rect 2655 2370 2659 2374
rect 2687 2370 2691 2374
rect 2743 2370 2747 2374
rect 2799 2370 2803 2374
rect 2839 2370 2843 2374
rect 2911 2370 2915 2374
rect 2935 2370 2939 2374
rect 3023 2370 3027 2374
rect 3463 2370 3467 2374
rect 111 2298 115 2302
rect 151 2298 155 2302
rect 271 2298 275 2302
rect 319 2298 323 2302
rect 391 2298 395 2302
rect 431 2298 435 2302
rect 519 2298 523 2302
rect 543 2298 547 2302
rect 647 2298 651 2302
rect 655 2298 659 2302
rect 767 2298 771 2302
rect 775 2298 779 2302
rect 879 2298 883 2302
rect 895 2298 899 2302
rect 991 2298 995 2302
rect 1015 2298 1019 2302
rect 1103 2298 1107 2302
rect 1143 2298 1147 2302
rect 1215 2298 1219 2302
rect 1271 2298 1275 2302
rect 1335 2298 1339 2302
rect 1767 2298 1771 2302
rect 1807 2298 1811 2302
rect 1887 2298 1891 2302
rect 2039 2298 2043 2302
rect 2167 2298 2171 2302
rect 2199 2298 2203 2302
rect 2263 2298 2267 2302
rect 2367 2298 2371 2302
rect 2375 2298 2379 2302
rect 2471 2298 2475 2302
rect 2551 2298 2555 2302
rect 2575 2298 2579 2302
rect 2687 2298 2691 2302
rect 2719 2298 2723 2302
rect 2799 2298 2803 2302
rect 2887 2298 2891 2302
rect 2911 2298 2915 2302
rect 3023 2298 3027 2302
rect 3055 2298 3059 2302
rect 3223 2298 3227 2302
rect 3367 2298 3371 2302
rect 3463 2298 3467 2302
rect 111 2230 115 2234
rect 135 2230 139 2234
rect 151 2230 155 2234
rect 247 2230 251 2234
rect 271 2230 275 2234
rect 391 2230 395 2234
rect 407 2230 411 2234
rect 519 2230 523 2234
rect 583 2230 587 2234
rect 647 2230 651 2234
rect 767 2230 771 2234
rect 775 2230 779 2234
rect 895 2230 899 2234
rect 951 2230 955 2234
rect 1015 2230 1019 2234
rect 1135 2230 1139 2234
rect 1143 2230 1147 2234
rect 1271 2230 1275 2234
rect 1319 2230 1323 2234
rect 1503 2230 1507 2234
rect 1671 2230 1675 2234
rect 1767 2230 1771 2234
rect 1807 2234 1811 2238
rect 1831 2234 1835 2238
rect 1887 2234 1891 2238
rect 1967 2234 1971 2238
rect 2039 2234 2043 2238
rect 2135 2234 2139 2238
rect 2199 2234 2203 2238
rect 2311 2234 2315 2238
rect 2375 2234 2379 2238
rect 2487 2234 2491 2238
rect 2551 2234 2555 2238
rect 2655 2234 2659 2238
rect 2719 2234 2723 2238
rect 2815 2234 2819 2238
rect 2887 2234 2891 2238
rect 2959 2234 2963 2238
rect 3055 2234 3059 2238
rect 3103 2234 3107 2238
rect 3223 2234 3227 2238
rect 3247 2234 3251 2238
rect 3367 2234 3371 2238
rect 3463 2234 3467 2238
rect 1807 2170 1811 2174
rect 1831 2170 1835 2174
rect 1967 2170 1971 2174
rect 2135 2170 2139 2174
rect 2311 2170 2315 2174
rect 2487 2170 2491 2174
rect 2655 2170 2659 2174
rect 2815 2170 2819 2174
rect 2927 2170 2931 2174
rect 2959 2170 2963 2174
rect 3015 2170 3019 2174
rect 3103 2170 3107 2174
rect 3191 2170 3195 2174
rect 3247 2170 3251 2174
rect 3279 2170 3283 2174
rect 3367 2170 3371 2174
rect 3463 2170 3467 2174
rect 111 2158 115 2162
rect 135 2158 139 2162
rect 247 2158 251 2162
rect 391 2158 395 2162
rect 407 2158 411 2162
rect 543 2158 547 2162
rect 583 2158 587 2162
rect 695 2158 699 2162
rect 767 2158 771 2162
rect 839 2158 843 2162
rect 951 2158 955 2162
rect 975 2158 979 2162
rect 1103 2158 1107 2162
rect 1135 2158 1139 2162
rect 1231 2158 1235 2162
rect 1319 2158 1323 2162
rect 1351 2158 1355 2162
rect 1463 2158 1467 2162
rect 1503 2158 1507 2162
rect 1575 2158 1579 2162
rect 1671 2158 1675 2162
rect 1767 2158 1771 2162
rect 1807 2098 1811 2102
rect 1831 2098 1835 2102
rect 1991 2098 1995 2102
rect 2167 2098 2171 2102
rect 2343 2098 2347 2102
rect 2503 2098 2507 2102
rect 2655 2098 2659 2102
rect 2791 2098 2795 2102
rect 2919 2098 2923 2102
rect 2927 2098 2931 2102
rect 3015 2098 3019 2102
rect 3039 2098 3043 2102
rect 3103 2098 3107 2102
rect 3159 2098 3163 2102
rect 3191 2098 3195 2102
rect 3271 2098 3275 2102
rect 3279 2098 3283 2102
rect 3367 2098 3371 2102
rect 3463 2098 3467 2102
rect 111 2090 115 2094
rect 135 2090 139 2094
rect 223 2090 227 2094
rect 247 2090 251 2094
rect 343 2090 347 2094
rect 391 2090 395 2094
rect 463 2090 467 2094
rect 543 2090 547 2094
rect 583 2090 587 2094
rect 695 2090 699 2094
rect 703 2090 707 2094
rect 823 2090 827 2094
rect 839 2090 843 2094
rect 935 2090 939 2094
rect 975 2090 979 2094
rect 1047 2090 1051 2094
rect 1103 2090 1107 2094
rect 1159 2090 1163 2094
rect 1231 2090 1235 2094
rect 1279 2090 1283 2094
rect 1351 2090 1355 2094
rect 1463 2090 1467 2094
rect 1575 2090 1579 2094
rect 1671 2090 1675 2094
rect 1767 2090 1771 2094
rect 1807 2030 1811 2034
rect 1831 2030 1835 2034
rect 1991 2030 1995 2034
rect 2015 2030 2019 2034
rect 2167 2030 2171 2034
rect 2223 2030 2227 2034
rect 2343 2030 2347 2034
rect 2431 2030 2435 2034
rect 2503 2030 2507 2034
rect 2631 2030 2635 2034
rect 2655 2030 2659 2034
rect 2791 2030 2795 2034
rect 2823 2030 2827 2034
rect 2919 2030 2923 2034
rect 3007 2030 3011 2034
rect 3039 2030 3043 2034
rect 3159 2030 3163 2034
rect 3199 2030 3203 2034
rect 3271 2030 3275 2034
rect 3367 2030 3371 2034
rect 3463 2030 3467 2034
rect 111 2018 115 2022
rect 135 2018 139 2022
rect 223 2018 227 2022
rect 239 2018 243 2022
rect 343 2018 347 2022
rect 367 2018 371 2022
rect 463 2018 467 2022
rect 503 2018 507 2022
rect 583 2018 587 2022
rect 639 2018 643 2022
rect 703 2018 707 2022
rect 775 2018 779 2022
rect 823 2018 827 2022
rect 911 2018 915 2022
rect 935 2018 939 2022
rect 1047 2018 1051 2022
rect 1159 2018 1163 2022
rect 1183 2018 1187 2022
rect 1279 2018 1283 2022
rect 1327 2018 1331 2022
rect 1767 2018 1771 2022
rect 1807 1962 1811 1966
rect 1831 1962 1835 1966
rect 1863 1962 1867 1966
rect 1999 1962 2003 1966
rect 2015 1962 2019 1966
rect 2143 1962 2147 1966
rect 2223 1962 2227 1966
rect 2287 1962 2291 1966
rect 2431 1962 2435 1966
rect 2575 1962 2579 1966
rect 2631 1962 2635 1966
rect 2711 1962 2715 1966
rect 2823 1962 2827 1966
rect 2831 1962 2835 1966
rect 2951 1962 2955 1966
rect 3007 1962 3011 1966
rect 3063 1962 3067 1966
rect 3167 1962 3171 1966
rect 3199 1962 3203 1966
rect 3279 1962 3283 1966
rect 3367 1962 3371 1966
rect 3463 1962 3467 1966
rect 111 1950 115 1954
rect 135 1950 139 1954
rect 239 1950 243 1954
rect 295 1950 299 1954
rect 367 1950 371 1954
rect 423 1950 427 1954
rect 503 1950 507 1954
rect 559 1950 563 1954
rect 639 1950 643 1954
rect 703 1950 707 1954
rect 775 1950 779 1954
rect 855 1950 859 1954
rect 911 1950 915 1954
rect 1007 1950 1011 1954
rect 1047 1950 1051 1954
rect 1159 1950 1163 1954
rect 1183 1950 1187 1954
rect 1311 1950 1315 1954
rect 1327 1950 1331 1954
rect 1471 1950 1475 1954
rect 1767 1950 1771 1954
rect 1807 1894 1811 1898
rect 1863 1894 1867 1898
rect 1999 1894 2003 1898
rect 2015 1894 2019 1898
rect 2111 1894 2115 1898
rect 2143 1894 2147 1898
rect 2215 1894 2219 1898
rect 2287 1894 2291 1898
rect 2327 1894 2331 1898
rect 2431 1894 2435 1898
rect 2439 1894 2443 1898
rect 2543 1894 2547 1898
rect 2575 1894 2579 1898
rect 2647 1894 2651 1898
rect 2711 1894 2715 1898
rect 2759 1894 2763 1898
rect 2831 1894 2835 1898
rect 2871 1894 2875 1898
rect 2951 1894 2955 1898
rect 2983 1894 2987 1898
rect 3063 1894 3067 1898
rect 3167 1894 3171 1898
rect 3279 1894 3283 1898
rect 3367 1894 3371 1898
rect 3463 1894 3467 1898
rect 111 1886 115 1890
rect 295 1886 299 1890
rect 423 1886 427 1890
rect 431 1886 435 1890
rect 559 1886 563 1890
rect 575 1886 579 1890
rect 703 1886 707 1890
rect 727 1886 731 1890
rect 855 1886 859 1890
rect 887 1886 891 1890
rect 1007 1886 1011 1890
rect 1047 1886 1051 1890
rect 1159 1886 1163 1890
rect 1199 1886 1203 1890
rect 1311 1886 1315 1890
rect 1351 1886 1355 1890
rect 1471 1886 1475 1890
rect 1511 1886 1515 1890
rect 1671 1886 1675 1890
rect 1767 1886 1771 1890
rect 111 1818 115 1822
rect 431 1818 435 1822
rect 511 1818 515 1822
rect 575 1818 579 1822
rect 631 1818 635 1822
rect 727 1818 731 1822
rect 759 1818 763 1822
rect 887 1818 891 1822
rect 1023 1818 1027 1822
rect 1047 1818 1051 1822
rect 1151 1818 1155 1822
rect 1199 1818 1203 1822
rect 1279 1818 1283 1822
rect 1351 1818 1355 1822
rect 1407 1818 1411 1822
rect 1511 1818 1515 1822
rect 1535 1818 1539 1822
rect 1671 1818 1675 1822
rect 1767 1818 1771 1822
rect 1807 1822 1811 1826
rect 2015 1822 2019 1826
rect 2103 1822 2107 1826
rect 2111 1822 2115 1826
rect 2191 1822 2195 1826
rect 2215 1822 2219 1826
rect 2279 1822 2283 1826
rect 2327 1822 2331 1826
rect 2367 1822 2371 1826
rect 2439 1822 2443 1826
rect 2455 1822 2459 1826
rect 2543 1822 2547 1826
rect 2631 1822 2635 1826
rect 2647 1822 2651 1826
rect 2719 1822 2723 1826
rect 2759 1822 2763 1826
rect 2807 1822 2811 1826
rect 2871 1822 2875 1826
rect 2895 1822 2899 1826
rect 2983 1822 2987 1826
rect 3463 1822 3467 1826
rect 111 1750 115 1754
rect 439 1750 443 1754
rect 511 1750 515 1754
rect 535 1750 539 1754
rect 631 1750 635 1754
rect 639 1750 643 1754
rect 743 1750 747 1754
rect 759 1750 763 1754
rect 847 1750 851 1754
rect 887 1750 891 1754
rect 951 1750 955 1754
rect 1023 1750 1027 1754
rect 1055 1750 1059 1754
rect 1151 1750 1155 1754
rect 1159 1750 1163 1754
rect 1271 1750 1275 1754
rect 1279 1750 1283 1754
rect 1383 1750 1387 1754
rect 1407 1750 1411 1754
rect 1535 1750 1539 1754
rect 1671 1750 1675 1754
rect 1767 1750 1771 1754
rect 1807 1746 1811 1750
rect 2103 1746 2107 1750
rect 2143 1746 2147 1750
rect 2191 1746 2195 1750
rect 2231 1746 2235 1750
rect 2279 1746 2283 1750
rect 2319 1746 2323 1750
rect 2367 1746 2371 1750
rect 2407 1746 2411 1750
rect 2455 1746 2459 1750
rect 2495 1746 2499 1750
rect 2543 1746 2547 1750
rect 2583 1746 2587 1750
rect 2631 1746 2635 1750
rect 2671 1746 2675 1750
rect 2719 1746 2723 1750
rect 2759 1746 2763 1750
rect 2807 1746 2811 1750
rect 2847 1746 2851 1750
rect 2895 1746 2899 1750
rect 3463 1746 3467 1750
rect 111 1682 115 1686
rect 399 1682 403 1686
rect 439 1682 443 1686
rect 487 1682 491 1686
rect 535 1682 539 1686
rect 575 1682 579 1686
rect 639 1682 643 1686
rect 663 1682 667 1686
rect 743 1682 747 1686
rect 759 1682 763 1686
rect 847 1682 851 1686
rect 855 1682 859 1686
rect 951 1682 955 1686
rect 1047 1682 1051 1686
rect 1055 1682 1059 1686
rect 1143 1682 1147 1686
rect 1159 1682 1163 1686
rect 1271 1682 1275 1686
rect 1383 1682 1387 1686
rect 1767 1682 1771 1686
rect 1807 1678 1811 1682
rect 2103 1678 2107 1682
rect 2143 1678 2147 1682
rect 2191 1678 2195 1682
rect 2231 1678 2235 1682
rect 2279 1678 2283 1682
rect 2319 1678 2323 1682
rect 2367 1678 2371 1682
rect 2407 1678 2411 1682
rect 2455 1678 2459 1682
rect 2495 1678 2499 1682
rect 2543 1678 2547 1682
rect 2583 1678 2587 1682
rect 2631 1678 2635 1682
rect 2671 1678 2675 1682
rect 2719 1678 2723 1682
rect 2759 1678 2763 1682
rect 2807 1678 2811 1682
rect 2847 1678 2851 1682
rect 2895 1678 2899 1682
rect 3463 1678 3467 1682
rect 111 1614 115 1618
rect 279 1614 283 1618
rect 383 1614 387 1618
rect 399 1614 403 1618
rect 487 1614 491 1618
rect 495 1614 499 1618
rect 575 1614 579 1618
rect 607 1614 611 1618
rect 663 1614 667 1618
rect 719 1614 723 1618
rect 759 1614 763 1618
rect 831 1614 835 1618
rect 855 1614 859 1618
rect 943 1614 947 1618
rect 951 1614 955 1618
rect 1047 1614 1051 1618
rect 1055 1614 1059 1618
rect 1143 1614 1147 1618
rect 1167 1614 1171 1618
rect 1279 1614 1283 1618
rect 1767 1614 1771 1618
rect 1807 1610 1811 1614
rect 2063 1610 2067 1614
rect 2103 1610 2107 1614
rect 2159 1610 2163 1614
rect 2191 1610 2195 1614
rect 2255 1610 2259 1614
rect 2279 1610 2283 1614
rect 2359 1610 2363 1614
rect 2367 1610 2371 1614
rect 2455 1610 2459 1614
rect 2463 1610 2467 1614
rect 2543 1610 2547 1614
rect 2567 1610 2571 1614
rect 2631 1610 2635 1614
rect 2671 1610 2675 1614
rect 2719 1610 2723 1614
rect 2775 1610 2779 1614
rect 2807 1610 2811 1614
rect 2887 1610 2891 1614
rect 2895 1610 2899 1614
rect 3463 1610 3467 1614
rect 111 1542 115 1546
rect 183 1542 187 1546
rect 279 1542 283 1546
rect 327 1542 331 1546
rect 383 1542 387 1546
rect 471 1542 475 1546
rect 495 1542 499 1546
rect 607 1542 611 1546
rect 623 1542 627 1546
rect 719 1542 723 1546
rect 767 1542 771 1546
rect 831 1542 835 1546
rect 911 1542 915 1546
rect 943 1542 947 1546
rect 1047 1542 1051 1546
rect 1055 1542 1059 1546
rect 1167 1542 1171 1546
rect 1175 1542 1179 1546
rect 1279 1542 1283 1546
rect 1311 1542 1315 1546
rect 1447 1542 1451 1546
rect 1767 1542 1771 1546
rect 1807 1546 1811 1550
rect 1919 1546 1923 1550
rect 2039 1546 2043 1550
rect 2063 1546 2067 1550
rect 2159 1546 2163 1550
rect 2167 1546 2171 1550
rect 2255 1546 2259 1550
rect 2295 1546 2299 1550
rect 2359 1546 2363 1550
rect 2423 1546 2427 1550
rect 2463 1546 2467 1550
rect 2551 1546 2555 1550
rect 2567 1546 2571 1550
rect 2671 1546 2675 1550
rect 2679 1546 2683 1550
rect 2775 1546 2779 1550
rect 2799 1546 2803 1550
rect 2887 1546 2891 1550
rect 2927 1546 2931 1550
rect 3055 1546 3059 1550
rect 3463 1546 3467 1550
rect 111 1474 115 1478
rect 159 1474 163 1478
rect 183 1474 187 1478
rect 327 1474 331 1478
rect 375 1474 379 1478
rect 471 1474 475 1478
rect 583 1474 587 1478
rect 623 1474 627 1478
rect 767 1474 771 1478
rect 783 1474 787 1478
rect 911 1474 915 1478
rect 959 1474 963 1478
rect 1047 1474 1051 1478
rect 1127 1474 1131 1478
rect 1175 1474 1179 1478
rect 1279 1474 1283 1478
rect 1311 1474 1315 1478
rect 1431 1474 1435 1478
rect 1447 1474 1451 1478
rect 1591 1474 1595 1478
rect 1767 1474 1771 1478
rect 1807 1474 1811 1478
rect 1831 1474 1835 1478
rect 1919 1474 1923 1478
rect 1951 1474 1955 1478
rect 2039 1474 2043 1478
rect 2111 1474 2115 1478
rect 2167 1474 2171 1478
rect 2271 1474 2275 1478
rect 2295 1474 2299 1478
rect 2423 1474 2427 1478
rect 2431 1474 2435 1478
rect 2551 1474 2555 1478
rect 2591 1474 2595 1478
rect 2679 1474 2683 1478
rect 2735 1474 2739 1478
rect 2799 1474 2803 1478
rect 2871 1474 2875 1478
rect 2927 1474 2931 1478
rect 3007 1474 3011 1478
rect 3055 1474 3059 1478
rect 3135 1474 3139 1478
rect 3263 1474 3267 1478
rect 3367 1474 3371 1478
rect 3463 1474 3467 1478
rect 111 1406 115 1410
rect 135 1406 139 1410
rect 159 1406 163 1410
rect 303 1406 307 1410
rect 375 1406 379 1410
rect 495 1406 499 1410
rect 583 1406 587 1410
rect 679 1406 683 1410
rect 783 1406 787 1410
rect 855 1406 859 1410
rect 959 1406 963 1410
rect 1015 1406 1019 1410
rect 1127 1406 1131 1410
rect 1167 1406 1171 1410
rect 1279 1406 1283 1410
rect 1303 1406 1307 1410
rect 1431 1406 1435 1410
rect 1559 1406 1563 1410
rect 1591 1406 1595 1410
rect 1671 1406 1675 1410
rect 1767 1406 1771 1410
rect 1807 1406 1811 1410
rect 1831 1406 1835 1410
rect 1951 1406 1955 1410
rect 2007 1406 2011 1410
rect 2111 1406 2115 1410
rect 2199 1406 2203 1410
rect 2271 1406 2275 1410
rect 2383 1406 2387 1410
rect 2431 1406 2435 1410
rect 2559 1406 2563 1410
rect 2591 1406 2595 1410
rect 2719 1406 2723 1410
rect 2735 1406 2739 1410
rect 2863 1406 2867 1410
rect 2871 1406 2875 1410
rect 2999 1406 3003 1410
rect 3007 1406 3011 1410
rect 3127 1406 3131 1410
rect 3135 1406 3139 1410
rect 3255 1406 3259 1410
rect 3263 1406 3267 1410
rect 3367 1406 3371 1410
rect 3463 1406 3467 1410
rect 111 1338 115 1342
rect 135 1338 139 1342
rect 247 1338 251 1342
rect 303 1338 307 1342
rect 399 1338 403 1342
rect 495 1338 499 1342
rect 559 1338 563 1342
rect 679 1338 683 1342
rect 727 1338 731 1342
rect 855 1338 859 1342
rect 895 1338 899 1342
rect 1015 1338 1019 1342
rect 1063 1338 1067 1342
rect 1167 1338 1171 1342
rect 1223 1338 1227 1342
rect 1303 1338 1307 1342
rect 1375 1338 1379 1342
rect 1431 1338 1435 1342
rect 1535 1338 1539 1342
rect 1559 1338 1563 1342
rect 1671 1338 1675 1342
rect 1767 1338 1771 1342
rect 1807 1334 1811 1338
rect 1831 1334 1835 1338
rect 1967 1334 1971 1338
rect 2007 1334 2011 1338
rect 2143 1334 2147 1338
rect 2199 1334 2203 1338
rect 2327 1334 2331 1338
rect 2383 1334 2387 1338
rect 2511 1334 2515 1338
rect 2559 1334 2563 1338
rect 2687 1334 2691 1338
rect 2719 1334 2723 1338
rect 2863 1334 2867 1338
rect 2999 1334 3003 1338
rect 3039 1334 3043 1338
rect 3127 1334 3131 1338
rect 3215 1334 3219 1338
rect 3255 1334 3259 1338
rect 3367 1334 3371 1338
rect 3463 1334 3467 1338
rect 111 1270 115 1274
rect 135 1270 139 1274
rect 223 1270 227 1274
rect 247 1270 251 1274
rect 319 1270 323 1274
rect 399 1270 403 1274
rect 431 1270 435 1274
rect 551 1270 555 1274
rect 559 1270 563 1274
rect 679 1270 683 1274
rect 727 1270 731 1274
rect 823 1270 827 1274
rect 895 1270 899 1274
rect 975 1270 979 1274
rect 1063 1270 1067 1274
rect 1143 1270 1147 1274
rect 1223 1270 1227 1274
rect 1319 1270 1323 1274
rect 1375 1270 1379 1274
rect 1503 1270 1507 1274
rect 1535 1270 1539 1274
rect 1671 1270 1675 1274
rect 1767 1270 1771 1274
rect 1807 1270 1811 1274
rect 1831 1270 1835 1274
rect 1967 1270 1971 1274
rect 2095 1270 2099 1274
rect 2143 1270 2147 1274
rect 2327 1270 2331 1274
rect 2359 1270 2363 1274
rect 2511 1270 2515 1274
rect 2599 1270 2603 1274
rect 2687 1270 2691 1274
rect 2807 1270 2811 1274
rect 2863 1270 2867 1274
rect 3007 1270 3011 1274
rect 3039 1270 3043 1274
rect 3199 1270 3203 1274
rect 3215 1270 3219 1274
rect 3367 1270 3371 1274
rect 3463 1270 3467 1274
rect 111 1198 115 1202
rect 135 1198 139 1202
rect 223 1198 227 1202
rect 231 1198 235 1202
rect 319 1198 323 1202
rect 359 1198 363 1202
rect 431 1198 435 1202
rect 487 1198 491 1202
rect 551 1198 555 1202
rect 615 1198 619 1202
rect 679 1198 683 1202
rect 743 1198 747 1202
rect 823 1198 827 1202
rect 871 1198 875 1202
rect 975 1198 979 1202
rect 991 1198 995 1202
rect 1119 1198 1123 1202
rect 1143 1198 1147 1202
rect 1247 1198 1251 1202
rect 1319 1198 1323 1202
rect 1503 1198 1507 1202
rect 1671 1198 1675 1202
rect 1767 1198 1771 1202
rect 1807 1198 1811 1202
rect 1831 1198 1835 1202
rect 1935 1198 1939 1202
rect 2039 1198 2043 1202
rect 2095 1198 2099 1202
rect 2159 1198 2163 1202
rect 2287 1198 2291 1202
rect 2359 1198 2363 1202
rect 2423 1198 2427 1202
rect 2567 1198 2571 1202
rect 2599 1198 2603 1202
rect 2703 1198 2707 1202
rect 2807 1198 2811 1202
rect 2839 1198 2843 1202
rect 2975 1198 2979 1202
rect 3007 1198 3011 1202
rect 3111 1198 3115 1202
rect 3199 1198 3203 1202
rect 3247 1198 3251 1202
rect 3367 1198 3371 1202
rect 3463 1198 3467 1202
rect 111 1130 115 1134
rect 135 1130 139 1134
rect 231 1130 235 1134
rect 247 1130 251 1134
rect 359 1130 363 1134
rect 367 1130 371 1134
rect 487 1130 491 1134
rect 495 1130 499 1134
rect 615 1130 619 1134
rect 623 1130 627 1134
rect 743 1130 747 1134
rect 759 1130 763 1134
rect 871 1130 875 1134
rect 887 1130 891 1134
rect 991 1130 995 1134
rect 1015 1130 1019 1134
rect 1119 1130 1123 1134
rect 1143 1130 1147 1134
rect 1247 1130 1251 1134
rect 1271 1130 1275 1134
rect 1399 1130 1403 1134
rect 1767 1130 1771 1134
rect 1807 1126 1811 1130
rect 1935 1126 1939 1130
rect 1943 1126 1947 1130
rect 2039 1126 2043 1130
rect 2063 1126 2067 1130
rect 2159 1126 2163 1130
rect 2191 1126 2195 1130
rect 2287 1126 2291 1130
rect 2319 1126 2323 1130
rect 2423 1126 2427 1130
rect 2455 1126 2459 1130
rect 2567 1126 2571 1130
rect 2599 1126 2603 1130
rect 2703 1126 2707 1130
rect 2751 1126 2755 1130
rect 2839 1126 2843 1130
rect 2903 1126 2907 1130
rect 2975 1126 2979 1130
rect 3063 1126 3067 1130
rect 3111 1126 3115 1130
rect 3223 1126 3227 1130
rect 3247 1126 3251 1130
rect 3367 1126 3371 1130
rect 3463 1126 3467 1130
rect 111 1062 115 1066
rect 247 1062 251 1066
rect 367 1062 371 1066
rect 431 1062 435 1066
rect 495 1062 499 1066
rect 543 1062 547 1066
rect 623 1062 627 1066
rect 663 1062 667 1066
rect 759 1062 763 1066
rect 791 1062 795 1066
rect 887 1062 891 1066
rect 919 1062 923 1066
rect 1015 1062 1019 1066
rect 1039 1062 1043 1066
rect 1143 1062 1147 1066
rect 1159 1062 1163 1066
rect 1271 1062 1275 1066
rect 1279 1062 1283 1066
rect 1399 1062 1403 1066
rect 1407 1062 1411 1066
rect 1535 1062 1539 1066
rect 1767 1062 1771 1066
rect 1807 1058 1811 1062
rect 1847 1058 1851 1062
rect 1943 1058 1947 1062
rect 1983 1058 1987 1062
rect 2063 1058 2067 1062
rect 2119 1058 2123 1062
rect 2191 1058 2195 1062
rect 2255 1058 2259 1062
rect 2319 1058 2323 1062
rect 2391 1058 2395 1062
rect 2455 1058 2459 1062
rect 2543 1058 2547 1062
rect 2599 1058 2603 1062
rect 2703 1058 2707 1062
rect 2751 1058 2755 1062
rect 2863 1058 2867 1062
rect 2903 1058 2907 1062
rect 3031 1058 3035 1062
rect 3063 1058 3067 1062
rect 3207 1058 3211 1062
rect 3223 1058 3227 1062
rect 3367 1058 3371 1062
rect 3463 1058 3467 1062
rect 111 990 115 994
rect 431 990 435 994
rect 543 990 547 994
rect 567 990 571 994
rect 663 990 667 994
rect 679 990 683 994
rect 791 990 795 994
rect 911 990 915 994
rect 919 990 923 994
rect 1031 990 1035 994
rect 1039 990 1043 994
rect 1143 990 1147 994
rect 1159 990 1163 994
rect 1255 990 1259 994
rect 1279 990 1283 994
rect 1359 990 1363 994
rect 1407 990 1411 994
rect 1471 990 1475 994
rect 1535 990 1539 994
rect 1583 990 1587 994
rect 1671 990 1675 994
rect 1767 990 1771 994
rect 1807 990 1811 994
rect 1831 990 1835 994
rect 1847 990 1851 994
rect 1975 990 1979 994
rect 1983 990 1987 994
rect 2119 990 2123 994
rect 2135 990 2139 994
rect 2255 990 2259 994
rect 2295 990 2299 994
rect 2391 990 2395 994
rect 2463 990 2467 994
rect 2543 990 2547 994
rect 2631 990 2635 994
rect 2703 990 2707 994
rect 2807 990 2811 994
rect 2863 990 2867 994
rect 2991 990 2995 994
rect 3031 990 3035 994
rect 3183 990 3187 994
rect 3207 990 3211 994
rect 3367 990 3371 994
rect 3463 990 3467 994
rect 111 922 115 926
rect 415 922 419 926
rect 559 922 563 926
rect 567 922 571 926
rect 679 922 683 926
rect 727 922 731 926
rect 791 922 795 926
rect 911 922 915 926
rect 1031 922 1035 926
rect 1119 922 1123 926
rect 1143 922 1147 926
rect 1255 922 1259 926
rect 1335 922 1339 926
rect 1359 922 1363 926
rect 1471 922 1475 926
rect 1559 922 1563 926
rect 1583 922 1587 926
rect 1671 922 1675 926
rect 1767 922 1771 926
rect 1807 926 1811 930
rect 1831 926 1835 930
rect 1975 926 1979 930
rect 2127 926 2131 930
rect 2135 926 2139 930
rect 2215 926 2219 930
rect 2295 926 2299 930
rect 2303 926 2307 930
rect 2391 926 2395 930
rect 2463 926 2467 930
rect 2479 926 2483 930
rect 2567 926 2571 930
rect 2631 926 2635 930
rect 2655 926 2659 930
rect 2743 926 2747 930
rect 2807 926 2811 930
rect 2831 926 2835 930
rect 2991 926 2995 930
rect 3183 926 3187 930
rect 3367 926 3371 930
rect 3463 926 3467 930
rect 111 854 115 858
rect 135 854 139 858
rect 231 854 235 858
rect 359 854 363 858
rect 415 854 419 858
rect 487 854 491 858
rect 559 854 563 858
rect 623 854 627 858
rect 727 854 731 858
rect 751 854 755 858
rect 879 854 883 858
rect 911 854 915 858
rect 1007 854 1011 858
rect 1119 854 1123 858
rect 1135 854 1139 858
rect 1271 854 1275 858
rect 1335 854 1339 858
rect 1559 854 1563 858
rect 1767 854 1771 858
rect 1807 854 1811 858
rect 2127 854 2131 858
rect 2159 854 2163 858
rect 2215 854 2219 858
rect 2247 854 2251 858
rect 2303 854 2307 858
rect 2335 854 2339 858
rect 2391 854 2395 858
rect 2423 854 2427 858
rect 2479 854 2483 858
rect 2527 854 2531 858
rect 2567 854 2571 858
rect 2639 854 2643 858
rect 2655 854 2659 858
rect 2743 854 2747 858
rect 2767 854 2771 858
rect 2831 854 2835 858
rect 2911 854 2915 858
rect 3063 854 3067 858
rect 3223 854 3227 858
rect 3367 854 3371 858
rect 3463 854 3467 858
rect 111 786 115 790
rect 135 786 139 790
rect 223 786 227 790
rect 231 786 235 790
rect 343 786 347 790
rect 359 786 363 790
rect 471 786 475 790
rect 487 786 491 790
rect 607 786 611 790
rect 623 786 627 790
rect 743 786 747 790
rect 751 786 755 790
rect 879 786 883 790
rect 887 786 891 790
rect 1007 786 1011 790
rect 1039 786 1043 790
rect 1135 786 1139 790
rect 1191 786 1195 790
rect 1271 786 1275 790
rect 1351 786 1355 790
rect 1767 786 1771 790
rect 1807 786 1811 790
rect 2063 786 2067 790
rect 2159 786 2163 790
rect 2175 786 2179 790
rect 2247 786 2251 790
rect 2295 786 2299 790
rect 2335 786 2339 790
rect 2423 786 2427 790
rect 2527 786 2531 790
rect 2559 786 2563 790
rect 2639 786 2643 790
rect 2711 786 2715 790
rect 2767 786 2771 790
rect 2871 786 2875 790
rect 2911 786 2915 790
rect 3039 786 3043 790
rect 3063 786 3067 790
rect 3215 786 3219 790
rect 3223 786 3227 790
rect 3367 786 3371 790
rect 3463 786 3467 790
rect 111 718 115 722
rect 135 718 139 722
rect 167 718 171 722
rect 223 718 227 722
rect 295 718 299 722
rect 343 718 347 722
rect 431 718 435 722
rect 471 718 475 722
rect 575 718 579 722
rect 607 718 611 722
rect 727 718 731 722
rect 743 718 747 722
rect 879 718 883 722
rect 887 718 891 722
rect 1031 718 1035 722
rect 1039 718 1043 722
rect 1183 718 1187 722
rect 1191 718 1195 722
rect 1343 718 1347 722
rect 1351 718 1355 722
rect 1503 718 1507 722
rect 1767 718 1771 722
rect 1807 722 1811 726
rect 1927 722 1931 726
rect 2063 722 2067 726
rect 2071 722 2075 726
rect 2175 722 2179 726
rect 2231 722 2235 726
rect 2295 722 2299 726
rect 2391 722 2395 726
rect 2423 722 2427 726
rect 2551 722 2555 726
rect 2559 722 2563 726
rect 2703 722 2707 726
rect 2711 722 2715 726
rect 2847 722 2851 726
rect 2871 722 2875 726
rect 2983 722 2987 726
rect 3039 722 3043 726
rect 3119 722 3123 726
rect 3215 722 3219 726
rect 3255 722 3259 726
rect 3367 722 3371 726
rect 3463 722 3467 726
rect 111 650 115 654
rect 167 650 171 654
rect 295 650 299 654
rect 431 650 435 654
rect 455 650 459 654
rect 559 650 563 654
rect 575 650 579 654
rect 679 650 683 654
rect 727 650 731 654
rect 799 650 803 654
rect 879 650 883 654
rect 927 650 931 654
rect 1031 650 1035 654
rect 1055 650 1059 654
rect 1183 650 1187 654
rect 1311 650 1315 654
rect 1343 650 1347 654
rect 1447 650 1451 654
rect 1503 650 1507 654
rect 1583 650 1587 654
rect 1767 650 1771 654
rect 1807 650 1811 654
rect 1831 650 1835 654
rect 1927 650 1931 654
rect 1967 650 1971 654
rect 2071 650 2075 654
rect 2135 650 2139 654
rect 2231 650 2235 654
rect 2311 650 2315 654
rect 2391 650 2395 654
rect 2487 650 2491 654
rect 2551 650 2555 654
rect 2655 650 2659 654
rect 2703 650 2707 654
rect 2815 650 2819 654
rect 2847 650 2851 654
rect 2959 650 2963 654
rect 2983 650 2987 654
rect 3103 650 3107 654
rect 3119 650 3123 654
rect 3247 650 3251 654
rect 3255 650 3259 654
rect 3367 650 3371 654
rect 3463 650 3467 654
rect 1807 586 1811 590
rect 1831 586 1835 590
rect 1967 586 1971 590
rect 2127 586 2131 590
rect 2135 586 2139 590
rect 2287 586 2291 590
rect 2311 586 2315 590
rect 2455 586 2459 590
rect 2487 586 2491 590
rect 2623 586 2627 590
rect 2655 586 2659 590
rect 2799 586 2803 590
rect 2815 586 2819 590
rect 2959 586 2963 590
rect 2983 586 2987 590
rect 3103 586 3107 590
rect 3167 586 3171 590
rect 3247 586 3251 590
rect 3359 586 3363 590
rect 3367 586 3371 590
rect 3463 586 3467 590
rect 111 578 115 582
rect 455 578 459 582
rect 559 578 563 582
rect 599 578 603 582
rect 679 578 683 582
rect 703 578 707 582
rect 799 578 803 582
rect 815 578 819 582
rect 927 578 931 582
rect 1039 578 1043 582
rect 1055 578 1059 582
rect 1151 578 1155 582
rect 1183 578 1187 582
rect 1255 578 1259 582
rect 1311 578 1315 582
rect 1359 578 1363 582
rect 1447 578 1451 582
rect 1471 578 1475 582
rect 1583 578 1587 582
rect 1671 578 1675 582
rect 1767 578 1771 582
rect 111 514 115 518
rect 303 514 307 518
rect 431 514 435 518
rect 567 514 571 518
rect 599 514 603 518
rect 703 514 707 518
rect 815 514 819 518
rect 847 514 851 518
rect 927 514 931 518
rect 983 514 987 518
rect 1039 514 1043 518
rect 1111 514 1115 518
rect 1151 514 1155 518
rect 1231 514 1235 518
rect 1255 514 1259 518
rect 1351 514 1355 518
rect 1359 514 1363 518
rect 1463 514 1467 518
rect 1471 514 1475 518
rect 1575 514 1579 518
rect 1583 514 1587 518
rect 1671 514 1675 518
rect 1767 514 1771 518
rect 1807 506 1811 510
rect 1831 506 1835 510
rect 1967 506 1971 510
rect 2127 506 2131 510
rect 2287 506 2291 510
rect 2295 506 2299 510
rect 2455 506 2459 510
rect 2479 506 2483 510
rect 2623 506 2627 510
rect 2679 506 2683 510
rect 2799 506 2803 510
rect 2887 506 2891 510
rect 2983 506 2987 510
rect 3111 506 3115 510
rect 3167 506 3171 510
rect 3335 506 3339 510
rect 3359 506 3363 510
rect 3463 506 3467 510
rect 111 442 115 446
rect 135 442 139 446
rect 255 442 259 446
rect 303 442 307 446
rect 415 442 419 446
rect 431 442 435 446
rect 567 442 571 446
rect 583 442 587 446
rect 703 442 707 446
rect 743 442 747 446
rect 847 442 851 446
rect 903 442 907 446
rect 983 442 987 446
rect 1047 442 1051 446
rect 1111 442 1115 446
rect 1183 442 1187 446
rect 1231 442 1235 446
rect 1311 442 1315 446
rect 1351 442 1355 446
rect 1439 442 1443 446
rect 1463 442 1467 446
rect 1567 442 1571 446
rect 1575 442 1579 446
rect 1671 442 1675 446
rect 1767 442 1771 446
rect 1807 442 1811 446
rect 1831 442 1835 446
rect 1959 442 1963 446
rect 1967 442 1971 446
rect 2111 442 2115 446
rect 2127 442 2131 446
rect 2271 442 2275 446
rect 2295 442 2299 446
rect 2455 442 2459 446
rect 2479 442 2483 446
rect 2655 442 2659 446
rect 2679 442 2683 446
rect 2871 442 2875 446
rect 2887 442 2891 446
rect 3103 442 3107 446
rect 3111 442 3115 446
rect 3335 442 3339 446
rect 3463 442 3467 446
rect 111 374 115 378
rect 135 374 139 378
rect 223 374 227 378
rect 255 374 259 378
rect 343 374 347 378
rect 415 374 419 378
rect 471 374 475 378
rect 583 374 587 378
rect 599 374 603 378
rect 719 374 723 378
rect 743 374 747 378
rect 839 374 843 378
rect 903 374 907 378
rect 959 374 963 378
rect 1047 374 1051 378
rect 1079 374 1083 378
rect 1183 374 1187 378
rect 1207 374 1211 378
rect 1311 374 1315 378
rect 1439 374 1443 378
rect 1567 374 1571 378
rect 1671 374 1675 378
rect 1767 374 1771 378
rect 1807 374 1811 378
rect 1831 374 1835 378
rect 1927 374 1931 378
rect 1959 374 1963 378
rect 2039 374 2043 378
rect 2111 374 2115 378
rect 2159 374 2163 378
rect 2271 374 2275 378
rect 2287 374 2291 378
rect 2423 374 2427 378
rect 2455 374 2459 378
rect 2583 374 2587 378
rect 2655 374 2659 378
rect 2759 374 2763 378
rect 2871 374 2875 378
rect 2951 374 2955 378
rect 3103 374 3107 378
rect 3151 374 3155 378
rect 3335 374 3339 378
rect 3359 374 3363 378
rect 3463 374 3467 378
rect 111 306 115 310
rect 135 306 139 310
rect 223 306 227 310
rect 263 306 267 310
rect 343 306 347 310
rect 375 306 379 310
rect 471 306 475 310
rect 487 306 491 310
rect 599 306 603 310
rect 711 306 715 310
rect 719 306 723 310
rect 815 306 819 310
rect 839 306 843 310
rect 919 306 923 310
rect 959 306 963 310
rect 1023 306 1027 310
rect 1079 306 1083 310
rect 1127 306 1131 310
rect 1207 306 1211 310
rect 1239 306 1243 310
rect 1767 306 1771 310
rect 1807 310 1811 314
rect 1927 310 1931 314
rect 2039 310 2043 314
rect 2159 310 2163 314
rect 2223 310 2227 314
rect 2287 310 2291 314
rect 2311 310 2315 314
rect 2399 310 2403 314
rect 2423 310 2427 314
rect 2487 310 2491 314
rect 2575 310 2579 314
rect 2583 310 2587 314
rect 2679 310 2683 314
rect 2759 310 2763 314
rect 2799 310 2803 314
rect 2927 310 2931 314
rect 2951 310 2955 314
rect 3071 310 3075 314
rect 3151 310 3155 314
rect 3223 310 3227 314
rect 3359 310 3363 314
rect 3367 310 3371 314
rect 3463 310 3467 314
rect 111 238 115 242
rect 263 238 267 242
rect 375 238 379 242
rect 447 238 451 242
rect 487 238 491 242
rect 535 238 539 242
rect 599 238 603 242
rect 623 238 627 242
rect 711 238 715 242
rect 807 238 811 242
rect 815 238 819 242
rect 903 238 907 242
rect 919 238 923 242
rect 999 238 1003 242
rect 1023 238 1027 242
rect 1103 238 1107 242
rect 1127 238 1131 242
rect 1207 238 1211 242
rect 1239 238 1243 242
rect 1311 238 1315 242
rect 1767 238 1771 242
rect 1807 238 1811 242
rect 2143 238 2147 242
rect 2223 238 2227 242
rect 2263 238 2267 242
rect 2311 238 2315 242
rect 2383 238 2387 242
rect 2399 238 2403 242
rect 2487 238 2491 242
rect 2511 238 2515 242
rect 2575 238 2579 242
rect 2639 238 2643 242
rect 2679 238 2683 242
rect 2767 238 2771 242
rect 2799 238 2803 242
rect 2895 238 2899 242
rect 2927 238 2931 242
rect 3015 238 3019 242
rect 3071 238 3075 242
rect 3135 238 3139 242
rect 3223 238 3227 242
rect 3263 238 3267 242
rect 3367 238 3371 242
rect 3463 238 3467 242
rect 111 146 115 150
rect 263 146 267 150
rect 351 146 355 150
rect 439 146 443 150
rect 447 146 451 150
rect 527 146 531 150
rect 535 146 539 150
rect 615 146 619 150
rect 623 146 627 150
rect 703 146 707 150
rect 711 146 715 150
rect 791 146 795 150
rect 807 146 811 150
rect 879 146 883 150
rect 903 146 907 150
rect 967 146 971 150
rect 999 146 1003 150
rect 1055 146 1059 150
rect 1103 146 1107 150
rect 1143 146 1147 150
rect 1207 146 1211 150
rect 1231 146 1235 150
rect 1311 146 1315 150
rect 1319 146 1323 150
rect 1407 146 1411 150
rect 1495 146 1499 150
rect 1583 146 1587 150
rect 1671 146 1675 150
rect 1767 146 1771 150
rect 1807 150 1811 154
rect 1831 150 1835 154
rect 1919 150 1923 154
rect 2007 150 2011 154
rect 2095 150 2099 154
rect 2143 150 2147 154
rect 2183 150 2187 154
rect 2263 150 2267 154
rect 2295 150 2299 154
rect 2383 150 2387 154
rect 2407 150 2411 154
rect 2511 150 2515 154
rect 2615 150 2619 154
rect 2639 150 2643 154
rect 2719 150 2723 154
rect 2767 150 2771 154
rect 2815 150 2819 154
rect 2895 150 2899 154
rect 2911 150 2915 154
rect 3007 150 3011 154
rect 3015 150 3019 154
rect 3103 150 3107 154
rect 3135 150 3139 154
rect 3191 150 3195 154
rect 3263 150 3267 154
rect 3279 150 3283 154
rect 3367 150 3371 154
rect 3463 150 3467 154
rect 111 82 115 86
rect 263 82 267 86
rect 351 82 355 86
rect 439 82 443 86
rect 527 82 531 86
rect 615 82 619 86
rect 703 82 707 86
rect 791 82 795 86
rect 879 82 883 86
rect 967 82 971 86
rect 1055 82 1059 86
rect 1143 82 1147 86
rect 1231 82 1235 86
rect 1319 82 1323 86
rect 1407 82 1411 86
rect 1495 82 1499 86
rect 1583 82 1587 86
rect 1671 82 1675 86
rect 1767 82 1771 86
rect 1807 86 1811 90
rect 1831 86 1835 90
rect 1919 86 1923 90
rect 2007 86 2011 90
rect 2095 86 2099 90
rect 2183 86 2187 90
rect 2295 86 2299 90
rect 2407 86 2411 90
rect 2511 86 2515 90
rect 2615 86 2619 90
rect 2719 86 2723 90
rect 2815 86 2819 90
rect 2911 86 2915 90
rect 3007 86 3011 90
rect 3103 86 3107 90
rect 3191 86 3195 90
rect 3279 86 3283 90
rect 3367 86 3371 90
rect 3463 86 3467 90
<< m4 >>
rect 96 3501 97 3507
rect 103 3506 1791 3507
rect 103 3502 111 3506
rect 115 3502 135 3506
rect 139 3502 271 3506
rect 275 3502 439 3506
rect 443 3502 615 3506
rect 619 3502 791 3506
rect 795 3502 959 3506
rect 963 3502 1119 3506
rect 1123 3502 1263 3506
rect 1267 3502 1407 3506
rect 1411 3502 1551 3506
rect 1555 3502 1671 3506
rect 1675 3502 1767 3506
rect 1771 3502 1791 3506
rect 103 3501 1791 3502
rect 1797 3501 1798 3507
rect 1790 3489 1791 3495
rect 1797 3494 3499 3495
rect 1797 3490 1807 3494
rect 1811 3490 1831 3494
rect 1835 3490 1975 3494
rect 1979 3490 2143 3494
rect 2147 3490 2311 3494
rect 2315 3490 2479 3494
rect 2483 3490 2639 3494
rect 2643 3490 2799 3494
rect 2803 3490 2967 3494
rect 2971 3490 3463 3494
rect 3467 3490 3499 3494
rect 1797 3489 3499 3490
rect 3505 3489 3506 3495
rect 84 3433 85 3439
rect 91 3438 1779 3439
rect 91 3434 111 3438
rect 115 3434 135 3438
rect 139 3434 255 3438
rect 259 3434 271 3438
rect 275 3434 415 3438
rect 419 3434 439 3438
rect 443 3434 575 3438
rect 579 3434 615 3438
rect 619 3434 735 3438
rect 739 3434 791 3438
rect 795 3434 895 3438
rect 899 3434 959 3438
rect 963 3434 1063 3438
rect 1067 3434 1119 3438
rect 1123 3434 1231 3438
rect 1235 3434 1263 3438
rect 1267 3434 1399 3438
rect 1403 3434 1407 3438
rect 1411 3434 1551 3438
rect 1555 3434 1671 3438
rect 1675 3434 1767 3438
rect 1771 3434 1779 3438
rect 91 3433 1779 3434
rect 1785 3433 1786 3439
rect 1778 3431 1786 3433
rect 1778 3425 1779 3431
rect 1785 3430 3487 3431
rect 1785 3426 1807 3430
rect 1811 3426 1831 3430
rect 1835 3426 1975 3430
rect 1979 3426 2031 3430
rect 2035 3426 2143 3430
rect 2147 3426 2151 3430
rect 2155 3426 2271 3430
rect 2275 3426 2311 3430
rect 2315 3426 2391 3430
rect 2395 3426 2479 3430
rect 2483 3426 2511 3430
rect 2515 3426 2623 3430
rect 2627 3426 2639 3430
rect 2643 3426 2727 3430
rect 2731 3426 2799 3430
rect 2803 3426 2831 3430
rect 2835 3426 2935 3430
rect 2939 3426 2967 3430
rect 2971 3426 3039 3430
rect 3043 3426 3151 3430
rect 3155 3426 3463 3430
rect 3467 3426 3487 3430
rect 1785 3425 3487 3426
rect 3493 3425 3494 3431
rect 96 3361 97 3367
rect 103 3366 1791 3367
rect 103 3362 111 3366
rect 115 3362 135 3366
rect 139 3362 255 3366
rect 259 3362 327 3366
rect 331 3362 415 3366
rect 419 3362 535 3366
rect 539 3362 575 3366
rect 579 3362 735 3366
rect 739 3362 743 3366
rect 747 3362 895 3366
rect 899 3362 935 3366
rect 939 3362 1063 3366
rect 1067 3362 1119 3366
rect 1123 3362 1231 3366
rect 1235 3362 1295 3366
rect 1299 3362 1399 3366
rect 1403 3362 1463 3366
rect 1467 3362 1639 3366
rect 1643 3362 1767 3366
rect 1771 3362 1791 3366
rect 103 3361 1791 3362
rect 1797 3363 1798 3367
rect 1797 3362 3506 3363
rect 1797 3361 1807 3362
rect 1790 3358 1807 3361
rect 1811 3358 2031 3362
rect 2035 3358 2151 3362
rect 2155 3358 2159 3362
rect 2163 3358 2271 3362
rect 2275 3358 2295 3362
rect 2299 3358 2391 3362
rect 2395 3358 2431 3362
rect 2435 3358 2511 3362
rect 2515 3358 2567 3362
rect 2571 3358 2623 3362
rect 2627 3358 2703 3362
rect 2707 3358 2727 3362
rect 2731 3358 2831 3362
rect 2835 3358 2839 3362
rect 2843 3358 2935 3362
rect 2939 3358 2975 3362
rect 2979 3358 3039 3362
rect 3043 3358 3119 3362
rect 3123 3358 3151 3362
rect 3155 3358 3463 3362
rect 3467 3358 3506 3362
rect 1790 3357 3506 3358
rect 1778 3298 3494 3299
rect 1778 3295 1807 3298
rect 84 3289 85 3295
rect 91 3294 1779 3295
rect 91 3290 111 3294
rect 115 3290 135 3294
rect 139 3290 279 3294
rect 283 3290 327 3294
rect 331 3290 463 3294
rect 467 3290 535 3294
rect 539 3290 647 3294
rect 651 3290 743 3294
rect 747 3290 831 3294
rect 835 3290 935 3294
rect 939 3290 1007 3294
rect 1011 3290 1119 3294
rect 1123 3290 1175 3294
rect 1179 3290 1295 3294
rect 1299 3290 1343 3294
rect 1347 3290 1463 3294
rect 1467 3290 1503 3294
rect 1507 3290 1639 3294
rect 1643 3290 1671 3294
rect 1675 3290 1767 3294
rect 1771 3290 1779 3294
rect 91 3289 1779 3290
rect 1785 3294 1807 3295
rect 1811 3294 2087 3298
rect 2091 3294 2159 3298
rect 2163 3294 2239 3298
rect 2243 3294 2295 3298
rect 2299 3294 2399 3298
rect 2403 3294 2431 3298
rect 2435 3294 2559 3298
rect 2563 3294 2567 3298
rect 2571 3294 2703 3298
rect 2707 3294 2719 3298
rect 2723 3294 2839 3298
rect 2843 3294 2879 3298
rect 2883 3294 2975 3298
rect 2979 3294 3039 3298
rect 3043 3294 3119 3298
rect 3123 3294 3199 3298
rect 3203 3294 3463 3298
rect 3467 3294 3494 3298
rect 1785 3293 3494 3294
rect 1785 3289 1786 3293
rect 1790 3225 1791 3231
rect 1797 3230 3499 3231
rect 1797 3226 1807 3230
rect 1811 3226 1911 3230
rect 1915 3226 2047 3230
rect 2051 3226 2087 3230
rect 2091 3226 2199 3230
rect 2203 3226 2239 3230
rect 2243 3226 2359 3230
rect 2363 3226 2399 3230
rect 2403 3226 2527 3230
rect 2531 3226 2559 3230
rect 2563 3226 2687 3230
rect 2691 3226 2719 3230
rect 2723 3226 2847 3230
rect 2851 3226 2879 3230
rect 2883 3226 3007 3230
rect 3011 3226 3039 3230
rect 3043 3226 3167 3230
rect 3171 3226 3199 3230
rect 3203 3226 3335 3230
rect 3339 3226 3463 3230
rect 3467 3226 3499 3230
rect 1797 3225 3499 3226
rect 3505 3225 3506 3231
rect 1790 3223 1798 3225
rect 96 3217 97 3223
rect 103 3222 1791 3223
rect 103 3218 111 3222
rect 115 3218 135 3222
rect 139 3218 183 3222
rect 187 3218 279 3222
rect 283 3218 327 3222
rect 331 3218 463 3222
rect 467 3218 487 3222
rect 491 3218 647 3222
rect 651 3218 807 3222
rect 811 3218 831 3222
rect 835 3218 967 3222
rect 971 3218 1007 3222
rect 1011 3218 1135 3222
rect 1139 3218 1175 3222
rect 1179 3218 1303 3222
rect 1307 3218 1343 3222
rect 1347 3218 1471 3222
rect 1475 3218 1503 3222
rect 1507 3218 1671 3222
rect 1675 3218 1767 3222
rect 1771 3218 1791 3222
rect 103 3217 1791 3218
rect 1797 3217 1798 3223
rect 1778 3161 1779 3167
rect 1785 3166 3487 3167
rect 1785 3162 1807 3166
rect 1811 3162 1831 3166
rect 1835 3162 1911 3166
rect 1915 3162 2007 3166
rect 2011 3162 2047 3166
rect 2051 3162 2199 3166
rect 2203 3162 2207 3166
rect 2211 3162 2359 3166
rect 2363 3162 2399 3166
rect 2403 3162 2527 3166
rect 2531 3162 2583 3166
rect 2587 3162 2687 3166
rect 2691 3162 2759 3166
rect 2763 3162 2847 3166
rect 2851 3162 2919 3166
rect 2923 3162 3007 3166
rect 3011 3162 3079 3166
rect 3083 3162 3167 3166
rect 3171 3162 3231 3166
rect 3235 3162 3335 3166
rect 3339 3162 3367 3166
rect 3371 3162 3463 3166
rect 3467 3162 3487 3166
rect 1785 3161 3487 3162
rect 3493 3161 3494 3167
rect 1778 3159 1786 3161
rect 84 3153 85 3159
rect 91 3158 1779 3159
rect 91 3154 111 3158
rect 115 3154 183 3158
rect 187 3154 327 3158
rect 331 3154 367 3158
rect 371 3154 487 3158
rect 491 3154 607 3158
rect 611 3154 647 3158
rect 651 3154 727 3158
rect 731 3154 807 3158
rect 811 3154 847 3158
rect 851 3154 967 3158
rect 971 3154 1079 3158
rect 1083 3154 1135 3158
rect 1139 3154 1199 3158
rect 1203 3154 1303 3158
rect 1307 3154 1319 3158
rect 1323 3154 1471 3158
rect 1475 3154 1767 3158
rect 1771 3154 1779 3158
rect 91 3153 1779 3154
rect 1785 3153 1786 3159
rect 1790 3094 3506 3095
rect 1790 3091 1807 3094
rect 96 3085 97 3091
rect 103 3090 1791 3091
rect 103 3086 111 3090
rect 115 3086 367 3090
rect 371 3086 439 3090
rect 443 3086 487 3090
rect 491 3086 527 3090
rect 531 3086 607 3090
rect 611 3086 615 3090
rect 619 3086 703 3090
rect 707 3086 727 3090
rect 731 3086 791 3090
rect 795 3086 847 3090
rect 851 3086 879 3090
rect 883 3086 967 3090
rect 971 3086 1055 3090
rect 1059 3086 1079 3090
rect 1083 3086 1143 3090
rect 1147 3086 1199 3090
rect 1203 3086 1319 3090
rect 1323 3086 1767 3090
rect 1771 3086 1791 3090
rect 103 3085 1791 3086
rect 1797 3090 1807 3091
rect 1811 3090 1831 3094
rect 1835 3090 1959 3094
rect 1963 3090 2007 3094
rect 2011 3090 2119 3094
rect 2123 3090 2207 3094
rect 2211 3090 2295 3094
rect 2299 3090 2399 3094
rect 2403 3090 2487 3094
rect 2491 3090 2583 3094
rect 2587 3090 2695 3094
rect 2699 3090 2759 3094
rect 2763 3090 2919 3094
rect 2923 3090 3079 3094
rect 3083 3090 3151 3094
rect 3155 3090 3231 3094
rect 3235 3090 3367 3094
rect 3371 3090 3463 3094
rect 3467 3090 3506 3094
rect 1797 3089 3506 3090
rect 1797 3085 1798 3089
rect 84 3013 85 3019
rect 91 3018 1779 3019
rect 91 3014 111 3018
rect 115 3014 439 3018
rect 443 3014 503 3018
rect 507 3014 527 3018
rect 531 3014 591 3018
rect 595 3014 615 3018
rect 619 3014 679 3018
rect 683 3014 703 3018
rect 707 3014 767 3018
rect 771 3014 791 3018
rect 795 3014 855 3018
rect 859 3014 879 3018
rect 883 3014 943 3018
rect 947 3014 967 3018
rect 971 3014 1031 3018
rect 1035 3014 1055 3018
rect 1059 3014 1119 3018
rect 1123 3014 1143 3018
rect 1147 3014 1207 3018
rect 1211 3014 1295 3018
rect 1299 3014 1767 3018
rect 1771 3014 1779 3018
rect 91 3013 1779 3014
rect 1785 3015 1786 3019
rect 1785 3014 3494 3015
rect 1785 3013 1807 3014
rect 1778 3010 1807 3013
rect 1811 3010 1831 3014
rect 1835 3010 1919 3014
rect 1923 3010 1959 3014
rect 1963 3010 2031 3014
rect 2035 3010 2119 3014
rect 2123 3010 2143 3014
rect 2147 3010 2247 3014
rect 2251 3010 2295 3014
rect 2299 3010 2359 3014
rect 2363 3010 2479 3014
rect 2483 3010 2487 3014
rect 2491 3010 2623 3014
rect 2627 3010 2695 3014
rect 2699 3010 2791 3014
rect 2795 3010 2919 3014
rect 2923 3010 2983 3014
rect 2987 3010 3151 3014
rect 3155 3010 3183 3014
rect 3187 3010 3367 3014
rect 3371 3010 3463 3014
rect 3467 3010 3494 3014
rect 1778 3009 3494 3010
rect 96 2937 97 2943
rect 103 2942 1791 2943
rect 103 2938 111 2942
rect 115 2938 327 2942
rect 331 2938 447 2942
rect 451 2938 503 2942
rect 507 2938 575 2942
rect 579 2938 591 2942
rect 595 2938 679 2942
rect 683 2938 711 2942
rect 715 2938 767 2942
rect 771 2938 847 2942
rect 851 2938 855 2942
rect 859 2938 943 2942
rect 947 2938 975 2942
rect 979 2938 1031 2942
rect 1035 2938 1103 2942
rect 1107 2938 1119 2942
rect 1123 2938 1207 2942
rect 1211 2938 1231 2942
rect 1235 2938 1295 2942
rect 1299 2938 1359 2942
rect 1363 2938 1495 2942
rect 1499 2938 1767 2942
rect 1771 2938 1791 2942
rect 103 2937 1791 2938
rect 1797 2939 1798 2943
rect 1797 2938 3506 2939
rect 1797 2937 1807 2938
rect 1790 2934 1807 2937
rect 1811 2934 1831 2938
rect 1835 2934 1919 2938
rect 1923 2934 2015 2938
rect 2019 2934 2031 2938
rect 2035 2934 2143 2938
rect 2147 2934 2215 2938
rect 2219 2934 2247 2938
rect 2251 2934 2359 2938
rect 2363 2934 2407 2938
rect 2411 2934 2479 2938
rect 2483 2934 2591 2938
rect 2595 2934 2623 2938
rect 2627 2934 2759 2938
rect 2763 2934 2791 2938
rect 2795 2934 2911 2938
rect 2915 2934 2983 2938
rect 2987 2934 3063 2938
rect 3067 2934 3183 2938
rect 3187 2934 3207 2938
rect 3211 2934 3359 2938
rect 3363 2934 3367 2938
rect 3371 2934 3463 2938
rect 3467 2934 3506 2938
rect 1790 2933 3506 2934
rect 1778 2874 3494 2875
rect 1778 2871 1807 2874
rect 84 2865 85 2871
rect 91 2870 1779 2871
rect 91 2866 111 2870
rect 115 2866 135 2870
rect 139 2866 255 2870
rect 259 2866 327 2870
rect 331 2866 415 2870
rect 419 2866 447 2870
rect 451 2866 575 2870
rect 579 2866 711 2870
rect 715 2866 735 2870
rect 739 2866 847 2870
rect 851 2866 895 2870
rect 899 2866 975 2870
rect 979 2866 1047 2870
rect 1051 2866 1103 2870
rect 1107 2866 1191 2870
rect 1195 2866 1231 2870
rect 1235 2866 1343 2870
rect 1347 2866 1359 2870
rect 1363 2866 1495 2870
rect 1499 2866 1767 2870
rect 1771 2866 1779 2870
rect 91 2865 1779 2866
rect 1785 2870 1807 2871
rect 1811 2870 1831 2874
rect 1835 2870 1999 2874
rect 2003 2870 2015 2874
rect 2019 2870 2191 2874
rect 2195 2870 2215 2874
rect 2219 2870 2383 2874
rect 2387 2870 2407 2874
rect 2411 2870 2567 2874
rect 2571 2870 2591 2874
rect 2595 2870 2735 2874
rect 2739 2870 2759 2874
rect 2763 2870 2903 2874
rect 2907 2870 2911 2874
rect 2915 2870 3063 2874
rect 3067 2870 3207 2874
rect 3211 2870 3223 2874
rect 3227 2870 3359 2874
rect 3363 2870 3367 2874
rect 3371 2870 3463 2874
rect 3467 2870 3494 2874
rect 1785 2869 3494 2870
rect 1785 2865 1786 2869
rect 1790 2801 1791 2807
rect 1797 2806 3499 2807
rect 1797 2802 1807 2806
rect 1811 2802 1831 2806
rect 1835 2802 1999 2806
rect 2003 2802 2015 2806
rect 2019 2802 2191 2806
rect 2195 2802 2215 2806
rect 2219 2802 2383 2806
rect 2387 2802 2407 2806
rect 2411 2802 2567 2806
rect 2571 2802 2583 2806
rect 2587 2802 2735 2806
rect 2739 2802 2751 2806
rect 2755 2802 2903 2806
rect 2907 2802 2911 2806
rect 2915 2802 3063 2806
rect 3067 2802 3071 2806
rect 3075 2802 3223 2806
rect 3227 2802 3231 2806
rect 3235 2802 3367 2806
rect 3371 2802 3463 2806
rect 3467 2802 3499 2806
rect 1797 2801 3499 2802
rect 3505 2801 3506 2807
rect 96 2789 97 2795
rect 103 2794 1791 2795
rect 103 2790 111 2794
rect 115 2790 135 2794
rect 139 2790 247 2794
rect 251 2790 255 2794
rect 259 2790 391 2794
rect 395 2790 415 2794
rect 419 2790 543 2794
rect 547 2790 575 2794
rect 579 2790 695 2794
rect 699 2790 735 2794
rect 739 2790 855 2794
rect 859 2790 895 2794
rect 899 2790 1023 2794
rect 1027 2790 1047 2794
rect 1051 2790 1191 2794
rect 1195 2790 1343 2794
rect 1347 2790 1359 2794
rect 1363 2790 1495 2794
rect 1499 2790 1527 2794
rect 1531 2790 1671 2794
rect 1675 2790 1767 2794
rect 1771 2790 1791 2794
rect 103 2789 1791 2790
rect 1797 2789 1798 2795
rect 1778 2726 3494 2727
rect 1778 2723 1807 2726
rect 84 2717 85 2723
rect 91 2722 1779 2723
rect 91 2718 111 2722
rect 115 2718 135 2722
rect 139 2718 247 2722
rect 251 2718 359 2722
rect 363 2718 391 2722
rect 395 2718 479 2722
rect 483 2718 543 2722
rect 547 2718 615 2722
rect 619 2718 695 2722
rect 699 2718 759 2722
rect 763 2718 855 2722
rect 859 2718 911 2722
rect 915 2718 1023 2722
rect 1027 2718 1063 2722
rect 1067 2718 1191 2722
rect 1195 2718 1215 2722
rect 1219 2718 1359 2722
rect 1363 2718 1375 2722
rect 1379 2718 1527 2722
rect 1531 2718 1535 2722
rect 1539 2718 1671 2722
rect 1675 2718 1767 2722
rect 1771 2718 1779 2722
rect 91 2717 1779 2718
rect 1785 2722 1807 2723
rect 1811 2722 1831 2726
rect 1835 2722 2015 2726
rect 2019 2722 2039 2726
rect 2043 2722 2159 2726
rect 2163 2722 2215 2726
rect 2219 2722 2279 2726
rect 2283 2722 2407 2726
rect 2411 2722 2543 2726
rect 2547 2722 2583 2726
rect 2587 2722 2687 2726
rect 2691 2722 2751 2726
rect 2755 2722 2847 2726
rect 2851 2722 2911 2726
rect 2915 2722 3023 2726
rect 3027 2722 3071 2726
rect 3075 2722 3207 2726
rect 3211 2722 3231 2726
rect 3235 2722 3367 2726
rect 3371 2722 3463 2726
rect 3467 2722 3494 2726
rect 1785 2721 3494 2722
rect 1785 2717 1786 2721
rect 96 2645 97 2651
rect 103 2650 1791 2651
rect 103 2646 111 2650
rect 115 2646 247 2650
rect 251 2646 359 2650
rect 363 2646 463 2650
rect 467 2646 479 2650
rect 483 2646 551 2650
rect 555 2646 615 2650
rect 619 2646 639 2650
rect 643 2646 743 2650
rect 747 2646 759 2650
rect 763 2646 855 2650
rect 859 2646 911 2650
rect 915 2646 983 2650
rect 987 2646 1063 2650
rect 1067 2646 1127 2650
rect 1131 2646 1215 2650
rect 1219 2646 1279 2650
rect 1283 2646 1375 2650
rect 1379 2646 1439 2650
rect 1443 2646 1535 2650
rect 1539 2646 1607 2650
rect 1611 2646 1671 2650
rect 1675 2646 1767 2650
rect 1771 2646 1791 2650
rect 103 2645 1791 2646
rect 1797 2650 3506 2651
rect 1797 2646 1807 2650
rect 1811 2646 1871 2650
rect 1875 2646 1967 2650
rect 1971 2646 2039 2650
rect 2043 2646 2071 2650
rect 2075 2646 2159 2650
rect 2163 2646 2183 2650
rect 2187 2646 2279 2650
rect 2283 2646 2295 2650
rect 2299 2646 2407 2650
rect 2411 2646 2431 2650
rect 2435 2646 2543 2650
rect 2547 2646 2583 2650
rect 2587 2646 2687 2650
rect 2691 2646 2759 2650
rect 2763 2646 2847 2650
rect 2851 2646 2959 2650
rect 2963 2646 3023 2650
rect 3027 2646 3167 2650
rect 3171 2646 3207 2650
rect 3211 2646 3367 2650
rect 3371 2646 3463 2650
rect 3467 2646 3506 2650
rect 1797 2645 3506 2646
rect 84 2573 85 2579
rect 91 2578 1779 2579
rect 91 2574 111 2578
rect 115 2574 463 2578
rect 467 2574 503 2578
rect 507 2574 551 2578
rect 555 2574 591 2578
rect 595 2574 639 2578
rect 643 2574 679 2578
rect 683 2574 743 2578
rect 747 2574 775 2578
rect 779 2574 855 2578
rect 859 2574 879 2578
rect 883 2574 983 2578
rect 987 2574 991 2578
rect 995 2574 1103 2578
rect 1107 2574 1127 2578
rect 1131 2574 1223 2578
rect 1227 2574 1279 2578
rect 1283 2574 1351 2578
rect 1355 2574 1439 2578
rect 1443 2574 1479 2578
rect 1483 2574 1607 2578
rect 1611 2574 1767 2578
rect 1771 2574 1779 2578
rect 91 2573 1779 2574
rect 1785 2575 1786 2579
rect 1785 2574 3494 2575
rect 1785 2573 1807 2574
rect 1778 2570 1807 2573
rect 1811 2570 1831 2574
rect 1835 2570 1871 2574
rect 1875 2570 1919 2574
rect 1923 2570 1967 2574
rect 1971 2570 2007 2574
rect 2011 2570 2071 2574
rect 2075 2570 2111 2574
rect 2115 2570 2183 2574
rect 2187 2570 2223 2574
rect 2227 2570 2295 2574
rect 2299 2570 2343 2574
rect 2347 2570 2431 2574
rect 2435 2570 2487 2574
rect 2491 2570 2583 2574
rect 2587 2570 2647 2574
rect 2651 2570 2759 2574
rect 2763 2570 2815 2574
rect 2819 2570 2959 2574
rect 2963 2570 2999 2574
rect 3003 2570 3167 2574
rect 3171 2570 3191 2574
rect 3195 2570 3367 2574
rect 3371 2570 3463 2574
rect 3467 2570 3494 2574
rect 1778 2569 3494 2570
rect 1790 2510 3506 2511
rect 1790 2507 1807 2510
rect 96 2501 97 2507
rect 103 2506 1791 2507
rect 103 2502 111 2506
rect 115 2502 503 2506
rect 507 2502 551 2506
rect 555 2502 591 2506
rect 595 2502 679 2506
rect 683 2502 735 2506
rect 739 2502 775 2506
rect 779 2502 879 2506
rect 883 2502 911 2506
rect 915 2502 991 2506
rect 995 2502 1079 2506
rect 1083 2502 1103 2506
rect 1107 2502 1223 2506
rect 1227 2502 1239 2506
rect 1243 2502 1351 2506
rect 1355 2502 1399 2506
rect 1403 2502 1479 2506
rect 1483 2502 1567 2506
rect 1571 2502 1607 2506
rect 1611 2502 1767 2506
rect 1771 2502 1791 2506
rect 103 2501 1791 2502
rect 1797 2506 1807 2507
rect 1811 2506 1831 2510
rect 1835 2506 1919 2510
rect 1923 2506 1951 2510
rect 1955 2506 2007 2510
rect 2011 2506 2039 2510
rect 2043 2506 2111 2510
rect 2115 2506 2135 2510
rect 2139 2506 2223 2510
rect 2227 2506 2239 2510
rect 2243 2506 2343 2510
rect 2347 2506 2367 2510
rect 2371 2506 2487 2510
rect 2491 2506 2527 2510
rect 2531 2506 2647 2510
rect 2651 2506 2711 2510
rect 2715 2506 2815 2510
rect 2819 2506 2919 2510
rect 2923 2506 2999 2510
rect 3003 2506 3143 2510
rect 3147 2506 3191 2510
rect 3195 2506 3367 2510
rect 3371 2506 3463 2510
rect 3467 2506 3506 2510
rect 1797 2505 3506 2506
rect 1797 2501 1798 2505
rect 84 2437 85 2443
rect 91 2442 1779 2443
rect 91 2438 111 2442
rect 115 2438 415 2442
rect 419 2438 503 2442
rect 507 2438 551 2442
rect 555 2438 599 2442
rect 603 2438 703 2442
rect 707 2438 735 2442
rect 739 2438 807 2442
rect 811 2438 911 2442
rect 915 2438 919 2442
rect 923 2438 1039 2442
rect 1043 2438 1079 2442
rect 1083 2438 1167 2442
rect 1171 2438 1239 2442
rect 1243 2438 1295 2442
rect 1299 2438 1399 2442
rect 1403 2438 1423 2442
rect 1427 2438 1567 2442
rect 1571 2438 1767 2442
rect 1771 2438 1779 2442
rect 91 2437 1779 2438
rect 1785 2439 1786 2443
rect 1785 2438 3494 2439
rect 1785 2437 1807 2438
rect 1778 2434 1807 2437
rect 1811 2434 1951 2438
rect 1955 2434 2039 2438
rect 2043 2434 2135 2438
rect 2139 2434 2215 2438
rect 2219 2434 2239 2438
rect 2243 2434 2303 2438
rect 2307 2434 2367 2438
rect 2371 2434 2391 2438
rect 2395 2434 2479 2438
rect 2483 2434 2527 2438
rect 2531 2434 2567 2438
rect 2571 2434 2655 2438
rect 2659 2434 2711 2438
rect 2715 2434 2743 2438
rect 2747 2434 2839 2438
rect 2843 2434 2919 2438
rect 2923 2434 2935 2438
rect 2939 2434 3143 2438
rect 3147 2434 3367 2438
rect 3371 2434 3463 2438
rect 3467 2434 3494 2438
rect 1778 2433 3494 2434
rect 96 2369 97 2375
rect 103 2374 1791 2375
rect 103 2370 111 2374
rect 115 2370 319 2374
rect 323 2370 415 2374
rect 419 2370 431 2374
rect 435 2370 503 2374
rect 507 2370 543 2374
rect 547 2370 599 2374
rect 603 2370 655 2374
rect 659 2370 703 2374
rect 707 2370 767 2374
rect 771 2370 807 2374
rect 811 2370 879 2374
rect 883 2370 919 2374
rect 923 2370 991 2374
rect 995 2370 1039 2374
rect 1043 2370 1103 2374
rect 1107 2370 1167 2374
rect 1171 2370 1215 2374
rect 1219 2370 1295 2374
rect 1299 2370 1335 2374
rect 1339 2370 1423 2374
rect 1427 2370 1767 2374
rect 1771 2370 1791 2374
rect 103 2369 1791 2370
rect 1797 2374 3506 2375
rect 1797 2370 1807 2374
rect 1811 2370 2167 2374
rect 2171 2370 2215 2374
rect 2219 2370 2263 2374
rect 2267 2370 2303 2374
rect 2307 2370 2367 2374
rect 2371 2370 2391 2374
rect 2395 2370 2471 2374
rect 2475 2370 2479 2374
rect 2483 2370 2567 2374
rect 2571 2370 2575 2374
rect 2579 2370 2655 2374
rect 2659 2370 2687 2374
rect 2691 2370 2743 2374
rect 2747 2370 2799 2374
rect 2803 2370 2839 2374
rect 2843 2370 2911 2374
rect 2915 2370 2935 2374
rect 2939 2370 3023 2374
rect 3027 2370 3463 2374
rect 3467 2370 3506 2374
rect 1797 2369 3506 2370
rect 84 2297 85 2303
rect 91 2302 1779 2303
rect 91 2298 111 2302
rect 115 2298 151 2302
rect 155 2298 271 2302
rect 275 2298 319 2302
rect 323 2298 391 2302
rect 395 2298 431 2302
rect 435 2298 519 2302
rect 523 2298 543 2302
rect 547 2298 647 2302
rect 651 2298 655 2302
rect 659 2298 767 2302
rect 771 2298 775 2302
rect 779 2298 879 2302
rect 883 2298 895 2302
rect 899 2298 991 2302
rect 995 2298 1015 2302
rect 1019 2298 1103 2302
rect 1107 2298 1143 2302
rect 1147 2298 1215 2302
rect 1219 2298 1271 2302
rect 1275 2298 1335 2302
rect 1339 2298 1767 2302
rect 1771 2298 1779 2302
rect 91 2297 1779 2298
rect 1785 2302 3494 2303
rect 1785 2298 1807 2302
rect 1811 2298 1887 2302
rect 1891 2298 2039 2302
rect 2043 2298 2167 2302
rect 2171 2298 2199 2302
rect 2203 2298 2263 2302
rect 2267 2298 2367 2302
rect 2371 2298 2375 2302
rect 2379 2298 2471 2302
rect 2475 2298 2551 2302
rect 2555 2298 2575 2302
rect 2579 2298 2687 2302
rect 2691 2298 2719 2302
rect 2723 2298 2799 2302
rect 2803 2298 2887 2302
rect 2891 2298 2911 2302
rect 2915 2298 3023 2302
rect 3027 2298 3055 2302
rect 3059 2298 3223 2302
rect 3227 2298 3367 2302
rect 3371 2298 3463 2302
rect 3467 2298 3494 2302
rect 1785 2297 3494 2298
rect 1790 2238 3506 2239
rect 1790 2235 1807 2238
rect 96 2229 97 2235
rect 103 2234 1791 2235
rect 103 2230 111 2234
rect 115 2230 135 2234
rect 139 2230 151 2234
rect 155 2230 247 2234
rect 251 2230 271 2234
rect 275 2230 391 2234
rect 395 2230 407 2234
rect 411 2230 519 2234
rect 523 2230 583 2234
rect 587 2230 647 2234
rect 651 2230 767 2234
rect 771 2230 775 2234
rect 779 2230 895 2234
rect 899 2230 951 2234
rect 955 2230 1015 2234
rect 1019 2230 1135 2234
rect 1139 2230 1143 2234
rect 1147 2230 1271 2234
rect 1275 2230 1319 2234
rect 1323 2230 1503 2234
rect 1507 2230 1671 2234
rect 1675 2230 1767 2234
rect 1771 2230 1791 2234
rect 103 2229 1791 2230
rect 1797 2234 1807 2235
rect 1811 2234 1831 2238
rect 1835 2234 1887 2238
rect 1891 2234 1967 2238
rect 1971 2234 2039 2238
rect 2043 2234 2135 2238
rect 2139 2234 2199 2238
rect 2203 2234 2311 2238
rect 2315 2234 2375 2238
rect 2379 2234 2487 2238
rect 2491 2234 2551 2238
rect 2555 2234 2655 2238
rect 2659 2234 2719 2238
rect 2723 2234 2815 2238
rect 2819 2234 2887 2238
rect 2891 2234 2959 2238
rect 2963 2234 3055 2238
rect 3059 2234 3103 2238
rect 3107 2234 3223 2238
rect 3227 2234 3247 2238
rect 3251 2234 3367 2238
rect 3371 2234 3463 2238
rect 3467 2234 3506 2238
rect 1797 2233 3506 2234
rect 1797 2229 1798 2233
rect 1778 2169 1779 2175
rect 1785 2174 3487 2175
rect 1785 2170 1807 2174
rect 1811 2170 1831 2174
rect 1835 2170 1967 2174
rect 1971 2170 2135 2174
rect 2139 2170 2311 2174
rect 2315 2170 2487 2174
rect 2491 2170 2655 2174
rect 2659 2170 2815 2174
rect 2819 2170 2927 2174
rect 2931 2170 2959 2174
rect 2963 2170 3015 2174
rect 3019 2170 3103 2174
rect 3107 2170 3191 2174
rect 3195 2170 3247 2174
rect 3251 2170 3279 2174
rect 3283 2170 3367 2174
rect 3371 2170 3463 2174
rect 3467 2170 3487 2174
rect 1785 2169 3487 2170
rect 3493 2169 3494 2175
rect 84 2157 85 2163
rect 91 2162 1779 2163
rect 91 2158 111 2162
rect 115 2158 135 2162
rect 139 2158 247 2162
rect 251 2158 391 2162
rect 395 2158 407 2162
rect 411 2158 543 2162
rect 547 2158 583 2162
rect 587 2158 695 2162
rect 699 2158 767 2162
rect 771 2158 839 2162
rect 843 2158 951 2162
rect 955 2158 975 2162
rect 979 2158 1103 2162
rect 1107 2158 1135 2162
rect 1139 2158 1231 2162
rect 1235 2158 1319 2162
rect 1323 2158 1351 2162
rect 1355 2158 1463 2162
rect 1467 2158 1503 2162
rect 1507 2158 1575 2162
rect 1579 2158 1671 2162
rect 1675 2158 1767 2162
rect 1771 2158 1779 2162
rect 91 2157 1779 2158
rect 1785 2157 1786 2163
rect 1790 2097 1791 2103
rect 1797 2102 3499 2103
rect 1797 2098 1807 2102
rect 1811 2098 1831 2102
rect 1835 2098 1991 2102
rect 1995 2098 2167 2102
rect 2171 2098 2343 2102
rect 2347 2098 2503 2102
rect 2507 2098 2655 2102
rect 2659 2098 2791 2102
rect 2795 2098 2919 2102
rect 2923 2098 2927 2102
rect 2931 2098 3015 2102
rect 3019 2098 3039 2102
rect 3043 2098 3103 2102
rect 3107 2098 3159 2102
rect 3163 2098 3191 2102
rect 3195 2098 3271 2102
rect 3275 2098 3279 2102
rect 3283 2098 3367 2102
rect 3371 2098 3463 2102
rect 3467 2098 3499 2102
rect 1797 2097 3499 2098
rect 3505 2097 3506 2103
rect 1790 2095 1798 2097
rect 96 2089 97 2095
rect 103 2094 1791 2095
rect 103 2090 111 2094
rect 115 2090 135 2094
rect 139 2090 223 2094
rect 227 2090 247 2094
rect 251 2090 343 2094
rect 347 2090 391 2094
rect 395 2090 463 2094
rect 467 2090 543 2094
rect 547 2090 583 2094
rect 587 2090 695 2094
rect 699 2090 703 2094
rect 707 2090 823 2094
rect 827 2090 839 2094
rect 843 2090 935 2094
rect 939 2090 975 2094
rect 979 2090 1047 2094
rect 1051 2090 1103 2094
rect 1107 2090 1159 2094
rect 1163 2090 1231 2094
rect 1235 2090 1279 2094
rect 1283 2090 1351 2094
rect 1355 2090 1463 2094
rect 1467 2090 1575 2094
rect 1579 2090 1671 2094
rect 1675 2090 1767 2094
rect 1771 2090 1791 2094
rect 103 2089 1791 2090
rect 1797 2089 1798 2095
rect 1778 2029 1779 2035
rect 1785 2034 3487 2035
rect 1785 2030 1807 2034
rect 1811 2030 1831 2034
rect 1835 2030 1991 2034
rect 1995 2030 2015 2034
rect 2019 2030 2167 2034
rect 2171 2030 2223 2034
rect 2227 2030 2343 2034
rect 2347 2030 2431 2034
rect 2435 2030 2503 2034
rect 2507 2030 2631 2034
rect 2635 2030 2655 2034
rect 2659 2030 2791 2034
rect 2795 2030 2823 2034
rect 2827 2030 2919 2034
rect 2923 2030 3007 2034
rect 3011 2030 3039 2034
rect 3043 2030 3159 2034
rect 3163 2030 3199 2034
rect 3203 2030 3271 2034
rect 3275 2030 3367 2034
rect 3371 2030 3463 2034
rect 3467 2030 3487 2034
rect 1785 2029 3487 2030
rect 3493 2029 3494 2035
rect 84 2017 85 2023
rect 91 2022 1779 2023
rect 91 2018 111 2022
rect 115 2018 135 2022
rect 139 2018 223 2022
rect 227 2018 239 2022
rect 243 2018 343 2022
rect 347 2018 367 2022
rect 371 2018 463 2022
rect 467 2018 503 2022
rect 507 2018 583 2022
rect 587 2018 639 2022
rect 643 2018 703 2022
rect 707 2018 775 2022
rect 779 2018 823 2022
rect 827 2018 911 2022
rect 915 2018 935 2022
rect 939 2018 1047 2022
rect 1051 2018 1159 2022
rect 1163 2018 1183 2022
rect 1187 2018 1279 2022
rect 1283 2018 1327 2022
rect 1331 2018 1767 2022
rect 1771 2018 1779 2022
rect 91 2017 1779 2018
rect 1785 2017 1786 2023
rect 1790 1961 1791 1967
rect 1797 1966 3499 1967
rect 1797 1962 1807 1966
rect 1811 1962 1831 1966
rect 1835 1962 1863 1966
rect 1867 1962 1999 1966
rect 2003 1962 2015 1966
rect 2019 1962 2143 1966
rect 2147 1962 2223 1966
rect 2227 1962 2287 1966
rect 2291 1962 2431 1966
rect 2435 1962 2575 1966
rect 2579 1962 2631 1966
rect 2635 1962 2711 1966
rect 2715 1962 2823 1966
rect 2827 1962 2831 1966
rect 2835 1962 2951 1966
rect 2955 1962 3007 1966
rect 3011 1962 3063 1966
rect 3067 1962 3167 1966
rect 3171 1962 3199 1966
rect 3203 1962 3279 1966
rect 3283 1962 3367 1966
rect 3371 1962 3463 1966
rect 3467 1962 3499 1966
rect 1797 1961 3499 1962
rect 3505 1961 3506 1967
rect 96 1949 97 1955
rect 103 1954 1791 1955
rect 103 1950 111 1954
rect 115 1950 135 1954
rect 139 1950 239 1954
rect 243 1950 295 1954
rect 299 1950 367 1954
rect 371 1950 423 1954
rect 427 1950 503 1954
rect 507 1950 559 1954
rect 563 1950 639 1954
rect 643 1950 703 1954
rect 707 1950 775 1954
rect 779 1950 855 1954
rect 859 1950 911 1954
rect 915 1950 1007 1954
rect 1011 1950 1047 1954
rect 1051 1950 1159 1954
rect 1163 1950 1183 1954
rect 1187 1950 1311 1954
rect 1315 1950 1327 1954
rect 1331 1950 1471 1954
rect 1475 1950 1767 1954
rect 1771 1950 1791 1954
rect 103 1949 1791 1950
rect 1797 1949 1798 1955
rect 1778 1893 1779 1899
rect 1785 1898 3487 1899
rect 1785 1894 1807 1898
rect 1811 1894 1863 1898
rect 1867 1894 1999 1898
rect 2003 1894 2015 1898
rect 2019 1894 2111 1898
rect 2115 1894 2143 1898
rect 2147 1894 2215 1898
rect 2219 1894 2287 1898
rect 2291 1894 2327 1898
rect 2331 1894 2431 1898
rect 2435 1894 2439 1898
rect 2443 1894 2543 1898
rect 2547 1894 2575 1898
rect 2579 1894 2647 1898
rect 2651 1894 2711 1898
rect 2715 1894 2759 1898
rect 2763 1894 2831 1898
rect 2835 1894 2871 1898
rect 2875 1894 2951 1898
rect 2955 1894 2983 1898
rect 2987 1894 3063 1898
rect 3067 1894 3167 1898
rect 3171 1894 3279 1898
rect 3283 1894 3367 1898
rect 3371 1894 3463 1898
rect 3467 1894 3487 1898
rect 1785 1893 3487 1894
rect 3493 1893 3494 1899
rect 1778 1891 1786 1893
rect 84 1885 85 1891
rect 91 1890 1779 1891
rect 91 1886 111 1890
rect 115 1886 295 1890
rect 299 1886 423 1890
rect 427 1886 431 1890
rect 435 1886 559 1890
rect 563 1886 575 1890
rect 579 1886 703 1890
rect 707 1886 727 1890
rect 731 1886 855 1890
rect 859 1886 887 1890
rect 891 1886 1007 1890
rect 1011 1886 1047 1890
rect 1051 1886 1159 1890
rect 1163 1886 1199 1890
rect 1203 1886 1311 1890
rect 1315 1886 1351 1890
rect 1355 1886 1471 1890
rect 1475 1886 1511 1890
rect 1515 1886 1671 1890
rect 1675 1886 1767 1890
rect 1771 1886 1779 1890
rect 91 1885 1779 1886
rect 1785 1885 1786 1891
rect 1790 1826 3506 1827
rect 1790 1823 1807 1826
rect 96 1817 97 1823
rect 103 1822 1791 1823
rect 103 1818 111 1822
rect 115 1818 431 1822
rect 435 1818 511 1822
rect 515 1818 575 1822
rect 579 1818 631 1822
rect 635 1818 727 1822
rect 731 1818 759 1822
rect 763 1818 887 1822
rect 891 1818 1023 1822
rect 1027 1818 1047 1822
rect 1051 1818 1151 1822
rect 1155 1818 1199 1822
rect 1203 1818 1279 1822
rect 1283 1818 1351 1822
rect 1355 1818 1407 1822
rect 1411 1818 1511 1822
rect 1515 1818 1535 1822
rect 1539 1818 1671 1822
rect 1675 1818 1767 1822
rect 1771 1818 1791 1822
rect 103 1817 1791 1818
rect 1797 1822 1807 1823
rect 1811 1822 2015 1826
rect 2019 1822 2103 1826
rect 2107 1822 2111 1826
rect 2115 1822 2191 1826
rect 2195 1822 2215 1826
rect 2219 1822 2279 1826
rect 2283 1822 2327 1826
rect 2331 1822 2367 1826
rect 2371 1822 2439 1826
rect 2443 1822 2455 1826
rect 2459 1822 2543 1826
rect 2547 1822 2631 1826
rect 2635 1822 2647 1826
rect 2651 1822 2719 1826
rect 2723 1822 2759 1826
rect 2763 1822 2807 1826
rect 2811 1822 2871 1826
rect 2875 1822 2895 1826
rect 2899 1822 2983 1826
rect 2987 1822 3463 1826
rect 3467 1822 3506 1826
rect 1797 1821 3506 1822
rect 1797 1817 1798 1821
rect 84 1749 85 1755
rect 91 1754 1779 1755
rect 91 1750 111 1754
rect 115 1750 439 1754
rect 443 1750 511 1754
rect 515 1750 535 1754
rect 539 1750 631 1754
rect 635 1750 639 1754
rect 643 1750 743 1754
rect 747 1750 759 1754
rect 763 1750 847 1754
rect 851 1750 887 1754
rect 891 1750 951 1754
rect 955 1750 1023 1754
rect 1027 1750 1055 1754
rect 1059 1750 1151 1754
rect 1155 1750 1159 1754
rect 1163 1750 1271 1754
rect 1275 1750 1279 1754
rect 1283 1750 1383 1754
rect 1387 1750 1407 1754
rect 1411 1750 1535 1754
rect 1539 1750 1671 1754
rect 1675 1750 1767 1754
rect 1771 1750 1779 1754
rect 91 1749 1779 1750
rect 1785 1751 1786 1755
rect 1785 1750 3494 1751
rect 1785 1749 1807 1750
rect 1778 1746 1807 1749
rect 1811 1746 2103 1750
rect 2107 1746 2143 1750
rect 2147 1746 2191 1750
rect 2195 1746 2231 1750
rect 2235 1746 2279 1750
rect 2283 1746 2319 1750
rect 2323 1746 2367 1750
rect 2371 1746 2407 1750
rect 2411 1746 2455 1750
rect 2459 1746 2495 1750
rect 2499 1746 2543 1750
rect 2547 1746 2583 1750
rect 2587 1746 2631 1750
rect 2635 1746 2671 1750
rect 2675 1746 2719 1750
rect 2723 1746 2759 1750
rect 2763 1746 2807 1750
rect 2811 1746 2847 1750
rect 2851 1746 2895 1750
rect 2899 1746 3463 1750
rect 3467 1746 3494 1750
rect 1778 1745 3494 1746
rect 96 1681 97 1687
rect 103 1686 1791 1687
rect 103 1682 111 1686
rect 115 1682 399 1686
rect 403 1682 439 1686
rect 443 1682 487 1686
rect 491 1682 535 1686
rect 539 1682 575 1686
rect 579 1682 639 1686
rect 643 1682 663 1686
rect 667 1682 743 1686
rect 747 1682 759 1686
rect 763 1682 847 1686
rect 851 1682 855 1686
rect 859 1682 951 1686
rect 955 1682 1047 1686
rect 1051 1682 1055 1686
rect 1059 1682 1143 1686
rect 1147 1682 1159 1686
rect 1163 1682 1271 1686
rect 1275 1682 1383 1686
rect 1387 1682 1767 1686
rect 1771 1682 1791 1686
rect 103 1681 1791 1682
rect 1797 1683 1798 1687
rect 1797 1682 3506 1683
rect 1797 1681 1807 1682
rect 1790 1678 1807 1681
rect 1811 1678 2103 1682
rect 2107 1678 2143 1682
rect 2147 1678 2191 1682
rect 2195 1678 2231 1682
rect 2235 1678 2279 1682
rect 2283 1678 2319 1682
rect 2323 1678 2367 1682
rect 2371 1678 2407 1682
rect 2411 1678 2455 1682
rect 2459 1678 2495 1682
rect 2499 1678 2543 1682
rect 2547 1678 2583 1682
rect 2587 1678 2631 1682
rect 2635 1678 2671 1682
rect 2675 1678 2719 1682
rect 2723 1678 2759 1682
rect 2763 1678 2807 1682
rect 2811 1678 2847 1682
rect 2851 1678 2895 1682
rect 2899 1678 3463 1682
rect 3467 1678 3506 1682
rect 1790 1677 3506 1678
rect 84 1613 85 1619
rect 91 1618 1779 1619
rect 91 1614 111 1618
rect 115 1614 279 1618
rect 283 1614 383 1618
rect 387 1614 399 1618
rect 403 1614 487 1618
rect 491 1614 495 1618
rect 499 1614 575 1618
rect 579 1614 607 1618
rect 611 1614 663 1618
rect 667 1614 719 1618
rect 723 1614 759 1618
rect 763 1614 831 1618
rect 835 1614 855 1618
rect 859 1614 943 1618
rect 947 1614 951 1618
rect 955 1614 1047 1618
rect 1051 1614 1055 1618
rect 1059 1614 1143 1618
rect 1147 1614 1167 1618
rect 1171 1614 1279 1618
rect 1283 1614 1767 1618
rect 1771 1614 1779 1618
rect 91 1613 1779 1614
rect 1785 1615 1786 1619
rect 1785 1614 3494 1615
rect 1785 1613 1807 1614
rect 1778 1610 1807 1613
rect 1811 1610 2063 1614
rect 2067 1610 2103 1614
rect 2107 1610 2159 1614
rect 2163 1610 2191 1614
rect 2195 1610 2255 1614
rect 2259 1610 2279 1614
rect 2283 1610 2359 1614
rect 2363 1610 2367 1614
rect 2371 1610 2455 1614
rect 2459 1610 2463 1614
rect 2467 1610 2543 1614
rect 2547 1610 2567 1614
rect 2571 1610 2631 1614
rect 2635 1610 2671 1614
rect 2675 1610 2719 1614
rect 2723 1610 2775 1614
rect 2779 1610 2807 1614
rect 2811 1610 2887 1614
rect 2891 1610 2895 1614
rect 2899 1610 3463 1614
rect 3467 1610 3494 1614
rect 1778 1609 3494 1610
rect 1790 1550 3506 1551
rect 1790 1547 1807 1550
rect 96 1541 97 1547
rect 103 1546 1791 1547
rect 103 1542 111 1546
rect 115 1542 183 1546
rect 187 1542 279 1546
rect 283 1542 327 1546
rect 331 1542 383 1546
rect 387 1542 471 1546
rect 475 1542 495 1546
rect 499 1542 607 1546
rect 611 1542 623 1546
rect 627 1542 719 1546
rect 723 1542 767 1546
rect 771 1542 831 1546
rect 835 1542 911 1546
rect 915 1542 943 1546
rect 947 1542 1047 1546
rect 1051 1542 1055 1546
rect 1059 1542 1167 1546
rect 1171 1542 1175 1546
rect 1179 1542 1279 1546
rect 1283 1542 1311 1546
rect 1315 1542 1447 1546
rect 1451 1542 1767 1546
rect 1771 1542 1791 1546
rect 103 1541 1791 1542
rect 1797 1546 1807 1547
rect 1811 1546 1919 1550
rect 1923 1546 2039 1550
rect 2043 1546 2063 1550
rect 2067 1546 2159 1550
rect 2163 1546 2167 1550
rect 2171 1546 2255 1550
rect 2259 1546 2295 1550
rect 2299 1546 2359 1550
rect 2363 1546 2423 1550
rect 2427 1546 2463 1550
rect 2467 1546 2551 1550
rect 2555 1546 2567 1550
rect 2571 1546 2671 1550
rect 2675 1546 2679 1550
rect 2683 1546 2775 1550
rect 2779 1546 2799 1550
rect 2803 1546 2887 1550
rect 2891 1546 2927 1550
rect 2931 1546 3055 1550
rect 3059 1546 3463 1550
rect 3467 1546 3506 1550
rect 1797 1545 3506 1546
rect 1797 1541 1798 1545
rect 84 1473 85 1479
rect 91 1478 1779 1479
rect 91 1474 111 1478
rect 115 1474 159 1478
rect 163 1474 183 1478
rect 187 1474 327 1478
rect 331 1474 375 1478
rect 379 1474 471 1478
rect 475 1474 583 1478
rect 587 1474 623 1478
rect 627 1474 767 1478
rect 771 1474 783 1478
rect 787 1474 911 1478
rect 915 1474 959 1478
rect 963 1474 1047 1478
rect 1051 1474 1127 1478
rect 1131 1474 1175 1478
rect 1179 1474 1279 1478
rect 1283 1474 1311 1478
rect 1315 1474 1431 1478
rect 1435 1474 1447 1478
rect 1451 1474 1591 1478
rect 1595 1474 1767 1478
rect 1771 1474 1779 1478
rect 91 1473 1779 1474
rect 1785 1478 3494 1479
rect 1785 1474 1807 1478
rect 1811 1474 1831 1478
rect 1835 1474 1919 1478
rect 1923 1474 1951 1478
rect 1955 1474 2039 1478
rect 2043 1474 2111 1478
rect 2115 1474 2167 1478
rect 2171 1474 2271 1478
rect 2275 1474 2295 1478
rect 2299 1474 2423 1478
rect 2427 1474 2431 1478
rect 2435 1474 2551 1478
rect 2555 1474 2591 1478
rect 2595 1474 2679 1478
rect 2683 1474 2735 1478
rect 2739 1474 2799 1478
rect 2803 1474 2871 1478
rect 2875 1474 2927 1478
rect 2931 1474 3007 1478
rect 3011 1474 3055 1478
rect 3059 1474 3135 1478
rect 3139 1474 3263 1478
rect 3267 1474 3367 1478
rect 3371 1474 3463 1478
rect 3467 1474 3494 1478
rect 1785 1473 3494 1474
rect 96 1405 97 1411
rect 103 1410 1791 1411
rect 103 1406 111 1410
rect 115 1406 135 1410
rect 139 1406 159 1410
rect 163 1406 303 1410
rect 307 1406 375 1410
rect 379 1406 495 1410
rect 499 1406 583 1410
rect 587 1406 679 1410
rect 683 1406 783 1410
rect 787 1406 855 1410
rect 859 1406 959 1410
rect 963 1406 1015 1410
rect 1019 1406 1127 1410
rect 1131 1406 1167 1410
rect 1171 1406 1279 1410
rect 1283 1406 1303 1410
rect 1307 1406 1431 1410
rect 1435 1406 1559 1410
rect 1563 1406 1591 1410
rect 1595 1406 1671 1410
rect 1675 1406 1767 1410
rect 1771 1406 1791 1410
rect 103 1405 1791 1406
rect 1797 1410 3506 1411
rect 1797 1406 1807 1410
rect 1811 1406 1831 1410
rect 1835 1406 1951 1410
rect 1955 1406 2007 1410
rect 2011 1406 2111 1410
rect 2115 1406 2199 1410
rect 2203 1406 2271 1410
rect 2275 1406 2383 1410
rect 2387 1406 2431 1410
rect 2435 1406 2559 1410
rect 2563 1406 2591 1410
rect 2595 1406 2719 1410
rect 2723 1406 2735 1410
rect 2739 1406 2863 1410
rect 2867 1406 2871 1410
rect 2875 1406 2999 1410
rect 3003 1406 3007 1410
rect 3011 1406 3127 1410
rect 3131 1406 3135 1410
rect 3139 1406 3255 1410
rect 3259 1406 3263 1410
rect 3267 1406 3367 1410
rect 3371 1406 3463 1410
rect 3467 1406 3506 1410
rect 1797 1405 3506 1406
rect 84 1337 85 1343
rect 91 1342 1779 1343
rect 91 1338 111 1342
rect 115 1338 135 1342
rect 139 1338 247 1342
rect 251 1338 303 1342
rect 307 1338 399 1342
rect 403 1338 495 1342
rect 499 1338 559 1342
rect 563 1338 679 1342
rect 683 1338 727 1342
rect 731 1338 855 1342
rect 859 1338 895 1342
rect 899 1338 1015 1342
rect 1019 1338 1063 1342
rect 1067 1338 1167 1342
rect 1171 1338 1223 1342
rect 1227 1338 1303 1342
rect 1307 1338 1375 1342
rect 1379 1338 1431 1342
rect 1435 1338 1535 1342
rect 1539 1338 1559 1342
rect 1563 1338 1671 1342
rect 1675 1338 1767 1342
rect 1771 1338 1779 1342
rect 91 1337 1779 1338
rect 1785 1339 1786 1343
rect 1785 1338 3494 1339
rect 1785 1337 1807 1338
rect 1778 1334 1807 1337
rect 1811 1334 1831 1338
rect 1835 1334 1967 1338
rect 1971 1334 2007 1338
rect 2011 1334 2143 1338
rect 2147 1334 2199 1338
rect 2203 1334 2327 1338
rect 2331 1334 2383 1338
rect 2387 1334 2511 1338
rect 2515 1334 2559 1338
rect 2563 1334 2687 1338
rect 2691 1334 2719 1338
rect 2723 1334 2863 1338
rect 2867 1334 2999 1338
rect 3003 1334 3039 1338
rect 3043 1334 3127 1338
rect 3131 1334 3215 1338
rect 3219 1334 3255 1338
rect 3259 1334 3367 1338
rect 3371 1334 3463 1338
rect 3467 1334 3494 1338
rect 1778 1333 3494 1334
rect 96 1269 97 1275
rect 103 1274 1791 1275
rect 103 1270 111 1274
rect 115 1270 135 1274
rect 139 1270 223 1274
rect 227 1270 247 1274
rect 251 1270 319 1274
rect 323 1270 399 1274
rect 403 1270 431 1274
rect 435 1270 551 1274
rect 555 1270 559 1274
rect 563 1270 679 1274
rect 683 1270 727 1274
rect 731 1270 823 1274
rect 827 1270 895 1274
rect 899 1270 975 1274
rect 979 1270 1063 1274
rect 1067 1270 1143 1274
rect 1147 1270 1223 1274
rect 1227 1270 1319 1274
rect 1323 1270 1375 1274
rect 1379 1270 1503 1274
rect 1507 1270 1535 1274
rect 1539 1270 1671 1274
rect 1675 1270 1767 1274
rect 1771 1270 1791 1274
rect 103 1269 1791 1270
rect 1797 1274 3506 1275
rect 1797 1270 1807 1274
rect 1811 1270 1831 1274
rect 1835 1270 1967 1274
rect 1971 1270 2095 1274
rect 2099 1270 2143 1274
rect 2147 1270 2327 1274
rect 2331 1270 2359 1274
rect 2363 1270 2511 1274
rect 2515 1270 2599 1274
rect 2603 1270 2687 1274
rect 2691 1270 2807 1274
rect 2811 1270 2863 1274
rect 2867 1270 3007 1274
rect 3011 1270 3039 1274
rect 3043 1270 3199 1274
rect 3203 1270 3215 1274
rect 3219 1270 3367 1274
rect 3371 1270 3463 1274
rect 3467 1270 3506 1274
rect 1797 1269 3506 1270
rect 84 1197 85 1203
rect 91 1202 1779 1203
rect 91 1198 111 1202
rect 115 1198 135 1202
rect 139 1198 223 1202
rect 227 1198 231 1202
rect 235 1198 319 1202
rect 323 1198 359 1202
rect 363 1198 431 1202
rect 435 1198 487 1202
rect 491 1198 551 1202
rect 555 1198 615 1202
rect 619 1198 679 1202
rect 683 1198 743 1202
rect 747 1198 823 1202
rect 827 1198 871 1202
rect 875 1198 975 1202
rect 979 1198 991 1202
rect 995 1198 1119 1202
rect 1123 1198 1143 1202
rect 1147 1198 1247 1202
rect 1251 1198 1319 1202
rect 1323 1198 1503 1202
rect 1507 1198 1671 1202
rect 1675 1198 1767 1202
rect 1771 1198 1779 1202
rect 91 1197 1779 1198
rect 1785 1202 3494 1203
rect 1785 1198 1807 1202
rect 1811 1198 1831 1202
rect 1835 1198 1935 1202
rect 1939 1198 2039 1202
rect 2043 1198 2095 1202
rect 2099 1198 2159 1202
rect 2163 1198 2287 1202
rect 2291 1198 2359 1202
rect 2363 1198 2423 1202
rect 2427 1198 2567 1202
rect 2571 1198 2599 1202
rect 2603 1198 2703 1202
rect 2707 1198 2807 1202
rect 2811 1198 2839 1202
rect 2843 1198 2975 1202
rect 2979 1198 3007 1202
rect 3011 1198 3111 1202
rect 3115 1198 3199 1202
rect 3203 1198 3247 1202
rect 3251 1198 3367 1202
rect 3371 1198 3463 1202
rect 3467 1198 3494 1202
rect 1785 1197 3494 1198
rect 96 1129 97 1135
rect 103 1134 1791 1135
rect 103 1130 111 1134
rect 115 1130 135 1134
rect 139 1130 231 1134
rect 235 1130 247 1134
rect 251 1130 359 1134
rect 363 1130 367 1134
rect 371 1130 487 1134
rect 491 1130 495 1134
rect 499 1130 615 1134
rect 619 1130 623 1134
rect 627 1130 743 1134
rect 747 1130 759 1134
rect 763 1130 871 1134
rect 875 1130 887 1134
rect 891 1130 991 1134
rect 995 1130 1015 1134
rect 1019 1130 1119 1134
rect 1123 1130 1143 1134
rect 1147 1130 1247 1134
rect 1251 1130 1271 1134
rect 1275 1130 1399 1134
rect 1403 1130 1767 1134
rect 1771 1130 1791 1134
rect 103 1129 1791 1130
rect 1797 1131 1798 1135
rect 1797 1130 3506 1131
rect 1797 1129 1807 1130
rect 1790 1126 1807 1129
rect 1811 1126 1935 1130
rect 1939 1126 1943 1130
rect 1947 1126 2039 1130
rect 2043 1126 2063 1130
rect 2067 1126 2159 1130
rect 2163 1126 2191 1130
rect 2195 1126 2287 1130
rect 2291 1126 2319 1130
rect 2323 1126 2423 1130
rect 2427 1126 2455 1130
rect 2459 1126 2567 1130
rect 2571 1126 2599 1130
rect 2603 1126 2703 1130
rect 2707 1126 2751 1130
rect 2755 1126 2839 1130
rect 2843 1126 2903 1130
rect 2907 1126 2975 1130
rect 2979 1126 3063 1130
rect 3067 1126 3111 1130
rect 3115 1126 3223 1130
rect 3227 1126 3247 1130
rect 3251 1126 3367 1130
rect 3371 1126 3463 1130
rect 3467 1126 3506 1130
rect 1790 1125 3506 1126
rect 84 1061 85 1067
rect 91 1066 1779 1067
rect 91 1062 111 1066
rect 115 1062 247 1066
rect 251 1062 367 1066
rect 371 1062 431 1066
rect 435 1062 495 1066
rect 499 1062 543 1066
rect 547 1062 623 1066
rect 627 1062 663 1066
rect 667 1062 759 1066
rect 763 1062 791 1066
rect 795 1062 887 1066
rect 891 1062 919 1066
rect 923 1062 1015 1066
rect 1019 1062 1039 1066
rect 1043 1062 1143 1066
rect 1147 1062 1159 1066
rect 1163 1062 1271 1066
rect 1275 1062 1279 1066
rect 1283 1062 1399 1066
rect 1403 1062 1407 1066
rect 1411 1062 1535 1066
rect 1539 1062 1767 1066
rect 1771 1062 1779 1066
rect 91 1061 1779 1062
rect 1785 1063 1786 1067
rect 1785 1062 3494 1063
rect 1785 1061 1807 1062
rect 1778 1058 1807 1061
rect 1811 1058 1847 1062
rect 1851 1058 1943 1062
rect 1947 1058 1983 1062
rect 1987 1058 2063 1062
rect 2067 1058 2119 1062
rect 2123 1058 2191 1062
rect 2195 1058 2255 1062
rect 2259 1058 2319 1062
rect 2323 1058 2391 1062
rect 2395 1058 2455 1062
rect 2459 1058 2543 1062
rect 2547 1058 2599 1062
rect 2603 1058 2703 1062
rect 2707 1058 2751 1062
rect 2755 1058 2863 1062
rect 2867 1058 2903 1062
rect 2907 1058 3031 1062
rect 3035 1058 3063 1062
rect 3067 1058 3207 1062
rect 3211 1058 3223 1062
rect 3227 1058 3367 1062
rect 3371 1058 3463 1062
rect 3467 1058 3494 1062
rect 1778 1057 3494 1058
rect 96 989 97 995
rect 103 994 1791 995
rect 103 990 111 994
rect 115 990 431 994
rect 435 990 543 994
rect 547 990 567 994
rect 571 990 663 994
rect 667 990 679 994
rect 683 990 791 994
rect 795 990 911 994
rect 915 990 919 994
rect 923 990 1031 994
rect 1035 990 1039 994
rect 1043 990 1143 994
rect 1147 990 1159 994
rect 1163 990 1255 994
rect 1259 990 1279 994
rect 1283 990 1359 994
rect 1363 990 1407 994
rect 1411 990 1471 994
rect 1475 990 1535 994
rect 1539 990 1583 994
rect 1587 990 1671 994
rect 1675 990 1767 994
rect 1771 990 1791 994
rect 103 989 1791 990
rect 1797 994 3506 995
rect 1797 990 1807 994
rect 1811 990 1831 994
rect 1835 990 1847 994
rect 1851 990 1975 994
rect 1979 990 1983 994
rect 1987 990 2119 994
rect 2123 990 2135 994
rect 2139 990 2255 994
rect 2259 990 2295 994
rect 2299 990 2391 994
rect 2395 990 2463 994
rect 2467 990 2543 994
rect 2547 990 2631 994
rect 2635 990 2703 994
rect 2707 990 2807 994
rect 2811 990 2863 994
rect 2867 990 2991 994
rect 2995 990 3031 994
rect 3035 990 3183 994
rect 3187 990 3207 994
rect 3211 990 3367 994
rect 3371 990 3463 994
rect 3467 990 3506 994
rect 1797 989 3506 990
rect 1778 930 3494 931
rect 1778 927 1807 930
rect 84 921 85 927
rect 91 926 1779 927
rect 91 922 111 926
rect 115 922 415 926
rect 419 922 559 926
rect 563 922 567 926
rect 571 922 679 926
rect 683 922 727 926
rect 731 922 791 926
rect 795 922 911 926
rect 915 922 1031 926
rect 1035 922 1119 926
rect 1123 922 1143 926
rect 1147 922 1255 926
rect 1259 922 1335 926
rect 1339 922 1359 926
rect 1363 922 1471 926
rect 1475 922 1559 926
rect 1563 922 1583 926
rect 1587 922 1671 926
rect 1675 922 1767 926
rect 1771 922 1779 926
rect 91 921 1779 922
rect 1785 926 1807 927
rect 1811 926 1831 930
rect 1835 926 1975 930
rect 1979 926 2127 930
rect 2131 926 2135 930
rect 2139 926 2215 930
rect 2219 926 2295 930
rect 2299 926 2303 930
rect 2307 926 2391 930
rect 2395 926 2463 930
rect 2467 926 2479 930
rect 2483 926 2567 930
rect 2571 926 2631 930
rect 2635 926 2655 930
rect 2659 926 2743 930
rect 2747 926 2807 930
rect 2811 926 2831 930
rect 2835 926 2991 930
rect 2995 926 3183 930
rect 3187 926 3367 930
rect 3371 926 3463 930
rect 3467 926 3494 930
rect 1785 925 3494 926
rect 1785 921 1786 925
rect 96 853 97 859
rect 103 858 1791 859
rect 103 854 111 858
rect 115 854 135 858
rect 139 854 231 858
rect 235 854 359 858
rect 363 854 415 858
rect 419 854 487 858
rect 491 854 559 858
rect 563 854 623 858
rect 627 854 727 858
rect 731 854 751 858
rect 755 854 879 858
rect 883 854 911 858
rect 915 854 1007 858
rect 1011 854 1119 858
rect 1123 854 1135 858
rect 1139 854 1271 858
rect 1275 854 1335 858
rect 1339 854 1559 858
rect 1563 854 1767 858
rect 1771 854 1791 858
rect 103 853 1791 854
rect 1797 858 3506 859
rect 1797 854 1807 858
rect 1811 854 2127 858
rect 2131 854 2159 858
rect 2163 854 2215 858
rect 2219 854 2247 858
rect 2251 854 2303 858
rect 2307 854 2335 858
rect 2339 854 2391 858
rect 2395 854 2423 858
rect 2427 854 2479 858
rect 2483 854 2527 858
rect 2531 854 2567 858
rect 2571 854 2639 858
rect 2643 854 2655 858
rect 2659 854 2743 858
rect 2747 854 2767 858
rect 2771 854 2831 858
rect 2835 854 2911 858
rect 2915 854 3063 858
rect 3067 854 3223 858
rect 3227 854 3367 858
rect 3371 854 3463 858
rect 3467 854 3506 858
rect 1797 853 3506 854
rect 84 785 85 791
rect 91 790 1779 791
rect 91 786 111 790
rect 115 786 135 790
rect 139 786 223 790
rect 227 786 231 790
rect 235 786 343 790
rect 347 786 359 790
rect 363 786 471 790
rect 475 786 487 790
rect 491 786 607 790
rect 611 786 623 790
rect 627 786 743 790
rect 747 786 751 790
rect 755 786 879 790
rect 883 786 887 790
rect 891 786 1007 790
rect 1011 786 1039 790
rect 1043 786 1135 790
rect 1139 786 1191 790
rect 1195 786 1271 790
rect 1275 786 1351 790
rect 1355 786 1767 790
rect 1771 786 1779 790
rect 91 785 1779 786
rect 1785 790 3494 791
rect 1785 786 1807 790
rect 1811 786 2063 790
rect 2067 786 2159 790
rect 2163 786 2175 790
rect 2179 786 2247 790
rect 2251 786 2295 790
rect 2299 786 2335 790
rect 2339 786 2423 790
rect 2427 786 2527 790
rect 2531 786 2559 790
rect 2563 786 2639 790
rect 2643 786 2711 790
rect 2715 786 2767 790
rect 2771 786 2871 790
rect 2875 786 2911 790
rect 2915 786 3039 790
rect 3043 786 3063 790
rect 3067 786 3215 790
rect 3219 786 3223 790
rect 3227 786 3367 790
rect 3371 786 3463 790
rect 3467 786 3494 790
rect 1785 785 3494 786
rect 1790 726 3506 727
rect 1790 723 1807 726
rect 96 717 97 723
rect 103 722 1791 723
rect 103 718 111 722
rect 115 718 135 722
rect 139 718 167 722
rect 171 718 223 722
rect 227 718 295 722
rect 299 718 343 722
rect 347 718 431 722
rect 435 718 471 722
rect 475 718 575 722
rect 579 718 607 722
rect 611 718 727 722
rect 731 718 743 722
rect 747 718 879 722
rect 883 718 887 722
rect 891 718 1031 722
rect 1035 718 1039 722
rect 1043 718 1183 722
rect 1187 718 1191 722
rect 1195 718 1343 722
rect 1347 718 1351 722
rect 1355 718 1503 722
rect 1507 718 1767 722
rect 1771 718 1791 722
rect 103 717 1791 718
rect 1797 722 1807 723
rect 1811 722 1927 726
rect 1931 722 2063 726
rect 2067 722 2071 726
rect 2075 722 2175 726
rect 2179 722 2231 726
rect 2235 722 2295 726
rect 2299 722 2391 726
rect 2395 722 2423 726
rect 2427 722 2551 726
rect 2555 722 2559 726
rect 2563 722 2703 726
rect 2707 722 2711 726
rect 2715 722 2847 726
rect 2851 722 2871 726
rect 2875 722 2983 726
rect 2987 722 3039 726
rect 3043 722 3119 726
rect 3123 722 3215 726
rect 3219 722 3255 726
rect 3259 722 3367 726
rect 3371 722 3463 726
rect 3467 722 3506 726
rect 1797 721 3506 722
rect 1797 717 1798 721
rect 84 649 85 655
rect 91 654 1779 655
rect 91 650 111 654
rect 115 650 167 654
rect 171 650 295 654
rect 299 650 431 654
rect 435 650 455 654
rect 459 650 559 654
rect 563 650 575 654
rect 579 650 679 654
rect 683 650 727 654
rect 731 650 799 654
rect 803 650 879 654
rect 883 650 927 654
rect 931 650 1031 654
rect 1035 650 1055 654
rect 1059 650 1183 654
rect 1187 650 1311 654
rect 1315 650 1343 654
rect 1347 650 1447 654
rect 1451 650 1503 654
rect 1507 650 1583 654
rect 1587 650 1767 654
rect 1771 650 1779 654
rect 91 649 1779 650
rect 1785 654 3494 655
rect 1785 650 1807 654
rect 1811 650 1831 654
rect 1835 650 1927 654
rect 1931 650 1967 654
rect 1971 650 2071 654
rect 2075 650 2135 654
rect 2139 650 2231 654
rect 2235 650 2311 654
rect 2315 650 2391 654
rect 2395 650 2487 654
rect 2491 650 2551 654
rect 2555 650 2655 654
rect 2659 650 2703 654
rect 2707 650 2815 654
rect 2819 650 2847 654
rect 2851 650 2959 654
rect 2963 650 2983 654
rect 2987 650 3103 654
rect 3107 650 3119 654
rect 3123 650 3247 654
rect 3251 650 3255 654
rect 3259 650 3367 654
rect 3371 650 3463 654
rect 3467 650 3494 654
rect 1785 649 3494 650
rect 1790 585 1791 591
rect 1797 590 3499 591
rect 1797 586 1807 590
rect 1811 586 1831 590
rect 1835 586 1967 590
rect 1971 586 2127 590
rect 2131 586 2135 590
rect 2139 586 2287 590
rect 2291 586 2311 590
rect 2315 586 2455 590
rect 2459 586 2487 590
rect 2491 586 2623 590
rect 2627 586 2655 590
rect 2659 586 2799 590
rect 2803 586 2815 590
rect 2819 586 2959 590
rect 2963 586 2983 590
rect 2987 586 3103 590
rect 3107 586 3167 590
rect 3171 586 3247 590
rect 3251 586 3359 590
rect 3363 586 3367 590
rect 3371 586 3463 590
rect 3467 586 3499 590
rect 1797 585 3499 586
rect 3505 585 3506 591
rect 1790 583 1798 585
rect 96 577 97 583
rect 103 582 1791 583
rect 103 578 111 582
rect 115 578 455 582
rect 459 578 559 582
rect 563 578 599 582
rect 603 578 679 582
rect 683 578 703 582
rect 707 578 799 582
rect 803 578 815 582
rect 819 578 927 582
rect 931 578 1039 582
rect 1043 578 1055 582
rect 1059 578 1151 582
rect 1155 578 1183 582
rect 1187 578 1255 582
rect 1259 578 1311 582
rect 1315 578 1359 582
rect 1363 578 1447 582
rect 1451 578 1471 582
rect 1475 578 1583 582
rect 1587 578 1671 582
rect 1675 578 1767 582
rect 1771 578 1791 582
rect 103 577 1791 578
rect 1797 577 1798 583
rect 84 513 85 519
rect 91 518 1779 519
rect 91 514 111 518
rect 115 514 303 518
rect 307 514 431 518
rect 435 514 567 518
rect 571 514 599 518
rect 603 514 703 518
rect 707 514 815 518
rect 819 514 847 518
rect 851 514 927 518
rect 931 514 983 518
rect 987 514 1039 518
rect 1043 514 1111 518
rect 1115 514 1151 518
rect 1155 514 1231 518
rect 1235 514 1255 518
rect 1259 514 1351 518
rect 1355 514 1359 518
rect 1363 514 1463 518
rect 1467 514 1471 518
rect 1475 514 1575 518
rect 1579 514 1583 518
rect 1587 514 1671 518
rect 1675 514 1767 518
rect 1771 514 1779 518
rect 91 513 1779 514
rect 1785 513 1786 519
rect 1778 511 1786 513
rect 1778 505 1779 511
rect 1785 510 3487 511
rect 1785 506 1807 510
rect 1811 506 1831 510
rect 1835 506 1967 510
rect 1971 506 2127 510
rect 2131 506 2287 510
rect 2291 506 2295 510
rect 2299 506 2455 510
rect 2459 506 2479 510
rect 2483 506 2623 510
rect 2627 506 2679 510
rect 2683 506 2799 510
rect 2803 506 2887 510
rect 2891 506 2983 510
rect 2987 506 3111 510
rect 3115 506 3167 510
rect 3171 506 3335 510
rect 3339 506 3359 510
rect 3363 506 3463 510
rect 3467 506 3487 510
rect 1785 505 3487 506
rect 3493 505 3494 511
rect 96 441 97 447
rect 103 446 1791 447
rect 103 442 111 446
rect 115 442 135 446
rect 139 442 255 446
rect 259 442 303 446
rect 307 442 415 446
rect 419 442 431 446
rect 435 442 567 446
rect 571 442 583 446
rect 587 442 703 446
rect 707 442 743 446
rect 747 442 847 446
rect 851 442 903 446
rect 907 442 983 446
rect 987 442 1047 446
rect 1051 442 1111 446
rect 1115 442 1183 446
rect 1187 442 1231 446
rect 1235 442 1311 446
rect 1315 442 1351 446
rect 1355 442 1439 446
rect 1443 442 1463 446
rect 1467 442 1567 446
rect 1571 442 1575 446
rect 1579 442 1671 446
rect 1675 442 1767 446
rect 1771 442 1791 446
rect 103 441 1791 442
rect 1797 446 3506 447
rect 1797 442 1807 446
rect 1811 442 1831 446
rect 1835 442 1959 446
rect 1963 442 1967 446
rect 1971 442 2111 446
rect 2115 442 2127 446
rect 2131 442 2271 446
rect 2275 442 2295 446
rect 2299 442 2455 446
rect 2459 442 2479 446
rect 2483 442 2655 446
rect 2659 442 2679 446
rect 2683 442 2871 446
rect 2875 442 2887 446
rect 2891 442 3103 446
rect 3107 442 3111 446
rect 3115 442 3335 446
rect 3339 442 3463 446
rect 3467 442 3506 446
rect 1797 441 3506 442
rect 84 373 85 379
rect 91 378 1779 379
rect 91 374 111 378
rect 115 374 135 378
rect 139 374 223 378
rect 227 374 255 378
rect 259 374 343 378
rect 347 374 415 378
rect 419 374 471 378
rect 475 374 583 378
rect 587 374 599 378
rect 603 374 719 378
rect 723 374 743 378
rect 747 374 839 378
rect 843 374 903 378
rect 907 374 959 378
rect 963 374 1047 378
rect 1051 374 1079 378
rect 1083 374 1183 378
rect 1187 374 1207 378
rect 1211 374 1311 378
rect 1315 374 1439 378
rect 1443 374 1567 378
rect 1571 374 1671 378
rect 1675 374 1767 378
rect 1771 374 1779 378
rect 91 373 1779 374
rect 1785 378 3494 379
rect 1785 374 1807 378
rect 1811 374 1831 378
rect 1835 374 1927 378
rect 1931 374 1959 378
rect 1963 374 2039 378
rect 2043 374 2111 378
rect 2115 374 2159 378
rect 2163 374 2271 378
rect 2275 374 2287 378
rect 2291 374 2423 378
rect 2427 374 2455 378
rect 2459 374 2583 378
rect 2587 374 2655 378
rect 2659 374 2759 378
rect 2763 374 2871 378
rect 2875 374 2951 378
rect 2955 374 3103 378
rect 3107 374 3151 378
rect 3155 374 3335 378
rect 3339 374 3359 378
rect 3363 374 3463 378
rect 3467 374 3494 378
rect 1785 373 3494 374
rect 1790 314 3506 315
rect 1790 311 1807 314
rect 96 305 97 311
rect 103 310 1791 311
rect 103 306 111 310
rect 115 306 135 310
rect 139 306 223 310
rect 227 306 263 310
rect 267 306 343 310
rect 347 306 375 310
rect 379 306 471 310
rect 475 306 487 310
rect 491 306 599 310
rect 603 306 711 310
rect 715 306 719 310
rect 723 306 815 310
rect 819 306 839 310
rect 843 306 919 310
rect 923 306 959 310
rect 963 306 1023 310
rect 1027 306 1079 310
rect 1083 306 1127 310
rect 1131 306 1207 310
rect 1211 306 1239 310
rect 1243 306 1767 310
rect 1771 306 1791 310
rect 103 305 1791 306
rect 1797 310 1807 311
rect 1811 310 1927 314
rect 1931 310 2039 314
rect 2043 310 2159 314
rect 2163 310 2223 314
rect 2227 310 2287 314
rect 2291 310 2311 314
rect 2315 310 2399 314
rect 2403 310 2423 314
rect 2427 310 2487 314
rect 2491 310 2575 314
rect 2579 310 2583 314
rect 2587 310 2679 314
rect 2683 310 2759 314
rect 2763 310 2799 314
rect 2803 310 2927 314
rect 2931 310 2951 314
rect 2955 310 3071 314
rect 3075 310 3151 314
rect 3155 310 3223 314
rect 3227 310 3359 314
rect 3363 310 3367 314
rect 3371 310 3463 314
rect 3467 310 3506 314
rect 1797 309 3506 310
rect 1797 305 1798 309
rect 84 237 85 243
rect 91 242 1779 243
rect 91 238 111 242
rect 115 238 263 242
rect 267 238 375 242
rect 379 238 447 242
rect 451 238 487 242
rect 491 238 535 242
rect 539 238 599 242
rect 603 238 623 242
rect 627 238 711 242
rect 715 238 807 242
rect 811 238 815 242
rect 819 238 903 242
rect 907 238 919 242
rect 923 238 999 242
rect 1003 238 1023 242
rect 1027 238 1103 242
rect 1107 238 1127 242
rect 1131 238 1207 242
rect 1211 238 1239 242
rect 1243 238 1311 242
rect 1315 238 1767 242
rect 1771 238 1779 242
rect 91 237 1779 238
rect 1785 242 3494 243
rect 1785 238 1807 242
rect 1811 238 2143 242
rect 2147 238 2223 242
rect 2227 238 2263 242
rect 2267 238 2311 242
rect 2315 238 2383 242
rect 2387 238 2399 242
rect 2403 238 2487 242
rect 2491 238 2511 242
rect 2515 238 2575 242
rect 2579 238 2639 242
rect 2643 238 2679 242
rect 2683 238 2767 242
rect 2771 238 2799 242
rect 2803 238 2895 242
rect 2899 238 2927 242
rect 2931 238 3015 242
rect 3019 238 3071 242
rect 3075 238 3135 242
rect 3139 238 3223 242
rect 3227 238 3263 242
rect 3267 238 3367 242
rect 3371 238 3463 242
rect 3467 238 3494 242
rect 1785 237 3494 238
rect 1790 154 3506 155
rect 1790 151 1807 154
rect 96 145 97 151
rect 103 150 1791 151
rect 103 146 111 150
rect 115 146 263 150
rect 267 146 351 150
rect 355 146 439 150
rect 443 146 447 150
rect 451 146 527 150
rect 531 146 535 150
rect 539 146 615 150
rect 619 146 623 150
rect 627 146 703 150
rect 707 146 711 150
rect 715 146 791 150
rect 795 146 807 150
rect 811 146 879 150
rect 883 146 903 150
rect 907 146 967 150
rect 971 146 999 150
rect 1003 146 1055 150
rect 1059 146 1103 150
rect 1107 146 1143 150
rect 1147 146 1207 150
rect 1211 146 1231 150
rect 1235 146 1311 150
rect 1315 146 1319 150
rect 1323 146 1407 150
rect 1411 146 1495 150
rect 1499 146 1583 150
rect 1587 146 1671 150
rect 1675 146 1767 150
rect 1771 146 1791 150
rect 103 145 1791 146
rect 1797 150 1807 151
rect 1811 150 1831 154
rect 1835 150 1919 154
rect 1923 150 2007 154
rect 2011 150 2095 154
rect 2099 150 2143 154
rect 2147 150 2183 154
rect 2187 150 2263 154
rect 2267 150 2295 154
rect 2299 150 2383 154
rect 2387 150 2407 154
rect 2411 150 2511 154
rect 2515 150 2615 154
rect 2619 150 2639 154
rect 2643 150 2719 154
rect 2723 150 2767 154
rect 2771 150 2815 154
rect 2819 150 2895 154
rect 2899 150 2911 154
rect 2915 150 3007 154
rect 3011 150 3015 154
rect 3019 150 3103 154
rect 3107 150 3135 154
rect 3139 150 3191 154
rect 3195 150 3263 154
rect 3267 150 3279 154
rect 3283 150 3367 154
rect 3371 150 3463 154
rect 3467 150 3506 154
rect 1797 149 3506 150
rect 1797 145 1798 149
rect 1778 90 3494 91
rect 1778 87 1807 90
rect 84 81 85 87
rect 91 86 1779 87
rect 91 82 111 86
rect 115 82 263 86
rect 267 82 351 86
rect 355 82 439 86
rect 443 82 527 86
rect 531 82 615 86
rect 619 82 703 86
rect 707 82 791 86
rect 795 82 879 86
rect 883 82 967 86
rect 971 82 1055 86
rect 1059 82 1143 86
rect 1147 82 1231 86
rect 1235 82 1319 86
rect 1323 82 1407 86
rect 1411 82 1495 86
rect 1499 82 1583 86
rect 1587 82 1671 86
rect 1675 82 1767 86
rect 1771 82 1779 86
rect 91 81 1779 82
rect 1785 86 1807 87
rect 1811 86 1831 90
rect 1835 86 1919 90
rect 1923 86 2007 90
rect 2011 86 2095 90
rect 2099 86 2183 90
rect 2187 86 2295 90
rect 2299 86 2407 90
rect 2411 86 2511 90
rect 2515 86 2615 90
rect 2619 86 2719 90
rect 2723 86 2815 90
rect 2819 86 2911 90
rect 2915 86 3007 90
rect 3011 86 3103 90
rect 3107 86 3191 90
rect 3195 86 3279 90
rect 3283 86 3367 90
rect 3371 86 3463 90
rect 3467 86 3494 90
rect 1785 85 3494 86
rect 1785 81 1786 85
<< m5c >>
rect 97 3501 103 3507
rect 1791 3501 1797 3507
rect 1791 3489 1797 3495
rect 3499 3489 3505 3495
rect 85 3433 91 3439
rect 1779 3433 1785 3439
rect 1779 3425 1785 3431
rect 3487 3425 3493 3431
rect 97 3361 103 3367
rect 1791 3361 1797 3367
rect 85 3289 91 3295
rect 1779 3289 1785 3295
rect 1791 3225 1797 3231
rect 3499 3225 3505 3231
rect 97 3217 103 3223
rect 1791 3217 1797 3223
rect 1779 3161 1785 3167
rect 3487 3161 3493 3167
rect 85 3153 91 3159
rect 1779 3153 1785 3159
rect 97 3085 103 3091
rect 1791 3085 1797 3091
rect 85 3013 91 3019
rect 1779 3013 1785 3019
rect 97 2937 103 2943
rect 1791 2937 1797 2943
rect 85 2865 91 2871
rect 1779 2865 1785 2871
rect 1791 2801 1797 2807
rect 3499 2801 3505 2807
rect 97 2789 103 2795
rect 1791 2789 1797 2795
rect 85 2717 91 2723
rect 1779 2717 1785 2723
rect 97 2645 103 2651
rect 1791 2645 1797 2651
rect 85 2573 91 2579
rect 1779 2573 1785 2579
rect 97 2501 103 2507
rect 1791 2501 1797 2507
rect 85 2437 91 2443
rect 1779 2437 1785 2443
rect 97 2369 103 2375
rect 1791 2369 1797 2375
rect 85 2297 91 2303
rect 1779 2297 1785 2303
rect 97 2229 103 2235
rect 1791 2229 1797 2235
rect 1779 2169 1785 2175
rect 3487 2169 3493 2175
rect 85 2157 91 2163
rect 1779 2157 1785 2163
rect 1791 2097 1797 2103
rect 3499 2097 3505 2103
rect 97 2089 103 2095
rect 1791 2089 1797 2095
rect 1779 2029 1785 2035
rect 3487 2029 3493 2035
rect 85 2017 91 2023
rect 1779 2017 1785 2023
rect 1791 1961 1797 1967
rect 3499 1961 3505 1967
rect 97 1949 103 1955
rect 1791 1949 1797 1955
rect 1779 1893 1785 1899
rect 3487 1893 3493 1899
rect 85 1885 91 1891
rect 1779 1885 1785 1891
rect 97 1817 103 1823
rect 1791 1817 1797 1823
rect 85 1749 91 1755
rect 1779 1749 1785 1755
rect 97 1681 103 1687
rect 1791 1681 1797 1687
rect 85 1613 91 1619
rect 1779 1613 1785 1619
rect 97 1541 103 1547
rect 1791 1541 1797 1547
rect 85 1473 91 1479
rect 1779 1473 1785 1479
rect 97 1405 103 1411
rect 1791 1405 1797 1411
rect 85 1337 91 1343
rect 1779 1337 1785 1343
rect 97 1269 103 1275
rect 1791 1269 1797 1275
rect 85 1197 91 1203
rect 1779 1197 1785 1203
rect 97 1129 103 1135
rect 1791 1129 1797 1135
rect 85 1061 91 1067
rect 1779 1061 1785 1067
rect 97 989 103 995
rect 1791 989 1797 995
rect 85 921 91 927
rect 1779 921 1785 927
rect 97 853 103 859
rect 1791 853 1797 859
rect 85 785 91 791
rect 1779 785 1785 791
rect 97 717 103 723
rect 1791 717 1797 723
rect 85 649 91 655
rect 1779 649 1785 655
rect 1791 585 1797 591
rect 3499 585 3505 591
rect 97 577 103 583
rect 1791 577 1797 583
rect 85 513 91 519
rect 1779 513 1785 519
rect 1779 505 1785 511
rect 3487 505 3493 511
rect 97 441 103 447
rect 1791 441 1797 447
rect 85 373 91 379
rect 1779 373 1785 379
rect 97 305 103 311
rect 1791 305 1797 311
rect 85 237 91 243
rect 1779 237 1785 243
rect 97 145 103 151
rect 1791 145 1797 151
rect 85 81 91 87
rect 1779 81 1785 87
<< m5 >>
rect 84 3439 92 3528
rect 84 3433 85 3439
rect 91 3433 92 3439
rect 84 3295 92 3433
rect 84 3289 85 3295
rect 91 3289 92 3295
rect 84 3159 92 3289
rect 84 3153 85 3159
rect 91 3153 92 3159
rect 84 3019 92 3153
rect 84 3013 85 3019
rect 91 3013 92 3019
rect 84 2871 92 3013
rect 84 2865 85 2871
rect 91 2865 92 2871
rect 84 2723 92 2865
rect 84 2717 85 2723
rect 91 2717 92 2723
rect 84 2579 92 2717
rect 84 2573 85 2579
rect 91 2573 92 2579
rect 84 2443 92 2573
rect 84 2437 85 2443
rect 91 2437 92 2443
rect 84 2303 92 2437
rect 84 2297 85 2303
rect 91 2297 92 2303
rect 84 2163 92 2297
rect 84 2157 85 2163
rect 91 2157 92 2163
rect 84 2023 92 2157
rect 84 2017 85 2023
rect 91 2017 92 2023
rect 84 1891 92 2017
rect 84 1885 85 1891
rect 91 1885 92 1891
rect 84 1755 92 1885
rect 84 1749 85 1755
rect 91 1749 92 1755
rect 84 1619 92 1749
rect 84 1613 85 1619
rect 91 1613 92 1619
rect 84 1479 92 1613
rect 84 1473 85 1479
rect 91 1473 92 1479
rect 84 1343 92 1473
rect 84 1337 85 1343
rect 91 1337 92 1343
rect 84 1203 92 1337
rect 84 1197 85 1203
rect 91 1197 92 1203
rect 84 1067 92 1197
rect 84 1061 85 1067
rect 91 1061 92 1067
rect 84 927 92 1061
rect 84 921 85 927
rect 91 921 92 927
rect 84 791 92 921
rect 84 785 85 791
rect 91 785 92 791
rect 84 655 92 785
rect 84 649 85 655
rect 91 649 92 655
rect 84 519 92 649
rect 84 513 85 519
rect 91 513 92 519
rect 84 379 92 513
rect 84 373 85 379
rect 91 373 92 379
rect 84 243 92 373
rect 84 237 85 243
rect 91 237 92 243
rect 84 87 92 237
rect 84 81 85 87
rect 91 81 92 87
rect 84 72 92 81
rect 96 3507 104 3528
rect 96 3501 97 3507
rect 103 3501 104 3507
rect 96 3367 104 3501
rect 96 3361 97 3367
rect 103 3361 104 3367
rect 96 3223 104 3361
rect 96 3217 97 3223
rect 103 3217 104 3223
rect 96 3091 104 3217
rect 96 3085 97 3091
rect 103 3085 104 3091
rect 96 2943 104 3085
rect 96 2937 97 2943
rect 103 2937 104 2943
rect 96 2795 104 2937
rect 96 2789 97 2795
rect 103 2789 104 2795
rect 96 2651 104 2789
rect 96 2645 97 2651
rect 103 2645 104 2651
rect 96 2507 104 2645
rect 96 2501 97 2507
rect 103 2501 104 2507
rect 96 2375 104 2501
rect 96 2369 97 2375
rect 103 2369 104 2375
rect 96 2235 104 2369
rect 96 2229 97 2235
rect 103 2229 104 2235
rect 96 2095 104 2229
rect 96 2089 97 2095
rect 103 2089 104 2095
rect 96 1955 104 2089
rect 96 1949 97 1955
rect 103 1949 104 1955
rect 96 1823 104 1949
rect 96 1817 97 1823
rect 103 1817 104 1823
rect 96 1687 104 1817
rect 96 1681 97 1687
rect 103 1681 104 1687
rect 96 1547 104 1681
rect 96 1541 97 1547
rect 103 1541 104 1547
rect 96 1411 104 1541
rect 96 1405 97 1411
rect 103 1405 104 1411
rect 96 1275 104 1405
rect 96 1269 97 1275
rect 103 1269 104 1275
rect 96 1135 104 1269
rect 96 1129 97 1135
rect 103 1129 104 1135
rect 96 995 104 1129
rect 96 989 97 995
rect 103 989 104 995
rect 96 859 104 989
rect 96 853 97 859
rect 103 853 104 859
rect 96 723 104 853
rect 96 717 97 723
rect 103 717 104 723
rect 96 583 104 717
rect 96 577 97 583
rect 103 577 104 583
rect 96 447 104 577
rect 96 441 97 447
rect 103 441 104 447
rect 96 311 104 441
rect 96 305 97 311
rect 103 305 104 311
rect 96 151 104 305
rect 96 145 97 151
rect 103 145 104 151
rect 96 72 104 145
rect 1778 3439 1786 3528
rect 1778 3433 1779 3439
rect 1785 3433 1786 3439
rect 1778 3431 1786 3433
rect 1778 3425 1779 3431
rect 1785 3425 1786 3431
rect 1778 3295 1786 3425
rect 1778 3289 1779 3295
rect 1785 3289 1786 3295
rect 1778 3167 1786 3289
rect 1778 3161 1779 3167
rect 1785 3161 1786 3167
rect 1778 3159 1786 3161
rect 1778 3153 1779 3159
rect 1785 3153 1786 3159
rect 1778 3019 1786 3153
rect 1778 3013 1779 3019
rect 1785 3013 1786 3019
rect 1778 2871 1786 3013
rect 1778 2865 1779 2871
rect 1785 2865 1786 2871
rect 1778 2723 1786 2865
rect 1778 2717 1779 2723
rect 1785 2717 1786 2723
rect 1778 2579 1786 2717
rect 1778 2573 1779 2579
rect 1785 2573 1786 2579
rect 1778 2443 1786 2573
rect 1778 2437 1779 2443
rect 1785 2437 1786 2443
rect 1778 2303 1786 2437
rect 1778 2297 1779 2303
rect 1785 2297 1786 2303
rect 1778 2175 1786 2297
rect 1778 2169 1779 2175
rect 1785 2169 1786 2175
rect 1778 2163 1786 2169
rect 1778 2157 1779 2163
rect 1785 2157 1786 2163
rect 1778 2035 1786 2157
rect 1778 2029 1779 2035
rect 1785 2029 1786 2035
rect 1778 2023 1786 2029
rect 1778 2017 1779 2023
rect 1785 2017 1786 2023
rect 1778 1899 1786 2017
rect 1778 1893 1779 1899
rect 1785 1893 1786 1899
rect 1778 1891 1786 1893
rect 1778 1885 1779 1891
rect 1785 1885 1786 1891
rect 1778 1755 1786 1885
rect 1778 1749 1779 1755
rect 1785 1749 1786 1755
rect 1778 1619 1786 1749
rect 1778 1613 1779 1619
rect 1785 1613 1786 1619
rect 1778 1479 1786 1613
rect 1778 1473 1779 1479
rect 1785 1473 1786 1479
rect 1778 1343 1786 1473
rect 1778 1337 1779 1343
rect 1785 1337 1786 1343
rect 1778 1203 1786 1337
rect 1778 1197 1779 1203
rect 1785 1197 1786 1203
rect 1778 1067 1786 1197
rect 1778 1061 1779 1067
rect 1785 1061 1786 1067
rect 1778 927 1786 1061
rect 1778 921 1779 927
rect 1785 921 1786 927
rect 1778 791 1786 921
rect 1778 785 1779 791
rect 1785 785 1786 791
rect 1778 655 1786 785
rect 1778 649 1779 655
rect 1785 649 1786 655
rect 1778 519 1786 649
rect 1778 513 1779 519
rect 1785 513 1786 519
rect 1778 511 1786 513
rect 1778 505 1779 511
rect 1785 505 1786 511
rect 1778 379 1786 505
rect 1778 373 1779 379
rect 1785 373 1786 379
rect 1778 243 1786 373
rect 1778 237 1779 243
rect 1785 237 1786 243
rect 1778 87 1786 237
rect 1778 81 1779 87
rect 1785 81 1786 87
rect 1778 72 1786 81
rect 1790 3507 1798 3528
rect 1790 3501 1791 3507
rect 1797 3501 1798 3507
rect 1790 3495 1798 3501
rect 1790 3489 1791 3495
rect 1797 3489 1798 3495
rect 1790 3367 1798 3489
rect 1790 3361 1791 3367
rect 1797 3361 1798 3367
rect 1790 3231 1798 3361
rect 1790 3225 1791 3231
rect 1797 3225 1798 3231
rect 1790 3223 1798 3225
rect 1790 3217 1791 3223
rect 1797 3217 1798 3223
rect 1790 3091 1798 3217
rect 1790 3085 1791 3091
rect 1797 3085 1798 3091
rect 1790 2943 1798 3085
rect 1790 2937 1791 2943
rect 1797 2937 1798 2943
rect 1790 2807 1798 2937
rect 1790 2801 1791 2807
rect 1797 2801 1798 2807
rect 1790 2795 1798 2801
rect 1790 2789 1791 2795
rect 1797 2789 1798 2795
rect 1790 2651 1798 2789
rect 1790 2645 1791 2651
rect 1797 2645 1798 2651
rect 1790 2507 1798 2645
rect 1790 2501 1791 2507
rect 1797 2501 1798 2507
rect 1790 2375 1798 2501
rect 1790 2369 1791 2375
rect 1797 2369 1798 2375
rect 1790 2235 1798 2369
rect 1790 2229 1791 2235
rect 1797 2229 1798 2235
rect 1790 2103 1798 2229
rect 1790 2097 1791 2103
rect 1797 2097 1798 2103
rect 1790 2095 1798 2097
rect 1790 2089 1791 2095
rect 1797 2089 1798 2095
rect 1790 1967 1798 2089
rect 1790 1961 1791 1967
rect 1797 1961 1798 1967
rect 1790 1955 1798 1961
rect 1790 1949 1791 1955
rect 1797 1949 1798 1955
rect 1790 1823 1798 1949
rect 1790 1817 1791 1823
rect 1797 1817 1798 1823
rect 1790 1687 1798 1817
rect 1790 1681 1791 1687
rect 1797 1681 1798 1687
rect 1790 1547 1798 1681
rect 1790 1541 1791 1547
rect 1797 1541 1798 1547
rect 1790 1411 1798 1541
rect 1790 1405 1791 1411
rect 1797 1405 1798 1411
rect 1790 1275 1798 1405
rect 1790 1269 1791 1275
rect 1797 1269 1798 1275
rect 1790 1135 1798 1269
rect 1790 1129 1791 1135
rect 1797 1129 1798 1135
rect 1790 995 1798 1129
rect 1790 989 1791 995
rect 1797 989 1798 995
rect 1790 859 1798 989
rect 1790 853 1791 859
rect 1797 853 1798 859
rect 1790 723 1798 853
rect 1790 717 1791 723
rect 1797 717 1798 723
rect 1790 591 1798 717
rect 1790 585 1791 591
rect 1797 585 1798 591
rect 1790 583 1798 585
rect 1790 577 1791 583
rect 1797 577 1798 583
rect 1790 447 1798 577
rect 1790 441 1791 447
rect 1797 441 1798 447
rect 1790 311 1798 441
rect 1790 305 1791 311
rect 1797 305 1798 311
rect 1790 151 1798 305
rect 1790 145 1791 151
rect 1797 145 1798 151
rect 1790 72 1798 145
rect 3486 3431 3494 3528
rect 3486 3425 3487 3431
rect 3493 3425 3494 3431
rect 3486 3167 3494 3425
rect 3486 3161 3487 3167
rect 3493 3161 3494 3167
rect 3486 2175 3494 3161
rect 3486 2169 3487 2175
rect 3493 2169 3494 2175
rect 3486 2035 3494 2169
rect 3486 2029 3487 2035
rect 3493 2029 3494 2035
rect 3486 1899 3494 2029
rect 3486 1893 3487 1899
rect 3493 1893 3494 1899
rect 3486 511 3494 1893
rect 3486 505 3487 511
rect 3493 505 3494 511
rect 3486 72 3494 505
rect 3498 3495 3506 3528
rect 3498 3489 3499 3495
rect 3505 3489 3506 3495
rect 3498 3231 3506 3489
rect 3498 3225 3499 3231
rect 3505 3225 3506 3231
rect 3498 2807 3506 3225
rect 3498 2801 3499 2807
rect 3505 2801 3506 2807
rect 3498 2103 3506 2801
rect 3498 2097 3499 2103
rect 3505 2097 3506 2103
rect 3498 1967 3506 2097
rect 3498 1961 3499 1967
rect 3505 1961 3506 1967
rect 3498 591 3506 1961
rect 3498 585 3499 591
rect 3505 585 3506 591
rect 3498 72 3506 585
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__195
timestamp 1731220323
transform 1 0 3456 0 1 3448
box 7 3 12 24
use welltap_svt  __well_tap__194
timestamp 1731220323
transform 1 0 1800 0 1 3448
box 7 3 12 24
use welltap_svt  __well_tap__193
timestamp 1731220323
transform 1 0 3456 0 -1 3408
box 7 3 12 24
use welltap_svt  __well_tap__192
timestamp 1731220323
transform 1 0 1800 0 -1 3408
box 7 3 12 24
use welltap_svt  __well_tap__191
timestamp 1731220323
transform 1 0 3456 0 1 3316
box 7 3 12 24
use welltap_svt  __well_tap__190
timestamp 1731220323
transform 1 0 1800 0 1 3316
box 7 3 12 24
use welltap_svt  __well_tap__189
timestamp 1731220323
transform 1 0 3456 0 -1 3276
box 7 3 12 24
use welltap_svt  __well_tap__188
timestamp 1731220323
transform 1 0 1800 0 -1 3276
box 7 3 12 24
use welltap_svt  __well_tap__187
timestamp 1731220323
transform 1 0 3456 0 1 3184
box 7 3 12 24
use welltap_svt  __well_tap__186
timestamp 1731220323
transform 1 0 1800 0 1 3184
box 7 3 12 24
use welltap_svt  __well_tap__185
timestamp 1731220323
transform 1 0 3456 0 -1 3144
box 7 3 12 24
use welltap_svt  __well_tap__184
timestamp 1731220323
transform 1 0 1800 0 -1 3144
box 7 3 12 24
use welltap_svt  __well_tap__183
timestamp 1731220323
transform 1 0 3456 0 1 3048
box 7 3 12 24
use welltap_svt  __well_tap__182
timestamp 1731220323
transform 1 0 1800 0 1 3048
box 7 3 12 24
use welltap_svt  __well_tap__181
timestamp 1731220323
transform 1 0 3456 0 -1 2992
box 7 3 12 24
use welltap_svt  __well_tap__180
timestamp 1731220323
transform 1 0 1800 0 -1 2992
box 7 3 12 24
use welltap_svt  __well_tap__179
timestamp 1731220323
transform 1 0 3456 0 1 2892
box 7 3 12 24
use welltap_svt  __well_tap__178
timestamp 1731220323
transform 1 0 1800 0 1 2892
box 7 3 12 24
use welltap_svt  __well_tap__177
timestamp 1731220323
transform 1 0 3456 0 -1 2852
box 7 3 12 24
use welltap_svt  __well_tap__176
timestamp 1731220323
transform 1 0 1800 0 -1 2852
box 7 3 12 24
use welltap_svt  __well_tap__175
timestamp 1731220323
transform 1 0 3456 0 1 2760
box 7 3 12 24
use welltap_svt  __well_tap__174
timestamp 1731220323
transform 1 0 1800 0 1 2760
box 7 3 12 24
use welltap_svt  __well_tap__173
timestamp 1731220323
transform 1 0 3456 0 -1 2704
box 7 3 12 24
use welltap_svt  __well_tap__172
timestamp 1731220323
transform 1 0 1800 0 -1 2704
box 7 3 12 24
use welltap_svt  __well_tap__171
timestamp 1731220323
transform 1 0 3456 0 1 2604
box 7 3 12 24
use welltap_svt  __well_tap__170
timestamp 1731220323
transform 1 0 1800 0 1 2604
box 7 3 12 24
use welltap_svt  __well_tap__169
timestamp 1731220323
transform 1 0 3456 0 -1 2552
box 7 3 12 24
use welltap_svt  __well_tap__168
timestamp 1731220323
transform 1 0 1800 0 -1 2552
box 7 3 12 24
use welltap_svt  __well_tap__167
timestamp 1731220323
transform 1 0 3456 0 1 2464
box 7 3 12 24
use welltap_svt  __well_tap__166
timestamp 1731220323
transform 1 0 1800 0 1 2464
box 7 3 12 24
use welltap_svt  __well_tap__165
timestamp 1731220323
transform 1 0 3456 0 -1 2416
box 7 3 12 24
use welltap_svt  __well_tap__164
timestamp 1731220323
transform 1 0 1800 0 -1 2416
box 7 3 12 24
use welltap_svt  __well_tap__163
timestamp 1731220323
transform 1 0 3456 0 1 2328
box 7 3 12 24
use welltap_svt  __well_tap__162
timestamp 1731220323
transform 1 0 1800 0 1 2328
box 7 3 12 24
use welltap_svt  __well_tap__161
timestamp 1731220323
transform 1 0 3456 0 -1 2280
box 7 3 12 24
use welltap_svt  __well_tap__160
timestamp 1731220323
transform 1 0 1800 0 -1 2280
box 7 3 12 24
use welltap_svt  __well_tap__159
timestamp 1731220323
transform 1 0 3456 0 1 2192
box 7 3 12 24
use welltap_svt  __well_tap__158
timestamp 1731220323
transform 1 0 1800 0 1 2192
box 7 3 12 24
use welltap_svt  __well_tap__157
timestamp 1731220323
transform 1 0 3456 0 -1 2152
box 7 3 12 24
use welltap_svt  __well_tap__156
timestamp 1731220323
transform 1 0 1800 0 -1 2152
box 7 3 12 24
use welltap_svt  __well_tap__155
timestamp 1731220323
transform 1 0 3456 0 1 2056
box 7 3 12 24
use welltap_svt  __well_tap__154
timestamp 1731220323
transform 1 0 1800 0 1 2056
box 7 3 12 24
use welltap_svt  __well_tap__153
timestamp 1731220323
transform 1 0 3456 0 -1 2012
box 7 3 12 24
use welltap_svt  __well_tap__152
timestamp 1731220323
transform 1 0 1800 0 -1 2012
box 7 3 12 24
use welltap_svt  __well_tap__151
timestamp 1731220323
transform 1 0 3456 0 1 1920
box 7 3 12 24
use welltap_svt  __well_tap__150
timestamp 1731220323
transform 1 0 1800 0 1 1920
box 7 3 12 24
use welltap_svt  __well_tap__149
timestamp 1731220323
transform 1 0 3456 0 -1 1876
box 7 3 12 24
use welltap_svt  __well_tap__148
timestamp 1731220323
transform 1 0 1800 0 -1 1876
box 7 3 12 24
use welltap_svt  __well_tap__147
timestamp 1731220323
transform 1 0 3456 0 1 1780
box 7 3 12 24
use welltap_svt  __well_tap__146
timestamp 1731220323
transform 1 0 1800 0 1 1780
box 7 3 12 24
use welltap_svt  __well_tap__145
timestamp 1731220323
transform 1 0 3456 0 -1 1728
box 7 3 12 24
use welltap_svt  __well_tap__144
timestamp 1731220323
transform 1 0 1800 0 -1 1728
box 7 3 12 24
use welltap_svt  __well_tap__143
timestamp 1731220323
transform 1 0 3456 0 1 1636
box 7 3 12 24
use welltap_svt  __well_tap__142
timestamp 1731220323
transform 1 0 1800 0 1 1636
box 7 3 12 24
use welltap_svt  __well_tap__141
timestamp 1731220323
transform 1 0 3456 0 -1 1592
box 7 3 12 24
use welltap_svt  __well_tap__140
timestamp 1731220323
transform 1 0 1800 0 -1 1592
box 7 3 12 24
use welltap_svt  __well_tap__139
timestamp 1731220323
transform 1 0 3456 0 1 1504
box 7 3 12 24
use welltap_svt  __well_tap__138
timestamp 1731220323
transform 1 0 1800 0 1 1504
box 7 3 12 24
use welltap_svt  __well_tap__137
timestamp 1731220323
transform 1 0 3456 0 -1 1456
box 7 3 12 24
use welltap_svt  __well_tap__136
timestamp 1731220323
transform 1 0 1800 0 -1 1456
box 7 3 12 24
use welltap_svt  __well_tap__135
timestamp 1731220323
transform 1 0 3456 0 1 1364
box 7 3 12 24
use welltap_svt  __well_tap__134
timestamp 1731220323
transform 1 0 1800 0 1 1364
box 7 3 12 24
use welltap_svt  __well_tap__133
timestamp 1731220323
transform 1 0 3456 0 -1 1316
box 7 3 12 24
use welltap_svt  __well_tap__132
timestamp 1731220323
transform 1 0 1800 0 -1 1316
box 7 3 12 24
use welltap_svt  __well_tap__131
timestamp 1731220323
transform 1 0 3456 0 1 1228
box 7 3 12 24
use welltap_svt  __well_tap__130
timestamp 1731220323
transform 1 0 1800 0 1 1228
box 7 3 12 24
use welltap_svt  __well_tap__129
timestamp 1731220323
transform 1 0 3456 0 -1 1180
box 7 3 12 24
use welltap_svt  __well_tap__128
timestamp 1731220323
transform 1 0 1800 0 -1 1180
box 7 3 12 24
use welltap_svt  __well_tap__127
timestamp 1731220323
transform 1 0 3456 0 1 1084
box 7 3 12 24
use welltap_svt  __well_tap__126
timestamp 1731220323
transform 1 0 1800 0 1 1084
box 7 3 12 24
use welltap_svt  __well_tap__125
timestamp 1731220323
transform 1 0 3456 0 -1 1040
box 7 3 12 24
use welltap_svt  __well_tap__124
timestamp 1731220323
transform 1 0 1800 0 -1 1040
box 7 3 12 24
use welltap_svt  __well_tap__123
timestamp 1731220323
transform 1 0 3456 0 1 948
box 7 3 12 24
use welltap_svt  __well_tap__122
timestamp 1731220323
transform 1 0 1800 0 1 948
box 7 3 12 24
use welltap_svt  __well_tap__121
timestamp 1731220323
transform 1 0 3456 0 -1 908
box 7 3 12 24
use welltap_svt  __well_tap__120
timestamp 1731220323
transform 1 0 1800 0 -1 908
box 7 3 12 24
use welltap_svt  __well_tap__119
timestamp 1731220323
transform 1 0 3456 0 1 812
box 7 3 12 24
use welltap_svt  __well_tap__118
timestamp 1731220323
transform 1 0 1800 0 1 812
box 7 3 12 24
use welltap_svt  __well_tap__117
timestamp 1731220323
transform 1 0 3456 0 -1 768
box 7 3 12 24
use welltap_svt  __well_tap__116
timestamp 1731220323
transform 1 0 1800 0 -1 768
box 7 3 12 24
use welltap_svt  __well_tap__115
timestamp 1731220323
transform 1 0 3456 0 1 680
box 7 3 12 24
use welltap_svt  __well_tap__114
timestamp 1731220323
transform 1 0 1800 0 1 680
box 7 3 12 24
use welltap_svt  __well_tap__113
timestamp 1731220323
transform 1 0 3456 0 -1 632
box 7 3 12 24
use welltap_svt  __well_tap__112
timestamp 1731220323
transform 1 0 1800 0 -1 632
box 7 3 12 24
use welltap_svt  __well_tap__111
timestamp 1731220323
transform 1 0 3456 0 1 544
box 7 3 12 24
use welltap_svt  __well_tap__110
timestamp 1731220323
transform 1 0 1800 0 1 544
box 7 3 12 24
use welltap_svt  __well_tap__109
timestamp 1731220323
transform 1 0 3456 0 -1 488
box 7 3 12 24
use welltap_svt  __well_tap__108
timestamp 1731220323
transform 1 0 1800 0 -1 488
box 7 3 12 24
use welltap_svt  __well_tap__107
timestamp 1731220323
transform 1 0 3456 0 1 400
box 7 3 12 24
use welltap_svt  __well_tap__106
timestamp 1731220323
transform 1 0 1800 0 1 400
box 7 3 12 24
use welltap_svt  __well_tap__105
timestamp 1731220323
transform 1 0 3456 0 -1 356
box 7 3 12 24
use welltap_svt  __well_tap__104
timestamp 1731220323
transform 1 0 1800 0 -1 356
box 7 3 12 24
use welltap_svt  __well_tap__103
timestamp 1731220323
transform 1 0 3456 0 1 268
box 7 3 12 24
use welltap_svt  __well_tap__102
timestamp 1731220323
transform 1 0 1800 0 1 268
box 7 3 12 24
use welltap_svt  __well_tap__101
timestamp 1731220323
transform 1 0 3456 0 -1 220
box 7 3 12 24
use welltap_svt  __well_tap__100
timestamp 1731220323
transform 1 0 1800 0 -1 220
box 7 3 12 24
use welltap_svt  __well_tap__99
timestamp 1731220323
transform 1 0 3456 0 1 108
box 7 3 12 24
use welltap_svt  __well_tap__98
timestamp 1731220323
transform 1 0 1800 0 1 108
box 7 3 12 24
use welltap_svt  __well_tap__97
timestamp 1731220323
transform 1 0 1760 0 1 3460
box 7 3 12 24
use welltap_svt  __well_tap__96
timestamp 1731220323
transform 1 0 104 0 1 3460
box 7 3 12 24
use welltap_svt  __well_tap__95
timestamp 1731220323
transform 1 0 1760 0 -1 3416
box 7 3 12 24
use welltap_svt  __well_tap__94
timestamp 1731220323
transform 1 0 104 0 -1 3416
box 7 3 12 24
use welltap_svt  __well_tap__93
timestamp 1731220323
transform 1 0 1760 0 1 3320
box 7 3 12 24
use welltap_svt  __well_tap__92
timestamp 1731220323
transform 1 0 104 0 1 3320
box 7 3 12 24
use welltap_svt  __well_tap__91
timestamp 1731220323
transform 1 0 1760 0 -1 3272
box 7 3 12 24
use welltap_svt  __well_tap__90
timestamp 1731220323
transform 1 0 104 0 -1 3272
box 7 3 12 24
use welltap_svt  __well_tap__89
timestamp 1731220323
transform 1 0 1760 0 1 3176
box 7 3 12 24
use welltap_svt  __well_tap__88
timestamp 1731220323
transform 1 0 104 0 1 3176
box 7 3 12 24
use welltap_svt  __well_tap__87
timestamp 1731220323
transform 1 0 1760 0 -1 3136
box 7 3 12 24
use welltap_svt  __well_tap__86
timestamp 1731220323
transform 1 0 104 0 -1 3136
box 7 3 12 24
use welltap_svt  __well_tap__85
timestamp 1731220323
transform 1 0 1760 0 1 3044
box 7 3 12 24
use welltap_svt  __well_tap__84
timestamp 1731220323
transform 1 0 104 0 1 3044
box 7 3 12 24
use welltap_svt  __well_tap__83
timestamp 1731220323
transform 1 0 1760 0 -1 2996
box 7 3 12 24
use welltap_svt  __well_tap__82
timestamp 1731220323
transform 1 0 104 0 -1 2996
box 7 3 12 24
use welltap_svt  __well_tap__81
timestamp 1731220323
transform 1 0 1760 0 1 2896
box 7 3 12 24
use welltap_svt  __well_tap__80
timestamp 1731220323
transform 1 0 104 0 1 2896
box 7 3 12 24
use welltap_svt  __well_tap__79
timestamp 1731220323
transform 1 0 1760 0 -1 2848
box 7 3 12 24
use welltap_svt  __well_tap__78
timestamp 1731220323
transform 1 0 104 0 -1 2848
box 7 3 12 24
use welltap_svt  __well_tap__77
timestamp 1731220323
transform 1 0 1760 0 1 2748
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220323
transform 1 0 104 0 1 2748
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220323
transform 1 0 1760 0 -1 2700
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220323
transform 1 0 104 0 -1 2700
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220323
transform 1 0 1760 0 1 2604
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220323
transform 1 0 104 0 1 2604
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220323
transform 1 0 1760 0 -1 2556
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220323
transform 1 0 104 0 -1 2556
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220323
transform 1 0 1760 0 1 2460
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220323
transform 1 0 104 0 1 2460
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220323
transform 1 0 1760 0 -1 2420
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220323
transform 1 0 104 0 -1 2420
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220323
transform 1 0 1760 0 1 2328
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220323
transform 1 0 104 0 1 2328
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220323
transform 1 0 1760 0 -1 2280
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220323
transform 1 0 104 0 -1 2280
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220323
transform 1 0 1760 0 1 2188
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220323
transform 1 0 104 0 1 2188
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220323
transform 1 0 1760 0 -1 2140
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220323
transform 1 0 104 0 -1 2140
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220323
transform 1 0 1760 0 1 2048
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220323
transform 1 0 104 0 1 2048
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220323
transform 1 0 1760 0 -1 2000
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220323
transform 1 0 104 0 -1 2000
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220323
transform 1 0 1760 0 1 1908
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220323
transform 1 0 104 0 1 1908
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220323
transform 1 0 1760 0 -1 1868
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220323
transform 1 0 104 0 -1 1868
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220323
transform 1 0 1760 0 1 1776
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220323
transform 1 0 104 0 1 1776
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220323
transform 1 0 1760 0 -1 1732
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220323
transform 1 0 104 0 -1 1732
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220323
transform 1 0 1760 0 1 1640
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220323
transform 1 0 104 0 1 1640
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220323
transform 1 0 1760 0 -1 1596
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220323
transform 1 0 104 0 -1 1596
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220323
transform 1 0 1760 0 1 1500
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220323
transform 1 0 104 0 1 1500
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220323
transform 1 0 1760 0 -1 1456
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220323
transform 1 0 104 0 -1 1456
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220323
transform 1 0 1760 0 1 1364
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220323
transform 1 0 104 0 1 1364
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220323
transform 1 0 1760 0 -1 1320
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220323
transform 1 0 104 0 -1 1320
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220323
transform 1 0 1760 0 1 1228
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220323
transform 1 0 104 0 1 1228
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220323
transform 1 0 1760 0 -1 1180
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220323
transform 1 0 104 0 -1 1180
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220323
transform 1 0 1760 0 1 1088
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220323
transform 1 0 104 0 1 1088
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220323
transform 1 0 1760 0 -1 1044
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220323
transform 1 0 104 0 -1 1044
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220323
transform 1 0 1760 0 1 948
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220323
transform 1 0 104 0 1 948
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220323
transform 1 0 1760 0 -1 904
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220323
transform 1 0 104 0 -1 904
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220323
transform 1 0 1760 0 1 812
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220323
transform 1 0 104 0 1 812
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220323
transform 1 0 1760 0 -1 768
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220323
transform 1 0 104 0 -1 768
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220323
transform 1 0 1760 0 1 676
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220323
transform 1 0 104 0 1 676
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220323
transform 1 0 1760 0 -1 632
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220323
transform 1 0 104 0 -1 632
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220323
transform 1 0 1760 0 1 536
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220323
transform 1 0 104 0 1 536
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220323
transform 1 0 1760 0 -1 496
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220323
transform 1 0 104 0 -1 496
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220323
transform 1 0 1760 0 1 400
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220323
transform 1 0 104 0 1 400
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220323
transform 1 0 1760 0 -1 356
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220323
transform 1 0 104 0 -1 356
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220323
transform 1 0 1760 0 1 264
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220323
transform 1 0 104 0 1 264
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220323
transform 1 0 1760 0 -1 220
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220323
transform 1 0 104 0 -1 220
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220323
transform 1 0 1760 0 1 104
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220323
transform 1 0 104 0 1 104
box 7 3 12 24
use _0_0cell_0_0gcelem2x0  tst_5999_6
timestamp 1731220323
transform 1 0 3272 0 1 88
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5998_6
timestamp 1731220323
transform 1 0 3360 0 1 88
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5997_6
timestamp 1731220323
transform 1 0 3360 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5996_6
timestamp 1731220323
transform 1 0 3360 0 1 248
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5995_6
timestamp 1731220323
transform 1 0 3352 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5994_6
timestamp 1731220323
transform 1 0 3328 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5993_6
timestamp 1731220323
transform 1 0 3256 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5992_6
timestamp 1731220323
transform 1 0 3128 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5991_6
timestamp 1731220323
transform 1 0 3184 0 1 88
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5990_6
timestamp 1731220323
transform 1 0 3096 0 1 88
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5989_6
timestamp 1731220323
transform 1 0 3000 0 1 88
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5988_6
timestamp 1731220323
transform 1 0 2904 0 1 88
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5987_6
timestamp 1731220323
transform 1 0 2808 0 1 88
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5986_6
timestamp 1731220323
transform 1 0 2712 0 1 88
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5985_6
timestamp 1731220323
transform 1 0 2608 0 1 88
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5984_6
timestamp 1731220323
transform 1 0 2504 0 1 88
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5983_6
timestamp 1731220323
transform 1 0 2760 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5982_6
timestamp 1731220323
transform 1 0 2888 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5981_6
timestamp 1731220323
transform 1 0 3008 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5980_6
timestamp 1731220323
transform 1 0 3216 0 1 248
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5979_6
timestamp 1731220323
transform 1 0 3064 0 1 248
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5978_6
timestamp 1731220323
transform 1 0 2920 0 1 248
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5977_6
timestamp 1731220323
transform 1 0 2792 0 1 248
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5976_6
timestamp 1731220323
transform 1 0 2672 0 1 248
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5975_6
timestamp 1731220323
transform 1 0 3144 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5974_6
timestamp 1731220323
transform 1 0 2944 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5973_6
timestamp 1731220323
transform 1 0 2752 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5972_6
timestamp 1731220323
transform 1 0 2576 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5971_6
timestamp 1731220323
transform 1 0 3096 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5970_6
timestamp 1731220323
transform 1 0 2864 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5969_6
timestamp 1731220323
transform 1 0 2648 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5968_6
timestamp 1731220323
transform 1 0 2448 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5967_6
timestamp 1731220323
transform 1 0 2264 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5966_6
timestamp 1731220323
transform 1 0 2288 0 -1 508
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5965_6
timestamp 1731220323
transform 1 0 2472 0 -1 508
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5964_6
timestamp 1731220323
transform 1 0 2672 0 -1 508
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5963_6
timestamp 1731220323
transform 1 0 3104 0 -1 508
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5962_6
timestamp 1731220323
transform 1 0 2880 0 -1 508
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5961_6
timestamp 1731220323
transform 1 0 2792 0 1 524
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5960_6
timestamp 1731220323
transform 1 0 2616 0 1 524
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5959_6
timestamp 1731220323
transform 1 0 2448 0 1 524
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5958_6
timestamp 1731220323
transform 1 0 2976 0 1 524
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5957_6
timestamp 1731220323
transform 1 0 3160 0 1 524
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5956_6
timestamp 1731220323
transform 1 0 3096 0 -1 652
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5955_6
timestamp 1731220323
transform 1 0 2952 0 -1 652
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5954_6
timestamp 1731220323
transform 1 0 2808 0 -1 652
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5953_6
timestamp 1731220323
transform 1 0 2648 0 -1 652
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5952_6
timestamp 1731220323
transform 1 0 2696 0 1 660
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5951_6
timestamp 1731220323
transform 1 0 2840 0 1 660
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5950_6
timestamp 1731220323
transform 1 0 2976 0 1 660
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5949_6
timestamp 1731220323
transform 1 0 3208 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5948_6
timestamp 1731220323
transform 1 0 3032 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5947_6
timestamp 1731220323
transform 1 0 2864 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5946_6
timestamp 1731220323
transform 1 0 2704 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5945_6
timestamp 1731220323
transform 1 0 3056 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5944_6
timestamp 1731220323
transform 1 0 2904 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5943_6
timestamp 1731220323
transform 1 0 2760 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5942_6
timestamp 1731220323
transform 1 0 2632 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5941_6
timestamp 1731220323
transform 1 0 2824 0 -1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5940_6
timestamp 1731220323
transform 1 0 2736 0 -1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5939_6
timestamp 1731220323
transform 1 0 2648 0 -1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5938_6
timestamp 1731220323
transform 1 0 2560 0 -1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5937_6
timestamp 1731220323
transform 1 0 2384 0 -1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5936_6
timestamp 1731220323
transform 1 0 2296 0 -1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5935_6
timestamp 1731220323
transform 1 0 2208 0 -1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5934_6
timestamp 1731220323
transform 1 0 2120 0 -1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5933_6
timestamp 1731220323
transform 1 0 2128 0 1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5932_6
timestamp 1731220323
transform 1 0 2456 0 1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5931_6
timestamp 1731220323
transform 1 0 2624 0 1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5930_6
timestamp 1731220323
transform 1 0 2984 0 1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5929_6
timestamp 1731220323
transform 1 0 2800 0 1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5928_6
timestamp 1731220323
transform 1 0 2696 0 -1 1060
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5927_6
timestamp 1731220323
transform 1 0 2536 0 -1 1060
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5926_6
timestamp 1731220323
transform 1 0 3024 0 -1 1060
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5925_6
timestamp 1731220323
transform 1 0 2856 0 -1 1060
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5924_6
timestamp 1731220323
transform 1 0 2744 0 1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5923_6
timestamp 1731220323
transform 1 0 2592 0 1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5922_6
timestamp 1731220323
transform 1 0 2896 0 1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5921_6
timestamp 1731220323
transform 1 0 3056 0 1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5920_6
timestamp 1731220323
transform 1 0 2968 0 -1 1200
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5919_6
timestamp 1731220323
transform 1 0 2832 0 -1 1200
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5918_6
timestamp 1731220323
transform 1 0 2696 0 -1 1200
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5917_6
timestamp 1731220323
transform 1 0 2592 0 1 1208
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5916_6
timestamp 1731220323
transform 1 0 2352 0 1 1208
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5915_6
timestamp 1731220323
transform 1 0 2800 0 1 1208
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5914_6
timestamp 1731220323
transform 1 0 2680 0 -1 1336
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5913_6
timestamp 1731220323
transform 1 0 2856 0 -1 1336
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5912_6
timestamp 1731220323
transform 1 0 3032 0 -1 1336
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5911_6
timestamp 1731220323
transform 1 0 3208 0 -1 1336
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5910_6
timestamp 1731220323
transform 1 0 3192 0 1 1208
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5909_6
timestamp 1731220323
transform 1 0 3000 0 1 1208
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5908_6
timestamp 1731220323
transform 1 0 3104 0 -1 1200
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5907_6
timestamp 1731220323
transform 1 0 3240 0 -1 1200
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5906_6
timestamp 1731220323
transform 1 0 3216 0 1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5905_6
timestamp 1731220323
transform 1 0 3200 0 -1 1060
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5904_6
timestamp 1731220323
transform 1 0 3176 0 1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5903_6
timestamp 1731220323
transform 1 0 3216 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5902_6
timestamp 1731220323
transform 1 0 3112 0 1 660
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5901_6
timestamp 1731220323
transform 1 0 3248 0 1 660
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5900_6
timestamp 1731220323
transform 1 0 3240 0 -1 652
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5899_6
timestamp 1731220323
transform 1 0 3328 0 -1 508
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5898_6
timestamp 1731220323
transform 1 0 3352 0 1 524
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5897_6
timestamp 1731220323
transform 1 0 3360 0 -1 652
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5896_6
timestamp 1731220323
transform 1 0 3360 0 1 660
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5895_6
timestamp 1731220323
transform 1 0 3360 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5894_6
timestamp 1731220323
transform 1 0 3360 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5893_6
timestamp 1731220323
transform 1 0 3360 0 1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5892_6
timestamp 1731220323
transform 1 0 3360 0 -1 1060
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5891_6
timestamp 1731220323
transform 1 0 3360 0 1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5890_6
timestamp 1731220323
transform 1 0 3360 0 -1 1200
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5889_6
timestamp 1731220323
transform 1 0 3360 0 1 1208
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5888_6
timestamp 1731220323
transform 1 0 3360 0 -1 1336
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5887_6
timestamp 1731220323
transform 1 0 3360 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5886_6
timestamp 1731220323
transform 1 0 3360 0 -1 1476
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5885_6
timestamp 1731220323
transform 1 0 3256 0 -1 1476
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5884_6
timestamp 1731220323
transform 1 0 3248 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5883_6
timestamp 1731220323
transform 1 0 3120 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5882_6
timestamp 1731220323
transform 1 0 2992 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5881_6
timestamp 1731220323
transform 1 0 2856 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5880_6
timestamp 1731220323
transform 1 0 2712 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5879_6
timestamp 1731220323
transform 1 0 2552 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5878_6
timestamp 1731220323
transform 1 0 3128 0 -1 1476
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5877_6
timestamp 1731220323
transform 1 0 3000 0 -1 1476
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5876_6
timestamp 1731220323
transform 1 0 2864 0 -1 1476
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5875_6
timestamp 1731220323
transform 1 0 2728 0 -1 1476
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5874_6
timestamp 1731220323
transform 1 0 2584 0 -1 1476
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5873_6
timestamp 1731220323
transform 1 0 3048 0 1 1484
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5872_6
timestamp 1731220323
transform 1 0 2920 0 1 1484
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5871_6
timestamp 1731220323
transform 1 0 2792 0 1 1484
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5870_6
timestamp 1731220323
transform 1 0 2672 0 1 1484
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5869_6
timestamp 1731220323
transform 1 0 2544 0 1 1484
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5868_6
timestamp 1731220323
transform 1 0 2880 0 -1 1612
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5867_6
timestamp 1731220323
transform 1 0 2768 0 -1 1612
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5866_6
timestamp 1731220323
transform 1 0 2664 0 -1 1612
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5865_6
timestamp 1731220323
transform 1 0 2560 0 -1 1612
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5864_6
timestamp 1731220323
transform 1 0 2888 0 1 1616
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5863_6
timestamp 1731220323
transform 1 0 2800 0 1 1616
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5862_6
timestamp 1731220323
transform 1 0 2712 0 1 1616
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5861_6
timestamp 1731220323
transform 1 0 2624 0 1 1616
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5860_6
timestamp 1731220323
transform 1 0 2536 0 1 1616
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5859_6
timestamp 1731220323
transform 1 0 2576 0 -1 1748
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5858_6
timestamp 1731220323
transform 1 0 2840 0 -1 1748
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5857_6
timestamp 1731220323
transform 1 0 2752 0 -1 1748
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5856_6
timestamp 1731220323
transform 1 0 2664 0 -1 1748
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5855_6
timestamp 1731220323
transform 1 0 2624 0 1 1760
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5854_6
timestamp 1731220323
transform 1 0 2536 0 1 1760
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5853_6
timestamp 1731220323
transform 1 0 2712 0 1 1760
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5852_6
timestamp 1731220323
transform 1 0 2800 0 1 1760
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5851_6
timestamp 1731220323
transform 1 0 2888 0 1 1760
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5850_6
timestamp 1731220323
transform 1 0 2976 0 -1 1896
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5849_6
timestamp 1731220323
transform 1 0 2864 0 -1 1896
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5848_6
timestamp 1731220323
transform 1 0 2752 0 -1 1896
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5847_6
timestamp 1731220323
transform 1 0 2640 0 -1 1896
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5846_6
timestamp 1731220323
transform 1 0 2536 0 -1 1896
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5845_6
timestamp 1731220323
transform 1 0 2568 0 1 1900
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5844_6
timestamp 1731220323
transform 1 0 2704 0 1 1900
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5843_6
timestamp 1731220323
transform 1 0 2824 0 1 1900
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5842_6
timestamp 1731220323
transform 1 0 2944 0 1 1900
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5841_6
timestamp 1731220323
transform 1 0 3000 0 -1 2032
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5840_6
timestamp 1731220323
transform 1 0 2816 0 -1 2032
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5839_6
timestamp 1731220323
transform 1 0 2624 0 -1 2032
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5838_6
timestamp 1731220323
transform 1 0 2496 0 1 2036
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5837_6
timestamp 1731220323
transform 1 0 2648 0 1 2036
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5836_6
timestamp 1731220323
transform 1 0 2784 0 1 2036
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5835_6
timestamp 1731220323
transform 1 0 2912 0 1 2036
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5834_6
timestamp 1731220323
transform 1 0 3184 0 -1 2172
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5833_6
timestamp 1731220323
transform 1 0 3264 0 1 2036
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5832_6
timestamp 1731220323
transform 1 0 3152 0 1 2036
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5831_6
timestamp 1731220323
transform 1 0 3032 0 1 2036
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5830_6
timestamp 1731220323
transform 1 0 3192 0 -1 2032
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5829_6
timestamp 1731220323
transform 1 0 3160 0 1 1900
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5828_6
timestamp 1731220323
transform 1 0 3056 0 1 1900
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5827_6
timestamp 1731220323
transform 1 0 3272 0 1 1900
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5826_6
timestamp 1731220323
transform 1 0 3360 0 1 1900
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5825_6
timestamp 1731220323
transform 1 0 3360 0 -1 2032
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5824_6
timestamp 1731220323
transform 1 0 3360 0 1 2036
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5823_6
timestamp 1731220323
transform 1 0 3272 0 -1 2172
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5822_6
timestamp 1731220323
transform 1 0 3360 0 -1 2172
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5821_6
timestamp 1731220323
transform 1 0 3360 0 1 2172
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5820_6
timestamp 1731220323
transform 1 0 3360 0 -1 2300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5819_6
timestamp 1731220323
transform 1 0 3216 0 -1 2300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5818_6
timestamp 1731220323
transform 1 0 3048 0 -1 2300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5817_6
timestamp 1731220323
transform 1 0 2952 0 1 2172
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5816_6
timestamp 1731220323
transform 1 0 3096 0 1 2172
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5815_6
timestamp 1731220323
transform 1 0 3240 0 1 2172
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5814_6
timestamp 1731220323
transform 1 0 3096 0 -1 2172
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5813_6
timestamp 1731220323
transform 1 0 3008 0 -1 2172
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5812_6
timestamp 1731220323
transform 1 0 2920 0 -1 2172
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5811_6
timestamp 1731220323
transform 1 0 2808 0 1 2172
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5810_6
timestamp 1731220323
transform 1 0 2648 0 1 2172
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5809_6
timestamp 1731220323
transform 1 0 2712 0 -1 2300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5808_6
timestamp 1731220323
transform 1 0 2880 0 -1 2300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5807_6
timestamp 1731220323
transform 1 0 3016 0 1 2308
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5806_6
timestamp 1731220323
transform 1 0 2904 0 1 2308
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5805_6
timestamp 1731220323
transform 1 0 2792 0 1 2308
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5804_6
timestamp 1731220323
transform 1 0 2680 0 1 2308
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5803_6
timestamp 1731220323
transform 1 0 2928 0 -1 2436
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5802_6
timestamp 1731220323
transform 1 0 2832 0 -1 2436
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5801_6
timestamp 1731220323
transform 1 0 2736 0 -1 2436
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5800_6
timestamp 1731220323
transform 1 0 2648 0 -1 2436
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5799_6
timestamp 1731220323
transform 1 0 2560 0 -1 2436
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5798_6
timestamp 1731220323
transform 1 0 3136 0 1 2444
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5797_6
timestamp 1731220323
transform 1 0 2912 0 1 2444
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5796_6
timestamp 1731220323
transform 1 0 2704 0 1 2444
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5795_6
timestamp 1731220323
transform 1 0 2520 0 1 2444
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5794_6
timestamp 1731220323
transform 1 0 2992 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5793_6
timestamp 1731220323
transform 1 0 2808 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5792_6
timestamp 1731220323
transform 1 0 2640 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5791_6
timestamp 1731220323
transform 1 0 2480 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5790_6
timestamp 1731220323
transform 1 0 2336 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5789_6
timestamp 1731220323
transform 1 0 2424 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5788_6
timestamp 1731220323
transform 1 0 2576 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5787_6
timestamp 1731220323
transform 1 0 3160 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5786_6
timestamp 1731220323
transform 1 0 2952 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5785_6
timestamp 1731220323
transform 1 0 2752 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5784_6
timestamp 1731220323
transform 1 0 2680 0 -1 2724
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5783_6
timestamp 1731220323
transform 1 0 2536 0 -1 2724
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5782_6
timestamp 1731220323
transform 1 0 2840 0 -1 2724
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5781_6
timestamp 1731220323
transform 1 0 3200 0 -1 2724
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5780_6
timestamp 1731220323
transform 1 0 3016 0 -1 2724
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5779_6
timestamp 1731220323
transform 1 0 2904 0 1 2740
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5778_6
timestamp 1731220323
transform 1 0 2744 0 1 2740
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5777_6
timestamp 1731220323
transform 1 0 2576 0 1 2740
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5776_6
timestamp 1731220323
transform 1 0 3064 0 1 2740
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5775_6
timestamp 1731220323
transform 1 0 3056 0 -1 2872
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5774_6
timestamp 1731220323
transform 1 0 2896 0 -1 2872
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5773_6
timestamp 1731220323
transform 1 0 2728 0 -1 2872
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5772_6
timestamp 1731220323
transform 1 0 2752 0 1 2872
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5771_6
timestamp 1731220323
transform 1 0 2904 0 1 2872
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5770_6
timestamp 1731220323
transform 1 0 3056 0 1 2872
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5769_6
timestamp 1731220323
transform 1 0 3200 0 1 2872
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5768_6
timestamp 1731220323
transform 1 0 3352 0 1 2872
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5767_6
timestamp 1731220323
transform 1 0 3216 0 -1 2872
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5766_6
timestamp 1731220323
transform 1 0 3224 0 1 2740
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5765_6
timestamp 1731220323
transform 1 0 3184 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5764_6
timestamp 1731220323
transform 1 0 3360 0 1 2444
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5763_6
timestamp 1731220323
transform 1 0 3360 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5762_6
timestamp 1731220323
transform 1 0 3360 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5761_6
timestamp 1731220323
transform 1 0 3360 0 -1 2724
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5760_6
timestamp 1731220323
transform 1 0 3360 0 1 2740
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5759_6
timestamp 1731220323
transform 1 0 3360 0 -1 2872
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5758_6
timestamp 1731220323
transform 1 0 3360 0 -1 3012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5757_6
timestamp 1731220323
transform 1 0 3360 0 1 3028
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5756_6
timestamp 1731220323
transform 1 0 3360 0 -1 3164
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5755_6
timestamp 1731220323
transform 1 0 3328 0 1 3164
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5754_6
timestamp 1731220323
transform 1 0 3224 0 -1 3164
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5753_6
timestamp 1731220323
transform 1 0 3072 0 -1 3164
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5752_6
timestamp 1731220323
transform 1 0 2912 0 -1 3164
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5751_6
timestamp 1731220323
transform 1 0 3000 0 1 3164
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5750_6
timestamp 1731220323
transform 1 0 3160 0 1 3164
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5749_6
timestamp 1731220323
transform 1 0 3192 0 -1 3296
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5748_6
timestamp 1731220323
transform 1 0 3032 0 -1 3296
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5747_6
timestamp 1731220323
transform 1 0 2872 0 -1 3296
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5746_6
timestamp 1731220323
transform 1 0 2832 0 1 3296
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5745_6
timestamp 1731220323
transform 1 0 2968 0 1 3296
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5744_6
timestamp 1731220323
transform 1 0 3112 0 1 3296
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5743_6
timestamp 1731220323
transform 1 0 3144 0 -1 3428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5742_6
timestamp 1731220323
transform 1 0 3032 0 -1 3428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5741_6
timestamp 1731220323
transform 1 0 2928 0 -1 3428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5740_6
timestamp 1731220323
transform 1 0 2824 0 -1 3428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5739_6
timestamp 1731220323
transform 1 0 2960 0 1 3428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5738_6
timestamp 1731220323
transform 1 0 2792 0 1 3428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5737_6
timestamp 1731220323
transform 1 0 2632 0 1 3428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5736_6
timestamp 1731220323
transform 1 0 2472 0 1 3428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5735_6
timestamp 1731220323
transform 1 0 2504 0 -1 3428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5734_6
timestamp 1731220323
transform 1 0 2616 0 -1 3428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5733_6
timestamp 1731220323
transform 1 0 2720 0 -1 3428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5732_6
timestamp 1731220323
transform 1 0 2696 0 1 3296
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5731_6
timestamp 1731220323
transform 1 0 2712 0 -1 3296
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5730_6
timestamp 1731220323
transform 1 0 2680 0 1 3164
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5729_6
timestamp 1731220323
transform 1 0 2840 0 1 3164
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5728_6
timestamp 1731220323
transform 1 0 2752 0 -1 3164
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5727_6
timestamp 1731220323
transform 1 0 2576 0 -1 3164
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5726_6
timestamp 1731220323
transform 1 0 3144 0 1 3028
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5725_6
timestamp 1731220323
transform 1 0 2912 0 1 3028
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5724_6
timestamp 1731220323
transform 1 0 2688 0 1 3028
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5723_6
timestamp 1731220323
transform 1 0 2480 0 1 3028
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5722_6
timestamp 1731220323
transform 1 0 3176 0 -1 3012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5721_6
timestamp 1731220323
transform 1 0 2976 0 -1 3012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5720_6
timestamp 1731220323
transform 1 0 2784 0 -1 3012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5719_6
timestamp 1731220323
transform 1 0 2616 0 -1 3012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5718_6
timestamp 1731220323
transform 1 0 2472 0 -1 3012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5717_6
timestamp 1731220323
transform 1 0 2352 0 -1 3012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5716_6
timestamp 1731220323
transform 1 0 2240 0 -1 3012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5715_6
timestamp 1731220323
transform 1 0 2136 0 -1 3012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5714_6
timestamp 1731220323
transform 1 0 2208 0 1 2872
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5713_6
timestamp 1731220323
transform 1 0 2400 0 1 2872
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5712_6
timestamp 1731220323
transform 1 0 2584 0 1 2872
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5711_6
timestamp 1731220323
transform 1 0 2560 0 -1 2872
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5710_6
timestamp 1731220323
transform 1 0 2376 0 -1 2872
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5709_6
timestamp 1731220323
transform 1 0 2184 0 -1 2872
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5708_6
timestamp 1731220323
transform 1 0 2008 0 1 2740
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5707_6
timestamp 1731220323
transform 1 0 2208 0 1 2740
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5706_6
timestamp 1731220323
transform 1 0 2400 0 1 2740
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5705_6
timestamp 1731220323
transform 1 0 2400 0 -1 2724
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5704_6
timestamp 1731220323
transform 1 0 2272 0 -1 2724
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5703_6
timestamp 1731220323
transform 1 0 2152 0 -1 2724
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5702_6
timestamp 1731220323
transform 1 0 2032 0 -1 2724
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5701_6
timestamp 1731220323
transform 1 0 2288 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5700_6
timestamp 1731220323
transform 1 0 2176 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5699_6
timestamp 1731220323
transform 1 0 2064 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5698_6
timestamp 1731220323
transform 1 0 1960 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5697_6
timestamp 1731220323
transform 1 0 1864 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5696_6
timestamp 1731220323
transform 1 0 1824 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5695_6
timestamp 1731220323
transform 1 0 1912 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5694_6
timestamp 1731220323
transform 1 0 2000 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5693_6
timestamp 1731220323
transform 1 0 2104 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5692_6
timestamp 1731220323
transform 1 0 2216 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5691_6
timestamp 1731220323
transform 1 0 2128 0 1 2444
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5690_6
timestamp 1731220323
transform 1 0 2032 0 1 2444
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5689_6
timestamp 1731220323
transform 1 0 1944 0 1 2444
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5688_6
timestamp 1731220323
transform 1 0 2232 0 1 2444
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5687_6
timestamp 1731220323
transform 1 0 2360 0 1 2444
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5686_6
timestamp 1731220323
transform 1 0 2296 0 -1 2436
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5685_6
timestamp 1731220323
transform 1 0 2208 0 -1 2436
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5684_6
timestamp 1731220323
transform 1 0 2384 0 -1 2436
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5683_6
timestamp 1731220323
transform 1 0 2472 0 -1 2436
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5682_6
timestamp 1731220323
transform 1 0 2568 0 1 2308
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5681_6
timestamp 1731220323
transform 1 0 2464 0 1 2308
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5680_6
timestamp 1731220323
transform 1 0 2360 0 1 2308
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5679_6
timestamp 1731220323
transform 1 0 2256 0 1 2308
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5678_6
timestamp 1731220323
transform 1 0 2160 0 1 2308
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5677_6
timestamp 1731220323
transform 1 0 2544 0 -1 2300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5676_6
timestamp 1731220323
transform 1 0 2368 0 -1 2300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5675_6
timestamp 1731220323
transform 1 0 2192 0 -1 2300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5674_6
timestamp 1731220323
transform 1 0 2032 0 -1 2300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5673_6
timestamp 1731220323
transform 1 0 1880 0 -1 2300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5672_6
timestamp 1731220323
transform 1 0 2480 0 1 2172
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5671_6
timestamp 1731220323
transform 1 0 2304 0 1 2172
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5670_6
timestamp 1731220323
transform 1 0 2128 0 1 2172
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5669_6
timestamp 1731220323
transform 1 0 1960 0 1 2172
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5668_6
timestamp 1731220323
transform 1 0 1824 0 1 2172
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5667_6
timestamp 1731220323
transform 1 0 1664 0 1 2168
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5666_6
timestamp 1731220323
transform 1 0 1496 0 1 2168
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5665_6
timestamp 1731220323
transform 1 0 1312 0 1 2168
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5664_6
timestamp 1731220323
transform 1 0 1224 0 -1 2160
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5663_6
timestamp 1731220323
transform 1 0 1096 0 -1 2160
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5662_6
timestamp 1731220323
transform 1 0 1344 0 -1 2160
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5661_6
timestamp 1731220323
transform 1 0 1456 0 -1 2160
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5660_6
timestamp 1731220323
transform 1 0 1568 0 -1 2160
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5659_6
timestamp 1731220323
transform 1 0 1664 0 -1 2160
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5658_6
timestamp 1731220323
transform 1 0 1824 0 1 2036
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5657_6
timestamp 1731220323
transform 1 0 1984 0 1 2036
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5656_6
timestamp 1731220323
transform 1 0 2160 0 1 2036
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5655_6
timestamp 1731220323
transform 1 0 2336 0 1 2036
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5654_6
timestamp 1731220323
transform 1 0 2424 0 -1 2032
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5653_6
timestamp 1731220323
transform 1 0 2216 0 -1 2032
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5652_6
timestamp 1731220323
transform 1 0 2008 0 -1 2032
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5651_6
timestamp 1731220323
transform 1 0 1824 0 -1 2032
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5650_6
timestamp 1731220323
transform 1 0 1856 0 1 1900
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5649_6
timestamp 1731220323
transform 1 0 1992 0 1 1900
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5648_6
timestamp 1731220323
transform 1 0 2136 0 1 1900
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5647_6
timestamp 1731220323
transform 1 0 2424 0 1 1900
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5646_6
timestamp 1731220323
transform 1 0 2280 0 1 1900
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5645_6
timestamp 1731220323
transform 1 0 2208 0 -1 1896
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5644_6
timestamp 1731220323
transform 1 0 2104 0 -1 1896
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5643_6
timestamp 1731220323
transform 1 0 2008 0 -1 1896
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5642_6
timestamp 1731220323
transform 1 0 2320 0 -1 1896
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5641_6
timestamp 1731220323
transform 1 0 2432 0 -1 1896
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5640_6
timestamp 1731220323
transform 1 0 2448 0 1 1760
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5639_6
timestamp 1731220323
transform 1 0 2360 0 1 1760
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5638_6
timestamp 1731220323
transform 1 0 2272 0 1 1760
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5637_6
timestamp 1731220323
transform 1 0 2184 0 1 1760
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5636_6
timestamp 1731220323
transform 1 0 2096 0 1 1760
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5635_6
timestamp 1731220323
transform 1 0 2136 0 -1 1748
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5634_6
timestamp 1731220323
transform 1 0 2224 0 -1 1748
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5633_6
timestamp 1731220323
transform 1 0 2312 0 -1 1748
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5632_6
timestamp 1731220323
transform 1 0 2400 0 -1 1748
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5631_6
timestamp 1731220323
transform 1 0 2488 0 -1 1748
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5630_6
timestamp 1731220323
transform 1 0 2448 0 1 1616
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5629_6
timestamp 1731220323
transform 1 0 2360 0 1 1616
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5628_6
timestamp 1731220323
transform 1 0 2272 0 1 1616
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5627_6
timestamp 1731220323
transform 1 0 2184 0 1 1616
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5626_6
timestamp 1731220323
transform 1 0 2096 0 1 1616
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5625_6
timestamp 1731220323
transform 1 0 2456 0 -1 1612
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5624_6
timestamp 1731220323
transform 1 0 2352 0 -1 1612
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5623_6
timestamp 1731220323
transform 1 0 2248 0 -1 1612
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5622_6
timestamp 1731220323
transform 1 0 2152 0 -1 1612
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5621_6
timestamp 1731220323
transform 1 0 2056 0 -1 1612
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5620_6
timestamp 1731220323
transform 1 0 2416 0 1 1484
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5619_6
timestamp 1731220323
transform 1 0 2288 0 1 1484
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5618_6
timestamp 1731220323
transform 1 0 2160 0 1 1484
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5617_6
timestamp 1731220323
transform 1 0 2032 0 1 1484
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5616_6
timestamp 1731220323
transform 1 0 1912 0 1 1484
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5615_6
timestamp 1731220323
transform 1 0 2424 0 -1 1476
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5614_6
timestamp 1731220323
transform 1 0 2264 0 -1 1476
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5613_6
timestamp 1731220323
transform 1 0 2104 0 -1 1476
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5612_6
timestamp 1731220323
transform 1 0 1944 0 -1 1476
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5611_6
timestamp 1731220323
transform 1 0 1824 0 -1 1476
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5610_6
timestamp 1731220323
transform 1 0 2376 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5609_6
timestamp 1731220323
transform 1 0 2192 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5608_6
timestamp 1731220323
transform 1 0 2000 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5607_6
timestamp 1731220323
transform 1 0 1664 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5606_6
timestamp 1731220323
transform 1 0 1824 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5605_6
timestamp 1731220323
transform 1 0 1824 0 -1 1336
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5604_6
timestamp 1731220323
transform 1 0 1960 0 -1 1336
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5603_6
timestamp 1731220323
transform 1 0 2504 0 -1 1336
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5602_6
timestamp 1731220323
transform 1 0 2320 0 -1 1336
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5601_6
timestamp 1731220323
transform 1 0 2136 0 -1 1336
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5600_6
timestamp 1731220323
transform 1 0 2088 0 1 1208
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5599_6
timestamp 1731220323
transform 1 0 1824 0 1 1208
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5598_6
timestamp 1731220323
transform 1 0 1664 0 1 1208
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5597_6
timestamp 1731220323
transform 1 0 1496 0 1 1208
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5596_6
timestamp 1731220323
transform 1 0 1664 0 -1 1340
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5595_6
timestamp 1731220323
transform 1 0 1528 0 -1 1340
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5594_6
timestamp 1731220323
transform 1 0 1368 0 -1 1340
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5593_6
timestamp 1731220323
transform 1 0 1216 0 -1 1340
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5592_6
timestamp 1731220323
transform 1 0 1552 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5591_6
timestamp 1731220323
transform 1 0 1424 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5590_6
timestamp 1731220323
transform 1 0 1296 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5589_6
timestamp 1731220323
transform 1 0 1160 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5588_6
timestamp 1731220323
transform 1 0 1008 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5587_6
timestamp 1731220323
transform 1 0 1584 0 -1 1476
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5586_6
timestamp 1731220323
transform 1 0 1424 0 -1 1476
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5585_6
timestamp 1731220323
transform 1 0 1272 0 -1 1476
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5584_6
timestamp 1731220323
transform 1 0 1120 0 -1 1476
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5583_6
timestamp 1731220323
transform 1 0 952 0 -1 1476
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5582_6
timestamp 1731220323
transform 1 0 1440 0 1 1480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5581_6
timestamp 1731220323
transform 1 0 1304 0 1 1480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5580_6
timestamp 1731220323
transform 1 0 1168 0 1 1480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5579_6
timestamp 1731220323
transform 1 0 1040 0 1 1480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5578_6
timestamp 1731220323
transform 1 0 904 0 1 1480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5577_6
timestamp 1731220323
transform 1 0 1272 0 -1 1616
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5576_6
timestamp 1731220323
transform 1 0 1160 0 -1 1616
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5575_6
timestamp 1731220323
transform 1 0 1048 0 -1 1616
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5574_6
timestamp 1731220323
transform 1 0 936 0 -1 1616
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5573_6
timestamp 1731220323
transform 1 0 824 0 -1 1616
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5572_6
timestamp 1731220323
transform 1 0 752 0 1 1620
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5571_6
timestamp 1731220323
transform 1 0 848 0 1 1620
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5570_6
timestamp 1731220323
transform 1 0 944 0 1 1620
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5569_6
timestamp 1731220323
transform 1 0 1136 0 1 1620
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5568_6
timestamp 1731220323
transform 1 0 1040 0 1 1620
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5567_6
timestamp 1731220323
transform 1 0 944 0 -1 1752
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5566_6
timestamp 1731220323
transform 1 0 1048 0 -1 1752
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5565_6
timestamp 1731220323
transform 1 0 1152 0 -1 1752
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5564_6
timestamp 1731220323
transform 1 0 1264 0 -1 1752
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5563_6
timestamp 1731220323
transform 1 0 1376 0 -1 1752
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5562_6
timestamp 1731220323
transform 1 0 1272 0 1 1756
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5561_6
timestamp 1731220323
transform 1 0 1144 0 1 1756
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5560_6
timestamp 1731220323
transform 1 0 1400 0 1 1756
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5559_6
timestamp 1731220323
transform 1 0 1528 0 1 1756
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5558_6
timestamp 1731220323
transform 1 0 1664 0 1 1756
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5557_6
timestamp 1731220323
transform 1 0 1664 0 -1 1888
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5556_6
timestamp 1731220323
transform 1 0 1504 0 -1 1888
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5555_6
timestamp 1731220323
transform 1 0 1344 0 -1 1888
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5554_6
timestamp 1731220323
transform 1 0 1192 0 -1 1888
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5553_6
timestamp 1731220323
transform 1 0 1152 0 1 1888
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5552_6
timestamp 1731220323
transform 1 0 1304 0 1 1888
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5551_6
timestamp 1731220323
transform 1 0 1464 0 1 1888
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5550_6
timestamp 1731220323
transform 1 0 1320 0 -1 2020
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5549_6
timestamp 1731220323
transform 1 0 1176 0 -1 2020
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5548_6
timestamp 1731220323
transform 1 0 1040 0 -1 2020
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5547_6
timestamp 1731220323
transform 1 0 1272 0 1 2028
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5546_6
timestamp 1731220323
transform 1 0 1152 0 1 2028
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5545_6
timestamp 1731220323
transform 1 0 1040 0 1 2028
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5544_6
timestamp 1731220323
transform 1 0 968 0 -1 2160
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5543_6
timestamp 1731220323
transform 1 0 832 0 -1 2160
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5542_6
timestamp 1731220323
transform 1 0 928 0 1 2028
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5541_6
timestamp 1731220323
transform 1 0 816 0 1 2028
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5540_6
timestamp 1731220323
transform 1 0 696 0 1 2028
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5539_6
timestamp 1731220323
transform 1 0 768 0 -1 2020
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5538_6
timestamp 1731220323
transform 1 0 904 0 -1 2020
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5537_6
timestamp 1731220323
transform 1 0 1000 0 1 1888
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5536_6
timestamp 1731220323
transform 1 0 848 0 1 1888
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5535_6
timestamp 1731220323
transform 1 0 880 0 -1 1888
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5534_6
timestamp 1731220323
transform 1 0 1040 0 -1 1888
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5533_6
timestamp 1731220323
transform 1 0 1016 0 1 1756
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5532_6
timestamp 1731220323
transform 1 0 880 0 1 1756
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5531_6
timestamp 1731220323
transform 1 0 752 0 1 1756
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5530_6
timestamp 1731220323
transform 1 0 840 0 -1 1752
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5529_6
timestamp 1731220323
transform 1 0 736 0 -1 1752
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5528_6
timestamp 1731220323
transform 1 0 656 0 1 1620
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5527_6
timestamp 1731220323
transform 1 0 568 0 1 1620
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5526_6
timestamp 1731220323
transform 1 0 600 0 -1 1616
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5525_6
timestamp 1731220323
transform 1 0 712 0 -1 1616
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5524_6
timestamp 1731220323
transform 1 0 616 0 1 1480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5523_6
timestamp 1731220323
transform 1 0 760 0 1 1480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5522_6
timestamp 1731220323
transform 1 0 776 0 -1 1476
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5521_6
timestamp 1731220323
transform 1 0 576 0 -1 1476
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5520_6
timestamp 1731220323
transform 1 0 672 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5519_6
timestamp 1731220323
transform 1 0 848 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5518_6
timestamp 1731220323
transform 1 0 1056 0 -1 1340
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5517_6
timestamp 1731220323
transform 1 0 888 0 -1 1340
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5516_6
timestamp 1731220323
transform 1 0 720 0 -1 1340
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5515_6
timestamp 1731220323
transform 1 0 672 0 1 1208
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5514_6
timestamp 1731220323
transform 1 0 816 0 1 1208
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5513_6
timestamp 1731220323
transform 1 0 968 0 1 1208
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5512_6
timestamp 1731220323
transform 1 0 1136 0 1 1208
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5511_6
timestamp 1731220323
transform 1 0 1312 0 1 1208
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5510_6
timestamp 1731220323
transform 1 0 1240 0 -1 1200
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5509_6
timestamp 1731220323
transform 1 0 1112 0 -1 1200
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5508_6
timestamp 1731220323
transform 1 0 984 0 -1 1200
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5507_6
timestamp 1731220323
transform 1 0 864 0 -1 1200
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5506_6
timestamp 1731220323
transform 1 0 736 0 -1 1200
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5505_6
timestamp 1731220323
transform 1 0 880 0 1 1068
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5504_6
timestamp 1731220323
transform 1 0 1008 0 1 1068
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5503_6
timestamp 1731220323
transform 1 0 1136 0 1 1068
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5502_6
timestamp 1731220323
transform 1 0 1264 0 1 1068
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5501_6
timestamp 1731220323
transform 1 0 1392 0 1 1068
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5500_6
timestamp 1731220323
transform 1 0 1272 0 -1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5499_6
timestamp 1731220323
transform 1 0 1152 0 -1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5498_6
timestamp 1731220323
transform 1 0 1032 0 -1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5497_6
timestamp 1731220323
transform 1 0 1528 0 -1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5496_6
timestamp 1731220323
transform 1 0 1400 0 -1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5495_6
timestamp 1731220323
transform 1 0 1352 0 1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5494_6
timestamp 1731220323
transform 1 0 1248 0 1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5493_6
timestamp 1731220323
transform 1 0 1136 0 1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5492_6
timestamp 1731220323
transform 1 0 1464 0 1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5491_6
timestamp 1731220323
transform 1 0 1552 0 -1 924
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5490_6
timestamp 1731220323
transform 1 0 1576 0 1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5489_6
timestamp 1731220323
transform 1 0 1664 0 1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5488_6
timestamp 1731220323
transform 1 0 1824 0 1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5487_6
timestamp 1731220323
transform 1 0 1968 0 1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5486_6
timestamp 1731220323
transform 1 0 1840 0 -1 1060
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5485_6
timestamp 1731220323
transform 1 0 1976 0 -1 1060
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5484_6
timestamp 1731220323
transform 1 0 2112 0 -1 1060
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5483_6
timestamp 1731220323
transform 1 0 2184 0 1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5482_6
timestamp 1731220323
transform 1 0 2056 0 1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5481_6
timestamp 1731220323
transform 1 0 1936 0 1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5480_6
timestamp 1731220323
transform 1 0 1928 0 -1 1200
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5479_6
timestamp 1731220323
transform 1 0 2032 0 -1 1200
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5478_6
timestamp 1731220323
transform 1 0 2152 0 -1 1200
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5477_6
timestamp 1731220323
transform 1 0 2280 0 -1 1200
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5476_6
timestamp 1731220323
transform 1 0 2416 0 -1 1200
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5475_6
timestamp 1731220323
transform 1 0 2560 0 -1 1200
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5474_6
timestamp 1731220323
transform 1 0 2448 0 1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5473_6
timestamp 1731220323
transform 1 0 2312 0 1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5472_6
timestamp 1731220323
transform 1 0 2384 0 -1 1060
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5471_6
timestamp 1731220323
transform 1 0 2248 0 -1 1060
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5470_6
timestamp 1731220323
transform 1 0 2288 0 1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5469_6
timestamp 1731220323
transform 1 0 2472 0 -1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5468_6
timestamp 1731220323
transform 1 0 2520 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5467_6
timestamp 1731220323
transform 1 0 2416 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5466_6
timestamp 1731220323
transform 1 0 2328 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5465_6
timestamp 1731220323
transform 1 0 2240 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5464_6
timestamp 1731220323
transform 1 0 2152 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5463_6
timestamp 1731220323
transform 1 0 2552 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5462_6
timestamp 1731220323
transform 1 0 2416 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5461_6
timestamp 1731220323
transform 1 0 2288 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5460_6
timestamp 1731220323
transform 1 0 2168 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5459_6
timestamp 1731220323
transform 1 0 2056 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5458_6
timestamp 1731220323
transform 1 0 2544 0 1 660
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5457_6
timestamp 1731220323
transform 1 0 2384 0 1 660
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5456_6
timestamp 1731220323
transform 1 0 2224 0 1 660
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5455_6
timestamp 1731220323
transform 1 0 2064 0 1 660
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5454_6
timestamp 1731220323
transform 1 0 1920 0 1 660
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5453_6
timestamp 1731220323
transform 1 0 2480 0 -1 652
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5452_6
timestamp 1731220323
transform 1 0 2304 0 -1 652
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5451_6
timestamp 1731220323
transform 1 0 2128 0 -1 652
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5450_6
timestamp 1731220323
transform 1 0 1960 0 -1 652
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5449_6
timestamp 1731220323
transform 1 0 1824 0 -1 652
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5448_6
timestamp 1731220323
transform 1 0 2280 0 1 524
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5447_6
timestamp 1731220323
transform 1 0 2120 0 1 524
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5446_6
timestamp 1731220323
transform 1 0 1960 0 1 524
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5445_6
timestamp 1731220323
transform 1 0 1824 0 1 524
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5444_6
timestamp 1731220323
transform 1 0 1664 0 1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5443_6
timestamp 1731220323
transform 1 0 1664 0 -1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5442_6
timestamp 1731220323
transform 1 0 1568 0 -1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5441_6
timestamp 1731220323
transform 1 0 1824 0 -1 508
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5440_6
timestamp 1731220323
transform 1 0 2120 0 -1 508
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5439_6
timestamp 1731220323
transform 1 0 1960 0 -1 508
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5438_6
timestamp 1731220323
transform 1 0 1952 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5437_6
timestamp 1731220323
transform 1 0 1824 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5436_6
timestamp 1731220323
transform 1 0 1664 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5435_6
timestamp 1731220323
transform 1 0 1560 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5434_6
timestamp 1731220323
transform 1 0 1432 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5433_6
timestamp 1731220323
transform 1 0 1304 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5432_6
timestamp 1731220323
transform 1 0 1224 0 -1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5431_6
timestamp 1731220323
transform 1 0 1344 0 -1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5430_6
timestamp 1731220323
transform 1 0 1456 0 -1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5429_6
timestamp 1731220323
transform 1 0 1352 0 1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5428_6
timestamp 1731220323
transform 1 0 1464 0 1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5427_6
timestamp 1731220323
transform 1 0 1576 0 1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5426_6
timestamp 1731220323
transform 1 0 1576 0 -1 652
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5425_6
timestamp 1731220323
transform 1 0 1440 0 -1 652
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5424_6
timestamp 1731220323
transform 1 0 1304 0 -1 652
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5423_6
timestamp 1731220323
transform 1 0 1176 0 1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5422_6
timestamp 1731220323
transform 1 0 1336 0 1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5421_6
timestamp 1731220323
transform 1 0 1496 0 1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5420_6
timestamp 1731220323
transform 1 0 1344 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5419_6
timestamp 1731220323
transform 1 0 1184 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5418_6
timestamp 1731220323
transform 1 0 1128 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5417_6
timestamp 1731220323
transform 1 0 1000 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5416_6
timestamp 1731220323
transform 1 0 1264 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5415_6
timestamp 1731220323
transform 1 0 1328 0 -1 924
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5414_6
timestamp 1731220323
transform 1 0 1112 0 -1 924
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5413_6
timestamp 1731220323
transform 1 0 872 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5412_6
timestamp 1731220323
transform 1 0 744 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5411_6
timestamp 1731220323
transform 1 0 736 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5410_6
timestamp 1731220323
transform 1 0 880 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5409_6
timestamp 1731220323
transform 1 0 1032 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5408_6
timestamp 1731220323
transform 1 0 1024 0 1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5407_6
timestamp 1731220323
transform 1 0 872 0 1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5406_6
timestamp 1731220323
transform 1 0 1048 0 -1 652
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5405_6
timestamp 1731220323
transform 1 0 1176 0 -1 652
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5404_6
timestamp 1731220323
transform 1 0 1248 0 1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5403_6
timestamp 1731220323
transform 1 0 1144 0 1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5402_6
timestamp 1731220323
transform 1 0 1104 0 -1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5401_6
timestamp 1731220323
transform 1 0 976 0 -1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5400_6
timestamp 1731220323
transform 1 0 896 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5399_6
timestamp 1731220323
transform 1 0 1040 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5398_6
timestamp 1731220323
transform 1 0 1176 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5397_6
timestamp 1731220323
transform 1 0 2104 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5396_6
timestamp 1731220323
transform 1 0 2032 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5395_6
timestamp 1731220323
transform 1 0 1920 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5394_6
timestamp 1731220323
transform 1 0 2152 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5393_6
timestamp 1731220323
transform 1 0 2280 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5392_6
timestamp 1731220323
transform 1 0 2416 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5391_6
timestamp 1731220323
transform 1 0 2392 0 1 248
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5390_6
timestamp 1731220323
transform 1 0 2304 0 1 248
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5389_6
timestamp 1731220323
transform 1 0 2216 0 1 248
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5388_6
timestamp 1731220323
transform 1 0 2480 0 1 248
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5387_6
timestamp 1731220323
transform 1 0 2568 0 1 248
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5386_6
timestamp 1731220323
transform 1 0 2632 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5385_6
timestamp 1731220323
transform 1 0 2504 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5384_6
timestamp 1731220323
transform 1 0 2376 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5383_6
timestamp 1731220323
transform 1 0 2256 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5382_6
timestamp 1731220323
transform 1 0 2136 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5381_6
timestamp 1731220323
transform 1 0 2400 0 1 88
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5380_6
timestamp 1731220323
transform 1 0 2288 0 1 88
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5379_6
timestamp 1731220323
transform 1 0 2176 0 1 88
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5378_6
timestamp 1731220323
transform 1 0 2088 0 1 88
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5377_6
timestamp 1731220323
transform 1 0 2000 0 1 88
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5376_6
timestamp 1731220323
transform 1 0 1912 0 1 88
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5375_6
timestamp 1731220323
transform 1 0 1824 0 1 88
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5374_6
timestamp 1731220323
transform 1 0 1664 0 1 84
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5373_6
timestamp 1731220323
transform 1 0 1576 0 1 84
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5372_6
timestamp 1731220323
transform 1 0 1488 0 1 84
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5371_6
timestamp 1731220323
transform 1 0 1400 0 1 84
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5370_6
timestamp 1731220323
transform 1 0 1312 0 1 84
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5369_6
timestamp 1731220323
transform 1 0 1224 0 1 84
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5368_6
timestamp 1731220323
transform 1 0 1136 0 1 84
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5367_6
timestamp 1731220323
transform 1 0 1048 0 1 84
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5366_6
timestamp 1731220323
transform 1 0 960 0 1 84
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5365_6
timestamp 1731220323
transform 1 0 1096 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5364_6
timestamp 1731220323
transform 1 0 1200 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5363_6
timestamp 1731220323
transform 1 0 1304 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5362_6
timestamp 1731220323
transform 1 0 1232 0 1 244
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5361_6
timestamp 1731220323
transform 1 0 1120 0 1 244
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5360_6
timestamp 1731220323
transform 1 0 1016 0 1 244
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5359_6
timestamp 1731220323
transform 1 0 1200 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5358_6
timestamp 1731220323
transform 1 0 1072 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5357_6
timestamp 1731220323
transform 1 0 952 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5356_6
timestamp 1731220323
transform 1 0 832 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5355_6
timestamp 1731220323
transform 1 0 712 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5354_6
timestamp 1731220323
transform 1 0 808 0 1 244
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5353_6
timestamp 1731220323
transform 1 0 912 0 1 244
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5352_6
timestamp 1731220323
transform 1 0 992 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5351_6
timestamp 1731220323
transform 1 0 800 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5350_6
timestamp 1731220323
transform 1 0 704 0 1 244
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5349_6
timestamp 1731220323
transform 1 0 704 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5348_6
timestamp 1731220323
transform 1 0 616 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5347_6
timestamp 1731220323
transform 1 0 896 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5346_6
timestamp 1731220323
transform 1 0 872 0 1 84
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5345_6
timestamp 1731220323
transform 1 0 784 0 1 84
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5344_6
timestamp 1731220323
transform 1 0 696 0 1 84
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5343_6
timestamp 1731220323
transform 1 0 608 0 1 84
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5342_6
timestamp 1731220323
transform 1 0 520 0 1 84
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5341_6
timestamp 1731220323
transform 1 0 432 0 1 84
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5340_6
timestamp 1731220323
transform 1 0 344 0 1 84
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5339_6
timestamp 1731220323
transform 1 0 256 0 1 84
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5338_6
timestamp 1731220323
transform 1 0 440 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5337_6
timestamp 1731220323
transform 1 0 528 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5336_6
timestamp 1731220323
transform 1 0 592 0 1 244
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5335_6
timestamp 1731220323
transform 1 0 480 0 1 244
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5334_6
timestamp 1731220323
transform 1 0 368 0 1 244
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5333_6
timestamp 1731220323
transform 1 0 256 0 1 244
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5332_6
timestamp 1731220323
transform 1 0 592 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5331_6
timestamp 1731220323
transform 1 0 464 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5330_6
timestamp 1731220323
transform 1 0 336 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5329_6
timestamp 1731220323
transform 1 0 216 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5328_6
timestamp 1731220323
transform 1 0 128 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5327_6
timestamp 1731220323
transform 1 0 128 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5326_6
timestamp 1731220323
transform 1 0 248 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5325_6
timestamp 1731220323
transform 1 0 408 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5324_6
timestamp 1731220323
transform 1 0 736 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5323_6
timestamp 1731220323
transform 1 0 576 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5322_6
timestamp 1731220323
transform 1 0 560 0 -1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5321_6
timestamp 1731220323
transform 1 0 424 0 -1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5320_6
timestamp 1731220323
transform 1 0 296 0 -1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5319_6
timestamp 1731220323
transform 1 0 696 0 -1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5318_6
timestamp 1731220323
transform 1 0 840 0 -1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5317_6
timestamp 1731220323
transform 1 0 808 0 1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5316_6
timestamp 1731220323
transform 1 0 696 0 1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5315_6
timestamp 1731220323
transform 1 0 592 0 1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5314_6
timestamp 1731220323
transform 1 0 1032 0 1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5313_6
timestamp 1731220323
transform 1 0 920 0 1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5312_6
timestamp 1731220323
transform 1 0 920 0 -1 652
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5311_6
timestamp 1731220323
transform 1 0 792 0 -1 652
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5310_6
timestamp 1731220323
transform 1 0 672 0 -1 652
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5309_6
timestamp 1731220323
transform 1 0 552 0 -1 652
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5308_6
timestamp 1731220323
transform 1 0 448 0 -1 652
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5307_6
timestamp 1731220323
transform 1 0 720 0 1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5306_6
timestamp 1731220323
transform 1 0 568 0 1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5305_6
timestamp 1731220323
transform 1 0 424 0 1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5304_6
timestamp 1731220323
transform 1 0 288 0 1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5303_6
timestamp 1731220323
transform 1 0 160 0 1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5302_6
timestamp 1731220323
transform 1 0 600 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5301_6
timestamp 1731220323
transform 1 0 464 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5300_6
timestamp 1731220323
transform 1 0 336 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5299_6
timestamp 1731220323
transform 1 0 216 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5298_6
timestamp 1731220323
transform 1 0 128 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5297_6
timestamp 1731220323
transform 1 0 128 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5296_6
timestamp 1731220323
transform 1 0 224 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5295_6
timestamp 1731220323
transform 1 0 352 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5294_6
timestamp 1731220323
transform 1 0 480 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5293_6
timestamp 1731220323
transform 1 0 616 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5292_6
timestamp 1731220323
transform 1 0 552 0 -1 924
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5291_6
timestamp 1731220323
transform 1 0 408 0 -1 924
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5290_6
timestamp 1731220323
transform 1 0 720 0 -1 924
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5289_6
timestamp 1731220323
transform 1 0 904 0 -1 924
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5288_6
timestamp 1731220323
transform 1 0 1024 0 1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5287_6
timestamp 1731220323
transform 1 0 904 0 1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5286_6
timestamp 1731220323
transform 1 0 784 0 1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5285_6
timestamp 1731220323
transform 1 0 672 0 1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5284_6
timestamp 1731220323
transform 1 0 560 0 1 928
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5283_6
timestamp 1731220323
transform 1 0 912 0 -1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5282_6
timestamp 1731220323
transform 1 0 784 0 -1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5281_6
timestamp 1731220323
transform 1 0 656 0 -1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5280_6
timestamp 1731220323
transform 1 0 536 0 -1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5279_6
timestamp 1731220323
transform 1 0 424 0 -1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5278_6
timestamp 1731220323
transform 1 0 752 0 1 1068
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5277_6
timestamp 1731220323
transform 1 0 616 0 1 1068
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5276_6
timestamp 1731220323
transform 1 0 488 0 1 1068
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5275_6
timestamp 1731220323
transform 1 0 360 0 1 1068
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5274_6
timestamp 1731220323
transform 1 0 240 0 1 1068
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5273_6
timestamp 1731220323
transform 1 0 608 0 -1 1200
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5272_6
timestamp 1731220323
transform 1 0 480 0 -1 1200
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5271_6
timestamp 1731220323
transform 1 0 352 0 -1 1200
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5270_6
timestamp 1731220323
transform 1 0 224 0 -1 1200
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5269_6
timestamp 1731220323
transform 1 0 128 0 -1 1200
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5268_6
timestamp 1731220323
transform 1 0 544 0 1 1208
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5267_6
timestamp 1731220323
transform 1 0 424 0 1 1208
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5266_6
timestamp 1731220323
transform 1 0 312 0 1 1208
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5265_6
timestamp 1731220323
transform 1 0 216 0 1 1208
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5264_6
timestamp 1731220323
transform 1 0 128 0 1 1208
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5263_6
timestamp 1731220323
transform 1 0 552 0 -1 1340
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5262_6
timestamp 1731220323
transform 1 0 392 0 -1 1340
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5261_6
timestamp 1731220323
transform 1 0 240 0 -1 1340
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5260_6
timestamp 1731220323
transform 1 0 128 0 -1 1340
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5259_6
timestamp 1731220323
transform 1 0 128 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5258_6
timestamp 1731220323
transform 1 0 296 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5257_6
timestamp 1731220323
transform 1 0 488 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5256_6
timestamp 1731220323
transform 1 0 368 0 -1 1476
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5255_6
timestamp 1731220323
transform 1 0 152 0 -1 1476
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5254_6
timestamp 1731220323
transform 1 0 176 0 1 1480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5253_6
timestamp 1731220323
transform 1 0 320 0 1 1480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5252_6
timestamp 1731220323
transform 1 0 464 0 1 1480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5251_6
timestamp 1731220323
transform 1 0 376 0 -1 1616
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5250_6
timestamp 1731220323
transform 1 0 272 0 -1 1616
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5249_6
timestamp 1731220323
transform 1 0 488 0 -1 1616
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5248_6
timestamp 1731220323
transform 1 0 480 0 1 1620
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5247_6
timestamp 1731220323
transform 1 0 392 0 1 1620
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5246_6
timestamp 1731220323
transform 1 0 432 0 -1 1752
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5245_6
timestamp 1731220323
transform 1 0 528 0 -1 1752
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5244_6
timestamp 1731220323
transform 1 0 632 0 -1 1752
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5243_6
timestamp 1731220323
transform 1 0 624 0 1 1756
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5242_6
timestamp 1731220323
transform 1 0 504 0 1 1756
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5241_6
timestamp 1731220323
transform 1 0 424 0 -1 1888
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5240_6
timestamp 1731220323
transform 1 0 568 0 -1 1888
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5239_6
timestamp 1731220323
transform 1 0 720 0 -1 1888
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5238_6
timestamp 1731220323
transform 1 0 696 0 1 1888
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5237_6
timestamp 1731220323
transform 1 0 552 0 1 1888
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5236_6
timestamp 1731220323
transform 1 0 416 0 1 1888
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5235_6
timestamp 1731220323
transform 1 0 288 0 1 1888
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5234_6
timestamp 1731220323
transform 1 0 632 0 -1 2020
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5233_6
timestamp 1731220323
transform 1 0 496 0 -1 2020
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5232_6
timestamp 1731220323
transform 1 0 360 0 -1 2020
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5231_6
timestamp 1731220323
transform 1 0 232 0 -1 2020
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5230_6
timestamp 1731220323
transform 1 0 128 0 -1 2020
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5229_6
timestamp 1731220323
transform 1 0 576 0 1 2028
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5228_6
timestamp 1731220323
transform 1 0 456 0 1 2028
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5227_6
timestamp 1731220323
transform 1 0 336 0 1 2028
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5226_6
timestamp 1731220323
transform 1 0 216 0 1 2028
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5225_6
timestamp 1731220323
transform 1 0 128 0 1 2028
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5224_6
timestamp 1731220323
transform 1 0 688 0 -1 2160
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5223_6
timestamp 1731220323
transform 1 0 536 0 -1 2160
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5222_6
timestamp 1731220323
transform 1 0 384 0 -1 2160
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5221_6
timestamp 1731220323
transform 1 0 240 0 -1 2160
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5220_6
timestamp 1731220323
transform 1 0 128 0 -1 2160
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5219_6
timestamp 1731220323
transform 1 0 128 0 1 2168
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5218_6
timestamp 1731220323
transform 1 0 240 0 1 2168
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5217_6
timestamp 1731220323
transform 1 0 760 0 1 2168
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5216_6
timestamp 1731220323
transform 1 0 576 0 1 2168
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5215_6
timestamp 1731220323
transform 1 0 400 0 1 2168
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5214_6
timestamp 1731220323
transform 1 0 264 0 -1 2300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5213_6
timestamp 1731220323
transform 1 0 144 0 -1 2300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5212_6
timestamp 1731220323
transform 1 0 640 0 -1 2300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5211_6
timestamp 1731220323
transform 1 0 512 0 -1 2300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5210_6
timestamp 1731220323
transform 1 0 384 0 -1 2300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5209_6
timestamp 1731220323
transform 1 0 312 0 1 2308
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5208_6
timestamp 1731220323
transform 1 0 424 0 1 2308
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5207_6
timestamp 1731220323
transform 1 0 648 0 1 2308
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5206_6
timestamp 1731220323
transform 1 0 536 0 1 2308
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5205_6
timestamp 1731220323
transform 1 0 496 0 -1 2440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5204_6
timestamp 1731220323
transform 1 0 408 0 -1 2440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5203_6
timestamp 1731220323
transform 1 0 592 0 -1 2440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5202_6
timestamp 1731220323
transform 1 0 544 0 1 2440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5201_6
timestamp 1731220323
transform 1 0 728 0 1 2440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5200_6
timestamp 1731220323
transform 1 0 904 0 1 2440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5199_6
timestamp 1731220323
transform 1 0 912 0 -1 2440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5198_6
timestamp 1731220323
transform 1 0 800 0 -1 2440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5197_6
timestamp 1731220323
transform 1 0 696 0 -1 2440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5196_6
timestamp 1731220323
transform 1 0 1032 0 -1 2440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5195_6
timestamp 1731220323
transform 1 0 984 0 1 2308
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5194_6
timestamp 1731220323
transform 1 0 872 0 1 2308
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5193_6
timestamp 1731220323
transform 1 0 760 0 1 2308
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5192_6
timestamp 1731220323
transform 1 0 768 0 -1 2300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5191_6
timestamp 1731220323
transform 1 0 888 0 -1 2300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5190_6
timestamp 1731220323
transform 1 0 944 0 1 2168
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5189_6
timestamp 1731220323
transform 1 0 1128 0 1 2168
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5188_6
timestamp 1731220323
transform 1 0 1264 0 -1 2300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5187_6
timestamp 1731220323
transform 1 0 1136 0 -1 2300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5186_6
timestamp 1731220323
transform 1 0 1008 0 -1 2300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5185_6
timestamp 1731220323
transform 1 0 1096 0 1 2308
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5184_6
timestamp 1731220323
transform 1 0 1208 0 1 2308
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5183_6
timestamp 1731220323
transform 1 0 1328 0 1 2308
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5182_6
timestamp 1731220323
transform 1 0 1416 0 -1 2440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5181_6
timestamp 1731220323
transform 1 0 1288 0 -1 2440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5180_6
timestamp 1731220323
transform 1 0 1160 0 -1 2440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5179_6
timestamp 1731220323
transform 1 0 1072 0 1 2440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5178_6
timestamp 1731220323
transform 1 0 1232 0 1 2440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5177_6
timestamp 1731220323
transform 1 0 1560 0 1 2440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5176_6
timestamp 1731220323
transform 1 0 1392 0 1 2440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5175_6
timestamp 1731220323
transform 1 0 1344 0 -1 2576
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5174_6
timestamp 1731220323
transform 1 0 1472 0 -1 2576
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5173_6
timestamp 1731220323
transform 1 0 1600 0 -1 2576
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5172_6
timestamp 1731220323
transform 1 0 1600 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5171_6
timestamp 1731220323
transform 1 0 1432 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5170_6
timestamp 1731220323
transform 1 0 1368 0 -1 2720
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5169_6
timestamp 1731220323
transform 1 0 1664 0 -1 2720
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5168_6
timestamp 1731220323
transform 1 0 1528 0 -1 2720
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5167_6
timestamp 1731220323
transform 1 0 1520 0 1 2728
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5166_6
timestamp 1731220323
transform 1 0 1664 0 1 2728
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5165_6
timestamp 1731220323
transform 1 0 1824 0 1 2740
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5164_6
timestamp 1731220323
transform 1 0 1824 0 -1 2872
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5163_6
timestamp 1731220323
transform 1 0 1992 0 -1 2872
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5162_6
timestamp 1731220323
transform 1 0 2008 0 1 2872
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5161_6
timestamp 1731220323
transform 1 0 1824 0 1 2872
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5160_6
timestamp 1731220323
transform 1 0 1824 0 -1 3012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5159_6
timestamp 1731220323
transform 1 0 1912 0 -1 3012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5158_6
timestamp 1731220323
transform 1 0 2024 0 -1 3012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5157_6
timestamp 1731220323
transform 1 0 2288 0 1 3028
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5156_6
timestamp 1731220323
transform 1 0 2112 0 1 3028
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5155_6
timestamp 1731220323
transform 1 0 1952 0 1 3028
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5154_6
timestamp 1731220323
transform 1 0 1824 0 1 3028
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5153_6
timestamp 1731220323
transform 1 0 1824 0 -1 3164
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5152_6
timestamp 1731220323
transform 1 0 2000 0 -1 3164
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5151_6
timestamp 1731220323
transform 1 0 2392 0 -1 3164
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5150_6
timestamp 1731220323
transform 1 0 2200 0 -1 3164
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5149_6
timestamp 1731220323
transform 1 0 2192 0 1 3164
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5148_6
timestamp 1731220323
transform 1 0 2040 0 1 3164
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5147_6
timestamp 1731220323
transform 1 0 1904 0 1 3164
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5146_6
timestamp 1731220323
transform 1 0 2520 0 1 3164
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5145_6
timestamp 1731220323
transform 1 0 2352 0 1 3164
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5144_6
timestamp 1731220323
transform 1 0 2232 0 -1 3296
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5143_6
timestamp 1731220323
transform 1 0 2080 0 -1 3296
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5142_6
timestamp 1731220323
transform 1 0 2392 0 -1 3296
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5141_6
timestamp 1731220323
transform 1 0 2552 0 -1 3296
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5140_6
timestamp 1731220323
transform 1 0 2560 0 1 3296
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5139_6
timestamp 1731220323
transform 1 0 2424 0 1 3296
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5138_6
timestamp 1731220323
transform 1 0 2288 0 1 3296
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5137_6
timestamp 1731220323
transform 1 0 2152 0 1 3296
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5136_6
timestamp 1731220323
transform 1 0 2384 0 -1 3428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5135_6
timestamp 1731220323
transform 1 0 2264 0 -1 3428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5134_6
timestamp 1731220323
transform 1 0 2144 0 -1 3428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5133_6
timestamp 1731220323
transform 1 0 2024 0 -1 3428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5132_6
timestamp 1731220323
transform 1 0 2304 0 1 3428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5131_6
timestamp 1731220323
transform 1 0 2136 0 1 3428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5130_6
timestamp 1731220323
transform 1 0 1968 0 1 3428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5129_6
timestamp 1731220323
transform 1 0 1824 0 1 3428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5128_6
timestamp 1731220323
transform 1 0 1664 0 1 3440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5127_6
timestamp 1731220323
transform 1 0 1544 0 1 3440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5126_6
timestamp 1731220323
transform 1 0 1400 0 1 3440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5125_6
timestamp 1731220323
transform 1 0 1256 0 1 3440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5124_6
timestamp 1731220323
transform 1 0 1112 0 1 3440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5123_6
timestamp 1731220323
transform 1 0 952 0 1 3440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5122_6
timestamp 1731220323
transform 1 0 1392 0 -1 3436
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5121_6
timestamp 1731220323
transform 1 0 1224 0 -1 3436
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5120_6
timestamp 1731220323
transform 1 0 1056 0 -1 3436
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5119_6
timestamp 1731220323
transform 1 0 888 0 -1 3436
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5118_6
timestamp 1731220323
transform 1 0 928 0 1 3300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5117_6
timestamp 1731220323
transform 1 0 1112 0 1 3300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5116_6
timestamp 1731220323
transform 1 0 1288 0 1 3300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5115_6
timestamp 1731220323
transform 1 0 1456 0 1 3300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5114_6
timestamp 1731220323
transform 1 0 1632 0 1 3300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5113_6
timestamp 1731220323
transform 1 0 1664 0 -1 3292
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5112_6
timestamp 1731220323
transform 1 0 1496 0 -1 3292
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5111_6
timestamp 1731220323
transform 1 0 1336 0 -1 3292
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5110_6
timestamp 1731220323
transform 1 0 1168 0 -1 3292
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5109_6
timestamp 1731220323
transform 1 0 1000 0 -1 3292
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5108_6
timestamp 1731220323
transform 1 0 1464 0 1 3156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5107_6
timestamp 1731220323
transform 1 0 1296 0 1 3156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5106_6
timestamp 1731220323
transform 1 0 1128 0 1 3156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5105_6
timestamp 1731220323
transform 1 0 960 0 1 3156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5104_6
timestamp 1731220323
transform 1 0 1312 0 -1 3156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5103_6
timestamp 1731220323
transform 1 0 1192 0 -1 3156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5102_6
timestamp 1731220323
transform 1 0 1072 0 -1 3156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5101_6
timestamp 1731220323
transform 1 0 960 0 -1 3156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5100_6
timestamp 1731220323
transform 1 0 840 0 -1 3156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_599_6
timestamp 1731220323
transform 1 0 1136 0 1 3024
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_598_6
timestamp 1731220323
transform 1 0 1048 0 1 3024
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_597_6
timestamp 1731220323
transform 1 0 960 0 1 3024
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_596_6
timestamp 1731220323
transform 1 0 872 0 1 3024
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_595_6
timestamp 1731220323
transform 1 0 936 0 -1 3016
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_594_6
timestamp 1731220323
transform 1 0 1024 0 -1 3016
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_593_6
timestamp 1731220323
transform 1 0 1288 0 -1 3016
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_592_6
timestamp 1731220323
transform 1 0 1200 0 -1 3016
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_591_6
timestamp 1731220323
transform 1 0 1112 0 -1 3016
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_590_6
timestamp 1731220323
transform 1 0 1096 0 1 2876
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_589_6
timestamp 1731220323
transform 1 0 968 0 1 2876
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_588_6
timestamp 1731220323
transform 1 0 1224 0 1 2876
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_587_6
timestamp 1731220323
transform 1 0 1352 0 1 2876
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_586_6
timestamp 1731220323
transform 1 0 1488 0 1 2876
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_585_6
timestamp 1731220323
transform 1 0 1488 0 -1 2868
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_584_6
timestamp 1731220323
transform 1 0 1336 0 -1 2868
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_583_6
timestamp 1731220323
transform 1 0 1184 0 -1 2868
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_582_6
timestamp 1731220323
transform 1 0 1040 0 -1 2868
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_581_6
timestamp 1731220323
transform 1 0 888 0 -1 2868
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_580_6
timestamp 1731220323
transform 1 0 1352 0 1 2728
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_579_6
timestamp 1731220323
transform 1 0 1184 0 1 2728
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_578_6
timestamp 1731220323
transform 1 0 1016 0 1 2728
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_577_6
timestamp 1731220323
transform 1 0 848 0 1 2728
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_576_6
timestamp 1731220323
transform 1 0 904 0 -1 2720
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_575_6
timestamp 1731220323
transform 1 0 1208 0 -1 2720
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_574_6
timestamp 1731220323
transform 1 0 1056 0 -1 2720
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_573_6
timestamp 1731220323
transform 1 0 976 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_572_6
timestamp 1731220323
transform 1 0 1120 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_571_6
timestamp 1731220323
transform 1 0 1272 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_570_6
timestamp 1731220323
transform 1 0 1216 0 -1 2576
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_569_6
timestamp 1731220323
transform 1 0 1096 0 -1 2576
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_568_6
timestamp 1731220323
transform 1 0 984 0 -1 2576
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_567_6
timestamp 1731220323
transform 1 0 872 0 -1 2576
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_566_6
timestamp 1731220323
transform 1 0 768 0 -1 2576
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_565_6
timestamp 1731220323
transform 1 0 672 0 -1 2576
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_564_6
timestamp 1731220323
transform 1 0 584 0 -1 2576
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_563_6
timestamp 1731220323
transform 1 0 496 0 -1 2576
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_562_6
timestamp 1731220323
transform 1 0 848 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_561_6
timestamp 1731220323
transform 1 0 736 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_560_6
timestamp 1731220323
transform 1 0 632 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_559_6
timestamp 1731220323
transform 1 0 544 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_558_6
timestamp 1731220323
transform 1 0 456 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_557_6
timestamp 1731220323
transform 1 0 752 0 -1 2720
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_556_6
timestamp 1731220323
transform 1 0 608 0 -1 2720
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_555_6
timestamp 1731220323
transform 1 0 472 0 -1 2720
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_554_6
timestamp 1731220323
transform 1 0 352 0 -1 2720
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_553_6
timestamp 1731220323
transform 1 0 240 0 -1 2720
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_552_6
timestamp 1731220323
transform 1 0 688 0 1 2728
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_551_6
timestamp 1731220323
transform 1 0 536 0 1 2728
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_550_6
timestamp 1731220323
transform 1 0 384 0 1 2728
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_549_6
timestamp 1731220323
transform 1 0 240 0 1 2728
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_548_6
timestamp 1731220323
transform 1 0 128 0 1 2728
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_547_6
timestamp 1731220323
transform 1 0 128 0 -1 2868
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_546_6
timestamp 1731220323
transform 1 0 248 0 -1 2868
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_545_6
timestamp 1731220323
transform 1 0 408 0 -1 2868
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_544_6
timestamp 1731220323
transform 1 0 728 0 -1 2868
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_543_6
timestamp 1731220323
transform 1 0 568 0 -1 2868
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_542_6
timestamp 1731220323
transform 1 0 568 0 1 2876
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_541_6
timestamp 1731220323
transform 1 0 440 0 1 2876
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_540_6
timestamp 1731220323
transform 1 0 320 0 1 2876
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_539_6
timestamp 1731220323
transform 1 0 840 0 1 2876
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_538_6
timestamp 1731220323
transform 1 0 704 0 1 2876
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_537_6
timestamp 1731220323
transform 1 0 672 0 -1 3016
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_536_6
timestamp 1731220323
transform 1 0 584 0 -1 3016
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_535_6
timestamp 1731220323
transform 1 0 496 0 -1 3016
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_534_6
timestamp 1731220323
transform 1 0 760 0 -1 3016
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_533_6
timestamp 1731220323
transform 1 0 848 0 -1 3016
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_532_6
timestamp 1731220323
transform 1 0 784 0 1 3024
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_531_6
timestamp 1731220323
transform 1 0 696 0 1 3024
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_530_6
timestamp 1731220323
transform 1 0 608 0 1 3024
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_529_6
timestamp 1731220323
transform 1 0 520 0 1 3024
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_528_6
timestamp 1731220323
transform 1 0 432 0 1 3024
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_527_6
timestamp 1731220323
transform 1 0 720 0 -1 3156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_526_6
timestamp 1731220323
transform 1 0 600 0 -1 3156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_525_6
timestamp 1731220323
transform 1 0 480 0 -1 3156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_524_6
timestamp 1731220323
transform 1 0 360 0 -1 3156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_523_6
timestamp 1731220323
transform 1 0 800 0 1 3156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_522_6
timestamp 1731220323
transform 1 0 640 0 1 3156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_521_6
timestamp 1731220323
transform 1 0 480 0 1 3156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_520_6
timestamp 1731220323
transform 1 0 320 0 1 3156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_519_6
timestamp 1731220323
transform 1 0 176 0 1 3156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_518_6
timestamp 1731220323
transform 1 0 824 0 -1 3292
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_517_6
timestamp 1731220323
transform 1 0 640 0 -1 3292
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_516_6
timestamp 1731220323
transform 1 0 456 0 -1 3292
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_515_6
timestamp 1731220323
transform 1 0 272 0 -1 3292
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_514_6
timestamp 1731220323
transform 1 0 128 0 -1 3292
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_513_6
timestamp 1731220323
transform 1 0 128 0 1 3300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_512_6
timestamp 1731220323
transform 1 0 320 0 1 3300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_511_6
timestamp 1731220323
transform 1 0 736 0 1 3300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_510_6
timestamp 1731220323
transform 1 0 528 0 1 3300
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_59_6
timestamp 1731220323
transform 1 0 408 0 -1 3436
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_58_6
timestamp 1731220323
transform 1 0 248 0 -1 3436
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_57_6
timestamp 1731220323
transform 1 0 128 0 -1 3436
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_56_6
timestamp 1731220323
transform 1 0 568 0 -1 3436
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_55_6
timestamp 1731220323
transform 1 0 728 0 -1 3436
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_54_6
timestamp 1731220323
transform 1 0 784 0 1 3440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_53_6
timestamp 1731220323
transform 1 0 608 0 1 3440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_52_6
timestamp 1731220323
transform 1 0 432 0 1 3440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_51_6
timestamp 1731220323
transform 1 0 264 0 1 3440
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_50_6
timestamp 1731220323
transform 1 0 128 0 1 3440
box 8 4 84 60
<< end >>
