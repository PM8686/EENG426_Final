magic
tech TSMC180
timestamp 1734143796
<< ndiffusion >>
rect 6 21 12 22
rect 6 19 7 21
rect 9 19 12 21
rect 6 12 12 19
rect 14 15 20 22
rect 14 13 17 15
rect 19 13 20 15
rect 14 12 20 13
rect 22 21 28 22
rect 22 19 25 21
rect 27 19 28 21
rect 22 12 28 19
rect 32 21 38 22
rect 32 19 35 21
rect 37 19 38 21
rect 32 12 38 19
rect 40 15 48 22
rect 40 13 43 15
rect 45 13 48 15
rect 40 12 48 13
rect 50 21 56 22
rect 50 19 53 21
rect 55 19 56 21
rect 50 12 56 19
rect 60 21 66 22
rect 60 19 61 21
rect 63 19 66 21
rect 60 12 66 19
rect 68 15 76 22
rect 68 13 69 15
rect 71 13 76 15
rect 68 12 76 13
rect 78 21 84 22
rect 78 19 79 21
rect 81 19 84 21
rect 78 12 84 19
<< ndcontact >>
rect 7 19 9 21
rect 17 13 19 15
rect 25 19 27 21
rect 35 19 37 21
rect 43 13 45 15
rect 53 19 55 21
rect 61 19 63 21
rect 69 13 71 15
rect 79 19 81 21
<< ntransistor >>
rect 12 12 14 22
rect 20 12 22 22
rect 38 12 40 22
rect 48 12 50 22
rect 66 12 68 22
rect 76 12 78 22
<< pdiffusion >>
rect 6 52 12 53
rect 6 50 7 52
rect 9 50 12 52
rect 6 38 12 50
rect 14 52 20 53
rect 14 50 17 52
rect 19 50 20 52
rect 14 38 20 50
rect 22 41 28 53
rect 44 48 48 58
rect 22 39 25 41
rect 27 39 28 41
rect 22 38 28 39
rect 32 41 38 48
rect 32 39 35 41
rect 37 39 38 41
rect 32 38 38 39
rect 40 41 48 48
rect 40 39 43 41
rect 45 39 48 41
rect 40 38 48 39
rect 50 57 56 58
rect 50 55 53 57
rect 55 55 56 57
rect 50 38 56 55
rect 72 57 76 58
rect 72 55 73 57
rect 75 55 76 57
rect 72 48 76 55
rect 60 41 66 48
rect 60 39 61 41
rect 63 39 66 41
rect 60 38 66 39
rect 68 38 76 48
rect 78 57 84 58
rect 78 55 80 57
rect 82 55 84 57
rect 78 38 84 55
<< pdcontact >>
rect 7 50 9 52
rect 17 50 19 52
rect 25 39 27 41
rect 35 39 37 41
rect 43 39 45 41
rect 53 55 55 57
rect 73 55 75 57
rect 61 39 63 41
rect 80 55 82 57
<< ptransistor >>
rect 12 38 14 53
rect 20 38 22 53
rect 38 38 40 48
rect 48 38 50 58
rect 66 38 68 48
rect 76 38 78 58
<< polysilicon >>
rect 48 58 50 61
rect 76 58 78 61
rect 30 57 34 58
rect 12 53 14 56
rect 20 55 31 57
rect 33 55 40 57
rect 20 53 22 55
rect 30 54 34 55
rect 38 48 40 55
rect 64 53 68 54
rect 64 51 65 53
rect 67 51 68 53
rect 64 50 68 51
rect 66 48 68 50
rect 12 22 14 38
rect 20 22 22 38
rect 38 22 40 38
rect 48 32 50 38
rect 48 31 52 32
rect 48 29 49 31
rect 51 29 52 31
rect 48 28 52 29
rect 48 22 50 28
rect 66 22 68 38
rect 76 34 78 38
rect 75 33 79 34
rect 75 31 76 33
rect 78 31 79 33
rect 75 30 79 31
rect 76 22 78 30
rect 12 6 14 12
rect 20 9 22 12
rect 38 9 40 12
rect 48 9 50 12
rect 66 9 68 12
rect 76 9 78 12
rect 9 5 14 6
rect 9 3 10 5
rect 12 3 14 5
rect 9 2 14 3
<< polycontact >>
rect 31 55 33 57
rect 65 51 67 53
rect 49 29 51 31
rect 76 31 78 33
rect 10 3 12 5
<< m1 >>
rect 6 53 9 70
rect 14 62 19 63
rect 14 59 15 62
rect 18 59 19 62
rect 14 58 19 59
rect 16 53 19 58
rect 30 58 33 70
rect 53 66 82 69
rect 53 58 56 66
rect 71 62 76 63
rect 71 59 72 62
rect 75 59 76 62
rect 71 58 76 59
rect 30 57 34 58
rect 30 55 31 57
rect 33 55 34 57
rect 30 54 34 55
rect 52 57 56 58
rect 52 55 53 57
rect 55 55 56 57
rect 52 54 56 55
rect 72 57 76 58
rect 72 55 73 57
rect 75 55 76 57
rect 72 54 76 55
rect 79 58 82 66
rect 79 57 83 58
rect 79 55 80 57
rect 82 55 83 57
rect 79 54 83 55
rect 63 53 68 54
rect 6 52 11 53
rect 6 49 7 52
rect 10 49 11 52
rect 16 52 20 53
rect 16 50 17 52
rect 19 50 20 52
rect 16 49 20 50
rect 63 52 65 53
rect 63 49 64 52
rect 67 49 68 53
rect 6 48 11 49
rect 63 48 68 49
rect 6 22 9 48
rect 34 42 39 43
rect 59 42 64 43
rect 24 41 28 42
rect 24 39 25 41
rect 27 39 28 41
rect 24 38 28 39
rect 34 39 35 42
rect 38 39 39 42
rect 34 38 39 39
rect 42 41 46 42
rect 42 39 43 41
rect 45 39 46 41
rect 42 38 46 39
rect 59 39 60 42
rect 63 39 64 42
rect 59 38 64 39
rect 25 33 28 38
rect 25 32 30 33
rect 25 29 26 32
rect 29 29 30 32
rect 25 28 30 29
rect 25 22 28 28
rect 6 21 10 22
rect 6 19 7 21
rect 9 19 10 21
rect 6 18 10 19
rect 24 21 28 22
rect 24 19 25 21
rect 27 19 28 21
rect 24 18 28 19
rect 34 22 39 23
rect 34 19 35 22
rect 38 19 39 22
rect 34 18 39 19
rect 42 16 45 38
rect 75 33 93 34
rect 48 32 53 33
rect 48 29 49 32
rect 52 29 53 32
rect 75 31 76 33
rect 78 31 93 33
rect 75 30 79 31
rect 48 28 53 29
rect 77 22 82 23
rect 52 21 64 22
rect 52 19 53 21
rect 55 19 61 21
rect 63 19 64 21
rect 52 18 64 19
rect 77 19 78 22
rect 81 19 82 22
rect 77 18 82 19
rect 16 15 20 16
rect 16 13 17 15
rect 19 13 20 15
rect 42 15 46 16
rect 42 13 43 15
rect 45 13 46 15
rect 68 15 72 16
rect 68 13 69 15
rect 71 13 72 15
rect 16 12 21 13
rect 16 9 17 12
rect 20 9 21 12
rect 16 8 21 9
rect 42 12 46 13
rect 67 12 72 13
rect 9 5 13 6
rect 42 5 45 12
rect 67 9 68 12
rect 71 9 72 12
rect 67 8 72 9
rect 9 3 10 5
rect 12 3 45 5
rect 9 2 45 3
<< m2c >>
rect 15 59 18 62
rect 72 59 75 62
rect 7 50 9 52
rect 9 50 10 52
rect 7 49 10 50
rect 64 51 65 52
rect 65 51 67 52
rect 64 49 67 51
rect 35 41 38 42
rect 35 39 37 41
rect 37 39 38 41
rect 60 41 63 42
rect 60 39 61 41
rect 61 39 63 41
rect 26 29 29 32
rect 35 21 38 22
rect 35 19 37 21
rect 37 19 38 21
rect 49 31 52 32
rect 49 29 51 31
rect 51 29 52 31
rect 78 21 81 22
rect 78 19 79 21
rect 79 19 81 21
rect 17 9 20 12
rect 68 9 71 12
<< m2 >>
rect 14 62 76 63
rect 14 59 15 62
rect 18 59 72 62
rect 75 59 76 62
rect 14 58 76 59
rect 6 52 68 53
rect 6 49 7 52
rect 10 49 64 52
rect 67 49 68 52
rect 6 48 68 49
rect 34 42 64 43
rect 34 39 35 42
rect 38 39 60 42
rect 63 39 64 42
rect 34 38 64 39
rect 25 32 53 33
rect 25 29 26 32
rect 29 29 49 32
rect 52 29 53 32
rect 25 28 53 29
rect 34 22 82 23
rect 34 19 35 22
rect 38 19 78 22
rect 81 19 82 22
rect 34 18 82 19
rect 16 12 72 13
rect 16 9 17 12
rect 20 9 68 12
rect 71 9 72 12
rect 16 8 72 9
<< labels >>
rlabel m1 s 33 55 34 57 6 CLK
port 1 nsew signal input
rlabel m1 s 31 55 33 57 6 CLK
port 1 nsew signal input
rlabel m1 s 30 54 34 55 6 CLK
port 1 nsew signal input
rlabel m1 s 30 55 31 57 6 CLK
port 1 nsew signal input
rlabel m1 s 30 57 34 58 6 CLK
port 1 nsew signal input
rlabel m1 s 30 58 33 70 6 CLK
port 1 nsew signal input
rlabel m1 s 78 31 93 33 6 D
port 2 nsew signal input
rlabel m1 s 76 31 78 33 6 D
port 2 nsew signal input
rlabel m1 s 75 30 79 31 6 D
port 2 nsew signal input
rlabel m1 s 75 31 76 33 6 D
port 2 nsew signal input
rlabel m1 s 75 33 93 34 6 D
port 2 nsew signal input
rlabel m2 s 67 49 68 52 6 Q
port 3 nsew signal output
rlabel m2 s 65 51 67 52 6 Q
port 3 nsew signal output
rlabel m2 s 64 49 67 51 6 Q
port 3 nsew signal output
rlabel m2 s 64 51 65 52 6 Q
port 3 nsew signal output
rlabel m2 s 10 49 64 52 6 Q
port 3 nsew signal output
rlabel m2 s 9 50 10 52 6 Q
port 3 nsew signal output
rlabel m2 s 7 49 10 50 6 Q
port 3 nsew signal output
rlabel m2 s 7 50 9 52 6 Q
port 3 nsew signal output
rlabel m2 s 6 48 68 49 6 Q
port 3 nsew signal output
rlabel m2 s 6 49 7 52 6 Q
port 3 nsew signal output
rlabel m2 s 6 52 68 53 6 Q
port 3 nsew signal output
rlabel m2c s 65 51 67 52 6 Q
port 3 nsew signal output
rlabel m2c s 64 49 67 51 6 Q
port 3 nsew signal output
rlabel m2c s 64 51 65 52 6 Q
port 3 nsew signal output
rlabel m2c s 9 50 10 52 6 Q
port 3 nsew signal output
rlabel m2c s 7 49 10 50 6 Q
port 3 nsew signal output
rlabel m2c s 7 50 9 52 6 Q
port 3 nsew signal output
rlabel m1 s 67 49 68 53 6 Q
port 3 nsew signal output
rlabel m1 s 65 51 67 52 6 Q
port 3 nsew signal output
rlabel m1 s 64 49 67 51 6 Q
port 3 nsew signal output
rlabel m1 s 64 51 65 52 6 Q
port 3 nsew signal output
rlabel m1 s 65 52 67 53 6 Q
port 3 nsew signal output
rlabel m1 s 63 48 68 49 6 Q
port 3 nsew signal output
rlabel m1 s 63 49 64 52 6 Q
port 3 nsew signal output
rlabel m1 s 63 52 65 53 6 Q
port 3 nsew signal output
rlabel m1 s 63 53 68 54 6 Q
port 3 nsew signal output
rlabel m1 s 9 19 10 21 6 Q
port 3 nsew signal output
rlabel m1 s 10 49 11 52 6 Q
port 3 nsew signal output
rlabel m1 s 9 50 10 52 6 Q
port 3 nsew signal output
rlabel m1 s 7 19 9 21 6 Q
port 3 nsew signal output
rlabel m1 s 7 49 10 50 6 Q
port 3 nsew signal output
rlabel m1 s 7 50 9 52 6 Q
port 3 nsew signal output
rlabel m1 s 6 18 10 19 6 Q
port 3 nsew signal output
rlabel m1 s 6 19 7 21 6 Q
port 3 nsew signal output
rlabel m1 s 6 21 10 22 6 Q
port 3 nsew signal output
rlabel m1 s 6 22 9 48 6 Q
port 3 nsew signal output
rlabel m1 s 6 48 11 49 6 Q
port 3 nsew signal output
rlabel m1 s 6 49 7 52 6 Q
port 3 nsew signal output
rlabel m1 s 6 52 11 53 6 Q
port 3 nsew signal output
rlabel m1 s 6 53 9 70 6 Q
port 3 nsew signal output
rlabel m2 s 75 59 76 62 6 Vdd
port 4 nsew power input
rlabel m2 s 72 59 75 62 6 Vdd
port 4 nsew power input
rlabel m2 s 18 59 72 62 6 Vdd
port 4 nsew power input
rlabel m2 s 15 59 18 62 6 Vdd
port 4 nsew power input
rlabel m2 s 14 58 76 59 6 Vdd
port 4 nsew power input
rlabel m2 s 14 59 15 62 6 Vdd
port 4 nsew power input
rlabel m2 s 14 62 76 63 6 Vdd
port 4 nsew power input
rlabel m2c s 72 59 75 62 6 Vdd
port 4 nsew power input
rlabel m2c s 15 59 18 62 6 Vdd
port 4 nsew power input
rlabel m1 s 75 55 76 57 6 Vdd
port 4 nsew power input
rlabel m1 s 73 55 75 57 6 Vdd
port 4 nsew power input
rlabel m1 s 72 54 76 55 6 Vdd
port 4 nsew power input
rlabel m1 s 72 55 73 57 6 Vdd
port 4 nsew power input
rlabel m1 s 72 57 76 58 6 Vdd
port 4 nsew power input
rlabel m1 s 75 59 76 62 6 Vdd
port 4 nsew power input
rlabel m1 s 72 59 75 62 6 Vdd
port 4 nsew power input
rlabel m1 s 71 58 76 59 6 Vdd
port 4 nsew power input
rlabel m1 s 71 59 72 62 6 Vdd
port 4 nsew power input
rlabel m1 s 71 62 76 63 6 Vdd
port 4 nsew power input
rlabel m1 s 19 50 20 52 6 Vdd
port 4 nsew power input
rlabel m1 s 17 50 19 52 6 Vdd
port 4 nsew power input
rlabel m1 s 16 49 20 50 6 Vdd
port 4 nsew power input
rlabel m1 s 16 50 17 52 6 Vdd
port 4 nsew power input
rlabel m1 s 16 52 20 53 6 Vdd
port 4 nsew power input
rlabel m1 s 16 53 19 58 6 Vdd
port 4 nsew power input
rlabel m1 s 18 59 19 62 6 Vdd
port 4 nsew power input
rlabel m1 s 15 59 18 62 6 Vdd
port 4 nsew power input
rlabel m1 s 14 58 19 59 6 Vdd
port 4 nsew power input
rlabel m1 s 14 59 15 62 6 Vdd
port 4 nsew power input
rlabel m1 s 14 62 19 63 6 Vdd
port 4 nsew power input
rlabel m2 s 71 9 72 12 6 GND
port 5 nsew ground input
rlabel m2 s 68 9 71 12 6 GND
port 5 nsew ground input
rlabel m2 s 20 9 68 12 6 GND
port 5 nsew ground input
rlabel m2 s 17 9 20 12 6 GND
port 5 nsew ground input
rlabel m2 s 16 8 72 9 6 GND
port 5 nsew ground input
rlabel m2 s 16 9 17 12 6 GND
port 5 nsew ground input
rlabel m2 s 16 12 72 13 6 GND
port 5 nsew ground input
rlabel m2c s 68 9 71 12 6 GND
port 5 nsew ground input
rlabel m2c s 17 9 20 12 6 GND
port 5 nsew ground input
rlabel m1 s 71 13 72 15 6 GND
port 5 nsew ground input
rlabel m1 s 69 13 71 15 6 GND
port 5 nsew ground input
rlabel m1 s 68 13 69 15 6 GND
port 5 nsew ground input
rlabel m1 s 68 15 72 16 6 GND
port 5 nsew ground input
rlabel m1 s 71 9 72 12 6 GND
port 5 nsew ground input
rlabel m1 s 68 9 71 12 6 GND
port 5 nsew ground input
rlabel m1 s 67 8 72 9 6 GND
port 5 nsew ground input
rlabel m1 s 67 9 68 12 6 GND
port 5 nsew ground input
rlabel m1 s 67 12 72 13 6 GND
port 5 nsew ground input
rlabel m1 s 20 9 21 12 6 GND
port 5 nsew ground input
rlabel m1 s 19 13 20 15 6 GND
port 5 nsew ground input
rlabel m1 s 17 9 20 12 6 GND
port 5 nsew ground input
rlabel m1 s 17 13 19 15 6 GND
port 5 nsew ground input
rlabel m1 s 16 8 21 9 6 GND
port 5 nsew ground input
rlabel m1 s 16 9 17 12 6 GND
port 5 nsew ground input
rlabel m1 s 16 12 21 13 6 GND
port 5 nsew ground input
rlabel m1 s 16 13 17 15 6 GND
port 5 nsew ground input
rlabel m1 s 16 15 20 16 6 GND
port 5 nsew ground input
rlabel space 0 0 96 80 1 prboundary
rlabel polysilicon 77 23 77 23 3 D
rlabel polysilicon 77 35 77 35 3 D
rlabel polysilicon 77 59 77 59 3 D
rlabel ndiffusion 79 13 79 13 3 #5
rlabel pdiffusion 79 39 79 39 3 #7
rlabel pdiffusion 79 56 79 56 3 #7
rlabel pdiffusion 79 58 79 58 3 #7
rlabel pdiffusion 73 49 73 49 3 Vdd
rlabel ntransistor 77 13 77 13 3 D
rlabel ptransistor 77 39 77 39 3 D
rlabel polysilicon 68 52 68 52 3 Q
rlabel ndiffusion 69 13 69 13 3 GND
rlabel ndiffusion 61 20 61 20 3 #10
rlabel pdiffusion 69 39 69 39 3 Vdd
rlabel polysilicon 67 49 67 49 3 Q
rlabel ntransistor 67 13 67 13 3 Q
rlabel polysilicon 67 23 67 23 3 Q
rlabel ptransistor 67 39 67 39 3 Q
rlabel polysilicon 65 51 65 51 3 Q
rlabel polysilicon 65 54 65 54 3 Q
rlabel polysilicon 77 10 77 10 3 D
rlabel ndiffusion 61 13 61 13 3 #10
rlabel ndiffusion 61 22 61 22 3 #10
rlabel pdiffusion 61 39 61 39 3 #8
rlabel polysilicon 49 23 49 23 3 _clk
rlabel polysilicon 49 32 49 32 3 _clk
rlabel polysilicon 49 59 49 59 3 _clk
rlabel pdiffusion 51 39 51 39 3 #7
rlabel pdiffusion 51 56 51 56 3 #7
rlabel pdiffusion 51 58 51 58 3 #7
rlabel pdiffusion 45 49 45 49 3 _q
rlabel polysilicon 67 10 67 10 3 Q
rlabel ndiffusion 51 13 51 13 3 #10
rlabel ndiffusion 51 20 51 20 3 #10
rlabel ndiffusion 51 22 51 22 3 #10
rlabel ptransistor 49 39 49 39 3 _clk
rlabel ntransistor 49 13 49 13 3 _clk
rlabel pdiffusion 41 39 41 39 3 _q
rlabel pdiffusion 41 40 41 40 3 _q
rlabel pdiffusion 41 42 41 42 3 _q
rlabel polysilicon 39 49 39 49 3 CLK
rlabel polysilicon 49 10 49 10 3 _clk
rlabel ndiffusion 41 13 41 13 3 _q
rlabel ndiffusion 41 14 41 14 3 _q
rlabel ndiffusion 41 16 41 16 3 _q
rlabel ndiffusion 33 20 33 20 3 #5
rlabel polysilicon 39 23 39 23 3 CLK
rlabel ptransistor 39 39 39 39 3 CLK
rlabel ntransistor 39 13 39 13 3 CLK
rlabel ndiffusion 33 22 33 22 3 #5
rlabel pdiffusion 33 39 33 39 3 #8
rlabel pdiffusion 33 40 33 40 3 #8
rlabel pdiffusion 33 42 33 42 3 #8
rlabel polysilicon 39 10 39 10 3 CLK
rlabel ndiffusion 33 13 33 13 3 #5
rlabel polysilicon 21 10 21 10 3 CLK
rlabel ndiffusion 23 13 23 13 3 _clk
rlabel ndiffusion 23 20 23 20 3 _clk
rlabel ndiffusion 23 22 23 22 3 _clk
rlabel pdiffusion 23 39 23 39 3 _clk
rlabel pdiffusion 23 40 23 40 3 _clk
rlabel pdiffusion 23 42 23 42 3 _clk
rlabel ntransistor 21 13 21 13 3 CLK
rlabel polysilicon 21 23 21 23 3 CLK
rlabel ptransistor 21 39 21 39 3 CLK
rlabel polysilicon 21 54 21 54 3 CLK
rlabel polysilicon 21 56 21 56 3 CLK
rlabel polysilicon 13 7 13 7 3 _q
rlabel ndiffusion 15 13 15 13 3 GND
rlabel ndiffusion 15 14 15 14 3 GND
rlabel ndiffusion 15 16 15 16 3 GND
rlabel pdiffusion 15 39 15 39 3 Vdd
rlabel pdiffusion 15 51 15 51 3 Vdd
rlabel pdiffusion 15 53 15 53 3 Vdd
rlabel ntransistor 13 13 13 13 3 _q
rlabel polysilicon 13 23 13 23 3 _q
rlabel ptransistor 13 39 13 39 3 _q
rlabel polysilicon 13 54 13 54 3 _q
rlabel ndiffusion 7 13 7 13 3 Q
rlabel pdiffusion 7 39 7 39 3 Q
rlabel pdiffusion 7 51 7 51 3 Q
rlabel m1 83 56 83 56 3 #7
rlabel pdcontact 81 56 81 56 3 #7
rlabel m1 80 56 80 56 3 #7
rlabel m1 80 55 80 55 3 #7
rlabel m1 76 56 76 56 3 Vdd
rlabel m1 80 58 80 58 3 #7
rlabel m1 78 20 78 20 3 #5
rlabel m1 78 23 78 23 3 #5
rlabel m1 79 32 79 32 3 D
port 2 e default input
rlabel pdcontact 74 56 74 56 3 Vdd
rlabel polycontact 77 32 77 32 3 D
port 2 e
rlabel m1 73 55 73 55 3 Vdd
rlabel m1 73 56 73 56 3 Vdd
rlabel m1 73 58 73 58 3 Vdd
rlabel m1 56 56 56 56 3 #7
rlabel m1 76 31 76 31 3 D
port 2 e
rlabel m1 76 32 76 32 3 D
port 2 e
rlabel m1 76 34 76 34 3 D
port 2 e
rlabel m1 80 59 80 59 3 #7
rlabel pdcontact 54 56 54 56 3 #7
rlabel m1 54 59 54 59 3 #7
rlabel m1 54 67 54 67 3 #7
rlabel m1 46 40 46 40 3 _q
rlabel m1 53 55 53 55 3 #7
rlabel m1 53 56 53 56 3 #7
rlabel m1 53 58 53 58 3 #7
rlabel m1 72 59 72 59 3 Vdd
rlabel m1 72 60 72 60 3 Vdd
rlabel m1 72 63 72 63 3 Vdd
rlabel pdcontact 44 40 44 40 3 _q
rlabel m1 66 53 66 53 3 Q
port 3 e default output
rlabel m1 43 40 43 40 3 _q
rlabel m1 43 42 43 42 3 _q
rlabel m1 64 49 64 49 3 Q
port 3 e default output
rlabel m1 64 50 64 50 3 Q
port 3 e default output
rlabel m1 64 53 64 53 3 Q
port 3 e default output
rlabel m1 64 54 64 54 3 Q
port 3 e default output
rlabel m1 64 20 64 20 3 #10
rlabel m1 72 14 72 14 3 GND
rlabel m1 78 19 78 19 3 #5
rlabel ndcontact 62 20 62 20 3 #10
rlabel m1 60 39 60 39 3 #8
rlabel m1 60 40 60 40 3 #8
rlabel m1 60 43 60 43 3 #8
rlabel m1 43 39 43 39 3 _q
rlabel ndcontact 70 14 70 14 3 GND
rlabel m1 56 20 56 20 3 #10
rlabel m1 69 14 69 14 3 GND
rlabel m1 69 16 69 16 3 GND
rlabel ndcontact 54 20 54 20 3 #10
rlabel m1 53 20 53 20 3 #10
rlabel m1 53 22 53 22 3 #10
rlabel m1 46 14 46 14 3 _q
rlabel m1 53 19 53 19 3 #10
rlabel m1 49 29 49 29 3 _clk
rlabel m1 49 30 49 30 3 _clk
rlabel m1 49 33 49 33 3 _clk
rlabel m1 34 56 34 56 3 CLK
port 1 e default input
rlabel ndcontact 44 14 44 14 3 _q
rlabel polycontact 32 56 32 56 3 CLK
port 1 e default input
rlabel m1 68 9 68 9 3 GND
rlabel m1 68 10 68 10 3 GND
rlabel m1 43 14 43 14 3 _q
rlabel m1 43 16 43 16 3 _q
rlabel m1 43 17 43 17 3 _q
rlabel m1 28 20 28 20 3 _clk
rlabel m1 28 40 28 40 3 _clk
rlabel m1 31 55 31 55 3 CLK
port 1 e default input
rlabel m1 31 56 31 56 3 CLK
port 1 e default input
rlabel m1 31 58 31 58 3 CLK
port 1 e default input
rlabel m1 31 59 31 59 3 CLK
port 1 e
rlabel m1 68 13 68 13 3 GND
rlabel ndcontact 26 20 26 20 3 _clk
rlabel m1 26 23 26 23 3 _clk
rlabel m1 26 34 26 34 3 _clk
rlabel pdcontact 26 40 26 40 3 _clk
rlabel m1 43 6 43 6 3 _q
rlabel m1 25 20 25 20 3 _clk
rlabel m1 25 22 25 22 3 _clk
rlabel m1 25 39 25 39 3 _clk
rlabel m1 25 40 25 40 3 _clk
rlabel m1 25 42 25 42 3 _clk
rlabel m1 20 51 20 51 3 Vdd
rlabel m1 43 13 43 13 3 _q
rlabel m1 20 14 20 14 3 GND
rlabel m1 25 19 25 19 3 _clk
rlabel pdcontact 18 51 18 51 3 Vdd
rlabel ndcontact 18 14 18 14 3 GND
rlabel m1 17 50 17 50 3 Vdd
rlabel m1 17 51 17 51 3 Vdd
rlabel m1 17 53 17 53 3 Vdd
rlabel m1 17 54 17 54 3 Vdd
rlabel m1 13 4 13 4 3 _q
rlabel m1 17 14 17 14 3 GND
rlabel m1 17 16 17 16 3 GND
rlabel polycontact 11 4 11 4 3 _q
rlabel m1 10 3 10 3 3 _q
rlabel m1 10 4 10 4 3 _q
rlabel m1 10 6 10 6 3 _q
rlabel m1 10 20 10 20 3 Q
port 3 e default output
rlabel ndcontact 8 20 8 20 3 Q
port 3 e default output
rlabel m1 7 19 7 19 3 Q
port 3 e default output
rlabel m1 7 20 7 20 3 Q
port 3 e default output
rlabel m1 7 22 7 22 3 Q
port 3 e default output
rlabel m1 7 23 7 23 3 Q
port 3 e default output
rlabel m1 7 54 7 54 3 Q
port 3 e default output
rlabel m2 64 40 64 40 3 #8
rlabel m2 82 20 82 20 3 #5
rlabel m2c 62 40 62 40 3 #8
rlabel m2c 80 20 80 20 3 #5
rlabel m2c 61 40 61 40 3 #8
rlabel m2 61 42 61 42 3 #8
rlabel m2c 79 20 79 20 3 #5
rlabel m2 79 22 79 22 3 #5
rlabel m2 39 40 39 40 3 #8
rlabel m2 39 20 39 20 3 #5
rlabel m2 53 30 53 30 3 _clk
rlabel m2 38 40 38 40 3 #8
rlabel m2 38 20 38 20 3 #5
rlabel m2 52 30 52 30 3 _clk
rlabel m2c 36 40 36 40 3 #8
rlabel m2 36 42 36 42 3 #8
rlabel m2c 36 20 36 20 3 #5
rlabel m2 36 22 36 22 3 #5
rlabel m2c 50 30 50 30 3 _clk
rlabel m2 50 32 50 32 3 _clk
rlabel m2 35 39 35 39 3 #8
rlabel m2 35 40 35 40 3 #8
rlabel m2 35 43 35 43 3 #8
rlabel m2 35 19 35 19 3 #5
rlabel m2 35 20 35 20 3 #5
rlabel m2 35 23 35 23 3 #5
rlabel m2 30 30 30 30 3 _clk
rlabel m2 76 60 76 60 3 Vdd
rlabel m2 72 10 72 10 3 GND
rlabel m2c 27 30 27 30 3 _clk
rlabel m2c 73 60 73 60 3 Vdd
rlabel m2c 69 10 69 10 3 GND
rlabel m2 26 29 26 29 3 _clk
rlabel m2 26 30 26 30 3 _clk
rlabel m2 26 33 26 33 3 _clk
rlabel m2 19 60 19 60 3 Vdd
rlabel m2 21 10 21 10 3 GND
rlabel m2c 16 60 16 60 3 Vdd
rlabel m2c 18 10 18 10 3 GND
rlabel m2 68 50 68 50 3 Q
port 3 e default output
rlabel m2 66 52 66 52 3 Q
port 3 e default output
rlabel m2 15 59 15 59 3 Vdd
rlabel m2 15 60 15 60 3 Vdd
rlabel m2 15 63 15 63 3 Vdd
rlabel m2 17 9 17 9 3 GND
rlabel m2 17 10 17 10 3 GND
rlabel m2 17 13 17 13 3 GND
rlabel m2c 65 50 65 50 3 Q
port 3 e default output
rlabel m2 65 52 65 52 3 Q
port 3 e default output
rlabel m2 11 50 11 50 3 Q
port 3 e
rlabel m2 10 51 10 51 3 Q
port 3 e
rlabel m2c 8 50 8 50 3 Q
port 3 e
rlabel m2c 8 51 8 51 3 Q
port 3 e
rlabel m2 7 49 7 49 3 Q
port 3 e
rlabel m2 7 50 7 50 3 Q
port 3 e
rlabel m2 7 53 7 53 3 Q
port 3 e
<< properties >>
string FIXED_BBOX 0 0 96 80
string LEFclass CORE
string LEFsite CoreSite
string LEFsymmetry X Y
string LEFview TRUE
<< end >>
