magic
tech sky130l
timestamp 1731220340
<< m2 >>
rect 110 4004 116 4005
rect 2006 4004 2012 4005
rect 110 4000 111 4004
rect 115 4000 116 4004
rect 110 3999 116 4000
rect 1518 4003 1524 4004
rect 1518 3999 1519 4003
rect 1523 3999 1524 4003
rect 1518 3998 1524 3999
rect 1614 4003 1620 4004
rect 1614 3999 1615 4003
rect 1619 3999 1620 4003
rect 1614 3998 1620 3999
rect 1710 4003 1716 4004
rect 1710 3999 1711 4003
rect 1715 3999 1716 4003
rect 1710 3998 1716 3999
rect 1806 4003 1812 4004
rect 1806 3999 1807 4003
rect 1811 3999 1812 4003
rect 1806 3998 1812 3999
rect 1902 4003 1908 4004
rect 1902 3999 1903 4003
rect 1907 3999 1908 4003
rect 2006 4000 2007 4004
rect 2011 4000 2012 4004
rect 2006 3999 2012 4000
rect 1902 3998 1908 3999
rect 2070 3988 2076 3989
rect 110 3987 116 3988
rect 110 3983 111 3987
rect 115 3983 116 3987
rect 2006 3987 2012 3988
rect 110 3982 116 3983
rect 1518 3984 1524 3985
rect 1518 3980 1519 3984
rect 1523 3980 1524 3984
rect 1518 3979 1524 3980
rect 1614 3984 1620 3985
rect 1614 3980 1615 3984
rect 1619 3980 1620 3984
rect 1614 3979 1620 3980
rect 1710 3984 1716 3985
rect 1710 3980 1711 3984
rect 1715 3980 1716 3984
rect 1710 3979 1716 3980
rect 1806 3984 1812 3985
rect 1806 3980 1807 3984
rect 1811 3980 1812 3984
rect 1806 3979 1812 3980
rect 1902 3984 1908 3985
rect 1902 3980 1903 3984
rect 1907 3980 1908 3984
rect 2006 3983 2007 3987
rect 2011 3983 2012 3987
rect 2006 3982 2012 3983
rect 2046 3985 2052 3986
rect 2046 3981 2047 3985
rect 2051 3981 2052 3985
rect 2070 3984 2071 3988
rect 2075 3984 2076 3988
rect 2070 3983 2076 3984
rect 2166 3988 2172 3989
rect 2166 3984 2167 3988
rect 2171 3984 2172 3988
rect 2166 3983 2172 3984
rect 2262 3988 2268 3989
rect 2262 3984 2263 3988
rect 2267 3984 2268 3988
rect 2262 3983 2268 3984
rect 3942 3985 3948 3986
rect 2046 3980 2052 3981
rect 3942 3981 3943 3985
rect 3947 3981 3948 3985
rect 3942 3980 3948 3981
rect 1902 3979 1908 3980
rect 2070 3969 2076 3970
rect 2046 3968 2052 3969
rect 2046 3964 2047 3968
rect 2051 3964 2052 3968
rect 2070 3965 2071 3969
rect 2075 3965 2076 3969
rect 2070 3964 2076 3965
rect 2166 3969 2172 3970
rect 2166 3965 2167 3969
rect 2171 3965 2172 3969
rect 2166 3964 2172 3965
rect 2262 3969 2268 3970
rect 2262 3965 2263 3969
rect 2267 3965 2268 3969
rect 2262 3964 2268 3965
rect 3942 3968 3948 3969
rect 3942 3964 3943 3968
rect 3947 3964 3948 3968
rect 2046 3963 2052 3964
rect 3942 3963 3948 3964
rect 198 3924 204 3925
rect 110 3921 116 3922
rect 110 3917 111 3921
rect 115 3917 116 3921
rect 198 3920 199 3924
rect 203 3920 204 3924
rect 198 3919 204 3920
rect 294 3924 300 3925
rect 294 3920 295 3924
rect 299 3920 300 3924
rect 294 3919 300 3920
rect 390 3924 396 3925
rect 390 3920 391 3924
rect 395 3920 396 3924
rect 390 3919 396 3920
rect 494 3924 500 3925
rect 494 3920 495 3924
rect 499 3920 500 3924
rect 494 3919 500 3920
rect 614 3924 620 3925
rect 614 3920 615 3924
rect 619 3920 620 3924
rect 614 3919 620 3920
rect 742 3924 748 3925
rect 742 3920 743 3924
rect 747 3920 748 3924
rect 742 3919 748 3920
rect 870 3924 876 3925
rect 870 3920 871 3924
rect 875 3920 876 3924
rect 870 3919 876 3920
rect 998 3924 1004 3925
rect 998 3920 999 3924
rect 1003 3920 1004 3924
rect 998 3919 1004 3920
rect 1126 3924 1132 3925
rect 1126 3920 1127 3924
rect 1131 3920 1132 3924
rect 1126 3919 1132 3920
rect 1254 3924 1260 3925
rect 1254 3920 1255 3924
rect 1259 3920 1260 3924
rect 1254 3919 1260 3920
rect 1382 3924 1388 3925
rect 1382 3920 1383 3924
rect 1387 3920 1388 3924
rect 1382 3919 1388 3920
rect 1510 3924 1516 3925
rect 1510 3920 1511 3924
rect 1515 3920 1516 3924
rect 1510 3919 1516 3920
rect 1646 3924 1652 3925
rect 1646 3920 1647 3924
rect 1651 3920 1652 3924
rect 1646 3919 1652 3920
rect 2006 3921 2012 3922
rect 110 3916 116 3917
rect 2006 3917 2007 3921
rect 2011 3917 2012 3921
rect 2006 3916 2012 3917
rect 2046 3916 2052 3917
rect 3942 3916 3948 3917
rect 2046 3912 2047 3916
rect 2051 3912 2052 3916
rect 2046 3911 2052 3912
rect 2158 3915 2164 3916
rect 2158 3911 2159 3915
rect 2163 3911 2164 3915
rect 2158 3910 2164 3911
rect 2286 3915 2292 3916
rect 2286 3911 2287 3915
rect 2291 3911 2292 3915
rect 2286 3910 2292 3911
rect 2414 3915 2420 3916
rect 2414 3911 2415 3915
rect 2419 3911 2420 3915
rect 2414 3910 2420 3911
rect 2550 3915 2556 3916
rect 2550 3911 2551 3915
rect 2555 3911 2556 3915
rect 2550 3910 2556 3911
rect 2686 3915 2692 3916
rect 2686 3911 2687 3915
rect 2691 3911 2692 3915
rect 2686 3910 2692 3911
rect 2822 3915 2828 3916
rect 2822 3911 2823 3915
rect 2827 3911 2828 3915
rect 2822 3910 2828 3911
rect 2950 3915 2956 3916
rect 2950 3911 2951 3915
rect 2955 3911 2956 3915
rect 2950 3910 2956 3911
rect 3070 3915 3076 3916
rect 3070 3911 3071 3915
rect 3075 3911 3076 3915
rect 3070 3910 3076 3911
rect 3190 3915 3196 3916
rect 3190 3911 3191 3915
rect 3195 3911 3196 3915
rect 3190 3910 3196 3911
rect 3302 3915 3308 3916
rect 3302 3911 3303 3915
rect 3307 3911 3308 3915
rect 3302 3910 3308 3911
rect 3406 3915 3412 3916
rect 3406 3911 3407 3915
rect 3411 3911 3412 3915
rect 3406 3910 3412 3911
rect 3518 3915 3524 3916
rect 3518 3911 3519 3915
rect 3523 3911 3524 3915
rect 3518 3910 3524 3911
rect 3630 3915 3636 3916
rect 3630 3911 3631 3915
rect 3635 3911 3636 3915
rect 3630 3910 3636 3911
rect 3742 3915 3748 3916
rect 3742 3911 3743 3915
rect 3747 3911 3748 3915
rect 3942 3912 3943 3916
rect 3947 3912 3948 3916
rect 3942 3911 3948 3912
rect 3742 3910 3748 3911
rect 198 3905 204 3906
rect 110 3904 116 3905
rect 110 3900 111 3904
rect 115 3900 116 3904
rect 198 3901 199 3905
rect 203 3901 204 3905
rect 198 3900 204 3901
rect 294 3905 300 3906
rect 294 3901 295 3905
rect 299 3901 300 3905
rect 294 3900 300 3901
rect 390 3905 396 3906
rect 390 3901 391 3905
rect 395 3901 396 3905
rect 390 3900 396 3901
rect 494 3905 500 3906
rect 494 3901 495 3905
rect 499 3901 500 3905
rect 494 3900 500 3901
rect 614 3905 620 3906
rect 614 3901 615 3905
rect 619 3901 620 3905
rect 614 3900 620 3901
rect 742 3905 748 3906
rect 742 3901 743 3905
rect 747 3901 748 3905
rect 742 3900 748 3901
rect 870 3905 876 3906
rect 870 3901 871 3905
rect 875 3901 876 3905
rect 870 3900 876 3901
rect 998 3905 1004 3906
rect 998 3901 999 3905
rect 1003 3901 1004 3905
rect 998 3900 1004 3901
rect 1126 3905 1132 3906
rect 1126 3901 1127 3905
rect 1131 3901 1132 3905
rect 1126 3900 1132 3901
rect 1254 3905 1260 3906
rect 1254 3901 1255 3905
rect 1259 3901 1260 3905
rect 1254 3900 1260 3901
rect 1382 3905 1388 3906
rect 1382 3901 1383 3905
rect 1387 3901 1388 3905
rect 1382 3900 1388 3901
rect 1510 3905 1516 3906
rect 1510 3901 1511 3905
rect 1515 3901 1516 3905
rect 1510 3900 1516 3901
rect 1646 3905 1652 3906
rect 1646 3901 1647 3905
rect 1651 3901 1652 3905
rect 1646 3900 1652 3901
rect 2006 3904 2012 3905
rect 2006 3900 2007 3904
rect 2011 3900 2012 3904
rect 110 3899 116 3900
rect 2006 3899 2012 3900
rect 2046 3899 2052 3900
rect 2046 3895 2047 3899
rect 2051 3895 2052 3899
rect 3942 3899 3948 3900
rect 2046 3894 2052 3895
rect 2158 3896 2164 3897
rect 2158 3892 2159 3896
rect 2163 3892 2164 3896
rect 2158 3891 2164 3892
rect 2286 3896 2292 3897
rect 2286 3892 2287 3896
rect 2291 3892 2292 3896
rect 2286 3891 2292 3892
rect 2414 3896 2420 3897
rect 2414 3892 2415 3896
rect 2419 3892 2420 3896
rect 2414 3891 2420 3892
rect 2550 3896 2556 3897
rect 2550 3892 2551 3896
rect 2555 3892 2556 3896
rect 2550 3891 2556 3892
rect 2686 3896 2692 3897
rect 2686 3892 2687 3896
rect 2691 3892 2692 3896
rect 2686 3891 2692 3892
rect 2822 3896 2828 3897
rect 2822 3892 2823 3896
rect 2827 3892 2828 3896
rect 2822 3891 2828 3892
rect 2950 3896 2956 3897
rect 2950 3892 2951 3896
rect 2955 3892 2956 3896
rect 2950 3891 2956 3892
rect 3070 3896 3076 3897
rect 3070 3892 3071 3896
rect 3075 3892 3076 3896
rect 3070 3891 3076 3892
rect 3190 3896 3196 3897
rect 3190 3892 3191 3896
rect 3195 3892 3196 3896
rect 3190 3891 3196 3892
rect 3302 3896 3308 3897
rect 3302 3892 3303 3896
rect 3307 3892 3308 3896
rect 3302 3891 3308 3892
rect 3406 3896 3412 3897
rect 3406 3892 3407 3896
rect 3411 3892 3412 3896
rect 3406 3891 3412 3892
rect 3518 3896 3524 3897
rect 3518 3892 3519 3896
rect 3523 3892 3524 3896
rect 3518 3891 3524 3892
rect 3630 3896 3636 3897
rect 3630 3892 3631 3896
rect 3635 3892 3636 3896
rect 3630 3891 3636 3892
rect 3742 3896 3748 3897
rect 3742 3892 3743 3896
rect 3747 3892 3748 3896
rect 3942 3895 3943 3899
rect 3947 3895 3948 3899
rect 3942 3894 3948 3895
rect 3742 3891 3748 3892
rect 110 3852 116 3853
rect 2006 3852 2012 3853
rect 110 3848 111 3852
rect 115 3848 116 3852
rect 110 3847 116 3848
rect 334 3851 340 3852
rect 334 3847 335 3851
rect 339 3847 340 3851
rect 334 3846 340 3847
rect 454 3851 460 3852
rect 454 3847 455 3851
rect 459 3847 460 3851
rect 454 3846 460 3847
rect 582 3851 588 3852
rect 582 3847 583 3851
rect 587 3847 588 3851
rect 582 3846 588 3847
rect 718 3851 724 3852
rect 718 3847 719 3851
rect 723 3847 724 3851
rect 718 3846 724 3847
rect 846 3851 852 3852
rect 846 3847 847 3851
rect 851 3847 852 3851
rect 846 3846 852 3847
rect 974 3851 980 3852
rect 974 3847 975 3851
rect 979 3847 980 3851
rect 974 3846 980 3847
rect 1102 3851 1108 3852
rect 1102 3847 1103 3851
rect 1107 3847 1108 3851
rect 1102 3846 1108 3847
rect 1230 3851 1236 3852
rect 1230 3847 1231 3851
rect 1235 3847 1236 3851
rect 1230 3846 1236 3847
rect 1358 3851 1364 3852
rect 1358 3847 1359 3851
rect 1363 3847 1364 3851
rect 1358 3846 1364 3847
rect 1486 3851 1492 3852
rect 1486 3847 1487 3851
rect 1491 3847 1492 3851
rect 2006 3848 2007 3852
rect 2011 3848 2012 3852
rect 2006 3847 2012 3848
rect 1486 3846 1492 3847
rect 110 3835 116 3836
rect 110 3831 111 3835
rect 115 3831 116 3835
rect 2006 3835 2012 3836
rect 110 3830 116 3831
rect 334 3832 340 3833
rect 334 3828 335 3832
rect 339 3828 340 3832
rect 334 3827 340 3828
rect 454 3832 460 3833
rect 454 3828 455 3832
rect 459 3828 460 3832
rect 454 3827 460 3828
rect 582 3832 588 3833
rect 582 3828 583 3832
rect 587 3828 588 3832
rect 582 3827 588 3828
rect 718 3832 724 3833
rect 718 3828 719 3832
rect 723 3828 724 3832
rect 718 3827 724 3828
rect 846 3832 852 3833
rect 846 3828 847 3832
rect 851 3828 852 3832
rect 846 3827 852 3828
rect 974 3832 980 3833
rect 974 3828 975 3832
rect 979 3828 980 3832
rect 974 3827 980 3828
rect 1102 3832 1108 3833
rect 1102 3828 1103 3832
rect 1107 3828 1108 3832
rect 1102 3827 1108 3828
rect 1230 3832 1236 3833
rect 1230 3828 1231 3832
rect 1235 3828 1236 3832
rect 1230 3827 1236 3828
rect 1358 3832 1364 3833
rect 1358 3828 1359 3832
rect 1363 3828 1364 3832
rect 1358 3827 1364 3828
rect 1486 3832 1492 3833
rect 1486 3828 1487 3832
rect 1491 3828 1492 3832
rect 2006 3831 2007 3835
rect 2011 3831 2012 3835
rect 2006 3830 2012 3831
rect 1486 3827 1492 3828
rect 2206 3828 2212 3829
rect 2046 3825 2052 3826
rect 2046 3821 2047 3825
rect 2051 3821 2052 3825
rect 2206 3824 2207 3828
rect 2211 3824 2212 3828
rect 2206 3823 2212 3824
rect 2342 3828 2348 3829
rect 2342 3824 2343 3828
rect 2347 3824 2348 3828
rect 2342 3823 2348 3824
rect 2486 3828 2492 3829
rect 2486 3824 2487 3828
rect 2491 3824 2492 3828
rect 2486 3823 2492 3824
rect 2646 3828 2652 3829
rect 2646 3824 2647 3828
rect 2651 3824 2652 3828
rect 2646 3823 2652 3824
rect 2822 3828 2828 3829
rect 2822 3824 2823 3828
rect 2827 3824 2828 3828
rect 2822 3823 2828 3824
rect 3014 3828 3020 3829
rect 3014 3824 3015 3828
rect 3019 3824 3020 3828
rect 3014 3823 3020 3824
rect 3222 3828 3228 3829
rect 3222 3824 3223 3828
rect 3227 3824 3228 3828
rect 3222 3823 3228 3824
rect 3438 3828 3444 3829
rect 3438 3824 3439 3828
rect 3443 3824 3444 3828
rect 3438 3823 3444 3824
rect 3654 3828 3660 3829
rect 3654 3824 3655 3828
rect 3659 3824 3660 3828
rect 3654 3823 3660 3824
rect 3942 3825 3948 3826
rect 2046 3820 2052 3821
rect 3942 3821 3943 3825
rect 3947 3821 3948 3825
rect 3942 3820 3948 3821
rect 2206 3809 2212 3810
rect 2046 3808 2052 3809
rect 2046 3804 2047 3808
rect 2051 3804 2052 3808
rect 2206 3805 2207 3809
rect 2211 3805 2212 3809
rect 2206 3804 2212 3805
rect 2342 3809 2348 3810
rect 2342 3805 2343 3809
rect 2347 3805 2348 3809
rect 2342 3804 2348 3805
rect 2486 3809 2492 3810
rect 2486 3805 2487 3809
rect 2491 3805 2492 3809
rect 2486 3804 2492 3805
rect 2646 3809 2652 3810
rect 2646 3805 2647 3809
rect 2651 3805 2652 3809
rect 2646 3804 2652 3805
rect 2822 3809 2828 3810
rect 2822 3805 2823 3809
rect 2827 3805 2828 3809
rect 2822 3804 2828 3805
rect 3014 3809 3020 3810
rect 3014 3805 3015 3809
rect 3019 3805 3020 3809
rect 3014 3804 3020 3805
rect 3222 3809 3228 3810
rect 3222 3805 3223 3809
rect 3227 3805 3228 3809
rect 3222 3804 3228 3805
rect 3438 3809 3444 3810
rect 3438 3805 3439 3809
rect 3443 3805 3444 3809
rect 3438 3804 3444 3805
rect 3654 3809 3660 3810
rect 3654 3805 3655 3809
rect 3659 3805 3660 3809
rect 3654 3804 3660 3805
rect 3942 3808 3948 3809
rect 3942 3804 3943 3808
rect 3947 3804 3948 3808
rect 2046 3803 2052 3804
rect 3942 3803 3948 3804
rect 502 3768 508 3769
rect 110 3765 116 3766
rect 110 3761 111 3765
rect 115 3761 116 3765
rect 502 3764 503 3768
rect 507 3764 508 3768
rect 502 3763 508 3764
rect 614 3768 620 3769
rect 614 3764 615 3768
rect 619 3764 620 3768
rect 614 3763 620 3764
rect 734 3768 740 3769
rect 734 3764 735 3768
rect 739 3764 740 3768
rect 734 3763 740 3764
rect 862 3768 868 3769
rect 862 3764 863 3768
rect 867 3764 868 3768
rect 862 3763 868 3764
rect 998 3768 1004 3769
rect 998 3764 999 3768
rect 1003 3764 1004 3768
rect 998 3763 1004 3764
rect 1142 3768 1148 3769
rect 1142 3764 1143 3768
rect 1147 3764 1148 3768
rect 1142 3763 1148 3764
rect 1286 3768 1292 3769
rect 1286 3764 1287 3768
rect 1291 3764 1292 3768
rect 1286 3763 1292 3764
rect 1430 3768 1436 3769
rect 1430 3764 1431 3768
rect 1435 3764 1436 3768
rect 1430 3763 1436 3764
rect 1582 3768 1588 3769
rect 1582 3764 1583 3768
rect 1587 3764 1588 3768
rect 1582 3763 1588 3764
rect 2006 3765 2012 3766
rect 110 3760 116 3761
rect 2006 3761 2007 3765
rect 2011 3761 2012 3765
rect 2006 3760 2012 3761
rect 2046 3756 2052 3757
rect 3942 3756 3948 3757
rect 2046 3752 2047 3756
rect 2051 3752 2052 3756
rect 2046 3751 2052 3752
rect 2190 3755 2196 3756
rect 2190 3751 2191 3755
rect 2195 3751 2196 3755
rect 2190 3750 2196 3751
rect 2374 3755 2380 3756
rect 2374 3751 2375 3755
rect 2379 3751 2380 3755
rect 2374 3750 2380 3751
rect 2558 3755 2564 3756
rect 2558 3751 2559 3755
rect 2563 3751 2564 3755
rect 2558 3750 2564 3751
rect 2742 3755 2748 3756
rect 2742 3751 2743 3755
rect 2747 3751 2748 3755
rect 2742 3750 2748 3751
rect 2934 3755 2940 3756
rect 2934 3751 2935 3755
rect 2939 3751 2940 3755
rect 2934 3750 2940 3751
rect 3126 3755 3132 3756
rect 3126 3751 3127 3755
rect 3131 3751 3132 3755
rect 3126 3750 3132 3751
rect 3318 3755 3324 3756
rect 3318 3751 3319 3755
rect 3323 3751 3324 3755
rect 3318 3750 3324 3751
rect 3510 3755 3516 3756
rect 3510 3751 3511 3755
rect 3515 3751 3516 3755
rect 3510 3750 3516 3751
rect 3710 3755 3716 3756
rect 3710 3751 3711 3755
rect 3715 3751 3716 3755
rect 3942 3752 3943 3756
rect 3947 3752 3948 3756
rect 3942 3751 3948 3752
rect 3710 3750 3716 3751
rect 502 3749 508 3750
rect 110 3748 116 3749
rect 110 3744 111 3748
rect 115 3744 116 3748
rect 502 3745 503 3749
rect 507 3745 508 3749
rect 502 3744 508 3745
rect 614 3749 620 3750
rect 614 3745 615 3749
rect 619 3745 620 3749
rect 614 3744 620 3745
rect 734 3749 740 3750
rect 734 3745 735 3749
rect 739 3745 740 3749
rect 734 3744 740 3745
rect 862 3749 868 3750
rect 862 3745 863 3749
rect 867 3745 868 3749
rect 862 3744 868 3745
rect 998 3749 1004 3750
rect 998 3745 999 3749
rect 1003 3745 1004 3749
rect 998 3744 1004 3745
rect 1142 3749 1148 3750
rect 1142 3745 1143 3749
rect 1147 3745 1148 3749
rect 1142 3744 1148 3745
rect 1286 3749 1292 3750
rect 1286 3745 1287 3749
rect 1291 3745 1292 3749
rect 1286 3744 1292 3745
rect 1430 3749 1436 3750
rect 1430 3745 1431 3749
rect 1435 3745 1436 3749
rect 1430 3744 1436 3745
rect 1582 3749 1588 3750
rect 1582 3745 1583 3749
rect 1587 3745 1588 3749
rect 1582 3744 1588 3745
rect 2006 3748 2012 3749
rect 2006 3744 2007 3748
rect 2011 3744 2012 3748
rect 110 3743 116 3744
rect 2006 3743 2012 3744
rect 2046 3739 2052 3740
rect 2046 3735 2047 3739
rect 2051 3735 2052 3739
rect 3942 3739 3948 3740
rect 2046 3734 2052 3735
rect 2190 3736 2196 3737
rect 2190 3732 2191 3736
rect 2195 3732 2196 3736
rect 2190 3731 2196 3732
rect 2374 3736 2380 3737
rect 2374 3732 2375 3736
rect 2379 3732 2380 3736
rect 2374 3731 2380 3732
rect 2558 3736 2564 3737
rect 2558 3732 2559 3736
rect 2563 3732 2564 3736
rect 2558 3731 2564 3732
rect 2742 3736 2748 3737
rect 2742 3732 2743 3736
rect 2747 3732 2748 3736
rect 2742 3731 2748 3732
rect 2934 3736 2940 3737
rect 2934 3732 2935 3736
rect 2939 3732 2940 3736
rect 2934 3731 2940 3732
rect 3126 3736 3132 3737
rect 3126 3732 3127 3736
rect 3131 3732 3132 3736
rect 3126 3731 3132 3732
rect 3318 3736 3324 3737
rect 3318 3732 3319 3736
rect 3323 3732 3324 3736
rect 3318 3731 3324 3732
rect 3510 3736 3516 3737
rect 3510 3732 3511 3736
rect 3515 3732 3516 3736
rect 3510 3731 3516 3732
rect 3710 3736 3716 3737
rect 3710 3732 3711 3736
rect 3715 3732 3716 3736
rect 3942 3735 3943 3739
rect 3947 3735 3948 3739
rect 3942 3734 3948 3735
rect 3710 3731 3716 3732
rect 110 3688 116 3689
rect 2006 3688 2012 3689
rect 110 3684 111 3688
rect 115 3684 116 3688
rect 110 3683 116 3684
rect 494 3687 500 3688
rect 494 3683 495 3687
rect 499 3683 500 3687
rect 494 3682 500 3683
rect 590 3687 596 3688
rect 590 3683 591 3687
rect 595 3683 596 3687
rect 590 3682 596 3683
rect 686 3687 692 3688
rect 686 3683 687 3687
rect 691 3683 692 3687
rect 686 3682 692 3683
rect 790 3687 796 3688
rect 790 3683 791 3687
rect 795 3683 796 3687
rect 790 3682 796 3683
rect 910 3687 916 3688
rect 910 3683 911 3687
rect 915 3683 916 3687
rect 910 3682 916 3683
rect 1038 3687 1044 3688
rect 1038 3683 1039 3687
rect 1043 3683 1044 3687
rect 1038 3682 1044 3683
rect 1182 3687 1188 3688
rect 1182 3683 1183 3687
rect 1187 3683 1188 3687
rect 1182 3682 1188 3683
rect 1334 3687 1340 3688
rect 1334 3683 1335 3687
rect 1339 3683 1340 3687
rect 1334 3682 1340 3683
rect 1494 3687 1500 3688
rect 1494 3683 1495 3687
rect 1499 3683 1500 3687
rect 1494 3682 1500 3683
rect 1654 3687 1660 3688
rect 1654 3683 1655 3687
rect 1659 3683 1660 3687
rect 2006 3684 2007 3688
rect 2011 3684 2012 3688
rect 2006 3683 2012 3684
rect 1654 3682 1660 3683
rect 2126 3672 2132 3673
rect 110 3671 116 3672
rect 110 3667 111 3671
rect 115 3667 116 3671
rect 2006 3671 2012 3672
rect 110 3666 116 3667
rect 494 3668 500 3669
rect 494 3664 495 3668
rect 499 3664 500 3668
rect 494 3663 500 3664
rect 590 3668 596 3669
rect 590 3664 591 3668
rect 595 3664 596 3668
rect 590 3663 596 3664
rect 686 3668 692 3669
rect 686 3664 687 3668
rect 691 3664 692 3668
rect 686 3663 692 3664
rect 790 3668 796 3669
rect 790 3664 791 3668
rect 795 3664 796 3668
rect 790 3663 796 3664
rect 910 3668 916 3669
rect 910 3664 911 3668
rect 915 3664 916 3668
rect 910 3663 916 3664
rect 1038 3668 1044 3669
rect 1038 3664 1039 3668
rect 1043 3664 1044 3668
rect 1038 3663 1044 3664
rect 1182 3668 1188 3669
rect 1182 3664 1183 3668
rect 1187 3664 1188 3668
rect 1182 3663 1188 3664
rect 1334 3668 1340 3669
rect 1334 3664 1335 3668
rect 1339 3664 1340 3668
rect 1334 3663 1340 3664
rect 1494 3668 1500 3669
rect 1494 3664 1495 3668
rect 1499 3664 1500 3668
rect 1494 3663 1500 3664
rect 1654 3668 1660 3669
rect 1654 3664 1655 3668
rect 1659 3664 1660 3668
rect 2006 3667 2007 3671
rect 2011 3667 2012 3671
rect 2006 3666 2012 3667
rect 2046 3669 2052 3670
rect 2046 3665 2047 3669
rect 2051 3665 2052 3669
rect 2126 3668 2127 3672
rect 2131 3668 2132 3672
rect 2126 3667 2132 3668
rect 2350 3672 2356 3673
rect 2350 3668 2351 3672
rect 2355 3668 2356 3672
rect 2350 3667 2356 3668
rect 2582 3672 2588 3673
rect 2582 3668 2583 3672
rect 2587 3668 2588 3672
rect 2582 3667 2588 3668
rect 2814 3672 2820 3673
rect 2814 3668 2815 3672
rect 2819 3668 2820 3672
rect 2814 3667 2820 3668
rect 3046 3672 3052 3673
rect 3046 3668 3047 3672
rect 3051 3668 3052 3672
rect 3046 3667 3052 3668
rect 3278 3672 3284 3673
rect 3278 3668 3279 3672
rect 3283 3668 3284 3672
rect 3278 3667 3284 3668
rect 3510 3672 3516 3673
rect 3510 3668 3511 3672
rect 3515 3668 3516 3672
rect 3510 3667 3516 3668
rect 3750 3672 3756 3673
rect 3750 3668 3751 3672
rect 3755 3668 3756 3672
rect 3750 3667 3756 3668
rect 3942 3669 3948 3670
rect 2046 3664 2052 3665
rect 3942 3665 3943 3669
rect 3947 3665 3948 3669
rect 3942 3664 3948 3665
rect 1654 3663 1660 3664
rect 2126 3653 2132 3654
rect 2046 3652 2052 3653
rect 2046 3648 2047 3652
rect 2051 3648 2052 3652
rect 2126 3649 2127 3653
rect 2131 3649 2132 3653
rect 2126 3648 2132 3649
rect 2350 3653 2356 3654
rect 2350 3649 2351 3653
rect 2355 3649 2356 3653
rect 2350 3648 2356 3649
rect 2582 3653 2588 3654
rect 2582 3649 2583 3653
rect 2587 3649 2588 3653
rect 2582 3648 2588 3649
rect 2814 3653 2820 3654
rect 2814 3649 2815 3653
rect 2819 3649 2820 3653
rect 2814 3648 2820 3649
rect 3046 3653 3052 3654
rect 3046 3649 3047 3653
rect 3051 3649 3052 3653
rect 3046 3648 3052 3649
rect 3278 3653 3284 3654
rect 3278 3649 3279 3653
rect 3283 3649 3284 3653
rect 3278 3648 3284 3649
rect 3510 3653 3516 3654
rect 3510 3649 3511 3653
rect 3515 3649 3516 3653
rect 3510 3648 3516 3649
rect 3750 3653 3756 3654
rect 3750 3649 3751 3653
rect 3755 3649 3756 3653
rect 3750 3648 3756 3649
rect 3942 3652 3948 3653
rect 3942 3648 3943 3652
rect 3947 3648 3948 3652
rect 2046 3647 2052 3648
rect 3942 3647 3948 3648
rect 334 3600 340 3601
rect 110 3597 116 3598
rect 110 3593 111 3597
rect 115 3593 116 3597
rect 334 3596 335 3600
rect 339 3596 340 3600
rect 334 3595 340 3596
rect 462 3600 468 3601
rect 462 3596 463 3600
rect 467 3596 468 3600
rect 462 3595 468 3596
rect 606 3600 612 3601
rect 606 3596 607 3600
rect 611 3596 612 3600
rect 606 3595 612 3596
rect 758 3600 764 3601
rect 758 3596 759 3600
rect 763 3596 764 3600
rect 758 3595 764 3596
rect 926 3600 932 3601
rect 926 3596 927 3600
rect 931 3596 932 3600
rect 926 3595 932 3596
rect 1094 3600 1100 3601
rect 1094 3596 1095 3600
rect 1099 3596 1100 3600
rect 1094 3595 1100 3596
rect 1262 3600 1268 3601
rect 1262 3596 1263 3600
rect 1267 3596 1268 3600
rect 1262 3595 1268 3596
rect 1438 3600 1444 3601
rect 1438 3596 1439 3600
rect 1443 3596 1444 3600
rect 1438 3595 1444 3596
rect 1614 3600 1620 3601
rect 1614 3596 1615 3600
rect 1619 3596 1620 3600
rect 1614 3595 1620 3596
rect 1790 3600 1796 3601
rect 1790 3596 1791 3600
rect 1795 3596 1796 3600
rect 1790 3595 1796 3596
rect 2006 3597 2012 3598
rect 110 3592 116 3593
rect 2006 3593 2007 3597
rect 2011 3593 2012 3597
rect 2006 3592 2012 3593
rect 2046 3592 2052 3593
rect 3942 3592 3948 3593
rect 2046 3588 2047 3592
rect 2051 3588 2052 3592
rect 2046 3587 2052 3588
rect 2190 3591 2196 3592
rect 2190 3587 2191 3591
rect 2195 3587 2196 3591
rect 2190 3586 2196 3587
rect 2326 3591 2332 3592
rect 2326 3587 2327 3591
rect 2331 3587 2332 3591
rect 2326 3586 2332 3587
rect 2454 3591 2460 3592
rect 2454 3587 2455 3591
rect 2459 3587 2460 3591
rect 2454 3586 2460 3587
rect 2582 3591 2588 3592
rect 2582 3587 2583 3591
rect 2587 3587 2588 3591
rect 2582 3586 2588 3587
rect 2718 3591 2724 3592
rect 2718 3587 2719 3591
rect 2723 3587 2724 3591
rect 2718 3586 2724 3587
rect 2854 3591 2860 3592
rect 2854 3587 2855 3591
rect 2859 3587 2860 3591
rect 2854 3586 2860 3587
rect 2998 3591 3004 3592
rect 2998 3587 2999 3591
rect 3003 3587 3004 3591
rect 2998 3586 3004 3587
rect 3142 3591 3148 3592
rect 3142 3587 3143 3591
rect 3147 3587 3148 3591
rect 3142 3586 3148 3587
rect 3294 3591 3300 3592
rect 3294 3587 3295 3591
rect 3299 3587 3300 3591
rect 3294 3586 3300 3587
rect 3454 3591 3460 3592
rect 3454 3587 3455 3591
rect 3459 3587 3460 3591
rect 3454 3586 3460 3587
rect 3622 3591 3628 3592
rect 3622 3587 3623 3591
rect 3627 3587 3628 3591
rect 3942 3588 3943 3592
rect 3947 3588 3948 3592
rect 3942 3587 3948 3588
rect 3622 3586 3628 3587
rect 334 3581 340 3582
rect 110 3580 116 3581
rect 110 3576 111 3580
rect 115 3576 116 3580
rect 334 3577 335 3581
rect 339 3577 340 3581
rect 334 3576 340 3577
rect 462 3581 468 3582
rect 462 3577 463 3581
rect 467 3577 468 3581
rect 462 3576 468 3577
rect 606 3581 612 3582
rect 606 3577 607 3581
rect 611 3577 612 3581
rect 606 3576 612 3577
rect 758 3581 764 3582
rect 758 3577 759 3581
rect 763 3577 764 3581
rect 758 3576 764 3577
rect 926 3581 932 3582
rect 926 3577 927 3581
rect 931 3577 932 3581
rect 926 3576 932 3577
rect 1094 3581 1100 3582
rect 1094 3577 1095 3581
rect 1099 3577 1100 3581
rect 1094 3576 1100 3577
rect 1262 3581 1268 3582
rect 1262 3577 1263 3581
rect 1267 3577 1268 3581
rect 1262 3576 1268 3577
rect 1438 3581 1444 3582
rect 1438 3577 1439 3581
rect 1443 3577 1444 3581
rect 1438 3576 1444 3577
rect 1614 3581 1620 3582
rect 1614 3577 1615 3581
rect 1619 3577 1620 3581
rect 1614 3576 1620 3577
rect 1790 3581 1796 3582
rect 1790 3577 1791 3581
rect 1795 3577 1796 3581
rect 1790 3576 1796 3577
rect 2006 3580 2012 3581
rect 2006 3576 2007 3580
rect 2011 3576 2012 3580
rect 110 3575 116 3576
rect 2006 3575 2012 3576
rect 2046 3575 2052 3576
rect 2046 3571 2047 3575
rect 2051 3571 2052 3575
rect 3942 3575 3948 3576
rect 2046 3570 2052 3571
rect 2190 3572 2196 3573
rect 2190 3568 2191 3572
rect 2195 3568 2196 3572
rect 2190 3567 2196 3568
rect 2326 3572 2332 3573
rect 2326 3568 2327 3572
rect 2331 3568 2332 3572
rect 2326 3567 2332 3568
rect 2454 3572 2460 3573
rect 2454 3568 2455 3572
rect 2459 3568 2460 3572
rect 2454 3567 2460 3568
rect 2582 3572 2588 3573
rect 2582 3568 2583 3572
rect 2587 3568 2588 3572
rect 2582 3567 2588 3568
rect 2718 3572 2724 3573
rect 2718 3568 2719 3572
rect 2723 3568 2724 3572
rect 2718 3567 2724 3568
rect 2854 3572 2860 3573
rect 2854 3568 2855 3572
rect 2859 3568 2860 3572
rect 2854 3567 2860 3568
rect 2998 3572 3004 3573
rect 2998 3568 2999 3572
rect 3003 3568 3004 3572
rect 2998 3567 3004 3568
rect 3142 3572 3148 3573
rect 3142 3568 3143 3572
rect 3147 3568 3148 3572
rect 3142 3567 3148 3568
rect 3294 3572 3300 3573
rect 3294 3568 3295 3572
rect 3299 3568 3300 3572
rect 3294 3567 3300 3568
rect 3454 3572 3460 3573
rect 3454 3568 3455 3572
rect 3459 3568 3460 3572
rect 3454 3567 3460 3568
rect 3622 3572 3628 3573
rect 3622 3568 3623 3572
rect 3627 3568 3628 3572
rect 3942 3571 3943 3575
rect 3947 3571 3948 3575
rect 3942 3570 3948 3571
rect 3622 3567 3628 3568
rect 110 3516 116 3517
rect 2006 3516 2012 3517
rect 110 3512 111 3516
rect 115 3512 116 3516
rect 110 3511 116 3512
rect 158 3515 164 3516
rect 158 3511 159 3515
rect 163 3511 164 3515
rect 158 3510 164 3511
rect 302 3515 308 3516
rect 302 3511 303 3515
rect 307 3511 308 3515
rect 302 3510 308 3511
rect 462 3515 468 3516
rect 462 3511 463 3515
rect 467 3511 468 3515
rect 462 3510 468 3511
rect 638 3515 644 3516
rect 638 3511 639 3515
rect 643 3511 644 3515
rect 638 3510 644 3511
rect 814 3515 820 3516
rect 814 3511 815 3515
rect 819 3511 820 3515
rect 814 3510 820 3511
rect 998 3515 1004 3516
rect 998 3511 999 3515
rect 1003 3511 1004 3515
rect 998 3510 1004 3511
rect 1174 3515 1180 3516
rect 1174 3511 1175 3515
rect 1179 3511 1180 3515
rect 1174 3510 1180 3511
rect 1350 3515 1356 3516
rect 1350 3511 1351 3515
rect 1355 3511 1356 3515
rect 1350 3510 1356 3511
rect 1526 3515 1532 3516
rect 1526 3511 1527 3515
rect 1531 3511 1532 3515
rect 1526 3510 1532 3511
rect 1702 3515 1708 3516
rect 1702 3511 1703 3515
rect 1707 3511 1708 3515
rect 1702 3510 1708 3511
rect 1878 3515 1884 3516
rect 1878 3511 1879 3515
rect 1883 3511 1884 3515
rect 2006 3512 2007 3516
rect 2011 3512 2012 3516
rect 2006 3511 2012 3512
rect 2102 3512 2108 3513
rect 1878 3510 1884 3511
rect 2046 3509 2052 3510
rect 2046 3505 2047 3509
rect 2051 3505 2052 3509
rect 2102 3508 2103 3512
rect 2107 3508 2108 3512
rect 2102 3507 2108 3508
rect 2270 3512 2276 3513
rect 2270 3508 2271 3512
rect 2275 3508 2276 3512
rect 2270 3507 2276 3508
rect 2446 3512 2452 3513
rect 2446 3508 2447 3512
rect 2451 3508 2452 3512
rect 2446 3507 2452 3508
rect 2630 3512 2636 3513
rect 2630 3508 2631 3512
rect 2635 3508 2636 3512
rect 2630 3507 2636 3508
rect 2814 3512 2820 3513
rect 2814 3508 2815 3512
rect 2819 3508 2820 3512
rect 2814 3507 2820 3508
rect 2998 3512 3004 3513
rect 2998 3508 2999 3512
rect 3003 3508 3004 3512
rect 2998 3507 3004 3508
rect 3174 3512 3180 3513
rect 3174 3508 3175 3512
rect 3179 3508 3180 3512
rect 3174 3507 3180 3508
rect 3350 3512 3356 3513
rect 3350 3508 3351 3512
rect 3355 3508 3356 3512
rect 3350 3507 3356 3508
rect 3518 3512 3524 3513
rect 3518 3508 3519 3512
rect 3523 3508 3524 3512
rect 3518 3507 3524 3508
rect 3686 3512 3692 3513
rect 3686 3508 3687 3512
rect 3691 3508 3692 3512
rect 3686 3507 3692 3508
rect 3838 3512 3844 3513
rect 3838 3508 3839 3512
rect 3843 3508 3844 3512
rect 3838 3507 3844 3508
rect 3942 3509 3948 3510
rect 2046 3504 2052 3505
rect 3942 3505 3943 3509
rect 3947 3505 3948 3509
rect 3942 3504 3948 3505
rect 110 3499 116 3500
rect 110 3495 111 3499
rect 115 3495 116 3499
rect 2006 3499 2012 3500
rect 110 3494 116 3495
rect 158 3496 164 3497
rect 158 3492 159 3496
rect 163 3492 164 3496
rect 158 3491 164 3492
rect 302 3496 308 3497
rect 302 3492 303 3496
rect 307 3492 308 3496
rect 302 3491 308 3492
rect 462 3496 468 3497
rect 462 3492 463 3496
rect 467 3492 468 3496
rect 462 3491 468 3492
rect 638 3496 644 3497
rect 638 3492 639 3496
rect 643 3492 644 3496
rect 638 3491 644 3492
rect 814 3496 820 3497
rect 814 3492 815 3496
rect 819 3492 820 3496
rect 814 3491 820 3492
rect 998 3496 1004 3497
rect 998 3492 999 3496
rect 1003 3492 1004 3496
rect 998 3491 1004 3492
rect 1174 3496 1180 3497
rect 1174 3492 1175 3496
rect 1179 3492 1180 3496
rect 1174 3491 1180 3492
rect 1350 3496 1356 3497
rect 1350 3492 1351 3496
rect 1355 3492 1356 3496
rect 1350 3491 1356 3492
rect 1526 3496 1532 3497
rect 1526 3492 1527 3496
rect 1531 3492 1532 3496
rect 1526 3491 1532 3492
rect 1702 3496 1708 3497
rect 1702 3492 1703 3496
rect 1707 3492 1708 3496
rect 1702 3491 1708 3492
rect 1878 3496 1884 3497
rect 1878 3492 1879 3496
rect 1883 3492 1884 3496
rect 2006 3495 2007 3499
rect 2011 3495 2012 3499
rect 2006 3494 2012 3495
rect 2102 3493 2108 3494
rect 1878 3491 1884 3492
rect 2046 3492 2052 3493
rect 2046 3488 2047 3492
rect 2051 3488 2052 3492
rect 2102 3489 2103 3493
rect 2107 3489 2108 3493
rect 2102 3488 2108 3489
rect 2270 3493 2276 3494
rect 2270 3489 2271 3493
rect 2275 3489 2276 3493
rect 2270 3488 2276 3489
rect 2446 3493 2452 3494
rect 2446 3489 2447 3493
rect 2451 3489 2452 3493
rect 2446 3488 2452 3489
rect 2630 3493 2636 3494
rect 2630 3489 2631 3493
rect 2635 3489 2636 3493
rect 2630 3488 2636 3489
rect 2814 3493 2820 3494
rect 2814 3489 2815 3493
rect 2819 3489 2820 3493
rect 2814 3488 2820 3489
rect 2998 3493 3004 3494
rect 2998 3489 2999 3493
rect 3003 3489 3004 3493
rect 2998 3488 3004 3489
rect 3174 3493 3180 3494
rect 3174 3489 3175 3493
rect 3179 3489 3180 3493
rect 3174 3488 3180 3489
rect 3350 3493 3356 3494
rect 3350 3489 3351 3493
rect 3355 3489 3356 3493
rect 3350 3488 3356 3489
rect 3518 3493 3524 3494
rect 3518 3489 3519 3493
rect 3523 3489 3524 3493
rect 3518 3488 3524 3489
rect 3686 3493 3692 3494
rect 3686 3489 3687 3493
rect 3691 3489 3692 3493
rect 3686 3488 3692 3489
rect 3838 3493 3844 3494
rect 3838 3489 3839 3493
rect 3843 3489 3844 3493
rect 3838 3488 3844 3489
rect 3942 3492 3948 3493
rect 3942 3488 3943 3492
rect 3947 3488 3948 3492
rect 2046 3487 2052 3488
rect 3942 3487 3948 3488
rect 2046 3436 2052 3437
rect 3942 3436 3948 3437
rect 2046 3432 2047 3436
rect 2051 3432 2052 3436
rect 2046 3431 2052 3432
rect 2126 3435 2132 3436
rect 2126 3431 2127 3435
rect 2131 3431 2132 3435
rect 2126 3430 2132 3431
rect 2310 3435 2316 3436
rect 2310 3431 2311 3435
rect 2315 3431 2316 3435
rect 2310 3430 2316 3431
rect 2494 3435 2500 3436
rect 2494 3431 2495 3435
rect 2499 3431 2500 3435
rect 2494 3430 2500 3431
rect 2678 3435 2684 3436
rect 2678 3431 2679 3435
rect 2683 3431 2684 3435
rect 2678 3430 2684 3431
rect 2862 3435 2868 3436
rect 2862 3431 2863 3435
rect 2867 3431 2868 3435
rect 2862 3430 2868 3431
rect 3046 3435 3052 3436
rect 3046 3431 3047 3435
rect 3051 3431 3052 3435
rect 3046 3430 3052 3431
rect 3222 3435 3228 3436
rect 3222 3431 3223 3435
rect 3227 3431 3228 3435
rect 3222 3430 3228 3431
rect 3406 3435 3412 3436
rect 3406 3431 3407 3435
rect 3411 3431 3412 3435
rect 3406 3430 3412 3431
rect 3590 3435 3596 3436
rect 3590 3431 3591 3435
rect 3595 3431 3596 3435
rect 3590 3430 3596 3431
rect 3774 3435 3780 3436
rect 3774 3431 3775 3435
rect 3779 3431 3780 3435
rect 3942 3432 3943 3436
rect 3947 3432 3948 3436
rect 3942 3431 3948 3432
rect 3774 3430 3780 3431
rect 134 3428 140 3429
rect 110 3425 116 3426
rect 110 3421 111 3425
rect 115 3421 116 3425
rect 134 3424 135 3428
rect 139 3424 140 3428
rect 134 3423 140 3424
rect 318 3428 324 3429
rect 318 3424 319 3428
rect 323 3424 324 3428
rect 318 3423 324 3424
rect 534 3428 540 3429
rect 534 3424 535 3428
rect 539 3424 540 3428
rect 534 3423 540 3424
rect 750 3428 756 3429
rect 750 3424 751 3428
rect 755 3424 756 3428
rect 750 3423 756 3424
rect 958 3428 964 3429
rect 958 3424 959 3428
rect 963 3424 964 3428
rect 958 3423 964 3424
rect 1158 3428 1164 3429
rect 1158 3424 1159 3428
rect 1163 3424 1164 3428
rect 1158 3423 1164 3424
rect 1350 3428 1356 3429
rect 1350 3424 1351 3428
rect 1355 3424 1356 3428
rect 1350 3423 1356 3424
rect 1534 3428 1540 3429
rect 1534 3424 1535 3428
rect 1539 3424 1540 3428
rect 1534 3423 1540 3424
rect 1718 3428 1724 3429
rect 1718 3424 1719 3428
rect 1723 3424 1724 3428
rect 1718 3423 1724 3424
rect 1902 3428 1908 3429
rect 1902 3424 1903 3428
rect 1907 3424 1908 3428
rect 1902 3423 1908 3424
rect 2006 3425 2012 3426
rect 110 3420 116 3421
rect 2006 3421 2007 3425
rect 2011 3421 2012 3425
rect 2006 3420 2012 3421
rect 2046 3419 2052 3420
rect 2046 3415 2047 3419
rect 2051 3415 2052 3419
rect 3942 3419 3948 3420
rect 2046 3414 2052 3415
rect 2126 3416 2132 3417
rect 2126 3412 2127 3416
rect 2131 3412 2132 3416
rect 2126 3411 2132 3412
rect 2310 3416 2316 3417
rect 2310 3412 2311 3416
rect 2315 3412 2316 3416
rect 2310 3411 2316 3412
rect 2494 3416 2500 3417
rect 2494 3412 2495 3416
rect 2499 3412 2500 3416
rect 2494 3411 2500 3412
rect 2678 3416 2684 3417
rect 2678 3412 2679 3416
rect 2683 3412 2684 3416
rect 2678 3411 2684 3412
rect 2862 3416 2868 3417
rect 2862 3412 2863 3416
rect 2867 3412 2868 3416
rect 2862 3411 2868 3412
rect 3046 3416 3052 3417
rect 3046 3412 3047 3416
rect 3051 3412 3052 3416
rect 3046 3411 3052 3412
rect 3222 3416 3228 3417
rect 3222 3412 3223 3416
rect 3227 3412 3228 3416
rect 3222 3411 3228 3412
rect 3406 3416 3412 3417
rect 3406 3412 3407 3416
rect 3411 3412 3412 3416
rect 3406 3411 3412 3412
rect 3590 3416 3596 3417
rect 3590 3412 3591 3416
rect 3595 3412 3596 3416
rect 3590 3411 3596 3412
rect 3774 3416 3780 3417
rect 3774 3412 3775 3416
rect 3779 3412 3780 3416
rect 3942 3415 3943 3419
rect 3947 3415 3948 3419
rect 3942 3414 3948 3415
rect 3774 3411 3780 3412
rect 134 3409 140 3410
rect 110 3408 116 3409
rect 110 3404 111 3408
rect 115 3404 116 3408
rect 134 3405 135 3409
rect 139 3405 140 3409
rect 134 3404 140 3405
rect 318 3409 324 3410
rect 318 3405 319 3409
rect 323 3405 324 3409
rect 318 3404 324 3405
rect 534 3409 540 3410
rect 534 3405 535 3409
rect 539 3405 540 3409
rect 534 3404 540 3405
rect 750 3409 756 3410
rect 750 3405 751 3409
rect 755 3405 756 3409
rect 750 3404 756 3405
rect 958 3409 964 3410
rect 958 3405 959 3409
rect 963 3405 964 3409
rect 958 3404 964 3405
rect 1158 3409 1164 3410
rect 1158 3405 1159 3409
rect 1163 3405 1164 3409
rect 1158 3404 1164 3405
rect 1350 3409 1356 3410
rect 1350 3405 1351 3409
rect 1355 3405 1356 3409
rect 1350 3404 1356 3405
rect 1534 3409 1540 3410
rect 1534 3405 1535 3409
rect 1539 3405 1540 3409
rect 1534 3404 1540 3405
rect 1718 3409 1724 3410
rect 1718 3405 1719 3409
rect 1723 3405 1724 3409
rect 1718 3404 1724 3405
rect 1902 3409 1908 3410
rect 1902 3405 1903 3409
rect 1907 3405 1908 3409
rect 1902 3404 1908 3405
rect 2006 3408 2012 3409
rect 2006 3404 2007 3408
rect 2011 3404 2012 3408
rect 110 3403 116 3404
rect 2006 3403 2012 3404
rect 110 3356 116 3357
rect 2006 3356 2012 3357
rect 110 3352 111 3356
rect 115 3352 116 3356
rect 110 3351 116 3352
rect 134 3355 140 3356
rect 134 3351 135 3355
rect 139 3351 140 3355
rect 134 3350 140 3351
rect 230 3355 236 3356
rect 230 3351 231 3355
rect 235 3351 236 3355
rect 230 3350 236 3351
rect 374 3355 380 3356
rect 374 3351 375 3355
rect 379 3351 380 3355
rect 374 3350 380 3351
rect 534 3355 540 3356
rect 534 3351 535 3355
rect 539 3351 540 3355
rect 534 3350 540 3351
rect 702 3355 708 3356
rect 702 3351 703 3355
rect 707 3351 708 3355
rect 702 3350 708 3351
rect 870 3355 876 3356
rect 870 3351 871 3355
rect 875 3351 876 3355
rect 870 3350 876 3351
rect 1046 3355 1052 3356
rect 1046 3351 1047 3355
rect 1051 3351 1052 3355
rect 1046 3350 1052 3351
rect 1214 3355 1220 3356
rect 1214 3351 1215 3355
rect 1219 3351 1220 3355
rect 1214 3350 1220 3351
rect 1382 3355 1388 3356
rect 1382 3351 1383 3355
rect 1387 3351 1388 3355
rect 1382 3350 1388 3351
rect 1542 3355 1548 3356
rect 1542 3351 1543 3355
rect 1547 3351 1548 3355
rect 1542 3350 1548 3351
rect 1702 3355 1708 3356
rect 1702 3351 1703 3355
rect 1707 3351 1708 3355
rect 1702 3350 1708 3351
rect 1870 3355 1876 3356
rect 1870 3351 1871 3355
rect 1875 3351 1876 3355
rect 2006 3352 2007 3356
rect 2011 3352 2012 3356
rect 2006 3351 2012 3352
rect 1870 3350 1876 3351
rect 2070 3340 2076 3341
rect 110 3339 116 3340
rect 110 3335 111 3339
rect 115 3335 116 3339
rect 2006 3339 2012 3340
rect 110 3334 116 3335
rect 134 3336 140 3337
rect 134 3332 135 3336
rect 139 3332 140 3336
rect 134 3331 140 3332
rect 230 3336 236 3337
rect 230 3332 231 3336
rect 235 3332 236 3336
rect 230 3331 236 3332
rect 374 3336 380 3337
rect 374 3332 375 3336
rect 379 3332 380 3336
rect 374 3331 380 3332
rect 534 3336 540 3337
rect 534 3332 535 3336
rect 539 3332 540 3336
rect 534 3331 540 3332
rect 702 3336 708 3337
rect 702 3332 703 3336
rect 707 3332 708 3336
rect 702 3331 708 3332
rect 870 3336 876 3337
rect 870 3332 871 3336
rect 875 3332 876 3336
rect 870 3331 876 3332
rect 1046 3336 1052 3337
rect 1046 3332 1047 3336
rect 1051 3332 1052 3336
rect 1046 3331 1052 3332
rect 1214 3336 1220 3337
rect 1214 3332 1215 3336
rect 1219 3332 1220 3336
rect 1214 3331 1220 3332
rect 1382 3336 1388 3337
rect 1382 3332 1383 3336
rect 1387 3332 1388 3336
rect 1382 3331 1388 3332
rect 1542 3336 1548 3337
rect 1542 3332 1543 3336
rect 1547 3332 1548 3336
rect 1542 3331 1548 3332
rect 1702 3336 1708 3337
rect 1702 3332 1703 3336
rect 1707 3332 1708 3336
rect 1702 3331 1708 3332
rect 1870 3336 1876 3337
rect 1870 3332 1871 3336
rect 1875 3332 1876 3336
rect 2006 3335 2007 3339
rect 2011 3335 2012 3339
rect 2006 3334 2012 3335
rect 2046 3337 2052 3338
rect 2046 3333 2047 3337
rect 2051 3333 2052 3337
rect 2070 3336 2071 3340
rect 2075 3336 2076 3340
rect 2070 3335 2076 3336
rect 2214 3340 2220 3341
rect 2214 3336 2215 3340
rect 2219 3336 2220 3340
rect 2214 3335 2220 3336
rect 2358 3340 2364 3341
rect 2358 3336 2359 3340
rect 2363 3336 2364 3340
rect 2358 3335 2364 3336
rect 2510 3340 2516 3341
rect 2510 3336 2511 3340
rect 2515 3336 2516 3340
rect 2510 3335 2516 3336
rect 2654 3340 2660 3341
rect 2654 3336 2655 3340
rect 2659 3336 2660 3340
rect 2654 3335 2660 3336
rect 2798 3340 2804 3341
rect 2798 3336 2799 3340
rect 2803 3336 2804 3340
rect 2798 3335 2804 3336
rect 2934 3340 2940 3341
rect 2934 3336 2935 3340
rect 2939 3336 2940 3340
rect 2934 3335 2940 3336
rect 3078 3340 3084 3341
rect 3078 3336 3079 3340
rect 3083 3336 3084 3340
rect 3078 3335 3084 3336
rect 3222 3340 3228 3341
rect 3222 3336 3223 3340
rect 3227 3336 3228 3340
rect 3222 3335 3228 3336
rect 3374 3340 3380 3341
rect 3374 3336 3375 3340
rect 3379 3336 3380 3340
rect 3374 3335 3380 3336
rect 3534 3340 3540 3341
rect 3534 3336 3535 3340
rect 3539 3336 3540 3340
rect 3534 3335 3540 3336
rect 3694 3340 3700 3341
rect 3694 3336 3695 3340
rect 3699 3336 3700 3340
rect 3694 3335 3700 3336
rect 3838 3340 3844 3341
rect 3838 3336 3839 3340
rect 3843 3336 3844 3340
rect 3838 3335 3844 3336
rect 3942 3337 3948 3338
rect 2046 3332 2052 3333
rect 3942 3333 3943 3337
rect 3947 3333 3948 3337
rect 3942 3332 3948 3333
rect 1870 3331 1876 3332
rect 2070 3321 2076 3322
rect 2046 3320 2052 3321
rect 2046 3316 2047 3320
rect 2051 3316 2052 3320
rect 2070 3317 2071 3321
rect 2075 3317 2076 3321
rect 2070 3316 2076 3317
rect 2214 3321 2220 3322
rect 2214 3317 2215 3321
rect 2219 3317 2220 3321
rect 2214 3316 2220 3317
rect 2358 3321 2364 3322
rect 2358 3317 2359 3321
rect 2363 3317 2364 3321
rect 2358 3316 2364 3317
rect 2510 3321 2516 3322
rect 2510 3317 2511 3321
rect 2515 3317 2516 3321
rect 2510 3316 2516 3317
rect 2654 3321 2660 3322
rect 2654 3317 2655 3321
rect 2659 3317 2660 3321
rect 2654 3316 2660 3317
rect 2798 3321 2804 3322
rect 2798 3317 2799 3321
rect 2803 3317 2804 3321
rect 2798 3316 2804 3317
rect 2934 3321 2940 3322
rect 2934 3317 2935 3321
rect 2939 3317 2940 3321
rect 2934 3316 2940 3317
rect 3078 3321 3084 3322
rect 3078 3317 3079 3321
rect 3083 3317 3084 3321
rect 3078 3316 3084 3317
rect 3222 3321 3228 3322
rect 3222 3317 3223 3321
rect 3227 3317 3228 3321
rect 3222 3316 3228 3317
rect 3374 3321 3380 3322
rect 3374 3317 3375 3321
rect 3379 3317 3380 3321
rect 3374 3316 3380 3317
rect 3534 3321 3540 3322
rect 3534 3317 3535 3321
rect 3539 3317 3540 3321
rect 3534 3316 3540 3317
rect 3694 3321 3700 3322
rect 3694 3317 3695 3321
rect 3699 3317 3700 3321
rect 3694 3316 3700 3317
rect 3838 3321 3844 3322
rect 3838 3317 3839 3321
rect 3843 3317 3844 3321
rect 3838 3316 3844 3317
rect 3942 3320 3948 3321
rect 3942 3316 3943 3320
rect 3947 3316 3948 3320
rect 2046 3315 2052 3316
rect 3942 3315 3948 3316
rect 134 3276 140 3277
rect 110 3273 116 3274
rect 110 3269 111 3273
rect 115 3269 116 3273
rect 134 3272 135 3276
rect 139 3272 140 3276
rect 134 3271 140 3272
rect 278 3276 284 3277
rect 278 3272 279 3276
rect 283 3272 284 3276
rect 278 3271 284 3272
rect 462 3276 468 3277
rect 462 3272 463 3276
rect 467 3272 468 3276
rect 462 3271 468 3272
rect 662 3276 668 3277
rect 662 3272 663 3276
rect 667 3272 668 3276
rect 662 3271 668 3272
rect 870 3276 876 3277
rect 870 3272 871 3276
rect 875 3272 876 3276
rect 870 3271 876 3272
rect 1078 3276 1084 3277
rect 1078 3272 1079 3276
rect 1083 3272 1084 3276
rect 1078 3271 1084 3272
rect 1294 3276 1300 3277
rect 1294 3272 1295 3276
rect 1299 3272 1300 3276
rect 1294 3271 1300 3272
rect 1518 3276 1524 3277
rect 1518 3272 1519 3276
rect 1523 3272 1524 3276
rect 1518 3271 1524 3272
rect 1742 3276 1748 3277
rect 1742 3272 1743 3276
rect 1747 3272 1748 3276
rect 1742 3271 1748 3272
rect 2006 3273 2012 3274
rect 110 3268 116 3269
rect 2006 3269 2007 3273
rect 2011 3269 2012 3273
rect 2006 3268 2012 3269
rect 2046 3260 2052 3261
rect 3942 3260 3948 3261
rect 134 3257 140 3258
rect 110 3256 116 3257
rect 110 3252 111 3256
rect 115 3252 116 3256
rect 134 3253 135 3257
rect 139 3253 140 3257
rect 134 3252 140 3253
rect 278 3257 284 3258
rect 278 3253 279 3257
rect 283 3253 284 3257
rect 278 3252 284 3253
rect 462 3257 468 3258
rect 462 3253 463 3257
rect 467 3253 468 3257
rect 462 3252 468 3253
rect 662 3257 668 3258
rect 662 3253 663 3257
rect 667 3253 668 3257
rect 662 3252 668 3253
rect 870 3257 876 3258
rect 870 3253 871 3257
rect 875 3253 876 3257
rect 870 3252 876 3253
rect 1078 3257 1084 3258
rect 1078 3253 1079 3257
rect 1083 3253 1084 3257
rect 1078 3252 1084 3253
rect 1294 3257 1300 3258
rect 1294 3253 1295 3257
rect 1299 3253 1300 3257
rect 1294 3252 1300 3253
rect 1518 3257 1524 3258
rect 1518 3253 1519 3257
rect 1523 3253 1524 3257
rect 1518 3252 1524 3253
rect 1742 3257 1748 3258
rect 1742 3253 1743 3257
rect 1747 3253 1748 3257
rect 1742 3252 1748 3253
rect 2006 3256 2012 3257
rect 2006 3252 2007 3256
rect 2011 3252 2012 3256
rect 2046 3256 2047 3260
rect 2051 3256 2052 3260
rect 2046 3255 2052 3256
rect 2110 3259 2116 3260
rect 2110 3255 2111 3259
rect 2115 3255 2116 3259
rect 2110 3254 2116 3255
rect 2246 3259 2252 3260
rect 2246 3255 2247 3259
rect 2251 3255 2252 3259
rect 2246 3254 2252 3255
rect 2398 3259 2404 3260
rect 2398 3255 2399 3259
rect 2403 3255 2404 3259
rect 2398 3254 2404 3255
rect 2574 3259 2580 3260
rect 2574 3255 2575 3259
rect 2579 3255 2580 3259
rect 2574 3254 2580 3255
rect 2782 3259 2788 3260
rect 2782 3255 2783 3259
rect 2787 3255 2788 3259
rect 2782 3254 2788 3255
rect 3014 3259 3020 3260
rect 3014 3255 3015 3259
rect 3019 3255 3020 3259
rect 3014 3254 3020 3255
rect 3262 3259 3268 3260
rect 3262 3255 3263 3259
rect 3267 3255 3268 3259
rect 3262 3254 3268 3255
rect 3526 3259 3532 3260
rect 3526 3255 3527 3259
rect 3531 3255 3532 3259
rect 3526 3254 3532 3255
rect 3790 3259 3796 3260
rect 3790 3255 3791 3259
rect 3795 3255 3796 3259
rect 3942 3256 3943 3260
rect 3947 3256 3948 3260
rect 3942 3255 3948 3256
rect 3790 3254 3796 3255
rect 110 3251 116 3252
rect 2006 3251 2012 3252
rect 2046 3243 2052 3244
rect 2046 3239 2047 3243
rect 2051 3239 2052 3243
rect 3942 3243 3948 3244
rect 2046 3238 2052 3239
rect 2110 3240 2116 3241
rect 2110 3236 2111 3240
rect 2115 3236 2116 3240
rect 2110 3235 2116 3236
rect 2246 3240 2252 3241
rect 2246 3236 2247 3240
rect 2251 3236 2252 3240
rect 2246 3235 2252 3236
rect 2398 3240 2404 3241
rect 2398 3236 2399 3240
rect 2403 3236 2404 3240
rect 2398 3235 2404 3236
rect 2574 3240 2580 3241
rect 2574 3236 2575 3240
rect 2579 3236 2580 3240
rect 2574 3235 2580 3236
rect 2782 3240 2788 3241
rect 2782 3236 2783 3240
rect 2787 3236 2788 3240
rect 2782 3235 2788 3236
rect 3014 3240 3020 3241
rect 3014 3236 3015 3240
rect 3019 3236 3020 3240
rect 3014 3235 3020 3236
rect 3262 3240 3268 3241
rect 3262 3236 3263 3240
rect 3267 3236 3268 3240
rect 3262 3235 3268 3236
rect 3526 3240 3532 3241
rect 3526 3236 3527 3240
rect 3531 3236 3532 3240
rect 3526 3235 3532 3236
rect 3790 3240 3796 3241
rect 3790 3236 3791 3240
rect 3795 3236 3796 3240
rect 3942 3239 3943 3243
rect 3947 3239 3948 3243
rect 3942 3238 3948 3239
rect 3790 3235 3796 3236
rect 110 3204 116 3205
rect 2006 3204 2012 3205
rect 110 3200 111 3204
rect 115 3200 116 3204
rect 110 3199 116 3200
rect 134 3203 140 3204
rect 134 3199 135 3203
rect 139 3199 140 3203
rect 134 3198 140 3199
rect 286 3203 292 3204
rect 286 3199 287 3203
rect 291 3199 292 3203
rect 286 3198 292 3199
rect 446 3203 452 3204
rect 446 3199 447 3203
rect 451 3199 452 3203
rect 446 3198 452 3199
rect 614 3203 620 3204
rect 614 3199 615 3203
rect 619 3199 620 3203
rect 614 3198 620 3199
rect 790 3203 796 3204
rect 790 3199 791 3203
rect 795 3199 796 3203
rect 790 3198 796 3199
rect 966 3203 972 3204
rect 966 3199 967 3203
rect 971 3199 972 3203
rect 966 3198 972 3199
rect 1142 3203 1148 3204
rect 1142 3199 1143 3203
rect 1147 3199 1148 3203
rect 1142 3198 1148 3199
rect 1326 3203 1332 3204
rect 1326 3199 1327 3203
rect 1331 3199 1332 3203
rect 1326 3198 1332 3199
rect 1510 3203 1516 3204
rect 1510 3199 1511 3203
rect 1515 3199 1516 3203
rect 1510 3198 1516 3199
rect 1694 3203 1700 3204
rect 1694 3199 1695 3203
rect 1699 3199 1700 3203
rect 2006 3200 2007 3204
rect 2011 3200 2012 3204
rect 2006 3199 2012 3200
rect 1694 3198 1700 3199
rect 110 3187 116 3188
rect 110 3183 111 3187
rect 115 3183 116 3187
rect 2006 3187 2012 3188
rect 110 3182 116 3183
rect 134 3184 140 3185
rect 134 3180 135 3184
rect 139 3180 140 3184
rect 134 3179 140 3180
rect 286 3184 292 3185
rect 286 3180 287 3184
rect 291 3180 292 3184
rect 286 3179 292 3180
rect 446 3184 452 3185
rect 446 3180 447 3184
rect 451 3180 452 3184
rect 446 3179 452 3180
rect 614 3184 620 3185
rect 614 3180 615 3184
rect 619 3180 620 3184
rect 614 3179 620 3180
rect 790 3184 796 3185
rect 790 3180 791 3184
rect 795 3180 796 3184
rect 790 3179 796 3180
rect 966 3184 972 3185
rect 966 3180 967 3184
rect 971 3180 972 3184
rect 966 3179 972 3180
rect 1142 3184 1148 3185
rect 1142 3180 1143 3184
rect 1147 3180 1148 3184
rect 1142 3179 1148 3180
rect 1326 3184 1332 3185
rect 1326 3180 1327 3184
rect 1331 3180 1332 3184
rect 1326 3179 1332 3180
rect 1510 3184 1516 3185
rect 1510 3180 1511 3184
rect 1515 3180 1516 3184
rect 1510 3179 1516 3180
rect 1694 3184 1700 3185
rect 1694 3180 1695 3184
rect 1699 3180 1700 3184
rect 2006 3183 2007 3187
rect 2011 3183 2012 3187
rect 2006 3182 2012 3183
rect 1694 3179 1700 3180
rect 2070 3180 2076 3181
rect 2046 3177 2052 3178
rect 2046 3173 2047 3177
rect 2051 3173 2052 3177
rect 2070 3176 2071 3180
rect 2075 3176 2076 3180
rect 2070 3175 2076 3176
rect 2166 3180 2172 3181
rect 2166 3176 2167 3180
rect 2171 3176 2172 3180
rect 2166 3175 2172 3176
rect 2262 3180 2268 3181
rect 2262 3176 2263 3180
rect 2267 3176 2268 3180
rect 2262 3175 2268 3176
rect 2358 3180 2364 3181
rect 2358 3176 2359 3180
rect 2363 3176 2364 3180
rect 2358 3175 2364 3176
rect 2454 3180 2460 3181
rect 2454 3176 2455 3180
rect 2459 3176 2460 3180
rect 2454 3175 2460 3176
rect 2550 3180 2556 3181
rect 2550 3176 2551 3180
rect 2555 3176 2556 3180
rect 2550 3175 2556 3176
rect 2646 3180 2652 3181
rect 2646 3176 2647 3180
rect 2651 3176 2652 3180
rect 2646 3175 2652 3176
rect 2742 3180 2748 3181
rect 2742 3176 2743 3180
rect 2747 3176 2748 3180
rect 2742 3175 2748 3176
rect 2838 3180 2844 3181
rect 2838 3176 2839 3180
rect 2843 3176 2844 3180
rect 2838 3175 2844 3176
rect 2934 3180 2940 3181
rect 2934 3176 2935 3180
rect 2939 3176 2940 3180
rect 2934 3175 2940 3176
rect 3030 3180 3036 3181
rect 3030 3176 3031 3180
rect 3035 3176 3036 3180
rect 3030 3175 3036 3176
rect 3126 3180 3132 3181
rect 3126 3176 3127 3180
rect 3131 3176 3132 3180
rect 3126 3175 3132 3176
rect 3222 3180 3228 3181
rect 3222 3176 3223 3180
rect 3227 3176 3228 3180
rect 3222 3175 3228 3176
rect 3318 3180 3324 3181
rect 3318 3176 3319 3180
rect 3323 3176 3324 3180
rect 3318 3175 3324 3176
rect 3438 3180 3444 3181
rect 3438 3176 3439 3180
rect 3443 3176 3444 3180
rect 3438 3175 3444 3176
rect 3574 3180 3580 3181
rect 3574 3176 3575 3180
rect 3579 3176 3580 3180
rect 3574 3175 3580 3176
rect 3718 3180 3724 3181
rect 3718 3176 3719 3180
rect 3723 3176 3724 3180
rect 3718 3175 3724 3176
rect 3838 3180 3844 3181
rect 3838 3176 3839 3180
rect 3843 3176 3844 3180
rect 3838 3175 3844 3176
rect 3942 3177 3948 3178
rect 2046 3172 2052 3173
rect 3942 3173 3943 3177
rect 3947 3173 3948 3177
rect 3942 3172 3948 3173
rect 2070 3161 2076 3162
rect 2046 3160 2052 3161
rect 2046 3156 2047 3160
rect 2051 3156 2052 3160
rect 2070 3157 2071 3161
rect 2075 3157 2076 3161
rect 2070 3156 2076 3157
rect 2166 3161 2172 3162
rect 2166 3157 2167 3161
rect 2171 3157 2172 3161
rect 2166 3156 2172 3157
rect 2262 3161 2268 3162
rect 2262 3157 2263 3161
rect 2267 3157 2268 3161
rect 2262 3156 2268 3157
rect 2358 3161 2364 3162
rect 2358 3157 2359 3161
rect 2363 3157 2364 3161
rect 2358 3156 2364 3157
rect 2454 3161 2460 3162
rect 2454 3157 2455 3161
rect 2459 3157 2460 3161
rect 2454 3156 2460 3157
rect 2550 3161 2556 3162
rect 2550 3157 2551 3161
rect 2555 3157 2556 3161
rect 2550 3156 2556 3157
rect 2646 3161 2652 3162
rect 2646 3157 2647 3161
rect 2651 3157 2652 3161
rect 2646 3156 2652 3157
rect 2742 3161 2748 3162
rect 2742 3157 2743 3161
rect 2747 3157 2748 3161
rect 2742 3156 2748 3157
rect 2838 3161 2844 3162
rect 2838 3157 2839 3161
rect 2843 3157 2844 3161
rect 2838 3156 2844 3157
rect 2934 3161 2940 3162
rect 2934 3157 2935 3161
rect 2939 3157 2940 3161
rect 2934 3156 2940 3157
rect 3030 3161 3036 3162
rect 3030 3157 3031 3161
rect 3035 3157 3036 3161
rect 3030 3156 3036 3157
rect 3126 3161 3132 3162
rect 3126 3157 3127 3161
rect 3131 3157 3132 3161
rect 3126 3156 3132 3157
rect 3222 3161 3228 3162
rect 3222 3157 3223 3161
rect 3227 3157 3228 3161
rect 3222 3156 3228 3157
rect 3318 3161 3324 3162
rect 3318 3157 3319 3161
rect 3323 3157 3324 3161
rect 3318 3156 3324 3157
rect 3438 3161 3444 3162
rect 3438 3157 3439 3161
rect 3443 3157 3444 3161
rect 3438 3156 3444 3157
rect 3574 3161 3580 3162
rect 3574 3157 3575 3161
rect 3579 3157 3580 3161
rect 3574 3156 3580 3157
rect 3718 3161 3724 3162
rect 3718 3157 3719 3161
rect 3723 3157 3724 3161
rect 3718 3156 3724 3157
rect 3838 3161 3844 3162
rect 3838 3157 3839 3161
rect 3843 3157 3844 3161
rect 3838 3156 3844 3157
rect 3942 3160 3948 3161
rect 3942 3156 3943 3160
rect 3947 3156 3948 3160
rect 2046 3155 2052 3156
rect 3942 3155 3948 3156
rect 310 3120 316 3121
rect 110 3117 116 3118
rect 110 3113 111 3117
rect 115 3113 116 3117
rect 310 3116 311 3120
rect 315 3116 316 3120
rect 310 3115 316 3116
rect 438 3120 444 3121
rect 438 3116 439 3120
rect 443 3116 444 3120
rect 438 3115 444 3116
rect 582 3120 588 3121
rect 582 3116 583 3120
rect 587 3116 588 3120
rect 582 3115 588 3116
rect 742 3120 748 3121
rect 742 3116 743 3120
rect 747 3116 748 3120
rect 742 3115 748 3116
rect 902 3120 908 3121
rect 902 3116 903 3120
rect 907 3116 908 3120
rect 902 3115 908 3116
rect 1062 3120 1068 3121
rect 1062 3116 1063 3120
rect 1067 3116 1068 3120
rect 1062 3115 1068 3116
rect 1222 3120 1228 3121
rect 1222 3116 1223 3120
rect 1227 3116 1228 3120
rect 1222 3115 1228 3116
rect 1390 3120 1396 3121
rect 1390 3116 1391 3120
rect 1395 3116 1396 3120
rect 1390 3115 1396 3116
rect 1558 3120 1564 3121
rect 1558 3116 1559 3120
rect 1563 3116 1564 3120
rect 1558 3115 1564 3116
rect 1726 3120 1732 3121
rect 1726 3116 1727 3120
rect 1731 3116 1732 3120
rect 1726 3115 1732 3116
rect 2006 3117 2012 3118
rect 110 3112 116 3113
rect 2006 3113 2007 3117
rect 2011 3113 2012 3117
rect 2006 3112 2012 3113
rect 310 3101 316 3102
rect 110 3100 116 3101
rect 110 3096 111 3100
rect 115 3096 116 3100
rect 310 3097 311 3101
rect 315 3097 316 3101
rect 310 3096 316 3097
rect 438 3101 444 3102
rect 438 3097 439 3101
rect 443 3097 444 3101
rect 438 3096 444 3097
rect 582 3101 588 3102
rect 582 3097 583 3101
rect 587 3097 588 3101
rect 582 3096 588 3097
rect 742 3101 748 3102
rect 742 3097 743 3101
rect 747 3097 748 3101
rect 742 3096 748 3097
rect 902 3101 908 3102
rect 902 3097 903 3101
rect 907 3097 908 3101
rect 902 3096 908 3097
rect 1062 3101 1068 3102
rect 1062 3097 1063 3101
rect 1067 3097 1068 3101
rect 1062 3096 1068 3097
rect 1222 3101 1228 3102
rect 1222 3097 1223 3101
rect 1227 3097 1228 3101
rect 1222 3096 1228 3097
rect 1390 3101 1396 3102
rect 1390 3097 1391 3101
rect 1395 3097 1396 3101
rect 1390 3096 1396 3097
rect 1558 3101 1564 3102
rect 1558 3097 1559 3101
rect 1563 3097 1564 3101
rect 1558 3096 1564 3097
rect 1726 3101 1732 3102
rect 1726 3097 1727 3101
rect 1731 3097 1732 3101
rect 1726 3096 1732 3097
rect 2006 3100 2012 3101
rect 2006 3096 2007 3100
rect 2011 3096 2012 3100
rect 110 3095 116 3096
rect 2006 3095 2012 3096
rect 2046 3096 2052 3097
rect 3942 3096 3948 3097
rect 2046 3092 2047 3096
rect 2051 3092 2052 3096
rect 2046 3091 2052 3092
rect 2070 3095 2076 3096
rect 2070 3091 2071 3095
rect 2075 3091 2076 3095
rect 2070 3090 2076 3091
rect 2334 3095 2340 3096
rect 2334 3091 2335 3095
rect 2339 3091 2340 3095
rect 2334 3090 2340 3091
rect 2622 3095 2628 3096
rect 2622 3091 2623 3095
rect 2627 3091 2628 3095
rect 2622 3090 2628 3091
rect 2910 3095 2916 3096
rect 2910 3091 2911 3095
rect 2915 3091 2916 3095
rect 2910 3090 2916 3091
rect 3206 3095 3212 3096
rect 3206 3091 3207 3095
rect 3211 3091 3212 3095
rect 3206 3090 3212 3091
rect 3502 3095 3508 3096
rect 3502 3091 3503 3095
rect 3507 3091 3508 3095
rect 3502 3090 3508 3091
rect 3798 3095 3804 3096
rect 3798 3091 3799 3095
rect 3803 3091 3804 3095
rect 3942 3092 3943 3096
rect 3947 3092 3948 3096
rect 3942 3091 3948 3092
rect 3798 3090 3804 3091
rect 2046 3079 2052 3080
rect 2046 3075 2047 3079
rect 2051 3075 2052 3079
rect 3942 3079 3948 3080
rect 2046 3074 2052 3075
rect 2070 3076 2076 3077
rect 2070 3072 2071 3076
rect 2075 3072 2076 3076
rect 2070 3071 2076 3072
rect 2334 3076 2340 3077
rect 2334 3072 2335 3076
rect 2339 3072 2340 3076
rect 2334 3071 2340 3072
rect 2622 3076 2628 3077
rect 2622 3072 2623 3076
rect 2627 3072 2628 3076
rect 2622 3071 2628 3072
rect 2910 3076 2916 3077
rect 2910 3072 2911 3076
rect 2915 3072 2916 3076
rect 2910 3071 2916 3072
rect 3206 3076 3212 3077
rect 3206 3072 3207 3076
rect 3211 3072 3212 3076
rect 3206 3071 3212 3072
rect 3502 3076 3508 3077
rect 3502 3072 3503 3076
rect 3507 3072 3508 3076
rect 3502 3071 3508 3072
rect 3798 3076 3804 3077
rect 3798 3072 3799 3076
rect 3803 3072 3804 3076
rect 3942 3075 3943 3079
rect 3947 3075 3948 3079
rect 3942 3074 3948 3075
rect 3798 3071 3804 3072
rect 110 3040 116 3041
rect 2006 3040 2012 3041
rect 110 3036 111 3040
rect 115 3036 116 3040
rect 110 3035 116 3036
rect 502 3039 508 3040
rect 502 3035 503 3039
rect 507 3035 508 3039
rect 502 3034 508 3035
rect 598 3039 604 3040
rect 598 3035 599 3039
rect 603 3035 604 3039
rect 598 3034 604 3035
rect 702 3039 708 3040
rect 702 3035 703 3039
rect 707 3035 708 3039
rect 702 3034 708 3035
rect 814 3039 820 3040
rect 814 3035 815 3039
rect 819 3035 820 3039
rect 814 3034 820 3035
rect 934 3039 940 3040
rect 934 3035 935 3039
rect 939 3035 940 3039
rect 934 3034 940 3035
rect 1070 3039 1076 3040
rect 1070 3035 1071 3039
rect 1075 3035 1076 3039
rect 1070 3034 1076 3035
rect 1222 3039 1228 3040
rect 1222 3035 1223 3039
rect 1227 3035 1228 3039
rect 1222 3034 1228 3035
rect 1382 3039 1388 3040
rect 1382 3035 1383 3039
rect 1387 3035 1388 3039
rect 1382 3034 1388 3035
rect 1550 3039 1556 3040
rect 1550 3035 1551 3039
rect 1555 3035 1556 3039
rect 1550 3034 1556 3035
rect 1718 3039 1724 3040
rect 1718 3035 1719 3039
rect 1723 3035 1724 3039
rect 2006 3036 2007 3040
rect 2011 3036 2012 3040
rect 2006 3035 2012 3036
rect 1718 3034 1724 3035
rect 110 3023 116 3024
rect 110 3019 111 3023
rect 115 3019 116 3023
rect 2006 3023 2012 3024
rect 110 3018 116 3019
rect 502 3020 508 3021
rect 502 3016 503 3020
rect 507 3016 508 3020
rect 502 3015 508 3016
rect 598 3020 604 3021
rect 598 3016 599 3020
rect 603 3016 604 3020
rect 598 3015 604 3016
rect 702 3020 708 3021
rect 702 3016 703 3020
rect 707 3016 708 3020
rect 702 3015 708 3016
rect 814 3020 820 3021
rect 814 3016 815 3020
rect 819 3016 820 3020
rect 814 3015 820 3016
rect 934 3020 940 3021
rect 934 3016 935 3020
rect 939 3016 940 3020
rect 934 3015 940 3016
rect 1070 3020 1076 3021
rect 1070 3016 1071 3020
rect 1075 3016 1076 3020
rect 1070 3015 1076 3016
rect 1222 3020 1228 3021
rect 1222 3016 1223 3020
rect 1227 3016 1228 3020
rect 1222 3015 1228 3016
rect 1382 3020 1388 3021
rect 1382 3016 1383 3020
rect 1387 3016 1388 3020
rect 1382 3015 1388 3016
rect 1550 3020 1556 3021
rect 1550 3016 1551 3020
rect 1555 3016 1556 3020
rect 1550 3015 1556 3016
rect 1718 3020 1724 3021
rect 1718 3016 1719 3020
rect 1723 3016 1724 3020
rect 2006 3019 2007 3023
rect 2011 3019 2012 3023
rect 2006 3018 2012 3019
rect 1718 3015 1724 3016
rect 2070 3016 2076 3017
rect 2046 3013 2052 3014
rect 2046 3009 2047 3013
rect 2051 3009 2052 3013
rect 2070 3012 2071 3016
rect 2075 3012 2076 3016
rect 2070 3011 2076 3012
rect 2382 3016 2388 3017
rect 2382 3012 2383 3016
rect 2387 3012 2388 3016
rect 2382 3011 2388 3012
rect 2702 3016 2708 3017
rect 2702 3012 2703 3016
rect 2707 3012 2708 3016
rect 2702 3011 2708 3012
rect 2998 3016 3004 3017
rect 2998 3012 2999 3016
rect 3003 3012 3004 3016
rect 2998 3011 3004 3012
rect 3286 3016 3292 3017
rect 3286 3012 3287 3016
rect 3291 3012 3292 3016
rect 3286 3011 3292 3012
rect 3574 3016 3580 3017
rect 3574 3012 3575 3016
rect 3579 3012 3580 3016
rect 3574 3011 3580 3012
rect 3838 3016 3844 3017
rect 3838 3012 3839 3016
rect 3843 3012 3844 3016
rect 3838 3011 3844 3012
rect 3942 3013 3948 3014
rect 2046 3008 2052 3009
rect 3942 3009 3943 3013
rect 3947 3009 3948 3013
rect 3942 3008 3948 3009
rect 2070 2997 2076 2998
rect 2046 2996 2052 2997
rect 2046 2992 2047 2996
rect 2051 2992 2052 2996
rect 2070 2993 2071 2997
rect 2075 2993 2076 2997
rect 2070 2992 2076 2993
rect 2382 2997 2388 2998
rect 2382 2993 2383 2997
rect 2387 2993 2388 2997
rect 2382 2992 2388 2993
rect 2702 2997 2708 2998
rect 2702 2993 2703 2997
rect 2707 2993 2708 2997
rect 2702 2992 2708 2993
rect 2998 2997 3004 2998
rect 2998 2993 2999 2997
rect 3003 2993 3004 2997
rect 2998 2992 3004 2993
rect 3286 2997 3292 2998
rect 3286 2993 3287 2997
rect 3291 2993 3292 2997
rect 3286 2992 3292 2993
rect 3574 2997 3580 2998
rect 3574 2993 3575 2997
rect 3579 2993 3580 2997
rect 3574 2992 3580 2993
rect 3838 2997 3844 2998
rect 3838 2993 3839 2997
rect 3843 2993 3844 2997
rect 3838 2992 3844 2993
rect 3942 2996 3948 2997
rect 3942 2992 3943 2996
rect 3947 2992 3948 2996
rect 2046 2991 2052 2992
rect 3942 2991 3948 2992
rect 550 2956 556 2957
rect 110 2953 116 2954
rect 110 2949 111 2953
rect 115 2949 116 2953
rect 550 2952 551 2956
rect 555 2952 556 2956
rect 550 2951 556 2952
rect 646 2956 652 2957
rect 646 2952 647 2956
rect 651 2952 652 2956
rect 646 2951 652 2952
rect 758 2956 764 2957
rect 758 2952 759 2956
rect 763 2952 764 2956
rect 758 2951 764 2952
rect 886 2956 892 2957
rect 886 2952 887 2956
rect 891 2952 892 2956
rect 886 2951 892 2952
rect 1022 2956 1028 2957
rect 1022 2952 1023 2956
rect 1027 2952 1028 2956
rect 1022 2951 1028 2952
rect 1174 2956 1180 2957
rect 1174 2952 1175 2956
rect 1179 2952 1180 2956
rect 1174 2951 1180 2952
rect 1326 2956 1332 2957
rect 1326 2952 1327 2956
rect 1331 2952 1332 2956
rect 1326 2951 1332 2952
rect 1486 2956 1492 2957
rect 1486 2952 1487 2956
rect 1491 2952 1492 2956
rect 1486 2951 1492 2952
rect 1654 2956 1660 2957
rect 1654 2952 1655 2956
rect 1659 2952 1660 2956
rect 1654 2951 1660 2952
rect 1822 2956 1828 2957
rect 1822 2952 1823 2956
rect 1827 2952 1828 2956
rect 1822 2951 1828 2952
rect 2006 2953 2012 2954
rect 110 2948 116 2949
rect 2006 2949 2007 2953
rect 2011 2949 2012 2953
rect 2006 2948 2012 2949
rect 2046 2940 2052 2941
rect 3942 2940 3948 2941
rect 550 2937 556 2938
rect 110 2936 116 2937
rect 110 2932 111 2936
rect 115 2932 116 2936
rect 550 2933 551 2937
rect 555 2933 556 2937
rect 550 2932 556 2933
rect 646 2937 652 2938
rect 646 2933 647 2937
rect 651 2933 652 2937
rect 646 2932 652 2933
rect 758 2937 764 2938
rect 758 2933 759 2937
rect 763 2933 764 2937
rect 758 2932 764 2933
rect 886 2937 892 2938
rect 886 2933 887 2937
rect 891 2933 892 2937
rect 886 2932 892 2933
rect 1022 2937 1028 2938
rect 1022 2933 1023 2937
rect 1027 2933 1028 2937
rect 1022 2932 1028 2933
rect 1174 2937 1180 2938
rect 1174 2933 1175 2937
rect 1179 2933 1180 2937
rect 1174 2932 1180 2933
rect 1326 2937 1332 2938
rect 1326 2933 1327 2937
rect 1331 2933 1332 2937
rect 1326 2932 1332 2933
rect 1486 2937 1492 2938
rect 1486 2933 1487 2937
rect 1491 2933 1492 2937
rect 1486 2932 1492 2933
rect 1654 2937 1660 2938
rect 1654 2933 1655 2937
rect 1659 2933 1660 2937
rect 1654 2932 1660 2933
rect 1822 2937 1828 2938
rect 1822 2933 1823 2937
rect 1827 2933 1828 2937
rect 1822 2932 1828 2933
rect 2006 2936 2012 2937
rect 2006 2932 2007 2936
rect 2011 2932 2012 2936
rect 2046 2936 2047 2940
rect 2051 2936 2052 2940
rect 2046 2935 2052 2936
rect 2070 2939 2076 2940
rect 2070 2935 2071 2939
rect 2075 2935 2076 2939
rect 2070 2934 2076 2935
rect 2390 2939 2396 2940
rect 2390 2935 2391 2939
rect 2395 2935 2396 2939
rect 2390 2934 2396 2935
rect 2702 2939 2708 2940
rect 2702 2935 2703 2939
rect 2707 2935 2708 2939
rect 2702 2934 2708 2935
rect 2974 2939 2980 2940
rect 2974 2935 2975 2939
rect 2979 2935 2980 2939
rect 2974 2934 2980 2935
rect 3214 2939 3220 2940
rect 3214 2935 3215 2939
rect 3219 2935 3220 2939
rect 3214 2934 3220 2935
rect 3438 2939 3444 2940
rect 3438 2935 3439 2939
rect 3443 2935 3444 2939
rect 3438 2934 3444 2935
rect 3646 2939 3652 2940
rect 3646 2935 3647 2939
rect 3651 2935 3652 2939
rect 3646 2934 3652 2935
rect 3838 2939 3844 2940
rect 3838 2935 3839 2939
rect 3843 2935 3844 2939
rect 3942 2936 3943 2940
rect 3947 2936 3948 2940
rect 3942 2935 3948 2936
rect 3838 2934 3844 2935
rect 110 2931 116 2932
rect 2006 2931 2012 2932
rect 2046 2923 2052 2924
rect 2046 2919 2047 2923
rect 2051 2919 2052 2923
rect 3942 2923 3948 2924
rect 2046 2918 2052 2919
rect 2070 2920 2076 2921
rect 2070 2916 2071 2920
rect 2075 2916 2076 2920
rect 2070 2915 2076 2916
rect 2390 2920 2396 2921
rect 2390 2916 2391 2920
rect 2395 2916 2396 2920
rect 2390 2915 2396 2916
rect 2702 2920 2708 2921
rect 2702 2916 2703 2920
rect 2707 2916 2708 2920
rect 2702 2915 2708 2916
rect 2974 2920 2980 2921
rect 2974 2916 2975 2920
rect 2979 2916 2980 2920
rect 2974 2915 2980 2916
rect 3214 2920 3220 2921
rect 3214 2916 3215 2920
rect 3219 2916 3220 2920
rect 3214 2915 3220 2916
rect 3438 2920 3444 2921
rect 3438 2916 3439 2920
rect 3443 2916 3444 2920
rect 3438 2915 3444 2916
rect 3646 2920 3652 2921
rect 3646 2916 3647 2920
rect 3651 2916 3652 2920
rect 3646 2915 3652 2916
rect 3838 2920 3844 2921
rect 3838 2916 3839 2920
rect 3843 2916 3844 2920
rect 3942 2919 3943 2923
rect 3947 2919 3948 2923
rect 3942 2918 3948 2919
rect 3838 2915 3844 2916
rect 110 2876 116 2877
rect 2006 2876 2012 2877
rect 110 2872 111 2876
rect 115 2872 116 2876
rect 110 2871 116 2872
rect 470 2875 476 2876
rect 470 2871 471 2875
rect 475 2871 476 2875
rect 470 2870 476 2871
rect 574 2875 580 2876
rect 574 2871 575 2875
rect 579 2871 580 2875
rect 574 2870 580 2871
rect 694 2875 700 2876
rect 694 2871 695 2875
rect 699 2871 700 2875
rect 694 2870 700 2871
rect 838 2875 844 2876
rect 838 2871 839 2875
rect 843 2871 844 2875
rect 838 2870 844 2871
rect 990 2875 996 2876
rect 990 2871 991 2875
rect 995 2871 996 2875
rect 990 2870 996 2871
rect 1150 2875 1156 2876
rect 1150 2871 1151 2875
rect 1155 2871 1156 2875
rect 1150 2870 1156 2871
rect 1318 2875 1324 2876
rect 1318 2871 1319 2875
rect 1323 2871 1324 2875
rect 1318 2870 1324 2871
rect 1494 2875 1500 2876
rect 1494 2871 1495 2875
rect 1499 2871 1500 2875
rect 1494 2870 1500 2871
rect 1670 2875 1676 2876
rect 1670 2871 1671 2875
rect 1675 2871 1676 2875
rect 1670 2870 1676 2871
rect 1846 2875 1852 2876
rect 1846 2871 1847 2875
rect 1851 2871 1852 2875
rect 2006 2872 2007 2876
rect 2011 2872 2012 2876
rect 2006 2871 2012 2872
rect 1846 2870 1852 2871
rect 2070 2860 2076 2861
rect 110 2859 116 2860
rect 110 2855 111 2859
rect 115 2855 116 2859
rect 2006 2859 2012 2860
rect 110 2854 116 2855
rect 470 2856 476 2857
rect 470 2852 471 2856
rect 475 2852 476 2856
rect 470 2851 476 2852
rect 574 2856 580 2857
rect 574 2852 575 2856
rect 579 2852 580 2856
rect 574 2851 580 2852
rect 694 2856 700 2857
rect 694 2852 695 2856
rect 699 2852 700 2856
rect 694 2851 700 2852
rect 838 2856 844 2857
rect 838 2852 839 2856
rect 843 2852 844 2856
rect 838 2851 844 2852
rect 990 2856 996 2857
rect 990 2852 991 2856
rect 995 2852 996 2856
rect 990 2851 996 2852
rect 1150 2856 1156 2857
rect 1150 2852 1151 2856
rect 1155 2852 1156 2856
rect 1150 2851 1156 2852
rect 1318 2856 1324 2857
rect 1318 2852 1319 2856
rect 1323 2852 1324 2856
rect 1318 2851 1324 2852
rect 1494 2856 1500 2857
rect 1494 2852 1495 2856
rect 1499 2852 1500 2856
rect 1494 2851 1500 2852
rect 1670 2856 1676 2857
rect 1670 2852 1671 2856
rect 1675 2852 1676 2856
rect 1670 2851 1676 2852
rect 1846 2856 1852 2857
rect 1846 2852 1847 2856
rect 1851 2852 1852 2856
rect 2006 2855 2007 2859
rect 2011 2855 2012 2859
rect 2006 2854 2012 2855
rect 2046 2857 2052 2858
rect 2046 2853 2047 2857
rect 2051 2853 2052 2857
rect 2070 2856 2071 2860
rect 2075 2856 2076 2860
rect 2070 2855 2076 2856
rect 2294 2860 2300 2861
rect 2294 2856 2295 2860
rect 2299 2856 2300 2860
rect 2294 2855 2300 2856
rect 2534 2860 2540 2861
rect 2534 2856 2535 2860
rect 2539 2856 2540 2860
rect 2534 2855 2540 2856
rect 2766 2860 2772 2861
rect 2766 2856 2767 2860
rect 2771 2856 2772 2860
rect 2766 2855 2772 2856
rect 2990 2860 2996 2861
rect 2990 2856 2991 2860
rect 2995 2856 2996 2860
rect 2990 2855 2996 2856
rect 3214 2860 3220 2861
rect 3214 2856 3215 2860
rect 3219 2856 3220 2860
rect 3214 2855 3220 2856
rect 3430 2860 3436 2861
rect 3430 2856 3431 2860
rect 3435 2856 3436 2860
rect 3430 2855 3436 2856
rect 3646 2860 3652 2861
rect 3646 2856 3647 2860
rect 3651 2856 3652 2860
rect 3646 2855 3652 2856
rect 3838 2860 3844 2861
rect 3838 2856 3839 2860
rect 3843 2856 3844 2860
rect 3838 2855 3844 2856
rect 3942 2857 3948 2858
rect 2046 2852 2052 2853
rect 3942 2853 3943 2857
rect 3947 2853 3948 2857
rect 3942 2852 3948 2853
rect 1846 2851 1852 2852
rect 2070 2841 2076 2842
rect 2046 2840 2052 2841
rect 2046 2836 2047 2840
rect 2051 2836 2052 2840
rect 2070 2837 2071 2841
rect 2075 2837 2076 2841
rect 2070 2836 2076 2837
rect 2294 2841 2300 2842
rect 2294 2837 2295 2841
rect 2299 2837 2300 2841
rect 2294 2836 2300 2837
rect 2534 2841 2540 2842
rect 2534 2837 2535 2841
rect 2539 2837 2540 2841
rect 2534 2836 2540 2837
rect 2766 2841 2772 2842
rect 2766 2837 2767 2841
rect 2771 2837 2772 2841
rect 2766 2836 2772 2837
rect 2990 2841 2996 2842
rect 2990 2837 2991 2841
rect 2995 2837 2996 2841
rect 2990 2836 2996 2837
rect 3214 2841 3220 2842
rect 3214 2837 3215 2841
rect 3219 2837 3220 2841
rect 3214 2836 3220 2837
rect 3430 2841 3436 2842
rect 3430 2837 3431 2841
rect 3435 2837 3436 2841
rect 3430 2836 3436 2837
rect 3646 2841 3652 2842
rect 3646 2837 3647 2841
rect 3651 2837 3652 2841
rect 3646 2836 3652 2837
rect 3838 2841 3844 2842
rect 3838 2837 3839 2841
rect 3843 2837 3844 2841
rect 3838 2836 3844 2837
rect 3942 2840 3948 2841
rect 3942 2836 3943 2840
rect 3947 2836 3948 2840
rect 2046 2835 2052 2836
rect 3942 2835 3948 2836
rect 478 2792 484 2793
rect 110 2789 116 2790
rect 110 2785 111 2789
rect 115 2785 116 2789
rect 478 2788 479 2792
rect 483 2788 484 2792
rect 478 2787 484 2788
rect 574 2792 580 2793
rect 574 2788 575 2792
rect 579 2788 580 2792
rect 574 2787 580 2788
rect 678 2792 684 2793
rect 678 2788 679 2792
rect 683 2788 684 2792
rect 678 2787 684 2788
rect 798 2792 804 2793
rect 798 2788 799 2792
rect 803 2788 804 2792
rect 798 2787 804 2788
rect 934 2792 940 2793
rect 934 2788 935 2792
rect 939 2788 940 2792
rect 934 2787 940 2788
rect 1078 2792 1084 2793
rect 1078 2788 1079 2792
rect 1083 2788 1084 2792
rect 1078 2787 1084 2788
rect 1238 2792 1244 2793
rect 1238 2788 1239 2792
rect 1243 2788 1244 2792
rect 1238 2787 1244 2788
rect 1414 2792 1420 2793
rect 1414 2788 1415 2792
rect 1419 2788 1420 2792
rect 1414 2787 1420 2788
rect 1598 2792 1604 2793
rect 1598 2788 1599 2792
rect 1603 2788 1604 2792
rect 1598 2787 1604 2788
rect 1782 2792 1788 2793
rect 1782 2788 1783 2792
rect 1787 2788 1788 2792
rect 1782 2787 1788 2788
rect 2006 2789 2012 2790
rect 110 2784 116 2785
rect 2006 2785 2007 2789
rect 2011 2785 2012 2789
rect 2006 2784 2012 2785
rect 2046 2784 2052 2785
rect 3942 2784 3948 2785
rect 2046 2780 2047 2784
rect 2051 2780 2052 2784
rect 2046 2779 2052 2780
rect 2070 2783 2076 2784
rect 2070 2779 2071 2783
rect 2075 2779 2076 2783
rect 2070 2778 2076 2779
rect 2198 2783 2204 2784
rect 2198 2779 2199 2783
rect 2203 2779 2204 2783
rect 2198 2778 2204 2779
rect 2366 2783 2372 2784
rect 2366 2779 2367 2783
rect 2371 2779 2372 2783
rect 2366 2778 2372 2779
rect 2550 2783 2556 2784
rect 2550 2779 2551 2783
rect 2555 2779 2556 2783
rect 2550 2778 2556 2779
rect 2734 2783 2740 2784
rect 2734 2779 2735 2783
rect 2739 2779 2740 2783
rect 2734 2778 2740 2779
rect 2926 2783 2932 2784
rect 2926 2779 2927 2783
rect 2931 2779 2932 2783
rect 2926 2778 2932 2779
rect 3110 2783 3116 2784
rect 3110 2779 3111 2783
rect 3115 2779 3116 2783
rect 3110 2778 3116 2779
rect 3294 2783 3300 2784
rect 3294 2779 3295 2783
rect 3299 2779 3300 2783
rect 3294 2778 3300 2779
rect 3478 2783 3484 2784
rect 3478 2779 3479 2783
rect 3483 2779 3484 2783
rect 3478 2778 3484 2779
rect 3670 2783 3676 2784
rect 3670 2779 3671 2783
rect 3675 2779 3676 2783
rect 3670 2778 3676 2779
rect 3838 2783 3844 2784
rect 3838 2779 3839 2783
rect 3843 2779 3844 2783
rect 3942 2780 3943 2784
rect 3947 2780 3948 2784
rect 3942 2779 3948 2780
rect 3838 2778 3844 2779
rect 478 2773 484 2774
rect 110 2772 116 2773
rect 110 2768 111 2772
rect 115 2768 116 2772
rect 478 2769 479 2773
rect 483 2769 484 2773
rect 478 2768 484 2769
rect 574 2773 580 2774
rect 574 2769 575 2773
rect 579 2769 580 2773
rect 574 2768 580 2769
rect 678 2773 684 2774
rect 678 2769 679 2773
rect 683 2769 684 2773
rect 678 2768 684 2769
rect 798 2773 804 2774
rect 798 2769 799 2773
rect 803 2769 804 2773
rect 798 2768 804 2769
rect 934 2773 940 2774
rect 934 2769 935 2773
rect 939 2769 940 2773
rect 934 2768 940 2769
rect 1078 2773 1084 2774
rect 1078 2769 1079 2773
rect 1083 2769 1084 2773
rect 1078 2768 1084 2769
rect 1238 2773 1244 2774
rect 1238 2769 1239 2773
rect 1243 2769 1244 2773
rect 1238 2768 1244 2769
rect 1414 2773 1420 2774
rect 1414 2769 1415 2773
rect 1419 2769 1420 2773
rect 1414 2768 1420 2769
rect 1598 2773 1604 2774
rect 1598 2769 1599 2773
rect 1603 2769 1604 2773
rect 1598 2768 1604 2769
rect 1782 2773 1788 2774
rect 1782 2769 1783 2773
rect 1787 2769 1788 2773
rect 1782 2768 1788 2769
rect 2006 2772 2012 2773
rect 2006 2768 2007 2772
rect 2011 2768 2012 2772
rect 110 2767 116 2768
rect 2006 2767 2012 2768
rect 2046 2767 2052 2768
rect 2046 2763 2047 2767
rect 2051 2763 2052 2767
rect 3942 2767 3948 2768
rect 2046 2762 2052 2763
rect 2070 2764 2076 2765
rect 2070 2760 2071 2764
rect 2075 2760 2076 2764
rect 2070 2759 2076 2760
rect 2198 2764 2204 2765
rect 2198 2760 2199 2764
rect 2203 2760 2204 2764
rect 2198 2759 2204 2760
rect 2366 2764 2372 2765
rect 2366 2760 2367 2764
rect 2371 2760 2372 2764
rect 2366 2759 2372 2760
rect 2550 2764 2556 2765
rect 2550 2760 2551 2764
rect 2555 2760 2556 2764
rect 2550 2759 2556 2760
rect 2734 2764 2740 2765
rect 2734 2760 2735 2764
rect 2739 2760 2740 2764
rect 2734 2759 2740 2760
rect 2926 2764 2932 2765
rect 2926 2760 2927 2764
rect 2931 2760 2932 2764
rect 2926 2759 2932 2760
rect 3110 2764 3116 2765
rect 3110 2760 3111 2764
rect 3115 2760 3116 2764
rect 3110 2759 3116 2760
rect 3294 2764 3300 2765
rect 3294 2760 3295 2764
rect 3299 2760 3300 2764
rect 3294 2759 3300 2760
rect 3478 2764 3484 2765
rect 3478 2760 3479 2764
rect 3483 2760 3484 2764
rect 3478 2759 3484 2760
rect 3670 2764 3676 2765
rect 3670 2760 3671 2764
rect 3675 2760 3676 2764
rect 3670 2759 3676 2760
rect 3838 2764 3844 2765
rect 3838 2760 3839 2764
rect 3843 2760 3844 2764
rect 3942 2763 3943 2767
rect 3947 2763 3948 2767
rect 3942 2762 3948 2763
rect 3838 2759 3844 2760
rect 110 2716 116 2717
rect 2006 2716 2012 2717
rect 110 2712 111 2716
rect 115 2712 116 2716
rect 110 2711 116 2712
rect 510 2715 516 2716
rect 510 2711 511 2715
rect 515 2711 516 2715
rect 510 2710 516 2711
rect 622 2715 628 2716
rect 622 2711 623 2715
rect 627 2711 628 2715
rect 622 2710 628 2711
rect 742 2715 748 2716
rect 742 2711 743 2715
rect 747 2711 748 2715
rect 742 2710 748 2711
rect 878 2715 884 2716
rect 878 2711 879 2715
rect 883 2711 884 2715
rect 878 2710 884 2711
rect 1014 2715 1020 2716
rect 1014 2711 1015 2715
rect 1019 2711 1020 2715
rect 1014 2710 1020 2711
rect 1158 2715 1164 2716
rect 1158 2711 1159 2715
rect 1163 2711 1164 2715
rect 1158 2710 1164 2711
rect 1310 2715 1316 2716
rect 1310 2711 1311 2715
rect 1315 2711 1316 2715
rect 1310 2710 1316 2711
rect 1462 2715 1468 2716
rect 1462 2711 1463 2715
rect 1467 2711 1468 2715
rect 1462 2710 1468 2711
rect 1622 2715 1628 2716
rect 1622 2711 1623 2715
rect 1627 2711 1628 2715
rect 1622 2710 1628 2711
rect 1782 2715 1788 2716
rect 1782 2711 1783 2715
rect 1787 2711 1788 2715
rect 2006 2712 2007 2716
rect 2011 2712 2012 2716
rect 2006 2711 2012 2712
rect 1782 2710 1788 2711
rect 2070 2700 2076 2701
rect 110 2699 116 2700
rect 110 2695 111 2699
rect 115 2695 116 2699
rect 2006 2699 2012 2700
rect 110 2694 116 2695
rect 510 2696 516 2697
rect 510 2692 511 2696
rect 515 2692 516 2696
rect 510 2691 516 2692
rect 622 2696 628 2697
rect 622 2692 623 2696
rect 627 2692 628 2696
rect 622 2691 628 2692
rect 742 2696 748 2697
rect 742 2692 743 2696
rect 747 2692 748 2696
rect 742 2691 748 2692
rect 878 2696 884 2697
rect 878 2692 879 2696
rect 883 2692 884 2696
rect 878 2691 884 2692
rect 1014 2696 1020 2697
rect 1014 2692 1015 2696
rect 1019 2692 1020 2696
rect 1014 2691 1020 2692
rect 1158 2696 1164 2697
rect 1158 2692 1159 2696
rect 1163 2692 1164 2696
rect 1158 2691 1164 2692
rect 1310 2696 1316 2697
rect 1310 2692 1311 2696
rect 1315 2692 1316 2696
rect 1310 2691 1316 2692
rect 1462 2696 1468 2697
rect 1462 2692 1463 2696
rect 1467 2692 1468 2696
rect 1462 2691 1468 2692
rect 1622 2696 1628 2697
rect 1622 2692 1623 2696
rect 1627 2692 1628 2696
rect 1622 2691 1628 2692
rect 1782 2696 1788 2697
rect 1782 2692 1783 2696
rect 1787 2692 1788 2696
rect 2006 2695 2007 2699
rect 2011 2695 2012 2699
rect 2006 2694 2012 2695
rect 2046 2697 2052 2698
rect 2046 2693 2047 2697
rect 2051 2693 2052 2697
rect 2070 2696 2071 2700
rect 2075 2696 2076 2700
rect 2070 2695 2076 2696
rect 2190 2700 2196 2701
rect 2190 2696 2191 2700
rect 2195 2696 2196 2700
rect 2190 2695 2196 2696
rect 2318 2700 2324 2701
rect 2318 2696 2319 2700
rect 2323 2696 2324 2700
rect 2318 2695 2324 2696
rect 2446 2700 2452 2701
rect 2446 2696 2447 2700
rect 2451 2696 2452 2700
rect 2446 2695 2452 2696
rect 2582 2700 2588 2701
rect 2582 2696 2583 2700
rect 2587 2696 2588 2700
rect 2582 2695 2588 2696
rect 2726 2700 2732 2701
rect 2726 2696 2727 2700
rect 2731 2696 2732 2700
rect 2726 2695 2732 2696
rect 2886 2700 2892 2701
rect 2886 2696 2887 2700
rect 2891 2696 2892 2700
rect 2886 2695 2892 2696
rect 3062 2700 3068 2701
rect 3062 2696 3063 2700
rect 3067 2696 3068 2700
rect 3062 2695 3068 2696
rect 3254 2700 3260 2701
rect 3254 2696 3255 2700
rect 3259 2696 3260 2700
rect 3254 2695 3260 2696
rect 3454 2700 3460 2701
rect 3454 2696 3455 2700
rect 3459 2696 3460 2700
rect 3454 2695 3460 2696
rect 3654 2700 3660 2701
rect 3654 2696 3655 2700
rect 3659 2696 3660 2700
rect 3654 2695 3660 2696
rect 3838 2700 3844 2701
rect 3838 2696 3839 2700
rect 3843 2696 3844 2700
rect 3838 2695 3844 2696
rect 3942 2697 3948 2698
rect 2046 2692 2052 2693
rect 3942 2693 3943 2697
rect 3947 2693 3948 2697
rect 3942 2692 3948 2693
rect 1782 2691 1788 2692
rect 2070 2681 2076 2682
rect 2046 2680 2052 2681
rect 2046 2676 2047 2680
rect 2051 2676 2052 2680
rect 2070 2677 2071 2681
rect 2075 2677 2076 2681
rect 2070 2676 2076 2677
rect 2190 2681 2196 2682
rect 2190 2677 2191 2681
rect 2195 2677 2196 2681
rect 2190 2676 2196 2677
rect 2318 2681 2324 2682
rect 2318 2677 2319 2681
rect 2323 2677 2324 2681
rect 2318 2676 2324 2677
rect 2446 2681 2452 2682
rect 2446 2677 2447 2681
rect 2451 2677 2452 2681
rect 2446 2676 2452 2677
rect 2582 2681 2588 2682
rect 2582 2677 2583 2681
rect 2587 2677 2588 2681
rect 2582 2676 2588 2677
rect 2726 2681 2732 2682
rect 2726 2677 2727 2681
rect 2731 2677 2732 2681
rect 2726 2676 2732 2677
rect 2886 2681 2892 2682
rect 2886 2677 2887 2681
rect 2891 2677 2892 2681
rect 2886 2676 2892 2677
rect 3062 2681 3068 2682
rect 3062 2677 3063 2681
rect 3067 2677 3068 2681
rect 3062 2676 3068 2677
rect 3254 2681 3260 2682
rect 3254 2677 3255 2681
rect 3259 2677 3260 2681
rect 3254 2676 3260 2677
rect 3454 2681 3460 2682
rect 3454 2677 3455 2681
rect 3459 2677 3460 2681
rect 3454 2676 3460 2677
rect 3654 2681 3660 2682
rect 3654 2677 3655 2681
rect 3659 2677 3660 2681
rect 3654 2676 3660 2677
rect 3838 2681 3844 2682
rect 3838 2677 3839 2681
rect 3843 2677 3844 2681
rect 3838 2676 3844 2677
rect 3942 2680 3948 2681
rect 3942 2676 3943 2680
rect 3947 2676 3948 2680
rect 2046 2675 2052 2676
rect 3942 2675 3948 2676
rect 366 2632 372 2633
rect 110 2629 116 2630
rect 110 2625 111 2629
rect 115 2625 116 2629
rect 366 2628 367 2632
rect 371 2628 372 2632
rect 366 2627 372 2628
rect 486 2632 492 2633
rect 486 2628 487 2632
rect 491 2628 492 2632
rect 486 2627 492 2628
rect 614 2632 620 2633
rect 614 2628 615 2632
rect 619 2628 620 2632
rect 614 2627 620 2628
rect 750 2632 756 2633
rect 750 2628 751 2632
rect 755 2628 756 2632
rect 750 2627 756 2628
rect 894 2632 900 2633
rect 894 2628 895 2632
rect 899 2628 900 2632
rect 894 2627 900 2628
rect 1030 2632 1036 2633
rect 1030 2628 1031 2632
rect 1035 2628 1036 2632
rect 1030 2627 1036 2628
rect 1166 2632 1172 2633
rect 1166 2628 1167 2632
rect 1171 2628 1172 2632
rect 1166 2627 1172 2628
rect 1302 2632 1308 2633
rect 1302 2628 1303 2632
rect 1307 2628 1308 2632
rect 1302 2627 1308 2628
rect 1430 2632 1436 2633
rect 1430 2628 1431 2632
rect 1435 2628 1436 2632
rect 1430 2627 1436 2628
rect 1566 2632 1572 2633
rect 1566 2628 1567 2632
rect 1571 2628 1572 2632
rect 1566 2627 1572 2628
rect 1702 2632 1708 2633
rect 1702 2628 1703 2632
rect 1707 2628 1708 2632
rect 1702 2627 1708 2628
rect 2006 2629 2012 2630
rect 110 2624 116 2625
rect 2006 2625 2007 2629
rect 2011 2625 2012 2629
rect 2006 2624 2012 2625
rect 2046 2620 2052 2621
rect 3942 2620 3948 2621
rect 2046 2616 2047 2620
rect 2051 2616 2052 2620
rect 2046 2615 2052 2616
rect 2230 2619 2236 2620
rect 2230 2615 2231 2619
rect 2235 2615 2236 2619
rect 2230 2614 2236 2615
rect 2334 2619 2340 2620
rect 2334 2615 2335 2619
rect 2339 2615 2340 2619
rect 2334 2614 2340 2615
rect 2446 2619 2452 2620
rect 2446 2615 2447 2619
rect 2451 2615 2452 2619
rect 2446 2614 2452 2615
rect 2558 2619 2564 2620
rect 2558 2615 2559 2619
rect 2563 2615 2564 2619
rect 2558 2614 2564 2615
rect 2670 2619 2676 2620
rect 2670 2615 2671 2619
rect 2675 2615 2676 2619
rect 2670 2614 2676 2615
rect 2790 2619 2796 2620
rect 2790 2615 2791 2619
rect 2795 2615 2796 2619
rect 2790 2614 2796 2615
rect 2910 2619 2916 2620
rect 2910 2615 2911 2619
rect 2915 2615 2916 2619
rect 2910 2614 2916 2615
rect 3030 2619 3036 2620
rect 3030 2615 3031 2619
rect 3035 2615 3036 2619
rect 3030 2614 3036 2615
rect 3150 2619 3156 2620
rect 3150 2615 3151 2619
rect 3155 2615 3156 2619
rect 3942 2616 3943 2620
rect 3947 2616 3948 2620
rect 3942 2615 3948 2616
rect 3150 2614 3156 2615
rect 366 2613 372 2614
rect 110 2612 116 2613
rect 110 2608 111 2612
rect 115 2608 116 2612
rect 366 2609 367 2613
rect 371 2609 372 2613
rect 366 2608 372 2609
rect 486 2613 492 2614
rect 486 2609 487 2613
rect 491 2609 492 2613
rect 486 2608 492 2609
rect 614 2613 620 2614
rect 614 2609 615 2613
rect 619 2609 620 2613
rect 614 2608 620 2609
rect 750 2613 756 2614
rect 750 2609 751 2613
rect 755 2609 756 2613
rect 750 2608 756 2609
rect 894 2613 900 2614
rect 894 2609 895 2613
rect 899 2609 900 2613
rect 894 2608 900 2609
rect 1030 2613 1036 2614
rect 1030 2609 1031 2613
rect 1035 2609 1036 2613
rect 1030 2608 1036 2609
rect 1166 2613 1172 2614
rect 1166 2609 1167 2613
rect 1171 2609 1172 2613
rect 1166 2608 1172 2609
rect 1302 2613 1308 2614
rect 1302 2609 1303 2613
rect 1307 2609 1308 2613
rect 1302 2608 1308 2609
rect 1430 2613 1436 2614
rect 1430 2609 1431 2613
rect 1435 2609 1436 2613
rect 1430 2608 1436 2609
rect 1566 2613 1572 2614
rect 1566 2609 1567 2613
rect 1571 2609 1572 2613
rect 1566 2608 1572 2609
rect 1702 2613 1708 2614
rect 1702 2609 1703 2613
rect 1707 2609 1708 2613
rect 1702 2608 1708 2609
rect 2006 2612 2012 2613
rect 2006 2608 2007 2612
rect 2011 2608 2012 2612
rect 110 2607 116 2608
rect 2006 2607 2012 2608
rect 2046 2603 2052 2604
rect 2046 2599 2047 2603
rect 2051 2599 2052 2603
rect 3942 2603 3948 2604
rect 2046 2598 2052 2599
rect 2230 2600 2236 2601
rect 2230 2596 2231 2600
rect 2235 2596 2236 2600
rect 2230 2595 2236 2596
rect 2334 2600 2340 2601
rect 2334 2596 2335 2600
rect 2339 2596 2340 2600
rect 2334 2595 2340 2596
rect 2446 2600 2452 2601
rect 2446 2596 2447 2600
rect 2451 2596 2452 2600
rect 2446 2595 2452 2596
rect 2558 2600 2564 2601
rect 2558 2596 2559 2600
rect 2563 2596 2564 2600
rect 2558 2595 2564 2596
rect 2670 2600 2676 2601
rect 2670 2596 2671 2600
rect 2675 2596 2676 2600
rect 2670 2595 2676 2596
rect 2790 2600 2796 2601
rect 2790 2596 2791 2600
rect 2795 2596 2796 2600
rect 2790 2595 2796 2596
rect 2910 2600 2916 2601
rect 2910 2596 2911 2600
rect 2915 2596 2916 2600
rect 2910 2595 2916 2596
rect 3030 2600 3036 2601
rect 3030 2596 3031 2600
rect 3035 2596 3036 2600
rect 3030 2595 3036 2596
rect 3150 2600 3156 2601
rect 3150 2596 3151 2600
rect 3155 2596 3156 2600
rect 3942 2599 3943 2603
rect 3947 2599 3948 2603
rect 3942 2598 3948 2599
rect 3150 2595 3156 2596
rect 110 2560 116 2561
rect 2006 2560 2012 2561
rect 110 2556 111 2560
rect 115 2556 116 2560
rect 110 2555 116 2556
rect 134 2559 140 2560
rect 134 2555 135 2559
rect 139 2555 140 2559
rect 134 2554 140 2555
rect 286 2559 292 2560
rect 286 2555 287 2559
rect 291 2555 292 2559
rect 286 2554 292 2555
rect 446 2559 452 2560
rect 446 2555 447 2559
rect 451 2555 452 2559
rect 446 2554 452 2555
rect 606 2559 612 2560
rect 606 2555 607 2559
rect 611 2555 612 2559
rect 606 2554 612 2555
rect 766 2559 772 2560
rect 766 2555 767 2559
rect 771 2555 772 2559
rect 766 2554 772 2555
rect 918 2559 924 2560
rect 918 2555 919 2559
rect 923 2555 924 2559
rect 918 2554 924 2555
rect 1062 2559 1068 2560
rect 1062 2555 1063 2559
rect 1067 2555 1068 2559
rect 1062 2554 1068 2555
rect 1198 2559 1204 2560
rect 1198 2555 1199 2559
rect 1203 2555 1204 2559
rect 1198 2554 1204 2555
rect 1334 2559 1340 2560
rect 1334 2555 1335 2559
rect 1339 2555 1340 2559
rect 1334 2554 1340 2555
rect 1462 2559 1468 2560
rect 1462 2555 1463 2559
rect 1467 2555 1468 2559
rect 1462 2554 1468 2555
rect 1590 2559 1596 2560
rect 1590 2555 1591 2559
rect 1595 2555 1596 2559
rect 1590 2554 1596 2555
rect 1726 2559 1732 2560
rect 1726 2555 1727 2559
rect 1731 2555 1732 2559
rect 2006 2556 2007 2560
rect 2011 2556 2012 2560
rect 2006 2555 2012 2556
rect 1726 2554 1732 2555
rect 110 2543 116 2544
rect 110 2539 111 2543
rect 115 2539 116 2543
rect 2006 2543 2012 2544
rect 110 2538 116 2539
rect 134 2540 140 2541
rect 134 2536 135 2540
rect 139 2536 140 2540
rect 134 2535 140 2536
rect 286 2540 292 2541
rect 286 2536 287 2540
rect 291 2536 292 2540
rect 286 2535 292 2536
rect 446 2540 452 2541
rect 446 2536 447 2540
rect 451 2536 452 2540
rect 446 2535 452 2536
rect 606 2540 612 2541
rect 606 2536 607 2540
rect 611 2536 612 2540
rect 606 2535 612 2536
rect 766 2540 772 2541
rect 766 2536 767 2540
rect 771 2536 772 2540
rect 766 2535 772 2536
rect 918 2540 924 2541
rect 918 2536 919 2540
rect 923 2536 924 2540
rect 918 2535 924 2536
rect 1062 2540 1068 2541
rect 1062 2536 1063 2540
rect 1067 2536 1068 2540
rect 1062 2535 1068 2536
rect 1198 2540 1204 2541
rect 1198 2536 1199 2540
rect 1203 2536 1204 2540
rect 1198 2535 1204 2536
rect 1334 2540 1340 2541
rect 1334 2536 1335 2540
rect 1339 2536 1340 2540
rect 1334 2535 1340 2536
rect 1462 2540 1468 2541
rect 1462 2536 1463 2540
rect 1467 2536 1468 2540
rect 1462 2535 1468 2536
rect 1590 2540 1596 2541
rect 1590 2536 1591 2540
rect 1595 2536 1596 2540
rect 1590 2535 1596 2536
rect 1726 2540 1732 2541
rect 1726 2536 1727 2540
rect 1731 2536 1732 2540
rect 2006 2539 2007 2543
rect 2011 2539 2012 2543
rect 2006 2538 2012 2539
rect 1726 2535 1732 2536
rect 2382 2536 2388 2537
rect 2046 2533 2052 2534
rect 2046 2529 2047 2533
rect 2051 2529 2052 2533
rect 2382 2532 2383 2536
rect 2387 2532 2388 2536
rect 2382 2531 2388 2532
rect 2494 2536 2500 2537
rect 2494 2532 2495 2536
rect 2499 2532 2500 2536
rect 2494 2531 2500 2532
rect 2614 2536 2620 2537
rect 2614 2532 2615 2536
rect 2619 2532 2620 2536
rect 2614 2531 2620 2532
rect 2742 2536 2748 2537
rect 2742 2532 2743 2536
rect 2747 2532 2748 2536
rect 2742 2531 2748 2532
rect 2870 2536 2876 2537
rect 2870 2532 2871 2536
rect 2875 2532 2876 2536
rect 2870 2531 2876 2532
rect 2990 2536 2996 2537
rect 2990 2532 2991 2536
rect 2995 2532 2996 2536
rect 2990 2531 2996 2532
rect 3110 2536 3116 2537
rect 3110 2532 3111 2536
rect 3115 2532 3116 2536
rect 3110 2531 3116 2532
rect 3230 2536 3236 2537
rect 3230 2532 3231 2536
rect 3235 2532 3236 2536
rect 3230 2531 3236 2532
rect 3358 2536 3364 2537
rect 3358 2532 3359 2536
rect 3363 2532 3364 2536
rect 3358 2531 3364 2532
rect 3486 2536 3492 2537
rect 3486 2532 3487 2536
rect 3491 2532 3492 2536
rect 3486 2531 3492 2532
rect 3942 2533 3948 2534
rect 2046 2528 2052 2529
rect 3942 2529 3943 2533
rect 3947 2529 3948 2533
rect 3942 2528 3948 2529
rect 2382 2517 2388 2518
rect 2046 2516 2052 2517
rect 2046 2512 2047 2516
rect 2051 2512 2052 2516
rect 2382 2513 2383 2517
rect 2387 2513 2388 2517
rect 2382 2512 2388 2513
rect 2494 2517 2500 2518
rect 2494 2513 2495 2517
rect 2499 2513 2500 2517
rect 2494 2512 2500 2513
rect 2614 2517 2620 2518
rect 2614 2513 2615 2517
rect 2619 2513 2620 2517
rect 2614 2512 2620 2513
rect 2742 2517 2748 2518
rect 2742 2513 2743 2517
rect 2747 2513 2748 2517
rect 2742 2512 2748 2513
rect 2870 2517 2876 2518
rect 2870 2513 2871 2517
rect 2875 2513 2876 2517
rect 2870 2512 2876 2513
rect 2990 2517 2996 2518
rect 2990 2513 2991 2517
rect 2995 2513 2996 2517
rect 2990 2512 2996 2513
rect 3110 2517 3116 2518
rect 3110 2513 3111 2517
rect 3115 2513 3116 2517
rect 3110 2512 3116 2513
rect 3230 2517 3236 2518
rect 3230 2513 3231 2517
rect 3235 2513 3236 2517
rect 3230 2512 3236 2513
rect 3358 2517 3364 2518
rect 3358 2513 3359 2517
rect 3363 2513 3364 2517
rect 3358 2512 3364 2513
rect 3486 2517 3492 2518
rect 3486 2513 3487 2517
rect 3491 2513 3492 2517
rect 3486 2512 3492 2513
rect 3942 2516 3948 2517
rect 3942 2512 3943 2516
rect 3947 2512 3948 2516
rect 2046 2511 2052 2512
rect 3942 2511 3948 2512
rect 134 2464 140 2465
rect 110 2461 116 2462
rect 110 2457 111 2461
rect 115 2457 116 2461
rect 134 2460 135 2464
rect 139 2460 140 2464
rect 134 2459 140 2460
rect 230 2464 236 2465
rect 230 2460 231 2464
rect 235 2460 236 2464
rect 230 2459 236 2460
rect 326 2464 332 2465
rect 326 2460 327 2464
rect 331 2460 332 2464
rect 326 2459 332 2460
rect 422 2464 428 2465
rect 422 2460 423 2464
rect 427 2460 428 2464
rect 422 2459 428 2460
rect 518 2464 524 2465
rect 518 2460 519 2464
rect 523 2460 524 2464
rect 518 2459 524 2460
rect 2006 2461 2012 2462
rect 110 2456 116 2457
rect 2006 2457 2007 2461
rect 2011 2457 2012 2461
rect 2006 2456 2012 2457
rect 2046 2460 2052 2461
rect 3942 2460 3948 2461
rect 2046 2456 2047 2460
rect 2051 2456 2052 2460
rect 2046 2455 2052 2456
rect 2534 2459 2540 2460
rect 2534 2455 2535 2459
rect 2539 2455 2540 2459
rect 2534 2454 2540 2455
rect 2710 2459 2716 2460
rect 2710 2455 2711 2459
rect 2715 2455 2716 2459
rect 2710 2454 2716 2455
rect 2878 2459 2884 2460
rect 2878 2455 2879 2459
rect 2883 2455 2884 2459
rect 2878 2454 2884 2455
rect 3046 2459 3052 2460
rect 3046 2455 3047 2459
rect 3051 2455 3052 2459
rect 3046 2454 3052 2455
rect 3206 2459 3212 2460
rect 3206 2455 3207 2459
rect 3211 2455 3212 2459
rect 3206 2454 3212 2455
rect 3358 2459 3364 2460
rect 3358 2455 3359 2459
rect 3363 2455 3364 2459
rect 3358 2454 3364 2455
rect 3502 2459 3508 2460
rect 3502 2455 3503 2459
rect 3507 2455 3508 2459
rect 3502 2454 3508 2455
rect 3654 2459 3660 2460
rect 3654 2455 3655 2459
rect 3659 2455 3660 2459
rect 3654 2454 3660 2455
rect 3806 2459 3812 2460
rect 3806 2455 3807 2459
rect 3811 2455 3812 2459
rect 3942 2456 3943 2460
rect 3947 2456 3948 2460
rect 3942 2455 3948 2456
rect 3806 2454 3812 2455
rect 134 2445 140 2446
rect 110 2444 116 2445
rect 110 2440 111 2444
rect 115 2440 116 2444
rect 134 2441 135 2445
rect 139 2441 140 2445
rect 134 2440 140 2441
rect 230 2445 236 2446
rect 230 2441 231 2445
rect 235 2441 236 2445
rect 230 2440 236 2441
rect 326 2445 332 2446
rect 326 2441 327 2445
rect 331 2441 332 2445
rect 326 2440 332 2441
rect 422 2445 428 2446
rect 422 2441 423 2445
rect 427 2441 428 2445
rect 422 2440 428 2441
rect 518 2445 524 2446
rect 518 2441 519 2445
rect 523 2441 524 2445
rect 518 2440 524 2441
rect 2006 2444 2012 2445
rect 2006 2440 2007 2444
rect 2011 2440 2012 2444
rect 110 2439 116 2440
rect 2006 2439 2012 2440
rect 2046 2443 2052 2444
rect 2046 2439 2047 2443
rect 2051 2439 2052 2443
rect 3942 2443 3948 2444
rect 2046 2438 2052 2439
rect 2534 2440 2540 2441
rect 2534 2436 2535 2440
rect 2539 2436 2540 2440
rect 2534 2435 2540 2436
rect 2710 2440 2716 2441
rect 2710 2436 2711 2440
rect 2715 2436 2716 2440
rect 2710 2435 2716 2436
rect 2878 2440 2884 2441
rect 2878 2436 2879 2440
rect 2883 2436 2884 2440
rect 2878 2435 2884 2436
rect 3046 2440 3052 2441
rect 3046 2436 3047 2440
rect 3051 2436 3052 2440
rect 3046 2435 3052 2436
rect 3206 2440 3212 2441
rect 3206 2436 3207 2440
rect 3211 2436 3212 2440
rect 3206 2435 3212 2436
rect 3358 2440 3364 2441
rect 3358 2436 3359 2440
rect 3363 2436 3364 2440
rect 3358 2435 3364 2436
rect 3502 2440 3508 2441
rect 3502 2436 3503 2440
rect 3507 2436 3508 2440
rect 3502 2435 3508 2436
rect 3654 2440 3660 2441
rect 3654 2436 3655 2440
rect 3659 2436 3660 2440
rect 3654 2435 3660 2436
rect 3806 2440 3812 2441
rect 3806 2436 3807 2440
rect 3811 2436 3812 2440
rect 3942 2439 3943 2443
rect 3947 2439 3948 2443
rect 3942 2438 3948 2439
rect 3806 2435 3812 2436
rect 110 2376 116 2377
rect 2006 2376 2012 2377
rect 110 2372 111 2376
rect 115 2372 116 2376
rect 110 2371 116 2372
rect 134 2375 140 2376
rect 134 2371 135 2375
rect 139 2371 140 2375
rect 134 2370 140 2371
rect 254 2375 260 2376
rect 254 2371 255 2375
rect 259 2371 260 2375
rect 254 2370 260 2371
rect 414 2375 420 2376
rect 414 2371 415 2375
rect 419 2371 420 2375
rect 414 2370 420 2371
rect 574 2375 580 2376
rect 574 2371 575 2375
rect 579 2371 580 2375
rect 574 2370 580 2371
rect 734 2375 740 2376
rect 734 2371 735 2375
rect 739 2371 740 2375
rect 734 2370 740 2371
rect 886 2375 892 2376
rect 886 2371 887 2375
rect 891 2371 892 2375
rect 886 2370 892 2371
rect 1038 2375 1044 2376
rect 1038 2371 1039 2375
rect 1043 2371 1044 2375
rect 1038 2370 1044 2371
rect 1182 2375 1188 2376
rect 1182 2371 1183 2375
rect 1187 2371 1188 2375
rect 1182 2370 1188 2371
rect 1326 2375 1332 2376
rect 1326 2371 1327 2375
rect 1331 2371 1332 2375
rect 1326 2370 1332 2371
rect 1478 2375 1484 2376
rect 1478 2371 1479 2375
rect 1483 2371 1484 2375
rect 2006 2372 2007 2376
rect 2011 2372 2012 2376
rect 2006 2371 2012 2372
rect 1478 2370 1484 2371
rect 2606 2368 2612 2369
rect 2046 2365 2052 2366
rect 2046 2361 2047 2365
rect 2051 2361 2052 2365
rect 2606 2364 2607 2368
rect 2611 2364 2612 2368
rect 2606 2363 2612 2364
rect 2814 2368 2820 2369
rect 2814 2364 2815 2368
rect 2819 2364 2820 2368
rect 2814 2363 2820 2364
rect 3006 2368 3012 2369
rect 3006 2364 3007 2368
rect 3011 2364 3012 2368
rect 3006 2363 3012 2364
rect 3190 2368 3196 2369
rect 3190 2364 3191 2368
rect 3195 2364 3196 2368
rect 3190 2363 3196 2364
rect 3358 2368 3364 2369
rect 3358 2364 3359 2368
rect 3363 2364 3364 2368
rect 3358 2363 3364 2364
rect 3518 2368 3524 2369
rect 3518 2364 3519 2368
rect 3523 2364 3524 2368
rect 3518 2363 3524 2364
rect 3678 2368 3684 2369
rect 3678 2364 3679 2368
rect 3683 2364 3684 2368
rect 3678 2363 3684 2364
rect 3838 2368 3844 2369
rect 3838 2364 3839 2368
rect 3843 2364 3844 2368
rect 3838 2363 3844 2364
rect 3942 2365 3948 2366
rect 2046 2360 2052 2361
rect 3942 2361 3943 2365
rect 3947 2361 3948 2365
rect 3942 2360 3948 2361
rect 110 2359 116 2360
rect 110 2355 111 2359
rect 115 2355 116 2359
rect 2006 2359 2012 2360
rect 110 2354 116 2355
rect 134 2356 140 2357
rect 134 2352 135 2356
rect 139 2352 140 2356
rect 134 2351 140 2352
rect 254 2356 260 2357
rect 254 2352 255 2356
rect 259 2352 260 2356
rect 254 2351 260 2352
rect 414 2356 420 2357
rect 414 2352 415 2356
rect 419 2352 420 2356
rect 414 2351 420 2352
rect 574 2356 580 2357
rect 574 2352 575 2356
rect 579 2352 580 2356
rect 574 2351 580 2352
rect 734 2356 740 2357
rect 734 2352 735 2356
rect 739 2352 740 2356
rect 734 2351 740 2352
rect 886 2356 892 2357
rect 886 2352 887 2356
rect 891 2352 892 2356
rect 886 2351 892 2352
rect 1038 2356 1044 2357
rect 1038 2352 1039 2356
rect 1043 2352 1044 2356
rect 1038 2351 1044 2352
rect 1182 2356 1188 2357
rect 1182 2352 1183 2356
rect 1187 2352 1188 2356
rect 1182 2351 1188 2352
rect 1326 2356 1332 2357
rect 1326 2352 1327 2356
rect 1331 2352 1332 2356
rect 1326 2351 1332 2352
rect 1478 2356 1484 2357
rect 1478 2352 1479 2356
rect 1483 2352 1484 2356
rect 2006 2355 2007 2359
rect 2011 2355 2012 2359
rect 2006 2354 2012 2355
rect 1478 2351 1484 2352
rect 2606 2349 2612 2350
rect 2046 2348 2052 2349
rect 2046 2344 2047 2348
rect 2051 2344 2052 2348
rect 2606 2345 2607 2349
rect 2611 2345 2612 2349
rect 2606 2344 2612 2345
rect 2814 2349 2820 2350
rect 2814 2345 2815 2349
rect 2819 2345 2820 2349
rect 2814 2344 2820 2345
rect 3006 2349 3012 2350
rect 3006 2345 3007 2349
rect 3011 2345 3012 2349
rect 3006 2344 3012 2345
rect 3190 2349 3196 2350
rect 3190 2345 3191 2349
rect 3195 2345 3196 2349
rect 3190 2344 3196 2345
rect 3358 2349 3364 2350
rect 3358 2345 3359 2349
rect 3363 2345 3364 2349
rect 3358 2344 3364 2345
rect 3518 2349 3524 2350
rect 3518 2345 3519 2349
rect 3523 2345 3524 2349
rect 3518 2344 3524 2345
rect 3678 2349 3684 2350
rect 3678 2345 3679 2349
rect 3683 2345 3684 2349
rect 3678 2344 3684 2345
rect 3838 2349 3844 2350
rect 3838 2345 3839 2349
rect 3843 2345 3844 2349
rect 3838 2344 3844 2345
rect 3942 2348 3948 2349
rect 3942 2344 3943 2348
rect 3947 2344 3948 2348
rect 2046 2343 2052 2344
rect 3942 2343 3948 2344
rect 134 2296 140 2297
rect 110 2293 116 2294
rect 110 2289 111 2293
rect 115 2289 116 2293
rect 134 2292 135 2296
rect 139 2292 140 2296
rect 134 2291 140 2292
rect 262 2296 268 2297
rect 262 2292 263 2296
rect 267 2292 268 2296
rect 262 2291 268 2292
rect 422 2296 428 2297
rect 422 2292 423 2296
rect 427 2292 428 2296
rect 422 2291 428 2292
rect 582 2296 588 2297
rect 582 2292 583 2296
rect 587 2292 588 2296
rect 582 2291 588 2292
rect 742 2296 748 2297
rect 742 2292 743 2296
rect 747 2292 748 2296
rect 742 2291 748 2292
rect 894 2296 900 2297
rect 894 2292 895 2296
rect 899 2292 900 2296
rect 894 2291 900 2292
rect 1046 2296 1052 2297
rect 1046 2292 1047 2296
rect 1051 2292 1052 2296
rect 1046 2291 1052 2292
rect 1198 2296 1204 2297
rect 1198 2292 1199 2296
rect 1203 2292 1204 2296
rect 1198 2291 1204 2292
rect 1350 2296 1356 2297
rect 1350 2292 1351 2296
rect 1355 2292 1356 2296
rect 1350 2291 1356 2292
rect 1502 2296 1508 2297
rect 1502 2292 1503 2296
rect 1507 2292 1508 2296
rect 1502 2291 1508 2292
rect 2006 2293 2012 2294
rect 110 2288 116 2289
rect 2006 2289 2007 2293
rect 2011 2289 2012 2293
rect 2006 2288 2012 2289
rect 2046 2280 2052 2281
rect 3942 2280 3948 2281
rect 134 2277 140 2278
rect 110 2276 116 2277
rect 110 2272 111 2276
rect 115 2272 116 2276
rect 134 2273 135 2277
rect 139 2273 140 2277
rect 134 2272 140 2273
rect 262 2277 268 2278
rect 262 2273 263 2277
rect 267 2273 268 2277
rect 262 2272 268 2273
rect 422 2277 428 2278
rect 422 2273 423 2277
rect 427 2273 428 2277
rect 422 2272 428 2273
rect 582 2277 588 2278
rect 582 2273 583 2277
rect 587 2273 588 2277
rect 582 2272 588 2273
rect 742 2277 748 2278
rect 742 2273 743 2277
rect 747 2273 748 2277
rect 742 2272 748 2273
rect 894 2277 900 2278
rect 894 2273 895 2277
rect 899 2273 900 2277
rect 894 2272 900 2273
rect 1046 2277 1052 2278
rect 1046 2273 1047 2277
rect 1051 2273 1052 2277
rect 1046 2272 1052 2273
rect 1198 2277 1204 2278
rect 1198 2273 1199 2277
rect 1203 2273 1204 2277
rect 1198 2272 1204 2273
rect 1350 2277 1356 2278
rect 1350 2273 1351 2277
rect 1355 2273 1356 2277
rect 1350 2272 1356 2273
rect 1502 2277 1508 2278
rect 1502 2273 1503 2277
rect 1507 2273 1508 2277
rect 1502 2272 1508 2273
rect 2006 2276 2012 2277
rect 2006 2272 2007 2276
rect 2011 2272 2012 2276
rect 2046 2276 2047 2280
rect 2051 2276 2052 2280
rect 2046 2275 2052 2276
rect 2070 2279 2076 2280
rect 2070 2275 2071 2279
rect 2075 2275 2076 2279
rect 2070 2274 2076 2275
rect 2166 2279 2172 2280
rect 2166 2275 2167 2279
rect 2171 2275 2172 2279
rect 2166 2274 2172 2275
rect 2270 2279 2276 2280
rect 2270 2275 2271 2279
rect 2275 2275 2276 2279
rect 2270 2274 2276 2275
rect 2414 2279 2420 2280
rect 2414 2275 2415 2279
rect 2419 2275 2420 2279
rect 2414 2274 2420 2275
rect 2574 2279 2580 2280
rect 2574 2275 2575 2279
rect 2579 2275 2580 2279
rect 2574 2274 2580 2275
rect 2742 2279 2748 2280
rect 2742 2275 2743 2279
rect 2747 2275 2748 2279
rect 2742 2274 2748 2275
rect 2910 2279 2916 2280
rect 2910 2275 2911 2279
rect 2915 2275 2916 2279
rect 2910 2274 2916 2275
rect 3070 2279 3076 2280
rect 3070 2275 3071 2279
rect 3075 2275 3076 2279
rect 3070 2274 3076 2275
rect 3230 2279 3236 2280
rect 3230 2275 3231 2279
rect 3235 2275 3236 2279
rect 3230 2274 3236 2275
rect 3382 2279 3388 2280
rect 3382 2275 3383 2279
rect 3387 2275 3388 2279
rect 3382 2274 3388 2275
rect 3534 2279 3540 2280
rect 3534 2275 3535 2279
rect 3539 2275 3540 2279
rect 3534 2274 3540 2275
rect 3694 2279 3700 2280
rect 3694 2275 3695 2279
rect 3699 2275 3700 2279
rect 3942 2276 3943 2280
rect 3947 2276 3948 2280
rect 3942 2275 3948 2276
rect 3694 2274 3700 2275
rect 110 2271 116 2272
rect 2006 2271 2012 2272
rect 2046 2263 2052 2264
rect 2046 2259 2047 2263
rect 2051 2259 2052 2263
rect 3942 2263 3948 2264
rect 2046 2258 2052 2259
rect 2070 2260 2076 2261
rect 2070 2256 2071 2260
rect 2075 2256 2076 2260
rect 2070 2255 2076 2256
rect 2166 2260 2172 2261
rect 2166 2256 2167 2260
rect 2171 2256 2172 2260
rect 2166 2255 2172 2256
rect 2270 2260 2276 2261
rect 2270 2256 2271 2260
rect 2275 2256 2276 2260
rect 2270 2255 2276 2256
rect 2414 2260 2420 2261
rect 2414 2256 2415 2260
rect 2419 2256 2420 2260
rect 2414 2255 2420 2256
rect 2574 2260 2580 2261
rect 2574 2256 2575 2260
rect 2579 2256 2580 2260
rect 2574 2255 2580 2256
rect 2742 2260 2748 2261
rect 2742 2256 2743 2260
rect 2747 2256 2748 2260
rect 2742 2255 2748 2256
rect 2910 2260 2916 2261
rect 2910 2256 2911 2260
rect 2915 2256 2916 2260
rect 2910 2255 2916 2256
rect 3070 2260 3076 2261
rect 3070 2256 3071 2260
rect 3075 2256 3076 2260
rect 3070 2255 3076 2256
rect 3230 2260 3236 2261
rect 3230 2256 3231 2260
rect 3235 2256 3236 2260
rect 3230 2255 3236 2256
rect 3382 2260 3388 2261
rect 3382 2256 3383 2260
rect 3387 2256 3388 2260
rect 3382 2255 3388 2256
rect 3534 2260 3540 2261
rect 3534 2256 3535 2260
rect 3539 2256 3540 2260
rect 3534 2255 3540 2256
rect 3694 2260 3700 2261
rect 3694 2256 3695 2260
rect 3699 2256 3700 2260
rect 3942 2259 3943 2263
rect 3947 2259 3948 2263
rect 3942 2258 3948 2259
rect 3694 2255 3700 2256
rect 110 2220 116 2221
rect 2006 2220 2012 2221
rect 110 2216 111 2220
rect 115 2216 116 2220
rect 110 2215 116 2216
rect 222 2219 228 2220
rect 222 2215 223 2219
rect 227 2215 228 2219
rect 222 2214 228 2215
rect 350 2219 356 2220
rect 350 2215 351 2219
rect 355 2215 356 2219
rect 350 2214 356 2215
rect 494 2219 500 2220
rect 494 2215 495 2219
rect 499 2215 500 2219
rect 494 2214 500 2215
rect 646 2219 652 2220
rect 646 2215 647 2219
rect 651 2215 652 2219
rect 646 2214 652 2215
rect 798 2219 804 2220
rect 798 2215 799 2219
rect 803 2215 804 2219
rect 798 2214 804 2215
rect 958 2219 964 2220
rect 958 2215 959 2219
rect 963 2215 964 2219
rect 958 2214 964 2215
rect 1118 2219 1124 2220
rect 1118 2215 1119 2219
rect 1123 2215 1124 2219
rect 1118 2214 1124 2215
rect 1278 2219 1284 2220
rect 1278 2215 1279 2219
rect 1283 2215 1284 2219
rect 1278 2214 1284 2215
rect 1438 2219 1444 2220
rect 1438 2215 1439 2219
rect 1443 2215 1444 2219
rect 1438 2214 1444 2215
rect 1598 2219 1604 2220
rect 1598 2215 1599 2219
rect 1603 2215 1604 2219
rect 2006 2216 2007 2220
rect 2011 2216 2012 2220
rect 2006 2215 2012 2216
rect 1598 2214 1604 2215
rect 110 2203 116 2204
rect 110 2199 111 2203
rect 115 2199 116 2203
rect 2006 2203 2012 2204
rect 110 2198 116 2199
rect 222 2200 228 2201
rect 222 2196 223 2200
rect 227 2196 228 2200
rect 222 2195 228 2196
rect 350 2200 356 2201
rect 350 2196 351 2200
rect 355 2196 356 2200
rect 350 2195 356 2196
rect 494 2200 500 2201
rect 494 2196 495 2200
rect 499 2196 500 2200
rect 494 2195 500 2196
rect 646 2200 652 2201
rect 646 2196 647 2200
rect 651 2196 652 2200
rect 646 2195 652 2196
rect 798 2200 804 2201
rect 798 2196 799 2200
rect 803 2196 804 2200
rect 798 2195 804 2196
rect 958 2200 964 2201
rect 958 2196 959 2200
rect 963 2196 964 2200
rect 958 2195 964 2196
rect 1118 2200 1124 2201
rect 1118 2196 1119 2200
rect 1123 2196 1124 2200
rect 1118 2195 1124 2196
rect 1278 2200 1284 2201
rect 1278 2196 1279 2200
rect 1283 2196 1284 2200
rect 1278 2195 1284 2196
rect 1438 2200 1444 2201
rect 1438 2196 1439 2200
rect 1443 2196 1444 2200
rect 1438 2195 1444 2196
rect 1598 2200 1604 2201
rect 1598 2196 1599 2200
rect 1603 2196 1604 2200
rect 2006 2199 2007 2203
rect 2011 2199 2012 2203
rect 2006 2198 2012 2199
rect 2070 2200 2076 2201
rect 1598 2195 1604 2196
rect 2046 2197 2052 2198
rect 2046 2193 2047 2197
rect 2051 2193 2052 2197
rect 2070 2196 2071 2200
rect 2075 2196 2076 2200
rect 2070 2195 2076 2196
rect 2174 2200 2180 2201
rect 2174 2196 2175 2200
rect 2179 2196 2180 2200
rect 2174 2195 2180 2196
rect 2318 2200 2324 2201
rect 2318 2196 2319 2200
rect 2323 2196 2324 2200
rect 2318 2195 2324 2196
rect 2470 2200 2476 2201
rect 2470 2196 2471 2200
rect 2475 2196 2476 2200
rect 2470 2195 2476 2196
rect 2622 2200 2628 2201
rect 2622 2196 2623 2200
rect 2627 2196 2628 2200
rect 2622 2195 2628 2196
rect 2782 2200 2788 2201
rect 2782 2196 2783 2200
rect 2787 2196 2788 2200
rect 2782 2195 2788 2196
rect 2934 2200 2940 2201
rect 2934 2196 2935 2200
rect 2939 2196 2940 2200
rect 2934 2195 2940 2196
rect 3078 2200 3084 2201
rect 3078 2196 3079 2200
rect 3083 2196 3084 2200
rect 3078 2195 3084 2196
rect 3222 2200 3228 2201
rect 3222 2196 3223 2200
rect 3227 2196 3228 2200
rect 3222 2195 3228 2196
rect 3366 2200 3372 2201
rect 3366 2196 3367 2200
rect 3371 2196 3372 2200
rect 3366 2195 3372 2196
rect 3518 2200 3524 2201
rect 3518 2196 3519 2200
rect 3523 2196 3524 2200
rect 3518 2195 3524 2196
rect 3942 2197 3948 2198
rect 2046 2192 2052 2193
rect 3942 2193 3943 2197
rect 3947 2193 3948 2197
rect 3942 2192 3948 2193
rect 2070 2181 2076 2182
rect 2046 2180 2052 2181
rect 2046 2176 2047 2180
rect 2051 2176 2052 2180
rect 2070 2177 2071 2181
rect 2075 2177 2076 2181
rect 2070 2176 2076 2177
rect 2174 2181 2180 2182
rect 2174 2177 2175 2181
rect 2179 2177 2180 2181
rect 2174 2176 2180 2177
rect 2318 2181 2324 2182
rect 2318 2177 2319 2181
rect 2323 2177 2324 2181
rect 2318 2176 2324 2177
rect 2470 2181 2476 2182
rect 2470 2177 2471 2181
rect 2475 2177 2476 2181
rect 2470 2176 2476 2177
rect 2622 2181 2628 2182
rect 2622 2177 2623 2181
rect 2627 2177 2628 2181
rect 2622 2176 2628 2177
rect 2782 2181 2788 2182
rect 2782 2177 2783 2181
rect 2787 2177 2788 2181
rect 2782 2176 2788 2177
rect 2934 2181 2940 2182
rect 2934 2177 2935 2181
rect 2939 2177 2940 2181
rect 2934 2176 2940 2177
rect 3078 2181 3084 2182
rect 3078 2177 3079 2181
rect 3083 2177 3084 2181
rect 3078 2176 3084 2177
rect 3222 2181 3228 2182
rect 3222 2177 3223 2181
rect 3227 2177 3228 2181
rect 3222 2176 3228 2177
rect 3366 2181 3372 2182
rect 3366 2177 3367 2181
rect 3371 2177 3372 2181
rect 3366 2176 3372 2177
rect 3518 2181 3524 2182
rect 3518 2177 3519 2181
rect 3523 2177 3524 2181
rect 3518 2176 3524 2177
rect 3942 2180 3948 2181
rect 3942 2176 3943 2180
rect 3947 2176 3948 2180
rect 2046 2175 2052 2176
rect 3942 2175 3948 2176
rect 470 2140 476 2141
rect 110 2137 116 2138
rect 110 2133 111 2137
rect 115 2133 116 2137
rect 470 2136 471 2140
rect 475 2136 476 2140
rect 470 2135 476 2136
rect 566 2140 572 2141
rect 566 2136 567 2140
rect 571 2136 572 2140
rect 566 2135 572 2136
rect 678 2140 684 2141
rect 678 2136 679 2140
rect 683 2136 684 2140
rect 678 2135 684 2136
rect 806 2140 812 2141
rect 806 2136 807 2140
rect 811 2136 812 2140
rect 806 2135 812 2136
rect 942 2140 948 2141
rect 942 2136 943 2140
rect 947 2136 948 2140
rect 942 2135 948 2136
rect 1078 2140 1084 2141
rect 1078 2136 1079 2140
rect 1083 2136 1084 2140
rect 1078 2135 1084 2136
rect 1222 2140 1228 2141
rect 1222 2136 1223 2140
rect 1227 2136 1228 2140
rect 1222 2135 1228 2136
rect 1366 2140 1372 2141
rect 1366 2136 1367 2140
rect 1371 2136 1372 2140
rect 1366 2135 1372 2136
rect 1502 2140 1508 2141
rect 1502 2136 1503 2140
rect 1507 2136 1508 2140
rect 1502 2135 1508 2136
rect 1638 2140 1644 2141
rect 1638 2136 1639 2140
rect 1643 2136 1644 2140
rect 1638 2135 1644 2136
rect 1782 2140 1788 2141
rect 1782 2136 1783 2140
rect 1787 2136 1788 2140
rect 1782 2135 1788 2136
rect 1902 2140 1908 2141
rect 1902 2136 1903 2140
rect 1907 2136 1908 2140
rect 1902 2135 1908 2136
rect 2006 2137 2012 2138
rect 110 2132 116 2133
rect 2006 2133 2007 2137
rect 2011 2133 2012 2137
rect 2006 2132 2012 2133
rect 470 2121 476 2122
rect 110 2120 116 2121
rect 110 2116 111 2120
rect 115 2116 116 2120
rect 470 2117 471 2121
rect 475 2117 476 2121
rect 470 2116 476 2117
rect 566 2121 572 2122
rect 566 2117 567 2121
rect 571 2117 572 2121
rect 566 2116 572 2117
rect 678 2121 684 2122
rect 678 2117 679 2121
rect 683 2117 684 2121
rect 678 2116 684 2117
rect 806 2121 812 2122
rect 806 2117 807 2121
rect 811 2117 812 2121
rect 806 2116 812 2117
rect 942 2121 948 2122
rect 942 2117 943 2121
rect 947 2117 948 2121
rect 942 2116 948 2117
rect 1078 2121 1084 2122
rect 1078 2117 1079 2121
rect 1083 2117 1084 2121
rect 1078 2116 1084 2117
rect 1222 2121 1228 2122
rect 1222 2117 1223 2121
rect 1227 2117 1228 2121
rect 1222 2116 1228 2117
rect 1366 2121 1372 2122
rect 1366 2117 1367 2121
rect 1371 2117 1372 2121
rect 1366 2116 1372 2117
rect 1502 2121 1508 2122
rect 1502 2117 1503 2121
rect 1507 2117 1508 2121
rect 1502 2116 1508 2117
rect 1638 2121 1644 2122
rect 1638 2117 1639 2121
rect 1643 2117 1644 2121
rect 1638 2116 1644 2117
rect 1782 2121 1788 2122
rect 1782 2117 1783 2121
rect 1787 2117 1788 2121
rect 1782 2116 1788 2117
rect 1902 2121 1908 2122
rect 1902 2117 1903 2121
rect 1907 2117 1908 2121
rect 1902 2116 1908 2117
rect 2006 2120 2012 2121
rect 2006 2116 2007 2120
rect 2011 2116 2012 2120
rect 110 2115 116 2116
rect 2006 2115 2012 2116
rect 2046 2108 2052 2109
rect 3942 2108 3948 2109
rect 2046 2104 2047 2108
rect 2051 2104 2052 2108
rect 2046 2103 2052 2104
rect 2278 2107 2284 2108
rect 2278 2103 2279 2107
rect 2283 2103 2284 2107
rect 2278 2102 2284 2103
rect 2390 2107 2396 2108
rect 2390 2103 2391 2107
rect 2395 2103 2396 2107
rect 2390 2102 2396 2103
rect 2510 2107 2516 2108
rect 2510 2103 2511 2107
rect 2515 2103 2516 2107
rect 2510 2102 2516 2103
rect 2630 2107 2636 2108
rect 2630 2103 2631 2107
rect 2635 2103 2636 2107
rect 2630 2102 2636 2103
rect 2758 2107 2764 2108
rect 2758 2103 2759 2107
rect 2763 2103 2764 2107
rect 2758 2102 2764 2103
rect 2894 2107 2900 2108
rect 2894 2103 2895 2107
rect 2899 2103 2900 2107
rect 2894 2102 2900 2103
rect 3038 2107 3044 2108
rect 3038 2103 3039 2107
rect 3043 2103 3044 2107
rect 3038 2102 3044 2103
rect 3190 2107 3196 2108
rect 3190 2103 3191 2107
rect 3195 2103 3196 2107
rect 3190 2102 3196 2103
rect 3350 2107 3356 2108
rect 3350 2103 3351 2107
rect 3355 2103 3356 2107
rect 3350 2102 3356 2103
rect 3518 2107 3524 2108
rect 3518 2103 3519 2107
rect 3523 2103 3524 2107
rect 3518 2102 3524 2103
rect 3686 2107 3692 2108
rect 3686 2103 3687 2107
rect 3691 2103 3692 2107
rect 3686 2102 3692 2103
rect 3838 2107 3844 2108
rect 3838 2103 3839 2107
rect 3843 2103 3844 2107
rect 3942 2104 3943 2108
rect 3947 2104 3948 2108
rect 3942 2103 3948 2104
rect 3838 2102 3844 2103
rect 2046 2091 2052 2092
rect 2046 2087 2047 2091
rect 2051 2087 2052 2091
rect 3942 2091 3948 2092
rect 2046 2086 2052 2087
rect 2278 2088 2284 2089
rect 2278 2084 2279 2088
rect 2283 2084 2284 2088
rect 2278 2083 2284 2084
rect 2390 2088 2396 2089
rect 2390 2084 2391 2088
rect 2395 2084 2396 2088
rect 2390 2083 2396 2084
rect 2510 2088 2516 2089
rect 2510 2084 2511 2088
rect 2515 2084 2516 2088
rect 2510 2083 2516 2084
rect 2630 2088 2636 2089
rect 2630 2084 2631 2088
rect 2635 2084 2636 2088
rect 2630 2083 2636 2084
rect 2758 2088 2764 2089
rect 2758 2084 2759 2088
rect 2763 2084 2764 2088
rect 2758 2083 2764 2084
rect 2894 2088 2900 2089
rect 2894 2084 2895 2088
rect 2899 2084 2900 2088
rect 2894 2083 2900 2084
rect 3038 2088 3044 2089
rect 3038 2084 3039 2088
rect 3043 2084 3044 2088
rect 3038 2083 3044 2084
rect 3190 2088 3196 2089
rect 3190 2084 3191 2088
rect 3195 2084 3196 2088
rect 3190 2083 3196 2084
rect 3350 2088 3356 2089
rect 3350 2084 3351 2088
rect 3355 2084 3356 2088
rect 3350 2083 3356 2084
rect 3518 2088 3524 2089
rect 3518 2084 3519 2088
rect 3523 2084 3524 2088
rect 3518 2083 3524 2084
rect 3686 2088 3692 2089
rect 3686 2084 3687 2088
rect 3691 2084 3692 2088
rect 3686 2083 3692 2084
rect 3838 2088 3844 2089
rect 3838 2084 3839 2088
rect 3843 2084 3844 2088
rect 3942 2087 3943 2091
rect 3947 2087 3948 2091
rect 3942 2086 3948 2087
rect 3838 2083 3844 2084
rect 110 2068 116 2069
rect 2006 2068 2012 2069
rect 110 2064 111 2068
rect 115 2064 116 2068
rect 110 2063 116 2064
rect 622 2067 628 2068
rect 622 2063 623 2067
rect 627 2063 628 2067
rect 622 2062 628 2063
rect 734 2067 740 2068
rect 734 2063 735 2067
rect 739 2063 740 2067
rect 734 2062 740 2063
rect 854 2067 860 2068
rect 854 2063 855 2067
rect 859 2063 860 2067
rect 854 2062 860 2063
rect 982 2067 988 2068
rect 982 2063 983 2067
rect 987 2063 988 2067
rect 982 2062 988 2063
rect 1118 2067 1124 2068
rect 1118 2063 1119 2067
rect 1123 2063 1124 2067
rect 1118 2062 1124 2063
rect 1254 2067 1260 2068
rect 1254 2063 1255 2067
rect 1259 2063 1260 2067
rect 1254 2062 1260 2063
rect 1390 2067 1396 2068
rect 1390 2063 1391 2067
rect 1395 2063 1396 2067
rect 1390 2062 1396 2063
rect 1526 2067 1532 2068
rect 1526 2063 1527 2067
rect 1531 2063 1532 2067
rect 1526 2062 1532 2063
rect 1654 2067 1660 2068
rect 1654 2063 1655 2067
rect 1659 2063 1660 2067
rect 1654 2062 1660 2063
rect 1790 2067 1796 2068
rect 1790 2063 1791 2067
rect 1795 2063 1796 2067
rect 1790 2062 1796 2063
rect 1902 2067 1908 2068
rect 1902 2063 1903 2067
rect 1907 2063 1908 2067
rect 2006 2064 2007 2068
rect 2011 2064 2012 2068
rect 2006 2063 2012 2064
rect 1902 2062 1908 2063
rect 110 2051 116 2052
rect 110 2047 111 2051
rect 115 2047 116 2051
rect 2006 2051 2012 2052
rect 110 2046 116 2047
rect 622 2048 628 2049
rect 622 2044 623 2048
rect 627 2044 628 2048
rect 622 2043 628 2044
rect 734 2048 740 2049
rect 734 2044 735 2048
rect 739 2044 740 2048
rect 734 2043 740 2044
rect 854 2048 860 2049
rect 854 2044 855 2048
rect 859 2044 860 2048
rect 854 2043 860 2044
rect 982 2048 988 2049
rect 982 2044 983 2048
rect 987 2044 988 2048
rect 982 2043 988 2044
rect 1118 2048 1124 2049
rect 1118 2044 1119 2048
rect 1123 2044 1124 2048
rect 1118 2043 1124 2044
rect 1254 2048 1260 2049
rect 1254 2044 1255 2048
rect 1259 2044 1260 2048
rect 1254 2043 1260 2044
rect 1390 2048 1396 2049
rect 1390 2044 1391 2048
rect 1395 2044 1396 2048
rect 1390 2043 1396 2044
rect 1526 2048 1532 2049
rect 1526 2044 1527 2048
rect 1531 2044 1532 2048
rect 1526 2043 1532 2044
rect 1654 2048 1660 2049
rect 1654 2044 1655 2048
rect 1659 2044 1660 2048
rect 1654 2043 1660 2044
rect 1790 2048 1796 2049
rect 1790 2044 1791 2048
rect 1795 2044 1796 2048
rect 1790 2043 1796 2044
rect 1902 2048 1908 2049
rect 1902 2044 1903 2048
rect 1907 2044 1908 2048
rect 2006 2047 2007 2051
rect 2011 2047 2012 2051
rect 2006 2046 2012 2047
rect 1902 2043 1908 2044
rect 2326 2020 2332 2021
rect 2046 2017 2052 2018
rect 2046 2013 2047 2017
rect 2051 2013 2052 2017
rect 2326 2016 2327 2020
rect 2331 2016 2332 2020
rect 2326 2015 2332 2016
rect 2430 2020 2436 2021
rect 2430 2016 2431 2020
rect 2435 2016 2436 2020
rect 2430 2015 2436 2016
rect 2534 2020 2540 2021
rect 2534 2016 2535 2020
rect 2539 2016 2540 2020
rect 2534 2015 2540 2016
rect 2646 2020 2652 2021
rect 2646 2016 2647 2020
rect 2651 2016 2652 2020
rect 2646 2015 2652 2016
rect 2774 2020 2780 2021
rect 2774 2016 2775 2020
rect 2779 2016 2780 2020
rect 2774 2015 2780 2016
rect 2918 2020 2924 2021
rect 2918 2016 2919 2020
rect 2923 2016 2924 2020
rect 2918 2015 2924 2016
rect 3078 2020 3084 2021
rect 3078 2016 3079 2020
rect 3083 2016 3084 2020
rect 3078 2015 3084 2016
rect 3262 2020 3268 2021
rect 3262 2016 3263 2020
rect 3267 2016 3268 2020
rect 3262 2015 3268 2016
rect 3454 2020 3460 2021
rect 3454 2016 3455 2020
rect 3459 2016 3460 2020
rect 3454 2015 3460 2016
rect 3654 2020 3660 2021
rect 3654 2016 3655 2020
rect 3659 2016 3660 2020
rect 3654 2015 3660 2016
rect 3838 2020 3844 2021
rect 3838 2016 3839 2020
rect 3843 2016 3844 2020
rect 3838 2015 3844 2016
rect 3942 2017 3948 2018
rect 2046 2012 2052 2013
rect 3942 2013 3943 2017
rect 3947 2013 3948 2017
rect 3942 2012 3948 2013
rect 2326 2001 2332 2002
rect 2046 2000 2052 2001
rect 2046 1996 2047 2000
rect 2051 1996 2052 2000
rect 2326 1997 2327 2001
rect 2331 1997 2332 2001
rect 2326 1996 2332 1997
rect 2430 2001 2436 2002
rect 2430 1997 2431 2001
rect 2435 1997 2436 2001
rect 2430 1996 2436 1997
rect 2534 2001 2540 2002
rect 2534 1997 2535 2001
rect 2539 1997 2540 2001
rect 2534 1996 2540 1997
rect 2646 2001 2652 2002
rect 2646 1997 2647 2001
rect 2651 1997 2652 2001
rect 2646 1996 2652 1997
rect 2774 2001 2780 2002
rect 2774 1997 2775 2001
rect 2779 1997 2780 2001
rect 2774 1996 2780 1997
rect 2918 2001 2924 2002
rect 2918 1997 2919 2001
rect 2923 1997 2924 2001
rect 2918 1996 2924 1997
rect 3078 2001 3084 2002
rect 3078 1997 3079 2001
rect 3083 1997 3084 2001
rect 3078 1996 3084 1997
rect 3262 2001 3268 2002
rect 3262 1997 3263 2001
rect 3267 1997 3268 2001
rect 3262 1996 3268 1997
rect 3454 2001 3460 2002
rect 3454 1997 3455 2001
rect 3459 1997 3460 2001
rect 3454 1996 3460 1997
rect 3654 2001 3660 2002
rect 3654 1997 3655 2001
rect 3659 1997 3660 2001
rect 3654 1996 3660 1997
rect 3838 2001 3844 2002
rect 3838 1997 3839 2001
rect 3843 1997 3844 2001
rect 3838 1996 3844 1997
rect 3942 2000 3948 2001
rect 3942 1996 3943 2000
rect 3947 1996 3948 2000
rect 2046 1995 2052 1996
rect 3942 1995 3948 1996
rect 446 1984 452 1985
rect 110 1981 116 1982
rect 110 1977 111 1981
rect 115 1977 116 1981
rect 446 1980 447 1984
rect 451 1980 452 1984
rect 446 1979 452 1980
rect 574 1984 580 1985
rect 574 1980 575 1984
rect 579 1980 580 1984
rect 574 1979 580 1980
rect 726 1984 732 1985
rect 726 1980 727 1984
rect 731 1980 732 1984
rect 726 1979 732 1980
rect 886 1984 892 1985
rect 886 1980 887 1984
rect 891 1980 892 1984
rect 886 1979 892 1980
rect 1054 1984 1060 1985
rect 1054 1980 1055 1984
rect 1059 1980 1060 1984
rect 1054 1979 1060 1980
rect 1230 1984 1236 1985
rect 1230 1980 1231 1984
rect 1235 1980 1236 1984
rect 1230 1979 1236 1980
rect 1398 1984 1404 1985
rect 1398 1980 1399 1984
rect 1403 1980 1404 1984
rect 1398 1979 1404 1980
rect 1574 1984 1580 1985
rect 1574 1980 1575 1984
rect 1579 1980 1580 1984
rect 1574 1979 1580 1980
rect 1750 1984 1756 1985
rect 1750 1980 1751 1984
rect 1755 1980 1756 1984
rect 1750 1979 1756 1980
rect 1902 1984 1908 1985
rect 1902 1980 1903 1984
rect 1907 1980 1908 1984
rect 1902 1979 1908 1980
rect 2006 1981 2012 1982
rect 110 1976 116 1977
rect 2006 1977 2007 1981
rect 2011 1977 2012 1981
rect 2006 1976 2012 1977
rect 446 1965 452 1966
rect 110 1964 116 1965
rect 110 1960 111 1964
rect 115 1960 116 1964
rect 446 1961 447 1965
rect 451 1961 452 1965
rect 446 1960 452 1961
rect 574 1965 580 1966
rect 574 1961 575 1965
rect 579 1961 580 1965
rect 574 1960 580 1961
rect 726 1965 732 1966
rect 726 1961 727 1965
rect 731 1961 732 1965
rect 726 1960 732 1961
rect 886 1965 892 1966
rect 886 1961 887 1965
rect 891 1961 892 1965
rect 886 1960 892 1961
rect 1054 1965 1060 1966
rect 1054 1961 1055 1965
rect 1059 1961 1060 1965
rect 1054 1960 1060 1961
rect 1230 1965 1236 1966
rect 1230 1961 1231 1965
rect 1235 1961 1236 1965
rect 1230 1960 1236 1961
rect 1398 1965 1404 1966
rect 1398 1961 1399 1965
rect 1403 1961 1404 1965
rect 1398 1960 1404 1961
rect 1574 1965 1580 1966
rect 1574 1961 1575 1965
rect 1579 1961 1580 1965
rect 1574 1960 1580 1961
rect 1750 1965 1756 1966
rect 1750 1961 1751 1965
rect 1755 1961 1756 1965
rect 1750 1960 1756 1961
rect 1902 1965 1908 1966
rect 1902 1961 1903 1965
rect 1907 1961 1908 1965
rect 1902 1960 1908 1961
rect 2006 1964 2012 1965
rect 2006 1960 2007 1964
rect 2011 1960 2012 1964
rect 110 1959 116 1960
rect 2006 1959 2012 1960
rect 2046 1944 2052 1945
rect 3942 1944 3948 1945
rect 2046 1940 2047 1944
rect 2051 1940 2052 1944
rect 2046 1939 2052 1940
rect 2254 1943 2260 1944
rect 2254 1939 2255 1943
rect 2259 1939 2260 1943
rect 2254 1938 2260 1939
rect 2350 1943 2356 1944
rect 2350 1939 2351 1943
rect 2355 1939 2356 1943
rect 2350 1938 2356 1939
rect 2446 1943 2452 1944
rect 2446 1939 2447 1943
rect 2451 1939 2452 1943
rect 2446 1938 2452 1939
rect 2542 1943 2548 1944
rect 2542 1939 2543 1943
rect 2547 1939 2548 1943
rect 2542 1938 2548 1939
rect 2646 1943 2652 1944
rect 2646 1939 2647 1943
rect 2651 1939 2652 1943
rect 2646 1938 2652 1939
rect 2766 1943 2772 1944
rect 2766 1939 2767 1943
rect 2771 1939 2772 1943
rect 2766 1938 2772 1939
rect 2918 1943 2924 1944
rect 2918 1939 2919 1943
rect 2923 1939 2924 1943
rect 2918 1938 2924 1939
rect 3102 1943 3108 1944
rect 3102 1939 3103 1943
rect 3107 1939 3108 1943
rect 3102 1938 3108 1939
rect 3318 1943 3324 1944
rect 3318 1939 3319 1943
rect 3323 1939 3324 1943
rect 3318 1938 3324 1939
rect 3542 1943 3548 1944
rect 3542 1939 3543 1943
rect 3547 1939 3548 1943
rect 3542 1938 3548 1939
rect 3774 1943 3780 1944
rect 3774 1939 3775 1943
rect 3779 1939 3780 1943
rect 3942 1940 3943 1944
rect 3947 1940 3948 1944
rect 3942 1939 3948 1940
rect 3774 1938 3780 1939
rect 2046 1927 2052 1928
rect 2046 1923 2047 1927
rect 2051 1923 2052 1927
rect 3942 1927 3948 1928
rect 2046 1922 2052 1923
rect 2254 1924 2260 1925
rect 2254 1920 2255 1924
rect 2259 1920 2260 1924
rect 2254 1919 2260 1920
rect 2350 1924 2356 1925
rect 2350 1920 2351 1924
rect 2355 1920 2356 1924
rect 2350 1919 2356 1920
rect 2446 1924 2452 1925
rect 2446 1920 2447 1924
rect 2451 1920 2452 1924
rect 2446 1919 2452 1920
rect 2542 1924 2548 1925
rect 2542 1920 2543 1924
rect 2547 1920 2548 1924
rect 2542 1919 2548 1920
rect 2646 1924 2652 1925
rect 2646 1920 2647 1924
rect 2651 1920 2652 1924
rect 2646 1919 2652 1920
rect 2766 1924 2772 1925
rect 2766 1920 2767 1924
rect 2771 1920 2772 1924
rect 2766 1919 2772 1920
rect 2918 1924 2924 1925
rect 2918 1920 2919 1924
rect 2923 1920 2924 1924
rect 2918 1919 2924 1920
rect 3102 1924 3108 1925
rect 3102 1920 3103 1924
rect 3107 1920 3108 1924
rect 3102 1919 3108 1920
rect 3318 1924 3324 1925
rect 3318 1920 3319 1924
rect 3323 1920 3324 1924
rect 3318 1919 3324 1920
rect 3542 1924 3548 1925
rect 3542 1920 3543 1924
rect 3547 1920 3548 1924
rect 3542 1919 3548 1920
rect 3774 1924 3780 1925
rect 3774 1920 3775 1924
rect 3779 1920 3780 1924
rect 3942 1923 3943 1927
rect 3947 1923 3948 1927
rect 3942 1922 3948 1923
rect 3774 1919 3780 1920
rect 110 1912 116 1913
rect 2006 1912 2012 1913
rect 110 1908 111 1912
rect 115 1908 116 1912
rect 110 1907 116 1908
rect 654 1911 660 1912
rect 654 1907 655 1911
rect 659 1907 660 1911
rect 654 1906 660 1907
rect 750 1911 756 1912
rect 750 1907 751 1911
rect 755 1907 756 1911
rect 750 1906 756 1907
rect 846 1911 852 1912
rect 846 1907 847 1911
rect 851 1907 852 1911
rect 846 1906 852 1907
rect 942 1911 948 1912
rect 942 1907 943 1911
rect 947 1907 948 1911
rect 942 1906 948 1907
rect 1038 1911 1044 1912
rect 1038 1907 1039 1911
rect 1043 1907 1044 1911
rect 1038 1906 1044 1907
rect 1134 1911 1140 1912
rect 1134 1907 1135 1911
rect 1139 1907 1140 1911
rect 1134 1906 1140 1907
rect 1230 1911 1236 1912
rect 1230 1907 1231 1911
rect 1235 1907 1236 1911
rect 1230 1906 1236 1907
rect 1326 1911 1332 1912
rect 1326 1907 1327 1911
rect 1331 1907 1332 1911
rect 1326 1906 1332 1907
rect 1422 1911 1428 1912
rect 1422 1907 1423 1911
rect 1427 1907 1428 1911
rect 2006 1908 2007 1912
rect 2011 1908 2012 1912
rect 2006 1907 2012 1908
rect 1422 1906 1428 1907
rect 110 1895 116 1896
rect 110 1891 111 1895
rect 115 1891 116 1895
rect 2006 1895 2012 1896
rect 110 1890 116 1891
rect 654 1892 660 1893
rect 654 1888 655 1892
rect 659 1888 660 1892
rect 654 1887 660 1888
rect 750 1892 756 1893
rect 750 1888 751 1892
rect 755 1888 756 1892
rect 750 1887 756 1888
rect 846 1892 852 1893
rect 846 1888 847 1892
rect 851 1888 852 1892
rect 846 1887 852 1888
rect 942 1892 948 1893
rect 942 1888 943 1892
rect 947 1888 948 1892
rect 942 1887 948 1888
rect 1038 1892 1044 1893
rect 1038 1888 1039 1892
rect 1043 1888 1044 1892
rect 1038 1887 1044 1888
rect 1134 1892 1140 1893
rect 1134 1888 1135 1892
rect 1139 1888 1140 1892
rect 1134 1887 1140 1888
rect 1230 1892 1236 1893
rect 1230 1888 1231 1892
rect 1235 1888 1236 1892
rect 1230 1887 1236 1888
rect 1326 1892 1332 1893
rect 1326 1888 1327 1892
rect 1331 1888 1332 1892
rect 1326 1887 1332 1888
rect 1422 1892 1428 1893
rect 1422 1888 1423 1892
rect 1427 1888 1428 1892
rect 2006 1891 2007 1895
rect 2011 1891 2012 1895
rect 2006 1890 2012 1891
rect 1422 1887 1428 1888
rect 2182 1852 2188 1853
rect 2046 1849 2052 1850
rect 2046 1845 2047 1849
rect 2051 1845 2052 1849
rect 2182 1848 2183 1852
rect 2187 1848 2188 1852
rect 2182 1847 2188 1848
rect 2278 1852 2284 1853
rect 2278 1848 2279 1852
rect 2283 1848 2284 1852
rect 2278 1847 2284 1848
rect 2382 1852 2388 1853
rect 2382 1848 2383 1852
rect 2387 1848 2388 1852
rect 2382 1847 2388 1848
rect 2486 1852 2492 1853
rect 2486 1848 2487 1852
rect 2491 1848 2492 1852
rect 2486 1847 2492 1848
rect 2590 1852 2596 1853
rect 2590 1848 2591 1852
rect 2595 1848 2596 1852
rect 2590 1847 2596 1848
rect 2702 1852 2708 1853
rect 2702 1848 2703 1852
rect 2707 1848 2708 1852
rect 2702 1847 2708 1848
rect 2830 1852 2836 1853
rect 2830 1848 2831 1852
rect 2835 1848 2836 1852
rect 2830 1847 2836 1848
rect 2990 1852 2996 1853
rect 2990 1848 2991 1852
rect 2995 1848 2996 1852
rect 2990 1847 2996 1848
rect 3182 1852 3188 1853
rect 3182 1848 3183 1852
rect 3187 1848 3188 1852
rect 3182 1847 3188 1848
rect 3398 1852 3404 1853
rect 3398 1848 3399 1852
rect 3403 1848 3404 1852
rect 3398 1847 3404 1848
rect 3630 1852 3636 1853
rect 3630 1848 3631 1852
rect 3635 1848 3636 1852
rect 3630 1847 3636 1848
rect 3838 1852 3844 1853
rect 3838 1848 3839 1852
rect 3843 1848 3844 1852
rect 3838 1847 3844 1848
rect 3942 1849 3948 1850
rect 2046 1844 2052 1845
rect 3942 1845 3943 1849
rect 3947 1845 3948 1849
rect 3942 1844 3948 1845
rect 2182 1833 2188 1834
rect 318 1832 324 1833
rect 110 1829 116 1830
rect 110 1825 111 1829
rect 115 1825 116 1829
rect 318 1828 319 1832
rect 323 1828 324 1832
rect 318 1827 324 1828
rect 446 1832 452 1833
rect 446 1828 447 1832
rect 451 1828 452 1832
rect 446 1827 452 1828
rect 582 1832 588 1833
rect 582 1828 583 1832
rect 587 1828 588 1832
rect 582 1827 588 1828
rect 718 1832 724 1833
rect 718 1828 719 1832
rect 723 1828 724 1832
rect 718 1827 724 1828
rect 854 1832 860 1833
rect 854 1828 855 1832
rect 859 1828 860 1832
rect 854 1827 860 1828
rect 990 1832 996 1833
rect 990 1828 991 1832
rect 995 1828 996 1832
rect 990 1827 996 1828
rect 1126 1832 1132 1833
rect 1126 1828 1127 1832
rect 1131 1828 1132 1832
rect 1126 1827 1132 1828
rect 1262 1832 1268 1833
rect 1262 1828 1263 1832
rect 1267 1828 1268 1832
rect 1262 1827 1268 1828
rect 1398 1832 1404 1833
rect 1398 1828 1399 1832
rect 1403 1828 1404 1832
rect 1398 1827 1404 1828
rect 1534 1832 1540 1833
rect 1534 1828 1535 1832
rect 1539 1828 1540 1832
rect 2046 1832 2052 1833
rect 1534 1827 1540 1828
rect 2006 1829 2012 1830
rect 110 1824 116 1825
rect 2006 1825 2007 1829
rect 2011 1825 2012 1829
rect 2046 1828 2047 1832
rect 2051 1828 2052 1832
rect 2182 1829 2183 1833
rect 2187 1829 2188 1833
rect 2182 1828 2188 1829
rect 2278 1833 2284 1834
rect 2278 1829 2279 1833
rect 2283 1829 2284 1833
rect 2278 1828 2284 1829
rect 2382 1833 2388 1834
rect 2382 1829 2383 1833
rect 2387 1829 2388 1833
rect 2382 1828 2388 1829
rect 2486 1833 2492 1834
rect 2486 1829 2487 1833
rect 2491 1829 2492 1833
rect 2486 1828 2492 1829
rect 2590 1833 2596 1834
rect 2590 1829 2591 1833
rect 2595 1829 2596 1833
rect 2590 1828 2596 1829
rect 2702 1833 2708 1834
rect 2702 1829 2703 1833
rect 2707 1829 2708 1833
rect 2702 1828 2708 1829
rect 2830 1833 2836 1834
rect 2830 1829 2831 1833
rect 2835 1829 2836 1833
rect 2830 1828 2836 1829
rect 2990 1833 2996 1834
rect 2990 1829 2991 1833
rect 2995 1829 2996 1833
rect 2990 1828 2996 1829
rect 3182 1833 3188 1834
rect 3182 1829 3183 1833
rect 3187 1829 3188 1833
rect 3182 1828 3188 1829
rect 3398 1833 3404 1834
rect 3398 1829 3399 1833
rect 3403 1829 3404 1833
rect 3398 1828 3404 1829
rect 3630 1833 3636 1834
rect 3630 1829 3631 1833
rect 3635 1829 3636 1833
rect 3630 1828 3636 1829
rect 3838 1833 3844 1834
rect 3838 1829 3839 1833
rect 3843 1829 3844 1833
rect 3838 1828 3844 1829
rect 3942 1832 3948 1833
rect 3942 1828 3943 1832
rect 3947 1828 3948 1832
rect 2046 1827 2052 1828
rect 3942 1827 3948 1828
rect 2006 1824 2012 1825
rect 318 1813 324 1814
rect 110 1812 116 1813
rect 110 1808 111 1812
rect 115 1808 116 1812
rect 318 1809 319 1813
rect 323 1809 324 1813
rect 318 1808 324 1809
rect 446 1813 452 1814
rect 446 1809 447 1813
rect 451 1809 452 1813
rect 446 1808 452 1809
rect 582 1813 588 1814
rect 582 1809 583 1813
rect 587 1809 588 1813
rect 582 1808 588 1809
rect 718 1813 724 1814
rect 718 1809 719 1813
rect 723 1809 724 1813
rect 718 1808 724 1809
rect 854 1813 860 1814
rect 854 1809 855 1813
rect 859 1809 860 1813
rect 854 1808 860 1809
rect 990 1813 996 1814
rect 990 1809 991 1813
rect 995 1809 996 1813
rect 990 1808 996 1809
rect 1126 1813 1132 1814
rect 1126 1809 1127 1813
rect 1131 1809 1132 1813
rect 1126 1808 1132 1809
rect 1262 1813 1268 1814
rect 1262 1809 1263 1813
rect 1267 1809 1268 1813
rect 1262 1808 1268 1809
rect 1398 1813 1404 1814
rect 1398 1809 1399 1813
rect 1403 1809 1404 1813
rect 1398 1808 1404 1809
rect 1534 1813 1540 1814
rect 1534 1809 1535 1813
rect 1539 1809 1540 1813
rect 1534 1808 1540 1809
rect 2006 1812 2012 1813
rect 2006 1808 2007 1812
rect 2011 1808 2012 1812
rect 110 1807 116 1808
rect 2006 1807 2012 1808
rect 2046 1776 2052 1777
rect 3942 1776 3948 1777
rect 2046 1772 2047 1776
rect 2051 1772 2052 1776
rect 2046 1771 2052 1772
rect 2126 1775 2132 1776
rect 2126 1771 2127 1775
rect 2131 1771 2132 1775
rect 2126 1770 2132 1771
rect 2310 1775 2316 1776
rect 2310 1771 2311 1775
rect 2315 1771 2316 1775
rect 2310 1770 2316 1771
rect 2494 1775 2500 1776
rect 2494 1771 2495 1775
rect 2499 1771 2500 1775
rect 2494 1770 2500 1771
rect 2686 1775 2692 1776
rect 2686 1771 2687 1775
rect 2691 1771 2692 1775
rect 2686 1770 2692 1771
rect 2878 1775 2884 1776
rect 2878 1771 2879 1775
rect 2883 1771 2884 1775
rect 2878 1770 2884 1771
rect 3070 1775 3076 1776
rect 3070 1771 3071 1775
rect 3075 1771 3076 1775
rect 3070 1770 3076 1771
rect 3262 1775 3268 1776
rect 3262 1771 3263 1775
rect 3267 1771 3268 1775
rect 3262 1770 3268 1771
rect 3462 1775 3468 1776
rect 3462 1771 3463 1775
rect 3467 1771 3468 1775
rect 3462 1770 3468 1771
rect 3662 1775 3668 1776
rect 3662 1771 3663 1775
rect 3667 1771 3668 1775
rect 3662 1770 3668 1771
rect 3838 1775 3844 1776
rect 3838 1771 3839 1775
rect 3843 1771 3844 1775
rect 3942 1772 3943 1776
rect 3947 1772 3948 1776
rect 3942 1771 3948 1772
rect 3838 1770 3844 1771
rect 2046 1759 2052 1760
rect 110 1756 116 1757
rect 2006 1756 2012 1757
rect 110 1752 111 1756
rect 115 1752 116 1756
rect 110 1751 116 1752
rect 254 1755 260 1756
rect 254 1751 255 1755
rect 259 1751 260 1755
rect 254 1750 260 1751
rect 390 1755 396 1756
rect 390 1751 391 1755
rect 395 1751 396 1755
rect 390 1750 396 1751
rect 534 1755 540 1756
rect 534 1751 535 1755
rect 539 1751 540 1755
rect 534 1750 540 1751
rect 694 1755 700 1756
rect 694 1751 695 1755
rect 699 1751 700 1755
rect 694 1750 700 1751
rect 862 1755 868 1756
rect 862 1751 863 1755
rect 867 1751 868 1755
rect 862 1750 868 1751
rect 1030 1755 1036 1756
rect 1030 1751 1031 1755
rect 1035 1751 1036 1755
rect 1030 1750 1036 1751
rect 1206 1755 1212 1756
rect 1206 1751 1207 1755
rect 1211 1751 1212 1755
rect 1206 1750 1212 1751
rect 1382 1755 1388 1756
rect 1382 1751 1383 1755
rect 1387 1751 1388 1755
rect 1382 1750 1388 1751
rect 1558 1755 1564 1756
rect 1558 1751 1559 1755
rect 1563 1751 1564 1755
rect 1558 1750 1564 1751
rect 1742 1755 1748 1756
rect 1742 1751 1743 1755
rect 1747 1751 1748 1755
rect 2006 1752 2007 1756
rect 2011 1752 2012 1756
rect 2046 1755 2047 1759
rect 2051 1755 2052 1759
rect 3942 1759 3948 1760
rect 2046 1754 2052 1755
rect 2126 1756 2132 1757
rect 2006 1751 2012 1752
rect 2126 1752 2127 1756
rect 2131 1752 2132 1756
rect 2126 1751 2132 1752
rect 2310 1756 2316 1757
rect 2310 1752 2311 1756
rect 2315 1752 2316 1756
rect 2310 1751 2316 1752
rect 2494 1756 2500 1757
rect 2494 1752 2495 1756
rect 2499 1752 2500 1756
rect 2494 1751 2500 1752
rect 2686 1756 2692 1757
rect 2686 1752 2687 1756
rect 2691 1752 2692 1756
rect 2686 1751 2692 1752
rect 2878 1756 2884 1757
rect 2878 1752 2879 1756
rect 2883 1752 2884 1756
rect 2878 1751 2884 1752
rect 3070 1756 3076 1757
rect 3070 1752 3071 1756
rect 3075 1752 3076 1756
rect 3070 1751 3076 1752
rect 3262 1756 3268 1757
rect 3262 1752 3263 1756
rect 3267 1752 3268 1756
rect 3262 1751 3268 1752
rect 3462 1756 3468 1757
rect 3462 1752 3463 1756
rect 3467 1752 3468 1756
rect 3462 1751 3468 1752
rect 3662 1756 3668 1757
rect 3662 1752 3663 1756
rect 3667 1752 3668 1756
rect 3662 1751 3668 1752
rect 3838 1756 3844 1757
rect 3838 1752 3839 1756
rect 3843 1752 3844 1756
rect 3942 1755 3943 1759
rect 3947 1755 3948 1759
rect 3942 1754 3948 1755
rect 3838 1751 3844 1752
rect 1742 1750 1748 1751
rect 110 1739 116 1740
rect 110 1735 111 1739
rect 115 1735 116 1739
rect 2006 1739 2012 1740
rect 110 1734 116 1735
rect 254 1736 260 1737
rect 254 1732 255 1736
rect 259 1732 260 1736
rect 254 1731 260 1732
rect 390 1736 396 1737
rect 390 1732 391 1736
rect 395 1732 396 1736
rect 390 1731 396 1732
rect 534 1736 540 1737
rect 534 1732 535 1736
rect 539 1732 540 1736
rect 534 1731 540 1732
rect 694 1736 700 1737
rect 694 1732 695 1736
rect 699 1732 700 1736
rect 694 1731 700 1732
rect 862 1736 868 1737
rect 862 1732 863 1736
rect 867 1732 868 1736
rect 862 1731 868 1732
rect 1030 1736 1036 1737
rect 1030 1732 1031 1736
rect 1035 1732 1036 1736
rect 1030 1731 1036 1732
rect 1206 1736 1212 1737
rect 1206 1732 1207 1736
rect 1211 1732 1212 1736
rect 1206 1731 1212 1732
rect 1382 1736 1388 1737
rect 1382 1732 1383 1736
rect 1387 1732 1388 1736
rect 1382 1731 1388 1732
rect 1558 1736 1564 1737
rect 1558 1732 1559 1736
rect 1563 1732 1564 1736
rect 1558 1731 1564 1732
rect 1742 1736 1748 1737
rect 1742 1732 1743 1736
rect 1747 1732 1748 1736
rect 2006 1735 2007 1739
rect 2011 1735 2012 1739
rect 2006 1734 2012 1735
rect 1742 1731 1748 1732
rect 2070 1692 2076 1693
rect 2046 1689 2052 1690
rect 2046 1685 2047 1689
rect 2051 1685 2052 1689
rect 2070 1688 2071 1692
rect 2075 1688 2076 1692
rect 2070 1687 2076 1688
rect 2190 1692 2196 1693
rect 2190 1688 2191 1692
rect 2195 1688 2196 1692
rect 2190 1687 2196 1688
rect 2342 1692 2348 1693
rect 2342 1688 2343 1692
rect 2347 1688 2348 1692
rect 2342 1687 2348 1688
rect 2510 1692 2516 1693
rect 2510 1688 2511 1692
rect 2515 1688 2516 1692
rect 2510 1687 2516 1688
rect 2686 1692 2692 1693
rect 2686 1688 2687 1692
rect 2691 1688 2692 1692
rect 2686 1687 2692 1688
rect 2870 1692 2876 1693
rect 2870 1688 2871 1692
rect 2875 1688 2876 1692
rect 2870 1687 2876 1688
rect 3062 1692 3068 1693
rect 3062 1688 3063 1692
rect 3067 1688 3068 1692
rect 3062 1687 3068 1688
rect 3254 1692 3260 1693
rect 3254 1688 3255 1692
rect 3259 1688 3260 1692
rect 3254 1687 3260 1688
rect 3446 1692 3452 1693
rect 3446 1688 3447 1692
rect 3451 1688 3452 1692
rect 3446 1687 3452 1688
rect 3646 1692 3652 1693
rect 3646 1688 3647 1692
rect 3651 1688 3652 1692
rect 3646 1687 3652 1688
rect 3838 1692 3844 1693
rect 3838 1688 3839 1692
rect 3843 1688 3844 1692
rect 3838 1687 3844 1688
rect 3942 1689 3948 1690
rect 2046 1684 2052 1685
rect 3942 1685 3943 1689
rect 3947 1685 3948 1689
rect 3942 1684 3948 1685
rect 134 1676 140 1677
rect 110 1673 116 1674
rect 110 1669 111 1673
rect 115 1669 116 1673
rect 134 1672 135 1676
rect 139 1672 140 1676
rect 134 1671 140 1672
rect 262 1676 268 1677
rect 262 1672 263 1676
rect 267 1672 268 1676
rect 262 1671 268 1672
rect 430 1676 436 1677
rect 430 1672 431 1676
rect 435 1672 436 1676
rect 430 1671 436 1672
rect 606 1676 612 1677
rect 606 1672 607 1676
rect 611 1672 612 1676
rect 606 1671 612 1672
rect 798 1676 804 1677
rect 798 1672 799 1676
rect 803 1672 804 1676
rect 798 1671 804 1672
rect 998 1676 1004 1677
rect 998 1672 999 1676
rect 1003 1672 1004 1676
rect 998 1671 1004 1672
rect 1198 1676 1204 1677
rect 1198 1672 1199 1676
rect 1203 1672 1204 1676
rect 1198 1671 1204 1672
rect 1406 1676 1412 1677
rect 1406 1672 1407 1676
rect 1411 1672 1412 1676
rect 1406 1671 1412 1672
rect 1622 1676 1628 1677
rect 1622 1672 1623 1676
rect 1627 1672 1628 1676
rect 1622 1671 1628 1672
rect 1838 1676 1844 1677
rect 1838 1672 1839 1676
rect 1843 1672 1844 1676
rect 1838 1671 1844 1672
rect 2006 1673 2012 1674
rect 2070 1673 2076 1674
rect 110 1668 116 1669
rect 2006 1669 2007 1673
rect 2011 1669 2012 1673
rect 2006 1668 2012 1669
rect 2046 1672 2052 1673
rect 2046 1668 2047 1672
rect 2051 1668 2052 1672
rect 2070 1669 2071 1673
rect 2075 1669 2076 1673
rect 2070 1668 2076 1669
rect 2190 1673 2196 1674
rect 2190 1669 2191 1673
rect 2195 1669 2196 1673
rect 2190 1668 2196 1669
rect 2342 1673 2348 1674
rect 2342 1669 2343 1673
rect 2347 1669 2348 1673
rect 2342 1668 2348 1669
rect 2510 1673 2516 1674
rect 2510 1669 2511 1673
rect 2515 1669 2516 1673
rect 2510 1668 2516 1669
rect 2686 1673 2692 1674
rect 2686 1669 2687 1673
rect 2691 1669 2692 1673
rect 2686 1668 2692 1669
rect 2870 1673 2876 1674
rect 2870 1669 2871 1673
rect 2875 1669 2876 1673
rect 2870 1668 2876 1669
rect 3062 1673 3068 1674
rect 3062 1669 3063 1673
rect 3067 1669 3068 1673
rect 3062 1668 3068 1669
rect 3254 1673 3260 1674
rect 3254 1669 3255 1673
rect 3259 1669 3260 1673
rect 3254 1668 3260 1669
rect 3446 1673 3452 1674
rect 3446 1669 3447 1673
rect 3451 1669 3452 1673
rect 3446 1668 3452 1669
rect 3646 1673 3652 1674
rect 3646 1669 3647 1673
rect 3651 1669 3652 1673
rect 3646 1668 3652 1669
rect 3838 1673 3844 1674
rect 3838 1669 3839 1673
rect 3843 1669 3844 1673
rect 3838 1668 3844 1669
rect 3942 1672 3948 1673
rect 3942 1668 3943 1672
rect 3947 1668 3948 1672
rect 2046 1667 2052 1668
rect 3942 1667 3948 1668
rect 134 1657 140 1658
rect 110 1656 116 1657
rect 110 1652 111 1656
rect 115 1652 116 1656
rect 134 1653 135 1657
rect 139 1653 140 1657
rect 134 1652 140 1653
rect 262 1657 268 1658
rect 262 1653 263 1657
rect 267 1653 268 1657
rect 262 1652 268 1653
rect 430 1657 436 1658
rect 430 1653 431 1657
rect 435 1653 436 1657
rect 430 1652 436 1653
rect 606 1657 612 1658
rect 606 1653 607 1657
rect 611 1653 612 1657
rect 606 1652 612 1653
rect 798 1657 804 1658
rect 798 1653 799 1657
rect 803 1653 804 1657
rect 798 1652 804 1653
rect 998 1657 1004 1658
rect 998 1653 999 1657
rect 1003 1653 1004 1657
rect 998 1652 1004 1653
rect 1198 1657 1204 1658
rect 1198 1653 1199 1657
rect 1203 1653 1204 1657
rect 1198 1652 1204 1653
rect 1406 1657 1412 1658
rect 1406 1653 1407 1657
rect 1411 1653 1412 1657
rect 1406 1652 1412 1653
rect 1622 1657 1628 1658
rect 1622 1653 1623 1657
rect 1627 1653 1628 1657
rect 1622 1652 1628 1653
rect 1838 1657 1844 1658
rect 1838 1653 1839 1657
rect 1843 1653 1844 1657
rect 1838 1652 1844 1653
rect 2006 1656 2012 1657
rect 2006 1652 2007 1656
rect 2011 1652 2012 1656
rect 110 1651 116 1652
rect 2006 1651 2012 1652
rect 2046 1620 2052 1621
rect 3942 1620 3948 1621
rect 2046 1616 2047 1620
rect 2051 1616 2052 1620
rect 2046 1615 2052 1616
rect 2070 1619 2076 1620
rect 2070 1615 2071 1619
rect 2075 1615 2076 1619
rect 2070 1614 2076 1615
rect 2334 1619 2340 1620
rect 2334 1615 2335 1619
rect 2339 1615 2340 1619
rect 2334 1614 2340 1615
rect 2598 1619 2604 1620
rect 2598 1615 2599 1619
rect 2603 1615 2604 1619
rect 2598 1614 2604 1615
rect 2838 1619 2844 1620
rect 2838 1615 2839 1619
rect 2843 1615 2844 1619
rect 2838 1614 2844 1615
rect 3046 1619 3052 1620
rect 3046 1615 3047 1619
rect 3051 1615 3052 1619
rect 3046 1614 3052 1615
rect 3230 1619 3236 1620
rect 3230 1615 3231 1619
rect 3235 1615 3236 1619
rect 3230 1614 3236 1615
rect 3398 1619 3404 1620
rect 3398 1615 3399 1619
rect 3403 1615 3404 1619
rect 3398 1614 3404 1615
rect 3550 1619 3556 1620
rect 3550 1615 3551 1619
rect 3555 1615 3556 1619
rect 3550 1614 3556 1615
rect 3694 1619 3700 1620
rect 3694 1615 3695 1619
rect 3699 1615 3700 1619
rect 3694 1614 3700 1615
rect 3838 1619 3844 1620
rect 3838 1615 3839 1619
rect 3843 1615 3844 1619
rect 3942 1616 3943 1620
rect 3947 1616 3948 1620
rect 3942 1615 3948 1616
rect 3838 1614 3844 1615
rect 110 1604 116 1605
rect 2006 1604 2012 1605
rect 110 1600 111 1604
rect 115 1600 116 1604
rect 110 1599 116 1600
rect 134 1603 140 1604
rect 134 1599 135 1603
rect 139 1599 140 1603
rect 134 1598 140 1599
rect 286 1603 292 1604
rect 286 1599 287 1603
rect 291 1599 292 1603
rect 286 1598 292 1599
rect 470 1603 476 1604
rect 470 1599 471 1603
rect 475 1599 476 1603
rect 470 1598 476 1599
rect 654 1603 660 1604
rect 654 1599 655 1603
rect 659 1599 660 1603
rect 654 1598 660 1599
rect 838 1603 844 1604
rect 838 1599 839 1603
rect 843 1599 844 1603
rect 838 1598 844 1599
rect 1014 1603 1020 1604
rect 1014 1599 1015 1603
rect 1019 1599 1020 1603
rect 1014 1598 1020 1599
rect 1182 1603 1188 1604
rect 1182 1599 1183 1603
rect 1187 1599 1188 1603
rect 1182 1598 1188 1599
rect 1342 1603 1348 1604
rect 1342 1599 1343 1603
rect 1347 1599 1348 1603
rect 1342 1598 1348 1599
rect 1494 1603 1500 1604
rect 1494 1599 1495 1603
rect 1499 1599 1500 1603
rect 1494 1598 1500 1599
rect 1638 1603 1644 1604
rect 1638 1599 1639 1603
rect 1643 1599 1644 1603
rect 1638 1598 1644 1599
rect 1782 1603 1788 1604
rect 1782 1599 1783 1603
rect 1787 1599 1788 1603
rect 1782 1598 1788 1599
rect 1902 1603 1908 1604
rect 1902 1599 1903 1603
rect 1907 1599 1908 1603
rect 2006 1600 2007 1604
rect 2011 1600 2012 1604
rect 2006 1599 2012 1600
rect 2046 1603 2052 1604
rect 2046 1599 2047 1603
rect 2051 1599 2052 1603
rect 3942 1603 3948 1604
rect 1902 1598 1908 1599
rect 2046 1598 2052 1599
rect 2070 1600 2076 1601
rect 2070 1596 2071 1600
rect 2075 1596 2076 1600
rect 2070 1595 2076 1596
rect 2334 1600 2340 1601
rect 2334 1596 2335 1600
rect 2339 1596 2340 1600
rect 2334 1595 2340 1596
rect 2598 1600 2604 1601
rect 2598 1596 2599 1600
rect 2603 1596 2604 1600
rect 2598 1595 2604 1596
rect 2838 1600 2844 1601
rect 2838 1596 2839 1600
rect 2843 1596 2844 1600
rect 2838 1595 2844 1596
rect 3046 1600 3052 1601
rect 3046 1596 3047 1600
rect 3051 1596 3052 1600
rect 3046 1595 3052 1596
rect 3230 1600 3236 1601
rect 3230 1596 3231 1600
rect 3235 1596 3236 1600
rect 3230 1595 3236 1596
rect 3398 1600 3404 1601
rect 3398 1596 3399 1600
rect 3403 1596 3404 1600
rect 3398 1595 3404 1596
rect 3550 1600 3556 1601
rect 3550 1596 3551 1600
rect 3555 1596 3556 1600
rect 3550 1595 3556 1596
rect 3694 1600 3700 1601
rect 3694 1596 3695 1600
rect 3699 1596 3700 1600
rect 3694 1595 3700 1596
rect 3838 1600 3844 1601
rect 3838 1596 3839 1600
rect 3843 1596 3844 1600
rect 3942 1599 3943 1603
rect 3947 1599 3948 1603
rect 3942 1598 3948 1599
rect 3838 1595 3844 1596
rect 110 1587 116 1588
rect 110 1583 111 1587
rect 115 1583 116 1587
rect 2006 1587 2012 1588
rect 110 1582 116 1583
rect 134 1584 140 1585
rect 134 1580 135 1584
rect 139 1580 140 1584
rect 134 1579 140 1580
rect 286 1584 292 1585
rect 286 1580 287 1584
rect 291 1580 292 1584
rect 286 1579 292 1580
rect 470 1584 476 1585
rect 470 1580 471 1584
rect 475 1580 476 1584
rect 470 1579 476 1580
rect 654 1584 660 1585
rect 654 1580 655 1584
rect 659 1580 660 1584
rect 654 1579 660 1580
rect 838 1584 844 1585
rect 838 1580 839 1584
rect 843 1580 844 1584
rect 838 1579 844 1580
rect 1014 1584 1020 1585
rect 1014 1580 1015 1584
rect 1019 1580 1020 1584
rect 1014 1579 1020 1580
rect 1182 1584 1188 1585
rect 1182 1580 1183 1584
rect 1187 1580 1188 1584
rect 1182 1579 1188 1580
rect 1342 1584 1348 1585
rect 1342 1580 1343 1584
rect 1347 1580 1348 1584
rect 1342 1579 1348 1580
rect 1494 1584 1500 1585
rect 1494 1580 1495 1584
rect 1499 1580 1500 1584
rect 1494 1579 1500 1580
rect 1638 1584 1644 1585
rect 1638 1580 1639 1584
rect 1643 1580 1644 1584
rect 1638 1579 1644 1580
rect 1782 1584 1788 1585
rect 1782 1580 1783 1584
rect 1787 1580 1788 1584
rect 1782 1579 1788 1580
rect 1902 1584 1908 1585
rect 1902 1580 1903 1584
rect 1907 1580 1908 1584
rect 2006 1583 2007 1587
rect 2011 1583 2012 1587
rect 2006 1582 2012 1583
rect 1902 1579 1908 1580
rect 2582 1536 2588 1537
rect 2046 1533 2052 1534
rect 2046 1529 2047 1533
rect 2051 1529 2052 1533
rect 2582 1532 2583 1536
rect 2587 1532 2588 1536
rect 2582 1531 2588 1532
rect 2742 1536 2748 1537
rect 2742 1532 2743 1536
rect 2747 1532 2748 1536
rect 2742 1531 2748 1532
rect 2902 1536 2908 1537
rect 2902 1532 2903 1536
rect 2907 1532 2908 1536
rect 2902 1531 2908 1532
rect 3062 1536 3068 1537
rect 3062 1532 3063 1536
rect 3067 1532 3068 1536
rect 3062 1531 3068 1532
rect 3222 1536 3228 1537
rect 3222 1532 3223 1536
rect 3227 1532 3228 1536
rect 3222 1531 3228 1532
rect 3382 1536 3388 1537
rect 3382 1532 3383 1536
rect 3387 1532 3388 1536
rect 3382 1531 3388 1532
rect 3542 1536 3548 1537
rect 3542 1532 3543 1536
rect 3547 1532 3548 1536
rect 3542 1531 3548 1532
rect 3702 1536 3708 1537
rect 3702 1532 3703 1536
rect 3707 1532 3708 1536
rect 3702 1531 3708 1532
rect 3942 1533 3948 1534
rect 2046 1528 2052 1529
rect 3942 1529 3943 1533
rect 3947 1529 3948 1533
rect 3942 1528 3948 1529
rect 134 1520 140 1521
rect 110 1517 116 1518
rect 110 1513 111 1517
rect 115 1513 116 1517
rect 134 1516 135 1520
rect 139 1516 140 1520
rect 134 1515 140 1516
rect 294 1520 300 1521
rect 294 1516 295 1520
rect 299 1516 300 1520
rect 294 1515 300 1516
rect 486 1520 492 1521
rect 486 1516 487 1520
rect 491 1516 492 1520
rect 486 1515 492 1516
rect 686 1520 692 1521
rect 686 1516 687 1520
rect 691 1516 692 1520
rect 686 1515 692 1516
rect 886 1520 892 1521
rect 886 1516 887 1520
rect 891 1516 892 1520
rect 886 1515 892 1516
rect 1078 1520 1084 1521
rect 1078 1516 1079 1520
rect 1083 1516 1084 1520
rect 1078 1515 1084 1516
rect 1262 1520 1268 1521
rect 1262 1516 1263 1520
rect 1267 1516 1268 1520
rect 1262 1515 1268 1516
rect 1446 1520 1452 1521
rect 1446 1516 1447 1520
rect 1451 1516 1452 1520
rect 1446 1515 1452 1516
rect 1622 1520 1628 1521
rect 1622 1516 1623 1520
rect 1627 1516 1628 1520
rect 1622 1515 1628 1516
rect 1806 1520 1812 1521
rect 1806 1516 1807 1520
rect 1811 1516 1812 1520
rect 1806 1515 1812 1516
rect 2006 1517 2012 1518
rect 2582 1517 2588 1518
rect 110 1512 116 1513
rect 2006 1513 2007 1517
rect 2011 1513 2012 1517
rect 2006 1512 2012 1513
rect 2046 1516 2052 1517
rect 2046 1512 2047 1516
rect 2051 1512 2052 1516
rect 2582 1513 2583 1517
rect 2587 1513 2588 1517
rect 2582 1512 2588 1513
rect 2742 1517 2748 1518
rect 2742 1513 2743 1517
rect 2747 1513 2748 1517
rect 2742 1512 2748 1513
rect 2902 1517 2908 1518
rect 2902 1513 2903 1517
rect 2907 1513 2908 1517
rect 2902 1512 2908 1513
rect 3062 1517 3068 1518
rect 3062 1513 3063 1517
rect 3067 1513 3068 1517
rect 3062 1512 3068 1513
rect 3222 1517 3228 1518
rect 3222 1513 3223 1517
rect 3227 1513 3228 1517
rect 3222 1512 3228 1513
rect 3382 1517 3388 1518
rect 3382 1513 3383 1517
rect 3387 1513 3388 1517
rect 3382 1512 3388 1513
rect 3542 1517 3548 1518
rect 3542 1513 3543 1517
rect 3547 1513 3548 1517
rect 3542 1512 3548 1513
rect 3702 1517 3708 1518
rect 3702 1513 3703 1517
rect 3707 1513 3708 1517
rect 3702 1512 3708 1513
rect 3942 1516 3948 1517
rect 3942 1512 3943 1516
rect 3947 1512 3948 1516
rect 2046 1511 2052 1512
rect 3942 1511 3948 1512
rect 134 1501 140 1502
rect 110 1500 116 1501
rect 110 1496 111 1500
rect 115 1496 116 1500
rect 134 1497 135 1501
rect 139 1497 140 1501
rect 134 1496 140 1497
rect 294 1501 300 1502
rect 294 1497 295 1501
rect 299 1497 300 1501
rect 294 1496 300 1497
rect 486 1501 492 1502
rect 486 1497 487 1501
rect 491 1497 492 1501
rect 486 1496 492 1497
rect 686 1501 692 1502
rect 686 1497 687 1501
rect 691 1497 692 1501
rect 686 1496 692 1497
rect 886 1501 892 1502
rect 886 1497 887 1501
rect 891 1497 892 1501
rect 886 1496 892 1497
rect 1078 1501 1084 1502
rect 1078 1497 1079 1501
rect 1083 1497 1084 1501
rect 1078 1496 1084 1497
rect 1262 1501 1268 1502
rect 1262 1497 1263 1501
rect 1267 1497 1268 1501
rect 1262 1496 1268 1497
rect 1446 1501 1452 1502
rect 1446 1497 1447 1501
rect 1451 1497 1452 1501
rect 1446 1496 1452 1497
rect 1622 1501 1628 1502
rect 1622 1497 1623 1501
rect 1627 1497 1628 1501
rect 1622 1496 1628 1497
rect 1806 1501 1812 1502
rect 1806 1497 1807 1501
rect 1811 1497 1812 1501
rect 1806 1496 1812 1497
rect 2006 1500 2012 1501
rect 2006 1496 2007 1500
rect 2011 1496 2012 1500
rect 110 1495 116 1496
rect 2006 1495 2012 1496
rect 2046 1464 2052 1465
rect 3942 1464 3948 1465
rect 2046 1460 2047 1464
rect 2051 1460 2052 1464
rect 2046 1459 2052 1460
rect 2414 1463 2420 1464
rect 2414 1459 2415 1463
rect 2419 1459 2420 1463
rect 2414 1458 2420 1459
rect 2510 1463 2516 1464
rect 2510 1459 2511 1463
rect 2515 1459 2516 1463
rect 2510 1458 2516 1459
rect 2606 1463 2612 1464
rect 2606 1459 2607 1463
rect 2611 1459 2612 1463
rect 2606 1458 2612 1459
rect 2702 1463 2708 1464
rect 2702 1459 2703 1463
rect 2707 1459 2708 1463
rect 2702 1458 2708 1459
rect 2798 1463 2804 1464
rect 2798 1459 2799 1463
rect 2803 1459 2804 1463
rect 2798 1458 2804 1459
rect 2918 1463 2924 1464
rect 2918 1459 2919 1463
rect 2923 1459 2924 1463
rect 2918 1458 2924 1459
rect 3062 1463 3068 1464
rect 3062 1459 3063 1463
rect 3067 1459 3068 1463
rect 3062 1458 3068 1459
rect 3230 1463 3236 1464
rect 3230 1459 3231 1463
rect 3235 1459 3236 1463
rect 3230 1458 3236 1459
rect 3414 1463 3420 1464
rect 3414 1459 3415 1463
rect 3419 1459 3420 1463
rect 3414 1458 3420 1459
rect 3614 1463 3620 1464
rect 3614 1459 3615 1463
rect 3619 1459 3620 1463
rect 3614 1458 3620 1459
rect 3814 1463 3820 1464
rect 3814 1459 3815 1463
rect 3819 1459 3820 1463
rect 3942 1460 3943 1464
rect 3947 1460 3948 1464
rect 3942 1459 3948 1460
rect 3814 1458 3820 1459
rect 110 1448 116 1449
rect 2006 1448 2012 1449
rect 110 1444 111 1448
rect 115 1444 116 1448
rect 110 1443 116 1444
rect 174 1447 180 1448
rect 174 1443 175 1447
rect 179 1443 180 1447
rect 174 1442 180 1443
rect 358 1447 364 1448
rect 358 1443 359 1447
rect 363 1443 364 1447
rect 358 1442 364 1443
rect 566 1447 572 1448
rect 566 1443 567 1447
rect 571 1443 572 1447
rect 566 1442 572 1443
rect 782 1447 788 1448
rect 782 1443 783 1447
rect 787 1443 788 1447
rect 782 1442 788 1443
rect 1006 1447 1012 1448
rect 1006 1443 1007 1447
rect 1011 1443 1012 1447
rect 1006 1442 1012 1443
rect 1230 1447 1236 1448
rect 1230 1443 1231 1447
rect 1235 1443 1236 1447
rect 1230 1442 1236 1443
rect 1462 1447 1468 1448
rect 1462 1443 1463 1447
rect 1467 1443 1468 1447
rect 1462 1442 1468 1443
rect 1694 1447 1700 1448
rect 1694 1443 1695 1447
rect 1699 1443 1700 1447
rect 1694 1442 1700 1443
rect 1902 1447 1908 1448
rect 1902 1443 1903 1447
rect 1907 1443 1908 1447
rect 2006 1444 2007 1448
rect 2011 1444 2012 1448
rect 2006 1443 2012 1444
rect 2046 1447 2052 1448
rect 2046 1443 2047 1447
rect 2051 1443 2052 1447
rect 3942 1447 3948 1448
rect 1902 1442 1908 1443
rect 2046 1442 2052 1443
rect 2414 1444 2420 1445
rect 2414 1440 2415 1444
rect 2419 1440 2420 1444
rect 2414 1439 2420 1440
rect 2510 1444 2516 1445
rect 2510 1440 2511 1444
rect 2515 1440 2516 1444
rect 2510 1439 2516 1440
rect 2606 1444 2612 1445
rect 2606 1440 2607 1444
rect 2611 1440 2612 1444
rect 2606 1439 2612 1440
rect 2702 1444 2708 1445
rect 2702 1440 2703 1444
rect 2707 1440 2708 1444
rect 2702 1439 2708 1440
rect 2798 1444 2804 1445
rect 2798 1440 2799 1444
rect 2803 1440 2804 1444
rect 2798 1439 2804 1440
rect 2918 1444 2924 1445
rect 2918 1440 2919 1444
rect 2923 1440 2924 1444
rect 2918 1439 2924 1440
rect 3062 1444 3068 1445
rect 3062 1440 3063 1444
rect 3067 1440 3068 1444
rect 3062 1439 3068 1440
rect 3230 1444 3236 1445
rect 3230 1440 3231 1444
rect 3235 1440 3236 1444
rect 3230 1439 3236 1440
rect 3414 1444 3420 1445
rect 3414 1440 3415 1444
rect 3419 1440 3420 1444
rect 3414 1439 3420 1440
rect 3614 1444 3620 1445
rect 3614 1440 3615 1444
rect 3619 1440 3620 1444
rect 3614 1439 3620 1440
rect 3814 1444 3820 1445
rect 3814 1440 3815 1444
rect 3819 1440 3820 1444
rect 3942 1443 3943 1447
rect 3947 1443 3948 1447
rect 3942 1442 3948 1443
rect 3814 1439 3820 1440
rect 110 1431 116 1432
rect 110 1427 111 1431
rect 115 1427 116 1431
rect 2006 1431 2012 1432
rect 110 1426 116 1427
rect 174 1428 180 1429
rect 174 1424 175 1428
rect 179 1424 180 1428
rect 174 1423 180 1424
rect 358 1428 364 1429
rect 358 1424 359 1428
rect 363 1424 364 1428
rect 358 1423 364 1424
rect 566 1428 572 1429
rect 566 1424 567 1428
rect 571 1424 572 1428
rect 566 1423 572 1424
rect 782 1428 788 1429
rect 782 1424 783 1428
rect 787 1424 788 1428
rect 782 1423 788 1424
rect 1006 1428 1012 1429
rect 1006 1424 1007 1428
rect 1011 1424 1012 1428
rect 1006 1423 1012 1424
rect 1230 1428 1236 1429
rect 1230 1424 1231 1428
rect 1235 1424 1236 1428
rect 1230 1423 1236 1424
rect 1462 1428 1468 1429
rect 1462 1424 1463 1428
rect 1467 1424 1468 1428
rect 1462 1423 1468 1424
rect 1694 1428 1700 1429
rect 1694 1424 1695 1428
rect 1699 1424 1700 1428
rect 1694 1423 1700 1424
rect 1902 1428 1908 1429
rect 1902 1424 1903 1428
rect 1907 1424 1908 1428
rect 2006 1427 2007 1431
rect 2011 1427 2012 1431
rect 2006 1426 2012 1427
rect 1902 1423 1908 1424
rect 326 1368 332 1369
rect 110 1365 116 1366
rect 110 1361 111 1365
rect 115 1361 116 1365
rect 326 1364 327 1368
rect 331 1364 332 1368
rect 326 1363 332 1364
rect 462 1368 468 1369
rect 462 1364 463 1368
rect 467 1364 468 1368
rect 462 1363 468 1364
rect 598 1368 604 1369
rect 598 1364 599 1368
rect 603 1364 604 1368
rect 598 1363 604 1364
rect 726 1368 732 1369
rect 726 1364 727 1368
rect 731 1364 732 1368
rect 726 1363 732 1364
rect 854 1368 860 1369
rect 854 1364 855 1368
rect 859 1364 860 1368
rect 854 1363 860 1364
rect 982 1368 988 1369
rect 982 1364 983 1368
rect 987 1364 988 1368
rect 982 1363 988 1364
rect 1118 1368 1124 1369
rect 1118 1364 1119 1368
rect 1123 1364 1124 1368
rect 1118 1363 1124 1364
rect 1262 1368 1268 1369
rect 1262 1364 1263 1368
rect 1267 1364 1268 1368
rect 1262 1363 1268 1364
rect 1422 1368 1428 1369
rect 1422 1364 1423 1368
rect 1427 1364 1428 1368
rect 1422 1363 1428 1364
rect 1582 1368 1588 1369
rect 1582 1364 1583 1368
rect 1587 1364 1588 1368
rect 1582 1363 1588 1364
rect 1750 1368 1756 1369
rect 1750 1364 1751 1368
rect 1755 1364 1756 1368
rect 1750 1363 1756 1364
rect 1902 1368 1908 1369
rect 1902 1364 1903 1368
rect 1907 1364 1908 1368
rect 1902 1363 1908 1364
rect 2006 1365 2012 1366
rect 110 1360 116 1361
rect 2006 1361 2007 1365
rect 2011 1361 2012 1365
rect 2070 1364 2076 1365
rect 2006 1360 2012 1361
rect 2046 1361 2052 1362
rect 2046 1357 2047 1361
rect 2051 1357 2052 1361
rect 2070 1360 2071 1364
rect 2075 1360 2076 1364
rect 2070 1359 2076 1360
rect 2302 1364 2308 1365
rect 2302 1360 2303 1364
rect 2307 1360 2308 1364
rect 2302 1359 2308 1360
rect 2558 1364 2564 1365
rect 2558 1360 2559 1364
rect 2563 1360 2564 1364
rect 2558 1359 2564 1360
rect 2806 1364 2812 1365
rect 2806 1360 2807 1364
rect 2811 1360 2812 1364
rect 2806 1359 2812 1360
rect 3054 1364 3060 1365
rect 3054 1360 3055 1364
rect 3059 1360 3060 1364
rect 3054 1359 3060 1360
rect 3302 1364 3308 1365
rect 3302 1360 3303 1364
rect 3307 1360 3308 1364
rect 3302 1359 3308 1360
rect 3558 1364 3564 1365
rect 3558 1360 3559 1364
rect 3563 1360 3564 1364
rect 3558 1359 3564 1360
rect 3814 1364 3820 1365
rect 3814 1360 3815 1364
rect 3819 1360 3820 1364
rect 3814 1359 3820 1360
rect 3942 1361 3948 1362
rect 2046 1356 2052 1357
rect 3942 1357 3943 1361
rect 3947 1357 3948 1361
rect 3942 1356 3948 1357
rect 326 1349 332 1350
rect 110 1348 116 1349
rect 110 1344 111 1348
rect 115 1344 116 1348
rect 326 1345 327 1349
rect 331 1345 332 1349
rect 326 1344 332 1345
rect 462 1349 468 1350
rect 462 1345 463 1349
rect 467 1345 468 1349
rect 462 1344 468 1345
rect 598 1349 604 1350
rect 598 1345 599 1349
rect 603 1345 604 1349
rect 598 1344 604 1345
rect 726 1349 732 1350
rect 726 1345 727 1349
rect 731 1345 732 1349
rect 726 1344 732 1345
rect 854 1349 860 1350
rect 854 1345 855 1349
rect 859 1345 860 1349
rect 854 1344 860 1345
rect 982 1349 988 1350
rect 982 1345 983 1349
rect 987 1345 988 1349
rect 982 1344 988 1345
rect 1118 1349 1124 1350
rect 1118 1345 1119 1349
rect 1123 1345 1124 1349
rect 1118 1344 1124 1345
rect 1262 1349 1268 1350
rect 1262 1345 1263 1349
rect 1267 1345 1268 1349
rect 1262 1344 1268 1345
rect 1422 1349 1428 1350
rect 1422 1345 1423 1349
rect 1427 1345 1428 1349
rect 1422 1344 1428 1345
rect 1582 1349 1588 1350
rect 1582 1345 1583 1349
rect 1587 1345 1588 1349
rect 1582 1344 1588 1345
rect 1750 1349 1756 1350
rect 1750 1345 1751 1349
rect 1755 1345 1756 1349
rect 1750 1344 1756 1345
rect 1902 1349 1908 1350
rect 1902 1345 1903 1349
rect 1907 1345 1908 1349
rect 1902 1344 1908 1345
rect 2006 1348 2012 1349
rect 2006 1344 2007 1348
rect 2011 1344 2012 1348
rect 2070 1345 2076 1346
rect 110 1343 116 1344
rect 2006 1343 2012 1344
rect 2046 1344 2052 1345
rect 2046 1340 2047 1344
rect 2051 1340 2052 1344
rect 2070 1341 2071 1345
rect 2075 1341 2076 1345
rect 2070 1340 2076 1341
rect 2302 1345 2308 1346
rect 2302 1341 2303 1345
rect 2307 1341 2308 1345
rect 2302 1340 2308 1341
rect 2558 1345 2564 1346
rect 2558 1341 2559 1345
rect 2563 1341 2564 1345
rect 2558 1340 2564 1341
rect 2806 1345 2812 1346
rect 2806 1341 2807 1345
rect 2811 1341 2812 1345
rect 2806 1340 2812 1341
rect 3054 1345 3060 1346
rect 3054 1341 3055 1345
rect 3059 1341 3060 1345
rect 3054 1340 3060 1341
rect 3302 1345 3308 1346
rect 3302 1341 3303 1345
rect 3307 1341 3308 1345
rect 3302 1340 3308 1341
rect 3558 1345 3564 1346
rect 3558 1341 3559 1345
rect 3563 1341 3564 1345
rect 3558 1340 3564 1341
rect 3814 1345 3820 1346
rect 3814 1341 3815 1345
rect 3819 1341 3820 1345
rect 3814 1340 3820 1341
rect 3942 1344 3948 1345
rect 3942 1340 3943 1344
rect 3947 1340 3948 1344
rect 2046 1339 2052 1340
rect 3942 1339 3948 1340
rect 110 1288 116 1289
rect 2006 1288 2012 1289
rect 110 1284 111 1288
rect 115 1284 116 1288
rect 110 1283 116 1284
rect 550 1287 556 1288
rect 550 1283 551 1287
rect 555 1283 556 1287
rect 550 1282 556 1283
rect 654 1287 660 1288
rect 654 1283 655 1287
rect 659 1283 660 1287
rect 654 1282 660 1283
rect 766 1287 772 1288
rect 766 1283 767 1287
rect 771 1283 772 1287
rect 766 1282 772 1283
rect 878 1287 884 1288
rect 878 1283 879 1287
rect 883 1283 884 1287
rect 878 1282 884 1283
rect 990 1287 996 1288
rect 990 1283 991 1287
rect 995 1283 996 1287
rect 990 1282 996 1283
rect 1102 1287 1108 1288
rect 1102 1283 1103 1287
rect 1107 1283 1108 1287
rect 1102 1282 1108 1283
rect 1214 1287 1220 1288
rect 1214 1283 1215 1287
rect 1219 1283 1220 1287
rect 1214 1282 1220 1283
rect 1326 1287 1332 1288
rect 1326 1283 1327 1287
rect 1331 1283 1332 1287
rect 1326 1282 1332 1283
rect 1438 1287 1444 1288
rect 1438 1283 1439 1287
rect 1443 1283 1444 1287
rect 1438 1282 1444 1283
rect 1558 1287 1564 1288
rect 1558 1283 1559 1287
rect 1563 1283 1564 1287
rect 2006 1284 2007 1288
rect 2011 1284 2012 1288
rect 2006 1283 2012 1284
rect 2046 1284 2052 1285
rect 3942 1284 3948 1285
rect 1558 1282 1564 1283
rect 2046 1280 2047 1284
rect 2051 1280 2052 1284
rect 2046 1279 2052 1280
rect 2070 1283 2076 1284
rect 2070 1279 2071 1283
rect 2075 1279 2076 1283
rect 2070 1278 2076 1279
rect 2222 1283 2228 1284
rect 2222 1279 2223 1283
rect 2227 1279 2228 1283
rect 2222 1278 2228 1279
rect 2414 1283 2420 1284
rect 2414 1279 2415 1283
rect 2419 1279 2420 1283
rect 2414 1278 2420 1279
rect 2614 1283 2620 1284
rect 2614 1279 2615 1283
rect 2619 1279 2620 1283
rect 2614 1278 2620 1279
rect 2814 1283 2820 1284
rect 2814 1279 2815 1283
rect 2819 1279 2820 1283
rect 2814 1278 2820 1279
rect 2998 1283 3004 1284
rect 2998 1279 2999 1283
rect 3003 1279 3004 1283
rect 2998 1278 3004 1279
rect 3174 1283 3180 1284
rect 3174 1279 3175 1283
rect 3179 1279 3180 1283
rect 3174 1278 3180 1279
rect 3342 1283 3348 1284
rect 3342 1279 3343 1283
rect 3347 1279 3348 1283
rect 3342 1278 3348 1279
rect 3502 1283 3508 1284
rect 3502 1279 3503 1283
rect 3507 1279 3508 1283
rect 3502 1278 3508 1279
rect 3662 1283 3668 1284
rect 3662 1279 3663 1283
rect 3667 1279 3668 1283
rect 3662 1278 3668 1279
rect 3830 1283 3836 1284
rect 3830 1279 3831 1283
rect 3835 1279 3836 1283
rect 3942 1280 3943 1284
rect 3947 1280 3948 1284
rect 3942 1279 3948 1280
rect 3830 1278 3836 1279
rect 110 1271 116 1272
rect 110 1267 111 1271
rect 115 1267 116 1271
rect 2006 1271 2012 1272
rect 110 1266 116 1267
rect 550 1268 556 1269
rect 550 1264 551 1268
rect 555 1264 556 1268
rect 550 1263 556 1264
rect 654 1268 660 1269
rect 654 1264 655 1268
rect 659 1264 660 1268
rect 654 1263 660 1264
rect 766 1268 772 1269
rect 766 1264 767 1268
rect 771 1264 772 1268
rect 766 1263 772 1264
rect 878 1268 884 1269
rect 878 1264 879 1268
rect 883 1264 884 1268
rect 878 1263 884 1264
rect 990 1268 996 1269
rect 990 1264 991 1268
rect 995 1264 996 1268
rect 990 1263 996 1264
rect 1102 1268 1108 1269
rect 1102 1264 1103 1268
rect 1107 1264 1108 1268
rect 1102 1263 1108 1264
rect 1214 1268 1220 1269
rect 1214 1264 1215 1268
rect 1219 1264 1220 1268
rect 1214 1263 1220 1264
rect 1326 1268 1332 1269
rect 1326 1264 1327 1268
rect 1331 1264 1332 1268
rect 1326 1263 1332 1264
rect 1438 1268 1444 1269
rect 1438 1264 1439 1268
rect 1443 1264 1444 1268
rect 1438 1263 1444 1264
rect 1558 1268 1564 1269
rect 1558 1264 1559 1268
rect 1563 1264 1564 1268
rect 2006 1267 2007 1271
rect 2011 1267 2012 1271
rect 2006 1266 2012 1267
rect 2046 1267 2052 1268
rect 1558 1263 1564 1264
rect 2046 1263 2047 1267
rect 2051 1263 2052 1267
rect 3942 1267 3948 1268
rect 2046 1262 2052 1263
rect 2070 1264 2076 1265
rect 2070 1260 2071 1264
rect 2075 1260 2076 1264
rect 2070 1259 2076 1260
rect 2222 1264 2228 1265
rect 2222 1260 2223 1264
rect 2227 1260 2228 1264
rect 2222 1259 2228 1260
rect 2414 1264 2420 1265
rect 2414 1260 2415 1264
rect 2419 1260 2420 1264
rect 2414 1259 2420 1260
rect 2614 1264 2620 1265
rect 2614 1260 2615 1264
rect 2619 1260 2620 1264
rect 2614 1259 2620 1260
rect 2814 1264 2820 1265
rect 2814 1260 2815 1264
rect 2819 1260 2820 1264
rect 2814 1259 2820 1260
rect 2998 1264 3004 1265
rect 2998 1260 2999 1264
rect 3003 1260 3004 1264
rect 2998 1259 3004 1260
rect 3174 1264 3180 1265
rect 3174 1260 3175 1264
rect 3179 1260 3180 1264
rect 3174 1259 3180 1260
rect 3342 1264 3348 1265
rect 3342 1260 3343 1264
rect 3347 1260 3348 1264
rect 3342 1259 3348 1260
rect 3502 1264 3508 1265
rect 3502 1260 3503 1264
rect 3507 1260 3508 1264
rect 3502 1259 3508 1260
rect 3662 1264 3668 1265
rect 3662 1260 3663 1264
rect 3667 1260 3668 1264
rect 3662 1259 3668 1260
rect 3830 1264 3836 1265
rect 3830 1260 3831 1264
rect 3835 1260 3836 1264
rect 3942 1263 3943 1267
rect 3947 1263 3948 1267
rect 3942 1262 3948 1263
rect 3830 1259 3836 1260
rect 390 1208 396 1209
rect 110 1205 116 1206
rect 110 1201 111 1205
rect 115 1201 116 1205
rect 390 1204 391 1208
rect 395 1204 396 1208
rect 390 1203 396 1204
rect 518 1208 524 1209
rect 518 1204 519 1208
rect 523 1204 524 1208
rect 518 1203 524 1204
rect 662 1208 668 1209
rect 662 1204 663 1208
rect 667 1204 668 1208
rect 662 1203 668 1204
rect 806 1208 812 1209
rect 806 1204 807 1208
rect 811 1204 812 1208
rect 806 1203 812 1204
rect 958 1208 964 1209
rect 958 1204 959 1208
rect 963 1204 964 1208
rect 958 1203 964 1204
rect 1110 1208 1116 1209
rect 1110 1204 1111 1208
rect 1115 1204 1116 1208
rect 1110 1203 1116 1204
rect 1254 1208 1260 1209
rect 1254 1204 1255 1208
rect 1259 1204 1260 1208
rect 1254 1203 1260 1204
rect 1406 1208 1412 1209
rect 1406 1204 1407 1208
rect 1411 1204 1412 1208
rect 1406 1203 1412 1204
rect 1558 1208 1564 1209
rect 1558 1204 1559 1208
rect 1563 1204 1564 1208
rect 1558 1203 1564 1204
rect 1710 1208 1716 1209
rect 1710 1204 1711 1208
rect 1715 1204 1716 1208
rect 1710 1203 1716 1204
rect 2006 1205 2012 1206
rect 110 1200 116 1201
rect 2006 1201 2007 1205
rect 2011 1201 2012 1205
rect 2006 1200 2012 1201
rect 2134 1196 2140 1197
rect 2046 1193 2052 1194
rect 390 1189 396 1190
rect 110 1188 116 1189
rect 110 1184 111 1188
rect 115 1184 116 1188
rect 390 1185 391 1189
rect 395 1185 396 1189
rect 390 1184 396 1185
rect 518 1189 524 1190
rect 518 1185 519 1189
rect 523 1185 524 1189
rect 518 1184 524 1185
rect 662 1189 668 1190
rect 662 1185 663 1189
rect 667 1185 668 1189
rect 662 1184 668 1185
rect 806 1189 812 1190
rect 806 1185 807 1189
rect 811 1185 812 1189
rect 806 1184 812 1185
rect 958 1189 964 1190
rect 958 1185 959 1189
rect 963 1185 964 1189
rect 958 1184 964 1185
rect 1110 1189 1116 1190
rect 1110 1185 1111 1189
rect 1115 1185 1116 1189
rect 1110 1184 1116 1185
rect 1254 1189 1260 1190
rect 1254 1185 1255 1189
rect 1259 1185 1260 1189
rect 1254 1184 1260 1185
rect 1406 1189 1412 1190
rect 1406 1185 1407 1189
rect 1411 1185 1412 1189
rect 1406 1184 1412 1185
rect 1558 1189 1564 1190
rect 1558 1185 1559 1189
rect 1563 1185 1564 1189
rect 1558 1184 1564 1185
rect 1710 1189 1716 1190
rect 2046 1189 2047 1193
rect 2051 1189 2052 1193
rect 2134 1192 2135 1196
rect 2139 1192 2140 1196
rect 2134 1191 2140 1192
rect 2310 1196 2316 1197
rect 2310 1192 2311 1196
rect 2315 1192 2316 1196
rect 2310 1191 2316 1192
rect 2502 1196 2508 1197
rect 2502 1192 2503 1196
rect 2507 1192 2508 1196
rect 2502 1191 2508 1192
rect 2694 1196 2700 1197
rect 2694 1192 2695 1196
rect 2699 1192 2700 1196
rect 2694 1191 2700 1192
rect 2886 1196 2892 1197
rect 2886 1192 2887 1196
rect 2891 1192 2892 1196
rect 2886 1191 2892 1192
rect 3070 1196 3076 1197
rect 3070 1192 3071 1196
rect 3075 1192 3076 1196
rect 3070 1191 3076 1192
rect 3238 1196 3244 1197
rect 3238 1192 3239 1196
rect 3243 1192 3244 1196
rect 3238 1191 3244 1192
rect 3398 1196 3404 1197
rect 3398 1192 3399 1196
rect 3403 1192 3404 1196
rect 3398 1191 3404 1192
rect 3550 1196 3556 1197
rect 3550 1192 3551 1196
rect 3555 1192 3556 1196
rect 3550 1191 3556 1192
rect 3702 1196 3708 1197
rect 3702 1192 3703 1196
rect 3707 1192 3708 1196
rect 3702 1191 3708 1192
rect 3838 1196 3844 1197
rect 3838 1192 3839 1196
rect 3843 1192 3844 1196
rect 3838 1191 3844 1192
rect 3942 1193 3948 1194
rect 1710 1185 1711 1189
rect 1715 1185 1716 1189
rect 1710 1184 1716 1185
rect 2006 1188 2012 1189
rect 2046 1188 2052 1189
rect 3942 1189 3943 1193
rect 3947 1189 3948 1193
rect 3942 1188 3948 1189
rect 2006 1184 2007 1188
rect 2011 1184 2012 1188
rect 110 1183 116 1184
rect 2006 1183 2012 1184
rect 2134 1177 2140 1178
rect 2046 1176 2052 1177
rect 2046 1172 2047 1176
rect 2051 1172 2052 1176
rect 2134 1173 2135 1177
rect 2139 1173 2140 1177
rect 2134 1172 2140 1173
rect 2310 1177 2316 1178
rect 2310 1173 2311 1177
rect 2315 1173 2316 1177
rect 2310 1172 2316 1173
rect 2502 1177 2508 1178
rect 2502 1173 2503 1177
rect 2507 1173 2508 1177
rect 2502 1172 2508 1173
rect 2694 1177 2700 1178
rect 2694 1173 2695 1177
rect 2699 1173 2700 1177
rect 2694 1172 2700 1173
rect 2886 1177 2892 1178
rect 2886 1173 2887 1177
rect 2891 1173 2892 1177
rect 2886 1172 2892 1173
rect 3070 1177 3076 1178
rect 3070 1173 3071 1177
rect 3075 1173 3076 1177
rect 3070 1172 3076 1173
rect 3238 1177 3244 1178
rect 3238 1173 3239 1177
rect 3243 1173 3244 1177
rect 3238 1172 3244 1173
rect 3398 1177 3404 1178
rect 3398 1173 3399 1177
rect 3403 1173 3404 1177
rect 3398 1172 3404 1173
rect 3550 1177 3556 1178
rect 3550 1173 3551 1177
rect 3555 1173 3556 1177
rect 3550 1172 3556 1173
rect 3702 1177 3708 1178
rect 3702 1173 3703 1177
rect 3707 1173 3708 1177
rect 3702 1172 3708 1173
rect 3838 1177 3844 1178
rect 3838 1173 3839 1177
rect 3843 1173 3844 1177
rect 3838 1172 3844 1173
rect 3942 1176 3948 1177
rect 3942 1172 3943 1176
rect 3947 1172 3948 1176
rect 2046 1171 2052 1172
rect 3942 1171 3948 1172
rect 110 1132 116 1133
rect 2006 1132 2012 1133
rect 110 1128 111 1132
rect 115 1128 116 1132
rect 110 1127 116 1128
rect 174 1131 180 1132
rect 174 1127 175 1131
rect 179 1127 180 1131
rect 174 1126 180 1127
rect 326 1131 332 1132
rect 326 1127 327 1131
rect 331 1127 332 1131
rect 326 1126 332 1127
rect 494 1131 500 1132
rect 494 1127 495 1131
rect 499 1127 500 1131
rect 494 1126 500 1127
rect 670 1131 676 1132
rect 670 1127 671 1131
rect 675 1127 676 1131
rect 670 1126 676 1127
rect 846 1131 852 1132
rect 846 1127 847 1131
rect 851 1127 852 1131
rect 846 1126 852 1127
rect 1030 1131 1036 1132
rect 1030 1127 1031 1131
rect 1035 1127 1036 1131
rect 1030 1126 1036 1127
rect 1206 1131 1212 1132
rect 1206 1127 1207 1131
rect 1211 1127 1212 1131
rect 1206 1126 1212 1127
rect 1382 1131 1388 1132
rect 1382 1127 1383 1131
rect 1387 1127 1388 1131
rect 1382 1126 1388 1127
rect 1566 1131 1572 1132
rect 1566 1127 1567 1131
rect 1571 1127 1572 1131
rect 1566 1126 1572 1127
rect 1750 1131 1756 1132
rect 1750 1127 1751 1131
rect 1755 1127 1756 1131
rect 2006 1128 2007 1132
rect 2011 1128 2012 1132
rect 2006 1127 2012 1128
rect 1750 1126 1756 1127
rect 2046 1116 2052 1117
rect 3942 1116 3948 1117
rect 110 1115 116 1116
rect 110 1111 111 1115
rect 115 1111 116 1115
rect 2006 1115 2012 1116
rect 110 1110 116 1111
rect 174 1112 180 1113
rect 174 1108 175 1112
rect 179 1108 180 1112
rect 174 1107 180 1108
rect 326 1112 332 1113
rect 326 1108 327 1112
rect 331 1108 332 1112
rect 326 1107 332 1108
rect 494 1112 500 1113
rect 494 1108 495 1112
rect 499 1108 500 1112
rect 494 1107 500 1108
rect 670 1112 676 1113
rect 670 1108 671 1112
rect 675 1108 676 1112
rect 670 1107 676 1108
rect 846 1112 852 1113
rect 846 1108 847 1112
rect 851 1108 852 1112
rect 846 1107 852 1108
rect 1030 1112 1036 1113
rect 1030 1108 1031 1112
rect 1035 1108 1036 1112
rect 1030 1107 1036 1108
rect 1206 1112 1212 1113
rect 1206 1108 1207 1112
rect 1211 1108 1212 1112
rect 1206 1107 1212 1108
rect 1382 1112 1388 1113
rect 1382 1108 1383 1112
rect 1387 1108 1388 1112
rect 1382 1107 1388 1108
rect 1566 1112 1572 1113
rect 1566 1108 1567 1112
rect 1571 1108 1572 1112
rect 1566 1107 1572 1108
rect 1750 1112 1756 1113
rect 1750 1108 1751 1112
rect 1755 1108 1756 1112
rect 2006 1111 2007 1115
rect 2011 1111 2012 1115
rect 2046 1112 2047 1116
rect 2051 1112 2052 1116
rect 2046 1111 2052 1112
rect 2294 1115 2300 1116
rect 2294 1111 2295 1115
rect 2299 1111 2300 1115
rect 2006 1110 2012 1111
rect 2294 1110 2300 1111
rect 2422 1115 2428 1116
rect 2422 1111 2423 1115
rect 2427 1111 2428 1115
rect 2422 1110 2428 1111
rect 2558 1115 2564 1116
rect 2558 1111 2559 1115
rect 2563 1111 2564 1115
rect 2558 1110 2564 1111
rect 2694 1115 2700 1116
rect 2694 1111 2695 1115
rect 2699 1111 2700 1115
rect 2694 1110 2700 1111
rect 2838 1115 2844 1116
rect 2838 1111 2839 1115
rect 2843 1111 2844 1115
rect 2838 1110 2844 1111
rect 2990 1115 2996 1116
rect 2990 1111 2991 1115
rect 2995 1111 2996 1115
rect 2990 1110 2996 1111
rect 3150 1115 3156 1116
rect 3150 1111 3151 1115
rect 3155 1111 3156 1115
rect 3150 1110 3156 1111
rect 3318 1115 3324 1116
rect 3318 1111 3319 1115
rect 3323 1111 3324 1115
rect 3318 1110 3324 1111
rect 3494 1115 3500 1116
rect 3494 1111 3495 1115
rect 3499 1111 3500 1115
rect 3494 1110 3500 1111
rect 3678 1115 3684 1116
rect 3678 1111 3679 1115
rect 3683 1111 3684 1115
rect 3678 1110 3684 1111
rect 3838 1115 3844 1116
rect 3838 1111 3839 1115
rect 3843 1111 3844 1115
rect 3942 1112 3943 1116
rect 3947 1112 3948 1116
rect 3942 1111 3948 1112
rect 3838 1110 3844 1111
rect 1750 1107 1756 1108
rect 2046 1099 2052 1100
rect 2046 1095 2047 1099
rect 2051 1095 2052 1099
rect 3942 1099 3948 1100
rect 2046 1094 2052 1095
rect 2294 1096 2300 1097
rect 2294 1092 2295 1096
rect 2299 1092 2300 1096
rect 2294 1091 2300 1092
rect 2422 1096 2428 1097
rect 2422 1092 2423 1096
rect 2427 1092 2428 1096
rect 2422 1091 2428 1092
rect 2558 1096 2564 1097
rect 2558 1092 2559 1096
rect 2563 1092 2564 1096
rect 2558 1091 2564 1092
rect 2694 1096 2700 1097
rect 2694 1092 2695 1096
rect 2699 1092 2700 1096
rect 2694 1091 2700 1092
rect 2838 1096 2844 1097
rect 2838 1092 2839 1096
rect 2843 1092 2844 1096
rect 2838 1091 2844 1092
rect 2990 1096 2996 1097
rect 2990 1092 2991 1096
rect 2995 1092 2996 1096
rect 2990 1091 2996 1092
rect 3150 1096 3156 1097
rect 3150 1092 3151 1096
rect 3155 1092 3156 1096
rect 3150 1091 3156 1092
rect 3318 1096 3324 1097
rect 3318 1092 3319 1096
rect 3323 1092 3324 1096
rect 3318 1091 3324 1092
rect 3494 1096 3500 1097
rect 3494 1092 3495 1096
rect 3499 1092 3500 1096
rect 3494 1091 3500 1092
rect 3678 1096 3684 1097
rect 3678 1092 3679 1096
rect 3683 1092 3684 1096
rect 3678 1091 3684 1092
rect 3838 1096 3844 1097
rect 3838 1092 3839 1096
rect 3843 1092 3844 1096
rect 3942 1095 3943 1099
rect 3947 1095 3948 1099
rect 3942 1094 3948 1095
rect 3838 1091 3844 1092
rect 134 1044 140 1045
rect 110 1041 116 1042
rect 110 1037 111 1041
rect 115 1037 116 1041
rect 134 1040 135 1044
rect 139 1040 140 1044
rect 134 1039 140 1040
rect 230 1044 236 1045
rect 230 1040 231 1044
rect 235 1040 236 1044
rect 230 1039 236 1040
rect 374 1044 380 1045
rect 374 1040 375 1044
rect 379 1040 380 1044
rect 374 1039 380 1040
rect 542 1044 548 1045
rect 542 1040 543 1044
rect 547 1040 548 1044
rect 542 1039 548 1040
rect 726 1044 732 1045
rect 726 1040 727 1044
rect 731 1040 732 1044
rect 726 1039 732 1040
rect 910 1044 916 1045
rect 910 1040 911 1044
rect 915 1040 916 1044
rect 910 1039 916 1040
rect 1094 1044 1100 1045
rect 1094 1040 1095 1044
rect 1099 1040 1100 1044
rect 1094 1039 1100 1040
rect 1278 1044 1284 1045
rect 1278 1040 1279 1044
rect 1283 1040 1284 1044
rect 1278 1039 1284 1040
rect 1462 1044 1468 1045
rect 1462 1040 1463 1044
rect 1467 1040 1468 1044
rect 1462 1039 1468 1040
rect 1646 1044 1652 1045
rect 1646 1040 1647 1044
rect 1651 1040 1652 1044
rect 1646 1039 1652 1040
rect 1830 1044 1836 1045
rect 1830 1040 1831 1044
rect 1835 1040 1836 1044
rect 1830 1039 1836 1040
rect 2006 1041 2012 1042
rect 110 1036 116 1037
rect 2006 1037 2007 1041
rect 2011 1037 2012 1041
rect 2006 1036 2012 1037
rect 2494 1032 2500 1033
rect 2046 1029 2052 1030
rect 134 1025 140 1026
rect 110 1024 116 1025
rect 110 1020 111 1024
rect 115 1020 116 1024
rect 134 1021 135 1025
rect 139 1021 140 1025
rect 134 1020 140 1021
rect 230 1025 236 1026
rect 230 1021 231 1025
rect 235 1021 236 1025
rect 230 1020 236 1021
rect 374 1025 380 1026
rect 374 1021 375 1025
rect 379 1021 380 1025
rect 374 1020 380 1021
rect 542 1025 548 1026
rect 542 1021 543 1025
rect 547 1021 548 1025
rect 542 1020 548 1021
rect 726 1025 732 1026
rect 726 1021 727 1025
rect 731 1021 732 1025
rect 726 1020 732 1021
rect 910 1025 916 1026
rect 910 1021 911 1025
rect 915 1021 916 1025
rect 910 1020 916 1021
rect 1094 1025 1100 1026
rect 1094 1021 1095 1025
rect 1099 1021 1100 1025
rect 1094 1020 1100 1021
rect 1278 1025 1284 1026
rect 1278 1021 1279 1025
rect 1283 1021 1284 1025
rect 1278 1020 1284 1021
rect 1462 1025 1468 1026
rect 1462 1021 1463 1025
rect 1467 1021 1468 1025
rect 1462 1020 1468 1021
rect 1646 1025 1652 1026
rect 1646 1021 1647 1025
rect 1651 1021 1652 1025
rect 1646 1020 1652 1021
rect 1830 1025 1836 1026
rect 2046 1025 2047 1029
rect 2051 1025 2052 1029
rect 2494 1028 2495 1032
rect 2499 1028 2500 1032
rect 2494 1027 2500 1028
rect 2598 1032 2604 1033
rect 2598 1028 2599 1032
rect 2603 1028 2604 1032
rect 2598 1027 2604 1028
rect 2710 1032 2716 1033
rect 2710 1028 2711 1032
rect 2715 1028 2716 1032
rect 2710 1027 2716 1028
rect 2846 1032 2852 1033
rect 2846 1028 2847 1032
rect 2851 1028 2852 1032
rect 2846 1027 2852 1028
rect 3006 1032 3012 1033
rect 3006 1028 3007 1032
rect 3011 1028 3012 1032
rect 3006 1027 3012 1028
rect 3198 1032 3204 1033
rect 3198 1028 3199 1032
rect 3203 1028 3204 1032
rect 3198 1027 3204 1028
rect 3406 1032 3412 1033
rect 3406 1028 3407 1032
rect 3411 1028 3412 1032
rect 3406 1027 3412 1028
rect 3630 1032 3636 1033
rect 3630 1028 3631 1032
rect 3635 1028 3636 1032
rect 3630 1027 3636 1028
rect 3838 1032 3844 1033
rect 3838 1028 3839 1032
rect 3843 1028 3844 1032
rect 3838 1027 3844 1028
rect 3942 1029 3948 1030
rect 1830 1021 1831 1025
rect 1835 1021 1836 1025
rect 1830 1020 1836 1021
rect 2006 1024 2012 1025
rect 2046 1024 2052 1025
rect 3942 1025 3943 1029
rect 3947 1025 3948 1029
rect 3942 1024 3948 1025
rect 2006 1020 2007 1024
rect 2011 1020 2012 1024
rect 110 1019 116 1020
rect 2006 1019 2012 1020
rect 2494 1013 2500 1014
rect 2046 1012 2052 1013
rect 2046 1008 2047 1012
rect 2051 1008 2052 1012
rect 2494 1009 2495 1013
rect 2499 1009 2500 1013
rect 2494 1008 2500 1009
rect 2598 1013 2604 1014
rect 2598 1009 2599 1013
rect 2603 1009 2604 1013
rect 2598 1008 2604 1009
rect 2710 1013 2716 1014
rect 2710 1009 2711 1013
rect 2715 1009 2716 1013
rect 2710 1008 2716 1009
rect 2846 1013 2852 1014
rect 2846 1009 2847 1013
rect 2851 1009 2852 1013
rect 2846 1008 2852 1009
rect 3006 1013 3012 1014
rect 3006 1009 3007 1013
rect 3011 1009 3012 1013
rect 3006 1008 3012 1009
rect 3198 1013 3204 1014
rect 3198 1009 3199 1013
rect 3203 1009 3204 1013
rect 3198 1008 3204 1009
rect 3406 1013 3412 1014
rect 3406 1009 3407 1013
rect 3411 1009 3412 1013
rect 3406 1008 3412 1009
rect 3630 1013 3636 1014
rect 3630 1009 3631 1013
rect 3635 1009 3636 1013
rect 3630 1008 3636 1009
rect 3838 1013 3844 1014
rect 3838 1009 3839 1013
rect 3843 1009 3844 1013
rect 3838 1008 3844 1009
rect 3942 1012 3948 1013
rect 3942 1008 3943 1012
rect 3947 1008 3948 1012
rect 2046 1007 2052 1008
rect 3942 1007 3948 1008
rect 110 972 116 973
rect 2006 972 2012 973
rect 110 968 111 972
rect 115 968 116 972
rect 110 967 116 968
rect 134 971 140 972
rect 134 967 135 971
rect 139 967 140 971
rect 134 966 140 967
rect 270 971 276 972
rect 270 967 271 971
rect 275 967 276 971
rect 270 966 276 967
rect 446 971 452 972
rect 446 967 447 971
rect 451 967 452 971
rect 446 966 452 967
rect 630 971 636 972
rect 630 967 631 971
rect 635 967 636 971
rect 630 966 636 967
rect 822 971 828 972
rect 822 967 823 971
rect 827 967 828 971
rect 822 966 828 967
rect 1006 971 1012 972
rect 1006 967 1007 971
rect 1011 967 1012 971
rect 1006 966 1012 967
rect 1174 971 1180 972
rect 1174 967 1175 971
rect 1179 967 1180 971
rect 1174 966 1180 967
rect 1334 971 1340 972
rect 1334 967 1335 971
rect 1339 967 1340 971
rect 1334 966 1340 967
rect 1486 971 1492 972
rect 1486 967 1487 971
rect 1491 967 1492 971
rect 1486 966 1492 967
rect 1630 971 1636 972
rect 1630 967 1631 971
rect 1635 967 1636 971
rect 1630 966 1636 967
rect 1774 971 1780 972
rect 1774 967 1775 971
rect 1779 967 1780 971
rect 1774 966 1780 967
rect 1902 971 1908 972
rect 1902 967 1903 971
rect 1907 967 1908 971
rect 2006 968 2007 972
rect 2011 968 2012 972
rect 2006 967 2012 968
rect 1902 966 1908 967
rect 2046 960 2052 961
rect 3942 960 3948 961
rect 2046 956 2047 960
rect 2051 956 2052 960
rect 110 955 116 956
rect 110 951 111 955
rect 115 951 116 955
rect 2006 955 2012 956
rect 2046 955 2052 956
rect 2646 959 2652 960
rect 2646 955 2647 959
rect 2651 955 2652 959
rect 110 950 116 951
rect 134 952 140 953
rect 134 948 135 952
rect 139 948 140 952
rect 134 947 140 948
rect 270 952 276 953
rect 270 948 271 952
rect 275 948 276 952
rect 270 947 276 948
rect 446 952 452 953
rect 446 948 447 952
rect 451 948 452 952
rect 446 947 452 948
rect 630 952 636 953
rect 630 948 631 952
rect 635 948 636 952
rect 630 947 636 948
rect 822 952 828 953
rect 822 948 823 952
rect 827 948 828 952
rect 822 947 828 948
rect 1006 952 1012 953
rect 1006 948 1007 952
rect 1011 948 1012 952
rect 1006 947 1012 948
rect 1174 952 1180 953
rect 1174 948 1175 952
rect 1179 948 1180 952
rect 1174 947 1180 948
rect 1334 952 1340 953
rect 1334 948 1335 952
rect 1339 948 1340 952
rect 1334 947 1340 948
rect 1486 952 1492 953
rect 1486 948 1487 952
rect 1491 948 1492 952
rect 1486 947 1492 948
rect 1630 952 1636 953
rect 1630 948 1631 952
rect 1635 948 1636 952
rect 1630 947 1636 948
rect 1774 952 1780 953
rect 1774 948 1775 952
rect 1779 948 1780 952
rect 1774 947 1780 948
rect 1902 952 1908 953
rect 1902 948 1903 952
rect 1907 948 1908 952
rect 2006 951 2007 955
rect 2011 951 2012 955
rect 2646 954 2652 955
rect 2742 959 2748 960
rect 2742 955 2743 959
rect 2747 955 2748 959
rect 2742 954 2748 955
rect 2846 959 2852 960
rect 2846 955 2847 959
rect 2851 955 2852 959
rect 2846 954 2852 955
rect 2966 959 2972 960
rect 2966 955 2967 959
rect 2971 955 2972 959
rect 2966 954 2972 955
rect 3110 959 3116 960
rect 3110 955 3111 959
rect 3115 955 3116 959
rect 3110 954 3116 955
rect 3278 959 3284 960
rect 3278 955 3279 959
rect 3283 955 3284 959
rect 3278 954 3284 955
rect 3462 959 3468 960
rect 3462 955 3463 959
rect 3467 955 3468 959
rect 3462 954 3468 955
rect 3662 959 3668 960
rect 3662 955 3663 959
rect 3667 955 3668 959
rect 3662 954 3668 955
rect 3838 959 3844 960
rect 3838 955 3839 959
rect 3843 955 3844 959
rect 3942 956 3943 960
rect 3947 956 3948 960
rect 3942 955 3948 956
rect 3838 954 3844 955
rect 2006 950 2012 951
rect 1902 947 1908 948
rect 2046 943 2052 944
rect 2046 939 2047 943
rect 2051 939 2052 943
rect 3942 943 3948 944
rect 2046 938 2052 939
rect 2646 940 2652 941
rect 2646 936 2647 940
rect 2651 936 2652 940
rect 2646 935 2652 936
rect 2742 940 2748 941
rect 2742 936 2743 940
rect 2747 936 2748 940
rect 2742 935 2748 936
rect 2846 940 2852 941
rect 2846 936 2847 940
rect 2851 936 2852 940
rect 2846 935 2852 936
rect 2966 940 2972 941
rect 2966 936 2967 940
rect 2971 936 2972 940
rect 2966 935 2972 936
rect 3110 940 3116 941
rect 3110 936 3111 940
rect 3115 936 3116 940
rect 3110 935 3116 936
rect 3278 940 3284 941
rect 3278 936 3279 940
rect 3283 936 3284 940
rect 3278 935 3284 936
rect 3462 940 3468 941
rect 3462 936 3463 940
rect 3467 936 3468 940
rect 3462 935 3468 936
rect 3662 940 3668 941
rect 3662 936 3663 940
rect 3667 936 3668 940
rect 3662 935 3668 936
rect 3838 940 3844 941
rect 3838 936 3839 940
rect 3843 936 3844 940
rect 3942 939 3943 943
rect 3947 939 3948 943
rect 3942 938 3948 939
rect 3838 935 3844 936
rect 134 892 140 893
rect 110 889 116 890
rect 110 885 111 889
rect 115 885 116 889
rect 134 888 135 892
rect 139 888 140 892
rect 134 887 140 888
rect 270 892 276 893
rect 270 888 271 892
rect 275 888 276 892
rect 270 887 276 888
rect 454 892 460 893
rect 454 888 455 892
rect 459 888 460 892
rect 454 887 460 888
rect 654 892 660 893
rect 654 888 655 892
rect 659 888 660 892
rect 654 887 660 888
rect 854 892 860 893
rect 854 888 855 892
rect 859 888 860 892
rect 854 887 860 888
rect 1054 892 1060 893
rect 1054 888 1055 892
rect 1059 888 1060 892
rect 1054 887 1060 888
rect 1238 892 1244 893
rect 1238 888 1239 892
rect 1243 888 1244 892
rect 1238 887 1244 888
rect 1414 892 1420 893
rect 1414 888 1415 892
rect 1419 888 1420 892
rect 1414 887 1420 888
rect 1582 892 1588 893
rect 1582 888 1583 892
rect 1587 888 1588 892
rect 1582 887 1588 888
rect 1750 892 1756 893
rect 1750 888 1751 892
rect 1755 888 1756 892
rect 1750 887 1756 888
rect 1902 892 1908 893
rect 1902 888 1903 892
rect 1907 888 1908 892
rect 1902 887 1908 888
rect 2006 889 2012 890
rect 110 884 116 885
rect 2006 885 2007 889
rect 2011 885 2012 889
rect 2006 884 2012 885
rect 134 873 140 874
rect 110 872 116 873
rect 110 868 111 872
rect 115 868 116 872
rect 134 869 135 873
rect 139 869 140 873
rect 134 868 140 869
rect 270 873 276 874
rect 270 869 271 873
rect 275 869 276 873
rect 270 868 276 869
rect 454 873 460 874
rect 454 869 455 873
rect 459 869 460 873
rect 454 868 460 869
rect 654 873 660 874
rect 654 869 655 873
rect 659 869 660 873
rect 654 868 660 869
rect 854 873 860 874
rect 854 869 855 873
rect 859 869 860 873
rect 854 868 860 869
rect 1054 873 1060 874
rect 1054 869 1055 873
rect 1059 869 1060 873
rect 1054 868 1060 869
rect 1238 873 1244 874
rect 1238 869 1239 873
rect 1243 869 1244 873
rect 1238 868 1244 869
rect 1414 873 1420 874
rect 1414 869 1415 873
rect 1419 869 1420 873
rect 1414 868 1420 869
rect 1582 873 1588 874
rect 1582 869 1583 873
rect 1587 869 1588 873
rect 1582 868 1588 869
rect 1750 873 1756 874
rect 1750 869 1751 873
rect 1755 869 1756 873
rect 1750 868 1756 869
rect 1902 873 1908 874
rect 1902 869 1903 873
rect 1907 869 1908 873
rect 1902 868 1908 869
rect 2006 872 2012 873
rect 2006 868 2007 872
rect 2011 868 2012 872
rect 110 867 116 868
rect 2006 867 2012 868
rect 2070 868 2076 869
rect 2046 865 2052 866
rect 2046 861 2047 865
rect 2051 861 2052 865
rect 2070 864 2071 868
rect 2075 864 2076 868
rect 2070 863 2076 864
rect 2254 868 2260 869
rect 2254 864 2255 868
rect 2259 864 2260 868
rect 2254 863 2260 864
rect 2462 868 2468 869
rect 2462 864 2463 868
rect 2467 864 2468 868
rect 2462 863 2468 864
rect 2678 868 2684 869
rect 2678 864 2679 868
rect 2683 864 2684 868
rect 2678 863 2684 864
rect 2894 868 2900 869
rect 2894 864 2895 868
rect 2899 864 2900 868
rect 2894 863 2900 864
rect 3126 868 3132 869
rect 3126 864 3127 868
rect 3131 864 3132 868
rect 3126 863 3132 864
rect 3366 868 3372 869
rect 3366 864 3367 868
rect 3371 864 3372 868
rect 3366 863 3372 864
rect 3614 868 3620 869
rect 3614 864 3615 868
rect 3619 864 3620 868
rect 3614 863 3620 864
rect 3838 868 3844 869
rect 3838 864 3839 868
rect 3843 864 3844 868
rect 3838 863 3844 864
rect 3942 865 3948 866
rect 2046 860 2052 861
rect 3942 861 3943 865
rect 3947 861 3948 865
rect 3942 860 3948 861
rect 2070 849 2076 850
rect 2046 848 2052 849
rect 2046 844 2047 848
rect 2051 844 2052 848
rect 2070 845 2071 849
rect 2075 845 2076 849
rect 2070 844 2076 845
rect 2254 849 2260 850
rect 2254 845 2255 849
rect 2259 845 2260 849
rect 2254 844 2260 845
rect 2462 849 2468 850
rect 2462 845 2463 849
rect 2467 845 2468 849
rect 2462 844 2468 845
rect 2678 849 2684 850
rect 2678 845 2679 849
rect 2683 845 2684 849
rect 2678 844 2684 845
rect 2894 849 2900 850
rect 2894 845 2895 849
rect 2899 845 2900 849
rect 2894 844 2900 845
rect 3126 849 3132 850
rect 3126 845 3127 849
rect 3131 845 3132 849
rect 3126 844 3132 845
rect 3366 849 3372 850
rect 3366 845 3367 849
rect 3371 845 3372 849
rect 3366 844 3372 845
rect 3614 849 3620 850
rect 3614 845 3615 849
rect 3619 845 3620 849
rect 3614 844 3620 845
rect 3838 849 3844 850
rect 3838 845 3839 849
rect 3843 845 3844 849
rect 3838 844 3844 845
rect 3942 848 3948 849
rect 3942 844 3943 848
rect 3947 844 3948 848
rect 2046 843 2052 844
rect 3942 843 3948 844
rect 110 820 116 821
rect 2006 820 2012 821
rect 110 816 111 820
rect 115 816 116 820
rect 110 815 116 816
rect 214 819 220 820
rect 214 815 215 819
rect 219 815 220 819
rect 214 814 220 815
rect 342 819 348 820
rect 342 815 343 819
rect 347 815 348 819
rect 342 814 348 815
rect 494 819 500 820
rect 494 815 495 819
rect 499 815 500 819
rect 494 814 500 815
rect 654 819 660 820
rect 654 815 655 819
rect 659 815 660 819
rect 654 814 660 815
rect 830 819 836 820
rect 830 815 831 819
rect 835 815 836 819
rect 830 814 836 815
rect 1006 819 1012 820
rect 1006 815 1007 819
rect 1011 815 1012 819
rect 1006 814 1012 815
rect 1182 819 1188 820
rect 1182 815 1183 819
rect 1187 815 1188 819
rect 1182 814 1188 815
rect 1358 819 1364 820
rect 1358 815 1359 819
rect 1363 815 1364 819
rect 1358 814 1364 815
rect 1534 819 1540 820
rect 1534 815 1535 819
rect 1539 815 1540 819
rect 1534 814 1540 815
rect 1718 819 1724 820
rect 1718 815 1719 819
rect 1723 815 1724 819
rect 2006 816 2007 820
rect 2011 816 2012 820
rect 2006 815 2012 816
rect 1718 814 1724 815
rect 110 803 116 804
rect 110 799 111 803
rect 115 799 116 803
rect 2006 803 2012 804
rect 110 798 116 799
rect 214 800 220 801
rect 214 796 215 800
rect 219 796 220 800
rect 214 795 220 796
rect 342 800 348 801
rect 342 796 343 800
rect 347 796 348 800
rect 342 795 348 796
rect 494 800 500 801
rect 494 796 495 800
rect 499 796 500 800
rect 494 795 500 796
rect 654 800 660 801
rect 654 796 655 800
rect 659 796 660 800
rect 654 795 660 796
rect 830 800 836 801
rect 830 796 831 800
rect 835 796 836 800
rect 830 795 836 796
rect 1006 800 1012 801
rect 1006 796 1007 800
rect 1011 796 1012 800
rect 1006 795 1012 796
rect 1182 800 1188 801
rect 1182 796 1183 800
rect 1187 796 1188 800
rect 1182 795 1188 796
rect 1358 800 1364 801
rect 1358 796 1359 800
rect 1363 796 1364 800
rect 1358 795 1364 796
rect 1534 800 1540 801
rect 1534 796 1535 800
rect 1539 796 1540 800
rect 1534 795 1540 796
rect 1718 800 1724 801
rect 1718 796 1719 800
rect 1723 796 1724 800
rect 2006 799 2007 803
rect 2011 799 2012 803
rect 2006 798 2012 799
rect 1718 795 1724 796
rect 2046 796 2052 797
rect 3942 796 3948 797
rect 2046 792 2047 796
rect 2051 792 2052 796
rect 2046 791 2052 792
rect 2214 795 2220 796
rect 2214 791 2215 795
rect 2219 791 2220 795
rect 2214 790 2220 791
rect 2326 795 2332 796
rect 2326 791 2327 795
rect 2331 791 2332 795
rect 2326 790 2332 791
rect 2446 795 2452 796
rect 2446 791 2447 795
rect 2451 791 2452 795
rect 2446 790 2452 791
rect 2582 795 2588 796
rect 2582 791 2583 795
rect 2587 791 2588 795
rect 2582 790 2588 791
rect 2734 795 2740 796
rect 2734 791 2735 795
rect 2739 791 2740 795
rect 2734 790 2740 791
rect 2894 795 2900 796
rect 2894 791 2895 795
rect 2899 791 2900 795
rect 2894 790 2900 791
rect 3062 795 3068 796
rect 3062 791 3063 795
rect 3067 791 3068 795
rect 3062 790 3068 791
rect 3246 795 3252 796
rect 3246 791 3247 795
rect 3251 791 3252 795
rect 3246 790 3252 791
rect 3446 795 3452 796
rect 3446 791 3447 795
rect 3451 791 3452 795
rect 3446 790 3452 791
rect 3654 795 3660 796
rect 3654 791 3655 795
rect 3659 791 3660 795
rect 3654 790 3660 791
rect 3838 795 3844 796
rect 3838 791 3839 795
rect 3843 791 3844 795
rect 3942 792 3943 796
rect 3947 792 3948 796
rect 3942 791 3948 792
rect 3838 790 3844 791
rect 2046 779 2052 780
rect 2046 775 2047 779
rect 2051 775 2052 779
rect 3942 779 3948 780
rect 2046 774 2052 775
rect 2214 776 2220 777
rect 2214 772 2215 776
rect 2219 772 2220 776
rect 2214 771 2220 772
rect 2326 776 2332 777
rect 2326 772 2327 776
rect 2331 772 2332 776
rect 2326 771 2332 772
rect 2446 776 2452 777
rect 2446 772 2447 776
rect 2451 772 2452 776
rect 2446 771 2452 772
rect 2582 776 2588 777
rect 2582 772 2583 776
rect 2587 772 2588 776
rect 2582 771 2588 772
rect 2734 776 2740 777
rect 2734 772 2735 776
rect 2739 772 2740 776
rect 2734 771 2740 772
rect 2894 776 2900 777
rect 2894 772 2895 776
rect 2899 772 2900 776
rect 2894 771 2900 772
rect 3062 776 3068 777
rect 3062 772 3063 776
rect 3067 772 3068 776
rect 3062 771 3068 772
rect 3246 776 3252 777
rect 3246 772 3247 776
rect 3251 772 3252 776
rect 3246 771 3252 772
rect 3446 776 3452 777
rect 3446 772 3447 776
rect 3451 772 3452 776
rect 3446 771 3452 772
rect 3654 776 3660 777
rect 3654 772 3655 776
rect 3659 772 3660 776
rect 3654 771 3660 772
rect 3838 776 3844 777
rect 3838 772 3839 776
rect 3843 772 3844 776
rect 3942 775 3943 779
rect 3947 775 3948 779
rect 3942 774 3948 775
rect 3838 771 3844 772
rect 374 740 380 741
rect 110 737 116 738
rect 110 733 111 737
rect 115 733 116 737
rect 374 736 375 740
rect 379 736 380 740
rect 374 735 380 736
rect 494 740 500 741
rect 494 736 495 740
rect 499 736 500 740
rect 494 735 500 736
rect 622 740 628 741
rect 622 736 623 740
rect 627 736 628 740
rect 622 735 628 736
rect 750 740 756 741
rect 750 736 751 740
rect 755 736 756 740
rect 750 735 756 736
rect 886 740 892 741
rect 886 736 887 740
rect 891 736 892 740
rect 886 735 892 736
rect 1022 740 1028 741
rect 1022 736 1023 740
rect 1027 736 1028 740
rect 1022 735 1028 736
rect 1166 740 1172 741
rect 1166 736 1167 740
rect 1171 736 1172 740
rect 1166 735 1172 736
rect 1310 740 1316 741
rect 1310 736 1311 740
rect 1315 736 1316 740
rect 1310 735 1316 736
rect 1454 740 1460 741
rect 1454 736 1455 740
rect 1459 736 1460 740
rect 1454 735 1460 736
rect 1598 740 1604 741
rect 1598 736 1599 740
rect 1603 736 1604 740
rect 1598 735 1604 736
rect 2006 737 2012 738
rect 110 732 116 733
rect 2006 733 2007 737
rect 2011 733 2012 737
rect 2006 732 2012 733
rect 374 721 380 722
rect 110 720 116 721
rect 110 716 111 720
rect 115 716 116 720
rect 374 717 375 721
rect 379 717 380 721
rect 374 716 380 717
rect 494 721 500 722
rect 494 717 495 721
rect 499 717 500 721
rect 494 716 500 717
rect 622 721 628 722
rect 622 717 623 721
rect 627 717 628 721
rect 622 716 628 717
rect 750 721 756 722
rect 750 717 751 721
rect 755 717 756 721
rect 750 716 756 717
rect 886 721 892 722
rect 886 717 887 721
rect 891 717 892 721
rect 886 716 892 717
rect 1022 721 1028 722
rect 1022 717 1023 721
rect 1027 717 1028 721
rect 1022 716 1028 717
rect 1166 721 1172 722
rect 1166 717 1167 721
rect 1171 717 1172 721
rect 1166 716 1172 717
rect 1310 721 1316 722
rect 1310 717 1311 721
rect 1315 717 1316 721
rect 1310 716 1316 717
rect 1454 721 1460 722
rect 1454 717 1455 721
rect 1459 717 1460 721
rect 1454 716 1460 717
rect 1598 721 1604 722
rect 1598 717 1599 721
rect 1603 717 1604 721
rect 1598 716 1604 717
rect 2006 720 2012 721
rect 2006 716 2007 720
rect 2011 716 2012 720
rect 110 715 116 716
rect 2006 715 2012 716
rect 2374 712 2380 713
rect 2046 709 2052 710
rect 2046 705 2047 709
rect 2051 705 2052 709
rect 2374 708 2375 712
rect 2379 708 2380 712
rect 2374 707 2380 708
rect 2494 712 2500 713
rect 2494 708 2495 712
rect 2499 708 2500 712
rect 2494 707 2500 708
rect 2622 712 2628 713
rect 2622 708 2623 712
rect 2627 708 2628 712
rect 2622 707 2628 708
rect 2766 712 2772 713
rect 2766 708 2767 712
rect 2771 708 2772 712
rect 2766 707 2772 708
rect 2910 712 2916 713
rect 2910 708 2911 712
rect 2915 708 2916 712
rect 2910 707 2916 708
rect 3062 712 3068 713
rect 3062 708 3063 712
rect 3067 708 3068 712
rect 3062 707 3068 708
rect 3214 712 3220 713
rect 3214 708 3215 712
rect 3219 708 3220 712
rect 3214 707 3220 708
rect 3366 712 3372 713
rect 3366 708 3367 712
rect 3371 708 3372 712
rect 3366 707 3372 708
rect 3518 712 3524 713
rect 3518 708 3519 712
rect 3523 708 3524 712
rect 3518 707 3524 708
rect 3678 712 3684 713
rect 3678 708 3679 712
rect 3683 708 3684 712
rect 3678 707 3684 708
rect 3838 712 3844 713
rect 3838 708 3839 712
rect 3843 708 3844 712
rect 3838 707 3844 708
rect 3942 709 3948 710
rect 2046 704 2052 705
rect 3942 705 3943 709
rect 3947 705 3948 709
rect 3942 704 3948 705
rect 2374 693 2380 694
rect 2046 692 2052 693
rect 2046 688 2047 692
rect 2051 688 2052 692
rect 2374 689 2375 693
rect 2379 689 2380 693
rect 2374 688 2380 689
rect 2494 693 2500 694
rect 2494 689 2495 693
rect 2499 689 2500 693
rect 2494 688 2500 689
rect 2622 693 2628 694
rect 2622 689 2623 693
rect 2627 689 2628 693
rect 2622 688 2628 689
rect 2766 693 2772 694
rect 2766 689 2767 693
rect 2771 689 2772 693
rect 2766 688 2772 689
rect 2910 693 2916 694
rect 2910 689 2911 693
rect 2915 689 2916 693
rect 2910 688 2916 689
rect 3062 693 3068 694
rect 3062 689 3063 693
rect 3067 689 3068 693
rect 3062 688 3068 689
rect 3214 693 3220 694
rect 3214 689 3215 693
rect 3219 689 3220 693
rect 3214 688 3220 689
rect 3366 693 3372 694
rect 3366 689 3367 693
rect 3371 689 3372 693
rect 3366 688 3372 689
rect 3518 693 3524 694
rect 3518 689 3519 693
rect 3523 689 3524 693
rect 3518 688 3524 689
rect 3678 693 3684 694
rect 3678 689 3679 693
rect 3683 689 3684 693
rect 3678 688 3684 689
rect 3838 693 3844 694
rect 3838 689 3839 693
rect 3843 689 3844 693
rect 3838 688 3844 689
rect 3942 692 3948 693
rect 3942 688 3943 692
rect 3947 688 3948 692
rect 2046 687 2052 688
rect 3942 687 3948 688
rect 110 668 116 669
rect 2006 668 2012 669
rect 110 664 111 668
rect 115 664 116 668
rect 110 663 116 664
rect 526 667 532 668
rect 526 663 527 667
rect 531 663 532 667
rect 526 662 532 663
rect 630 667 636 668
rect 630 663 631 667
rect 635 663 636 667
rect 630 662 636 663
rect 742 667 748 668
rect 742 663 743 667
rect 747 663 748 667
rect 742 662 748 663
rect 854 667 860 668
rect 854 663 855 667
rect 859 663 860 667
rect 854 662 860 663
rect 966 667 972 668
rect 966 663 967 667
rect 971 663 972 667
rect 966 662 972 663
rect 1070 667 1076 668
rect 1070 663 1071 667
rect 1075 663 1076 667
rect 1070 662 1076 663
rect 1182 667 1188 668
rect 1182 663 1183 667
rect 1187 663 1188 667
rect 1182 662 1188 663
rect 1294 667 1300 668
rect 1294 663 1295 667
rect 1299 663 1300 667
rect 1294 662 1300 663
rect 1406 667 1412 668
rect 1406 663 1407 667
rect 1411 663 1412 667
rect 1406 662 1412 663
rect 1518 667 1524 668
rect 1518 663 1519 667
rect 1523 663 1524 667
rect 2006 664 2007 668
rect 2011 664 2012 668
rect 2006 663 2012 664
rect 1518 662 1524 663
rect 110 651 116 652
rect 110 647 111 651
rect 115 647 116 651
rect 2006 651 2012 652
rect 110 646 116 647
rect 526 648 532 649
rect 526 644 527 648
rect 531 644 532 648
rect 526 643 532 644
rect 630 648 636 649
rect 630 644 631 648
rect 635 644 636 648
rect 630 643 636 644
rect 742 648 748 649
rect 742 644 743 648
rect 747 644 748 648
rect 742 643 748 644
rect 854 648 860 649
rect 854 644 855 648
rect 859 644 860 648
rect 854 643 860 644
rect 966 648 972 649
rect 966 644 967 648
rect 971 644 972 648
rect 966 643 972 644
rect 1070 648 1076 649
rect 1070 644 1071 648
rect 1075 644 1076 648
rect 1070 643 1076 644
rect 1182 648 1188 649
rect 1182 644 1183 648
rect 1187 644 1188 648
rect 1182 643 1188 644
rect 1294 648 1300 649
rect 1294 644 1295 648
rect 1299 644 1300 648
rect 1294 643 1300 644
rect 1406 648 1412 649
rect 1406 644 1407 648
rect 1411 644 1412 648
rect 1406 643 1412 644
rect 1518 648 1524 649
rect 1518 644 1519 648
rect 1523 644 1524 648
rect 2006 647 2007 651
rect 2011 647 2012 651
rect 2006 646 2012 647
rect 1518 643 1524 644
rect 2046 632 2052 633
rect 3942 632 3948 633
rect 2046 628 2047 632
rect 2051 628 2052 632
rect 2046 627 2052 628
rect 2110 631 2116 632
rect 2110 627 2111 631
rect 2115 627 2116 631
rect 2110 626 2116 627
rect 2246 631 2252 632
rect 2246 627 2247 631
rect 2251 627 2252 631
rect 2246 626 2252 627
rect 2398 631 2404 632
rect 2398 627 2399 631
rect 2403 627 2404 631
rect 2398 626 2404 627
rect 2574 631 2580 632
rect 2574 627 2575 631
rect 2579 627 2580 631
rect 2574 626 2580 627
rect 2758 631 2764 632
rect 2758 627 2759 631
rect 2763 627 2764 631
rect 2758 626 2764 627
rect 2942 631 2948 632
rect 2942 627 2943 631
rect 2947 627 2948 631
rect 2942 626 2948 627
rect 3126 631 3132 632
rect 3126 627 3127 631
rect 3131 627 3132 631
rect 3126 626 3132 627
rect 3302 631 3308 632
rect 3302 627 3303 631
rect 3307 627 3308 631
rect 3302 626 3308 627
rect 3478 631 3484 632
rect 3478 627 3479 631
rect 3483 627 3484 631
rect 3478 626 3484 627
rect 3654 631 3660 632
rect 3654 627 3655 631
rect 3659 627 3660 631
rect 3654 626 3660 627
rect 3830 631 3836 632
rect 3830 627 3831 631
rect 3835 627 3836 631
rect 3942 628 3943 632
rect 3947 628 3948 632
rect 3942 627 3948 628
rect 3830 626 3836 627
rect 2046 615 2052 616
rect 2046 611 2047 615
rect 2051 611 2052 615
rect 3942 615 3948 616
rect 2046 610 2052 611
rect 2110 612 2116 613
rect 2110 608 2111 612
rect 2115 608 2116 612
rect 2110 607 2116 608
rect 2246 612 2252 613
rect 2246 608 2247 612
rect 2251 608 2252 612
rect 2246 607 2252 608
rect 2398 612 2404 613
rect 2398 608 2399 612
rect 2403 608 2404 612
rect 2398 607 2404 608
rect 2574 612 2580 613
rect 2574 608 2575 612
rect 2579 608 2580 612
rect 2574 607 2580 608
rect 2758 612 2764 613
rect 2758 608 2759 612
rect 2763 608 2764 612
rect 2758 607 2764 608
rect 2942 612 2948 613
rect 2942 608 2943 612
rect 2947 608 2948 612
rect 2942 607 2948 608
rect 3126 612 3132 613
rect 3126 608 3127 612
rect 3131 608 3132 612
rect 3126 607 3132 608
rect 3302 612 3308 613
rect 3302 608 3303 612
rect 3307 608 3308 612
rect 3302 607 3308 608
rect 3478 612 3484 613
rect 3478 608 3479 612
rect 3483 608 3484 612
rect 3478 607 3484 608
rect 3654 612 3660 613
rect 3654 608 3655 612
rect 3659 608 3660 612
rect 3654 607 3660 608
rect 3830 612 3836 613
rect 3830 608 3831 612
rect 3835 608 3836 612
rect 3942 611 3943 615
rect 3947 611 3948 615
rect 3942 610 3948 611
rect 3830 607 3836 608
rect 686 588 692 589
rect 110 585 116 586
rect 110 581 111 585
rect 115 581 116 585
rect 686 584 687 588
rect 691 584 692 588
rect 686 583 692 584
rect 782 588 788 589
rect 782 584 783 588
rect 787 584 788 588
rect 782 583 788 584
rect 878 588 884 589
rect 878 584 879 588
rect 883 584 884 588
rect 878 583 884 584
rect 974 588 980 589
rect 974 584 975 588
rect 979 584 980 588
rect 974 583 980 584
rect 1070 588 1076 589
rect 1070 584 1071 588
rect 1075 584 1076 588
rect 1070 583 1076 584
rect 1166 588 1172 589
rect 1166 584 1167 588
rect 1171 584 1172 588
rect 1166 583 1172 584
rect 1262 588 1268 589
rect 1262 584 1263 588
rect 1267 584 1268 588
rect 1262 583 1268 584
rect 1358 588 1364 589
rect 1358 584 1359 588
rect 1363 584 1364 588
rect 1358 583 1364 584
rect 1454 588 1460 589
rect 1454 584 1455 588
rect 1459 584 1460 588
rect 1454 583 1460 584
rect 2006 585 2012 586
rect 110 580 116 581
rect 2006 581 2007 585
rect 2011 581 2012 585
rect 2006 580 2012 581
rect 686 569 692 570
rect 110 568 116 569
rect 110 564 111 568
rect 115 564 116 568
rect 686 565 687 569
rect 691 565 692 569
rect 686 564 692 565
rect 782 569 788 570
rect 782 565 783 569
rect 787 565 788 569
rect 782 564 788 565
rect 878 569 884 570
rect 878 565 879 569
rect 883 565 884 569
rect 878 564 884 565
rect 974 569 980 570
rect 974 565 975 569
rect 979 565 980 569
rect 974 564 980 565
rect 1070 569 1076 570
rect 1070 565 1071 569
rect 1075 565 1076 569
rect 1070 564 1076 565
rect 1166 569 1172 570
rect 1166 565 1167 569
rect 1171 565 1172 569
rect 1166 564 1172 565
rect 1262 569 1268 570
rect 1262 565 1263 569
rect 1267 565 1268 569
rect 1262 564 1268 565
rect 1358 569 1364 570
rect 1358 565 1359 569
rect 1363 565 1364 569
rect 1358 564 1364 565
rect 1454 569 1460 570
rect 1454 565 1455 569
rect 1459 565 1460 569
rect 1454 564 1460 565
rect 2006 568 2012 569
rect 2006 564 2007 568
rect 2011 564 2012 568
rect 110 563 116 564
rect 2006 563 2012 564
rect 2070 548 2076 549
rect 2046 545 2052 546
rect 2046 541 2047 545
rect 2051 541 2052 545
rect 2070 544 2071 548
rect 2075 544 2076 548
rect 2070 543 2076 544
rect 2182 548 2188 549
rect 2182 544 2183 548
rect 2187 544 2188 548
rect 2182 543 2188 544
rect 2334 548 2340 549
rect 2334 544 2335 548
rect 2339 544 2340 548
rect 2334 543 2340 544
rect 2502 548 2508 549
rect 2502 544 2503 548
rect 2507 544 2508 548
rect 2502 543 2508 544
rect 2686 548 2692 549
rect 2686 544 2687 548
rect 2691 544 2692 548
rect 2686 543 2692 544
rect 2878 548 2884 549
rect 2878 544 2879 548
rect 2883 544 2884 548
rect 2878 543 2884 544
rect 3070 548 3076 549
rect 3070 544 3071 548
rect 3075 544 3076 548
rect 3070 543 3076 544
rect 3262 548 3268 549
rect 3262 544 3263 548
rect 3267 544 3268 548
rect 3262 543 3268 544
rect 3454 548 3460 549
rect 3454 544 3455 548
rect 3459 544 3460 548
rect 3454 543 3460 544
rect 3646 548 3652 549
rect 3646 544 3647 548
rect 3651 544 3652 548
rect 3646 543 3652 544
rect 3838 548 3844 549
rect 3838 544 3839 548
rect 3843 544 3844 548
rect 3838 543 3844 544
rect 3942 545 3948 546
rect 2046 540 2052 541
rect 3942 541 3943 545
rect 3947 541 3948 545
rect 3942 540 3948 541
rect 2070 529 2076 530
rect 2046 528 2052 529
rect 2046 524 2047 528
rect 2051 524 2052 528
rect 2070 525 2071 529
rect 2075 525 2076 529
rect 2070 524 2076 525
rect 2182 529 2188 530
rect 2182 525 2183 529
rect 2187 525 2188 529
rect 2182 524 2188 525
rect 2334 529 2340 530
rect 2334 525 2335 529
rect 2339 525 2340 529
rect 2334 524 2340 525
rect 2502 529 2508 530
rect 2502 525 2503 529
rect 2507 525 2508 529
rect 2502 524 2508 525
rect 2686 529 2692 530
rect 2686 525 2687 529
rect 2691 525 2692 529
rect 2686 524 2692 525
rect 2878 529 2884 530
rect 2878 525 2879 529
rect 2883 525 2884 529
rect 2878 524 2884 525
rect 3070 529 3076 530
rect 3070 525 3071 529
rect 3075 525 3076 529
rect 3070 524 3076 525
rect 3262 529 3268 530
rect 3262 525 3263 529
rect 3267 525 3268 529
rect 3262 524 3268 525
rect 3454 529 3460 530
rect 3454 525 3455 529
rect 3459 525 3460 529
rect 3454 524 3460 525
rect 3646 529 3652 530
rect 3646 525 3647 529
rect 3651 525 3652 529
rect 3646 524 3652 525
rect 3838 529 3844 530
rect 3838 525 3839 529
rect 3843 525 3844 529
rect 3838 524 3844 525
rect 3942 528 3948 529
rect 3942 524 3943 528
rect 3947 524 3948 528
rect 2046 523 2052 524
rect 3942 523 3948 524
rect 110 496 116 497
rect 2006 496 2012 497
rect 110 492 111 496
rect 115 492 116 496
rect 110 491 116 492
rect 382 495 388 496
rect 382 491 383 495
rect 387 491 388 495
rect 382 490 388 491
rect 478 495 484 496
rect 478 491 479 495
rect 483 491 484 495
rect 478 490 484 491
rect 574 495 580 496
rect 574 491 575 495
rect 579 491 580 495
rect 574 490 580 491
rect 670 495 676 496
rect 670 491 671 495
rect 675 491 676 495
rect 670 490 676 491
rect 766 495 772 496
rect 766 491 767 495
rect 771 491 772 495
rect 766 490 772 491
rect 862 495 868 496
rect 862 491 863 495
rect 867 491 868 495
rect 862 490 868 491
rect 958 495 964 496
rect 958 491 959 495
rect 963 491 964 495
rect 958 490 964 491
rect 1054 495 1060 496
rect 1054 491 1055 495
rect 1059 491 1060 495
rect 1054 490 1060 491
rect 1150 495 1156 496
rect 1150 491 1151 495
rect 1155 491 1156 495
rect 1150 490 1156 491
rect 1246 495 1252 496
rect 1246 491 1247 495
rect 1251 491 1252 495
rect 1246 490 1252 491
rect 1342 495 1348 496
rect 1342 491 1343 495
rect 1347 491 1348 495
rect 1342 490 1348 491
rect 1438 495 1444 496
rect 1438 491 1439 495
rect 1443 491 1444 495
rect 1438 490 1444 491
rect 1534 495 1540 496
rect 1534 491 1535 495
rect 1539 491 1540 495
rect 2006 492 2007 496
rect 2011 492 2012 496
rect 2006 491 2012 492
rect 1534 490 1540 491
rect 110 479 116 480
rect 110 475 111 479
rect 115 475 116 479
rect 2006 479 2012 480
rect 110 474 116 475
rect 382 476 388 477
rect 382 472 383 476
rect 387 472 388 476
rect 382 471 388 472
rect 478 476 484 477
rect 478 472 479 476
rect 483 472 484 476
rect 478 471 484 472
rect 574 476 580 477
rect 574 472 575 476
rect 579 472 580 476
rect 574 471 580 472
rect 670 476 676 477
rect 670 472 671 476
rect 675 472 676 476
rect 670 471 676 472
rect 766 476 772 477
rect 766 472 767 476
rect 771 472 772 476
rect 766 471 772 472
rect 862 476 868 477
rect 862 472 863 476
rect 867 472 868 476
rect 862 471 868 472
rect 958 476 964 477
rect 958 472 959 476
rect 963 472 964 476
rect 958 471 964 472
rect 1054 476 1060 477
rect 1054 472 1055 476
rect 1059 472 1060 476
rect 1054 471 1060 472
rect 1150 476 1156 477
rect 1150 472 1151 476
rect 1155 472 1156 476
rect 1150 471 1156 472
rect 1246 476 1252 477
rect 1246 472 1247 476
rect 1251 472 1252 476
rect 1246 471 1252 472
rect 1342 476 1348 477
rect 1342 472 1343 476
rect 1347 472 1348 476
rect 1342 471 1348 472
rect 1438 476 1444 477
rect 1438 472 1439 476
rect 1443 472 1444 476
rect 1438 471 1444 472
rect 1534 476 1540 477
rect 1534 472 1535 476
rect 1539 472 1540 476
rect 2006 475 2007 479
rect 2011 475 2012 479
rect 2006 474 2012 475
rect 2046 476 2052 477
rect 3942 476 3948 477
rect 1534 471 1540 472
rect 2046 472 2047 476
rect 2051 472 2052 476
rect 2046 471 2052 472
rect 2182 475 2188 476
rect 2182 471 2183 475
rect 2187 471 2188 475
rect 2182 470 2188 471
rect 2318 475 2324 476
rect 2318 471 2319 475
rect 2323 471 2324 475
rect 2318 470 2324 471
rect 2462 475 2468 476
rect 2462 471 2463 475
rect 2467 471 2468 475
rect 2462 470 2468 471
rect 2614 475 2620 476
rect 2614 471 2615 475
rect 2619 471 2620 475
rect 2614 470 2620 471
rect 2774 475 2780 476
rect 2774 471 2775 475
rect 2779 471 2780 475
rect 2774 470 2780 471
rect 2958 475 2964 476
rect 2958 471 2959 475
rect 2963 471 2964 475
rect 2958 470 2964 471
rect 3158 475 3164 476
rect 3158 471 3159 475
rect 3163 471 3164 475
rect 3158 470 3164 471
rect 3366 475 3372 476
rect 3366 471 3367 475
rect 3371 471 3372 475
rect 3366 470 3372 471
rect 3582 475 3588 476
rect 3582 471 3583 475
rect 3587 471 3588 475
rect 3582 470 3588 471
rect 3806 475 3812 476
rect 3806 471 3807 475
rect 3811 471 3812 475
rect 3942 472 3943 476
rect 3947 472 3948 476
rect 3942 471 3948 472
rect 3806 470 3812 471
rect 2046 459 2052 460
rect 2046 455 2047 459
rect 2051 455 2052 459
rect 3942 459 3948 460
rect 2046 454 2052 455
rect 2182 456 2188 457
rect 2182 452 2183 456
rect 2187 452 2188 456
rect 2182 451 2188 452
rect 2318 456 2324 457
rect 2318 452 2319 456
rect 2323 452 2324 456
rect 2318 451 2324 452
rect 2462 456 2468 457
rect 2462 452 2463 456
rect 2467 452 2468 456
rect 2462 451 2468 452
rect 2614 456 2620 457
rect 2614 452 2615 456
rect 2619 452 2620 456
rect 2614 451 2620 452
rect 2774 456 2780 457
rect 2774 452 2775 456
rect 2779 452 2780 456
rect 2774 451 2780 452
rect 2958 456 2964 457
rect 2958 452 2959 456
rect 2963 452 2964 456
rect 2958 451 2964 452
rect 3158 456 3164 457
rect 3158 452 3159 456
rect 3163 452 3164 456
rect 3158 451 3164 452
rect 3366 456 3372 457
rect 3366 452 3367 456
rect 3371 452 3372 456
rect 3366 451 3372 452
rect 3582 456 3588 457
rect 3582 452 3583 456
rect 3587 452 3588 456
rect 3582 451 3588 452
rect 3806 456 3812 457
rect 3806 452 3807 456
rect 3811 452 3812 456
rect 3942 455 3943 459
rect 3947 455 3948 459
rect 3942 454 3948 455
rect 3806 451 3812 452
rect 486 404 492 405
rect 110 401 116 402
rect 110 397 111 401
rect 115 397 116 401
rect 486 400 487 404
rect 491 400 492 404
rect 486 399 492 400
rect 582 404 588 405
rect 582 400 583 404
rect 587 400 588 404
rect 582 399 588 400
rect 686 404 692 405
rect 686 400 687 404
rect 691 400 692 404
rect 686 399 692 400
rect 790 404 796 405
rect 790 400 791 404
rect 795 400 796 404
rect 790 399 796 400
rect 894 404 900 405
rect 894 400 895 404
rect 899 400 900 404
rect 894 399 900 400
rect 998 404 1004 405
rect 998 400 999 404
rect 1003 400 1004 404
rect 998 399 1004 400
rect 1102 404 1108 405
rect 1102 400 1103 404
rect 1107 400 1108 404
rect 1102 399 1108 400
rect 1206 404 1212 405
rect 1206 400 1207 404
rect 1211 400 1212 404
rect 1206 399 1212 400
rect 1318 404 1324 405
rect 1318 400 1319 404
rect 1323 400 1324 404
rect 1318 399 1324 400
rect 1430 404 1436 405
rect 1430 400 1431 404
rect 1435 400 1436 404
rect 1430 399 1436 400
rect 2006 401 2012 402
rect 110 396 116 397
rect 2006 397 2007 401
rect 2011 397 2012 401
rect 2006 396 2012 397
rect 2342 396 2348 397
rect 2046 393 2052 394
rect 2046 389 2047 393
rect 2051 389 2052 393
rect 2342 392 2343 396
rect 2347 392 2348 396
rect 2342 391 2348 392
rect 2486 396 2492 397
rect 2486 392 2487 396
rect 2491 392 2492 396
rect 2486 391 2492 392
rect 2638 396 2644 397
rect 2638 392 2639 396
rect 2643 392 2644 396
rect 2638 391 2644 392
rect 2798 396 2804 397
rect 2798 392 2799 396
rect 2803 392 2804 396
rect 2798 391 2804 392
rect 2958 396 2964 397
rect 2958 392 2959 396
rect 2963 392 2964 396
rect 2958 391 2964 392
rect 3110 396 3116 397
rect 3110 392 3111 396
rect 3115 392 3116 396
rect 3110 391 3116 392
rect 3262 396 3268 397
rect 3262 392 3263 396
rect 3267 392 3268 396
rect 3262 391 3268 392
rect 3414 396 3420 397
rect 3414 392 3415 396
rect 3419 392 3420 396
rect 3414 391 3420 392
rect 3558 396 3564 397
rect 3558 392 3559 396
rect 3563 392 3564 396
rect 3558 391 3564 392
rect 3710 396 3716 397
rect 3710 392 3711 396
rect 3715 392 3716 396
rect 3710 391 3716 392
rect 3838 396 3844 397
rect 3838 392 3839 396
rect 3843 392 3844 396
rect 3838 391 3844 392
rect 3942 393 3948 394
rect 2046 388 2052 389
rect 3942 389 3943 393
rect 3947 389 3948 393
rect 3942 388 3948 389
rect 486 385 492 386
rect 110 384 116 385
rect 110 380 111 384
rect 115 380 116 384
rect 486 381 487 385
rect 491 381 492 385
rect 486 380 492 381
rect 582 385 588 386
rect 582 381 583 385
rect 587 381 588 385
rect 582 380 588 381
rect 686 385 692 386
rect 686 381 687 385
rect 691 381 692 385
rect 686 380 692 381
rect 790 385 796 386
rect 790 381 791 385
rect 795 381 796 385
rect 790 380 796 381
rect 894 385 900 386
rect 894 381 895 385
rect 899 381 900 385
rect 894 380 900 381
rect 998 385 1004 386
rect 998 381 999 385
rect 1003 381 1004 385
rect 998 380 1004 381
rect 1102 385 1108 386
rect 1102 381 1103 385
rect 1107 381 1108 385
rect 1102 380 1108 381
rect 1206 385 1212 386
rect 1206 381 1207 385
rect 1211 381 1212 385
rect 1206 380 1212 381
rect 1318 385 1324 386
rect 1318 381 1319 385
rect 1323 381 1324 385
rect 1318 380 1324 381
rect 1430 385 1436 386
rect 1430 381 1431 385
rect 1435 381 1436 385
rect 1430 380 1436 381
rect 2006 384 2012 385
rect 2006 380 2007 384
rect 2011 380 2012 384
rect 110 379 116 380
rect 2006 379 2012 380
rect 2342 377 2348 378
rect 2046 376 2052 377
rect 2046 372 2047 376
rect 2051 372 2052 376
rect 2342 373 2343 377
rect 2347 373 2348 377
rect 2342 372 2348 373
rect 2486 377 2492 378
rect 2486 373 2487 377
rect 2491 373 2492 377
rect 2486 372 2492 373
rect 2638 377 2644 378
rect 2638 373 2639 377
rect 2643 373 2644 377
rect 2638 372 2644 373
rect 2798 377 2804 378
rect 2798 373 2799 377
rect 2803 373 2804 377
rect 2798 372 2804 373
rect 2958 377 2964 378
rect 2958 373 2959 377
rect 2963 373 2964 377
rect 2958 372 2964 373
rect 3110 377 3116 378
rect 3110 373 3111 377
rect 3115 373 3116 377
rect 3110 372 3116 373
rect 3262 377 3268 378
rect 3262 373 3263 377
rect 3267 373 3268 377
rect 3262 372 3268 373
rect 3414 377 3420 378
rect 3414 373 3415 377
rect 3419 373 3420 377
rect 3414 372 3420 373
rect 3558 377 3564 378
rect 3558 373 3559 377
rect 3563 373 3564 377
rect 3558 372 3564 373
rect 3710 377 3716 378
rect 3710 373 3711 377
rect 3715 373 3716 377
rect 3710 372 3716 373
rect 3838 377 3844 378
rect 3838 373 3839 377
rect 3843 373 3844 377
rect 3838 372 3844 373
rect 3942 376 3948 377
rect 3942 372 3943 376
rect 3947 372 3948 376
rect 2046 371 2052 372
rect 3942 371 3948 372
rect 110 328 116 329
rect 2006 328 2012 329
rect 110 324 111 328
rect 115 324 116 328
rect 110 323 116 324
rect 326 327 332 328
rect 326 323 327 327
rect 331 323 332 327
rect 326 322 332 323
rect 462 327 468 328
rect 462 323 463 327
rect 467 323 468 327
rect 462 322 468 323
rect 614 327 620 328
rect 614 323 615 327
rect 619 323 620 327
rect 614 322 620 323
rect 766 327 772 328
rect 766 323 767 327
rect 771 323 772 327
rect 766 322 772 323
rect 918 327 924 328
rect 918 323 919 327
rect 923 323 924 327
rect 918 322 924 323
rect 1062 327 1068 328
rect 1062 323 1063 327
rect 1067 323 1068 327
rect 1062 322 1068 323
rect 1206 327 1212 328
rect 1206 323 1207 327
rect 1211 323 1212 327
rect 1206 322 1212 323
rect 1350 327 1356 328
rect 1350 323 1351 327
rect 1355 323 1356 327
rect 1350 322 1356 323
rect 1494 327 1500 328
rect 1494 323 1495 327
rect 1499 323 1500 327
rect 1494 322 1500 323
rect 1638 327 1644 328
rect 1638 323 1639 327
rect 1643 323 1644 327
rect 2006 324 2007 328
rect 2011 324 2012 328
rect 2006 323 2012 324
rect 1638 322 1644 323
rect 2046 320 2052 321
rect 3942 320 3948 321
rect 2046 316 2047 320
rect 2051 316 2052 320
rect 2046 315 2052 316
rect 2494 319 2500 320
rect 2494 315 2495 319
rect 2499 315 2500 319
rect 2494 314 2500 315
rect 2638 319 2644 320
rect 2638 315 2639 319
rect 2643 315 2644 319
rect 2638 314 2644 315
rect 2798 319 2804 320
rect 2798 315 2799 319
rect 2803 315 2804 319
rect 2798 314 2804 315
rect 2958 319 2964 320
rect 2958 315 2959 319
rect 2963 315 2964 319
rect 2958 314 2964 315
rect 3118 319 3124 320
rect 3118 315 3119 319
rect 3123 315 3124 319
rect 3118 314 3124 315
rect 3270 319 3276 320
rect 3270 315 3271 319
rect 3275 315 3276 319
rect 3270 314 3276 315
rect 3422 319 3428 320
rect 3422 315 3423 319
rect 3427 315 3428 319
rect 3422 314 3428 315
rect 3566 319 3572 320
rect 3566 315 3567 319
rect 3571 315 3572 319
rect 3566 314 3572 315
rect 3710 319 3716 320
rect 3710 315 3711 319
rect 3715 315 3716 319
rect 3710 314 3716 315
rect 3838 319 3844 320
rect 3838 315 3839 319
rect 3843 315 3844 319
rect 3942 316 3943 320
rect 3947 316 3948 320
rect 3942 315 3948 316
rect 3838 314 3844 315
rect 110 311 116 312
rect 110 307 111 311
rect 115 307 116 311
rect 2006 311 2012 312
rect 110 306 116 307
rect 326 308 332 309
rect 326 304 327 308
rect 331 304 332 308
rect 326 303 332 304
rect 462 308 468 309
rect 462 304 463 308
rect 467 304 468 308
rect 462 303 468 304
rect 614 308 620 309
rect 614 304 615 308
rect 619 304 620 308
rect 614 303 620 304
rect 766 308 772 309
rect 766 304 767 308
rect 771 304 772 308
rect 766 303 772 304
rect 918 308 924 309
rect 918 304 919 308
rect 923 304 924 308
rect 918 303 924 304
rect 1062 308 1068 309
rect 1062 304 1063 308
rect 1067 304 1068 308
rect 1062 303 1068 304
rect 1206 308 1212 309
rect 1206 304 1207 308
rect 1211 304 1212 308
rect 1206 303 1212 304
rect 1350 308 1356 309
rect 1350 304 1351 308
rect 1355 304 1356 308
rect 1350 303 1356 304
rect 1494 308 1500 309
rect 1494 304 1495 308
rect 1499 304 1500 308
rect 1494 303 1500 304
rect 1638 308 1644 309
rect 1638 304 1639 308
rect 1643 304 1644 308
rect 2006 307 2007 311
rect 2011 307 2012 311
rect 2006 306 2012 307
rect 1638 303 1644 304
rect 2046 303 2052 304
rect 2046 299 2047 303
rect 2051 299 2052 303
rect 3942 303 3948 304
rect 2046 298 2052 299
rect 2494 300 2500 301
rect 2494 296 2495 300
rect 2499 296 2500 300
rect 2494 295 2500 296
rect 2638 300 2644 301
rect 2638 296 2639 300
rect 2643 296 2644 300
rect 2638 295 2644 296
rect 2798 300 2804 301
rect 2798 296 2799 300
rect 2803 296 2804 300
rect 2798 295 2804 296
rect 2958 300 2964 301
rect 2958 296 2959 300
rect 2963 296 2964 300
rect 2958 295 2964 296
rect 3118 300 3124 301
rect 3118 296 3119 300
rect 3123 296 3124 300
rect 3118 295 3124 296
rect 3270 300 3276 301
rect 3270 296 3271 300
rect 3275 296 3276 300
rect 3270 295 3276 296
rect 3422 300 3428 301
rect 3422 296 3423 300
rect 3427 296 3428 300
rect 3422 295 3428 296
rect 3566 300 3572 301
rect 3566 296 3567 300
rect 3571 296 3572 300
rect 3566 295 3572 296
rect 3710 300 3716 301
rect 3710 296 3711 300
rect 3715 296 3716 300
rect 3710 295 3716 296
rect 3838 300 3844 301
rect 3838 296 3839 300
rect 3843 296 3844 300
rect 3942 299 3943 303
rect 3947 299 3948 303
rect 3942 298 3948 299
rect 3838 295 3844 296
rect 166 240 172 241
rect 110 237 116 238
rect 110 233 111 237
rect 115 233 116 237
rect 166 236 167 240
rect 171 236 172 240
rect 166 235 172 236
rect 326 240 332 241
rect 326 236 327 240
rect 331 236 332 240
rect 326 235 332 236
rect 502 240 508 241
rect 502 236 503 240
rect 507 236 508 240
rect 502 235 508 236
rect 686 240 692 241
rect 686 236 687 240
rect 691 236 692 240
rect 686 235 692 236
rect 870 240 876 241
rect 870 236 871 240
rect 875 236 876 240
rect 870 235 876 236
rect 1046 240 1052 241
rect 1046 236 1047 240
rect 1051 236 1052 240
rect 1046 235 1052 236
rect 1214 240 1220 241
rect 1214 236 1215 240
rect 1219 236 1220 240
rect 1214 235 1220 236
rect 1366 240 1372 241
rect 1366 236 1367 240
rect 1371 236 1372 240
rect 1366 235 1372 236
rect 1510 240 1516 241
rect 1510 236 1511 240
rect 1515 236 1516 240
rect 1510 235 1516 236
rect 1646 240 1652 241
rect 1646 236 1647 240
rect 1651 236 1652 240
rect 1646 235 1652 236
rect 1782 240 1788 241
rect 1782 236 1783 240
rect 1787 236 1788 240
rect 1782 235 1788 236
rect 1902 240 1908 241
rect 1902 236 1903 240
rect 1907 236 1908 240
rect 2070 240 2076 241
rect 1902 235 1908 236
rect 2006 237 2012 238
rect 110 232 116 233
rect 2006 233 2007 237
rect 2011 233 2012 237
rect 2006 232 2012 233
rect 2046 237 2052 238
rect 2046 233 2047 237
rect 2051 233 2052 237
rect 2070 236 2071 240
rect 2075 236 2076 240
rect 2070 235 2076 236
rect 2270 240 2276 241
rect 2270 236 2271 240
rect 2275 236 2276 240
rect 2270 235 2276 236
rect 2494 240 2500 241
rect 2494 236 2495 240
rect 2499 236 2500 240
rect 2494 235 2500 236
rect 2702 240 2708 241
rect 2702 236 2703 240
rect 2707 236 2708 240
rect 2702 235 2708 236
rect 2902 240 2908 241
rect 2902 236 2903 240
rect 2907 236 2908 240
rect 2902 235 2908 236
rect 3094 240 3100 241
rect 3094 236 3095 240
rect 3099 236 3100 240
rect 3094 235 3100 236
rect 3286 240 3292 241
rect 3286 236 3287 240
rect 3291 236 3292 240
rect 3286 235 3292 236
rect 3478 240 3484 241
rect 3478 236 3479 240
rect 3483 236 3484 240
rect 3478 235 3484 236
rect 3670 240 3676 241
rect 3670 236 3671 240
rect 3675 236 3676 240
rect 3670 235 3676 236
rect 3838 240 3844 241
rect 3838 236 3839 240
rect 3843 236 3844 240
rect 3838 235 3844 236
rect 3942 237 3948 238
rect 2046 232 2052 233
rect 3942 233 3943 237
rect 3947 233 3948 237
rect 3942 232 3948 233
rect 166 221 172 222
rect 110 220 116 221
rect 110 216 111 220
rect 115 216 116 220
rect 166 217 167 221
rect 171 217 172 221
rect 166 216 172 217
rect 326 221 332 222
rect 326 217 327 221
rect 331 217 332 221
rect 326 216 332 217
rect 502 221 508 222
rect 502 217 503 221
rect 507 217 508 221
rect 502 216 508 217
rect 686 221 692 222
rect 686 217 687 221
rect 691 217 692 221
rect 686 216 692 217
rect 870 221 876 222
rect 870 217 871 221
rect 875 217 876 221
rect 870 216 876 217
rect 1046 221 1052 222
rect 1046 217 1047 221
rect 1051 217 1052 221
rect 1046 216 1052 217
rect 1214 221 1220 222
rect 1214 217 1215 221
rect 1219 217 1220 221
rect 1214 216 1220 217
rect 1366 221 1372 222
rect 1366 217 1367 221
rect 1371 217 1372 221
rect 1366 216 1372 217
rect 1510 221 1516 222
rect 1510 217 1511 221
rect 1515 217 1516 221
rect 1510 216 1516 217
rect 1646 221 1652 222
rect 1646 217 1647 221
rect 1651 217 1652 221
rect 1646 216 1652 217
rect 1782 221 1788 222
rect 1782 217 1783 221
rect 1787 217 1788 221
rect 1782 216 1788 217
rect 1902 221 1908 222
rect 2070 221 2076 222
rect 1902 217 1903 221
rect 1907 217 1908 221
rect 1902 216 1908 217
rect 2006 220 2012 221
rect 2006 216 2007 220
rect 2011 216 2012 220
rect 110 215 116 216
rect 2006 215 2012 216
rect 2046 220 2052 221
rect 2046 216 2047 220
rect 2051 216 2052 220
rect 2070 217 2071 221
rect 2075 217 2076 221
rect 2070 216 2076 217
rect 2270 221 2276 222
rect 2270 217 2271 221
rect 2275 217 2276 221
rect 2270 216 2276 217
rect 2494 221 2500 222
rect 2494 217 2495 221
rect 2499 217 2500 221
rect 2494 216 2500 217
rect 2702 221 2708 222
rect 2702 217 2703 221
rect 2707 217 2708 221
rect 2702 216 2708 217
rect 2902 221 2908 222
rect 2902 217 2903 221
rect 2907 217 2908 221
rect 2902 216 2908 217
rect 3094 221 3100 222
rect 3094 217 3095 221
rect 3099 217 3100 221
rect 3094 216 3100 217
rect 3286 221 3292 222
rect 3286 217 3287 221
rect 3291 217 3292 221
rect 3286 216 3292 217
rect 3478 221 3484 222
rect 3478 217 3479 221
rect 3483 217 3484 221
rect 3478 216 3484 217
rect 3670 221 3676 222
rect 3670 217 3671 221
rect 3675 217 3676 221
rect 3670 216 3676 217
rect 3838 221 3844 222
rect 3838 217 3839 221
rect 3843 217 3844 221
rect 3838 216 3844 217
rect 3942 220 3948 221
rect 3942 216 3943 220
rect 3947 216 3948 220
rect 2046 215 2052 216
rect 3942 215 3948 216
rect 2046 144 2052 145
rect 3942 144 3948 145
rect 110 140 116 141
rect 2006 140 2012 141
rect 110 136 111 140
rect 115 136 116 140
rect 110 135 116 136
rect 134 139 140 140
rect 134 135 135 139
rect 139 135 140 139
rect 134 134 140 135
rect 230 139 236 140
rect 230 135 231 139
rect 235 135 236 139
rect 230 134 236 135
rect 326 139 332 140
rect 326 135 327 139
rect 331 135 332 139
rect 326 134 332 135
rect 422 139 428 140
rect 422 135 423 139
rect 427 135 428 139
rect 422 134 428 135
rect 526 139 532 140
rect 526 135 527 139
rect 531 135 532 139
rect 526 134 532 135
rect 646 139 652 140
rect 646 135 647 139
rect 651 135 652 139
rect 646 134 652 135
rect 774 139 780 140
rect 774 135 775 139
rect 779 135 780 139
rect 774 134 780 135
rect 902 139 908 140
rect 902 135 903 139
rect 907 135 908 139
rect 902 134 908 135
rect 1030 139 1036 140
rect 1030 135 1031 139
rect 1035 135 1036 139
rect 1030 134 1036 135
rect 1150 139 1156 140
rect 1150 135 1151 139
rect 1155 135 1156 139
rect 1150 134 1156 135
rect 1270 139 1276 140
rect 1270 135 1271 139
rect 1275 135 1276 139
rect 1270 134 1276 135
rect 1382 139 1388 140
rect 1382 135 1383 139
rect 1387 135 1388 139
rect 1382 134 1388 135
rect 1486 139 1492 140
rect 1486 135 1487 139
rect 1491 135 1492 139
rect 1486 134 1492 135
rect 1590 139 1596 140
rect 1590 135 1591 139
rect 1595 135 1596 139
rect 1590 134 1596 135
rect 1702 139 1708 140
rect 1702 135 1703 139
rect 1707 135 1708 139
rect 1702 134 1708 135
rect 1806 139 1812 140
rect 1806 135 1807 139
rect 1811 135 1812 139
rect 1806 134 1812 135
rect 1902 139 1908 140
rect 1902 135 1903 139
rect 1907 135 1908 139
rect 2006 136 2007 140
rect 2011 136 2012 140
rect 2046 140 2047 144
rect 2051 140 2052 144
rect 2046 139 2052 140
rect 2070 143 2076 144
rect 2070 139 2071 143
rect 2075 139 2076 143
rect 2070 138 2076 139
rect 2166 143 2172 144
rect 2166 139 2167 143
rect 2171 139 2172 143
rect 2166 138 2172 139
rect 2262 143 2268 144
rect 2262 139 2263 143
rect 2267 139 2268 143
rect 2262 138 2268 139
rect 2358 143 2364 144
rect 2358 139 2359 143
rect 2363 139 2364 143
rect 2358 138 2364 139
rect 2454 143 2460 144
rect 2454 139 2455 143
rect 2459 139 2460 143
rect 2454 138 2460 139
rect 2550 143 2556 144
rect 2550 139 2551 143
rect 2555 139 2556 143
rect 2550 138 2556 139
rect 2654 143 2660 144
rect 2654 139 2655 143
rect 2659 139 2660 143
rect 2654 138 2660 139
rect 2758 143 2764 144
rect 2758 139 2759 143
rect 2763 139 2764 143
rect 2758 138 2764 139
rect 2862 143 2868 144
rect 2862 139 2863 143
rect 2867 139 2868 143
rect 2862 138 2868 139
rect 2974 143 2980 144
rect 2974 139 2975 143
rect 2979 139 2980 143
rect 2974 138 2980 139
rect 3102 143 3108 144
rect 3102 139 3103 143
rect 3107 139 3108 143
rect 3102 138 3108 139
rect 3238 143 3244 144
rect 3238 139 3239 143
rect 3243 139 3244 143
rect 3238 138 3244 139
rect 3382 143 3388 144
rect 3382 139 3383 143
rect 3387 139 3388 143
rect 3382 138 3388 139
rect 3534 143 3540 144
rect 3534 139 3535 143
rect 3539 139 3540 143
rect 3534 138 3540 139
rect 3694 143 3700 144
rect 3694 139 3695 143
rect 3699 139 3700 143
rect 3694 138 3700 139
rect 3838 143 3844 144
rect 3838 139 3839 143
rect 3843 139 3844 143
rect 3942 140 3943 144
rect 3947 140 3948 144
rect 3942 139 3948 140
rect 3838 138 3844 139
rect 2006 135 2012 136
rect 1902 134 1908 135
rect 2046 127 2052 128
rect 110 123 116 124
rect 110 119 111 123
rect 115 119 116 123
rect 2006 123 2012 124
rect 110 118 116 119
rect 134 120 140 121
rect 134 116 135 120
rect 139 116 140 120
rect 134 115 140 116
rect 230 120 236 121
rect 230 116 231 120
rect 235 116 236 120
rect 230 115 236 116
rect 326 120 332 121
rect 326 116 327 120
rect 331 116 332 120
rect 326 115 332 116
rect 422 120 428 121
rect 422 116 423 120
rect 427 116 428 120
rect 422 115 428 116
rect 526 120 532 121
rect 526 116 527 120
rect 531 116 532 120
rect 526 115 532 116
rect 646 120 652 121
rect 646 116 647 120
rect 651 116 652 120
rect 646 115 652 116
rect 774 120 780 121
rect 774 116 775 120
rect 779 116 780 120
rect 774 115 780 116
rect 902 120 908 121
rect 902 116 903 120
rect 907 116 908 120
rect 902 115 908 116
rect 1030 120 1036 121
rect 1030 116 1031 120
rect 1035 116 1036 120
rect 1030 115 1036 116
rect 1150 120 1156 121
rect 1150 116 1151 120
rect 1155 116 1156 120
rect 1150 115 1156 116
rect 1270 120 1276 121
rect 1270 116 1271 120
rect 1275 116 1276 120
rect 1270 115 1276 116
rect 1382 120 1388 121
rect 1382 116 1383 120
rect 1387 116 1388 120
rect 1382 115 1388 116
rect 1486 120 1492 121
rect 1486 116 1487 120
rect 1491 116 1492 120
rect 1486 115 1492 116
rect 1590 120 1596 121
rect 1590 116 1591 120
rect 1595 116 1596 120
rect 1590 115 1596 116
rect 1702 120 1708 121
rect 1702 116 1703 120
rect 1707 116 1708 120
rect 1702 115 1708 116
rect 1806 120 1812 121
rect 1806 116 1807 120
rect 1811 116 1812 120
rect 1806 115 1812 116
rect 1902 120 1908 121
rect 1902 116 1903 120
rect 1907 116 1908 120
rect 2006 119 2007 123
rect 2011 119 2012 123
rect 2046 123 2047 127
rect 2051 123 2052 127
rect 3942 127 3948 128
rect 2046 122 2052 123
rect 2070 124 2076 125
rect 2070 120 2071 124
rect 2075 120 2076 124
rect 2070 119 2076 120
rect 2166 124 2172 125
rect 2166 120 2167 124
rect 2171 120 2172 124
rect 2166 119 2172 120
rect 2262 124 2268 125
rect 2262 120 2263 124
rect 2267 120 2268 124
rect 2262 119 2268 120
rect 2358 124 2364 125
rect 2358 120 2359 124
rect 2363 120 2364 124
rect 2358 119 2364 120
rect 2454 124 2460 125
rect 2454 120 2455 124
rect 2459 120 2460 124
rect 2454 119 2460 120
rect 2550 124 2556 125
rect 2550 120 2551 124
rect 2555 120 2556 124
rect 2550 119 2556 120
rect 2654 124 2660 125
rect 2654 120 2655 124
rect 2659 120 2660 124
rect 2654 119 2660 120
rect 2758 124 2764 125
rect 2758 120 2759 124
rect 2763 120 2764 124
rect 2758 119 2764 120
rect 2862 124 2868 125
rect 2862 120 2863 124
rect 2867 120 2868 124
rect 2862 119 2868 120
rect 2974 124 2980 125
rect 2974 120 2975 124
rect 2979 120 2980 124
rect 2974 119 2980 120
rect 3102 124 3108 125
rect 3102 120 3103 124
rect 3107 120 3108 124
rect 3102 119 3108 120
rect 3238 124 3244 125
rect 3238 120 3239 124
rect 3243 120 3244 124
rect 3238 119 3244 120
rect 3382 124 3388 125
rect 3382 120 3383 124
rect 3387 120 3388 124
rect 3382 119 3388 120
rect 3534 124 3540 125
rect 3534 120 3535 124
rect 3539 120 3540 124
rect 3534 119 3540 120
rect 3694 124 3700 125
rect 3694 120 3695 124
rect 3699 120 3700 124
rect 3694 119 3700 120
rect 3838 124 3844 125
rect 3838 120 3839 124
rect 3843 120 3844 124
rect 3942 123 3943 127
rect 3947 123 3948 127
rect 3942 122 3948 123
rect 3838 119 3844 120
rect 2006 118 2012 119
rect 1902 115 1908 116
<< m3c >>
rect 111 4000 115 4004
rect 1519 3999 1523 4003
rect 1615 3999 1619 4003
rect 1711 3999 1715 4003
rect 1807 3999 1811 4003
rect 1903 3999 1907 4003
rect 2007 4000 2011 4004
rect 111 3983 115 3987
rect 1519 3980 1523 3984
rect 1615 3980 1619 3984
rect 1711 3980 1715 3984
rect 1807 3980 1811 3984
rect 1903 3980 1907 3984
rect 2007 3983 2011 3987
rect 2047 3981 2051 3985
rect 2071 3984 2075 3988
rect 2167 3984 2171 3988
rect 2263 3984 2267 3988
rect 3943 3981 3947 3985
rect 2047 3964 2051 3968
rect 2071 3965 2075 3969
rect 2167 3965 2171 3969
rect 2263 3965 2267 3969
rect 3943 3964 3947 3968
rect 111 3917 115 3921
rect 199 3920 203 3924
rect 295 3920 299 3924
rect 391 3920 395 3924
rect 495 3920 499 3924
rect 615 3920 619 3924
rect 743 3920 747 3924
rect 871 3920 875 3924
rect 999 3920 1003 3924
rect 1127 3920 1131 3924
rect 1255 3920 1259 3924
rect 1383 3920 1387 3924
rect 1511 3920 1515 3924
rect 1647 3920 1651 3924
rect 2007 3917 2011 3921
rect 2047 3912 2051 3916
rect 2159 3911 2163 3915
rect 2287 3911 2291 3915
rect 2415 3911 2419 3915
rect 2551 3911 2555 3915
rect 2687 3911 2691 3915
rect 2823 3911 2827 3915
rect 2951 3911 2955 3915
rect 3071 3911 3075 3915
rect 3191 3911 3195 3915
rect 3303 3911 3307 3915
rect 3407 3911 3411 3915
rect 3519 3911 3523 3915
rect 3631 3911 3635 3915
rect 3743 3911 3747 3915
rect 3943 3912 3947 3916
rect 111 3900 115 3904
rect 199 3901 203 3905
rect 295 3901 299 3905
rect 391 3901 395 3905
rect 495 3901 499 3905
rect 615 3901 619 3905
rect 743 3901 747 3905
rect 871 3901 875 3905
rect 999 3901 1003 3905
rect 1127 3901 1131 3905
rect 1255 3901 1259 3905
rect 1383 3901 1387 3905
rect 1511 3901 1515 3905
rect 1647 3901 1651 3905
rect 2007 3900 2011 3904
rect 2047 3895 2051 3899
rect 2159 3892 2163 3896
rect 2287 3892 2291 3896
rect 2415 3892 2419 3896
rect 2551 3892 2555 3896
rect 2687 3892 2691 3896
rect 2823 3892 2827 3896
rect 2951 3892 2955 3896
rect 3071 3892 3075 3896
rect 3191 3892 3195 3896
rect 3303 3892 3307 3896
rect 3407 3892 3411 3896
rect 3519 3892 3523 3896
rect 3631 3892 3635 3896
rect 3743 3892 3747 3896
rect 3943 3895 3947 3899
rect 111 3848 115 3852
rect 335 3847 339 3851
rect 455 3847 459 3851
rect 583 3847 587 3851
rect 719 3847 723 3851
rect 847 3847 851 3851
rect 975 3847 979 3851
rect 1103 3847 1107 3851
rect 1231 3847 1235 3851
rect 1359 3847 1363 3851
rect 1487 3847 1491 3851
rect 2007 3848 2011 3852
rect 111 3831 115 3835
rect 335 3828 339 3832
rect 455 3828 459 3832
rect 583 3828 587 3832
rect 719 3828 723 3832
rect 847 3828 851 3832
rect 975 3828 979 3832
rect 1103 3828 1107 3832
rect 1231 3828 1235 3832
rect 1359 3828 1363 3832
rect 1487 3828 1491 3832
rect 2007 3831 2011 3835
rect 2047 3821 2051 3825
rect 2207 3824 2211 3828
rect 2343 3824 2347 3828
rect 2487 3824 2491 3828
rect 2647 3824 2651 3828
rect 2823 3824 2827 3828
rect 3015 3824 3019 3828
rect 3223 3824 3227 3828
rect 3439 3824 3443 3828
rect 3655 3824 3659 3828
rect 3943 3821 3947 3825
rect 2047 3804 2051 3808
rect 2207 3805 2211 3809
rect 2343 3805 2347 3809
rect 2487 3805 2491 3809
rect 2647 3805 2651 3809
rect 2823 3805 2827 3809
rect 3015 3805 3019 3809
rect 3223 3805 3227 3809
rect 3439 3805 3443 3809
rect 3655 3805 3659 3809
rect 3943 3804 3947 3808
rect 111 3761 115 3765
rect 503 3764 507 3768
rect 615 3764 619 3768
rect 735 3764 739 3768
rect 863 3764 867 3768
rect 999 3764 1003 3768
rect 1143 3764 1147 3768
rect 1287 3764 1291 3768
rect 1431 3764 1435 3768
rect 1583 3764 1587 3768
rect 2007 3761 2011 3765
rect 2047 3752 2051 3756
rect 2191 3751 2195 3755
rect 2375 3751 2379 3755
rect 2559 3751 2563 3755
rect 2743 3751 2747 3755
rect 2935 3751 2939 3755
rect 3127 3751 3131 3755
rect 3319 3751 3323 3755
rect 3511 3751 3515 3755
rect 3711 3751 3715 3755
rect 3943 3752 3947 3756
rect 111 3744 115 3748
rect 503 3745 507 3749
rect 615 3745 619 3749
rect 735 3745 739 3749
rect 863 3745 867 3749
rect 999 3745 1003 3749
rect 1143 3745 1147 3749
rect 1287 3745 1291 3749
rect 1431 3745 1435 3749
rect 1583 3745 1587 3749
rect 2007 3744 2011 3748
rect 2047 3735 2051 3739
rect 2191 3732 2195 3736
rect 2375 3732 2379 3736
rect 2559 3732 2563 3736
rect 2743 3732 2747 3736
rect 2935 3732 2939 3736
rect 3127 3732 3131 3736
rect 3319 3732 3323 3736
rect 3511 3732 3515 3736
rect 3711 3732 3715 3736
rect 3943 3735 3947 3739
rect 111 3684 115 3688
rect 495 3683 499 3687
rect 591 3683 595 3687
rect 687 3683 691 3687
rect 791 3683 795 3687
rect 911 3683 915 3687
rect 1039 3683 1043 3687
rect 1183 3683 1187 3687
rect 1335 3683 1339 3687
rect 1495 3683 1499 3687
rect 1655 3683 1659 3687
rect 2007 3684 2011 3688
rect 111 3667 115 3671
rect 495 3664 499 3668
rect 591 3664 595 3668
rect 687 3664 691 3668
rect 791 3664 795 3668
rect 911 3664 915 3668
rect 1039 3664 1043 3668
rect 1183 3664 1187 3668
rect 1335 3664 1339 3668
rect 1495 3664 1499 3668
rect 1655 3664 1659 3668
rect 2007 3667 2011 3671
rect 2047 3665 2051 3669
rect 2127 3668 2131 3672
rect 2351 3668 2355 3672
rect 2583 3668 2587 3672
rect 2815 3668 2819 3672
rect 3047 3668 3051 3672
rect 3279 3668 3283 3672
rect 3511 3668 3515 3672
rect 3751 3668 3755 3672
rect 3943 3665 3947 3669
rect 2047 3648 2051 3652
rect 2127 3649 2131 3653
rect 2351 3649 2355 3653
rect 2583 3649 2587 3653
rect 2815 3649 2819 3653
rect 3047 3649 3051 3653
rect 3279 3649 3283 3653
rect 3511 3649 3515 3653
rect 3751 3649 3755 3653
rect 3943 3648 3947 3652
rect 111 3593 115 3597
rect 335 3596 339 3600
rect 463 3596 467 3600
rect 607 3596 611 3600
rect 759 3596 763 3600
rect 927 3596 931 3600
rect 1095 3596 1099 3600
rect 1263 3596 1267 3600
rect 1439 3596 1443 3600
rect 1615 3596 1619 3600
rect 1791 3596 1795 3600
rect 2007 3593 2011 3597
rect 2047 3588 2051 3592
rect 2191 3587 2195 3591
rect 2327 3587 2331 3591
rect 2455 3587 2459 3591
rect 2583 3587 2587 3591
rect 2719 3587 2723 3591
rect 2855 3587 2859 3591
rect 2999 3587 3003 3591
rect 3143 3587 3147 3591
rect 3295 3587 3299 3591
rect 3455 3587 3459 3591
rect 3623 3587 3627 3591
rect 3943 3588 3947 3592
rect 111 3576 115 3580
rect 335 3577 339 3581
rect 463 3577 467 3581
rect 607 3577 611 3581
rect 759 3577 763 3581
rect 927 3577 931 3581
rect 1095 3577 1099 3581
rect 1263 3577 1267 3581
rect 1439 3577 1443 3581
rect 1615 3577 1619 3581
rect 1791 3577 1795 3581
rect 2007 3576 2011 3580
rect 2047 3571 2051 3575
rect 2191 3568 2195 3572
rect 2327 3568 2331 3572
rect 2455 3568 2459 3572
rect 2583 3568 2587 3572
rect 2719 3568 2723 3572
rect 2855 3568 2859 3572
rect 2999 3568 3003 3572
rect 3143 3568 3147 3572
rect 3295 3568 3299 3572
rect 3455 3568 3459 3572
rect 3623 3568 3627 3572
rect 3943 3571 3947 3575
rect 111 3512 115 3516
rect 159 3511 163 3515
rect 303 3511 307 3515
rect 463 3511 467 3515
rect 639 3511 643 3515
rect 815 3511 819 3515
rect 999 3511 1003 3515
rect 1175 3511 1179 3515
rect 1351 3511 1355 3515
rect 1527 3511 1531 3515
rect 1703 3511 1707 3515
rect 1879 3511 1883 3515
rect 2007 3512 2011 3516
rect 2047 3505 2051 3509
rect 2103 3508 2107 3512
rect 2271 3508 2275 3512
rect 2447 3508 2451 3512
rect 2631 3508 2635 3512
rect 2815 3508 2819 3512
rect 2999 3508 3003 3512
rect 3175 3508 3179 3512
rect 3351 3508 3355 3512
rect 3519 3508 3523 3512
rect 3687 3508 3691 3512
rect 3839 3508 3843 3512
rect 3943 3505 3947 3509
rect 111 3495 115 3499
rect 159 3492 163 3496
rect 303 3492 307 3496
rect 463 3492 467 3496
rect 639 3492 643 3496
rect 815 3492 819 3496
rect 999 3492 1003 3496
rect 1175 3492 1179 3496
rect 1351 3492 1355 3496
rect 1527 3492 1531 3496
rect 1703 3492 1707 3496
rect 1879 3492 1883 3496
rect 2007 3495 2011 3499
rect 2047 3488 2051 3492
rect 2103 3489 2107 3493
rect 2271 3489 2275 3493
rect 2447 3489 2451 3493
rect 2631 3489 2635 3493
rect 2815 3489 2819 3493
rect 2999 3489 3003 3493
rect 3175 3489 3179 3493
rect 3351 3489 3355 3493
rect 3519 3489 3523 3493
rect 3687 3489 3691 3493
rect 3839 3489 3843 3493
rect 3943 3488 3947 3492
rect 2047 3432 2051 3436
rect 2127 3431 2131 3435
rect 2311 3431 2315 3435
rect 2495 3431 2499 3435
rect 2679 3431 2683 3435
rect 2863 3431 2867 3435
rect 3047 3431 3051 3435
rect 3223 3431 3227 3435
rect 3407 3431 3411 3435
rect 3591 3431 3595 3435
rect 3775 3431 3779 3435
rect 3943 3432 3947 3436
rect 111 3421 115 3425
rect 135 3424 139 3428
rect 319 3424 323 3428
rect 535 3424 539 3428
rect 751 3424 755 3428
rect 959 3424 963 3428
rect 1159 3424 1163 3428
rect 1351 3424 1355 3428
rect 1535 3424 1539 3428
rect 1719 3424 1723 3428
rect 1903 3424 1907 3428
rect 2007 3421 2011 3425
rect 2047 3415 2051 3419
rect 2127 3412 2131 3416
rect 2311 3412 2315 3416
rect 2495 3412 2499 3416
rect 2679 3412 2683 3416
rect 2863 3412 2867 3416
rect 3047 3412 3051 3416
rect 3223 3412 3227 3416
rect 3407 3412 3411 3416
rect 3591 3412 3595 3416
rect 3775 3412 3779 3416
rect 3943 3415 3947 3419
rect 111 3404 115 3408
rect 135 3405 139 3409
rect 319 3405 323 3409
rect 535 3405 539 3409
rect 751 3405 755 3409
rect 959 3405 963 3409
rect 1159 3405 1163 3409
rect 1351 3405 1355 3409
rect 1535 3405 1539 3409
rect 1719 3405 1723 3409
rect 1903 3405 1907 3409
rect 2007 3404 2011 3408
rect 111 3352 115 3356
rect 135 3351 139 3355
rect 231 3351 235 3355
rect 375 3351 379 3355
rect 535 3351 539 3355
rect 703 3351 707 3355
rect 871 3351 875 3355
rect 1047 3351 1051 3355
rect 1215 3351 1219 3355
rect 1383 3351 1387 3355
rect 1543 3351 1547 3355
rect 1703 3351 1707 3355
rect 1871 3351 1875 3355
rect 2007 3352 2011 3356
rect 111 3335 115 3339
rect 135 3332 139 3336
rect 231 3332 235 3336
rect 375 3332 379 3336
rect 535 3332 539 3336
rect 703 3332 707 3336
rect 871 3332 875 3336
rect 1047 3332 1051 3336
rect 1215 3332 1219 3336
rect 1383 3332 1387 3336
rect 1543 3332 1547 3336
rect 1703 3332 1707 3336
rect 1871 3332 1875 3336
rect 2007 3335 2011 3339
rect 2047 3333 2051 3337
rect 2071 3336 2075 3340
rect 2215 3336 2219 3340
rect 2359 3336 2363 3340
rect 2511 3336 2515 3340
rect 2655 3336 2659 3340
rect 2799 3336 2803 3340
rect 2935 3336 2939 3340
rect 3079 3336 3083 3340
rect 3223 3336 3227 3340
rect 3375 3336 3379 3340
rect 3535 3336 3539 3340
rect 3695 3336 3699 3340
rect 3839 3336 3843 3340
rect 3943 3333 3947 3337
rect 2047 3316 2051 3320
rect 2071 3317 2075 3321
rect 2215 3317 2219 3321
rect 2359 3317 2363 3321
rect 2511 3317 2515 3321
rect 2655 3317 2659 3321
rect 2799 3317 2803 3321
rect 2935 3317 2939 3321
rect 3079 3317 3083 3321
rect 3223 3317 3227 3321
rect 3375 3317 3379 3321
rect 3535 3317 3539 3321
rect 3695 3317 3699 3321
rect 3839 3317 3843 3321
rect 3943 3316 3947 3320
rect 111 3269 115 3273
rect 135 3272 139 3276
rect 279 3272 283 3276
rect 463 3272 467 3276
rect 663 3272 667 3276
rect 871 3272 875 3276
rect 1079 3272 1083 3276
rect 1295 3272 1299 3276
rect 1519 3272 1523 3276
rect 1743 3272 1747 3276
rect 2007 3269 2011 3273
rect 111 3252 115 3256
rect 135 3253 139 3257
rect 279 3253 283 3257
rect 463 3253 467 3257
rect 663 3253 667 3257
rect 871 3253 875 3257
rect 1079 3253 1083 3257
rect 1295 3253 1299 3257
rect 1519 3253 1523 3257
rect 1743 3253 1747 3257
rect 2007 3252 2011 3256
rect 2047 3256 2051 3260
rect 2111 3255 2115 3259
rect 2247 3255 2251 3259
rect 2399 3255 2403 3259
rect 2575 3255 2579 3259
rect 2783 3255 2787 3259
rect 3015 3255 3019 3259
rect 3263 3255 3267 3259
rect 3527 3255 3531 3259
rect 3791 3255 3795 3259
rect 3943 3256 3947 3260
rect 2047 3239 2051 3243
rect 2111 3236 2115 3240
rect 2247 3236 2251 3240
rect 2399 3236 2403 3240
rect 2575 3236 2579 3240
rect 2783 3236 2787 3240
rect 3015 3236 3019 3240
rect 3263 3236 3267 3240
rect 3527 3236 3531 3240
rect 3791 3236 3795 3240
rect 3943 3239 3947 3243
rect 111 3200 115 3204
rect 135 3199 139 3203
rect 287 3199 291 3203
rect 447 3199 451 3203
rect 615 3199 619 3203
rect 791 3199 795 3203
rect 967 3199 971 3203
rect 1143 3199 1147 3203
rect 1327 3199 1331 3203
rect 1511 3199 1515 3203
rect 1695 3199 1699 3203
rect 2007 3200 2011 3204
rect 111 3183 115 3187
rect 135 3180 139 3184
rect 287 3180 291 3184
rect 447 3180 451 3184
rect 615 3180 619 3184
rect 791 3180 795 3184
rect 967 3180 971 3184
rect 1143 3180 1147 3184
rect 1327 3180 1331 3184
rect 1511 3180 1515 3184
rect 1695 3180 1699 3184
rect 2007 3183 2011 3187
rect 2047 3173 2051 3177
rect 2071 3176 2075 3180
rect 2167 3176 2171 3180
rect 2263 3176 2267 3180
rect 2359 3176 2363 3180
rect 2455 3176 2459 3180
rect 2551 3176 2555 3180
rect 2647 3176 2651 3180
rect 2743 3176 2747 3180
rect 2839 3176 2843 3180
rect 2935 3176 2939 3180
rect 3031 3176 3035 3180
rect 3127 3176 3131 3180
rect 3223 3176 3227 3180
rect 3319 3176 3323 3180
rect 3439 3176 3443 3180
rect 3575 3176 3579 3180
rect 3719 3176 3723 3180
rect 3839 3176 3843 3180
rect 3943 3173 3947 3177
rect 2047 3156 2051 3160
rect 2071 3157 2075 3161
rect 2167 3157 2171 3161
rect 2263 3157 2267 3161
rect 2359 3157 2363 3161
rect 2455 3157 2459 3161
rect 2551 3157 2555 3161
rect 2647 3157 2651 3161
rect 2743 3157 2747 3161
rect 2839 3157 2843 3161
rect 2935 3157 2939 3161
rect 3031 3157 3035 3161
rect 3127 3157 3131 3161
rect 3223 3157 3227 3161
rect 3319 3157 3323 3161
rect 3439 3157 3443 3161
rect 3575 3157 3579 3161
rect 3719 3157 3723 3161
rect 3839 3157 3843 3161
rect 3943 3156 3947 3160
rect 111 3113 115 3117
rect 311 3116 315 3120
rect 439 3116 443 3120
rect 583 3116 587 3120
rect 743 3116 747 3120
rect 903 3116 907 3120
rect 1063 3116 1067 3120
rect 1223 3116 1227 3120
rect 1391 3116 1395 3120
rect 1559 3116 1563 3120
rect 1727 3116 1731 3120
rect 2007 3113 2011 3117
rect 111 3096 115 3100
rect 311 3097 315 3101
rect 439 3097 443 3101
rect 583 3097 587 3101
rect 743 3097 747 3101
rect 903 3097 907 3101
rect 1063 3097 1067 3101
rect 1223 3097 1227 3101
rect 1391 3097 1395 3101
rect 1559 3097 1563 3101
rect 1727 3097 1731 3101
rect 2007 3096 2011 3100
rect 2047 3092 2051 3096
rect 2071 3091 2075 3095
rect 2335 3091 2339 3095
rect 2623 3091 2627 3095
rect 2911 3091 2915 3095
rect 3207 3091 3211 3095
rect 3503 3091 3507 3095
rect 3799 3091 3803 3095
rect 3943 3092 3947 3096
rect 2047 3075 2051 3079
rect 2071 3072 2075 3076
rect 2335 3072 2339 3076
rect 2623 3072 2627 3076
rect 2911 3072 2915 3076
rect 3207 3072 3211 3076
rect 3503 3072 3507 3076
rect 3799 3072 3803 3076
rect 3943 3075 3947 3079
rect 111 3036 115 3040
rect 503 3035 507 3039
rect 599 3035 603 3039
rect 703 3035 707 3039
rect 815 3035 819 3039
rect 935 3035 939 3039
rect 1071 3035 1075 3039
rect 1223 3035 1227 3039
rect 1383 3035 1387 3039
rect 1551 3035 1555 3039
rect 1719 3035 1723 3039
rect 2007 3036 2011 3040
rect 111 3019 115 3023
rect 503 3016 507 3020
rect 599 3016 603 3020
rect 703 3016 707 3020
rect 815 3016 819 3020
rect 935 3016 939 3020
rect 1071 3016 1075 3020
rect 1223 3016 1227 3020
rect 1383 3016 1387 3020
rect 1551 3016 1555 3020
rect 1719 3016 1723 3020
rect 2007 3019 2011 3023
rect 2047 3009 2051 3013
rect 2071 3012 2075 3016
rect 2383 3012 2387 3016
rect 2703 3012 2707 3016
rect 2999 3012 3003 3016
rect 3287 3012 3291 3016
rect 3575 3012 3579 3016
rect 3839 3012 3843 3016
rect 3943 3009 3947 3013
rect 2047 2992 2051 2996
rect 2071 2993 2075 2997
rect 2383 2993 2387 2997
rect 2703 2993 2707 2997
rect 2999 2993 3003 2997
rect 3287 2993 3291 2997
rect 3575 2993 3579 2997
rect 3839 2993 3843 2997
rect 3943 2992 3947 2996
rect 111 2949 115 2953
rect 551 2952 555 2956
rect 647 2952 651 2956
rect 759 2952 763 2956
rect 887 2952 891 2956
rect 1023 2952 1027 2956
rect 1175 2952 1179 2956
rect 1327 2952 1331 2956
rect 1487 2952 1491 2956
rect 1655 2952 1659 2956
rect 1823 2952 1827 2956
rect 2007 2949 2011 2953
rect 111 2932 115 2936
rect 551 2933 555 2937
rect 647 2933 651 2937
rect 759 2933 763 2937
rect 887 2933 891 2937
rect 1023 2933 1027 2937
rect 1175 2933 1179 2937
rect 1327 2933 1331 2937
rect 1487 2933 1491 2937
rect 1655 2933 1659 2937
rect 1823 2933 1827 2937
rect 2007 2932 2011 2936
rect 2047 2936 2051 2940
rect 2071 2935 2075 2939
rect 2391 2935 2395 2939
rect 2703 2935 2707 2939
rect 2975 2935 2979 2939
rect 3215 2935 3219 2939
rect 3439 2935 3443 2939
rect 3647 2935 3651 2939
rect 3839 2935 3843 2939
rect 3943 2936 3947 2940
rect 2047 2919 2051 2923
rect 2071 2916 2075 2920
rect 2391 2916 2395 2920
rect 2703 2916 2707 2920
rect 2975 2916 2979 2920
rect 3215 2916 3219 2920
rect 3439 2916 3443 2920
rect 3647 2916 3651 2920
rect 3839 2916 3843 2920
rect 3943 2919 3947 2923
rect 111 2872 115 2876
rect 471 2871 475 2875
rect 575 2871 579 2875
rect 695 2871 699 2875
rect 839 2871 843 2875
rect 991 2871 995 2875
rect 1151 2871 1155 2875
rect 1319 2871 1323 2875
rect 1495 2871 1499 2875
rect 1671 2871 1675 2875
rect 1847 2871 1851 2875
rect 2007 2872 2011 2876
rect 111 2855 115 2859
rect 471 2852 475 2856
rect 575 2852 579 2856
rect 695 2852 699 2856
rect 839 2852 843 2856
rect 991 2852 995 2856
rect 1151 2852 1155 2856
rect 1319 2852 1323 2856
rect 1495 2852 1499 2856
rect 1671 2852 1675 2856
rect 1847 2852 1851 2856
rect 2007 2855 2011 2859
rect 2047 2853 2051 2857
rect 2071 2856 2075 2860
rect 2295 2856 2299 2860
rect 2535 2856 2539 2860
rect 2767 2856 2771 2860
rect 2991 2856 2995 2860
rect 3215 2856 3219 2860
rect 3431 2856 3435 2860
rect 3647 2856 3651 2860
rect 3839 2856 3843 2860
rect 3943 2853 3947 2857
rect 2047 2836 2051 2840
rect 2071 2837 2075 2841
rect 2295 2837 2299 2841
rect 2535 2837 2539 2841
rect 2767 2837 2771 2841
rect 2991 2837 2995 2841
rect 3215 2837 3219 2841
rect 3431 2837 3435 2841
rect 3647 2837 3651 2841
rect 3839 2837 3843 2841
rect 3943 2836 3947 2840
rect 111 2785 115 2789
rect 479 2788 483 2792
rect 575 2788 579 2792
rect 679 2788 683 2792
rect 799 2788 803 2792
rect 935 2788 939 2792
rect 1079 2788 1083 2792
rect 1239 2788 1243 2792
rect 1415 2788 1419 2792
rect 1599 2788 1603 2792
rect 1783 2788 1787 2792
rect 2007 2785 2011 2789
rect 2047 2780 2051 2784
rect 2071 2779 2075 2783
rect 2199 2779 2203 2783
rect 2367 2779 2371 2783
rect 2551 2779 2555 2783
rect 2735 2779 2739 2783
rect 2927 2779 2931 2783
rect 3111 2779 3115 2783
rect 3295 2779 3299 2783
rect 3479 2779 3483 2783
rect 3671 2779 3675 2783
rect 3839 2779 3843 2783
rect 3943 2780 3947 2784
rect 111 2768 115 2772
rect 479 2769 483 2773
rect 575 2769 579 2773
rect 679 2769 683 2773
rect 799 2769 803 2773
rect 935 2769 939 2773
rect 1079 2769 1083 2773
rect 1239 2769 1243 2773
rect 1415 2769 1419 2773
rect 1599 2769 1603 2773
rect 1783 2769 1787 2773
rect 2007 2768 2011 2772
rect 2047 2763 2051 2767
rect 2071 2760 2075 2764
rect 2199 2760 2203 2764
rect 2367 2760 2371 2764
rect 2551 2760 2555 2764
rect 2735 2760 2739 2764
rect 2927 2760 2931 2764
rect 3111 2760 3115 2764
rect 3295 2760 3299 2764
rect 3479 2760 3483 2764
rect 3671 2760 3675 2764
rect 3839 2760 3843 2764
rect 3943 2763 3947 2767
rect 111 2712 115 2716
rect 511 2711 515 2715
rect 623 2711 627 2715
rect 743 2711 747 2715
rect 879 2711 883 2715
rect 1015 2711 1019 2715
rect 1159 2711 1163 2715
rect 1311 2711 1315 2715
rect 1463 2711 1467 2715
rect 1623 2711 1627 2715
rect 1783 2711 1787 2715
rect 2007 2712 2011 2716
rect 111 2695 115 2699
rect 511 2692 515 2696
rect 623 2692 627 2696
rect 743 2692 747 2696
rect 879 2692 883 2696
rect 1015 2692 1019 2696
rect 1159 2692 1163 2696
rect 1311 2692 1315 2696
rect 1463 2692 1467 2696
rect 1623 2692 1627 2696
rect 1783 2692 1787 2696
rect 2007 2695 2011 2699
rect 2047 2693 2051 2697
rect 2071 2696 2075 2700
rect 2191 2696 2195 2700
rect 2319 2696 2323 2700
rect 2447 2696 2451 2700
rect 2583 2696 2587 2700
rect 2727 2696 2731 2700
rect 2887 2696 2891 2700
rect 3063 2696 3067 2700
rect 3255 2696 3259 2700
rect 3455 2696 3459 2700
rect 3655 2696 3659 2700
rect 3839 2696 3843 2700
rect 3943 2693 3947 2697
rect 2047 2676 2051 2680
rect 2071 2677 2075 2681
rect 2191 2677 2195 2681
rect 2319 2677 2323 2681
rect 2447 2677 2451 2681
rect 2583 2677 2587 2681
rect 2727 2677 2731 2681
rect 2887 2677 2891 2681
rect 3063 2677 3067 2681
rect 3255 2677 3259 2681
rect 3455 2677 3459 2681
rect 3655 2677 3659 2681
rect 3839 2677 3843 2681
rect 3943 2676 3947 2680
rect 111 2625 115 2629
rect 367 2628 371 2632
rect 487 2628 491 2632
rect 615 2628 619 2632
rect 751 2628 755 2632
rect 895 2628 899 2632
rect 1031 2628 1035 2632
rect 1167 2628 1171 2632
rect 1303 2628 1307 2632
rect 1431 2628 1435 2632
rect 1567 2628 1571 2632
rect 1703 2628 1707 2632
rect 2007 2625 2011 2629
rect 2047 2616 2051 2620
rect 2231 2615 2235 2619
rect 2335 2615 2339 2619
rect 2447 2615 2451 2619
rect 2559 2615 2563 2619
rect 2671 2615 2675 2619
rect 2791 2615 2795 2619
rect 2911 2615 2915 2619
rect 3031 2615 3035 2619
rect 3151 2615 3155 2619
rect 3943 2616 3947 2620
rect 111 2608 115 2612
rect 367 2609 371 2613
rect 487 2609 491 2613
rect 615 2609 619 2613
rect 751 2609 755 2613
rect 895 2609 899 2613
rect 1031 2609 1035 2613
rect 1167 2609 1171 2613
rect 1303 2609 1307 2613
rect 1431 2609 1435 2613
rect 1567 2609 1571 2613
rect 1703 2609 1707 2613
rect 2007 2608 2011 2612
rect 2047 2599 2051 2603
rect 2231 2596 2235 2600
rect 2335 2596 2339 2600
rect 2447 2596 2451 2600
rect 2559 2596 2563 2600
rect 2671 2596 2675 2600
rect 2791 2596 2795 2600
rect 2911 2596 2915 2600
rect 3031 2596 3035 2600
rect 3151 2596 3155 2600
rect 3943 2599 3947 2603
rect 111 2556 115 2560
rect 135 2555 139 2559
rect 287 2555 291 2559
rect 447 2555 451 2559
rect 607 2555 611 2559
rect 767 2555 771 2559
rect 919 2555 923 2559
rect 1063 2555 1067 2559
rect 1199 2555 1203 2559
rect 1335 2555 1339 2559
rect 1463 2555 1467 2559
rect 1591 2555 1595 2559
rect 1727 2555 1731 2559
rect 2007 2556 2011 2560
rect 111 2539 115 2543
rect 135 2536 139 2540
rect 287 2536 291 2540
rect 447 2536 451 2540
rect 607 2536 611 2540
rect 767 2536 771 2540
rect 919 2536 923 2540
rect 1063 2536 1067 2540
rect 1199 2536 1203 2540
rect 1335 2536 1339 2540
rect 1463 2536 1467 2540
rect 1591 2536 1595 2540
rect 1727 2536 1731 2540
rect 2007 2539 2011 2543
rect 2047 2529 2051 2533
rect 2383 2532 2387 2536
rect 2495 2532 2499 2536
rect 2615 2532 2619 2536
rect 2743 2532 2747 2536
rect 2871 2532 2875 2536
rect 2991 2532 2995 2536
rect 3111 2532 3115 2536
rect 3231 2532 3235 2536
rect 3359 2532 3363 2536
rect 3487 2532 3491 2536
rect 3943 2529 3947 2533
rect 2047 2512 2051 2516
rect 2383 2513 2387 2517
rect 2495 2513 2499 2517
rect 2615 2513 2619 2517
rect 2743 2513 2747 2517
rect 2871 2513 2875 2517
rect 2991 2513 2995 2517
rect 3111 2513 3115 2517
rect 3231 2513 3235 2517
rect 3359 2513 3363 2517
rect 3487 2513 3491 2517
rect 3943 2512 3947 2516
rect 111 2457 115 2461
rect 135 2460 139 2464
rect 231 2460 235 2464
rect 327 2460 331 2464
rect 423 2460 427 2464
rect 519 2460 523 2464
rect 2007 2457 2011 2461
rect 2047 2456 2051 2460
rect 2535 2455 2539 2459
rect 2711 2455 2715 2459
rect 2879 2455 2883 2459
rect 3047 2455 3051 2459
rect 3207 2455 3211 2459
rect 3359 2455 3363 2459
rect 3503 2455 3507 2459
rect 3655 2455 3659 2459
rect 3807 2455 3811 2459
rect 3943 2456 3947 2460
rect 111 2440 115 2444
rect 135 2441 139 2445
rect 231 2441 235 2445
rect 327 2441 331 2445
rect 423 2441 427 2445
rect 519 2441 523 2445
rect 2007 2440 2011 2444
rect 2047 2439 2051 2443
rect 2535 2436 2539 2440
rect 2711 2436 2715 2440
rect 2879 2436 2883 2440
rect 3047 2436 3051 2440
rect 3207 2436 3211 2440
rect 3359 2436 3363 2440
rect 3503 2436 3507 2440
rect 3655 2436 3659 2440
rect 3807 2436 3811 2440
rect 3943 2439 3947 2443
rect 111 2372 115 2376
rect 135 2371 139 2375
rect 255 2371 259 2375
rect 415 2371 419 2375
rect 575 2371 579 2375
rect 735 2371 739 2375
rect 887 2371 891 2375
rect 1039 2371 1043 2375
rect 1183 2371 1187 2375
rect 1327 2371 1331 2375
rect 1479 2371 1483 2375
rect 2007 2372 2011 2376
rect 2047 2361 2051 2365
rect 2607 2364 2611 2368
rect 2815 2364 2819 2368
rect 3007 2364 3011 2368
rect 3191 2364 3195 2368
rect 3359 2364 3363 2368
rect 3519 2364 3523 2368
rect 3679 2364 3683 2368
rect 3839 2364 3843 2368
rect 3943 2361 3947 2365
rect 111 2355 115 2359
rect 135 2352 139 2356
rect 255 2352 259 2356
rect 415 2352 419 2356
rect 575 2352 579 2356
rect 735 2352 739 2356
rect 887 2352 891 2356
rect 1039 2352 1043 2356
rect 1183 2352 1187 2356
rect 1327 2352 1331 2356
rect 1479 2352 1483 2356
rect 2007 2355 2011 2359
rect 2047 2344 2051 2348
rect 2607 2345 2611 2349
rect 2815 2345 2819 2349
rect 3007 2345 3011 2349
rect 3191 2345 3195 2349
rect 3359 2345 3363 2349
rect 3519 2345 3523 2349
rect 3679 2345 3683 2349
rect 3839 2345 3843 2349
rect 3943 2344 3947 2348
rect 111 2289 115 2293
rect 135 2292 139 2296
rect 263 2292 267 2296
rect 423 2292 427 2296
rect 583 2292 587 2296
rect 743 2292 747 2296
rect 895 2292 899 2296
rect 1047 2292 1051 2296
rect 1199 2292 1203 2296
rect 1351 2292 1355 2296
rect 1503 2292 1507 2296
rect 2007 2289 2011 2293
rect 111 2272 115 2276
rect 135 2273 139 2277
rect 263 2273 267 2277
rect 423 2273 427 2277
rect 583 2273 587 2277
rect 743 2273 747 2277
rect 895 2273 899 2277
rect 1047 2273 1051 2277
rect 1199 2273 1203 2277
rect 1351 2273 1355 2277
rect 1503 2273 1507 2277
rect 2007 2272 2011 2276
rect 2047 2276 2051 2280
rect 2071 2275 2075 2279
rect 2167 2275 2171 2279
rect 2271 2275 2275 2279
rect 2415 2275 2419 2279
rect 2575 2275 2579 2279
rect 2743 2275 2747 2279
rect 2911 2275 2915 2279
rect 3071 2275 3075 2279
rect 3231 2275 3235 2279
rect 3383 2275 3387 2279
rect 3535 2275 3539 2279
rect 3695 2275 3699 2279
rect 3943 2276 3947 2280
rect 2047 2259 2051 2263
rect 2071 2256 2075 2260
rect 2167 2256 2171 2260
rect 2271 2256 2275 2260
rect 2415 2256 2419 2260
rect 2575 2256 2579 2260
rect 2743 2256 2747 2260
rect 2911 2256 2915 2260
rect 3071 2256 3075 2260
rect 3231 2256 3235 2260
rect 3383 2256 3387 2260
rect 3535 2256 3539 2260
rect 3695 2256 3699 2260
rect 3943 2259 3947 2263
rect 111 2216 115 2220
rect 223 2215 227 2219
rect 351 2215 355 2219
rect 495 2215 499 2219
rect 647 2215 651 2219
rect 799 2215 803 2219
rect 959 2215 963 2219
rect 1119 2215 1123 2219
rect 1279 2215 1283 2219
rect 1439 2215 1443 2219
rect 1599 2215 1603 2219
rect 2007 2216 2011 2220
rect 111 2199 115 2203
rect 223 2196 227 2200
rect 351 2196 355 2200
rect 495 2196 499 2200
rect 647 2196 651 2200
rect 799 2196 803 2200
rect 959 2196 963 2200
rect 1119 2196 1123 2200
rect 1279 2196 1283 2200
rect 1439 2196 1443 2200
rect 1599 2196 1603 2200
rect 2007 2199 2011 2203
rect 2047 2193 2051 2197
rect 2071 2196 2075 2200
rect 2175 2196 2179 2200
rect 2319 2196 2323 2200
rect 2471 2196 2475 2200
rect 2623 2196 2627 2200
rect 2783 2196 2787 2200
rect 2935 2196 2939 2200
rect 3079 2196 3083 2200
rect 3223 2196 3227 2200
rect 3367 2196 3371 2200
rect 3519 2196 3523 2200
rect 3943 2193 3947 2197
rect 2047 2176 2051 2180
rect 2071 2177 2075 2181
rect 2175 2177 2179 2181
rect 2319 2177 2323 2181
rect 2471 2177 2475 2181
rect 2623 2177 2627 2181
rect 2783 2177 2787 2181
rect 2935 2177 2939 2181
rect 3079 2177 3083 2181
rect 3223 2177 3227 2181
rect 3367 2177 3371 2181
rect 3519 2177 3523 2181
rect 3943 2176 3947 2180
rect 111 2133 115 2137
rect 471 2136 475 2140
rect 567 2136 571 2140
rect 679 2136 683 2140
rect 807 2136 811 2140
rect 943 2136 947 2140
rect 1079 2136 1083 2140
rect 1223 2136 1227 2140
rect 1367 2136 1371 2140
rect 1503 2136 1507 2140
rect 1639 2136 1643 2140
rect 1783 2136 1787 2140
rect 1903 2136 1907 2140
rect 2007 2133 2011 2137
rect 111 2116 115 2120
rect 471 2117 475 2121
rect 567 2117 571 2121
rect 679 2117 683 2121
rect 807 2117 811 2121
rect 943 2117 947 2121
rect 1079 2117 1083 2121
rect 1223 2117 1227 2121
rect 1367 2117 1371 2121
rect 1503 2117 1507 2121
rect 1639 2117 1643 2121
rect 1783 2117 1787 2121
rect 1903 2117 1907 2121
rect 2007 2116 2011 2120
rect 2047 2104 2051 2108
rect 2279 2103 2283 2107
rect 2391 2103 2395 2107
rect 2511 2103 2515 2107
rect 2631 2103 2635 2107
rect 2759 2103 2763 2107
rect 2895 2103 2899 2107
rect 3039 2103 3043 2107
rect 3191 2103 3195 2107
rect 3351 2103 3355 2107
rect 3519 2103 3523 2107
rect 3687 2103 3691 2107
rect 3839 2103 3843 2107
rect 3943 2104 3947 2108
rect 2047 2087 2051 2091
rect 2279 2084 2283 2088
rect 2391 2084 2395 2088
rect 2511 2084 2515 2088
rect 2631 2084 2635 2088
rect 2759 2084 2763 2088
rect 2895 2084 2899 2088
rect 3039 2084 3043 2088
rect 3191 2084 3195 2088
rect 3351 2084 3355 2088
rect 3519 2084 3523 2088
rect 3687 2084 3691 2088
rect 3839 2084 3843 2088
rect 3943 2087 3947 2091
rect 111 2064 115 2068
rect 623 2063 627 2067
rect 735 2063 739 2067
rect 855 2063 859 2067
rect 983 2063 987 2067
rect 1119 2063 1123 2067
rect 1255 2063 1259 2067
rect 1391 2063 1395 2067
rect 1527 2063 1531 2067
rect 1655 2063 1659 2067
rect 1791 2063 1795 2067
rect 1903 2063 1907 2067
rect 2007 2064 2011 2068
rect 111 2047 115 2051
rect 623 2044 627 2048
rect 735 2044 739 2048
rect 855 2044 859 2048
rect 983 2044 987 2048
rect 1119 2044 1123 2048
rect 1255 2044 1259 2048
rect 1391 2044 1395 2048
rect 1527 2044 1531 2048
rect 1655 2044 1659 2048
rect 1791 2044 1795 2048
rect 1903 2044 1907 2048
rect 2007 2047 2011 2051
rect 2047 2013 2051 2017
rect 2327 2016 2331 2020
rect 2431 2016 2435 2020
rect 2535 2016 2539 2020
rect 2647 2016 2651 2020
rect 2775 2016 2779 2020
rect 2919 2016 2923 2020
rect 3079 2016 3083 2020
rect 3263 2016 3267 2020
rect 3455 2016 3459 2020
rect 3655 2016 3659 2020
rect 3839 2016 3843 2020
rect 3943 2013 3947 2017
rect 2047 1996 2051 2000
rect 2327 1997 2331 2001
rect 2431 1997 2435 2001
rect 2535 1997 2539 2001
rect 2647 1997 2651 2001
rect 2775 1997 2779 2001
rect 2919 1997 2923 2001
rect 3079 1997 3083 2001
rect 3263 1997 3267 2001
rect 3455 1997 3459 2001
rect 3655 1997 3659 2001
rect 3839 1997 3843 2001
rect 3943 1996 3947 2000
rect 111 1977 115 1981
rect 447 1980 451 1984
rect 575 1980 579 1984
rect 727 1980 731 1984
rect 887 1980 891 1984
rect 1055 1980 1059 1984
rect 1231 1980 1235 1984
rect 1399 1980 1403 1984
rect 1575 1980 1579 1984
rect 1751 1980 1755 1984
rect 1903 1980 1907 1984
rect 2007 1977 2011 1981
rect 111 1960 115 1964
rect 447 1961 451 1965
rect 575 1961 579 1965
rect 727 1961 731 1965
rect 887 1961 891 1965
rect 1055 1961 1059 1965
rect 1231 1961 1235 1965
rect 1399 1961 1403 1965
rect 1575 1961 1579 1965
rect 1751 1961 1755 1965
rect 1903 1961 1907 1965
rect 2007 1960 2011 1964
rect 2047 1940 2051 1944
rect 2255 1939 2259 1943
rect 2351 1939 2355 1943
rect 2447 1939 2451 1943
rect 2543 1939 2547 1943
rect 2647 1939 2651 1943
rect 2767 1939 2771 1943
rect 2919 1939 2923 1943
rect 3103 1939 3107 1943
rect 3319 1939 3323 1943
rect 3543 1939 3547 1943
rect 3775 1939 3779 1943
rect 3943 1940 3947 1944
rect 2047 1923 2051 1927
rect 2255 1920 2259 1924
rect 2351 1920 2355 1924
rect 2447 1920 2451 1924
rect 2543 1920 2547 1924
rect 2647 1920 2651 1924
rect 2767 1920 2771 1924
rect 2919 1920 2923 1924
rect 3103 1920 3107 1924
rect 3319 1920 3323 1924
rect 3543 1920 3547 1924
rect 3775 1920 3779 1924
rect 3943 1923 3947 1927
rect 111 1908 115 1912
rect 655 1907 659 1911
rect 751 1907 755 1911
rect 847 1907 851 1911
rect 943 1907 947 1911
rect 1039 1907 1043 1911
rect 1135 1907 1139 1911
rect 1231 1907 1235 1911
rect 1327 1907 1331 1911
rect 1423 1907 1427 1911
rect 2007 1908 2011 1912
rect 111 1891 115 1895
rect 655 1888 659 1892
rect 751 1888 755 1892
rect 847 1888 851 1892
rect 943 1888 947 1892
rect 1039 1888 1043 1892
rect 1135 1888 1139 1892
rect 1231 1888 1235 1892
rect 1327 1888 1331 1892
rect 1423 1888 1427 1892
rect 2007 1891 2011 1895
rect 2047 1845 2051 1849
rect 2183 1848 2187 1852
rect 2279 1848 2283 1852
rect 2383 1848 2387 1852
rect 2487 1848 2491 1852
rect 2591 1848 2595 1852
rect 2703 1848 2707 1852
rect 2831 1848 2835 1852
rect 2991 1848 2995 1852
rect 3183 1848 3187 1852
rect 3399 1848 3403 1852
rect 3631 1848 3635 1852
rect 3839 1848 3843 1852
rect 3943 1845 3947 1849
rect 111 1825 115 1829
rect 319 1828 323 1832
rect 447 1828 451 1832
rect 583 1828 587 1832
rect 719 1828 723 1832
rect 855 1828 859 1832
rect 991 1828 995 1832
rect 1127 1828 1131 1832
rect 1263 1828 1267 1832
rect 1399 1828 1403 1832
rect 1535 1828 1539 1832
rect 2007 1825 2011 1829
rect 2047 1828 2051 1832
rect 2183 1829 2187 1833
rect 2279 1829 2283 1833
rect 2383 1829 2387 1833
rect 2487 1829 2491 1833
rect 2591 1829 2595 1833
rect 2703 1829 2707 1833
rect 2831 1829 2835 1833
rect 2991 1829 2995 1833
rect 3183 1829 3187 1833
rect 3399 1829 3403 1833
rect 3631 1829 3635 1833
rect 3839 1829 3843 1833
rect 3943 1828 3947 1832
rect 111 1808 115 1812
rect 319 1809 323 1813
rect 447 1809 451 1813
rect 583 1809 587 1813
rect 719 1809 723 1813
rect 855 1809 859 1813
rect 991 1809 995 1813
rect 1127 1809 1131 1813
rect 1263 1809 1267 1813
rect 1399 1809 1403 1813
rect 1535 1809 1539 1813
rect 2007 1808 2011 1812
rect 2047 1772 2051 1776
rect 2127 1771 2131 1775
rect 2311 1771 2315 1775
rect 2495 1771 2499 1775
rect 2687 1771 2691 1775
rect 2879 1771 2883 1775
rect 3071 1771 3075 1775
rect 3263 1771 3267 1775
rect 3463 1771 3467 1775
rect 3663 1771 3667 1775
rect 3839 1771 3843 1775
rect 3943 1772 3947 1776
rect 111 1752 115 1756
rect 255 1751 259 1755
rect 391 1751 395 1755
rect 535 1751 539 1755
rect 695 1751 699 1755
rect 863 1751 867 1755
rect 1031 1751 1035 1755
rect 1207 1751 1211 1755
rect 1383 1751 1387 1755
rect 1559 1751 1563 1755
rect 1743 1751 1747 1755
rect 2007 1752 2011 1756
rect 2047 1755 2051 1759
rect 2127 1752 2131 1756
rect 2311 1752 2315 1756
rect 2495 1752 2499 1756
rect 2687 1752 2691 1756
rect 2879 1752 2883 1756
rect 3071 1752 3075 1756
rect 3263 1752 3267 1756
rect 3463 1752 3467 1756
rect 3663 1752 3667 1756
rect 3839 1752 3843 1756
rect 3943 1755 3947 1759
rect 111 1735 115 1739
rect 255 1732 259 1736
rect 391 1732 395 1736
rect 535 1732 539 1736
rect 695 1732 699 1736
rect 863 1732 867 1736
rect 1031 1732 1035 1736
rect 1207 1732 1211 1736
rect 1383 1732 1387 1736
rect 1559 1732 1563 1736
rect 1743 1732 1747 1736
rect 2007 1735 2011 1739
rect 2047 1685 2051 1689
rect 2071 1688 2075 1692
rect 2191 1688 2195 1692
rect 2343 1688 2347 1692
rect 2511 1688 2515 1692
rect 2687 1688 2691 1692
rect 2871 1688 2875 1692
rect 3063 1688 3067 1692
rect 3255 1688 3259 1692
rect 3447 1688 3451 1692
rect 3647 1688 3651 1692
rect 3839 1688 3843 1692
rect 3943 1685 3947 1689
rect 111 1669 115 1673
rect 135 1672 139 1676
rect 263 1672 267 1676
rect 431 1672 435 1676
rect 607 1672 611 1676
rect 799 1672 803 1676
rect 999 1672 1003 1676
rect 1199 1672 1203 1676
rect 1407 1672 1411 1676
rect 1623 1672 1627 1676
rect 1839 1672 1843 1676
rect 2007 1669 2011 1673
rect 2047 1668 2051 1672
rect 2071 1669 2075 1673
rect 2191 1669 2195 1673
rect 2343 1669 2347 1673
rect 2511 1669 2515 1673
rect 2687 1669 2691 1673
rect 2871 1669 2875 1673
rect 3063 1669 3067 1673
rect 3255 1669 3259 1673
rect 3447 1669 3451 1673
rect 3647 1669 3651 1673
rect 3839 1669 3843 1673
rect 3943 1668 3947 1672
rect 111 1652 115 1656
rect 135 1653 139 1657
rect 263 1653 267 1657
rect 431 1653 435 1657
rect 607 1653 611 1657
rect 799 1653 803 1657
rect 999 1653 1003 1657
rect 1199 1653 1203 1657
rect 1407 1653 1411 1657
rect 1623 1653 1627 1657
rect 1839 1653 1843 1657
rect 2007 1652 2011 1656
rect 2047 1616 2051 1620
rect 2071 1615 2075 1619
rect 2335 1615 2339 1619
rect 2599 1615 2603 1619
rect 2839 1615 2843 1619
rect 3047 1615 3051 1619
rect 3231 1615 3235 1619
rect 3399 1615 3403 1619
rect 3551 1615 3555 1619
rect 3695 1615 3699 1619
rect 3839 1615 3843 1619
rect 3943 1616 3947 1620
rect 111 1600 115 1604
rect 135 1599 139 1603
rect 287 1599 291 1603
rect 471 1599 475 1603
rect 655 1599 659 1603
rect 839 1599 843 1603
rect 1015 1599 1019 1603
rect 1183 1599 1187 1603
rect 1343 1599 1347 1603
rect 1495 1599 1499 1603
rect 1639 1599 1643 1603
rect 1783 1599 1787 1603
rect 1903 1599 1907 1603
rect 2007 1600 2011 1604
rect 2047 1599 2051 1603
rect 2071 1596 2075 1600
rect 2335 1596 2339 1600
rect 2599 1596 2603 1600
rect 2839 1596 2843 1600
rect 3047 1596 3051 1600
rect 3231 1596 3235 1600
rect 3399 1596 3403 1600
rect 3551 1596 3555 1600
rect 3695 1596 3699 1600
rect 3839 1596 3843 1600
rect 3943 1599 3947 1603
rect 111 1583 115 1587
rect 135 1580 139 1584
rect 287 1580 291 1584
rect 471 1580 475 1584
rect 655 1580 659 1584
rect 839 1580 843 1584
rect 1015 1580 1019 1584
rect 1183 1580 1187 1584
rect 1343 1580 1347 1584
rect 1495 1580 1499 1584
rect 1639 1580 1643 1584
rect 1783 1580 1787 1584
rect 1903 1580 1907 1584
rect 2007 1583 2011 1587
rect 2047 1529 2051 1533
rect 2583 1532 2587 1536
rect 2743 1532 2747 1536
rect 2903 1532 2907 1536
rect 3063 1532 3067 1536
rect 3223 1532 3227 1536
rect 3383 1532 3387 1536
rect 3543 1532 3547 1536
rect 3703 1532 3707 1536
rect 3943 1529 3947 1533
rect 111 1513 115 1517
rect 135 1516 139 1520
rect 295 1516 299 1520
rect 487 1516 491 1520
rect 687 1516 691 1520
rect 887 1516 891 1520
rect 1079 1516 1083 1520
rect 1263 1516 1267 1520
rect 1447 1516 1451 1520
rect 1623 1516 1627 1520
rect 1807 1516 1811 1520
rect 2007 1513 2011 1517
rect 2047 1512 2051 1516
rect 2583 1513 2587 1517
rect 2743 1513 2747 1517
rect 2903 1513 2907 1517
rect 3063 1513 3067 1517
rect 3223 1513 3227 1517
rect 3383 1513 3387 1517
rect 3543 1513 3547 1517
rect 3703 1513 3707 1517
rect 3943 1512 3947 1516
rect 111 1496 115 1500
rect 135 1497 139 1501
rect 295 1497 299 1501
rect 487 1497 491 1501
rect 687 1497 691 1501
rect 887 1497 891 1501
rect 1079 1497 1083 1501
rect 1263 1497 1267 1501
rect 1447 1497 1451 1501
rect 1623 1497 1627 1501
rect 1807 1497 1811 1501
rect 2007 1496 2011 1500
rect 2047 1460 2051 1464
rect 2415 1459 2419 1463
rect 2511 1459 2515 1463
rect 2607 1459 2611 1463
rect 2703 1459 2707 1463
rect 2799 1459 2803 1463
rect 2919 1459 2923 1463
rect 3063 1459 3067 1463
rect 3231 1459 3235 1463
rect 3415 1459 3419 1463
rect 3615 1459 3619 1463
rect 3815 1459 3819 1463
rect 3943 1460 3947 1464
rect 111 1444 115 1448
rect 175 1443 179 1447
rect 359 1443 363 1447
rect 567 1443 571 1447
rect 783 1443 787 1447
rect 1007 1443 1011 1447
rect 1231 1443 1235 1447
rect 1463 1443 1467 1447
rect 1695 1443 1699 1447
rect 1903 1443 1907 1447
rect 2007 1444 2011 1448
rect 2047 1443 2051 1447
rect 2415 1440 2419 1444
rect 2511 1440 2515 1444
rect 2607 1440 2611 1444
rect 2703 1440 2707 1444
rect 2799 1440 2803 1444
rect 2919 1440 2923 1444
rect 3063 1440 3067 1444
rect 3231 1440 3235 1444
rect 3415 1440 3419 1444
rect 3615 1440 3619 1444
rect 3815 1440 3819 1444
rect 3943 1443 3947 1447
rect 111 1427 115 1431
rect 175 1424 179 1428
rect 359 1424 363 1428
rect 567 1424 571 1428
rect 783 1424 787 1428
rect 1007 1424 1011 1428
rect 1231 1424 1235 1428
rect 1463 1424 1467 1428
rect 1695 1424 1699 1428
rect 1903 1424 1907 1428
rect 2007 1427 2011 1431
rect 111 1361 115 1365
rect 327 1364 331 1368
rect 463 1364 467 1368
rect 599 1364 603 1368
rect 727 1364 731 1368
rect 855 1364 859 1368
rect 983 1364 987 1368
rect 1119 1364 1123 1368
rect 1263 1364 1267 1368
rect 1423 1364 1427 1368
rect 1583 1364 1587 1368
rect 1751 1364 1755 1368
rect 1903 1364 1907 1368
rect 2007 1361 2011 1365
rect 2047 1357 2051 1361
rect 2071 1360 2075 1364
rect 2303 1360 2307 1364
rect 2559 1360 2563 1364
rect 2807 1360 2811 1364
rect 3055 1360 3059 1364
rect 3303 1360 3307 1364
rect 3559 1360 3563 1364
rect 3815 1360 3819 1364
rect 3943 1357 3947 1361
rect 111 1344 115 1348
rect 327 1345 331 1349
rect 463 1345 467 1349
rect 599 1345 603 1349
rect 727 1345 731 1349
rect 855 1345 859 1349
rect 983 1345 987 1349
rect 1119 1345 1123 1349
rect 1263 1345 1267 1349
rect 1423 1345 1427 1349
rect 1583 1345 1587 1349
rect 1751 1345 1755 1349
rect 1903 1345 1907 1349
rect 2007 1344 2011 1348
rect 2047 1340 2051 1344
rect 2071 1341 2075 1345
rect 2303 1341 2307 1345
rect 2559 1341 2563 1345
rect 2807 1341 2811 1345
rect 3055 1341 3059 1345
rect 3303 1341 3307 1345
rect 3559 1341 3563 1345
rect 3815 1341 3819 1345
rect 3943 1340 3947 1344
rect 111 1284 115 1288
rect 551 1283 555 1287
rect 655 1283 659 1287
rect 767 1283 771 1287
rect 879 1283 883 1287
rect 991 1283 995 1287
rect 1103 1283 1107 1287
rect 1215 1283 1219 1287
rect 1327 1283 1331 1287
rect 1439 1283 1443 1287
rect 1559 1283 1563 1287
rect 2007 1284 2011 1288
rect 2047 1280 2051 1284
rect 2071 1279 2075 1283
rect 2223 1279 2227 1283
rect 2415 1279 2419 1283
rect 2615 1279 2619 1283
rect 2815 1279 2819 1283
rect 2999 1279 3003 1283
rect 3175 1279 3179 1283
rect 3343 1279 3347 1283
rect 3503 1279 3507 1283
rect 3663 1279 3667 1283
rect 3831 1279 3835 1283
rect 3943 1280 3947 1284
rect 111 1267 115 1271
rect 551 1264 555 1268
rect 655 1264 659 1268
rect 767 1264 771 1268
rect 879 1264 883 1268
rect 991 1264 995 1268
rect 1103 1264 1107 1268
rect 1215 1264 1219 1268
rect 1327 1264 1331 1268
rect 1439 1264 1443 1268
rect 1559 1264 1563 1268
rect 2007 1267 2011 1271
rect 2047 1263 2051 1267
rect 2071 1260 2075 1264
rect 2223 1260 2227 1264
rect 2415 1260 2419 1264
rect 2615 1260 2619 1264
rect 2815 1260 2819 1264
rect 2999 1260 3003 1264
rect 3175 1260 3179 1264
rect 3343 1260 3347 1264
rect 3503 1260 3507 1264
rect 3663 1260 3667 1264
rect 3831 1260 3835 1264
rect 3943 1263 3947 1267
rect 111 1201 115 1205
rect 391 1204 395 1208
rect 519 1204 523 1208
rect 663 1204 667 1208
rect 807 1204 811 1208
rect 959 1204 963 1208
rect 1111 1204 1115 1208
rect 1255 1204 1259 1208
rect 1407 1204 1411 1208
rect 1559 1204 1563 1208
rect 1711 1204 1715 1208
rect 2007 1201 2011 1205
rect 111 1184 115 1188
rect 391 1185 395 1189
rect 519 1185 523 1189
rect 663 1185 667 1189
rect 807 1185 811 1189
rect 959 1185 963 1189
rect 1111 1185 1115 1189
rect 1255 1185 1259 1189
rect 1407 1185 1411 1189
rect 1559 1185 1563 1189
rect 2047 1189 2051 1193
rect 2135 1192 2139 1196
rect 2311 1192 2315 1196
rect 2503 1192 2507 1196
rect 2695 1192 2699 1196
rect 2887 1192 2891 1196
rect 3071 1192 3075 1196
rect 3239 1192 3243 1196
rect 3399 1192 3403 1196
rect 3551 1192 3555 1196
rect 3703 1192 3707 1196
rect 3839 1192 3843 1196
rect 1711 1185 1715 1189
rect 3943 1189 3947 1193
rect 2007 1184 2011 1188
rect 2047 1172 2051 1176
rect 2135 1173 2139 1177
rect 2311 1173 2315 1177
rect 2503 1173 2507 1177
rect 2695 1173 2699 1177
rect 2887 1173 2891 1177
rect 3071 1173 3075 1177
rect 3239 1173 3243 1177
rect 3399 1173 3403 1177
rect 3551 1173 3555 1177
rect 3703 1173 3707 1177
rect 3839 1173 3843 1177
rect 3943 1172 3947 1176
rect 111 1128 115 1132
rect 175 1127 179 1131
rect 327 1127 331 1131
rect 495 1127 499 1131
rect 671 1127 675 1131
rect 847 1127 851 1131
rect 1031 1127 1035 1131
rect 1207 1127 1211 1131
rect 1383 1127 1387 1131
rect 1567 1127 1571 1131
rect 1751 1127 1755 1131
rect 2007 1128 2011 1132
rect 111 1111 115 1115
rect 175 1108 179 1112
rect 327 1108 331 1112
rect 495 1108 499 1112
rect 671 1108 675 1112
rect 847 1108 851 1112
rect 1031 1108 1035 1112
rect 1207 1108 1211 1112
rect 1383 1108 1387 1112
rect 1567 1108 1571 1112
rect 1751 1108 1755 1112
rect 2007 1111 2011 1115
rect 2047 1112 2051 1116
rect 2295 1111 2299 1115
rect 2423 1111 2427 1115
rect 2559 1111 2563 1115
rect 2695 1111 2699 1115
rect 2839 1111 2843 1115
rect 2991 1111 2995 1115
rect 3151 1111 3155 1115
rect 3319 1111 3323 1115
rect 3495 1111 3499 1115
rect 3679 1111 3683 1115
rect 3839 1111 3843 1115
rect 3943 1112 3947 1116
rect 2047 1095 2051 1099
rect 2295 1092 2299 1096
rect 2423 1092 2427 1096
rect 2559 1092 2563 1096
rect 2695 1092 2699 1096
rect 2839 1092 2843 1096
rect 2991 1092 2995 1096
rect 3151 1092 3155 1096
rect 3319 1092 3323 1096
rect 3495 1092 3499 1096
rect 3679 1092 3683 1096
rect 3839 1092 3843 1096
rect 3943 1095 3947 1099
rect 111 1037 115 1041
rect 135 1040 139 1044
rect 231 1040 235 1044
rect 375 1040 379 1044
rect 543 1040 547 1044
rect 727 1040 731 1044
rect 911 1040 915 1044
rect 1095 1040 1099 1044
rect 1279 1040 1283 1044
rect 1463 1040 1467 1044
rect 1647 1040 1651 1044
rect 1831 1040 1835 1044
rect 2007 1037 2011 1041
rect 111 1020 115 1024
rect 135 1021 139 1025
rect 231 1021 235 1025
rect 375 1021 379 1025
rect 543 1021 547 1025
rect 727 1021 731 1025
rect 911 1021 915 1025
rect 1095 1021 1099 1025
rect 1279 1021 1283 1025
rect 1463 1021 1467 1025
rect 1647 1021 1651 1025
rect 2047 1025 2051 1029
rect 2495 1028 2499 1032
rect 2599 1028 2603 1032
rect 2711 1028 2715 1032
rect 2847 1028 2851 1032
rect 3007 1028 3011 1032
rect 3199 1028 3203 1032
rect 3407 1028 3411 1032
rect 3631 1028 3635 1032
rect 3839 1028 3843 1032
rect 1831 1021 1835 1025
rect 3943 1025 3947 1029
rect 2007 1020 2011 1024
rect 2047 1008 2051 1012
rect 2495 1009 2499 1013
rect 2599 1009 2603 1013
rect 2711 1009 2715 1013
rect 2847 1009 2851 1013
rect 3007 1009 3011 1013
rect 3199 1009 3203 1013
rect 3407 1009 3411 1013
rect 3631 1009 3635 1013
rect 3839 1009 3843 1013
rect 3943 1008 3947 1012
rect 111 968 115 972
rect 135 967 139 971
rect 271 967 275 971
rect 447 967 451 971
rect 631 967 635 971
rect 823 967 827 971
rect 1007 967 1011 971
rect 1175 967 1179 971
rect 1335 967 1339 971
rect 1487 967 1491 971
rect 1631 967 1635 971
rect 1775 967 1779 971
rect 1903 967 1907 971
rect 2007 968 2011 972
rect 2047 956 2051 960
rect 111 951 115 955
rect 2647 955 2651 959
rect 135 948 139 952
rect 271 948 275 952
rect 447 948 451 952
rect 631 948 635 952
rect 823 948 827 952
rect 1007 948 1011 952
rect 1175 948 1179 952
rect 1335 948 1339 952
rect 1487 948 1491 952
rect 1631 948 1635 952
rect 1775 948 1779 952
rect 1903 948 1907 952
rect 2007 951 2011 955
rect 2743 955 2747 959
rect 2847 955 2851 959
rect 2967 955 2971 959
rect 3111 955 3115 959
rect 3279 955 3283 959
rect 3463 955 3467 959
rect 3663 955 3667 959
rect 3839 955 3843 959
rect 3943 956 3947 960
rect 2047 939 2051 943
rect 2647 936 2651 940
rect 2743 936 2747 940
rect 2847 936 2851 940
rect 2967 936 2971 940
rect 3111 936 3115 940
rect 3279 936 3283 940
rect 3463 936 3467 940
rect 3663 936 3667 940
rect 3839 936 3843 940
rect 3943 939 3947 943
rect 111 885 115 889
rect 135 888 139 892
rect 271 888 275 892
rect 455 888 459 892
rect 655 888 659 892
rect 855 888 859 892
rect 1055 888 1059 892
rect 1239 888 1243 892
rect 1415 888 1419 892
rect 1583 888 1587 892
rect 1751 888 1755 892
rect 1903 888 1907 892
rect 2007 885 2011 889
rect 111 868 115 872
rect 135 869 139 873
rect 271 869 275 873
rect 455 869 459 873
rect 655 869 659 873
rect 855 869 859 873
rect 1055 869 1059 873
rect 1239 869 1243 873
rect 1415 869 1419 873
rect 1583 869 1587 873
rect 1751 869 1755 873
rect 1903 869 1907 873
rect 2007 868 2011 872
rect 2047 861 2051 865
rect 2071 864 2075 868
rect 2255 864 2259 868
rect 2463 864 2467 868
rect 2679 864 2683 868
rect 2895 864 2899 868
rect 3127 864 3131 868
rect 3367 864 3371 868
rect 3615 864 3619 868
rect 3839 864 3843 868
rect 3943 861 3947 865
rect 2047 844 2051 848
rect 2071 845 2075 849
rect 2255 845 2259 849
rect 2463 845 2467 849
rect 2679 845 2683 849
rect 2895 845 2899 849
rect 3127 845 3131 849
rect 3367 845 3371 849
rect 3615 845 3619 849
rect 3839 845 3843 849
rect 3943 844 3947 848
rect 111 816 115 820
rect 215 815 219 819
rect 343 815 347 819
rect 495 815 499 819
rect 655 815 659 819
rect 831 815 835 819
rect 1007 815 1011 819
rect 1183 815 1187 819
rect 1359 815 1363 819
rect 1535 815 1539 819
rect 1719 815 1723 819
rect 2007 816 2011 820
rect 111 799 115 803
rect 215 796 219 800
rect 343 796 347 800
rect 495 796 499 800
rect 655 796 659 800
rect 831 796 835 800
rect 1007 796 1011 800
rect 1183 796 1187 800
rect 1359 796 1363 800
rect 1535 796 1539 800
rect 1719 796 1723 800
rect 2007 799 2011 803
rect 2047 792 2051 796
rect 2215 791 2219 795
rect 2327 791 2331 795
rect 2447 791 2451 795
rect 2583 791 2587 795
rect 2735 791 2739 795
rect 2895 791 2899 795
rect 3063 791 3067 795
rect 3247 791 3251 795
rect 3447 791 3451 795
rect 3655 791 3659 795
rect 3839 791 3843 795
rect 3943 792 3947 796
rect 2047 775 2051 779
rect 2215 772 2219 776
rect 2327 772 2331 776
rect 2447 772 2451 776
rect 2583 772 2587 776
rect 2735 772 2739 776
rect 2895 772 2899 776
rect 3063 772 3067 776
rect 3247 772 3251 776
rect 3447 772 3451 776
rect 3655 772 3659 776
rect 3839 772 3843 776
rect 3943 775 3947 779
rect 111 733 115 737
rect 375 736 379 740
rect 495 736 499 740
rect 623 736 627 740
rect 751 736 755 740
rect 887 736 891 740
rect 1023 736 1027 740
rect 1167 736 1171 740
rect 1311 736 1315 740
rect 1455 736 1459 740
rect 1599 736 1603 740
rect 2007 733 2011 737
rect 111 716 115 720
rect 375 717 379 721
rect 495 717 499 721
rect 623 717 627 721
rect 751 717 755 721
rect 887 717 891 721
rect 1023 717 1027 721
rect 1167 717 1171 721
rect 1311 717 1315 721
rect 1455 717 1459 721
rect 1599 717 1603 721
rect 2007 716 2011 720
rect 2047 705 2051 709
rect 2375 708 2379 712
rect 2495 708 2499 712
rect 2623 708 2627 712
rect 2767 708 2771 712
rect 2911 708 2915 712
rect 3063 708 3067 712
rect 3215 708 3219 712
rect 3367 708 3371 712
rect 3519 708 3523 712
rect 3679 708 3683 712
rect 3839 708 3843 712
rect 3943 705 3947 709
rect 2047 688 2051 692
rect 2375 689 2379 693
rect 2495 689 2499 693
rect 2623 689 2627 693
rect 2767 689 2771 693
rect 2911 689 2915 693
rect 3063 689 3067 693
rect 3215 689 3219 693
rect 3367 689 3371 693
rect 3519 689 3523 693
rect 3679 689 3683 693
rect 3839 689 3843 693
rect 3943 688 3947 692
rect 111 664 115 668
rect 527 663 531 667
rect 631 663 635 667
rect 743 663 747 667
rect 855 663 859 667
rect 967 663 971 667
rect 1071 663 1075 667
rect 1183 663 1187 667
rect 1295 663 1299 667
rect 1407 663 1411 667
rect 1519 663 1523 667
rect 2007 664 2011 668
rect 111 647 115 651
rect 527 644 531 648
rect 631 644 635 648
rect 743 644 747 648
rect 855 644 859 648
rect 967 644 971 648
rect 1071 644 1075 648
rect 1183 644 1187 648
rect 1295 644 1299 648
rect 1407 644 1411 648
rect 1519 644 1523 648
rect 2007 647 2011 651
rect 2047 628 2051 632
rect 2111 627 2115 631
rect 2247 627 2251 631
rect 2399 627 2403 631
rect 2575 627 2579 631
rect 2759 627 2763 631
rect 2943 627 2947 631
rect 3127 627 3131 631
rect 3303 627 3307 631
rect 3479 627 3483 631
rect 3655 627 3659 631
rect 3831 627 3835 631
rect 3943 628 3947 632
rect 2047 611 2051 615
rect 2111 608 2115 612
rect 2247 608 2251 612
rect 2399 608 2403 612
rect 2575 608 2579 612
rect 2759 608 2763 612
rect 2943 608 2947 612
rect 3127 608 3131 612
rect 3303 608 3307 612
rect 3479 608 3483 612
rect 3655 608 3659 612
rect 3831 608 3835 612
rect 3943 611 3947 615
rect 111 581 115 585
rect 687 584 691 588
rect 783 584 787 588
rect 879 584 883 588
rect 975 584 979 588
rect 1071 584 1075 588
rect 1167 584 1171 588
rect 1263 584 1267 588
rect 1359 584 1363 588
rect 1455 584 1459 588
rect 2007 581 2011 585
rect 111 564 115 568
rect 687 565 691 569
rect 783 565 787 569
rect 879 565 883 569
rect 975 565 979 569
rect 1071 565 1075 569
rect 1167 565 1171 569
rect 1263 565 1267 569
rect 1359 565 1363 569
rect 1455 565 1459 569
rect 2007 564 2011 568
rect 2047 541 2051 545
rect 2071 544 2075 548
rect 2183 544 2187 548
rect 2335 544 2339 548
rect 2503 544 2507 548
rect 2687 544 2691 548
rect 2879 544 2883 548
rect 3071 544 3075 548
rect 3263 544 3267 548
rect 3455 544 3459 548
rect 3647 544 3651 548
rect 3839 544 3843 548
rect 3943 541 3947 545
rect 2047 524 2051 528
rect 2071 525 2075 529
rect 2183 525 2187 529
rect 2335 525 2339 529
rect 2503 525 2507 529
rect 2687 525 2691 529
rect 2879 525 2883 529
rect 3071 525 3075 529
rect 3263 525 3267 529
rect 3455 525 3459 529
rect 3647 525 3651 529
rect 3839 525 3843 529
rect 3943 524 3947 528
rect 111 492 115 496
rect 383 491 387 495
rect 479 491 483 495
rect 575 491 579 495
rect 671 491 675 495
rect 767 491 771 495
rect 863 491 867 495
rect 959 491 963 495
rect 1055 491 1059 495
rect 1151 491 1155 495
rect 1247 491 1251 495
rect 1343 491 1347 495
rect 1439 491 1443 495
rect 1535 491 1539 495
rect 2007 492 2011 496
rect 111 475 115 479
rect 383 472 387 476
rect 479 472 483 476
rect 575 472 579 476
rect 671 472 675 476
rect 767 472 771 476
rect 863 472 867 476
rect 959 472 963 476
rect 1055 472 1059 476
rect 1151 472 1155 476
rect 1247 472 1251 476
rect 1343 472 1347 476
rect 1439 472 1443 476
rect 1535 472 1539 476
rect 2007 475 2011 479
rect 2047 472 2051 476
rect 2183 471 2187 475
rect 2319 471 2323 475
rect 2463 471 2467 475
rect 2615 471 2619 475
rect 2775 471 2779 475
rect 2959 471 2963 475
rect 3159 471 3163 475
rect 3367 471 3371 475
rect 3583 471 3587 475
rect 3807 471 3811 475
rect 3943 472 3947 476
rect 2047 455 2051 459
rect 2183 452 2187 456
rect 2319 452 2323 456
rect 2463 452 2467 456
rect 2615 452 2619 456
rect 2775 452 2779 456
rect 2959 452 2963 456
rect 3159 452 3163 456
rect 3367 452 3371 456
rect 3583 452 3587 456
rect 3807 452 3811 456
rect 3943 455 3947 459
rect 111 397 115 401
rect 487 400 491 404
rect 583 400 587 404
rect 687 400 691 404
rect 791 400 795 404
rect 895 400 899 404
rect 999 400 1003 404
rect 1103 400 1107 404
rect 1207 400 1211 404
rect 1319 400 1323 404
rect 1431 400 1435 404
rect 2007 397 2011 401
rect 2047 389 2051 393
rect 2343 392 2347 396
rect 2487 392 2491 396
rect 2639 392 2643 396
rect 2799 392 2803 396
rect 2959 392 2963 396
rect 3111 392 3115 396
rect 3263 392 3267 396
rect 3415 392 3419 396
rect 3559 392 3563 396
rect 3711 392 3715 396
rect 3839 392 3843 396
rect 3943 389 3947 393
rect 111 380 115 384
rect 487 381 491 385
rect 583 381 587 385
rect 687 381 691 385
rect 791 381 795 385
rect 895 381 899 385
rect 999 381 1003 385
rect 1103 381 1107 385
rect 1207 381 1211 385
rect 1319 381 1323 385
rect 1431 381 1435 385
rect 2007 380 2011 384
rect 2047 372 2051 376
rect 2343 373 2347 377
rect 2487 373 2491 377
rect 2639 373 2643 377
rect 2799 373 2803 377
rect 2959 373 2963 377
rect 3111 373 3115 377
rect 3263 373 3267 377
rect 3415 373 3419 377
rect 3559 373 3563 377
rect 3711 373 3715 377
rect 3839 373 3843 377
rect 3943 372 3947 376
rect 111 324 115 328
rect 327 323 331 327
rect 463 323 467 327
rect 615 323 619 327
rect 767 323 771 327
rect 919 323 923 327
rect 1063 323 1067 327
rect 1207 323 1211 327
rect 1351 323 1355 327
rect 1495 323 1499 327
rect 1639 323 1643 327
rect 2007 324 2011 328
rect 2047 316 2051 320
rect 2495 315 2499 319
rect 2639 315 2643 319
rect 2799 315 2803 319
rect 2959 315 2963 319
rect 3119 315 3123 319
rect 3271 315 3275 319
rect 3423 315 3427 319
rect 3567 315 3571 319
rect 3711 315 3715 319
rect 3839 315 3843 319
rect 3943 316 3947 320
rect 111 307 115 311
rect 327 304 331 308
rect 463 304 467 308
rect 615 304 619 308
rect 767 304 771 308
rect 919 304 923 308
rect 1063 304 1067 308
rect 1207 304 1211 308
rect 1351 304 1355 308
rect 1495 304 1499 308
rect 1639 304 1643 308
rect 2007 307 2011 311
rect 2047 299 2051 303
rect 2495 296 2499 300
rect 2639 296 2643 300
rect 2799 296 2803 300
rect 2959 296 2963 300
rect 3119 296 3123 300
rect 3271 296 3275 300
rect 3423 296 3427 300
rect 3567 296 3571 300
rect 3711 296 3715 300
rect 3839 296 3843 300
rect 3943 299 3947 303
rect 111 233 115 237
rect 167 236 171 240
rect 327 236 331 240
rect 503 236 507 240
rect 687 236 691 240
rect 871 236 875 240
rect 1047 236 1051 240
rect 1215 236 1219 240
rect 1367 236 1371 240
rect 1511 236 1515 240
rect 1647 236 1651 240
rect 1783 236 1787 240
rect 1903 236 1907 240
rect 2007 233 2011 237
rect 2047 233 2051 237
rect 2071 236 2075 240
rect 2271 236 2275 240
rect 2495 236 2499 240
rect 2703 236 2707 240
rect 2903 236 2907 240
rect 3095 236 3099 240
rect 3287 236 3291 240
rect 3479 236 3483 240
rect 3671 236 3675 240
rect 3839 236 3843 240
rect 3943 233 3947 237
rect 111 216 115 220
rect 167 217 171 221
rect 327 217 331 221
rect 503 217 507 221
rect 687 217 691 221
rect 871 217 875 221
rect 1047 217 1051 221
rect 1215 217 1219 221
rect 1367 217 1371 221
rect 1511 217 1515 221
rect 1647 217 1651 221
rect 1783 217 1787 221
rect 1903 217 1907 221
rect 2007 216 2011 220
rect 2047 216 2051 220
rect 2071 217 2075 221
rect 2271 217 2275 221
rect 2495 217 2499 221
rect 2703 217 2707 221
rect 2903 217 2907 221
rect 3095 217 3099 221
rect 3287 217 3291 221
rect 3479 217 3483 221
rect 3671 217 3675 221
rect 3839 217 3843 221
rect 3943 216 3947 220
rect 111 136 115 140
rect 135 135 139 139
rect 231 135 235 139
rect 327 135 331 139
rect 423 135 427 139
rect 527 135 531 139
rect 647 135 651 139
rect 775 135 779 139
rect 903 135 907 139
rect 1031 135 1035 139
rect 1151 135 1155 139
rect 1271 135 1275 139
rect 1383 135 1387 139
rect 1487 135 1491 139
rect 1591 135 1595 139
rect 1703 135 1707 139
rect 1807 135 1811 139
rect 1903 135 1907 139
rect 2007 136 2011 140
rect 2047 140 2051 144
rect 2071 139 2075 143
rect 2167 139 2171 143
rect 2263 139 2267 143
rect 2359 139 2363 143
rect 2455 139 2459 143
rect 2551 139 2555 143
rect 2655 139 2659 143
rect 2759 139 2763 143
rect 2863 139 2867 143
rect 2975 139 2979 143
rect 3103 139 3107 143
rect 3239 139 3243 143
rect 3383 139 3387 143
rect 3535 139 3539 143
rect 3695 139 3699 143
rect 3839 139 3843 143
rect 3943 140 3947 144
rect 111 119 115 123
rect 135 116 139 120
rect 231 116 235 120
rect 327 116 331 120
rect 423 116 427 120
rect 527 116 531 120
rect 647 116 651 120
rect 775 116 779 120
rect 903 116 907 120
rect 1031 116 1035 120
rect 1151 116 1155 120
rect 1271 116 1275 120
rect 1383 116 1387 120
rect 1487 116 1491 120
rect 1591 116 1595 120
rect 1703 116 1707 120
rect 1807 116 1811 120
rect 1903 116 1907 120
rect 2007 119 2011 123
rect 2047 123 2051 127
rect 2071 120 2075 124
rect 2167 120 2171 124
rect 2263 120 2267 124
rect 2359 120 2363 124
rect 2455 120 2459 124
rect 2551 120 2555 124
rect 2655 120 2659 124
rect 2759 120 2763 124
rect 2863 120 2867 124
rect 2975 120 2979 124
rect 3103 120 3107 124
rect 3239 120 3243 124
rect 3383 120 3387 124
rect 3535 120 3539 124
rect 3695 120 3699 124
rect 3839 120 3843 124
rect 3943 123 3947 127
<< m3 >>
rect 111 4030 115 4031
rect 111 4025 115 4026
rect 1519 4030 1523 4031
rect 1519 4025 1523 4026
rect 1615 4030 1619 4031
rect 1615 4025 1619 4026
rect 1711 4030 1715 4031
rect 1711 4025 1715 4026
rect 1807 4030 1811 4031
rect 1807 4025 1811 4026
rect 1903 4030 1907 4031
rect 1903 4025 1907 4026
rect 2007 4030 2011 4031
rect 2007 4025 2011 4026
rect 112 4005 114 4025
rect 110 4004 116 4005
rect 1520 4004 1522 4025
rect 1616 4004 1618 4025
rect 1712 4004 1714 4025
rect 1808 4004 1810 4025
rect 1904 4004 1906 4025
rect 2008 4005 2010 4025
rect 2047 4018 2051 4019
rect 2047 4013 2051 4014
rect 2071 4018 2075 4019
rect 2071 4013 2075 4014
rect 2167 4018 2171 4019
rect 2167 4013 2171 4014
rect 2263 4018 2267 4019
rect 2263 4013 2267 4014
rect 3943 4018 3947 4019
rect 3943 4013 3947 4014
rect 2006 4004 2012 4005
rect 110 4000 111 4004
rect 115 4000 116 4004
rect 110 3999 116 4000
rect 1518 4003 1524 4004
rect 1518 3999 1519 4003
rect 1523 3999 1524 4003
rect 1518 3998 1524 3999
rect 1614 4003 1620 4004
rect 1614 3999 1615 4003
rect 1619 3999 1620 4003
rect 1614 3998 1620 3999
rect 1710 4003 1716 4004
rect 1710 3999 1711 4003
rect 1715 3999 1716 4003
rect 1710 3998 1716 3999
rect 1806 4003 1812 4004
rect 1806 3999 1807 4003
rect 1811 3999 1812 4003
rect 1806 3998 1812 3999
rect 1902 4003 1908 4004
rect 1902 3999 1903 4003
rect 1907 3999 1908 4003
rect 2006 4000 2007 4004
rect 2011 4000 2012 4004
rect 2006 3999 2012 4000
rect 1902 3998 1908 3999
rect 110 3987 116 3988
rect 110 3983 111 3987
rect 115 3983 116 3987
rect 2006 3987 2012 3988
rect 110 3982 116 3983
rect 1518 3984 1524 3985
rect 112 3955 114 3982
rect 1518 3980 1519 3984
rect 1523 3980 1524 3984
rect 1518 3979 1524 3980
rect 1614 3984 1620 3985
rect 1614 3980 1615 3984
rect 1619 3980 1620 3984
rect 1614 3979 1620 3980
rect 1710 3984 1716 3985
rect 1710 3980 1711 3984
rect 1715 3980 1716 3984
rect 1710 3979 1716 3980
rect 1806 3984 1812 3985
rect 1806 3980 1807 3984
rect 1811 3980 1812 3984
rect 1806 3979 1812 3980
rect 1902 3984 1908 3985
rect 1902 3980 1903 3984
rect 1907 3980 1908 3984
rect 2006 3983 2007 3987
rect 2011 3983 2012 3987
rect 2048 3986 2050 4013
rect 2072 3989 2074 4013
rect 2168 3989 2170 4013
rect 2264 3989 2266 4013
rect 2070 3988 2076 3989
rect 2006 3982 2012 3983
rect 2046 3985 2052 3986
rect 1902 3979 1908 3980
rect 1520 3955 1522 3979
rect 1616 3955 1618 3979
rect 1712 3955 1714 3979
rect 1808 3955 1810 3979
rect 1904 3955 1906 3979
rect 2008 3955 2010 3982
rect 2046 3981 2047 3985
rect 2051 3981 2052 3985
rect 2070 3984 2071 3988
rect 2075 3984 2076 3988
rect 2070 3983 2076 3984
rect 2166 3988 2172 3989
rect 2166 3984 2167 3988
rect 2171 3984 2172 3988
rect 2166 3983 2172 3984
rect 2262 3988 2268 3989
rect 2262 3984 2263 3988
rect 2267 3984 2268 3988
rect 3944 3986 3946 4013
rect 2262 3983 2268 3984
rect 3942 3985 3948 3986
rect 2046 3980 2052 3981
rect 3942 3981 3943 3985
rect 3947 3981 3948 3985
rect 3942 3980 3948 3981
rect 2070 3969 2076 3970
rect 2046 3968 2052 3969
rect 2046 3964 2047 3968
rect 2051 3964 2052 3968
rect 2070 3965 2071 3969
rect 2075 3965 2076 3969
rect 2070 3964 2076 3965
rect 2166 3969 2172 3970
rect 2166 3965 2167 3969
rect 2171 3965 2172 3969
rect 2166 3964 2172 3965
rect 2262 3969 2268 3970
rect 2262 3965 2263 3969
rect 2267 3965 2268 3969
rect 2262 3964 2268 3965
rect 3942 3968 3948 3969
rect 3942 3964 3943 3968
rect 3947 3964 3948 3968
rect 2046 3963 2052 3964
rect 111 3954 115 3955
rect 111 3949 115 3950
rect 199 3954 203 3955
rect 199 3949 203 3950
rect 295 3954 299 3955
rect 295 3949 299 3950
rect 391 3954 395 3955
rect 391 3949 395 3950
rect 495 3954 499 3955
rect 495 3949 499 3950
rect 615 3954 619 3955
rect 615 3949 619 3950
rect 743 3954 747 3955
rect 743 3949 747 3950
rect 871 3954 875 3955
rect 871 3949 875 3950
rect 999 3954 1003 3955
rect 999 3949 1003 3950
rect 1127 3954 1131 3955
rect 1127 3949 1131 3950
rect 1255 3954 1259 3955
rect 1255 3949 1259 3950
rect 1383 3954 1387 3955
rect 1383 3949 1387 3950
rect 1511 3954 1515 3955
rect 1511 3949 1515 3950
rect 1519 3954 1523 3955
rect 1519 3949 1523 3950
rect 1615 3954 1619 3955
rect 1615 3949 1619 3950
rect 1647 3954 1651 3955
rect 1647 3949 1651 3950
rect 1711 3954 1715 3955
rect 1711 3949 1715 3950
rect 1807 3954 1811 3955
rect 1807 3949 1811 3950
rect 1903 3954 1907 3955
rect 1903 3949 1907 3950
rect 2007 3954 2011 3955
rect 2007 3949 2011 3950
rect 112 3922 114 3949
rect 200 3925 202 3949
rect 296 3925 298 3949
rect 392 3925 394 3949
rect 496 3925 498 3949
rect 616 3925 618 3949
rect 744 3925 746 3949
rect 872 3925 874 3949
rect 1000 3925 1002 3949
rect 1128 3925 1130 3949
rect 1256 3925 1258 3949
rect 1384 3925 1386 3949
rect 1512 3925 1514 3949
rect 1648 3925 1650 3949
rect 198 3924 204 3925
rect 110 3921 116 3922
rect 110 3917 111 3921
rect 115 3917 116 3921
rect 198 3920 199 3924
rect 203 3920 204 3924
rect 198 3919 204 3920
rect 294 3924 300 3925
rect 294 3920 295 3924
rect 299 3920 300 3924
rect 294 3919 300 3920
rect 390 3924 396 3925
rect 390 3920 391 3924
rect 395 3920 396 3924
rect 390 3919 396 3920
rect 494 3924 500 3925
rect 494 3920 495 3924
rect 499 3920 500 3924
rect 494 3919 500 3920
rect 614 3924 620 3925
rect 614 3920 615 3924
rect 619 3920 620 3924
rect 614 3919 620 3920
rect 742 3924 748 3925
rect 742 3920 743 3924
rect 747 3920 748 3924
rect 742 3919 748 3920
rect 870 3924 876 3925
rect 870 3920 871 3924
rect 875 3920 876 3924
rect 870 3919 876 3920
rect 998 3924 1004 3925
rect 998 3920 999 3924
rect 1003 3920 1004 3924
rect 998 3919 1004 3920
rect 1126 3924 1132 3925
rect 1126 3920 1127 3924
rect 1131 3920 1132 3924
rect 1126 3919 1132 3920
rect 1254 3924 1260 3925
rect 1254 3920 1255 3924
rect 1259 3920 1260 3924
rect 1254 3919 1260 3920
rect 1382 3924 1388 3925
rect 1382 3920 1383 3924
rect 1387 3920 1388 3924
rect 1382 3919 1388 3920
rect 1510 3924 1516 3925
rect 1510 3920 1511 3924
rect 1515 3920 1516 3924
rect 1510 3919 1516 3920
rect 1646 3924 1652 3925
rect 1646 3920 1647 3924
rect 1651 3920 1652 3924
rect 2008 3922 2010 3949
rect 2048 3943 2050 3963
rect 2072 3943 2074 3964
rect 2168 3943 2170 3964
rect 2264 3943 2266 3964
rect 3942 3963 3948 3964
rect 3944 3943 3946 3963
rect 2047 3942 2051 3943
rect 2047 3937 2051 3938
rect 2071 3942 2075 3943
rect 2071 3937 2075 3938
rect 2159 3942 2163 3943
rect 2159 3937 2163 3938
rect 2167 3942 2171 3943
rect 2167 3937 2171 3938
rect 2263 3942 2267 3943
rect 2263 3937 2267 3938
rect 2287 3942 2291 3943
rect 2287 3937 2291 3938
rect 2415 3942 2419 3943
rect 2415 3937 2419 3938
rect 2551 3942 2555 3943
rect 2551 3937 2555 3938
rect 2687 3942 2691 3943
rect 2687 3937 2691 3938
rect 2823 3942 2827 3943
rect 2823 3937 2827 3938
rect 2951 3942 2955 3943
rect 2951 3937 2955 3938
rect 3071 3942 3075 3943
rect 3071 3937 3075 3938
rect 3191 3942 3195 3943
rect 3191 3937 3195 3938
rect 3303 3942 3307 3943
rect 3303 3937 3307 3938
rect 3407 3942 3411 3943
rect 3407 3937 3411 3938
rect 3519 3942 3523 3943
rect 3519 3937 3523 3938
rect 3631 3942 3635 3943
rect 3631 3937 3635 3938
rect 3743 3942 3747 3943
rect 3743 3937 3747 3938
rect 3943 3942 3947 3943
rect 3943 3937 3947 3938
rect 1646 3919 1652 3920
rect 2006 3921 2012 3922
rect 110 3916 116 3917
rect 2006 3917 2007 3921
rect 2011 3917 2012 3921
rect 2048 3917 2050 3937
rect 2006 3916 2012 3917
rect 2046 3916 2052 3917
rect 2160 3916 2162 3937
rect 2288 3916 2290 3937
rect 2416 3916 2418 3937
rect 2552 3916 2554 3937
rect 2688 3916 2690 3937
rect 2824 3916 2826 3937
rect 2952 3916 2954 3937
rect 3072 3916 3074 3937
rect 3192 3916 3194 3937
rect 3304 3916 3306 3937
rect 3408 3916 3410 3937
rect 3520 3916 3522 3937
rect 3632 3916 3634 3937
rect 3744 3916 3746 3937
rect 3944 3917 3946 3937
rect 3942 3916 3948 3917
rect 2046 3912 2047 3916
rect 2051 3912 2052 3916
rect 2046 3911 2052 3912
rect 2158 3915 2164 3916
rect 2158 3911 2159 3915
rect 2163 3911 2164 3915
rect 2158 3910 2164 3911
rect 2286 3915 2292 3916
rect 2286 3911 2287 3915
rect 2291 3911 2292 3915
rect 2286 3910 2292 3911
rect 2414 3915 2420 3916
rect 2414 3911 2415 3915
rect 2419 3911 2420 3915
rect 2414 3910 2420 3911
rect 2550 3915 2556 3916
rect 2550 3911 2551 3915
rect 2555 3911 2556 3915
rect 2550 3910 2556 3911
rect 2686 3915 2692 3916
rect 2686 3911 2687 3915
rect 2691 3911 2692 3915
rect 2686 3910 2692 3911
rect 2822 3915 2828 3916
rect 2822 3911 2823 3915
rect 2827 3911 2828 3915
rect 2822 3910 2828 3911
rect 2950 3915 2956 3916
rect 2950 3911 2951 3915
rect 2955 3911 2956 3915
rect 2950 3910 2956 3911
rect 3070 3915 3076 3916
rect 3070 3911 3071 3915
rect 3075 3911 3076 3915
rect 3070 3910 3076 3911
rect 3190 3915 3196 3916
rect 3190 3911 3191 3915
rect 3195 3911 3196 3915
rect 3190 3910 3196 3911
rect 3302 3915 3308 3916
rect 3302 3911 3303 3915
rect 3307 3911 3308 3915
rect 3302 3910 3308 3911
rect 3406 3915 3412 3916
rect 3406 3911 3407 3915
rect 3411 3911 3412 3915
rect 3406 3910 3412 3911
rect 3518 3915 3524 3916
rect 3518 3911 3519 3915
rect 3523 3911 3524 3915
rect 3518 3910 3524 3911
rect 3630 3915 3636 3916
rect 3630 3911 3631 3915
rect 3635 3911 3636 3915
rect 3630 3910 3636 3911
rect 3742 3915 3748 3916
rect 3742 3911 3743 3915
rect 3747 3911 3748 3915
rect 3942 3912 3943 3916
rect 3947 3912 3948 3916
rect 3942 3911 3948 3912
rect 3742 3910 3748 3911
rect 198 3905 204 3906
rect 110 3904 116 3905
rect 110 3900 111 3904
rect 115 3900 116 3904
rect 198 3901 199 3905
rect 203 3901 204 3905
rect 198 3900 204 3901
rect 294 3905 300 3906
rect 294 3901 295 3905
rect 299 3901 300 3905
rect 294 3900 300 3901
rect 390 3905 396 3906
rect 390 3901 391 3905
rect 395 3901 396 3905
rect 390 3900 396 3901
rect 494 3905 500 3906
rect 494 3901 495 3905
rect 499 3901 500 3905
rect 494 3900 500 3901
rect 614 3905 620 3906
rect 614 3901 615 3905
rect 619 3901 620 3905
rect 614 3900 620 3901
rect 742 3905 748 3906
rect 742 3901 743 3905
rect 747 3901 748 3905
rect 742 3900 748 3901
rect 870 3905 876 3906
rect 870 3901 871 3905
rect 875 3901 876 3905
rect 870 3900 876 3901
rect 998 3905 1004 3906
rect 998 3901 999 3905
rect 1003 3901 1004 3905
rect 998 3900 1004 3901
rect 1126 3905 1132 3906
rect 1126 3901 1127 3905
rect 1131 3901 1132 3905
rect 1126 3900 1132 3901
rect 1254 3905 1260 3906
rect 1254 3901 1255 3905
rect 1259 3901 1260 3905
rect 1254 3900 1260 3901
rect 1382 3905 1388 3906
rect 1382 3901 1383 3905
rect 1387 3901 1388 3905
rect 1382 3900 1388 3901
rect 1510 3905 1516 3906
rect 1510 3901 1511 3905
rect 1515 3901 1516 3905
rect 1510 3900 1516 3901
rect 1646 3905 1652 3906
rect 1646 3901 1647 3905
rect 1651 3901 1652 3905
rect 1646 3900 1652 3901
rect 2006 3904 2012 3905
rect 2006 3900 2007 3904
rect 2011 3900 2012 3904
rect 110 3899 116 3900
rect 112 3879 114 3899
rect 200 3879 202 3900
rect 296 3879 298 3900
rect 392 3879 394 3900
rect 496 3879 498 3900
rect 616 3879 618 3900
rect 744 3879 746 3900
rect 872 3879 874 3900
rect 1000 3879 1002 3900
rect 1128 3879 1130 3900
rect 1256 3879 1258 3900
rect 1384 3879 1386 3900
rect 1512 3879 1514 3900
rect 1648 3879 1650 3900
rect 2006 3899 2012 3900
rect 2046 3899 2052 3900
rect 2008 3879 2010 3899
rect 2046 3895 2047 3899
rect 2051 3895 2052 3899
rect 3942 3899 3948 3900
rect 2046 3894 2052 3895
rect 2158 3896 2164 3897
rect 111 3878 115 3879
rect 111 3873 115 3874
rect 199 3878 203 3879
rect 199 3873 203 3874
rect 295 3878 299 3879
rect 295 3873 299 3874
rect 335 3878 339 3879
rect 335 3873 339 3874
rect 391 3878 395 3879
rect 391 3873 395 3874
rect 455 3878 459 3879
rect 455 3873 459 3874
rect 495 3878 499 3879
rect 495 3873 499 3874
rect 583 3878 587 3879
rect 583 3873 587 3874
rect 615 3878 619 3879
rect 615 3873 619 3874
rect 719 3878 723 3879
rect 719 3873 723 3874
rect 743 3878 747 3879
rect 743 3873 747 3874
rect 847 3878 851 3879
rect 847 3873 851 3874
rect 871 3878 875 3879
rect 871 3873 875 3874
rect 975 3878 979 3879
rect 975 3873 979 3874
rect 999 3878 1003 3879
rect 999 3873 1003 3874
rect 1103 3878 1107 3879
rect 1103 3873 1107 3874
rect 1127 3878 1131 3879
rect 1127 3873 1131 3874
rect 1231 3878 1235 3879
rect 1231 3873 1235 3874
rect 1255 3878 1259 3879
rect 1255 3873 1259 3874
rect 1359 3878 1363 3879
rect 1359 3873 1363 3874
rect 1383 3878 1387 3879
rect 1383 3873 1387 3874
rect 1487 3878 1491 3879
rect 1487 3873 1491 3874
rect 1511 3878 1515 3879
rect 1511 3873 1515 3874
rect 1647 3878 1651 3879
rect 1647 3873 1651 3874
rect 2007 3878 2011 3879
rect 2007 3873 2011 3874
rect 112 3853 114 3873
rect 110 3852 116 3853
rect 336 3852 338 3873
rect 456 3852 458 3873
rect 584 3852 586 3873
rect 720 3852 722 3873
rect 848 3852 850 3873
rect 976 3852 978 3873
rect 1104 3852 1106 3873
rect 1232 3852 1234 3873
rect 1360 3852 1362 3873
rect 1488 3852 1490 3873
rect 2008 3853 2010 3873
rect 2048 3859 2050 3894
rect 2158 3892 2159 3896
rect 2163 3892 2164 3896
rect 2158 3891 2164 3892
rect 2286 3896 2292 3897
rect 2286 3892 2287 3896
rect 2291 3892 2292 3896
rect 2286 3891 2292 3892
rect 2414 3896 2420 3897
rect 2414 3892 2415 3896
rect 2419 3892 2420 3896
rect 2414 3891 2420 3892
rect 2550 3896 2556 3897
rect 2550 3892 2551 3896
rect 2555 3892 2556 3896
rect 2550 3891 2556 3892
rect 2686 3896 2692 3897
rect 2686 3892 2687 3896
rect 2691 3892 2692 3896
rect 2686 3891 2692 3892
rect 2822 3896 2828 3897
rect 2822 3892 2823 3896
rect 2827 3892 2828 3896
rect 2822 3891 2828 3892
rect 2950 3896 2956 3897
rect 2950 3892 2951 3896
rect 2955 3892 2956 3896
rect 2950 3891 2956 3892
rect 3070 3896 3076 3897
rect 3070 3892 3071 3896
rect 3075 3892 3076 3896
rect 3070 3891 3076 3892
rect 3190 3896 3196 3897
rect 3190 3892 3191 3896
rect 3195 3892 3196 3896
rect 3190 3891 3196 3892
rect 3302 3896 3308 3897
rect 3302 3892 3303 3896
rect 3307 3892 3308 3896
rect 3302 3891 3308 3892
rect 3406 3896 3412 3897
rect 3406 3892 3407 3896
rect 3411 3892 3412 3896
rect 3406 3891 3412 3892
rect 3518 3896 3524 3897
rect 3518 3892 3519 3896
rect 3523 3892 3524 3896
rect 3518 3891 3524 3892
rect 3630 3896 3636 3897
rect 3630 3892 3631 3896
rect 3635 3892 3636 3896
rect 3630 3891 3636 3892
rect 3742 3896 3748 3897
rect 3742 3892 3743 3896
rect 3747 3892 3748 3896
rect 3942 3895 3943 3899
rect 3947 3895 3948 3899
rect 3942 3894 3948 3895
rect 3742 3891 3748 3892
rect 2160 3859 2162 3891
rect 2288 3859 2290 3891
rect 2416 3859 2418 3891
rect 2552 3859 2554 3891
rect 2688 3859 2690 3891
rect 2824 3859 2826 3891
rect 2952 3859 2954 3891
rect 3072 3859 3074 3891
rect 3192 3859 3194 3891
rect 3304 3859 3306 3891
rect 3408 3859 3410 3891
rect 3520 3859 3522 3891
rect 3632 3859 3634 3891
rect 3744 3859 3746 3891
rect 3944 3859 3946 3894
rect 2047 3858 2051 3859
rect 2047 3853 2051 3854
rect 2159 3858 2163 3859
rect 2159 3853 2163 3854
rect 2207 3858 2211 3859
rect 2207 3853 2211 3854
rect 2287 3858 2291 3859
rect 2287 3853 2291 3854
rect 2343 3858 2347 3859
rect 2343 3853 2347 3854
rect 2415 3858 2419 3859
rect 2415 3853 2419 3854
rect 2487 3858 2491 3859
rect 2487 3853 2491 3854
rect 2551 3858 2555 3859
rect 2551 3853 2555 3854
rect 2647 3858 2651 3859
rect 2647 3853 2651 3854
rect 2687 3858 2691 3859
rect 2687 3853 2691 3854
rect 2823 3858 2827 3859
rect 2823 3853 2827 3854
rect 2951 3858 2955 3859
rect 2951 3853 2955 3854
rect 3015 3858 3019 3859
rect 3015 3853 3019 3854
rect 3071 3858 3075 3859
rect 3071 3853 3075 3854
rect 3191 3858 3195 3859
rect 3191 3853 3195 3854
rect 3223 3858 3227 3859
rect 3223 3853 3227 3854
rect 3303 3858 3307 3859
rect 3303 3853 3307 3854
rect 3407 3858 3411 3859
rect 3407 3853 3411 3854
rect 3439 3858 3443 3859
rect 3439 3853 3443 3854
rect 3519 3858 3523 3859
rect 3519 3853 3523 3854
rect 3631 3858 3635 3859
rect 3631 3853 3635 3854
rect 3655 3858 3659 3859
rect 3655 3853 3659 3854
rect 3743 3858 3747 3859
rect 3743 3853 3747 3854
rect 3943 3858 3947 3859
rect 3943 3853 3947 3854
rect 2006 3852 2012 3853
rect 110 3848 111 3852
rect 115 3848 116 3852
rect 110 3847 116 3848
rect 334 3851 340 3852
rect 334 3847 335 3851
rect 339 3847 340 3851
rect 334 3846 340 3847
rect 454 3851 460 3852
rect 454 3847 455 3851
rect 459 3847 460 3851
rect 454 3846 460 3847
rect 582 3851 588 3852
rect 582 3847 583 3851
rect 587 3847 588 3851
rect 582 3846 588 3847
rect 718 3851 724 3852
rect 718 3847 719 3851
rect 723 3847 724 3851
rect 718 3846 724 3847
rect 846 3851 852 3852
rect 846 3847 847 3851
rect 851 3847 852 3851
rect 846 3846 852 3847
rect 974 3851 980 3852
rect 974 3847 975 3851
rect 979 3847 980 3851
rect 974 3846 980 3847
rect 1102 3851 1108 3852
rect 1102 3847 1103 3851
rect 1107 3847 1108 3851
rect 1102 3846 1108 3847
rect 1230 3851 1236 3852
rect 1230 3847 1231 3851
rect 1235 3847 1236 3851
rect 1230 3846 1236 3847
rect 1358 3851 1364 3852
rect 1358 3847 1359 3851
rect 1363 3847 1364 3851
rect 1358 3846 1364 3847
rect 1486 3851 1492 3852
rect 1486 3847 1487 3851
rect 1491 3847 1492 3851
rect 2006 3848 2007 3852
rect 2011 3848 2012 3852
rect 2006 3847 2012 3848
rect 1486 3846 1492 3847
rect 110 3835 116 3836
rect 110 3831 111 3835
rect 115 3831 116 3835
rect 2006 3835 2012 3836
rect 110 3830 116 3831
rect 334 3832 340 3833
rect 112 3799 114 3830
rect 334 3828 335 3832
rect 339 3828 340 3832
rect 334 3827 340 3828
rect 454 3832 460 3833
rect 454 3828 455 3832
rect 459 3828 460 3832
rect 454 3827 460 3828
rect 582 3832 588 3833
rect 582 3828 583 3832
rect 587 3828 588 3832
rect 582 3827 588 3828
rect 718 3832 724 3833
rect 718 3828 719 3832
rect 723 3828 724 3832
rect 718 3827 724 3828
rect 846 3832 852 3833
rect 846 3828 847 3832
rect 851 3828 852 3832
rect 846 3827 852 3828
rect 974 3832 980 3833
rect 974 3828 975 3832
rect 979 3828 980 3832
rect 974 3827 980 3828
rect 1102 3832 1108 3833
rect 1102 3828 1103 3832
rect 1107 3828 1108 3832
rect 1102 3827 1108 3828
rect 1230 3832 1236 3833
rect 1230 3828 1231 3832
rect 1235 3828 1236 3832
rect 1230 3827 1236 3828
rect 1358 3832 1364 3833
rect 1358 3828 1359 3832
rect 1363 3828 1364 3832
rect 1358 3827 1364 3828
rect 1486 3832 1492 3833
rect 1486 3828 1487 3832
rect 1491 3828 1492 3832
rect 2006 3831 2007 3835
rect 2011 3831 2012 3835
rect 2006 3830 2012 3831
rect 1486 3827 1492 3828
rect 336 3799 338 3827
rect 456 3799 458 3827
rect 584 3799 586 3827
rect 720 3799 722 3827
rect 848 3799 850 3827
rect 976 3799 978 3827
rect 1104 3799 1106 3827
rect 1232 3799 1234 3827
rect 1360 3799 1362 3827
rect 1488 3799 1490 3827
rect 2008 3799 2010 3830
rect 2048 3826 2050 3853
rect 2208 3829 2210 3853
rect 2344 3829 2346 3853
rect 2488 3829 2490 3853
rect 2648 3829 2650 3853
rect 2824 3829 2826 3853
rect 3016 3829 3018 3853
rect 3224 3829 3226 3853
rect 3440 3829 3442 3853
rect 3656 3829 3658 3853
rect 2206 3828 2212 3829
rect 2046 3825 2052 3826
rect 2046 3821 2047 3825
rect 2051 3821 2052 3825
rect 2206 3824 2207 3828
rect 2211 3824 2212 3828
rect 2206 3823 2212 3824
rect 2342 3828 2348 3829
rect 2342 3824 2343 3828
rect 2347 3824 2348 3828
rect 2342 3823 2348 3824
rect 2486 3828 2492 3829
rect 2486 3824 2487 3828
rect 2491 3824 2492 3828
rect 2486 3823 2492 3824
rect 2646 3828 2652 3829
rect 2646 3824 2647 3828
rect 2651 3824 2652 3828
rect 2646 3823 2652 3824
rect 2822 3828 2828 3829
rect 2822 3824 2823 3828
rect 2827 3824 2828 3828
rect 2822 3823 2828 3824
rect 3014 3828 3020 3829
rect 3014 3824 3015 3828
rect 3019 3824 3020 3828
rect 3014 3823 3020 3824
rect 3222 3828 3228 3829
rect 3222 3824 3223 3828
rect 3227 3824 3228 3828
rect 3222 3823 3228 3824
rect 3438 3828 3444 3829
rect 3438 3824 3439 3828
rect 3443 3824 3444 3828
rect 3438 3823 3444 3824
rect 3654 3828 3660 3829
rect 3654 3824 3655 3828
rect 3659 3824 3660 3828
rect 3944 3826 3946 3853
rect 3654 3823 3660 3824
rect 3942 3825 3948 3826
rect 2046 3820 2052 3821
rect 3942 3821 3943 3825
rect 3947 3821 3948 3825
rect 3942 3820 3948 3821
rect 2206 3809 2212 3810
rect 2046 3808 2052 3809
rect 2046 3804 2047 3808
rect 2051 3804 2052 3808
rect 2206 3805 2207 3809
rect 2211 3805 2212 3809
rect 2206 3804 2212 3805
rect 2342 3809 2348 3810
rect 2342 3805 2343 3809
rect 2347 3805 2348 3809
rect 2342 3804 2348 3805
rect 2486 3809 2492 3810
rect 2486 3805 2487 3809
rect 2491 3805 2492 3809
rect 2486 3804 2492 3805
rect 2646 3809 2652 3810
rect 2646 3805 2647 3809
rect 2651 3805 2652 3809
rect 2646 3804 2652 3805
rect 2822 3809 2828 3810
rect 2822 3805 2823 3809
rect 2827 3805 2828 3809
rect 2822 3804 2828 3805
rect 3014 3809 3020 3810
rect 3014 3805 3015 3809
rect 3019 3805 3020 3809
rect 3014 3804 3020 3805
rect 3222 3809 3228 3810
rect 3222 3805 3223 3809
rect 3227 3805 3228 3809
rect 3222 3804 3228 3805
rect 3438 3809 3444 3810
rect 3438 3805 3439 3809
rect 3443 3805 3444 3809
rect 3438 3804 3444 3805
rect 3654 3809 3660 3810
rect 3654 3805 3655 3809
rect 3659 3805 3660 3809
rect 3654 3804 3660 3805
rect 3942 3808 3948 3809
rect 3942 3804 3943 3808
rect 3947 3804 3948 3808
rect 2046 3803 2052 3804
rect 111 3798 115 3799
rect 111 3793 115 3794
rect 335 3798 339 3799
rect 335 3793 339 3794
rect 455 3798 459 3799
rect 455 3793 459 3794
rect 503 3798 507 3799
rect 503 3793 507 3794
rect 583 3798 587 3799
rect 583 3793 587 3794
rect 615 3798 619 3799
rect 615 3793 619 3794
rect 719 3798 723 3799
rect 719 3793 723 3794
rect 735 3798 739 3799
rect 735 3793 739 3794
rect 847 3798 851 3799
rect 847 3793 851 3794
rect 863 3798 867 3799
rect 863 3793 867 3794
rect 975 3798 979 3799
rect 975 3793 979 3794
rect 999 3798 1003 3799
rect 999 3793 1003 3794
rect 1103 3798 1107 3799
rect 1103 3793 1107 3794
rect 1143 3798 1147 3799
rect 1143 3793 1147 3794
rect 1231 3798 1235 3799
rect 1231 3793 1235 3794
rect 1287 3798 1291 3799
rect 1287 3793 1291 3794
rect 1359 3798 1363 3799
rect 1359 3793 1363 3794
rect 1431 3798 1435 3799
rect 1431 3793 1435 3794
rect 1487 3798 1491 3799
rect 1487 3793 1491 3794
rect 1583 3798 1587 3799
rect 1583 3793 1587 3794
rect 2007 3798 2011 3799
rect 2007 3793 2011 3794
rect 112 3766 114 3793
rect 504 3769 506 3793
rect 616 3769 618 3793
rect 736 3769 738 3793
rect 864 3769 866 3793
rect 1000 3769 1002 3793
rect 1144 3769 1146 3793
rect 1288 3769 1290 3793
rect 1432 3769 1434 3793
rect 1584 3769 1586 3793
rect 502 3768 508 3769
rect 110 3765 116 3766
rect 110 3761 111 3765
rect 115 3761 116 3765
rect 502 3764 503 3768
rect 507 3764 508 3768
rect 502 3763 508 3764
rect 614 3768 620 3769
rect 614 3764 615 3768
rect 619 3764 620 3768
rect 614 3763 620 3764
rect 734 3768 740 3769
rect 734 3764 735 3768
rect 739 3764 740 3768
rect 734 3763 740 3764
rect 862 3768 868 3769
rect 862 3764 863 3768
rect 867 3764 868 3768
rect 862 3763 868 3764
rect 998 3768 1004 3769
rect 998 3764 999 3768
rect 1003 3764 1004 3768
rect 998 3763 1004 3764
rect 1142 3768 1148 3769
rect 1142 3764 1143 3768
rect 1147 3764 1148 3768
rect 1142 3763 1148 3764
rect 1286 3768 1292 3769
rect 1286 3764 1287 3768
rect 1291 3764 1292 3768
rect 1286 3763 1292 3764
rect 1430 3768 1436 3769
rect 1430 3764 1431 3768
rect 1435 3764 1436 3768
rect 1430 3763 1436 3764
rect 1582 3768 1588 3769
rect 1582 3764 1583 3768
rect 1587 3764 1588 3768
rect 2008 3766 2010 3793
rect 2048 3783 2050 3803
rect 2208 3783 2210 3804
rect 2344 3783 2346 3804
rect 2488 3783 2490 3804
rect 2648 3783 2650 3804
rect 2824 3783 2826 3804
rect 3016 3783 3018 3804
rect 3224 3783 3226 3804
rect 3440 3783 3442 3804
rect 3656 3783 3658 3804
rect 3942 3803 3948 3804
rect 3944 3783 3946 3803
rect 2047 3782 2051 3783
rect 2047 3777 2051 3778
rect 2191 3782 2195 3783
rect 2191 3777 2195 3778
rect 2207 3782 2211 3783
rect 2207 3777 2211 3778
rect 2343 3782 2347 3783
rect 2343 3777 2347 3778
rect 2375 3782 2379 3783
rect 2375 3777 2379 3778
rect 2487 3782 2491 3783
rect 2487 3777 2491 3778
rect 2559 3782 2563 3783
rect 2559 3777 2563 3778
rect 2647 3782 2651 3783
rect 2647 3777 2651 3778
rect 2743 3782 2747 3783
rect 2743 3777 2747 3778
rect 2823 3782 2827 3783
rect 2823 3777 2827 3778
rect 2935 3782 2939 3783
rect 2935 3777 2939 3778
rect 3015 3782 3019 3783
rect 3015 3777 3019 3778
rect 3127 3782 3131 3783
rect 3127 3777 3131 3778
rect 3223 3782 3227 3783
rect 3223 3777 3227 3778
rect 3319 3782 3323 3783
rect 3319 3777 3323 3778
rect 3439 3782 3443 3783
rect 3439 3777 3443 3778
rect 3511 3782 3515 3783
rect 3511 3777 3515 3778
rect 3655 3782 3659 3783
rect 3655 3777 3659 3778
rect 3711 3782 3715 3783
rect 3711 3777 3715 3778
rect 3943 3782 3947 3783
rect 3943 3777 3947 3778
rect 1582 3763 1588 3764
rect 2006 3765 2012 3766
rect 110 3760 116 3761
rect 2006 3761 2007 3765
rect 2011 3761 2012 3765
rect 2006 3760 2012 3761
rect 2048 3757 2050 3777
rect 2046 3756 2052 3757
rect 2192 3756 2194 3777
rect 2376 3756 2378 3777
rect 2560 3756 2562 3777
rect 2744 3756 2746 3777
rect 2936 3756 2938 3777
rect 3128 3756 3130 3777
rect 3320 3756 3322 3777
rect 3512 3756 3514 3777
rect 3712 3756 3714 3777
rect 3944 3757 3946 3777
rect 3942 3756 3948 3757
rect 2046 3752 2047 3756
rect 2051 3752 2052 3756
rect 2046 3751 2052 3752
rect 2190 3755 2196 3756
rect 2190 3751 2191 3755
rect 2195 3751 2196 3755
rect 2190 3750 2196 3751
rect 2374 3755 2380 3756
rect 2374 3751 2375 3755
rect 2379 3751 2380 3755
rect 2374 3750 2380 3751
rect 2558 3755 2564 3756
rect 2558 3751 2559 3755
rect 2563 3751 2564 3755
rect 2558 3750 2564 3751
rect 2742 3755 2748 3756
rect 2742 3751 2743 3755
rect 2747 3751 2748 3755
rect 2742 3750 2748 3751
rect 2934 3755 2940 3756
rect 2934 3751 2935 3755
rect 2939 3751 2940 3755
rect 2934 3750 2940 3751
rect 3126 3755 3132 3756
rect 3126 3751 3127 3755
rect 3131 3751 3132 3755
rect 3126 3750 3132 3751
rect 3318 3755 3324 3756
rect 3318 3751 3319 3755
rect 3323 3751 3324 3755
rect 3318 3750 3324 3751
rect 3510 3755 3516 3756
rect 3510 3751 3511 3755
rect 3515 3751 3516 3755
rect 3510 3750 3516 3751
rect 3710 3755 3716 3756
rect 3710 3751 3711 3755
rect 3715 3751 3716 3755
rect 3942 3752 3943 3756
rect 3947 3752 3948 3756
rect 3942 3751 3948 3752
rect 3710 3750 3716 3751
rect 502 3749 508 3750
rect 110 3748 116 3749
rect 110 3744 111 3748
rect 115 3744 116 3748
rect 502 3745 503 3749
rect 507 3745 508 3749
rect 502 3744 508 3745
rect 614 3749 620 3750
rect 614 3745 615 3749
rect 619 3745 620 3749
rect 614 3744 620 3745
rect 734 3749 740 3750
rect 734 3745 735 3749
rect 739 3745 740 3749
rect 734 3744 740 3745
rect 862 3749 868 3750
rect 862 3745 863 3749
rect 867 3745 868 3749
rect 862 3744 868 3745
rect 998 3749 1004 3750
rect 998 3745 999 3749
rect 1003 3745 1004 3749
rect 998 3744 1004 3745
rect 1142 3749 1148 3750
rect 1142 3745 1143 3749
rect 1147 3745 1148 3749
rect 1142 3744 1148 3745
rect 1286 3749 1292 3750
rect 1286 3745 1287 3749
rect 1291 3745 1292 3749
rect 1286 3744 1292 3745
rect 1430 3749 1436 3750
rect 1430 3745 1431 3749
rect 1435 3745 1436 3749
rect 1430 3744 1436 3745
rect 1582 3749 1588 3750
rect 1582 3745 1583 3749
rect 1587 3745 1588 3749
rect 1582 3744 1588 3745
rect 2006 3748 2012 3749
rect 2006 3744 2007 3748
rect 2011 3744 2012 3748
rect 110 3743 116 3744
rect 112 3715 114 3743
rect 504 3715 506 3744
rect 616 3715 618 3744
rect 736 3715 738 3744
rect 864 3715 866 3744
rect 1000 3715 1002 3744
rect 1144 3715 1146 3744
rect 1288 3715 1290 3744
rect 1432 3715 1434 3744
rect 1584 3715 1586 3744
rect 2006 3743 2012 3744
rect 2008 3715 2010 3743
rect 2046 3739 2052 3740
rect 2046 3735 2047 3739
rect 2051 3735 2052 3739
rect 3942 3739 3948 3740
rect 2046 3734 2052 3735
rect 2190 3736 2196 3737
rect 111 3714 115 3715
rect 111 3709 115 3710
rect 495 3714 499 3715
rect 495 3709 499 3710
rect 503 3714 507 3715
rect 503 3709 507 3710
rect 591 3714 595 3715
rect 591 3709 595 3710
rect 615 3714 619 3715
rect 615 3709 619 3710
rect 687 3714 691 3715
rect 687 3709 691 3710
rect 735 3714 739 3715
rect 735 3709 739 3710
rect 791 3714 795 3715
rect 791 3709 795 3710
rect 863 3714 867 3715
rect 863 3709 867 3710
rect 911 3714 915 3715
rect 911 3709 915 3710
rect 999 3714 1003 3715
rect 999 3709 1003 3710
rect 1039 3714 1043 3715
rect 1039 3709 1043 3710
rect 1143 3714 1147 3715
rect 1143 3709 1147 3710
rect 1183 3714 1187 3715
rect 1183 3709 1187 3710
rect 1287 3714 1291 3715
rect 1287 3709 1291 3710
rect 1335 3714 1339 3715
rect 1335 3709 1339 3710
rect 1431 3714 1435 3715
rect 1431 3709 1435 3710
rect 1495 3714 1499 3715
rect 1495 3709 1499 3710
rect 1583 3714 1587 3715
rect 1583 3709 1587 3710
rect 1655 3714 1659 3715
rect 1655 3709 1659 3710
rect 2007 3714 2011 3715
rect 2007 3709 2011 3710
rect 112 3689 114 3709
rect 110 3688 116 3689
rect 496 3688 498 3709
rect 592 3688 594 3709
rect 688 3688 690 3709
rect 792 3688 794 3709
rect 912 3688 914 3709
rect 1040 3688 1042 3709
rect 1184 3688 1186 3709
rect 1336 3688 1338 3709
rect 1496 3688 1498 3709
rect 1656 3688 1658 3709
rect 2008 3689 2010 3709
rect 2048 3703 2050 3734
rect 2190 3732 2191 3736
rect 2195 3732 2196 3736
rect 2190 3731 2196 3732
rect 2374 3736 2380 3737
rect 2374 3732 2375 3736
rect 2379 3732 2380 3736
rect 2374 3731 2380 3732
rect 2558 3736 2564 3737
rect 2558 3732 2559 3736
rect 2563 3732 2564 3736
rect 2558 3731 2564 3732
rect 2742 3736 2748 3737
rect 2742 3732 2743 3736
rect 2747 3732 2748 3736
rect 2742 3731 2748 3732
rect 2934 3736 2940 3737
rect 2934 3732 2935 3736
rect 2939 3732 2940 3736
rect 2934 3731 2940 3732
rect 3126 3736 3132 3737
rect 3126 3732 3127 3736
rect 3131 3732 3132 3736
rect 3126 3731 3132 3732
rect 3318 3736 3324 3737
rect 3318 3732 3319 3736
rect 3323 3732 3324 3736
rect 3318 3731 3324 3732
rect 3510 3736 3516 3737
rect 3510 3732 3511 3736
rect 3515 3732 3516 3736
rect 3510 3731 3516 3732
rect 3710 3736 3716 3737
rect 3710 3732 3711 3736
rect 3715 3732 3716 3736
rect 3942 3735 3943 3739
rect 3947 3735 3948 3739
rect 3942 3734 3948 3735
rect 3710 3731 3716 3732
rect 2192 3703 2194 3731
rect 2376 3703 2378 3731
rect 2560 3703 2562 3731
rect 2744 3703 2746 3731
rect 2936 3703 2938 3731
rect 3128 3703 3130 3731
rect 3320 3703 3322 3731
rect 3512 3703 3514 3731
rect 3712 3703 3714 3731
rect 3944 3703 3946 3734
rect 2047 3702 2051 3703
rect 2047 3697 2051 3698
rect 2127 3702 2131 3703
rect 2127 3697 2131 3698
rect 2191 3702 2195 3703
rect 2191 3697 2195 3698
rect 2351 3702 2355 3703
rect 2351 3697 2355 3698
rect 2375 3702 2379 3703
rect 2375 3697 2379 3698
rect 2559 3702 2563 3703
rect 2559 3697 2563 3698
rect 2583 3702 2587 3703
rect 2583 3697 2587 3698
rect 2743 3702 2747 3703
rect 2743 3697 2747 3698
rect 2815 3702 2819 3703
rect 2815 3697 2819 3698
rect 2935 3702 2939 3703
rect 2935 3697 2939 3698
rect 3047 3702 3051 3703
rect 3047 3697 3051 3698
rect 3127 3702 3131 3703
rect 3127 3697 3131 3698
rect 3279 3702 3283 3703
rect 3279 3697 3283 3698
rect 3319 3702 3323 3703
rect 3319 3697 3323 3698
rect 3511 3702 3515 3703
rect 3511 3697 3515 3698
rect 3711 3702 3715 3703
rect 3711 3697 3715 3698
rect 3751 3702 3755 3703
rect 3751 3697 3755 3698
rect 3943 3702 3947 3703
rect 3943 3697 3947 3698
rect 2006 3688 2012 3689
rect 110 3684 111 3688
rect 115 3684 116 3688
rect 110 3683 116 3684
rect 494 3687 500 3688
rect 494 3683 495 3687
rect 499 3683 500 3687
rect 494 3682 500 3683
rect 590 3687 596 3688
rect 590 3683 591 3687
rect 595 3683 596 3687
rect 590 3682 596 3683
rect 686 3687 692 3688
rect 686 3683 687 3687
rect 691 3683 692 3687
rect 686 3682 692 3683
rect 790 3687 796 3688
rect 790 3683 791 3687
rect 795 3683 796 3687
rect 790 3682 796 3683
rect 910 3687 916 3688
rect 910 3683 911 3687
rect 915 3683 916 3687
rect 910 3682 916 3683
rect 1038 3687 1044 3688
rect 1038 3683 1039 3687
rect 1043 3683 1044 3687
rect 1038 3682 1044 3683
rect 1182 3687 1188 3688
rect 1182 3683 1183 3687
rect 1187 3683 1188 3687
rect 1182 3682 1188 3683
rect 1334 3687 1340 3688
rect 1334 3683 1335 3687
rect 1339 3683 1340 3687
rect 1334 3682 1340 3683
rect 1494 3687 1500 3688
rect 1494 3683 1495 3687
rect 1499 3683 1500 3687
rect 1494 3682 1500 3683
rect 1654 3687 1660 3688
rect 1654 3683 1655 3687
rect 1659 3683 1660 3687
rect 2006 3684 2007 3688
rect 2011 3684 2012 3688
rect 2006 3683 2012 3684
rect 1654 3682 1660 3683
rect 110 3671 116 3672
rect 110 3667 111 3671
rect 115 3667 116 3671
rect 2006 3671 2012 3672
rect 110 3666 116 3667
rect 494 3668 500 3669
rect 112 3631 114 3666
rect 494 3664 495 3668
rect 499 3664 500 3668
rect 494 3663 500 3664
rect 590 3668 596 3669
rect 590 3664 591 3668
rect 595 3664 596 3668
rect 590 3663 596 3664
rect 686 3668 692 3669
rect 686 3664 687 3668
rect 691 3664 692 3668
rect 686 3663 692 3664
rect 790 3668 796 3669
rect 790 3664 791 3668
rect 795 3664 796 3668
rect 790 3663 796 3664
rect 910 3668 916 3669
rect 910 3664 911 3668
rect 915 3664 916 3668
rect 910 3663 916 3664
rect 1038 3668 1044 3669
rect 1038 3664 1039 3668
rect 1043 3664 1044 3668
rect 1038 3663 1044 3664
rect 1182 3668 1188 3669
rect 1182 3664 1183 3668
rect 1187 3664 1188 3668
rect 1182 3663 1188 3664
rect 1334 3668 1340 3669
rect 1334 3664 1335 3668
rect 1339 3664 1340 3668
rect 1334 3663 1340 3664
rect 1494 3668 1500 3669
rect 1494 3664 1495 3668
rect 1499 3664 1500 3668
rect 1494 3663 1500 3664
rect 1654 3668 1660 3669
rect 1654 3664 1655 3668
rect 1659 3664 1660 3668
rect 2006 3667 2007 3671
rect 2011 3667 2012 3671
rect 2048 3670 2050 3697
rect 2128 3673 2130 3697
rect 2352 3673 2354 3697
rect 2584 3673 2586 3697
rect 2816 3673 2818 3697
rect 3048 3673 3050 3697
rect 3280 3673 3282 3697
rect 3512 3673 3514 3697
rect 3752 3673 3754 3697
rect 2126 3672 2132 3673
rect 2006 3666 2012 3667
rect 2046 3669 2052 3670
rect 1654 3663 1660 3664
rect 496 3631 498 3663
rect 592 3631 594 3663
rect 688 3631 690 3663
rect 792 3631 794 3663
rect 912 3631 914 3663
rect 1040 3631 1042 3663
rect 1184 3631 1186 3663
rect 1336 3631 1338 3663
rect 1496 3631 1498 3663
rect 1656 3631 1658 3663
rect 2008 3631 2010 3666
rect 2046 3665 2047 3669
rect 2051 3665 2052 3669
rect 2126 3668 2127 3672
rect 2131 3668 2132 3672
rect 2126 3667 2132 3668
rect 2350 3672 2356 3673
rect 2350 3668 2351 3672
rect 2355 3668 2356 3672
rect 2350 3667 2356 3668
rect 2582 3672 2588 3673
rect 2582 3668 2583 3672
rect 2587 3668 2588 3672
rect 2582 3667 2588 3668
rect 2814 3672 2820 3673
rect 2814 3668 2815 3672
rect 2819 3668 2820 3672
rect 2814 3667 2820 3668
rect 3046 3672 3052 3673
rect 3046 3668 3047 3672
rect 3051 3668 3052 3672
rect 3046 3667 3052 3668
rect 3278 3672 3284 3673
rect 3278 3668 3279 3672
rect 3283 3668 3284 3672
rect 3278 3667 3284 3668
rect 3510 3672 3516 3673
rect 3510 3668 3511 3672
rect 3515 3668 3516 3672
rect 3510 3667 3516 3668
rect 3750 3672 3756 3673
rect 3750 3668 3751 3672
rect 3755 3668 3756 3672
rect 3944 3670 3946 3697
rect 3750 3667 3756 3668
rect 3942 3669 3948 3670
rect 2046 3664 2052 3665
rect 3942 3665 3943 3669
rect 3947 3665 3948 3669
rect 3942 3664 3948 3665
rect 2126 3653 2132 3654
rect 2046 3652 2052 3653
rect 2046 3648 2047 3652
rect 2051 3648 2052 3652
rect 2126 3649 2127 3653
rect 2131 3649 2132 3653
rect 2126 3648 2132 3649
rect 2350 3653 2356 3654
rect 2350 3649 2351 3653
rect 2355 3649 2356 3653
rect 2350 3648 2356 3649
rect 2582 3653 2588 3654
rect 2582 3649 2583 3653
rect 2587 3649 2588 3653
rect 2582 3648 2588 3649
rect 2814 3653 2820 3654
rect 2814 3649 2815 3653
rect 2819 3649 2820 3653
rect 2814 3648 2820 3649
rect 3046 3653 3052 3654
rect 3046 3649 3047 3653
rect 3051 3649 3052 3653
rect 3046 3648 3052 3649
rect 3278 3653 3284 3654
rect 3278 3649 3279 3653
rect 3283 3649 3284 3653
rect 3278 3648 3284 3649
rect 3510 3653 3516 3654
rect 3510 3649 3511 3653
rect 3515 3649 3516 3653
rect 3510 3648 3516 3649
rect 3750 3653 3756 3654
rect 3750 3649 3751 3653
rect 3755 3649 3756 3653
rect 3750 3648 3756 3649
rect 3942 3652 3948 3653
rect 3942 3648 3943 3652
rect 3947 3648 3948 3652
rect 2046 3647 2052 3648
rect 111 3630 115 3631
rect 111 3625 115 3626
rect 335 3630 339 3631
rect 335 3625 339 3626
rect 463 3630 467 3631
rect 463 3625 467 3626
rect 495 3630 499 3631
rect 495 3625 499 3626
rect 591 3630 595 3631
rect 591 3625 595 3626
rect 607 3630 611 3631
rect 607 3625 611 3626
rect 687 3630 691 3631
rect 687 3625 691 3626
rect 759 3630 763 3631
rect 759 3625 763 3626
rect 791 3630 795 3631
rect 791 3625 795 3626
rect 911 3630 915 3631
rect 911 3625 915 3626
rect 927 3630 931 3631
rect 927 3625 931 3626
rect 1039 3630 1043 3631
rect 1039 3625 1043 3626
rect 1095 3630 1099 3631
rect 1095 3625 1099 3626
rect 1183 3630 1187 3631
rect 1183 3625 1187 3626
rect 1263 3630 1267 3631
rect 1263 3625 1267 3626
rect 1335 3630 1339 3631
rect 1335 3625 1339 3626
rect 1439 3630 1443 3631
rect 1439 3625 1443 3626
rect 1495 3630 1499 3631
rect 1495 3625 1499 3626
rect 1615 3630 1619 3631
rect 1615 3625 1619 3626
rect 1655 3630 1659 3631
rect 1655 3625 1659 3626
rect 1791 3630 1795 3631
rect 1791 3625 1795 3626
rect 2007 3630 2011 3631
rect 2007 3625 2011 3626
rect 112 3598 114 3625
rect 336 3601 338 3625
rect 464 3601 466 3625
rect 608 3601 610 3625
rect 760 3601 762 3625
rect 928 3601 930 3625
rect 1096 3601 1098 3625
rect 1264 3601 1266 3625
rect 1440 3601 1442 3625
rect 1616 3601 1618 3625
rect 1792 3601 1794 3625
rect 334 3600 340 3601
rect 110 3597 116 3598
rect 110 3593 111 3597
rect 115 3593 116 3597
rect 334 3596 335 3600
rect 339 3596 340 3600
rect 334 3595 340 3596
rect 462 3600 468 3601
rect 462 3596 463 3600
rect 467 3596 468 3600
rect 462 3595 468 3596
rect 606 3600 612 3601
rect 606 3596 607 3600
rect 611 3596 612 3600
rect 606 3595 612 3596
rect 758 3600 764 3601
rect 758 3596 759 3600
rect 763 3596 764 3600
rect 758 3595 764 3596
rect 926 3600 932 3601
rect 926 3596 927 3600
rect 931 3596 932 3600
rect 926 3595 932 3596
rect 1094 3600 1100 3601
rect 1094 3596 1095 3600
rect 1099 3596 1100 3600
rect 1094 3595 1100 3596
rect 1262 3600 1268 3601
rect 1262 3596 1263 3600
rect 1267 3596 1268 3600
rect 1262 3595 1268 3596
rect 1438 3600 1444 3601
rect 1438 3596 1439 3600
rect 1443 3596 1444 3600
rect 1438 3595 1444 3596
rect 1614 3600 1620 3601
rect 1614 3596 1615 3600
rect 1619 3596 1620 3600
rect 1614 3595 1620 3596
rect 1790 3600 1796 3601
rect 1790 3596 1791 3600
rect 1795 3596 1796 3600
rect 2008 3598 2010 3625
rect 2048 3619 2050 3647
rect 2128 3619 2130 3648
rect 2352 3619 2354 3648
rect 2584 3619 2586 3648
rect 2816 3619 2818 3648
rect 3048 3619 3050 3648
rect 3280 3619 3282 3648
rect 3512 3619 3514 3648
rect 3752 3619 3754 3648
rect 3942 3647 3948 3648
rect 3944 3619 3946 3647
rect 2047 3618 2051 3619
rect 2047 3613 2051 3614
rect 2127 3618 2131 3619
rect 2127 3613 2131 3614
rect 2191 3618 2195 3619
rect 2191 3613 2195 3614
rect 2327 3618 2331 3619
rect 2327 3613 2331 3614
rect 2351 3618 2355 3619
rect 2351 3613 2355 3614
rect 2455 3618 2459 3619
rect 2455 3613 2459 3614
rect 2583 3618 2587 3619
rect 2583 3613 2587 3614
rect 2719 3618 2723 3619
rect 2719 3613 2723 3614
rect 2815 3618 2819 3619
rect 2815 3613 2819 3614
rect 2855 3618 2859 3619
rect 2855 3613 2859 3614
rect 2999 3618 3003 3619
rect 2999 3613 3003 3614
rect 3047 3618 3051 3619
rect 3047 3613 3051 3614
rect 3143 3618 3147 3619
rect 3143 3613 3147 3614
rect 3279 3618 3283 3619
rect 3279 3613 3283 3614
rect 3295 3618 3299 3619
rect 3295 3613 3299 3614
rect 3455 3618 3459 3619
rect 3455 3613 3459 3614
rect 3511 3618 3515 3619
rect 3511 3613 3515 3614
rect 3623 3618 3627 3619
rect 3623 3613 3627 3614
rect 3751 3618 3755 3619
rect 3751 3613 3755 3614
rect 3943 3618 3947 3619
rect 3943 3613 3947 3614
rect 1790 3595 1796 3596
rect 2006 3597 2012 3598
rect 110 3592 116 3593
rect 2006 3593 2007 3597
rect 2011 3593 2012 3597
rect 2048 3593 2050 3613
rect 2006 3592 2012 3593
rect 2046 3592 2052 3593
rect 2192 3592 2194 3613
rect 2328 3592 2330 3613
rect 2456 3592 2458 3613
rect 2584 3592 2586 3613
rect 2720 3592 2722 3613
rect 2856 3592 2858 3613
rect 3000 3592 3002 3613
rect 3144 3592 3146 3613
rect 3296 3592 3298 3613
rect 3456 3592 3458 3613
rect 3624 3592 3626 3613
rect 3944 3593 3946 3613
rect 3942 3592 3948 3593
rect 2046 3588 2047 3592
rect 2051 3588 2052 3592
rect 2046 3587 2052 3588
rect 2190 3591 2196 3592
rect 2190 3587 2191 3591
rect 2195 3587 2196 3591
rect 2190 3586 2196 3587
rect 2326 3591 2332 3592
rect 2326 3587 2327 3591
rect 2331 3587 2332 3591
rect 2326 3586 2332 3587
rect 2454 3591 2460 3592
rect 2454 3587 2455 3591
rect 2459 3587 2460 3591
rect 2454 3586 2460 3587
rect 2582 3591 2588 3592
rect 2582 3587 2583 3591
rect 2587 3587 2588 3591
rect 2582 3586 2588 3587
rect 2718 3591 2724 3592
rect 2718 3587 2719 3591
rect 2723 3587 2724 3591
rect 2718 3586 2724 3587
rect 2854 3591 2860 3592
rect 2854 3587 2855 3591
rect 2859 3587 2860 3591
rect 2854 3586 2860 3587
rect 2998 3591 3004 3592
rect 2998 3587 2999 3591
rect 3003 3587 3004 3591
rect 2998 3586 3004 3587
rect 3142 3591 3148 3592
rect 3142 3587 3143 3591
rect 3147 3587 3148 3591
rect 3142 3586 3148 3587
rect 3294 3591 3300 3592
rect 3294 3587 3295 3591
rect 3299 3587 3300 3591
rect 3294 3586 3300 3587
rect 3454 3591 3460 3592
rect 3454 3587 3455 3591
rect 3459 3587 3460 3591
rect 3454 3586 3460 3587
rect 3622 3591 3628 3592
rect 3622 3587 3623 3591
rect 3627 3587 3628 3591
rect 3942 3588 3943 3592
rect 3947 3588 3948 3592
rect 3942 3587 3948 3588
rect 3622 3586 3628 3587
rect 334 3581 340 3582
rect 110 3580 116 3581
rect 110 3576 111 3580
rect 115 3576 116 3580
rect 334 3577 335 3581
rect 339 3577 340 3581
rect 334 3576 340 3577
rect 462 3581 468 3582
rect 462 3577 463 3581
rect 467 3577 468 3581
rect 462 3576 468 3577
rect 606 3581 612 3582
rect 606 3577 607 3581
rect 611 3577 612 3581
rect 606 3576 612 3577
rect 758 3581 764 3582
rect 758 3577 759 3581
rect 763 3577 764 3581
rect 758 3576 764 3577
rect 926 3581 932 3582
rect 926 3577 927 3581
rect 931 3577 932 3581
rect 926 3576 932 3577
rect 1094 3581 1100 3582
rect 1094 3577 1095 3581
rect 1099 3577 1100 3581
rect 1094 3576 1100 3577
rect 1262 3581 1268 3582
rect 1262 3577 1263 3581
rect 1267 3577 1268 3581
rect 1262 3576 1268 3577
rect 1438 3581 1444 3582
rect 1438 3577 1439 3581
rect 1443 3577 1444 3581
rect 1438 3576 1444 3577
rect 1614 3581 1620 3582
rect 1614 3577 1615 3581
rect 1619 3577 1620 3581
rect 1614 3576 1620 3577
rect 1790 3581 1796 3582
rect 1790 3577 1791 3581
rect 1795 3577 1796 3581
rect 1790 3576 1796 3577
rect 2006 3580 2012 3581
rect 2006 3576 2007 3580
rect 2011 3576 2012 3580
rect 110 3575 116 3576
rect 112 3543 114 3575
rect 336 3543 338 3576
rect 464 3543 466 3576
rect 608 3543 610 3576
rect 760 3543 762 3576
rect 928 3543 930 3576
rect 1096 3543 1098 3576
rect 1264 3543 1266 3576
rect 1440 3543 1442 3576
rect 1616 3543 1618 3576
rect 1792 3543 1794 3576
rect 2006 3575 2012 3576
rect 2046 3575 2052 3576
rect 2008 3543 2010 3575
rect 2046 3571 2047 3575
rect 2051 3571 2052 3575
rect 3942 3575 3948 3576
rect 2046 3570 2052 3571
rect 2190 3572 2196 3573
rect 2048 3543 2050 3570
rect 2190 3568 2191 3572
rect 2195 3568 2196 3572
rect 2190 3567 2196 3568
rect 2326 3572 2332 3573
rect 2326 3568 2327 3572
rect 2331 3568 2332 3572
rect 2326 3567 2332 3568
rect 2454 3572 2460 3573
rect 2454 3568 2455 3572
rect 2459 3568 2460 3572
rect 2454 3567 2460 3568
rect 2582 3572 2588 3573
rect 2582 3568 2583 3572
rect 2587 3568 2588 3572
rect 2582 3567 2588 3568
rect 2718 3572 2724 3573
rect 2718 3568 2719 3572
rect 2723 3568 2724 3572
rect 2718 3567 2724 3568
rect 2854 3572 2860 3573
rect 2854 3568 2855 3572
rect 2859 3568 2860 3572
rect 2854 3567 2860 3568
rect 2998 3572 3004 3573
rect 2998 3568 2999 3572
rect 3003 3568 3004 3572
rect 2998 3567 3004 3568
rect 3142 3572 3148 3573
rect 3142 3568 3143 3572
rect 3147 3568 3148 3572
rect 3142 3567 3148 3568
rect 3294 3572 3300 3573
rect 3294 3568 3295 3572
rect 3299 3568 3300 3572
rect 3294 3567 3300 3568
rect 3454 3572 3460 3573
rect 3454 3568 3455 3572
rect 3459 3568 3460 3572
rect 3454 3567 3460 3568
rect 3622 3572 3628 3573
rect 3622 3568 3623 3572
rect 3627 3568 3628 3572
rect 3942 3571 3943 3575
rect 3947 3571 3948 3575
rect 3942 3570 3948 3571
rect 3622 3567 3628 3568
rect 2192 3543 2194 3567
rect 2328 3543 2330 3567
rect 2456 3543 2458 3567
rect 2584 3543 2586 3567
rect 2720 3543 2722 3567
rect 2856 3543 2858 3567
rect 3000 3543 3002 3567
rect 3144 3543 3146 3567
rect 3296 3543 3298 3567
rect 3456 3543 3458 3567
rect 3624 3543 3626 3567
rect 3944 3543 3946 3570
rect 111 3542 115 3543
rect 111 3537 115 3538
rect 159 3542 163 3543
rect 159 3537 163 3538
rect 303 3542 307 3543
rect 303 3537 307 3538
rect 335 3542 339 3543
rect 335 3537 339 3538
rect 463 3542 467 3543
rect 463 3537 467 3538
rect 607 3542 611 3543
rect 607 3537 611 3538
rect 639 3542 643 3543
rect 639 3537 643 3538
rect 759 3542 763 3543
rect 759 3537 763 3538
rect 815 3542 819 3543
rect 815 3537 819 3538
rect 927 3542 931 3543
rect 927 3537 931 3538
rect 999 3542 1003 3543
rect 999 3537 1003 3538
rect 1095 3542 1099 3543
rect 1095 3537 1099 3538
rect 1175 3542 1179 3543
rect 1175 3537 1179 3538
rect 1263 3542 1267 3543
rect 1263 3537 1267 3538
rect 1351 3542 1355 3543
rect 1351 3537 1355 3538
rect 1439 3542 1443 3543
rect 1439 3537 1443 3538
rect 1527 3542 1531 3543
rect 1527 3537 1531 3538
rect 1615 3542 1619 3543
rect 1615 3537 1619 3538
rect 1703 3542 1707 3543
rect 1703 3537 1707 3538
rect 1791 3542 1795 3543
rect 1791 3537 1795 3538
rect 1879 3542 1883 3543
rect 1879 3537 1883 3538
rect 2007 3542 2011 3543
rect 2007 3537 2011 3538
rect 2047 3542 2051 3543
rect 2047 3537 2051 3538
rect 2103 3542 2107 3543
rect 2103 3537 2107 3538
rect 2191 3542 2195 3543
rect 2191 3537 2195 3538
rect 2271 3542 2275 3543
rect 2271 3537 2275 3538
rect 2327 3542 2331 3543
rect 2327 3537 2331 3538
rect 2447 3542 2451 3543
rect 2447 3537 2451 3538
rect 2455 3542 2459 3543
rect 2455 3537 2459 3538
rect 2583 3542 2587 3543
rect 2583 3537 2587 3538
rect 2631 3542 2635 3543
rect 2631 3537 2635 3538
rect 2719 3542 2723 3543
rect 2719 3537 2723 3538
rect 2815 3542 2819 3543
rect 2815 3537 2819 3538
rect 2855 3542 2859 3543
rect 2855 3537 2859 3538
rect 2999 3542 3003 3543
rect 2999 3537 3003 3538
rect 3143 3542 3147 3543
rect 3143 3537 3147 3538
rect 3175 3542 3179 3543
rect 3175 3537 3179 3538
rect 3295 3542 3299 3543
rect 3295 3537 3299 3538
rect 3351 3542 3355 3543
rect 3351 3537 3355 3538
rect 3455 3542 3459 3543
rect 3455 3537 3459 3538
rect 3519 3542 3523 3543
rect 3519 3537 3523 3538
rect 3623 3542 3627 3543
rect 3623 3537 3627 3538
rect 3687 3542 3691 3543
rect 3687 3537 3691 3538
rect 3839 3542 3843 3543
rect 3839 3537 3843 3538
rect 3943 3542 3947 3543
rect 3943 3537 3947 3538
rect 112 3517 114 3537
rect 110 3516 116 3517
rect 160 3516 162 3537
rect 304 3516 306 3537
rect 464 3516 466 3537
rect 640 3516 642 3537
rect 816 3516 818 3537
rect 1000 3516 1002 3537
rect 1176 3516 1178 3537
rect 1352 3516 1354 3537
rect 1528 3516 1530 3537
rect 1704 3516 1706 3537
rect 1880 3516 1882 3537
rect 2008 3517 2010 3537
rect 2006 3516 2012 3517
rect 110 3512 111 3516
rect 115 3512 116 3516
rect 110 3511 116 3512
rect 158 3515 164 3516
rect 158 3511 159 3515
rect 163 3511 164 3515
rect 158 3510 164 3511
rect 302 3515 308 3516
rect 302 3511 303 3515
rect 307 3511 308 3515
rect 302 3510 308 3511
rect 462 3515 468 3516
rect 462 3511 463 3515
rect 467 3511 468 3515
rect 462 3510 468 3511
rect 638 3515 644 3516
rect 638 3511 639 3515
rect 643 3511 644 3515
rect 638 3510 644 3511
rect 814 3515 820 3516
rect 814 3511 815 3515
rect 819 3511 820 3515
rect 814 3510 820 3511
rect 998 3515 1004 3516
rect 998 3511 999 3515
rect 1003 3511 1004 3515
rect 998 3510 1004 3511
rect 1174 3515 1180 3516
rect 1174 3511 1175 3515
rect 1179 3511 1180 3515
rect 1174 3510 1180 3511
rect 1350 3515 1356 3516
rect 1350 3511 1351 3515
rect 1355 3511 1356 3515
rect 1350 3510 1356 3511
rect 1526 3515 1532 3516
rect 1526 3511 1527 3515
rect 1531 3511 1532 3515
rect 1526 3510 1532 3511
rect 1702 3515 1708 3516
rect 1702 3511 1703 3515
rect 1707 3511 1708 3515
rect 1702 3510 1708 3511
rect 1878 3515 1884 3516
rect 1878 3511 1879 3515
rect 1883 3511 1884 3515
rect 2006 3512 2007 3516
rect 2011 3512 2012 3516
rect 2006 3511 2012 3512
rect 1878 3510 1884 3511
rect 2048 3510 2050 3537
rect 2104 3513 2106 3537
rect 2272 3513 2274 3537
rect 2448 3513 2450 3537
rect 2632 3513 2634 3537
rect 2816 3513 2818 3537
rect 3000 3513 3002 3537
rect 3176 3513 3178 3537
rect 3352 3513 3354 3537
rect 3520 3513 3522 3537
rect 3688 3513 3690 3537
rect 3840 3513 3842 3537
rect 2102 3512 2108 3513
rect 2046 3509 2052 3510
rect 2046 3505 2047 3509
rect 2051 3505 2052 3509
rect 2102 3508 2103 3512
rect 2107 3508 2108 3512
rect 2102 3507 2108 3508
rect 2270 3512 2276 3513
rect 2270 3508 2271 3512
rect 2275 3508 2276 3512
rect 2270 3507 2276 3508
rect 2446 3512 2452 3513
rect 2446 3508 2447 3512
rect 2451 3508 2452 3512
rect 2446 3507 2452 3508
rect 2630 3512 2636 3513
rect 2630 3508 2631 3512
rect 2635 3508 2636 3512
rect 2630 3507 2636 3508
rect 2814 3512 2820 3513
rect 2814 3508 2815 3512
rect 2819 3508 2820 3512
rect 2814 3507 2820 3508
rect 2998 3512 3004 3513
rect 2998 3508 2999 3512
rect 3003 3508 3004 3512
rect 2998 3507 3004 3508
rect 3174 3512 3180 3513
rect 3174 3508 3175 3512
rect 3179 3508 3180 3512
rect 3174 3507 3180 3508
rect 3350 3512 3356 3513
rect 3350 3508 3351 3512
rect 3355 3508 3356 3512
rect 3350 3507 3356 3508
rect 3518 3512 3524 3513
rect 3518 3508 3519 3512
rect 3523 3508 3524 3512
rect 3518 3507 3524 3508
rect 3686 3512 3692 3513
rect 3686 3508 3687 3512
rect 3691 3508 3692 3512
rect 3686 3507 3692 3508
rect 3838 3512 3844 3513
rect 3838 3508 3839 3512
rect 3843 3508 3844 3512
rect 3944 3510 3946 3537
rect 3838 3507 3844 3508
rect 3942 3509 3948 3510
rect 2046 3504 2052 3505
rect 3942 3505 3943 3509
rect 3947 3505 3948 3509
rect 3942 3504 3948 3505
rect 110 3499 116 3500
rect 110 3495 111 3499
rect 115 3495 116 3499
rect 2006 3499 2012 3500
rect 110 3494 116 3495
rect 158 3496 164 3497
rect 112 3459 114 3494
rect 158 3492 159 3496
rect 163 3492 164 3496
rect 158 3491 164 3492
rect 302 3496 308 3497
rect 302 3492 303 3496
rect 307 3492 308 3496
rect 302 3491 308 3492
rect 462 3496 468 3497
rect 462 3492 463 3496
rect 467 3492 468 3496
rect 462 3491 468 3492
rect 638 3496 644 3497
rect 638 3492 639 3496
rect 643 3492 644 3496
rect 638 3491 644 3492
rect 814 3496 820 3497
rect 814 3492 815 3496
rect 819 3492 820 3496
rect 814 3491 820 3492
rect 998 3496 1004 3497
rect 998 3492 999 3496
rect 1003 3492 1004 3496
rect 998 3491 1004 3492
rect 1174 3496 1180 3497
rect 1174 3492 1175 3496
rect 1179 3492 1180 3496
rect 1174 3491 1180 3492
rect 1350 3496 1356 3497
rect 1350 3492 1351 3496
rect 1355 3492 1356 3496
rect 1350 3491 1356 3492
rect 1526 3496 1532 3497
rect 1526 3492 1527 3496
rect 1531 3492 1532 3496
rect 1526 3491 1532 3492
rect 1702 3496 1708 3497
rect 1702 3492 1703 3496
rect 1707 3492 1708 3496
rect 1702 3491 1708 3492
rect 1878 3496 1884 3497
rect 1878 3492 1879 3496
rect 1883 3492 1884 3496
rect 2006 3495 2007 3499
rect 2011 3495 2012 3499
rect 2006 3494 2012 3495
rect 1878 3491 1884 3492
rect 160 3459 162 3491
rect 304 3459 306 3491
rect 464 3459 466 3491
rect 640 3459 642 3491
rect 816 3459 818 3491
rect 1000 3459 1002 3491
rect 1176 3459 1178 3491
rect 1352 3459 1354 3491
rect 1528 3459 1530 3491
rect 1704 3459 1706 3491
rect 1880 3459 1882 3491
rect 2008 3459 2010 3494
rect 2102 3493 2108 3494
rect 2046 3492 2052 3493
rect 2046 3488 2047 3492
rect 2051 3488 2052 3492
rect 2102 3489 2103 3493
rect 2107 3489 2108 3493
rect 2102 3488 2108 3489
rect 2270 3493 2276 3494
rect 2270 3489 2271 3493
rect 2275 3489 2276 3493
rect 2270 3488 2276 3489
rect 2446 3493 2452 3494
rect 2446 3489 2447 3493
rect 2451 3489 2452 3493
rect 2446 3488 2452 3489
rect 2630 3493 2636 3494
rect 2630 3489 2631 3493
rect 2635 3489 2636 3493
rect 2630 3488 2636 3489
rect 2814 3493 2820 3494
rect 2814 3489 2815 3493
rect 2819 3489 2820 3493
rect 2814 3488 2820 3489
rect 2998 3493 3004 3494
rect 2998 3489 2999 3493
rect 3003 3489 3004 3493
rect 2998 3488 3004 3489
rect 3174 3493 3180 3494
rect 3174 3489 3175 3493
rect 3179 3489 3180 3493
rect 3174 3488 3180 3489
rect 3350 3493 3356 3494
rect 3350 3489 3351 3493
rect 3355 3489 3356 3493
rect 3350 3488 3356 3489
rect 3518 3493 3524 3494
rect 3518 3489 3519 3493
rect 3523 3489 3524 3493
rect 3518 3488 3524 3489
rect 3686 3493 3692 3494
rect 3686 3489 3687 3493
rect 3691 3489 3692 3493
rect 3686 3488 3692 3489
rect 3838 3493 3844 3494
rect 3838 3489 3839 3493
rect 3843 3489 3844 3493
rect 3838 3488 3844 3489
rect 3942 3492 3948 3493
rect 3942 3488 3943 3492
rect 3947 3488 3948 3492
rect 2046 3487 2052 3488
rect 2048 3463 2050 3487
rect 2104 3463 2106 3488
rect 2272 3463 2274 3488
rect 2448 3463 2450 3488
rect 2632 3463 2634 3488
rect 2816 3463 2818 3488
rect 3000 3463 3002 3488
rect 3176 3463 3178 3488
rect 3352 3463 3354 3488
rect 3520 3463 3522 3488
rect 3688 3463 3690 3488
rect 3840 3463 3842 3488
rect 3942 3487 3948 3488
rect 3944 3463 3946 3487
rect 2047 3462 2051 3463
rect 111 3458 115 3459
rect 111 3453 115 3454
rect 135 3458 139 3459
rect 135 3453 139 3454
rect 159 3458 163 3459
rect 159 3453 163 3454
rect 303 3458 307 3459
rect 303 3453 307 3454
rect 319 3458 323 3459
rect 319 3453 323 3454
rect 463 3458 467 3459
rect 463 3453 467 3454
rect 535 3458 539 3459
rect 535 3453 539 3454
rect 639 3458 643 3459
rect 639 3453 643 3454
rect 751 3458 755 3459
rect 751 3453 755 3454
rect 815 3458 819 3459
rect 815 3453 819 3454
rect 959 3458 963 3459
rect 959 3453 963 3454
rect 999 3458 1003 3459
rect 999 3453 1003 3454
rect 1159 3458 1163 3459
rect 1159 3453 1163 3454
rect 1175 3458 1179 3459
rect 1175 3453 1179 3454
rect 1351 3458 1355 3459
rect 1351 3453 1355 3454
rect 1527 3458 1531 3459
rect 1527 3453 1531 3454
rect 1535 3458 1539 3459
rect 1535 3453 1539 3454
rect 1703 3458 1707 3459
rect 1703 3453 1707 3454
rect 1719 3458 1723 3459
rect 1719 3453 1723 3454
rect 1879 3458 1883 3459
rect 1879 3453 1883 3454
rect 1903 3458 1907 3459
rect 1903 3453 1907 3454
rect 2007 3458 2011 3459
rect 2047 3457 2051 3458
rect 2103 3462 2107 3463
rect 2103 3457 2107 3458
rect 2127 3462 2131 3463
rect 2127 3457 2131 3458
rect 2271 3462 2275 3463
rect 2271 3457 2275 3458
rect 2311 3462 2315 3463
rect 2311 3457 2315 3458
rect 2447 3462 2451 3463
rect 2447 3457 2451 3458
rect 2495 3462 2499 3463
rect 2495 3457 2499 3458
rect 2631 3462 2635 3463
rect 2631 3457 2635 3458
rect 2679 3462 2683 3463
rect 2679 3457 2683 3458
rect 2815 3462 2819 3463
rect 2815 3457 2819 3458
rect 2863 3462 2867 3463
rect 2863 3457 2867 3458
rect 2999 3462 3003 3463
rect 2999 3457 3003 3458
rect 3047 3462 3051 3463
rect 3047 3457 3051 3458
rect 3175 3462 3179 3463
rect 3175 3457 3179 3458
rect 3223 3462 3227 3463
rect 3223 3457 3227 3458
rect 3351 3462 3355 3463
rect 3351 3457 3355 3458
rect 3407 3462 3411 3463
rect 3407 3457 3411 3458
rect 3519 3462 3523 3463
rect 3519 3457 3523 3458
rect 3591 3462 3595 3463
rect 3591 3457 3595 3458
rect 3687 3462 3691 3463
rect 3687 3457 3691 3458
rect 3775 3462 3779 3463
rect 3775 3457 3779 3458
rect 3839 3462 3843 3463
rect 3839 3457 3843 3458
rect 3943 3462 3947 3463
rect 3943 3457 3947 3458
rect 2007 3453 2011 3454
rect 112 3426 114 3453
rect 136 3429 138 3453
rect 320 3429 322 3453
rect 536 3429 538 3453
rect 752 3429 754 3453
rect 960 3429 962 3453
rect 1160 3429 1162 3453
rect 1352 3429 1354 3453
rect 1536 3429 1538 3453
rect 1720 3429 1722 3453
rect 1904 3429 1906 3453
rect 134 3428 140 3429
rect 110 3425 116 3426
rect 110 3421 111 3425
rect 115 3421 116 3425
rect 134 3424 135 3428
rect 139 3424 140 3428
rect 134 3423 140 3424
rect 318 3428 324 3429
rect 318 3424 319 3428
rect 323 3424 324 3428
rect 318 3423 324 3424
rect 534 3428 540 3429
rect 534 3424 535 3428
rect 539 3424 540 3428
rect 534 3423 540 3424
rect 750 3428 756 3429
rect 750 3424 751 3428
rect 755 3424 756 3428
rect 750 3423 756 3424
rect 958 3428 964 3429
rect 958 3424 959 3428
rect 963 3424 964 3428
rect 958 3423 964 3424
rect 1158 3428 1164 3429
rect 1158 3424 1159 3428
rect 1163 3424 1164 3428
rect 1158 3423 1164 3424
rect 1350 3428 1356 3429
rect 1350 3424 1351 3428
rect 1355 3424 1356 3428
rect 1350 3423 1356 3424
rect 1534 3428 1540 3429
rect 1534 3424 1535 3428
rect 1539 3424 1540 3428
rect 1534 3423 1540 3424
rect 1718 3428 1724 3429
rect 1718 3424 1719 3428
rect 1723 3424 1724 3428
rect 1718 3423 1724 3424
rect 1902 3428 1908 3429
rect 1902 3424 1903 3428
rect 1907 3424 1908 3428
rect 2008 3426 2010 3453
rect 2048 3437 2050 3457
rect 2046 3436 2052 3437
rect 2128 3436 2130 3457
rect 2312 3436 2314 3457
rect 2496 3436 2498 3457
rect 2680 3436 2682 3457
rect 2864 3436 2866 3457
rect 3048 3436 3050 3457
rect 3224 3436 3226 3457
rect 3408 3436 3410 3457
rect 3592 3436 3594 3457
rect 3776 3436 3778 3457
rect 3944 3437 3946 3457
rect 3942 3436 3948 3437
rect 2046 3432 2047 3436
rect 2051 3432 2052 3436
rect 2046 3431 2052 3432
rect 2126 3435 2132 3436
rect 2126 3431 2127 3435
rect 2131 3431 2132 3435
rect 2126 3430 2132 3431
rect 2310 3435 2316 3436
rect 2310 3431 2311 3435
rect 2315 3431 2316 3435
rect 2310 3430 2316 3431
rect 2494 3435 2500 3436
rect 2494 3431 2495 3435
rect 2499 3431 2500 3435
rect 2494 3430 2500 3431
rect 2678 3435 2684 3436
rect 2678 3431 2679 3435
rect 2683 3431 2684 3435
rect 2678 3430 2684 3431
rect 2862 3435 2868 3436
rect 2862 3431 2863 3435
rect 2867 3431 2868 3435
rect 2862 3430 2868 3431
rect 3046 3435 3052 3436
rect 3046 3431 3047 3435
rect 3051 3431 3052 3435
rect 3046 3430 3052 3431
rect 3222 3435 3228 3436
rect 3222 3431 3223 3435
rect 3227 3431 3228 3435
rect 3222 3430 3228 3431
rect 3406 3435 3412 3436
rect 3406 3431 3407 3435
rect 3411 3431 3412 3435
rect 3406 3430 3412 3431
rect 3590 3435 3596 3436
rect 3590 3431 3591 3435
rect 3595 3431 3596 3435
rect 3590 3430 3596 3431
rect 3774 3435 3780 3436
rect 3774 3431 3775 3435
rect 3779 3431 3780 3435
rect 3942 3432 3943 3436
rect 3947 3432 3948 3436
rect 3942 3431 3948 3432
rect 3774 3430 3780 3431
rect 1902 3423 1908 3424
rect 2006 3425 2012 3426
rect 110 3420 116 3421
rect 2006 3421 2007 3425
rect 2011 3421 2012 3425
rect 2006 3420 2012 3421
rect 2046 3419 2052 3420
rect 2046 3415 2047 3419
rect 2051 3415 2052 3419
rect 3942 3419 3948 3420
rect 2046 3414 2052 3415
rect 2126 3416 2132 3417
rect 134 3409 140 3410
rect 110 3408 116 3409
rect 110 3404 111 3408
rect 115 3404 116 3408
rect 134 3405 135 3409
rect 139 3405 140 3409
rect 134 3404 140 3405
rect 318 3409 324 3410
rect 318 3405 319 3409
rect 323 3405 324 3409
rect 318 3404 324 3405
rect 534 3409 540 3410
rect 534 3405 535 3409
rect 539 3405 540 3409
rect 534 3404 540 3405
rect 750 3409 756 3410
rect 750 3405 751 3409
rect 755 3405 756 3409
rect 750 3404 756 3405
rect 958 3409 964 3410
rect 958 3405 959 3409
rect 963 3405 964 3409
rect 958 3404 964 3405
rect 1158 3409 1164 3410
rect 1158 3405 1159 3409
rect 1163 3405 1164 3409
rect 1158 3404 1164 3405
rect 1350 3409 1356 3410
rect 1350 3405 1351 3409
rect 1355 3405 1356 3409
rect 1350 3404 1356 3405
rect 1534 3409 1540 3410
rect 1534 3405 1535 3409
rect 1539 3405 1540 3409
rect 1534 3404 1540 3405
rect 1718 3409 1724 3410
rect 1718 3405 1719 3409
rect 1723 3405 1724 3409
rect 1718 3404 1724 3405
rect 1902 3409 1908 3410
rect 1902 3405 1903 3409
rect 1907 3405 1908 3409
rect 1902 3404 1908 3405
rect 2006 3408 2012 3409
rect 2006 3404 2007 3408
rect 2011 3404 2012 3408
rect 110 3403 116 3404
rect 112 3383 114 3403
rect 136 3383 138 3404
rect 320 3383 322 3404
rect 536 3383 538 3404
rect 752 3383 754 3404
rect 960 3383 962 3404
rect 1160 3383 1162 3404
rect 1352 3383 1354 3404
rect 1536 3383 1538 3404
rect 1720 3383 1722 3404
rect 1904 3383 1906 3404
rect 2006 3403 2012 3404
rect 2008 3383 2010 3403
rect 111 3382 115 3383
rect 111 3377 115 3378
rect 135 3382 139 3383
rect 135 3377 139 3378
rect 231 3382 235 3383
rect 231 3377 235 3378
rect 319 3382 323 3383
rect 319 3377 323 3378
rect 375 3382 379 3383
rect 375 3377 379 3378
rect 535 3382 539 3383
rect 535 3377 539 3378
rect 703 3382 707 3383
rect 703 3377 707 3378
rect 751 3382 755 3383
rect 751 3377 755 3378
rect 871 3382 875 3383
rect 871 3377 875 3378
rect 959 3382 963 3383
rect 959 3377 963 3378
rect 1047 3382 1051 3383
rect 1047 3377 1051 3378
rect 1159 3382 1163 3383
rect 1159 3377 1163 3378
rect 1215 3382 1219 3383
rect 1215 3377 1219 3378
rect 1351 3382 1355 3383
rect 1351 3377 1355 3378
rect 1383 3382 1387 3383
rect 1383 3377 1387 3378
rect 1535 3382 1539 3383
rect 1535 3377 1539 3378
rect 1543 3382 1547 3383
rect 1543 3377 1547 3378
rect 1703 3382 1707 3383
rect 1703 3377 1707 3378
rect 1719 3382 1723 3383
rect 1719 3377 1723 3378
rect 1871 3382 1875 3383
rect 1871 3377 1875 3378
rect 1903 3382 1907 3383
rect 1903 3377 1907 3378
rect 2007 3382 2011 3383
rect 2007 3377 2011 3378
rect 112 3357 114 3377
rect 110 3356 116 3357
rect 136 3356 138 3377
rect 232 3356 234 3377
rect 376 3356 378 3377
rect 536 3356 538 3377
rect 704 3356 706 3377
rect 872 3356 874 3377
rect 1048 3356 1050 3377
rect 1216 3356 1218 3377
rect 1384 3356 1386 3377
rect 1544 3356 1546 3377
rect 1704 3356 1706 3377
rect 1872 3356 1874 3377
rect 2008 3357 2010 3377
rect 2048 3371 2050 3414
rect 2126 3412 2127 3416
rect 2131 3412 2132 3416
rect 2126 3411 2132 3412
rect 2310 3416 2316 3417
rect 2310 3412 2311 3416
rect 2315 3412 2316 3416
rect 2310 3411 2316 3412
rect 2494 3416 2500 3417
rect 2494 3412 2495 3416
rect 2499 3412 2500 3416
rect 2494 3411 2500 3412
rect 2678 3416 2684 3417
rect 2678 3412 2679 3416
rect 2683 3412 2684 3416
rect 2678 3411 2684 3412
rect 2862 3416 2868 3417
rect 2862 3412 2863 3416
rect 2867 3412 2868 3416
rect 2862 3411 2868 3412
rect 3046 3416 3052 3417
rect 3046 3412 3047 3416
rect 3051 3412 3052 3416
rect 3046 3411 3052 3412
rect 3222 3416 3228 3417
rect 3222 3412 3223 3416
rect 3227 3412 3228 3416
rect 3222 3411 3228 3412
rect 3406 3416 3412 3417
rect 3406 3412 3407 3416
rect 3411 3412 3412 3416
rect 3406 3411 3412 3412
rect 3590 3416 3596 3417
rect 3590 3412 3591 3416
rect 3595 3412 3596 3416
rect 3590 3411 3596 3412
rect 3774 3416 3780 3417
rect 3774 3412 3775 3416
rect 3779 3412 3780 3416
rect 3942 3415 3943 3419
rect 3947 3415 3948 3419
rect 3942 3414 3948 3415
rect 3774 3411 3780 3412
rect 2128 3371 2130 3411
rect 2312 3371 2314 3411
rect 2496 3371 2498 3411
rect 2680 3371 2682 3411
rect 2864 3371 2866 3411
rect 3048 3371 3050 3411
rect 3224 3371 3226 3411
rect 3408 3371 3410 3411
rect 3592 3371 3594 3411
rect 3776 3371 3778 3411
rect 3944 3371 3946 3414
rect 2047 3370 2051 3371
rect 2047 3365 2051 3366
rect 2071 3370 2075 3371
rect 2071 3365 2075 3366
rect 2127 3370 2131 3371
rect 2127 3365 2131 3366
rect 2215 3370 2219 3371
rect 2215 3365 2219 3366
rect 2311 3370 2315 3371
rect 2311 3365 2315 3366
rect 2359 3370 2363 3371
rect 2359 3365 2363 3366
rect 2495 3370 2499 3371
rect 2495 3365 2499 3366
rect 2511 3370 2515 3371
rect 2511 3365 2515 3366
rect 2655 3370 2659 3371
rect 2655 3365 2659 3366
rect 2679 3370 2683 3371
rect 2679 3365 2683 3366
rect 2799 3370 2803 3371
rect 2799 3365 2803 3366
rect 2863 3370 2867 3371
rect 2863 3365 2867 3366
rect 2935 3370 2939 3371
rect 2935 3365 2939 3366
rect 3047 3370 3051 3371
rect 3047 3365 3051 3366
rect 3079 3370 3083 3371
rect 3079 3365 3083 3366
rect 3223 3370 3227 3371
rect 3223 3365 3227 3366
rect 3375 3370 3379 3371
rect 3375 3365 3379 3366
rect 3407 3370 3411 3371
rect 3407 3365 3411 3366
rect 3535 3370 3539 3371
rect 3535 3365 3539 3366
rect 3591 3370 3595 3371
rect 3591 3365 3595 3366
rect 3695 3370 3699 3371
rect 3695 3365 3699 3366
rect 3775 3370 3779 3371
rect 3775 3365 3779 3366
rect 3839 3370 3843 3371
rect 3839 3365 3843 3366
rect 3943 3370 3947 3371
rect 3943 3365 3947 3366
rect 2006 3356 2012 3357
rect 110 3352 111 3356
rect 115 3352 116 3356
rect 110 3351 116 3352
rect 134 3355 140 3356
rect 134 3351 135 3355
rect 139 3351 140 3355
rect 134 3350 140 3351
rect 230 3355 236 3356
rect 230 3351 231 3355
rect 235 3351 236 3355
rect 230 3350 236 3351
rect 374 3355 380 3356
rect 374 3351 375 3355
rect 379 3351 380 3355
rect 374 3350 380 3351
rect 534 3355 540 3356
rect 534 3351 535 3355
rect 539 3351 540 3355
rect 534 3350 540 3351
rect 702 3355 708 3356
rect 702 3351 703 3355
rect 707 3351 708 3355
rect 702 3350 708 3351
rect 870 3355 876 3356
rect 870 3351 871 3355
rect 875 3351 876 3355
rect 870 3350 876 3351
rect 1046 3355 1052 3356
rect 1046 3351 1047 3355
rect 1051 3351 1052 3355
rect 1046 3350 1052 3351
rect 1214 3355 1220 3356
rect 1214 3351 1215 3355
rect 1219 3351 1220 3355
rect 1214 3350 1220 3351
rect 1382 3355 1388 3356
rect 1382 3351 1383 3355
rect 1387 3351 1388 3355
rect 1382 3350 1388 3351
rect 1542 3355 1548 3356
rect 1542 3351 1543 3355
rect 1547 3351 1548 3355
rect 1542 3350 1548 3351
rect 1702 3355 1708 3356
rect 1702 3351 1703 3355
rect 1707 3351 1708 3355
rect 1702 3350 1708 3351
rect 1870 3355 1876 3356
rect 1870 3351 1871 3355
rect 1875 3351 1876 3355
rect 2006 3352 2007 3356
rect 2011 3352 2012 3356
rect 2006 3351 2012 3352
rect 1870 3350 1876 3351
rect 110 3339 116 3340
rect 110 3335 111 3339
rect 115 3335 116 3339
rect 2006 3339 2012 3340
rect 110 3334 116 3335
rect 134 3336 140 3337
rect 112 3307 114 3334
rect 134 3332 135 3336
rect 139 3332 140 3336
rect 134 3331 140 3332
rect 230 3336 236 3337
rect 230 3332 231 3336
rect 235 3332 236 3336
rect 230 3331 236 3332
rect 374 3336 380 3337
rect 374 3332 375 3336
rect 379 3332 380 3336
rect 374 3331 380 3332
rect 534 3336 540 3337
rect 534 3332 535 3336
rect 539 3332 540 3336
rect 534 3331 540 3332
rect 702 3336 708 3337
rect 702 3332 703 3336
rect 707 3332 708 3336
rect 702 3331 708 3332
rect 870 3336 876 3337
rect 870 3332 871 3336
rect 875 3332 876 3336
rect 870 3331 876 3332
rect 1046 3336 1052 3337
rect 1046 3332 1047 3336
rect 1051 3332 1052 3336
rect 1046 3331 1052 3332
rect 1214 3336 1220 3337
rect 1214 3332 1215 3336
rect 1219 3332 1220 3336
rect 1214 3331 1220 3332
rect 1382 3336 1388 3337
rect 1382 3332 1383 3336
rect 1387 3332 1388 3336
rect 1382 3331 1388 3332
rect 1542 3336 1548 3337
rect 1542 3332 1543 3336
rect 1547 3332 1548 3336
rect 1542 3331 1548 3332
rect 1702 3336 1708 3337
rect 1702 3332 1703 3336
rect 1707 3332 1708 3336
rect 1702 3331 1708 3332
rect 1870 3336 1876 3337
rect 1870 3332 1871 3336
rect 1875 3332 1876 3336
rect 2006 3335 2007 3339
rect 2011 3335 2012 3339
rect 2048 3338 2050 3365
rect 2072 3341 2074 3365
rect 2216 3341 2218 3365
rect 2360 3341 2362 3365
rect 2512 3341 2514 3365
rect 2656 3341 2658 3365
rect 2800 3341 2802 3365
rect 2936 3341 2938 3365
rect 3080 3341 3082 3365
rect 3224 3341 3226 3365
rect 3376 3341 3378 3365
rect 3536 3341 3538 3365
rect 3696 3341 3698 3365
rect 3840 3341 3842 3365
rect 2070 3340 2076 3341
rect 2006 3334 2012 3335
rect 2046 3337 2052 3338
rect 1870 3331 1876 3332
rect 136 3307 138 3331
rect 232 3307 234 3331
rect 376 3307 378 3331
rect 536 3307 538 3331
rect 704 3307 706 3331
rect 872 3307 874 3331
rect 1048 3307 1050 3331
rect 1216 3307 1218 3331
rect 1384 3307 1386 3331
rect 1544 3307 1546 3331
rect 1704 3307 1706 3331
rect 1872 3307 1874 3331
rect 2008 3307 2010 3334
rect 2046 3333 2047 3337
rect 2051 3333 2052 3337
rect 2070 3336 2071 3340
rect 2075 3336 2076 3340
rect 2070 3335 2076 3336
rect 2214 3340 2220 3341
rect 2214 3336 2215 3340
rect 2219 3336 2220 3340
rect 2214 3335 2220 3336
rect 2358 3340 2364 3341
rect 2358 3336 2359 3340
rect 2363 3336 2364 3340
rect 2358 3335 2364 3336
rect 2510 3340 2516 3341
rect 2510 3336 2511 3340
rect 2515 3336 2516 3340
rect 2510 3335 2516 3336
rect 2654 3340 2660 3341
rect 2654 3336 2655 3340
rect 2659 3336 2660 3340
rect 2654 3335 2660 3336
rect 2798 3340 2804 3341
rect 2798 3336 2799 3340
rect 2803 3336 2804 3340
rect 2798 3335 2804 3336
rect 2934 3340 2940 3341
rect 2934 3336 2935 3340
rect 2939 3336 2940 3340
rect 2934 3335 2940 3336
rect 3078 3340 3084 3341
rect 3078 3336 3079 3340
rect 3083 3336 3084 3340
rect 3078 3335 3084 3336
rect 3222 3340 3228 3341
rect 3222 3336 3223 3340
rect 3227 3336 3228 3340
rect 3222 3335 3228 3336
rect 3374 3340 3380 3341
rect 3374 3336 3375 3340
rect 3379 3336 3380 3340
rect 3374 3335 3380 3336
rect 3534 3340 3540 3341
rect 3534 3336 3535 3340
rect 3539 3336 3540 3340
rect 3534 3335 3540 3336
rect 3694 3340 3700 3341
rect 3694 3336 3695 3340
rect 3699 3336 3700 3340
rect 3694 3335 3700 3336
rect 3838 3340 3844 3341
rect 3838 3336 3839 3340
rect 3843 3336 3844 3340
rect 3944 3338 3946 3365
rect 3838 3335 3844 3336
rect 3942 3337 3948 3338
rect 2046 3332 2052 3333
rect 3942 3333 3943 3337
rect 3947 3333 3948 3337
rect 3942 3332 3948 3333
rect 2070 3321 2076 3322
rect 2046 3320 2052 3321
rect 2046 3316 2047 3320
rect 2051 3316 2052 3320
rect 2070 3317 2071 3321
rect 2075 3317 2076 3321
rect 2070 3316 2076 3317
rect 2214 3321 2220 3322
rect 2214 3317 2215 3321
rect 2219 3317 2220 3321
rect 2214 3316 2220 3317
rect 2358 3321 2364 3322
rect 2358 3317 2359 3321
rect 2363 3317 2364 3321
rect 2358 3316 2364 3317
rect 2510 3321 2516 3322
rect 2510 3317 2511 3321
rect 2515 3317 2516 3321
rect 2510 3316 2516 3317
rect 2654 3321 2660 3322
rect 2654 3317 2655 3321
rect 2659 3317 2660 3321
rect 2654 3316 2660 3317
rect 2798 3321 2804 3322
rect 2798 3317 2799 3321
rect 2803 3317 2804 3321
rect 2798 3316 2804 3317
rect 2934 3321 2940 3322
rect 2934 3317 2935 3321
rect 2939 3317 2940 3321
rect 2934 3316 2940 3317
rect 3078 3321 3084 3322
rect 3078 3317 3079 3321
rect 3083 3317 3084 3321
rect 3078 3316 3084 3317
rect 3222 3321 3228 3322
rect 3222 3317 3223 3321
rect 3227 3317 3228 3321
rect 3222 3316 3228 3317
rect 3374 3321 3380 3322
rect 3374 3317 3375 3321
rect 3379 3317 3380 3321
rect 3374 3316 3380 3317
rect 3534 3321 3540 3322
rect 3534 3317 3535 3321
rect 3539 3317 3540 3321
rect 3534 3316 3540 3317
rect 3694 3321 3700 3322
rect 3694 3317 3695 3321
rect 3699 3317 3700 3321
rect 3694 3316 3700 3317
rect 3838 3321 3844 3322
rect 3838 3317 3839 3321
rect 3843 3317 3844 3321
rect 3838 3316 3844 3317
rect 3942 3320 3948 3321
rect 3942 3316 3943 3320
rect 3947 3316 3948 3320
rect 2046 3315 2052 3316
rect 111 3306 115 3307
rect 111 3301 115 3302
rect 135 3306 139 3307
rect 135 3301 139 3302
rect 231 3306 235 3307
rect 231 3301 235 3302
rect 279 3306 283 3307
rect 279 3301 283 3302
rect 375 3306 379 3307
rect 375 3301 379 3302
rect 463 3306 467 3307
rect 463 3301 467 3302
rect 535 3306 539 3307
rect 535 3301 539 3302
rect 663 3306 667 3307
rect 663 3301 667 3302
rect 703 3306 707 3307
rect 703 3301 707 3302
rect 871 3306 875 3307
rect 871 3301 875 3302
rect 1047 3306 1051 3307
rect 1047 3301 1051 3302
rect 1079 3306 1083 3307
rect 1079 3301 1083 3302
rect 1215 3306 1219 3307
rect 1215 3301 1219 3302
rect 1295 3306 1299 3307
rect 1295 3301 1299 3302
rect 1383 3306 1387 3307
rect 1383 3301 1387 3302
rect 1519 3306 1523 3307
rect 1519 3301 1523 3302
rect 1543 3306 1547 3307
rect 1543 3301 1547 3302
rect 1703 3306 1707 3307
rect 1703 3301 1707 3302
rect 1743 3306 1747 3307
rect 1743 3301 1747 3302
rect 1871 3306 1875 3307
rect 1871 3301 1875 3302
rect 2007 3306 2011 3307
rect 2007 3301 2011 3302
rect 112 3274 114 3301
rect 136 3277 138 3301
rect 280 3277 282 3301
rect 464 3277 466 3301
rect 664 3277 666 3301
rect 872 3277 874 3301
rect 1080 3277 1082 3301
rect 1296 3277 1298 3301
rect 1520 3277 1522 3301
rect 1744 3277 1746 3301
rect 134 3276 140 3277
rect 110 3273 116 3274
rect 110 3269 111 3273
rect 115 3269 116 3273
rect 134 3272 135 3276
rect 139 3272 140 3276
rect 134 3271 140 3272
rect 278 3276 284 3277
rect 278 3272 279 3276
rect 283 3272 284 3276
rect 278 3271 284 3272
rect 462 3276 468 3277
rect 462 3272 463 3276
rect 467 3272 468 3276
rect 462 3271 468 3272
rect 662 3276 668 3277
rect 662 3272 663 3276
rect 667 3272 668 3276
rect 662 3271 668 3272
rect 870 3276 876 3277
rect 870 3272 871 3276
rect 875 3272 876 3276
rect 870 3271 876 3272
rect 1078 3276 1084 3277
rect 1078 3272 1079 3276
rect 1083 3272 1084 3276
rect 1078 3271 1084 3272
rect 1294 3276 1300 3277
rect 1294 3272 1295 3276
rect 1299 3272 1300 3276
rect 1294 3271 1300 3272
rect 1518 3276 1524 3277
rect 1518 3272 1519 3276
rect 1523 3272 1524 3276
rect 1518 3271 1524 3272
rect 1742 3276 1748 3277
rect 1742 3272 1743 3276
rect 1747 3272 1748 3276
rect 2008 3274 2010 3301
rect 2048 3287 2050 3315
rect 2072 3287 2074 3316
rect 2216 3287 2218 3316
rect 2360 3287 2362 3316
rect 2512 3287 2514 3316
rect 2656 3287 2658 3316
rect 2800 3287 2802 3316
rect 2936 3287 2938 3316
rect 3080 3287 3082 3316
rect 3224 3287 3226 3316
rect 3376 3287 3378 3316
rect 3536 3287 3538 3316
rect 3696 3287 3698 3316
rect 3840 3287 3842 3316
rect 3942 3315 3948 3316
rect 3944 3287 3946 3315
rect 2047 3286 2051 3287
rect 2047 3281 2051 3282
rect 2071 3286 2075 3287
rect 2071 3281 2075 3282
rect 2111 3286 2115 3287
rect 2111 3281 2115 3282
rect 2215 3286 2219 3287
rect 2215 3281 2219 3282
rect 2247 3286 2251 3287
rect 2247 3281 2251 3282
rect 2359 3286 2363 3287
rect 2359 3281 2363 3282
rect 2399 3286 2403 3287
rect 2399 3281 2403 3282
rect 2511 3286 2515 3287
rect 2511 3281 2515 3282
rect 2575 3286 2579 3287
rect 2575 3281 2579 3282
rect 2655 3286 2659 3287
rect 2655 3281 2659 3282
rect 2783 3286 2787 3287
rect 2783 3281 2787 3282
rect 2799 3286 2803 3287
rect 2799 3281 2803 3282
rect 2935 3286 2939 3287
rect 2935 3281 2939 3282
rect 3015 3286 3019 3287
rect 3015 3281 3019 3282
rect 3079 3286 3083 3287
rect 3079 3281 3083 3282
rect 3223 3286 3227 3287
rect 3223 3281 3227 3282
rect 3263 3286 3267 3287
rect 3263 3281 3267 3282
rect 3375 3286 3379 3287
rect 3375 3281 3379 3282
rect 3527 3286 3531 3287
rect 3527 3281 3531 3282
rect 3535 3286 3539 3287
rect 3535 3281 3539 3282
rect 3695 3286 3699 3287
rect 3695 3281 3699 3282
rect 3791 3286 3795 3287
rect 3791 3281 3795 3282
rect 3839 3286 3843 3287
rect 3839 3281 3843 3282
rect 3943 3286 3947 3287
rect 3943 3281 3947 3282
rect 1742 3271 1748 3272
rect 2006 3273 2012 3274
rect 110 3268 116 3269
rect 2006 3269 2007 3273
rect 2011 3269 2012 3273
rect 2006 3268 2012 3269
rect 2048 3261 2050 3281
rect 2046 3260 2052 3261
rect 2112 3260 2114 3281
rect 2248 3260 2250 3281
rect 2400 3260 2402 3281
rect 2576 3260 2578 3281
rect 2784 3260 2786 3281
rect 3016 3260 3018 3281
rect 3264 3260 3266 3281
rect 3528 3260 3530 3281
rect 3792 3260 3794 3281
rect 3944 3261 3946 3281
rect 3942 3260 3948 3261
rect 134 3257 140 3258
rect 110 3256 116 3257
rect 110 3252 111 3256
rect 115 3252 116 3256
rect 134 3253 135 3257
rect 139 3253 140 3257
rect 134 3252 140 3253
rect 278 3257 284 3258
rect 278 3253 279 3257
rect 283 3253 284 3257
rect 278 3252 284 3253
rect 462 3257 468 3258
rect 462 3253 463 3257
rect 467 3253 468 3257
rect 462 3252 468 3253
rect 662 3257 668 3258
rect 662 3253 663 3257
rect 667 3253 668 3257
rect 662 3252 668 3253
rect 870 3257 876 3258
rect 870 3253 871 3257
rect 875 3253 876 3257
rect 870 3252 876 3253
rect 1078 3257 1084 3258
rect 1078 3253 1079 3257
rect 1083 3253 1084 3257
rect 1078 3252 1084 3253
rect 1294 3257 1300 3258
rect 1294 3253 1295 3257
rect 1299 3253 1300 3257
rect 1294 3252 1300 3253
rect 1518 3257 1524 3258
rect 1518 3253 1519 3257
rect 1523 3253 1524 3257
rect 1518 3252 1524 3253
rect 1742 3257 1748 3258
rect 1742 3253 1743 3257
rect 1747 3253 1748 3257
rect 1742 3252 1748 3253
rect 2006 3256 2012 3257
rect 2006 3252 2007 3256
rect 2011 3252 2012 3256
rect 2046 3256 2047 3260
rect 2051 3256 2052 3260
rect 2046 3255 2052 3256
rect 2110 3259 2116 3260
rect 2110 3255 2111 3259
rect 2115 3255 2116 3259
rect 2110 3254 2116 3255
rect 2246 3259 2252 3260
rect 2246 3255 2247 3259
rect 2251 3255 2252 3259
rect 2246 3254 2252 3255
rect 2398 3259 2404 3260
rect 2398 3255 2399 3259
rect 2403 3255 2404 3259
rect 2398 3254 2404 3255
rect 2574 3259 2580 3260
rect 2574 3255 2575 3259
rect 2579 3255 2580 3259
rect 2574 3254 2580 3255
rect 2782 3259 2788 3260
rect 2782 3255 2783 3259
rect 2787 3255 2788 3259
rect 2782 3254 2788 3255
rect 3014 3259 3020 3260
rect 3014 3255 3015 3259
rect 3019 3255 3020 3259
rect 3014 3254 3020 3255
rect 3262 3259 3268 3260
rect 3262 3255 3263 3259
rect 3267 3255 3268 3259
rect 3262 3254 3268 3255
rect 3526 3259 3532 3260
rect 3526 3255 3527 3259
rect 3531 3255 3532 3259
rect 3526 3254 3532 3255
rect 3790 3259 3796 3260
rect 3790 3255 3791 3259
rect 3795 3255 3796 3259
rect 3942 3256 3943 3260
rect 3947 3256 3948 3260
rect 3942 3255 3948 3256
rect 3790 3254 3796 3255
rect 110 3251 116 3252
rect 112 3231 114 3251
rect 136 3231 138 3252
rect 280 3231 282 3252
rect 464 3231 466 3252
rect 664 3231 666 3252
rect 872 3231 874 3252
rect 1080 3231 1082 3252
rect 1296 3231 1298 3252
rect 1520 3231 1522 3252
rect 1744 3231 1746 3252
rect 2006 3251 2012 3252
rect 2008 3231 2010 3251
rect 2046 3243 2052 3244
rect 2046 3239 2047 3243
rect 2051 3239 2052 3243
rect 3942 3243 3948 3244
rect 2046 3238 2052 3239
rect 2110 3240 2116 3241
rect 111 3230 115 3231
rect 111 3225 115 3226
rect 135 3230 139 3231
rect 135 3225 139 3226
rect 279 3230 283 3231
rect 279 3225 283 3226
rect 287 3230 291 3231
rect 287 3225 291 3226
rect 447 3230 451 3231
rect 447 3225 451 3226
rect 463 3230 467 3231
rect 463 3225 467 3226
rect 615 3230 619 3231
rect 615 3225 619 3226
rect 663 3230 667 3231
rect 663 3225 667 3226
rect 791 3230 795 3231
rect 791 3225 795 3226
rect 871 3230 875 3231
rect 871 3225 875 3226
rect 967 3230 971 3231
rect 967 3225 971 3226
rect 1079 3230 1083 3231
rect 1079 3225 1083 3226
rect 1143 3230 1147 3231
rect 1143 3225 1147 3226
rect 1295 3230 1299 3231
rect 1295 3225 1299 3226
rect 1327 3230 1331 3231
rect 1327 3225 1331 3226
rect 1511 3230 1515 3231
rect 1511 3225 1515 3226
rect 1519 3230 1523 3231
rect 1519 3225 1523 3226
rect 1695 3230 1699 3231
rect 1695 3225 1699 3226
rect 1743 3230 1747 3231
rect 1743 3225 1747 3226
rect 2007 3230 2011 3231
rect 2007 3225 2011 3226
rect 112 3205 114 3225
rect 110 3204 116 3205
rect 136 3204 138 3225
rect 288 3204 290 3225
rect 448 3204 450 3225
rect 616 3204 618 3225
rect 792 3204 794 3225
rect 968 3204 970 3225
rect 1144 3204 1146 3225
rect 1328 3204 1330 3225
rect 1512 3204 1514 3225
rect 1696 3204 1698 3225
rect 2008 3205 2010 3225
rect 2048 3211 2050 3238
rect 2110 3236 2111 3240
rect 2115 3236 2116 3240
rect 2110 3235 2116 3236
rect 2246 3240 2252 3241
rect 2246 3236 2247 3240
rect 2251 3236 2252 3240
rect 2246 3235 2252 3236
rect 2398 3240 2404 3241
rect 2398 3236 2399 3240
rect 2403 3236 2404 3240
rect 2398 3235 2404 3236
rect 2574 3240 2580 3241
rect 2574 3236 2575 3240
rect 2579 3236 2580 3240
rect 2574 3235 2580 3236
rect 2782 3240 2788 3241
rect 2782 3236 2783 3240
rect 2787 3236 2788 3240
rect 2782 3235 2788 3236
rect 3014 3240 3020 3241
rect 3014 3236 3015 3240
rect 3019 3236 3020 3240
rect 3014 3235 3020 3236
rect 3262 3240 3268 3241
rect 3262 3236 3263 3240
rect 3267 3236 3268 3240
rect 3262 3235 3268 3236
rect 3526 3240 3532 3241
rect 3526 3236 3527 3240
rect 3531 3236 3532 3240
rect 3526 3235 3532 3236
rect 3790 3240 3796 3241
rect 3790 3236 3791 3240
rect 3795 3236 3796 3240
rect 3942 3239 3943 3243
rect 3947 3239 3948 3243
rect 3942 3238 3948 3239
rect 3790 3235 3796 3236
rect 2112 3211 2114 3235
rect 2248 3211 2250 3235
rect 2400 3211 2402 3235
rect 2576 3211 2578 3235
rect 2784 3211 2786 3235
rect 3016 3211 3018 3235
rect 3264 3211 3266 3235
rect 3528 3211 3530 3235
rect 3792 3211 3794 3235
rect 3944 3211 3946 3238
rect 2047 3210 2051 3211
rect 2047 3205 2051 3206
rect 2071 3210 2075 3211
rect 2071 3205 2075 3206
rect 2111 3210 2115 3211
rect 2111 3205 2115 3206
rect 2167 3210 2171 3211
rect 2167 3205 2171 3206
rect 2247 3210 2251 3211
rect 2247 3205 2251 3206
rect 2263 3210 2267 3211
rect 2263 3205 2267 3206
rect 2359 3210 2363 3211
rect 2359 3205 2363 3206
rect 2399 3210 2403 3211
rect 2399 3205 2403 3206
rect 2455 3210 2459 3211
rect 2455 3205 2459 3206
rect 2551 3210 2555 3211
rect 2551 3205 2555 3206
rect 2575 3210 2579 3211
rect 2575 3205 2579 3206
rect 2647 3210 2651 3211
rect 2647 3205 2651 3206
rect 2743 3210 2747 3211
rect 2743 3205 2747 3206
rect 2783 3210 2787 3211
rect 2783 3205 2787 3206
rect 2839 3210 2843 3211
rect 2839 3205 2843 3206
rect 2935 3210 2939 3211
rect 2935 3205 2939 3206
rect 3015 3210 3019 3211
rect 3015 3205 3019 3206
rect 3031 3210 3035 3211
rect 3031 3205 3035 3206
rect 3127 3210 3131 3211
rect 3127 3205 3131 3206
rect 3223 3210 3227 3211
rect 3223 3205 3227 3206
rect 3263 3210 3267 3211
rect 3263 3205 3267 3206
rect 3319 3210 3323 3211
rect 3319 3205 3323 3206
rect 3439 3210 3443 3211
rect 3439 3205 3443 3206
rect 3527 3210 3531 3211
rect 3527 3205 3531 3206
rect 3575 3210 3579 3211
rect 3575 3205 3579 3206
rect 3719 3210 3723 3211
rect 3719 3205 3723 3206
rect 3791 3210 3795 3211
rect 3791 3205 3795 3206
rect 3839 3210 3843 3211
rect 3839 3205 3843 3206
rect 3943 3210 3947 3211
rect 3943 3205 3947 3206
rect 2006 3204 2012 3205
rect 110 3200 111 3204
rect 115 3200 116 3204
rect 110 3199 116 3200
rect 134 3203 140 3204
rect 134 3199 135 3203
rect 139 3199 140 3203
rect 134 3198 140 3199
rect 286 3203 292 3204
rect 286 3199 287 3203
rect 291 3199 292 3203
rect 286 3198 292 3199
rect 446 3203 452 3204
rect 446 3199 447 3203
rect 451 3199 452 3203
rect 446 3198 452 3199
rect 614 3203 620 3204
rect 614 3199 615 3203
rect 619 3199 620 3203
rect 614 3198 620 3199
rect 790 3203 796 3204
rect 790 3199 791 3203
rect 795 3199 796 3203
rect 790 3198 796 3199
rect 966 3203 972 3204
rect 966 3199 967 3203
rect 971 3199 972 3203
rect 966 3198 972 3199
rect 1142 3203 1148 3204
rect 1142 3199 1143 3203
rect 1147 3199 1148 3203
rect 1142 3198 1148 3199
rect 1326 3203 1332 3204
rect 1326 3199 1327 3203
rect 1331 3199 1332 3203
rect 1326 3198 1332 3199
rect 1510 3203 1516 3204
rect 1510 3199 1511 3203
rect 1515 3199 1516 3203
rect 1510 3198 1516 3199
rect 1694 3203 1700 3204
rect 1694 3199 1695 3203
rect 1699 3199 1700 3203
rect 2006 3200 2007 3204
rect 2011 3200 2012 3204
rect 2006 3199 2012 3200
rect 1694 3198 1700 3199
rect 110 3187 116 3188
rect 110 3183 111 3187
rect 115 3183 116 3187
rect 2006 3187 2012 3188
rect 110 3182 116 3183
rect 134 3184 140 3185
rect 112 3151 114 3182
rect 134 3180 135 3184
rect 139 3180 140 3184
rect 134 3179 140 3180
rect 286 3184 292 3185
rect 286 3180 287 3184
rect 291 3180 292 3184
rect 286 3179 292 3180
rect 446 3184 452 3185
rect 446 3180 447 3184
rect 451 3180 452 3184
rect 446 3179 452 3180
rect 614 3184 620 3185
rect 614 3180 615 3184
rect 619 3180 620 3184
rect 614 3179 620 3180
rect 790 3184 796 3185
rect 790 3180 791 3184
rect 795 3180 796 3184
rect 790 3179 796 3180
rect 966 3184 972 3185
rect 966 3180 967 3184
rect 971 3180 972 3184
rect 966 3179 972 3180
rect 1142 3184 1148 3185
rect 1142 3180 1143 3184
rect 1147 3180 1148 3184
rect 1142 3179 1148 3180
rect 1326 3184 1332 3185
rect 1326 3180 1327 3184
rect 1331 3180 1332 3184
rect 1326 3179 1332 3180
rect 1510 3184 1516 3185
rect 1510 3180 1511 3184
rect 1515 3180 1516 3184
rect 1510 3179 1516 3180
rect 1694 3184 1700 3185
rect 1694 3180 1695 3184
rect 1699 3180 1700 3184
rect 2006 3183 2007 3187
rect 2011 3183 2012 3187
rect 2006 3182 2012 3183
rect 1694 3179 1700 3180
rect 136 3151 138 3179
rect 288 3151 290 3179
rect 448 3151 450 3179
rect 616 3151 618 3179
rect 792 3151 794 3179
rect 968 3151 970 3179
rect 1144 3151 1146 3179
rect 1328 3151 1330 3179
rect 1512 3151 1514 3179
rect 1696 3151 1698 3179
rect 2008 3151 2010 3182
rect 2048 3178 2050 3205
rect 2072 3181 2074 3205
rect 2168 3181 2170 3205
rect 2264 3181 2266 3205
rect 2360 3181 2362 3205
rect 2456 3181 2458 3205
rect 2552 3181 2554 3205
rect 2648 3181 2650 3205
rect 2744 3181 2746 3205
rect 2840 3181 2842 3205
rect 2936 3181 2938 3205
rect 3032 3181 3034 3205
rect 3128 3181 3130 3205
rect 3224 3181 3226 3205
rect 3320 3181 3322 3205
rect 3440 3181 3442 3205
rect 3576 3181 3578 3205
rect 3720 3181 3722 3205
rect 3840 3181 3842 3205
rect 2070 3180 2076 3181
rect 2046 3177 2052 3178
rect 2046 3173 2047 3177
rect 2051 3173 2052 3177
rect 2070 3176 2071 3180
rect 2075 3176 2076 3180
rect 2070 3175 2076 3176
rect 2166 3180 2172 3181
rect 2166 3176 2167 3180
rect 2171 3176 2172 3180
rect 2166 3175 2172 3176
rect 2262 3180 2268 3181
rect 2262 3176 2263 3180
rect 2267 3176 2268 3180
rect 2262 3175 2268 3176
rect 2358 3180 2364 3181
rect 2358 3176 2359 3180
rect 2363 3176 2364 3180
rect 2358 3175 2364 3176
rect 2454 3180 2460 3181
rect 2454 3176 2455 3180
rect 2459 3176 2460 3180
rect 2454 3175 2460 3176
rect 2550 3180 2556 3181
rect 2550 3176 2551 3180
rect 2555 3176 2556 3180
rect 2550 3175 2556 3176
rect 2646 3180 2652 3181
rect 2646 3176 2647 3180
rect 2651 3176 2652 3180
rect 2646 3175 2652 3176
rect 2742 3180 2748 3181
rect 2742 3176 2743 3180
rect 2747 3176 2748 3180
rect 2742 3175 2748 3176
rect 2838 3180 2844 3181
rect 2838 3176 2839 3180
rect 2843 3176 2844 3180
rect 2838 3175 2844 3176
rect 2934 3180 2940 3181
rect 2934 3176 2935 3180
rect 2939 3176 2940 3180
rect 2934 3175 2940 3176
rect 3030 3180 3036 3181
rect 3030 3176 3031 3180
rect 3035 3176 3036 3180
rect 3030 3175 3036 3176
rect 3126 3180 3132 3181
rect 3126 3176 3127 3180
rect 3131 3176 3132 3180
rect 3126 3175 3132 3176
rect 3222 3180 3228 3181
rect 3222 3176 3223 3180
rect 3227 3176 3228 3180
rect 3222 3175 3228 3176
rect 3318 3180 3324 3181
rect 3318 3176 3319 3180
rect 3323 3176 3324 3180
rect 3318 3175 3324 3176
rect 3438 3180 3444 3181
rect 3438 3176 3439 3180
rect 3443 3176 3444 3180
rect 3438 3175 3444 3176
rect 3574 3180 3580 3181
rect 3574 3176 3575 3180
rect 3579 3176 3580 3180
rect 3574 3175 3580 3176
rect 3718 3180 3724 3181
rect 3718 3176 3719 3180
rect 3723 3176 3724 3180
rect 3718 3175 3724 3176
rect 3838 3180 3844 3181
rect 3838 3176 3839 3180
rect 3843 3176 3844 3180
rect 3944 3178 3946 3205
rect 3838 3175 3844 3176
rect 3942 3177 3948 3178
rect 2046 3172 2052 3173
rect 3942 3173 3943 3177
rect 3947 3173 3948 3177
rect 3942 3172 3948 3173
rect 2070 3161 2076 3162
rect 2046 3160 2052 3161
rect 2046 3156 2047 3160
rect 2051 3156 2052 3160
rect 2070 3157 2071 3161
rect 2075 3157 2076 3161
rect 2070 3156 2076 3157
rect 2166 3161 2172 3162
rect 2166 3157 2167 3161
rect 2171 3157 2172 3161
rect 2166 3156 2172 3157
rect 2262 3161 2268 3162
rect 2262 3157 2263 3161
rect 2267 3157 2268 3161
rect 2262 3156 2268 3157
rect 2358 3161 2364 3162
rect 2358 3157 2359 3161
rect 2363 3157 2364 3161
rect 2358 3156 2364 3157
rect 2454 3161 2460 3162
rect 2454 3157 2455 3161
rect 2459 3157 2460 3161
rect 2454 3156 2460 3157
rect 2550 3161 2556 3162
rect 2550 3157 2551 3161
rect 2555 3157 2556 3161
rect 2550 3156 2556 3157
rect 2646 3161 2652 3162
rect 2646 3157 2647 3161
rect 2651 3157 2652 3161
rect 2646 3156 2652 3157
rect 2742 3161 2748 3162
rect 2742 3157 2743 3161
rect 2747 3157 2748 3161
rect 2742 3156 2748 3157
rect 2838 3161 2844 3162
rect 2838 3157 2839 3161
rect 2843 3157 2844 3161
rect 2838 3156 2844 3157
rect 2934 3161 2940 3162
rect 2934 3157 2935 3161
rect 2939 3157 2940 3161
rect 2934 3156 2940 3157
rect 3030 3161 3036 3162
rect 3030 3157 3031 3161
rect 3035 3157 3036 3161
rect 3030 3156 3036 3157
rect 3126 3161 3132 3162
rect 3126 3157 3127 3161
rect 3131 3157 3132 3161
rect 3126 3156 3132 3157
rect 3222 3161 3228 3162
rect 3222 3157 3223 3161
rect 3227 3157 3228 3161
rect 3222 3156 3228 3157
rect 3318 3161 3324 3162
rect 3318 3157 3319 3161
rect 3323 3157 3324 3161
rect 3318 3156 3324 3157
rect 3438 3161 3444 3162
rect 3438 3157 3439 3161
rect 3443 3157 3444 3161
rect 3438 3156 3444 3157
rect 3574 3161 3580 3162
rect 3574 3157 3575 3161
rect 3579 3157 3580 3161
rect 3574 3156 3580 3157
rect 3718 3161 3724 3162
rect 3718 3157 3719 3161
rect 3723 3157 3724 3161
rect 3718 3156 3724 3157
rect 3838 3161 3844 3162
rect 3838 3157 3839 3161
rect 3843 3157 3844 3161
rect 3838 3156 3844 3157
rect 3942 3160 3948 3161
rect 3942 3156 3943 3160
rect 3947 3156 3948 3160
rect 2046 3155 2052 3156
rect 111 3150 115 3151
rect 111 3145 115 3146
rect 135 3150 139 3151
rect 135 3145 139 3146
rect 287 3150 291 3151
rect 287 3145 291 3146
rect 311 3150 315 3151
rect 311 3145 315 3146
rect 439 3150 443 3151
rect 439 3145 443 3146
rect 447 3150 451 3151
rect 447 3145 451 3146
rect 583 3150 587 3151
rect 583 3145 587 3146
rect 615 3150 619 3151
rect 615 3145 619 3146
rect 743 3150 747 3151
rect 743 3145 747 3146
rect 791 3150 795 3151
rect 791 3145 795 3146
rect 903 3150 907 3151
rect 903 3145 907 3146
rect 967 3150 971 3151
rect 967 3145 971 3146
rect 1063 3150 1067 3151
rect 1063 3145 1067 3146
rect 1143 3150 1147 3151
rect 1143 3145 1147 3146
rect 1223 3150 1227 3151
rect 1223 3145 1227 3146
rect 1327 3150 1331 3151
rect 1327 3145 1331 3146
rect 1391 3150 1395 3151
rect 1391 3145 1395 3146
rect 1511 3150 1515 3151
rect 1511 3145 1515 3146
rect 1559 3150 1563 3151
rect 1559 3145 1563 3146
rect 1695 3150 1699 3151
rect 1695 3145 1699 3146
rect 1727 3150 1731 3151
rect 1727 3145 1731 3146
rect 2007 3150 2011 3151
rect 2007 3145 2011 3146
rect 112 3118 114 3145
rect 312 3121 314 3145
rect 440 3121 442 3145
rect 584 3121 586 3145
rect 744 3121 746 3145
rect 904 3121 906 3145
rect 1064 3121 1066 3145
rect 1224 3121 1226 3145
rect 1392 3121 1394 3145
rect 1560 3121 1562 3145
rect 1728 3121 1730 3145
rect 310 3120 316 3121
rect 110 3117 116 3118
rect 110 3113 111 3117
rect 115 3113 116 3117
rect 310 3116 311 3120
rect 315 3116 316 3120
rect 310 3115 316 3116
rect 438 3120 444 3121
rect 438 3116 439 3120
rect 443 3116 444 3120
rect 438 3115 444 3116
rect 582 3120 588 3121
rect 582 3116 583 3120
rect 587 3116 588 3120
rect 582 3115 588 3116
rect 742 3120 748 3121
rect 742 3116 743 3120
rect 747 3116 748 3120
rect 742 3115 748 3116
rect 902 3120 908 3121
rect 902 3116 903 3120
rect 907 3116 908 3120
rect 902 3115 908 3116
rect 1062 3120 1068 3121
rect 1062 3116 1063 3120
rect 1067 3116 1068 3120
rect 1062 3115 1068 3116
rect 1222 3120 1228 3121
rect 1222 3116 1223 3120
rect 1227 3116 1228 3120
rect 1222 3115 1228 3116
rect 1390 3120 1396 3121
rect 1390 3116 1391 3120
rect 1395 3116 1396 3120
rect 1390 3115 1396 3116
rect 1558 3120 1564 3121
rect 1558 3116 1559 3120
rect 1563 3116 1564 3120
rect 1558 3115 1564 3116
rect 1726 3120 1732 3121
rect 1726 3116 1727 3120
rect 1731 3116 1732 3120
rect 2008 3118 2010 3145
rect 2048 3123 2050 3155
rect 2072 3123 2074 3156
rect 2168 3123 2170 3156
rect 2264 3123 2266 3156
rect 2360 3123 2362 3156
rect 2456 3123 2458 3156
rect 2552 3123 2554 3156
rect 2648 3123 2650 3156
rect 2744 3123 2746 3156
rect 2840 3123 2842 3156
rect 2936 3123 2938 3156
rect 3032 3123 3034 3156
rect 3128 3123 3130 3156
rect 3224 3123 3226 3156
rect 3320 3123 3322 3156
rect 3440 3123 3442 3156
rect 3576 3123 3578 3156
rect 3720 3123 3722 3156
rect 3840 3123 3842 3156
rect 3942 3155 3948 3156
rect 3944 3123 3946 3155
rect 2047 3122 2051 3123
rect 1726 3115 1732 3116
rect 2006 3117 2012 3118
rect 2047 3117 2051 3118
rect 2071 3122 2075 3123
rect 2071 3117 2075 3118
rect 2167 3122 2171 3123
rect 2167 3117 2171 3118
rect 2263 3122 2267 3123
rect 2263 3117 2267 3118
rect 2335 3122 2339 3123
rect 2335 3117 2339 3118
rect 2359 3122 2363 3123
rect 2359 3117 2363 3118
rect 2455 3122 2459 3123
rect 2455 3117 2459 3118
rect 2551 3122 2555 3123
rect 2551 3117 2555 3118
rect 2623 3122 2627 3123
rect 2623 3117 2627 3118
rect 2647 3122 2651 3123
rect 2647 3117 2651 3118
rect 2743 3122 2747 3123
rect 2743 3117 2747 3118
rect 2839 3122 2843 3123
rect 2839 3117 2843 3118
rect 2911 3122 2915 3123
rect 2911 3117 2915 3118
rect 2935 3122 2939 3123
rect 2935 3117 2939 3118
rect 3031 3122 3035 3123
rect 3031 3117 3035 3118
rect 3127 3122 3131 3123
rect 3127 3117 3131 3118
rect 3207 3122 3211 3123
rect 3207 3117 3211 3118
rect 3223 3122 3227 3123
rect 3223 3117 3227 3118
rect 3319 3122 3323 3123
rect 3319 3117 3323 3118
rect 3439 3122 3443 3123
rect 3439 3117 3443 3118
rect 3503 3122 3507 3123
rect 3503 3117 3507 3118
rect 3575 3122 3579 3123
rect 3575 3117 3579 3118
rect 3719 3122 3723 3123
rect 3719 3117 3723 3118
rect 3799 3122 3803 3123
rect 3799 3117 3803 3118
rect 3839 3122 3843 3123
rect 3839 3117 3843 3118
rect 3943 3122 3947 3123
rect 3943 3117 3947 3118
rect 110 3112 116 3113
rect 2006 3113 2007 3117
rect 2011 3113 2012 3117
rect 2006 3112 2012 3113
rect 310 3101 316 3102
rect 110 3100 116 3101
rect 110 3096 111 3100
rect 115 3096 116 3100
rect 310 3097 311 3101
rect 315 3097 316 3101
rect 310 3096 316 3097
rect 438 3101 444 3102
rect 438 3097 439 3101
rect 443 3097 444 3101
rect 438 3096 444 3097
rect 582 3101 588 3102
rect 582 3097 583 3101
rect 587 3097 588 3101
rect 582 3096 588 3097
rect 742 3101 748 3102
rect 742 3097 743 3101
rect 747 3097 748 3101
rect 742 3096 748 3097
rect 902 3101 908 3102
rect 902 3097 903 3101
rect 907 3097 908 3101
rect 902 3096 908 3097
rect 1062 3101 1068 3102
rect 1062 3097 1063 3101
rect 1067 3097 1068 3101
rect 1062 3096 1068 3097
rect 1222 3101 1228 3102
rect 1222 3097 1223 3101
rect 1227 3097 1228 3101
rect 1222 3096 1228 3097
rect 1390 3101 1396 3102
rect 1390 3097 1391 3101
rect 1395 3097 1396 3101
rect 1390 3096 1396 3097
rect 1558 3101 1564 3102
rect 1558 3097 1559 3101
rect 1563 3097 1564 3101
rect 1558 3096 1564 3097
rect 1726 3101 1732 3102
rect 1726 3097 1727 3101
rect 1731 3097 1732 3101
rect 1726 3096 1732 3097
rect 2006 3100 2012 3101
rect 2006 3096 2007 3100
rect 2011 3096 2012 3100
rect 2048 3097 2050 3117
rect 110 3095 116 3096
rect 112 3067 114 3095
rect 312 3067 314 3096
rect 440 3067 442 3096
rect 584 3067 586 3096
rect 744 3067 746 3096
rect 904 3067 906 3096
rect 1064 3067 1066 3096
rect 1224 3067 1226 3096
rect 1392 3067 1394 3096
rect 1560 3067 1562 3096
rect 1728 3067 1730 3096
rect 2006 3095 2012 3096
rect 2046 3096 2052 3097
rect 2072 3096 2074 3117
rect 2336 3096 2338 3117
rect 2624 3096 2626 3117
rect 2912 3096 2914 3117
rect 3208 3096 3210 3117
rect 3504 3096 3506 3117
rect 3800 3096 3802 3117
rect 3944 3097 3946 3117
rect 3942 3096 3948 3097
rect 2008 3067 2010 3095
rect 2046 3092 2047 3096
rect 2051 3092 2052 3096
rect 2046 3091 2052 3092
rect 2070 3095 2076 3096
rect 2070 3091 2071 3095
rect 2075 3091 2076 3095
rect 2070 3090 2076 3091
rect 2334 3095 2340 3096
rect 2334 3091 2335 3095
rect 2339 3091 2340 3095
rect 2334 3090 2340 3091
rect 2622 3095 2628 3096
rect 2622 3091 2623 3095
rect 2627 3091 2628 3095
rect 2622 3090 2628 3091
rect 2910 3095 2916 3096
rect 2910 3091 2911 3095
rect 2915 3091 2916 3095
rect 2910 3090 2916 3091
rect 3206 3095 3212 3096
rect 3206 3091 3207 3095
rect 3211 3091 3212 3095
rect 3206 3090 3212 3091
rect 3502 3095 3508 3096
rect 3502 3091 3503 3095
rect 3507 3091 3508 3095
rect 3502 3090 3508 3091
rect 3798 3095 3804 3096
rect 3798 3091 3799 3095
rect 3803 3091 3804 3095
rect 3942 3092 3943 3096
rect 3947 3092 3948 3096
rect 3942 3091 3948 3092
rect 3798 3090 3804 3091
rect 2046 3079 2052 3080
rect 2046 3075 2047 3079
rect 2051 3075 2052 3079
rect 3942 3079 3948 3080
rect 2046 3074 2052 3075
rect 2070 3076 2076 3077
rect 111 3066 115 3067
rect 111 3061 115 3062
rect 311 3066 315 3067
rect 311 3061 315 3062
rect 439 3066 443 3067
rect 439 3061 443 3062
rect 503 3066 507 3067
rect 503 3061 507 3062
rect 583 3066 587 3067
rect 583 3061 587 3062
rect 599 3066 603 3067
rect 599 3061 603 3062
rect 703 3066 707 3067
rect 703 3061 707 3062
rect 743 3066 747 3067
rect 743 3061 747 3062
rect 815 3066 819 3067
rect 815 3061 819 3062
rect 903 3066 907 3067
rect 903 3061 907 3062
rect 935 3066 939 3067
rect 935 3061 939 3062
rect 1063 3066 1067 3067
rect 1063 3061 1067 3062
rect 1071 3066 1075 3067
rect 1071 3061 1075 3062
rect 1223 3066 1227 3067
rect 1223 3061 1227 3062
rect 1383 3066 1387 3067
rect 1383 3061 1387 3062
rect 1391 3066 1395 3067
rect 1391 3061 1395 3062
rect 1551 3066 1555 3067
rect 1551 3061 1555 3062
rect 1559 3066 1563 3067
rect 1559 3061 1563 3062
rect 1719 3066 1723 3067
rect 1719 3061 1723 3062
rect 1727 3066 1731 3067
rect 1727 3061 1731 3062
rect 2007 3066 2011 3067
rect 2007 3061 2011 3062
rect 112 3041 114 3061
rect 110 3040 116 3041
rect 504 3040 506 3061
rect 600 3040 602 3061
rect 704 3040 706 3061
rect 816 3040 818 3061
rect 936 3040 938 3061
rect 1072 3040 1074 3061
rect 1224 3040 1226 3061
rect 1384 3040 1386 3061
rect 1552 3040 1554 3061
rect 1720 3040 1722 3061
rect 2008 3041 2010 3061
rect 2048 3047 2050 3074
rect 2070 3072 2071 3076
rect 2075 3072 2076 3076
rect 2070 3071 2076 3072
rect 2334 3076 2340 3077
rect 2334 3072 2335 3076
rect 2339 3072 2340 3076
rect 2334 3071 2340 3072
rect 2622 3076 2628 3077
rect 2622 3072 2623 3076
rect 2627 3072 2628 3076
rect 2622 3071 2628 3072
rect 2910 3076 2916 3077
rect 2910 3072 2911 3076
rect 2915 3072 2916 3076
rect 2910 3071 2916 3072
rect 3206 3076 3212 3077
rect 3206 3072 3207 3076
rect 3211 3072 3212 3076
rect 3206 3071 3212 3072
rect 3502 3076 3508 3077
rect 3502 3072 3503 3076
rect 3507 3072 3508 3076
rect 3502 3071 3508 3072
rect 3798 3076 3804 3077
rect 3798 3072 3799 3076
rect 3803 3072 3804 3076
rect 3942 3075 3943 3079
rect 3947 3075 3948 3079
rect 3942 3074 3948 3075
rect 3798 3071 3804 3072
rect 2072 3047 2074 3071
rect 2336 3047 2338 3071
rect 2624 3047 2626 3071
rect 2912 3047 2914 3071
rect 3208 3047 3210 3071
rect 3504 3047 3506 3071
rect 3800 3047 3802 3071
rect 3944 3047 3946 3074
rect 2047 3046 2051 3047
rect 2047 3041 2051 3042
rect 2071 3046 2075 3047
rect 2071 3041 2075 3042
rect 2335 3046 2339 3047
rect 2335 3041 2339 3042
rect 2383 3046 2387 3047
rect 2383 3041 2387 3042
rect 2623 3046 2627 3047
rect 2623 3041 2627 3042
rect 2703 3046 2707 3047
rect 2703 3041 2707 3042
rect 2911 3046 2915 3047
rect 2911 3041 2915 3042
rect 2999 3046 3003 3047
rect 2999 3041 3003 3042
rect 3207 3046 3211 3047
rect 3207 3041 3211 3042
rect 3287 3046 3291 3047
rect 3287 3041 3291 3042
rect 3503 3046 3507 3047
rect 3503 3041 3507 3042
rect 3575 3046 3579 3047
rect 3575 3041 3579 3042
rect 3799 3046 3803 3047
rect 3799 3041 3803 3042
rect 3839 3046 3843 3047
rect 3839 3041 3843 3042
rect 3943 3046 3947 3047
rect 3943 3041 3947 3042
rect 2006 3040 2012 3041
rect 110 3036 111 3040
rect 115 3036 116 3040
rect 110 3035 116 3036
rect 502 3039 508 3040
rect 502 3035 503 3039
rect 507 3035 508 3039
rect 502 3034 508 3035
rect 598 3039 604 3040
rect 598 3035 599 3039
rect 603 3035 604 3039
rect 598 3034 604 3035
rect 702 3039 708 3040
rect 702 3035 703 3039
rect 707 3035 708 3039
rect 702 3034 708 3035
rect 814 3039 820 3040
rect 814 3035 815 3039
rect 819 3035 820 3039
rect 814 3034 820 3035
rect 934 3039 940 3040
rect 934 3035 935 3039
rect 939 3035 940 3039
rect 934 3034 940 3035
rect 1070 3039 1076 3040
rect 1070 3035 1071 3039
rect 1075 3035 1076 3039
rect 1070 3034 1076 3035
rect 1222 3039 1228 3040
rect 1222 3035 1223 3039
rect 1227 3035 1228 3039
rect 1222 3034 1228 3035
rect 1382 3039 1388 3040
rect 1382 3035 1383 3039
rect 1387 3035 1388 3039
rect 1382 3034 1388 3035
rect 1550 3039 1556 3040
rect 1550 3035 1551 3039
rect 1555 3035 1556 3039
rect 1550 3034 1556 3035
rect 1718 3039 1724 3040
rect 1718 3035 1719 3039
rect 1723 3035 1724 3039
rect 2006 3036 2007 3040
rect 2011 3036 2012 3040
rect 2006 3035 2012 3036
rect 1718 3034 1724 3035
rect 110 3023 116 3024
rect 110 3019 111 3023
rect 115 3019 116 3023
rect 2006 3023 2012 3024
rect 110 3018 116 3019
rect 502 3020 508 3021
rect 112 2987 114 3018
rect 502 3016 503 3020
rect 507 3016 508 3020
rect 502 3015 508 3016
rect 598 3020 604 3021
rect 598 3016 599 3020
rect 603 3016 604 3020
rect 598 3015 604 3016
rect 702 3020 708 3021
rect 702 3016 703 3020
rect 707 3016 708 3020
rect 702 3015 708 3016
rect 814 3020 820 3021
rect 814 3016 815 3020
rect 819 3016 820 3020
rect 814 3015 820 3016
rect 934 3020 940 3021
rect 934 3016 935 3020
rect 939 3016 940 3020
rect 934 3015 940 3016
rect 1070 3020 1076 3021
rect 1070 3016 1071 3020
rect 1075 3016 1076 3020
rect 1070 3015 1076 3016
rect 1222 3020 1228 3021
rect 1222 3016 1223 3020
rect 1227 3016 1228 3020
rect 1222 3015 1228 3016
rect 1382 3020 1388 3021
rect 1382 3016 1383 3020
rect 1387 3016 1388 3020
rect 1382 3015 1388 3016
rect 1550 3020 1556 3021
rect 1550 3016 1551 3020
rect 1555 3016 1556 3020
rect 1550 3015 1556 3016
rect 1718 3020 1724 3021
rect 1718 3016 1719 3020
rect 1723 3016 1724 3020
rect 2006 3019 2007 3023
rect 2011 3019 2012 3023
rect 2006 3018 2012 3019
rect 1718 3015 1724 3016
rect 504 2987 506 3015
rect 600 2987 602 3015
rect 704 2987 706 3015
rect 816 2987 818 3015
rect 936 2987 938 3015
rect 1072 2987 1074 3015
rect 1224 2987 1226 3015
rect 1384 2987 1386 3015
rect 1552 2987 1554 3015
rect 1720 2987 1722 3015
rect 2008 2987 2010 3018
rect 2048 3014 2050 3041
rect 2072 3017 2074 3041
rect 2384 3017 2386 3041
rect 2704 3017 2706 3041
rect 3000 3017 3002 3041
rect 3288 3017 3290 3041
rect 3576 3017 3578 3041
rect 3840 3017 3842 3041
rect 2070 3016 2076 3017
rect 2046 3013 2052 3014
rect 2046 3009 2047 3013
rect 2051 3009 2052 3013
rect 2070 3012 2071 3016
rect 2075 3012 2076 3016
rect 2070 3011 2076 3012
rect 2382 3016 2388 3017
rect 2382 3012 2383 3016
rect 2387 3012 2388 3016
rect 2382 3011 2388 3012
rect 2702 3016 2708 3017
rect 2702 3012 2703 3016
rect 2707 3012 2708 3016
rect 2702 3011 2708 3012
rect 2998 3016 3004 3017
rect 2998 3012 2999 3016
rect 3003 3012 3004 3016
rect 2998 3011 3004 3012
rect 3286 3016 3292 3017
rect 3286 3012 3287 3016
rect 3291 3012 3292 3016
rect 3286 3011 3292 3012
rect 3574 3016 3580 3017
rect 3574 3012 3575 3016
rect 3579 3012 3580 3016
rect 3574 3011 3580 3012
rect 3838 3016 3844 3017
rect 3838 3012 3839 3016
rect 3843 3012 3844 3016
rect 3944 3014 3946 3041
rect 3838 3011 3844 3012
rect 3942 3013 3948 3014
rect 2046 3008 2052 3009
rect 3942 3009 3943 3013
rect 3947 3009 3948 3013
rect 3942 3008 3948 3009
rect 2070 2997 2076 2998
rect 2046 2996 2052 2997
rect 2046 2992 2047 2996
rect 2051 2992 2052 2996
rect 2070 2993 2071 2997
rect 2075 2993 2076 2997
rect 2070 2992 2076 2993
rect 2382 2997 2388 2998
rect 2382 2993 2383 2997
rect 2387 2993 2388 2997
rect 2382 2992 2388 2993
rect 2702 2997 2708 2998
rect 2702 2993 2703 2997
rect 2707 2993 2708 2997
rect 2702 2992 2708 2993
rect 2998 2997 3004 2998
rect 2998 2993 2999 2997
rect 3003 2993 3004 2997
rect 2998 2992 3004 2993
rect 3286 2997 3292 2998
rect 3286 2993 3287 2997
rect 3291 2993 3292 2997
rect 3286 2992 3292 2993
rect 3574 2997 3580 2998
rect 3574 2993 3575 2997
rect 3579 2993 3580 2997
rect 3574 2992 3580 2993
rect 3838 2997 3844 2998
rect 3838 2993 3839 2997
rect 3843 2993 3844 2997
rect 3838 2992 3844 2993
rect 3942 2996 3948 2997
rect 3942 2992 3943 2996
rect 3947 2992 3948 2996
rect 2046 2991 2052 2992
rect 111 2986 115 2987
rect 111 2981 115 2982
rect 503 2986 507 2987
rect 503 2981 507 2982
rect 551 2986 555 2987
rect 551 2981 555 2982
rect 599 2986 603 2987
rect 599 2981 603 2982
rect 647 2986 651 2987
rect 647 2981 651 2982
rect 703 2986 707 2987
rect 703 2981 707 2982
rect 759 2986 763 2987
rect 759 2981 763 2982
rect 815 2986 819 2987
rect 815 2981 819 2982
rect 887 2986 891 2987
rect 887 2981 891 2982
rect 935 2986 939 2987
rect 935 2981 939 2982
rect 1023 2986 1027 2987
rect 1023 2981 1027 2982
rect 1071 2986 1075 2987
rect 1071 2981 1075 2982
rect 1175 2986 1179 2987
rect 1175 2981 1179 2982
rect 1223 2986 1227 2987
rect 1223 2981 1227 2982
rect 1327 2986 1331 2987
rect 1327 2981 1331 2982
rect 1383 2986 1387 2987
rect 1383 2981 1387 2982
rect 1487 2986 1491 2987
rect 1487 2981 1491 2982
rect 1551 2986 1555 2987
rect 1551 2981 1555 2982
rect 1655 2986 1659 2987
rect 1655 2981 1659 2982
rect 1719 2986 1723 2987
rect 1719 2981 1723 2982
rect 1823 2986 1827 2987
rect 1823 2981 1827 2982
rect 2007 2986 2011 2987
rect 2007 2981 2011 2982
rect 112 2954 114 2981
rect 552 2957 554 2981
rect 648 2957 650 2981
rect 760 2957 762 2981
rect 888 2957 890 2981
rect 1024 2957 1026 2981
rect 1176 2957 1178 2981
rect 1328 2957 1330 2981
rect 1488 2957 1490 2981
rect 1656 2957 1658 2981
rect 1824 2957 1826 2981
rect 550 2956 556 2957
rect 110 2953 116 2954
rect 110 2949 111 2953
rect 115 2949 116 2953
rect 550 2952 551 2956
rect 555 2952 556 2956
rect 550 2951 556 2952
rect 646 2956 652 2957
rect 646 2952 647 2956
rect 651 2952 652 2956
rect 646 2951 652 2952
rect 758 2956 764 2957
rect 758 2952 759 2956
rect 763 2952 764 2956
rect 758 2951 764 2952
rect 886 2956 892 2957
rect 886 2952 887 2956
rect 891 2952 892 2956
rect 886 2951 892 2952
rect 1022 2956 1028 2957
rect 1022 2952 1023 2956
rect 1027 2952 1028 2956
rect 1022 2951 1028 2952
rect 1174 2956 1180 2957
rect 1174 2952 1175 2956
rect 1179 2952 1180 2956
rect 1174 2951 1180 2952
rect 1326 2956 1332 2957
rect 1326 2952 1327 2956
rect 1331 2952 1332 2956
rect 1326 2951 1332 2952
rect 1486 2956 1492 2957
rect 1486 2952 1487 2956
rect 1491 2952 1492 2956
rect 1486 2951 1492 2952
rect 1654 2956 1660 2957
rect 1654 2952 1655 2956
rect 1659 2952 1660 2956
rect 1654 2951 1660 2952
rect 1822 2956 1828 2957
rect 1822 2952 1823 2956
rect 1827 2952 1828 2956
rect 2008 2954 2010 2981
rect 2048 2967 2050 2991
rect 2072 2967 2074 2992
rect 2384 2967 2386 2992
rect 2704 2967 2706 2992
rect 3000 2967 3002 2992
rect 3288 2967 3290 2992
rect 3576 2967 3578 2992
rect 3840 2967 3842 2992
rect 3942 2991 3948 2992
rect 3944 2967 3946 2991
rect 2047 2966 2051 2967
rect 2047 2961 2051 2962
rect 2071 2966 2075 2967
rect 2071 2961 2075 2962
rect 2383 2966 2387 2967
rect 2383 2961 2387 2962
rect 2391 2966 2395 2967
rect 2391 2961 2395 2962
rect 2703 2966 2707 2967
rect 2703 2961 2707 2962
rect 2975 2966 2979 2967
rect 2975 2961 2979 2962
rect 2999 2966 3003 2967
rect 2999 2961 3003 2962
rect 3215 2966 3219 2967
rect 3215 2961 3219 2962
rect 3287 2966 3291 2967
rect 3287 2961 3291 2962
rect 3439 2966 3443 2967
rect 3439 2961 3443 2962
rect 3575 2966 3579 2967
rect 3575 2961 3579 2962
rect 3647 2966 3651 2967
rect 3647 2961 3651 2962
rect 3839 2966 3843 2967
rect 3839 2961 3843 2962
rect 3943 2966 3947 2967
rect 3943 2961 3947 2962
rect 1822 2951 1828 2952
rect 2006 2953 2012 2954
rect 110 2948 116 2949
rect 2006 2949 2007 2953
rect 2011 2949 2012 2953
rect 2006 2948 2012 2949
rect 2048 2941 2050 2961
rect 2046 2940 2052 2941
rect 2072 2940 2074 2961
rect 2392 2940 2394 2961
rect 2704 2940 2706 2961
rect 2976 2940 2978 2961
rect 3216 2940 3218 2961
rect 3440 2940 3442 2961
rect 3648 2940 3650 2961
rect 3840 2940 3842 2961
rect 3944 2941 3946 2961
rect 3942 2940 3948 2941
rect 550 2937 556 2938
rect 110 2936 116 2937
rect 110 2932 111 2936
rect 115 2932 116 2936
rect 550 2933 551 2937
rect 555 2933 556 2937
rect 550 2932 556 2933
rect 646 2937 652 2938
rect 646 2933 647 2937
rect 651 2933 652 2937
rect 646 2932 652 2933
rect 758 2937 764 2938
rect 758 2933 759 2937
rect 763 2933 764 2937
rect 758 2932 764 2933
rect 886 2937 892 2938
rect 886 2933 887 2937
rect 891 2933 892 2937
rect 886 2932 892 2933
rect 1022 2937 1028 2938
rect 1022 2933 1023 2937
rect 1027 2933 1028 2937
rect 1022 2932 1028 2933
rect 1174 2937 1180 2938
rect 1174 2933 1175 2937
rect 1179 2933 1180 2937
rect 1174 2932 1180 2933
rect 1326 2937 1332 2938
rect 1326 2933 1327 2937
rect 1331 2933 1332 2937
rect 1326 2932 1332 2933
rect 1486 2937 1492 2938
rect 1486 2933 1487 2937
rect 1491 2933 1492 2937
rect 1486 2932 1492 2933
rect 1654 2937 1660 2938
rect 1654 2933 1655 2937
rect 1659 2933 1660 2937
rect 1654 2932 1660 2933
rect 1822 2937 1828 2938
rect 1822 2933 1823 2937
rect 1827 2933 1828 2937
rect 1822 2932 1828 2933
rect 2006 2936 2012 2937
rect 2006 2932 2007 2936
rect 2011 2932 2012 2936
rect 2046 2936 2047 2940
rect 2051 2936 2052 2940
rect 2046 2935 2052 2936
rect 2070 2939 2076 2940
rect 2070 2935 2071 2939
rect 2075 2935 2076 2939
rect 2070 2934 2076 2935
rect 2390 2939 2396 2940
rect 2390 2935 2391 2939
rect 2395 2935 2396 2939
rect 2390 2934 2396 2935
rect 2702 2939 2708 2940
rect 2702 2935 2703 2939
rect 2707 2935 2708 2939
rect 2702 2934 2708 2935
rect 2974 2939 2980 2940
rect 2974 2935 2975 2939
rect 2979 2935 2980 2939
rect 2974 2934 2980 2935
rect 3214 2939 3220 2940
rect 3214 2935 3215 2939
rect 3219 2935 3220 2939
rect 3214 2934 3220 2935
rect 3438 2939 3444 2940
rect 3438 2935 3439 2939
rect 3443 2935 3444 2939
rect 3438 2934 3444 2935
rect 3646 2939 3652 2940
rect 3646 2935 3647 2939
rect 3651 2935 3652 2939
rect 3646 2934 3652 2935
rect 3838 2939 3844 2940
rect 3838 2935 3839 2939
rect 3843 2935 3844 2939
rect 3942 2936 3943 2940
rect 3947 2936 3948 2940
rect 3942 2935 3948 2936
rect 3838 2934 3844 2935
rect 110 2931 116 2932
rect 112 2903 114 2931
rect 552 2903 554 2932
rect 648 2903 650 2932
rect 760 2903 762 2932
rect 888 2903 890 2932
rect 1024 2903 1026 2932
rect 1176 2903 1178 2932
rect 1328 2903 1330 2932
rect 1488 2903 1490 2932
rect 1656 2903 1658 2932
rect 1824 2903 1826 2932
rect 2006 2931 2012 2932
rect 2008 2903 2010 2931
rect 2046 2923 2052 2924
rect 2046 2919 2047 2923
rect 2051 2919 2052 2923
rect 3942 2923 3948 2924
rect 2046 2918 2052 2919
rect 2070 2920 2076 2921
rect 111 2902 115 2903
rect 111 2897 115 2898
rect 471 2902 475 2903
rect 471 2897 475 2898
rect 551 2902 555 2903
rect 551 2897 555 2898
rect 575 2902 579 2903
rect 575 2897 579 2898
rect 647 2902 651 2903
rect 647 2897 651 2898
rect 695 2902 699 2903
rect 695 2897 699 2898
rect 759 2902 763 2903
rect 759 2897 763 2898
rect 839 2902 843 2903
rect 839 2897 843 2898
rect 887 2902 891 2903
rect 887 2897 891 2898
rect 991 2902 995 2903
rect 991 2897 995 2898
rect 1023 2902 1027 2903
rect 1023 2897 1027 2898
rect 1151 2902 1155 2903
rect 1151 2897 1155 2898
rect 1175 2902 1179 2903
rect 1175 2897 1179 2898
rect 1319 2902 1323 2903
rect 1319 2897 1323 2898
rect 1327 2902 1331 2903
rect 1327 2897 1331 2898
rect 1487 2902 1491 2903
rect 1487 2897 1491 2898
rect 1495 2902 1499 2903
rect 1495 2897 1499 2898
rect 1655 2902 1659 2903
rect 1655 2897 1659 2898
rect 1671 2902 1675 2903
rect 1671 2897 1675 2898
rect 1823 2902 1827 2903
rect 1823 2897 1827 2898
rect 1847 2902 1851 2903
rect 1847 2897 1851 2898
rect 2007 2902 2011 2903
rect 2007 2897 2011 2898
rect 112 2877 114 2897
rect 110 2876 116 2877
rect 472 2876 474 2897
rect 576 2876 578 2897
rect 696 2876 698 2897
rect 840 2876 842 2897
rect 992 2876 994 2897
rect 1152 2876 1154 2897
rect 1320 2876 1322 2897
rect 1496 2876 1498 2897
rect 1672 2876 1674 2897
rect 1848 2876 1850 2897
rect 2008 2877 2010 2897
rect 2048 2891 2050 2918
rect 2070 2916 2071 2920
rect 2075 2916 2076 2920
rect 2070 2915 2076 2916
rect 2390 2920 2396 2921
rect 2390 2916 2391 2920
rect 2395 2916 2396 2920
rect 2390 2915 2396 2916
rect 2702 2920 2708 2921
rect 2702 2916 2703 2920
rect 2707 2916 2708 2920
rect 2702 2915 2708 2916
rect 2974 2920 2980 2921
rect 2974 2916 2975 2920
rect 2979 2916 2980 2920
rect 2974 2915 2980 2916
rect 3214 2920 3220 2921
rect 3214 2916 3215 2920
rect 3219 2916 3220 2920
rect 3214 2915 3220 2916
rect 3438 2920 3444 2921
rect 3438 2916 3439 2920
rect 3443 2916 3444 2920
rect 3438 2915 3444 2916
rect 3646 2920 3652 2921
rect 3646 2916 3647 2920
rect 3651 2916 3652 2920
rect 3646 2915 3652 2916
rect 3838 2920 3844 2921
rect 3838 2916 3839 2920
rect 3843 2916 3844 2920
rect 3942 2919 3943 2923
rect 3947 2919 3948 2923
rect 3942 2918 3948 2919
rect 3838 2915 3844 2916
rect 2072 2891 2074 2915
rect 2392 2891 2394 2915
rect 2704 2891 2706 2915
rect 2976 2891 2978 2915
rect 3216 2891 3218 2915
rect 3440 2891 3442 2915
rect 3648 2891 3650 2915
rect 3840 2891 3842 2915
rect 3944 2891 3946 2918
rect 2047 2890 2051 2891
rect 2047 2885 2051 2886
rect 2071 2890 2075 2891
rect 2071 2885 2075 2886
rect 2295 2890 2299 2891
rect 2295 2885 2299 2886
rect 2391 2890 2395 2891
rect 2391 2885 2395 2886
rect 2535 2890 2539 2891
rect 2535 2885 2539 2886
rect 2703 2890 2707 2891
rect 2703 2885 2707 2886
rect 2767 2890 2771 2891
rect 2767 2885 2771 2886
rect 2975 2890 2979 2891
rect 2975 2885 2979 2886
rect 2991 2890 2995 2891
rect 2991 2885 2995 2886
rect 3215 2890 3219 2891
rect 3215 2885 3219 2886
rect 3431 2890 3435 2891
rect 3431 2885 3435 2886
rect 3439 2890 3443 2891
rect 3439 2885 3443 2886
rect 3647 2890 3651 2891
rect 3647 2885 3651 2886
rect 3839 2890 3843 2891
rect 3839 2885 3843 2886
rect 3943 2890 3947 2891
rect 3943 2885 3947 2886
rect 2006 2876 2012 2877
rect 110 2872 111 2876
rect 115 2872 116 2876
rect 110 2871 116 2872
rect 470 2875 476 2876
rect 470 2871 471 2875
rect 475 2871 476 2875
rect 470 2870 476 2871
rect 574 2875 580 2876
rect 574 2871 575 2875
rect 579 2871 580 2875
rect 574 2870 580 2871
rect 694 2875 700 2876
rect 694 2871 695 2875
rect 699 2871 700 2875
rect 694 2870 700 2871
rect 838 2875 844 2876
rect 838 2871 839 2875
rect 843 2871 844 2875
rect 838 2870 844 2871
rect 990 2875 996 2876
rect 990 2871 991 2875
rect 995 2871 996 2875
rect 990 2870 996 2871
rect 1150 2875 1156 2876
rect 1150 2871 1151 2875
rect 1155 2871 1156 2875
rect 1150 2870 1156 2871
rect 1318 2875 1324 2876
rect 1318 2871 1319 2875
rect 1323 2871 1324 2875
rect 1318 2870 1324 2871
rect 1494 2875 1500 2876
rect 1494 2871 1495 2875
rect 1499 2871 1500 2875
rect 1494 2870 1500 2871
rect 1670 2875 1676 2876
rect 1670 2871 1671 2875
rect 1675 2871 1676 2875
rect 1670 2870 1676 2871
rect 1846 2875 1852 2876
rect 1846 2871 1847 2875
rect 1851 2871 1852 2875
rect 2006 2872 2007 2876
rect 2011 2872 2012 2876
rect 2006 2871 2012 2872
rect 1846 2870 1852 2871
rect 110 2859 116 2860
rect 110 2855 111 2859
rect 115 2855 116 2859
rect 2006 2859 2012 2860
rect 110 2854 116 2855
rect 470 2856 476 2857
rect 112 2823 114 2854
rect 470 2852 471 2856
rect 475 2852 476 2856
rect 470 2851 476 2852
rect 574 2856 580 2857
rect 574 2852 575 2856
rect 579 2852 580 2856
rect 574 2851 580 2852
rect 694 2856 700 2857
rect 694 2852 695 2856
rect 699 2852 700 2856
rect 694 2851 700 2852
rect 838 2856 844 2857
rect 838 2852 839 2856
rect 843 2852 844 2856
rect 838 2851 844 2852
rect 990 2856 996 2857
rect 990 2852 991 2856
rect 995 2852 996 2856
rect 990 2851 996 2852
rect 1150 2856 1156 2857
rect 1150 2852 1151 2856
rect 1155 2852 1156 2856
rect 1150 2851 1156 2852
rect 1318 2856 1324 2857
rect 1318 2852 1319 2856
rect 1323 2852 1324 2856
rect 1318 2851 1324 2852
rect 1494 2856 1500 2857
rect 1494 2852 1495 2856
rect 1499 2852 1500 2856
rect 1494 2851 1500 2852
rect 1670 2856 1676 2857
rect 1670 2852 1671 2856
rect 1675 2852 1676 2856
rect 1670 2851 1676 2852
rect 1846 2856 1852 2857
rect 1846 2852 1847 2856
rect 1851 2852 1852 2856
rect 2006 2855 2007 2859
rect 2011 2855 2012 2859
rect 2048 2858 2050 2885
rect 2072 2861 2074 2885
rect 2296 2861 2298 2885
rect 2536 2861 2538 2885
rect 2768 2861 2770 2885
rect 2992 2861 2994 2885
rect 3216 2861 3218 2885
rect 3432 2861 3434 2885
rect 3648 2861 3650 2885
rect 3840 2861 3842 2885
rect 2070 2860 2076 2861
rect 2006 2854 2012 2855
rect 2046 2857 2052 2858
rect 1846 2851 1852 2852
rect 472 2823 474 2851
rect 576 2823 578 2851
rect 696 2823 698 2851
rect 840 2823 842 2851
rect 992 2823 994 2851
rect 1152 2823 1154 2851
rect 1320 2823 1322 2851
rect 1496 2823 1498 2851
rect 1672 2823 1674 2851
rect 1848 2823 1850 2851
rect 2008 2823 2010 2854
rect 2046 2853 2047 2857
rect 2051 2853 2052 2857
rect 2070 2856 2071 2860
rect 2075 2856 2076 2860
rect 2070 2855 2076 2856
rect 2294 2860 2300 2861
rect 2294 2856 2295 2860
rect 2299 2856 2300 2860
rect 2294 2855 2300 2856
rect 2534 2860 2540 2861
rect 2534 2856 2535 2860
rect 2539 2856 2540 2860
rect 2534 2855 2540 2856
rect 2766 2860 2772 2861
rect 2766 2856 2767 2860
rect 2771 2856 2772 2860
rect 2766 2855 2772 2856
rect 2990 2860 2996 2861
rect 2990 2856 2991 2860
rect 2995 2856 2996 2860
rect 2990 2855 2996 2856
rect 3214 2860 3220 2861
rect 3214 2856 3215 2860
rect 3219 2856 3220 2860
rect 3214 2855 3220 2856
rect 3430 2860 3436 2861
rect 3430 2856 3431 2860
rect 3435 2856 3436 2860
rect 3430 2855 3436 2856
rect 3646 2860 3652 2861
rect 3646 2856 3647 2860
rect 3651 2856 3652 2860
rect 3646 2855 3652 2856
rect 3838 2860 3844 2861
rect 3838 2856 3839 2860
rect 3843 2856 3844 2860
rect 3944 2858 3946 2885
rect 3838 2855 3844 2856
rect 3942 2857 3948 2858
rect 2046 2852 2052 2853
rect 3942 2853 3943 2857
rect 3947 2853 3948 2857
rect 3942 2852 3948 2853
rect 2070 2841 2076 2842
rect 2046 2840 2052 2841
rect 2046 2836 2047 2840
rect 2051 2836 2052 2840
rect 2070 2837 2071 2841
rect 2075 2837 2076 2841
rect 2070 2836 2076 2837
rect 2294 2841 2300 2842
rect 2294 2837 2295 2841
rect 2299 2837 2300 2841
rect 2294 2836 2300 2837
rect 2534 2841 2540 2842
rect 2534 2837 2535 2841
rect 2539 2837 2540 2841
rect 2534 2836 2540 2837
rect 2766 2841 2772 2842
rect 2766 2837 2767 2841
rect 2771 2837 2772 2841
rect 2766 2836 2772 2837
rect 2990 2841 2996 2842
rect 2990 2837 2991 2841
rect 2995 2837 2996 2841
rect 2990 2836 2996 2837
rect 3214 2841 3220 2842
rect 3214 2837 3215 2841
rect 3219 2837 3220 2841
rect 3214 2836 3220 2837
rect 3430 2841 3436 2842
rect 3430 2837 3431 2841
rect 3435 2837 3436 2841
rect 3430 2836 3436 2837
rect 3646 2841 3652 2842
rect 3646 2837 3647 2841
rect 3651 2837 3652 2841
rect 3646 2836 3652 2837
rect 3838 2841 3844 2842
rect 3838 2837 3839 2841
rect 3843 2837 3844 2841
rect 3838 2836 3844 2837
rect 3942 2840 3948 2841
rect 3942 2836 3943 2840
rect 3947 2836 3948 2840
rect 2046 2835 2052 2836
rect 111 2822 115 2823
rect 111 2817 115 2818
rect 471 2822 475 2823
rect 471 2817 475 2818
rect 479 2822 483 2823
rect 479 2817 483 2818
rect 575 2822 579 2823
rect 575 2817 579 2818
rect 679 2822 683 2823
rect 679 2817 683 2818
rect 695 2822 699 2823
rect 695 2817 699 2818
rect 799 2822 803 2823
rect 799 2817 803 2818
rect 839 2822 843 2823
rect 839 2817 843 2818
rect 935 2822 939 2823
rect 935 2817 939 2818
rect 991 2822 995 2823
rect 991 2817 995 2818
rect 1079 2822 1083 2823
rect 1079 2817 1083 2818
rect 1151 2822 1155 2823
rect 1151 2817 1155 2818
rect 1239 2822 1243 2823
rect 1239 2817 1243 2818
rect 1319 2822 1323 2823
rect 1319 2817 1323 2818
rect 1415 2822 1419 2823
rect 1415 2817 1419 2818
rect 1495 2822 1499 2823
rect 1495 2817 1499 2818
rect 1599 2822 1603 2823
rect 1599 2817 1603 2818
rect 1671 2822 1675 2823
rect 1671 2817 1675 2818
rect 1783 2822 1787 2823
rect 1783 2817 1787 2818
rect 1847 2822 1851 2823
rect 1847 2817 1851 2818
rect 2007 2822 2011 2823
rect 2007 2817 2011 2818
rect 112 2790 114 2817
rect 480 2793 482 2817
rect 576 2793 578 2817
rect 680 2793 682 2817
rect 800 2793 802 2817
rect 936 2793 938 2817
rect 1080 2793 1082 2817
rect 1240 2793 1242 2817
rect 1416 2793 1418 2817
rect 1600 2793 1602 2817
rect 1784 2793 1786 2817
rect 478 2792 484 2793
rect 110 2789 116 2790
rect 110 2785 111 2789
rect 115 2785 116 2789
rect 478 2788 479 2792
rect 483 2788 484 2792
rect 478 2787 484 2788
rect 574 2792 580 2793
rect 574 2788 575 2792
rect 579 2788 580 2792
rect 574 2787 580 2788
rect 678 2792 684 2793
rect 678 2788 679 2792
rect 683 2788 684 2792
rect 678 2787 684 2788
rect 798 2792 804 2793
rect 798 2788 799 2792
rect 803 2788 804 2792
rect 798 2787 804 2788
rect 934 2792 940 2793
rect 934 2788 935 2792
rect 939 2788 940 2792
rect 934 2787 940 2788
rect 1078 2792 1084 2793
rect 1078 2788 1079 2792
rect 1083 2788 1084 2792
rect 1078 2787 1084 2788
rect 1238 2792 1244 2793
rect 1238 2788 1239 2792
rect 1243 2788 1244 2792
rect 1238 2787 1244 2788
rect 1414 2792 1420 2793
rect 1414 2788 1415 2792
rect 1419 2788 1420 2792
rect 1414 2787 1420 2788
rect 1598 2792 1604 2793
rect 1598 2788 1599 2792
rect 1603 2788 1604 2792
rect 1598 2787 1604 2788
rect 1782 2792 1788 2793
rect 1782 2788 1783 2792
rect 1787 2788 1788 2792
rect 2008 2790 2010 2817
rect 2048 2811 2050 2835
rect 2072 2811 2074 2836
rect 2296 2811 2298 2836
rect 2536 2811 2538 2836
rect 2768 2811 2770 2836
rect 2992 2811 2994 2836
rect 3216 2811 3218 2836
rect 3432 2811 3434 2836
rect 3648 2811 3650 2836
rect 3840 2811 3842 2836
rect 3942 2835 3948 2836
rect 3944 2811 3946 2835
rect 2047 2810 2051 2811
rect 2047 2805 2051 2806
rect 2071 2810 2075 2811
rect 2071 2805 2075 2806
rect 2199 2810 2203 2811
rect 2199 2805 2203 2806
rect 2295 2810 2299 2811
rect 2295 2805 2299 2806
rect 2367 2810 2371 2811
rect 2367 2805 2371 2806
rect 2535 2810 2539 2811
rect 2535 2805 2539 2806
rect 2551 2810 2555 2811
rect 2551 2805 2555 2806
rect 2735 2810 2739 2811
rect 2735 2805 2739 2806
rect 2767 2810 2771 2811
rect 2767 2805 2771 2806
rect 2927 2810 2931 2811
rect 2927 2805 2931 2806
rect 2991 2810 2995 2811
rect 2991 2805 2995 2806
rect 3111 2810 3115 2811
rect 3111 2805 3115 2806
rect 3215 2810 3219 2811
rect 3215 2805 3219 2806
rect 3295 2810 3299 2811
rect 3295 2805 3299 2806
rect 3431 2810 3435 2811
rect 3431 2805 3435 2806
rect 3479 2810 3483 2811
rect 3479 2805 3483 2806
rect 3647 2810 3651 2811
rect 3647 2805 3651 2806
rect 3671 2810 3675 2811
rect 3671 2805 3675 2806
rect 3839 2810 3843 2811
rect 3839 2805 3843 2806
rect 3943 2810 3947 2811
rect 3943 2805 3947 2806
rect 1782 2787 1788 2788
rect 2006 2789 2012 2790
rect 110 2784 116 2785
rect 2006 2785 2007 2789
rect 2011 2785 2012 2789
rect 2048 2785 2050 2805
rect 2006 2784 2012 2785
rect 2046 2784 2052 2785
rect 2072 2784 2074 2805
rect 2200 2784 2202 2805
rect 2368 2784 2370 2805
rect 2552 2784 2554 2805
rect 2736 2784 2738 2805
rect 2928 2784 2930 2805
rect 3112 2784 3114 2805
rect 3296 2784 3298 2805
rect 3480 2784 3482 2805
rect 3672 2784 3674 2805
rect 3840 2784 3842 2805
rect 3944 2785 3946 2805
rect 3942 2784 3948 2785
rect 2046 2780 2047 2784
rect 2051 2780 2052 2784
rect 2046 2779 2052 2780
rect 2070 2783 2076 2784
rect 2070 2779 2071 2783
rect 2075 2779 2076 2783
rect 2070 2778 2076 2779
rect 2198 2783 2204 2784
rect 2198 2779 2199 2783
rect 2203 2779 2204 2783
rect 2198 2778 2204 2779
rect 2366 2783 2372 2784
rect 2366 2779 2367 2783
rect 2371 2779 2372 2783
rect 2366 2778 2372 2779
rect 2550 2783 2556 2784
rect 2550 2779 2551 2783
rect 2555 2779 2556 2783
rect 2550 2778 2556 2779
rect 2734 2783 2740 2784
rect 2734 2779 2735 2783
rect 2739 2779 2740 2783
rect 2734 2778 2740 2779
rect 2926 2783 2932 2784
rect 2926 2779 2927 2783
rect 2931 2779 2932 2783
rect 2926 2778 2932 2779
rect 3110 2783 3116 2784
rect 3110 2779 3111 2783
rect 3115 2779 3116 2783
rect 3110 2778 3116 2779
rect 3294 2783 3300 2784
rect 3294 2779 3295 2783
rect 3299 2779 3300 2783
rect 3294 2778 3300 2779
rect 3478 2783 3484 2784
rect 3478 2779 3479 2783
rect 3483 2779 3484 2783
rect 3478 2778 3484 2779
rect 3670 2783 3676 2784
rect 3670 2779 3671 2783
rect 3675 2779 3676 2783
rect 3670 2778 3676 2779
rect 3838 2783 3844 2784
rect 3838 2779 3839 2783
rect 3843 2779 3844 2783
rect 3942 2780 3943 2784
rect 3947 2780 3948 2784
rect 3942 2779 3948 2780
rect 3838 2778 3844 2779
rect 478 2773 484 2774
rect 110 2772 116 2773
rect 110 2768 111 2772
rect 115 2768 116 2772
rect 478 2769 479 2773
rect 483 2769 484 2773
rect 478 2768 484 2769
rect 574 2773 580 2774
rect 574 2769 575 2773
rect 579 2769 580 2773
rect 574 2768 580 2769
rect 678 2773 684 2774
rect 678 2769 679 2773
rect 683 2769 684 2773
rect 678 2768 684 2769
rect 798 2773 804 2774
rect 798 2769 799 2773
rect 803 2769 804 2773
rect 798 2768 804 2769
rect 934 2773 940 2774
rect 934 2769 935 2773
rect 939 2769 940 2773
rect 934 2768 940 2769
rect 1078 2773 1084 2774
rect 1078 2769 1079 2773
rect 1083 2769 1084 2773
rect 1078 2768 1084 2769
rect 1238 2773 1244 2774
rect 1238 2769 1239 2773
rect 1243 2769 1244 2773
rect 1238 2768 1244 2769
rect 1414 2773 1420 2774
rect 1414 2769 1415 2773
rect 1419 2769 1420 2773
rect 1414 2768 1420 2769
rect 1598 2773 1604 2774
rect 1598 2769 1599 2773
rect 1603 2769 1604 2773
rect 1598 2768 1604 2769
rect 1782 2773 1788 2774
rect 1782 2769 1783 2773
rect 1787 2769 1788 2773
rect 1782 2768 1788 2769
rect 2006 2772 2012 2773
rect 2006 2768 2007 2772
rect 2011 2768 2012 2772
rect 110 2767 116 2768
rect 112 2743 114 2767
rect 480 2743 482 2768
rect 576 2743 578 2768
rect 680 2743 682 2768
rect 800 2743 802 2768
rect 936 2743 938 2768
rect 1080 2743 1082 2768
rect 1240 2743 1242 2768
rect 1416 2743 1418 2768
rect 1600 2743 1602 2768
rect 1784 2743 1786 2768
rect 2006 2767 2012 2768
rect 2046 2767 2052 2768
rect 2008 2743 2010 2767
rect 2046 2763 2047 2767
rect 2051 2763 2052 2767
rect 3942 2767 3948 2768
rect 2046 2762 2052 2763
rect 2070 2764 2076 2765
rect 111 2742 115 2743
rect 111 2737 115 2738
rect 479 2742 483 2743
rect 479 2737 483 2738
rect 511 2742 515 2743
rect 511 2737 515 2738
rect 575 2742 579 2743
rect 575 2737 579 2738
rect 623 2742 627 2743
rect 623 2737 627 2738
rect 679 2742 683 2743
rect 679 2737 683 2738
rect 743 2742 747 2743
rect 743 2737 747 2738
rect 799 2742 803 2743
rect 799 2737 803 2738
rect 879 2742 883 2743
rect 879 2737 883 2738
rect 935 2742 939 2743
rect 935 2737 939 2738
rect 1015 2742 1019 2743
rect 1015 2737 1019 2738
rect 1079 2742 1083 2743
rect 1079 2737 1083 2738
rect 1159 2742 1163 2743
rect 1159 2737 1163 2738
rect 1239 2742 1243 2743
rect 1239 2737 1243 2738
rect 1311 2742 1315 2743
rect 1311 2737 1315 2738
rect 1415 2742 1419 2743
rect 1415 2737 1419 2738
rect 1463 2742 1467 2743
rect 1463 2737 1467 2738
rect 1599 2742 1603 2743
rect 1599 2737 1603 2738
rect 1623 2742 1627 2743
rect 1623 2737 1627 2738
rect 1783 2742 1787 2743
rect 1783 2737 1787 2738
rect 2007 2742 2011 2743
rect 2007 2737 2011 2738
rect 112 2717 114 2737
rect 110 2716 116 2717
rect 512 2716 514 2737
rect 624 2716 626 2737
rect 744 2716 746 2737
rect 880 2716 882 2737
rect 1016 2716 1018 2737
rect 1160 2716 1162 2737
rect 1312 2716 1314 2737
rect 1464 2716 1466 2737
rect 1624 2716 1626 2737
rect 1784 2716 1786 2737
rect 2008 2717 2010 2737
rect 2048 2731 2050 2762
rect 2070 2760 2071 2764
rect 2075 2760 2076 2764
rect 2070 2759 2076 2760
rect 2198 2764 2204 2765
rect 2198 2760 2199 2764
rect 2203 2760 2204 2764
rect 2198 2759 2204 2760
rect 2366 2764 2372 2765
rect 2366 2760 2367 2764
rect 2371 2760 2372 2764
rect 2366 2759 2372 2760
rect 2550 2764 2556 2765
rect 2550 2760 2551 2764
rect 2555 2760 2556 2764
rect 2550 2759 2556 2760
rect 2734 2764 2740 2765
rect 2734 2760 2735 2764
rect 2739 2760 2740 2764
rect 2734 2759 2740 2760
rect 2926 2764 2932 2765
rect 2926 2760 2927 2764
rect 2931 2760 2932 2764
rect 2926 2759 2932 2760
rect 3110 2764 3116 2765
rect 3110 2760 3111 2764
rect 3115 2760 3116 2764
rect 3110 2759 3116 2760
rect 3294 2764 3300 2765
rect 3294 2760 3295 2764
rect 3299 2760 3300 2764
rect 3294 2759 3300 2760
rect 3478 2764 3484 2765
rect 3478 2760 3479 2764
rect 3483 2760 3484 2764
rect 3478 2759 3484 2760
rect 3670 2764 3676 2765
rect 3670 2760 3671 2764
rect 3675 2760 3676 2764
rect 3670 2759 3676 2760
rect 3838 2764 3844 2765
rect 3838 2760 3839 2764
rect 3843 2760 3844 2764
rect 3942 2763 3943 2767
rect 3947 2763 3948 2767
rect 3942 2762 3948 2763
rect 3838 2759 3844 2760
rect 2072 2731 2074 2759
rect 2200 2731 2202 2759
rect 2368 2731 2370 2759
rect 2552 2731 2554 2759
rect 2736 2731 2738 2759
rect 2928 2731 2930 2759
rect 3112 2731 3114 2759
rect 3296 2731 3298 2759
rect 3480 2731 3482 2759
rect 3672 2731 3674 2759
rect 3840 2731 3842 2759
rect 3944 2731 3946 2762
rect 2047 2730 2051 2731
rect 2047 2725 2051 2726
rect 2071 2730 2075 2731
rect 2071 2725 2075 2726
rect 2191 2730 2195 2731
rect 2191 2725 2195 2726
rect 2199 2730 2203 2731
rect 2199 2725 2203 2726
rect 2319 2730 2323 2731
rect 2319 2725 2323 2726
rect 2367 2730 2371 2731
rect 2367 2725 2371 2726
rect 2447 2730 2451 2731
rect 2447 2725 2451 2726
rect 2551 2730 2555 2731
rect 2551 2725 2555 2726
rect 2583 2730 2587 2731
rect 2583 2725 2587 2726
rect 2727 2730 2731 2731
rect 2727 2725 2731 2726
rect 2735 2730 2739 2731
rect 2735 2725 2739 2726
rect 2887 2730 2891 2731
rect 2887 2725 2891 2726
rect 2927 2730 2931 2731
rect 2927 2725 2931 2726
rect 3063 2730 3067 2731
rect 3063 2725 3067 2726
rect 3111 2730 3115 2731
rect 3111 2725 3115 2726
rect 3255 2730 3259 2731
rect 3255 2725 3259 2726
rect 3295 2730 3299 2731
rect 3295 2725 3299 2726
rect 3455 2730 3459 2731
rect 3455 2725 3459 2726
rect 3479 2730 3483 2731
rect 3479 2725 3483 2726
rect 3655 2730 3659 2731
rect 3655 2725 3659 2726
rect 3671 2730 3675 2731
rect 3671 2725 3675 2726
rect 3839 2730 3843 2731
rect 3839 2725 3843 2726
rect 3943 2730 3947 2731
rect 3943 2725 3947 2726
rect 2006 2716 2012 2717
rect 110 2712 111 2716
rect 115 2712 116 2716
rect 110 2711 116 2712
rect 510 2715 516 2716
rect 510 2711 511 2715
rect 515 2711 516 2715
rect 510 2710 516 2711
rect 622 2715 628 2716
rect 622 2711 623 2715
rect 627 2711 628 2715
rect 622 2710 628 2711
rect 742 2715 748 2716
rect 742 2711 743 2715
rect 747 2711 748 2715
rect 742 2710 748 2711
rect 878 2715 884 2716
rect 878 2711 879 2715
rect 883 2711 884 2715
rect 878 2710 884 2711
rect 1014 2715 1020 2716
rect 1014 2711 1015 2715
rect 1019 2711 1020 2715
rect 1014 2710 1020 2711
rect 1158 2715 1164 2716
rect 1158 2711 1159 2715
rect 1163 2711 1164 2715
rect 1158 2710 1164 2711
rect 1310 2715 1316 2716
rect 1310 2711 1311 2715
rect 1315 2711 1316 2715
rect 1310 2710 1316 2711
rect 1462 2715 1468 2716
rect 1462 2711 1463 2715
rect 1467 2711 1468 2715
rect 1462 2710 1468 2711
rect 1622 2715 1628 2716
rect 1622 2711 1623 2715
rect 1627 2711 1628 2715
rect 1622 2710 1628 2711
rect 1782 2715 1788 2716
rect 1782 2711 1783 2715
rect 1787 2711 1788 2715
rect 2006 2712 2007 2716
rect 2011 2712 2012 2716
rect 2006 2711 2012 2712
rect 1782 2710 1788 2711
rect 110 2699 116 2700
rect 110 2695 111 2699
rect 115 2695 116 2699
rect 2006 2699 2012 2700
rect 110 2694 116 2695
rect 510 2696 516 2697
rect 112 2663 114 2694
rect 510 2692 511 2696
rect 515 2692 516 2696
rect 510 2691 516 2692
rect 622 2696 628 2697
rect 622 2692 623 2696
rect 627 2692 628 2696
rect 622 2691 628 2692
rect 742 2696 748 2697
rect 742 2692 743 2696
rect 747 2692 748 2696
rect 742 2691 748 2692
rect 878 2696 884 2697
rect 878 2692 879 2696
rect 883 2692 884 2696
rect 878 2691 884 2692
rect 1014 2696 1020 2697
rect 1014 2692 1015 2696
rect 1019 2692 1020 2696
rect 1014 2691 1020 2692
rect 1158 2696 1164 2697
rect 1158 2692 1159 2696
rect 1163 2692 1164 2696
rect 1158 2691 1164 2692
rect 1310 2696 1316 2697
rect 1310 2692 1311 2696
rect 1315 2692 1316 2696
rect 1310 2691 1316 2692
rect 1462 2696 1468 2697
rect 1462 2692 1463 2696
rect 1467 2692 1468 2696
rect 1462 2691 1468 2692
rect 1622 2696 1628 2697
rect 1622 2692 1623 2696
rect 1627 2692 1628 2696
rect 1622 2691 1628 2692
rect 1782 2696 1788 2697
rect 1782 2692 1783 2696
rect 1787 2692 1788 2696
rect 2006 2695 2007 2699
rect 2011 2695 2012 2699
rect 2048 2698 2050 2725
rect 2072 2701 2074 2725
rect 2192 2701 2194 2725
rect 2320 2701 2322 2725
rect 2448 2701 2450 2725
rect 2584 2701 2586 2725
rect 2728 2701 2730 2725
rect 2888 2701 2890 2725
rect 3064 2701 3066 2725
rect 3256 2701 3258 2725
rect 3456 2701 3458 2725
rect 3656 2701 3658 2725
rect 3840 2701 3842 2725
rect 2070 2700 2076 2701
rect 2006 2694 2012 2695
rect 2046 2697 2052 2698
rect 1782 2691 1788 2692
rect 512 2663 514 2691
rect 624 2663 626 2691
rect 744 2663 746 2691
rect 880 2663 882 2691
rect 1016 2663 1018 2691
rect 1160 2663 1162 2691
rect 1312 2663 1314 2691
rect 1464 2663 1466 2691
rect 1624 2663 1626 2691
rect 1784 2663 1786 2691
rect 2008 2663 2010 2694
rect 2046 2693 2047 2697
rect 2051 2693 2052 2697
rect 2070 2696 2071 2700
rect 2075 2696 2076 2700
rect 2070 2695 2076 2696
rect 2190 2700 2196 2701
rect 2190 2696 2191 2700
rect 2195 2696 2196 2700
rect 2190 2695 2196 2696
rect 2318 2700 2324 2701
rect 2318 2696 2319 2700
rect 2323 2696 2324 2700
rect 2318 2695 2324 2696
rect 2446 2700 2452 2701
rect 2446 2696 2447 2700
rect 2451 2696 2452 2700
rect 2446 2695 2452 2696
rect 2582 2700 2588 2701
rect 2582 2696 2583 2700
rect 2587 2696 2588 2700
rect 2582 2695 2588 2696
rect 2726 2700 2732 2701
rect 2726 2696 2727 2700
rect 2731 2696 2732 2700
rect 2726 2695 2732 2696
rect 2886 2700 2892 2701
rect 2886 2696 2887 2700
rect 2891 2696 2892 2700
rect 2886 2695 2892 2696
rect 3062 2700 3068 2701
rect 3062 2696 3063 2700
rect 3067 2696 3068 2700
rect 3062 2695 3068 2696
rect 3254 2700 3260 2701
rect 3254 2696 3255 2700
rect 3259 2696 3260 2700
rect 3254 2695 3260 2696
rect 3454 2700 3460 2701
rect 3454 2696 3455 2700
rect 3459 2696 3460 2700
rect 3454 2695 3460 2696
rect 3654 2700 3660 2701
rect 3654 2696 3655 2700
rect 3659 2696 3660 2700
rect 3654 2695 3660 2696
rect 3838 2700 3844 2701
rect 3838 2696 3839 2700
rect 3843 2696 3844 2700
rect 3944 2698 3946 2725
rect 3838 2695 3844 2696
rect 3942 2697 3948 2698
rect 2046 2692 2052 2693
rect 3942 2693 3943 2697
rect 3947 2693 3948 2697
rect 3942 2692 3948 2693
rect 2070 2681 2076 2682
rect 2046 2680 2052 2681
rect 2046 2676 2047 2680
rect 2051 2676 2052 2680
rect 2070 2677 2071 2681
rect 2075 2677 2076 2681
rect 2070 2676 2076 2677
rect 2190 2681 2196 2682
rect 2190 2677 2191 2681
rect 2195 2677 2196 2681
rect 2190 2676 2196 2677
rect 2318 2681 2324 2682
rect 2318 2677 2319 2681
rect 2323 2677 2324 2681
rect 2318 2676 2324 2677
rect 2446 2681 2452 2682
rect 2446 2677 2447 2681
rect 2451 2677 2452 2681
rect 2446 2676 2452 2677
rect 2582 2681 2588 2682
rect 2582 2677 2583 2681
rect 2587 2677 2588 2681
rect 2582 2676 2588 2677
rect 2726 2681 2732 2682
rect 2726 2677 2727 2681
rect 2731 2677 2732 2681
rect 2726 2676 2732 2677
rect 2886 2681 2892 2682
rect 2886 2677 2887 2681
rect 2891 2677 2892 2681
rect 2886 2676 2892 2677
rect 3062 2681 3068 2682
rect 3062 2677 3063 2681
rect 3067 2677 3068 2681
rect 3062 2676 3068 2677
rect 3254 2681 3260 2682
rect 3254 2677 3255 2681
rect 3259 2677 3260 2681
rect 3254 2676 3260 2677
rect 3454 2681 3460 2682
rect 3454 2677 3455 2681
rect 3459 2677 3460 2681
rect 3454 2676 3460 2677
rect 3654 2681 3660 2682
rect 3654 2677 3655 2681
rect 3659 2677 3660 2681
rect 3654 2676 3660 2677
rect 3838 2681 3844 2682
rect 3838 2677 3839 2681
rect 3843 2677 3844 2681
rect 3838 2676 3844 2677
rect 3942 2680 3948 2681
rect 3942 2676 3943 2680
rect 3947 2676 3948 2680
rect 2046 2675 2052 2676
rect 111 2662 115 2663
rect 111 2657 115 2658
rect 367 2662 371 2663
rect 367 2657 371 2658
rect 487 2662 491 2663
rect 487 2657 491 2658
rect 511 2662 515 2663
rect 511 2657 515 2658
rect 615 2662 619 2663
rect 615 2657 619 2658
rect 623 2662 627 2663
rect 623 2657 627 2658
rect 743 2662 747 2663
rect 743 2657 747 2658
rect 751 2662 755 2663
rect 751 2657 755 2658
rect 879 2662 883 2663
rect 879 2657 883 2658
rect 895 2662 899 2663
rect 895 2657 899 2658
rect 1015 2662 1019 2663
rect 1015 2657 1019 2658
rect 1031 2662 1035 2663
rect 1031 2657 1035 2658
rect 1159 2662 1163 2663
rect 1159 2657 1163 2658
rect 1167 2662 1171 2663
rect 1167 2657 1171 2658
rect 1303 2662 1307 2663
rect 1303 2657 1307 2658
rect 1311 2662 1315 2663
rect 1311 2657 1315 2658
rect 1431 2662 1435 2663
rect 1431 2657 1435 2658
rect 1463 2662 1467 2663
rect 1463 2657 1467 2658
rect 1567 2662 1571 2663
rect 1567 2657 1571 2658
rect 1623 2662 1627 2663
rect 1623 2657 1627 2658
rect 1703 2662 1707 2663
rect 1703 2657 1707 2658
rect 1783 2662 1787 2663
rect 1783 2657 1787 2658
rect 2007 2662 2011 2663
rect 2007 2657 2011 2658
rect 112 2630 114 2657
rect 368 2633 370 2657
rect 488 2633 490 2657
rect 616 2633 618 2657
rect 752 2633 754 2657
rect 896 2633 898 2657
rect 1032 2633 1034 2657
rect 1168 2633 1170 2657
rect 1304 2633 1306 2657
rect 1432 2633 1434 2657
rect 1568 2633 1570 2657
rect 1704 2633 1706 2657
rect 366 2632 372 2633
rect 110 2629 116 2630
rect 110 2625 111 2629
rect 115 2625 116 2629
rect 366 2628 367 2632
rect 371 2628 372 2632
rect 366 2627 372 2628
rect 486 2632 492 2633
rect 486 2628 487 2632
rect 491 2628 492 2632
rect 486 2627 492 2628
rect 614 2632 620 2633
rect 614 2628 615 2632
rect 619 2628 620 2632
rect 614 2627 620 2628
rect 750 2632 756 2633
rect 750 2628 751 2632
rect 755 2628 756 2632
rect 750 2627 756 2628
rect 894 2632 900 2633
rect 894 2628 895 2632
rect 899 2628 900 2632
rect 894 2627 900 2628
rect 1030 2632 1036 2633
rect 1030 2628 1031 2632
rect 1035 2628 1036 2632
rect 1030 2627 1036 2628
rect 1166 2632 1172 2633
rect 1166 2628 1167 2632
rect 1171 2628 1172 2632
rect 1166 2627 1172 2628
rect 1302 2632 1308 2633
rect 1302 2628 1303 2632
rect 1307 2628 1308 2632
rect 1302 2627 1308 2628
rect 1430 2632 1436 2633
rect 1430 2628 1431 2632
rect 1435 2628 1436 2632
rect 1430 2627 1436 2628
rect 1566 2632 1572 2633
rect 1566 2628 1567 2632
rect 1571 2628 1572 2632
rect 1566 2627 1572 2628
rect 1702 2632 1708 2633
rect 1702 2628 1703 2632
rect 1707 2628 1708 2632
rect 2008 2630 2010 2657
rect 2048 2647 2050 2675
rect 2072 2647 2074 2676
rect 2192 2647 2194 2676
rect 2320 2647 2322 2676
rect 2448 2647 2450 2676
rect 2584 2647 2586 2676
rect 2728 2647 2730 2676
rect 2888 2647 2890 2676
rect 3064 2647 3066 2676
rect 3256 2647 3258 2676
rect 3456 2647 3458 2676
rect 3656 2647 3658 2676
rect 3840 2647 3842 2676
rect 3942 2675 3948 2676
rect 3944 2647 3946 2675
rect 2047 2646 2051 2647
rect 2047 2641 2051 2642
rect 2071 2646 2075 2647
rect 2071 2641 2075 2642
rect 2191 2646 2195 2647
rect 2191 2641 2195 2642
rect 2231 2646 2235 2647
rect 2231 2641 2235 2642
rect 2319 2646 2323 2647
rect 2319 2641 2323 2642
rect 2335 2646 2339 2647
rect 2335 2641 2339 2642
rect 2447 2646 2451 2647
rect 2447 2641 2451 2642
rect 2559 2646 2563 2647
rect 2559 2641 2563 2642
rect 2583 2646 2587 2647
rect 2583 2641 2587 2642
rect 2671 2646 2675 2647
rect 2671 2641 2675 2642
rect 2727 2646 2731 2647
rect 2727 2641 2731 2642
rect 2791 2646 2795 2647
rect 2791 2641 2795 2642
rect 2887 2646 2891 2647
rect 2887 2641 2891 2642
rect 2911 2646 2915 2647
rect 2911 2641 2915 2642
rect 3031 2646 3035 2647
rect 3031 2641 3035 2642
rect 3063 2646 3067 2647
rect 3063 2641 3067 2642
rect 3151 2646 3155 2647
rect 3151 2641 3155 2642
rect 3255 2646 3259 2647
rect 3255 2641 3259 2642
rect 3455 2646 3459 2647
rect 3455 2641 3459 2642
rect 3655 2646 3659 2647
rect 3655 2641 3659 2642
rect 3839 2646 3843 2647
rect 3839 2641 3843 2642
rect 3943 2646 3947 2647
rect 3943 2641 3947 2642
rect 1702 2627 1708 2628
rect 2006 2629 2012 2630
rect 110 2624 116 2625
rect 2006 2625 2007 2629
rect 2011 2625 2012 2629
rect 2006 2624 2012 2625
rect 2048 2621 2050 2641
rect 2046 2620 2052 2621
rect 2232 2620 2234 2641
rect 2336 2620 2338 2641
rect 2448 2620 2450 2641
rect 2560 2620 2562 2641
rect 2672 2620 2674 2641
rect 2792 2620 2794 2641
rect 2912 2620 2914 2641
rect 3032 2620 3034 2641
rect 3152 2620 3154 2641
rect 3944 2621 3946 2641
rect 3942 2620 3948 2621
rect 2046 2616 2047 2620
rect 2051 2616 2052 2620
rect 2046 2615 2052 2616
rect 2230 2619 2236 2620
rect 2230 2615 2231 2619
rect 2235 2615 2236 2619
rect 2230 2614 2236 2615
rect 2334 2619 2340 2620
rect 2334 2615 2335 2619
rect 2339 2615 2340 2619
rect 2334 2614 2340 2615
rect 2446 2619 2452 2620
rect 2446 2615 2447 2619
rect 2451 2615 2452 2619
rect 2446 2614 2452 2615
rect 2558 2619 2564 2620
rect 2558 2615 2559 2619
rect 2563 2615 2564 2619
rect 2558 2614 2564 2615
rect 2670 2619 2676 2620
rect 2670 2615 2671 2619
rect 2675 2615 2676 2619
rect 2670 2614 2676 2615
rect 2790 2619 2796 2620
rect 2790 2615 2791 2619
rect 2795 2615 2796 2619
rect 2790 2614 2796 2615
rect 2910 2619 2916 2620
rect 2910 2615 2911 2619
rect 2915 2615 2916 2619
rect 2910 2614 2916 2615
rect 3030 2619 3036 2620
rect 3030 2615 3031 2619
rect 3035 2615 3036 2619
rect 3030 2614 3036 2615
rect 3150 2619 3156 2620
rect 3150 2615 3151 2619
rect 3155 2615 3156 2619
rect 3942 2616 3943 2620
rect 3947 2616 3948 2620
rect 3942 2615 3948 2616
rect 3150 2614 3156 2615
rect 366 2613 372 2614
rect 110 2612 116 2613
rect 110 2608 111 2612
rect 115 2608 116 2612
rect 366 2609 367 2613
rect 371 2609 372 2613
rect 366 2608 372 2609
rect 486 2613 492 2614
rect 486 2609 487 2613
rect 491 2609 492 2613
rect 486 2608 492 2609
rect 614 2613 620 2614
rect 614 2609 615 2613
rect 619 2609 620 2613
rect 614 2608 620 2609
rect 750 2613 756 2614
rect 750 2609 751 2613
rect 755 2609 756 2613
rect 750 2608 756 2609
rect 894 2613 900 2614
rect 894 2609 895 2613
rect 899 2609 900 2613
rect 894 2608 900 2609
rect 1030 2613 1036 2614
rect 1030 2609 1031 2613
rect 1035 2609 1036 2613
rect 1030 2608 1036 2609
rect 1166 2613 1172 2614
rect 1166 2609 1167 2613
rect 1171 2609 1172 2613
rect 1166 2608 1172 2609
rect 1302 2613 1308 2614
rect 1302 2609 1303 2613
rect 1307 2609 1308 2613
rect 1302 2608 1308 2609
rect 1430 2613 1436 2614
rect 1430 2609 1431 2613
rect 1435 2609 1436 2613
rect 1430 2608 1436 2609
rect 1566 2613 1572 2614
rect 1566 2609 1567 2613
rect 1571 2609 1572 2613
rect 1566 2608 1572 2609
rect 1702 2613 1708 2614
rect 1702 2609 1703 2613
rect 1707 2609 1708 2613
rect 1702 2608 1708 2609
rect 2006 2612 2012 2613
rect 2006 2608 2007 2612
rect 2011 2608 2012 2612
rect 110 2607 116 2608
rect 112 2587 114 2607
rect 368 2587 370 2608
rect 488 2587 490 2608
rect 616 2587 618 2608
rect 752 2587 754 2608
rect 896 2587 898 2608
rect 1032 2587 1034 2608
rect 1168 2587 1170 2608
rect 1304 2587 1306 2608
rect 1432 2587 1434 2608
rect 1568 2587 1570 2608
rect 1704 2587 1706 2608
rect 2006 2607 2012 2608
rect 2008 2587 2010 2607
rect 2046 2603 2052 2604
rect 2046 2599 2047 2603
rect 2051 2599 2052 2603
rect 3942 2603 3948 2604
rect 2046 2598 2052 2599
rect 2230 2600 2236 2601
rect 111 2586 115 2587
rect 111 2581 115 2582
rect 135 2586 139 2587
rect 135 2581 139 2582
rect 287 2586 291 2587
rect 287 2581 291 2582
rect 367 2586 371 2587
rect 367 2581 371 2582
rect 447 2586 451 2587
rect 447 2581 451 2582
rect 487 2586 491 2587
rect 487 2581 491 2582
rect 607 2586 611 2587
rect 607 2581 611 2582
rect 615 2586 619 2587
rect 615 2581 619 2582
rect 751 2586 755 2587
rect 751 2581 755 2582
rect 767 2586 771 2587
rect 767 2581 771 2582
rect 895 2586 899 2587
rect 895 2581 899 2582
rect 919 2586 923 2587
rect 919 2581 923 2582
rect 1031 2586 1035 2587
rect 1031 2581 1035 2582
rect 1063 2586 1067 2587
rect 1063 2581 1067 2582
rect 1167 2586 1171 2587
rect 1167 2581 1171 2582
rect 1199 2586 1203 2587
rect 1199 2581 1203 2582
rect 1303 2586 1307 2587
rect 1303 2581 1307 2582
rect 1335 2586 1339 2587
rect 1335 2581 1339 2582
rect 1431 2586 1435 2587
rect 1431 2581 1435 2582
rect 1463 2586 1467 2587
rect 1463 2581 1467 2582
rect 1567 2586 1571 2587
rect 1567 2581 1571 2582
rect 1591 2586 1595 2587
rect 1591 2581 1595 2582
rect 1703 2586 1707 2587
rect 1703 2581 1707 2582
rect 1727 2586 1731 2587
rect 1727 2581 1731 2582
rect 2007 2586 2011 2587
rect 2007 2581 2011 2582
rect 112 2561 114 2581
rect 110 2560 116 2561
rect 136 2560 138 2581
rect 288 2560 290 2581
rect 448 2560 450 2581
rect 608 2560 610 2581
rect 768 2560 770 2581
rect 920 2560 922 2581
rect 1064 2560 1066 2581
rect 1200 2560 1202 2581
rect 1336 2560 1338 2581
rect 1464 2560 1466 2581
rect 1592 2560 1594 2581
rect 1728 2560 1730 2581
rect 2008 2561 2010 2581
rect 2048 2567 2050 2598
rect 2230 2596 2231 2600
rect 2235 2596 2236 2600
rect 2230 2595 2236 2596
rect 2334 2600 2340 2601
rect 2334 2596 2335 2600
rect 2339 2596 2340 2600
rect 2334 2595 2340 2596
rect 2446 2600 2452 2601
rect 2446 2596 2447 2600
rect 2451 2596 2452 2600
rect 2446 2595 2452 2596
rect 2558 2600 2564 2601
rect 2558 2596 2559 2600
rect 2563 2596 2564 2600
rect 2558 2595 2564 2596
rect 2670 2600 2676 2601
rect 2670 2596 2671 2600
rect 2675 2596 2676 2600
rect 2670 2595 2676 2596
rect 2790 2600 2796 2601
rect 2790 2596 2791 2600
rect 2795 2596 2796 2600
rect 2790 2595 2796 2596
rect 2910 2600 2916 2601
rect 2910 2596 2911 2600
rect 2915 2596 2916 2600
rect 2910 2595 2916 2596
rect 3030 2600 3036 2601
rect 3030 2596 3031 2600
rect 3035 2596 3036 2600
rect 3030 2595 3036 2596
rect 3150 2600 3156 2601
rect 3150 2596 3151 2600
rect 3155 2596 3156 2600
rect 3942 2599 3943 2603
rect 3947 2599 3948 2603
rect 3942 2598 3948 2599
rect 3150 2595 3156 2596
rect 2232 2567 2234 2595
rect 2336 2567 2338 2595
rect 2448 2567 2450 2595
rect 2560 2567 2562 2595
rect 2672 2567 2674 2595
rect 2792 2567 2794 2595
rect 2912 2567 2914 2595
rect 3032 2567 3034 2595
rect 3152 2567 3154 2595
rect 3944 2567 3946 2598
rect 2047 2566 2051 2567
rect 2047 2561 2051 2562
rect 2231 2566 2235 2567
rect 2231 2561 2235 2562
rect 2335 2566 2339 2567
rect 2335 2561 2339 2562
rect 2383 2566 2387 2567
rect 2383 2561 2387 2562
rect 2447 2566 2451 2567
rect 2447 2561 2451 2562
rect 2495 2566 2499 2567
rect 2495 2561 2499 2562
rect 2559 2566 2563 2567
rect 2559 2561 2563 2562
rect 2615 2566 2619 2567
rect 2615 2561 2619 2562
rect 2671 2566 2675 2567
rect 2671 2561 2675 2562
rect 2743 2566 2747 2567
rect 2743 2561 2747 2562
rect 2791 2566 2795 2567
rect 2791 2561 2795 2562
rect 2871 2566 2875 2567
rect 2871 2561 2875 2562
rect 2911 2566 2915 2567
rect 2911 2561 2915 2562
rect 2991 2566 2995 2567
rect 2991 2561 2995 2562
rect 3031 2566 3035 2567
rect 3031 2561 3035 2562
rect 3111 2566 3115 2567
rect 3111 2561 3115 2562
rect 3151 2566 3155 2567
rect 3151 2561 3155 2562
rect 3231 2566 3235 2567
rect 3231 2561 3235 2562
rect 3359 2566 3363 2567
rect 3359 2561 3363 2562
rect 3487 2566 3491 2567
rect 3487 2561 3491 2562
rect 3943 2566 3947 2567
rect 3943 2561 3947 2562
rect 2006 2560 2012 2561
rect 110 2556 111 2560
rect 115 2556 116 2560
rect 110 2555 116 2556
rect 134 2559 140 2560
rect 134 2555 135 2559
rect 139 2555 140 2559
rect 134 2554 140 2555
rect 286 2559 292 2560
rect 286 2555 287 2559
rect 291 2555 292 2559
rect 286 2554 292 2555
rect 446 2559 452 2560
rect 446 2555 447 2559
rect 451 2555 452 2559
rect 446 2554 452 2555
rect 606 2559 612 2560
rect 606 2555 607 2559
rect 611 2555 612 2559
rect 606 2554 612 2555
rect 766 2559 772 2560
rect 766 2555 767 2559
rect 771 2555 772 2559
rect 766 2554 772 2555
rect 918 2559 924 2560
rect 918 2555 919 2559
rect 923 2555 924 2559
rect 918 2554 924 2555
rect 1062 2559 1068 2560
rect 1062 2555 1063 2559
rect 1067 2555 1068 2559
rect 1062 2554 1068 2555
rect 1198 2559 1204 2560
rect 1198 2555 1199 2559
rect 1203 2555 1204 2559
rect 1198 2554 1204 2555
rect 1334 2559 1340 2560
rect 1334 2555 1335 2559
rect 1339 2555 1340 2559
rect 1334 2554 1340 2555
rect 1462 2559 1468 2560
rect 1462 2555 1463 2559
rect 1467 2555 1468 2559
rect 1462 2554 1468 2555
rect 1590 2559 1596 2560
rect 1590 2555 1591 2559
rect 1595 2555 1596 2559
rect 1590 2554 1596 2555
rect 1726 2559 1732 2560
rect 1726 2555 1727 2559
rect 1731 2555 1732 2559
rect 2006 2556 2007 2560
rect 2011 2556 2012 2560
rect 2006 2555 2012 2556
rect 1726 2554 1732 2555
rect 110 2543 116 2544
rect 110 2539 111 2543
rect 115 2539 116 2543
rect 2006 2543 2012 2544
rect 110 2538 116 2539
rect 134 2540 140 2541
rect 112 2495 114 2538
rect 134 2536 135 2540
rect 139 2536 140 2540
rect 134 2535 140 2536
rect 286 2540 292 2541
rect 286 2536 287 2540
rect 291 2536 292 2540
rect 286 2535 292 2536
rect 446 2540 452 2541
rect 446 2536 447 2540
rect 451 2536 452 2540
rect 446 2535 452 2536
rect 606 2540 612 2541
rect 606 2536 607 2540
rect 611 2536 612 2540
rect 606 2535 612 2536
rect 766 2540 772 2541
rect 766 2536 767 2540
rect 771 2536 772 2540
rect 766 2535 772 2536
rect 918 2540 924 2541
rect 918 2536 919 2540
rect 923 2536 924 2540
rect 918 2535 924 2536
rect 1062 2540 1068 2541
rect 1062 2536 1063 2540
rect 1067 2536 1068 2540
rect 1062 2535 1068 2536
rect 1198 2540 1204 2541
rect 1198 2536 1199 2540
rect 1203 2536 1204 2540
rect 1198 2535 1204 2536
rect 1334 2540 1340 2541
rect 1334 2536 1335 2540
rect 1339 2536 1340 2540
rect 1334 2535 1340 2536
rect 1462 2540 1468 2541
rect 1462 2536 1463 2540
rect 1467 2536 1468 2540
rect 1462 2535 1468 2536
rect 1590 2540 1596 2541
rect 1590 2536 1591 2540
rect 1595 2536 1596 2540
rect 1590 2535 1596 2536
rect 1726 2540 1732 2541
rect 1726 2536 1727 2540
rect 1731 2536 1732 2540
rect 2006 2539 2007 2543
rect 2011 2539 2012 2543
rect 2006 2538 2012 2539
rect 1726 2535 1732 2536
rect 136 2495 138 2535
rect 288 2495 290 2535
rect 448 2495 450 2535
rect 608 2495 610 2535
rect 768 2495 770 2535
rect 920 2495 922 2535
rect 1064 2495 1066 2535
rect 1200 2495 1202 2535
rect 1336 2495 1338 2535
rect 1464 2495 1466 2535
rect 1592 2495 1594 2535
rect 1728 2495 1730 2535
rect 2008 2495 2010 2538
rect 2048 2534 2050 2561
rect 2384 2537 2386 2561
rect 2496 2537 2498 2561
rect 2616 2537 2618 2561
rect 2744 2537 2746 2561
rect 2872 2537 2874 2561
rect 2992 2537 2994 2561
rect 3112 2537 3114 2561
rect 3232 2537 3234 2561
rect 3360 2537 3362 2561
rect 3488 2537 3490 2561
rect 2382 2536 2388 2537
rect 2046 2533 2052 2534
rect 2046 2529 2047 2533
rect 2051 2529 2052 2533
rect 2382 2532 2383 2536
rect 2387 2532 2388 2536
rect 2382 2531 2388 2532
rect 2494 2536 2500 2537
rect 2494 2532 2495 2536
rect 2499 2532 2500 2536
rect 2494 2531 2500 2532
rect 2614 2536 2620 2537
rect 2614 2532 2615 2536
rect 2619 2532 2620 2536
rect 2614 2531 2620 2532
rect 2742 2536 2748 2537
rect 2742 2532 2743 2536
rect 2747 2532 2748 2536
rect 2742 2531 2748 2532
rect 2870 2536 2876 2537
rect 2870 2532 2871 2536
rect 2875 2532 2876 2536
rect 2870 2531 2876 2532
rect 2990 2536 2996 2537
rect 2990 2532 2991 2536
rect 2995 2532 2996 2536
rect 2990 2531 2996 2532
rect 3110 2536 3116 2537
rect 3110 2532 3111 2536
rect 3115 2532 3116 2536
rect 3110 2531 3116 2532
rect 3230 2536 3236 2537
rect 3230 2532 3231 2536
rect 3235 2532 3236 2536
rect 3230 2531 3236 2532
rect 3358 2536 3364 2537
rect 3358 2532 3359 2536
rect 3363 2532 3364 2536
rect 3358 2531 3364 2532
rect 3486 2536 3492 2537
rect 3486 2532 3487 2536
rect 3491 2532 3492 2536
rect 3944 2534 3946 2561
rect 3486 2531 3492 2532
rect 3942 2533 3948 2534
rect 2046 2528 2052 2529
rect 3942 2529 3943 2533
rect 3947 2529 3948 2533
rect 3942 2528 3948 2529
rect 2382 2517 2388 2518
rect 2046 2516 2052 2517
rect 2046 2512 2047 2516
rect 2051 2512 2052 2516
rect 2382 2513 2383 2517
rect 2387 2513 2388 2517
rect 2382 2512 2388 2513
rect 2494 2517 2500 2518
rect 2494 2513 2495 2517
rect 2499 2513 2500 2517
rect 2494 2512 2500 2513
rect 2614 2517 2620 2518
rect 2614 2513 2615 2517
rect 2619 2513 2620 2517
rect 2614 2512 2620 2513
rect 2742 2517 2748 2518
rect 2742 2513 2743 2517
rect 2747 2513 2748 2517
rect 2742 2512 2748 2513
rect 2870 2517 2876 2518
rect 2870 2513 2871 2517
rect 2875 2513 2876 2517
rect 2870 2512 2876 2513
rect 2990 2517 2996 2518
rect 2990 2513 2991 2517
rect 2995 2513 2996 2517
rect 2990 2512 2996 2513
rect 3110 2517 3116 2518
rect 3110 2513 3111 2517
rect 3115 2513 3116 2517
rect 3110 2512 3116 2513
rect 3230 2517 3236 2518
rect 3230 2513 3231 2517
rect 3235 2513 3236 2517
rect 3230 2512 3236 2513
rect 3358 2517 3364 2518
rect 3358 2513 3359 2517
rect 3363 2513 3364 2517
rect 3358 2512 3364 2513
rect 3486 2517 3492 2518
rect 3486 2513 3487 2517
rect 3491 2513 3492 2517
rect 3486 2512 3492 2513
rect 3942 2516 3948 2517
rect 3942 2512 3943 2516
rect 3947 2512 3948 2516
rect 2046 2511 2052 2512
rect 111 2494 115 2495
rect 111 2489 115 2490
rect 135 2494 139 2495
rect 135 2489 139 2490
rect 231 2494 235 2495
rect 231 2489 235 2490
rect 287 2494 291 2495
rect 287 2489 291 2490
rect 327 2494 331 2495
rect 327 2489 331 2490
rect 423 2494 427 2495
rect 423 2489 427 2490
rect 447 2494 451 2495
rect 447 2489 451 2490
rect 519 2494 523 2495
rect 519 2489 523 2490
rect 607 2494 611 2495
rect 607 2489 611 2490
rect 767 2494 771 2495
rect 767 2489 771 2490
rect 919 2494 923 2495
rect 919 2489 923 2490
rect 1063 2494 1067 2495
rect 1063 2489 1067 2490
rect 1199 2494 1203 2495
rect 1199 2489 1203 2490
rect 1335 2494 1339 2495
rect 1335 2489 1339 2490
rect 1463 2494 1467 2495
rect 1463 2489 1467 2490
rect 1591 2494 1595 2495
rect 1591 2489 1595 2490
rect 1727 2494 1731 2495
rect 1727 2489 1731 2490
rect 2007 2494 2011 2495
rect 2007 2489 2011 2490
rect 112 2462 114 2489
rect 136 2465 138 2489
rect 232 2465 234 2489
rect 328 2465 330 2489
rect 424 2465 426 2489
rect 520 2465 522 2489
rect 134 2464 140 2465
rect 110 2461 116 2462
rect 110 2457 111 2461
rect 115 2457 116 2461
rect 134 2460 135 2464
rect 139 2460 140 2464
rect 134 2459 140 2460
rect 230 2464 236 2465
rect 230 2460 231 2464
rect 235 2460 236 2464
rect 230 2459 236 2460
rect 326 2464 332 2465
rect 326 2460 327 2464
rect 331 2460 332 2464
rect 326 2459 332 2460
rect 422 2464 428 2465
rect 422 2460 423 2464
rect 427 2460 428 2464
rect 422 2459 428 2460
rect 518 2464 524 2465
rect 518 2460 519 2464
rect 523 2460 524 2464
rect 2008 2462 2010 2489
rect 2048 2487 2050 2511
rect 2384 2487 2386 2512
rect 2496 2487 2498 2512
rect 2616 2487 2618 2512
rect 2744 2487 2746 2512
rect 2872 2487 2874 2512
rect 2992 2487 2994 2512
rect 3112 2487 3114 2512
rect 3232 2487 3234 2512
rect 3360 2487 3362 2512
rect 3488 2487 3490 2512
rect 3942 2511 3948 2512
rect 3944 2487 3946 2511
rect 2047 2486 2051 2487
rect 2047 2481 2051 2482
rect 2383 2486 2387 2487
rect 2383 2481 2387 2482
rect 2495 2486 2499 2487
rect 2495 2481 2499 2482
rect 2535 2486 2539 2487
rect 2535 2481 2539 2482
rect 2615 2486 2619 2487
rect 2615 2481 2619 2482
rect 2711 2486 2715 2487
rect 2711 2481 2715 2482
rect 2743 2486 2747 2487
rect 2743 2481 2747 2482
rect 2871 2486 2875 2487
rect 2871 2481 2875 2482
rect 2879 2486 2883 2487
rect 2879 2481 2883 2482
rect 2991 2486 2995 2487
rect 2991 2481 2995 2482
rect 3047 2486 3051 2487
rect 3047 2481 3051 2482
rect 3111 2486 3115 2487
rect 3111 2481 3115 2482
rect 3207 2486 3211 2487
rect 3207 2481 3211 2482
rect 3231 2486 3235 2487
rect 3231 2481 3235 2482
rect 3359 2486 3363 2487
rect 3359 2481 3363 2482
rect 3487 2486 3491 2487
rect 3487 2481 3491 2482
rect 3503 2486 3507 2487
rect 3503 2481 3507 2482
rect 3655 2486 3659 2487
rect 3655 2481 3659 2482
rect 3807 2486 3811 2487
rect 3807 2481 3811 2482
rect 3943 2486 3947 2487
rect 3943 2481 3947 2482
rect 518 2459 524 2460
rect 2006 2461 2012 2462
rect 2048 2461 2050 2481
rect 110 2456 116 2457
rect 2006 2457 2007 2461
rect 2011 2457 2012 2461
rect 2006 2456 2012 2457
rect 2046 2460 2052 2461
rect 2536 2460 2538 2481
rect 2712 2460 2714 2481
rect 2880 2460 2882 2481
rect 3048 2460 3050 2481
rect 3208 2460 3210 2481
rect 3360 2460 3362 2481
rect 3504 2460 3506 2481
rect 3656 2460 3658 2481
rect 3808 2460 3810 2481
rect 3944 2461 3946 2481
rect 3942 2460 3948 2461
rect 2046 2456 2047 2460
rect 2051 2456 2052 2460
rect 2046 2455 2052 2456
rect 2534 2459 2540 2460
rect 2534 2455 2535 2459
rect 2539 2455 2540 2459
rect 2534 2454 2540 2455
rect 2710 2459 2716 2460
rect 2710 2455 2711 2459
rect 2715 2455 2716 2459
rect 2710 2454 2716 2455
rect 2878 2459 2884 2460
rect 2878 2455 2879 2459
rect 2883 2455 2884 2459
rect 2878 2454 2884 2455
rect 3046 2459 3052 2460
rect 3046 2455 3047 2459
rect 3051 2455 3052 2459
rect 3046 2454 3052 2455
rect 3206 2459 3212 2460
rect 3206 2455 3207 2459
rect 3211 2455 3212 2459
rect 3206 2454 3212 2455
rect 3358 2459 3364 2460
rect 3358 2455 3359 2459
rect 3363 2455 3364 2459
rect 3358 2454 3364 2455
rect 3502 2459 3508 2460
rect 3502 2455 3503 2459
rect 3507 2455 3508 2459
rect 3502 2454 3508 2455
rect 3654 2459 3660 2460
rect 3654 2455 3655 2459
rect 3659 2455 3660 2459
rect 3654 2454 3660 2455
rect 3806 2459 3812 2460
rect 3806 2455 3807 2459
rect 3811 2455 3812 2459
rect 3942 2456 3943 2460
rect 3947 2456 3948 2460
rect 3942 2455 3948 2456
rect 3806 2454 3812 2455
rect 134 2445 140 2446
rect 110 2444 116 2445
rect 110 2440 111 2444
rect 115 2440 116 2444
rect 134 2441 135 2445
rect 139 2441 140 2445
rect 134 2440 140 2441
rect 230 2445 236 2446
rect 230 2441 231 2445
rect 235 2441 236 2445
rect 230 2440 236 2441
rect 326 2445 332 2446
rect 326 2441 327 2445
rect 331 2441 332 2445
rect 326 2440 332 2441
rect 422 2445 428 2446
rect 422 2441 423 2445
rect 427 2441 428 2445
rect 422 2440 428 2441
rect 518 2445 524 2446
rect 518 2441 519 2445
rect 523 2441 524 2445
rect 518 2440 524 2441
rect 2006 2444 2012 2445
rect 2006 2440 2007 2444
rect 2011 2440 2012 2444
rect 110 2439 116 2440
rect 112 2403 114 2439
rect 136 2403 138 2440
rect 232 2403 234 2440
rect 328 2403 330 2440
rect 424 2403 426 2440
rect 520 2403 522 2440
rect 2006 2439 2012 2440
rect 2046 2443 2052 2444
rect 2046 2439 2047 2443
rect 2051 2439 2052 2443
rect 3942 2443 3948 2444
rect 2008 2403 2010 2439
rect 2046 2438 2052 2439
rect 2534 2440 2540 2441
rect 111 2402 115 2403
rect 111 2397 115 2398
rect 135 2402 139 2403
rect 135 2397 139 2398
rect 231 2402 235 2403
rect 231 2397 235 2398
rect 255 2402 259 2403
rect 255 2397 259 2398
rect 327 2402 331 2403
rect 327 2397 331 2398
rect 415 2402 419 2403
rect 415 2397 419 2398
rect 423 2402 427 2403
rect 423 2397 427 2398
rect 519 2402 523 2403
rect 519 2397 523 2398
rect 575 2402 579 2403
rect 575 2397 579 2398
rect 735 2402 739 2403
rect 735 2397 739 2398
rect 887 2402 891 2403
rect 887 2397 891 2398
rect 1039 2402 1043 2403
rect 1039 2397 1043 2398
rect 1183 2402 1187 2403
rect 1183 2397 1187 2398
rect 1327 2402 1331 2403
rect 1327 2397 1331 2398
rect 1479 2402 1483 2403
rect 1479 2397 1483 2398
rect 2007 2402 2011 2403
rect 2048 2399 2050 2438
rect 2534 2436 2535 2440
rect 2539 2436 2540 2440
rect 2534 2435 2540 2436
rect 2710 2440 2716 2441
rect 2710 2436 2711 2440
rect 2715 2436 2716 2440
rect 2710 2435 2716 2436
rect 2878 2440 2884 2441
rect 2878 2436 2879 2440
rect 2883 2436 2884 2440
rect 2878 2435 2884 2436
rect 3046 2440 3052 2441
rect 3046 2436 3047 2440
rect 3051 2436 3052 2440
rect 3046 2435 3052 2436
rect 3206 2440 3212 2441
rect 3206 2436 3207 2440
rect 3211 2436 3212 2440
rect 3206 2435 3212 2436
rect 3358 2440 3364 2441
rect 3358 2436 3359 2440
rect 3363 2436 3364 2440
rect 3358 2435 3364 2436
rect 3502 2440 3508 2441
rect 3502 2436 3503 2440
rect 3507 2436 3508 2440
rect 3502 2435 3508 2436
rect 3654 2440 3660 2441
rect 3654 2436 3655 2440
rect 3659 2436 3660 2440
rect 3654 2435 3660 2436
rect 3806 2440 3812 2441
rect 3806 2436 3807 2440
rect 3811 2436 3812 2440
rect 3942 2439 3943 2443
rect 3947 2439 3948 2443
rect 3942 2438 3948 2439
rect 3806 2435 3812 2436
rect 2536 2399 2538 2435
rect 2712 2399 2714 2435
rect 2880 2399 2882 2435
rect 3048 2399 3050 2435
rect 3208 2399 3210 2435
rect 3360 2399 3362 2435
rect 3504 2399 3506 2435
rect 3656 2399 3658 2435
rect 3808 2399 3810 2435
rect 3944 2399 3946 2438
rect 2007 2397 2011 2398
rect 2047 2398 2051 2399
rect 112 2377 114 2397
rect 110 2376 116 2377
rect 136 2376 138 2397
rect 256 2376 258 2397
rect 416 2376 418 2397
rect 576 2376 578 2397
rect 736 2376 738 2397
rect 888 2376 890 2397
rect 1040 2376 1042 2397
rect 1184 2376 1186 2397
rect 1328 2376 1330 2397
rect 1480 2376 1482 2397
rect 2008 2377 2010 2397
rect 2047 2393 2051 2394
rect 2535 2398 2539 2399
rect 2535 2393 2539 2394
rect 2607 2398 2611 2399
rect 2607 2393 2611 2394
rect 2711 2398 2715 2399
rect 2711 2393 2715 2394
rect 2815 2398 2819 2399
rect 2815 2393 2819 2394
rect 2879 2398 2883 2399
rect 2879 2393 2883 2394
rect 3007 2398 3011 2399
rect 3007 2393 3011 2394
rect 3047 2398 3051 2399
rect 3047 2393 3051 2394
rect 3191 2398 3195 2399
rect 3191 2393 3195 2394
rect 3207 2398 3211 2399
rect 3207 2393 3211 2394
rect 3359 2398 3363 2399
rect 3359 2393 3363 2394
rect 3503 2398 3507 2399
rect 3503 2393 3507 2394
rect 3519 2398 3523 2399
rect 3519 2393 3523 2394
rect 3655 2398 3659 2399
rect 3655 2393 3659 2394
rect 3679 2398 3683 2399
rect 3679 2393 3683 2394
rect 3807 2398 3811 2399
rect 3807 2393 3811 2394
rect 3839 2398 3843 2399
rect 3839 2393 3843 2394
rect 3943 2398 3947 2399
rect 3943 2393 3947 2394
rect 2006 2376 2012 2377
rect 110 2372 111 2376
rect 115 2372 116 2376
rect 110 2371 116 2372
rect 134 2375 140 2376
rect 134 2371 135 2375
rect 139 2371 140 2375
rect 134 2370 140 2371
rect 254 2375 260 2376
rect 254 2371 255 2375
rect 259 2371 260 2375
rect 254 2370 260 2371
rect 414 2375 420 2376
rect 414 2371 415 2375
rect 419 2371 420 2375
rect 414 2370 420 2371
rect 574 2375 580 2376
rect 574 2371 575 2375
rect 579 2371 580 2375
rect 574 2370 580 2371
rect 734 2375 740 2376
rect 734 2371 735 2375
rect 739 2371 740 2375
rect 734 2370 740 2371
rect 886 2375 892 2376
rect 886 2371 887 2375
rect 891 2371 892 2375
rect 886 2370 892 2371
rect 1038 2375 1044 2376
rect 1038 2371 1039 2375
rect 1043 2371 1044 2375
rect 1038 2370 1044 2371
rect 1182 2375 1188 2376
rect 1182 2371 1183 2375
rect 1187 2371 1188 2375
rect 1182 2370 1188 2371
rect 1326 2375 1332 2376
rect 1326 2371 1327 2375
rect 1331 2371 1332 2375
rect 1326 2370 1332 2371
rect 1478 2375 1484 2376
rect 1478 2371 1479 2375
rect 1483 2371 1484 2375
rect 2006 2372 2007 2376
rect 2011 2372 2012 2376
rect 2006 2371 2012 2372
rect 1478 2370 1484 2371
rect 2048 2366 2050 2393
rect 2608 2369 2610 2393
rect 2816 2369 2818 2393
rect 3008 2369 3010 2393
rect 3192 2369 3194 2393
rect 3360 2369 3362 2393
rect 3520 2369 3522 2393
rect 3680 2369 3682 2393
rect 3840 2369 3842 2393
rect 2606 2368 2612 2369
rect 2046 2365 2052 2366
rect 2046 2361 2047 2365
rect 2051 2361 2052 2365
rect 2606 2364 2607 2368
rect 2611 2364 2612 2368
rect 2606 2363 2612 2364
rect 2814 2368 2820 2369
rect 2814 2364 2815 2368
rect 2819 2364 2820 2368
rect 2814 2363 2820 2364
rect 3006 2368 3012 2369
rect 3006 2364 3007 2368
rect 3011 2364 3012 2368
rect 3006 2363 3012 2364
rect 3190 2368 3196 2369
rect 3190 2364 3191 2368
rect 3195 2364 3196 2368
rect 3190 2363 3196 2364
rect 3358 2368 3364 2369
rect 3358 2364 3359 2368
rect 3363 2364 3364 2368
rect 3358 2363 3364 2364
rect 3518 2368 3524 2369
rect 3518 2364 3519 2368
rect 3523 2364 3524 2368
rect 3518 2363 3524 2364
rect 3678 2368 3684 2369
rect 3678 2364 3679 2368
rect 3683 2364 3684 2368
rect 3678 2363 3684 2364
rect 3838 2368 3844 2369
rect 3838 2364 3839 2368
rect 3843 2364 3844 2368
rect 3944 2366 3946 2393
rect 3838 2363 3844 2364
rect 3942 2365 3948 2366
rect 2046 2360 2052 2361
rect 3942 2361 3943 2365
rect 3947 2361 3948 2365
rect 3942 2360 3948 2361
rect 110 2359 116 2360
rect 110 2355 111 2359
rect 115 2355 116 2359
rect 2006 2359 2012 2360
rect 110 2354 116 2355
rect 134 2356 140 2357
rect 112 2327 114 2354
rect 134 2352 135 2356
rect 139 2352 140 2356
rect 134 2351 140 2352
rect 254 2356 260 2357
rect 254 2352 255 2356
rect 259 2352 260 2356
rect 254 2351 260 2352
rect 414 2356 420 2357
rect 414 2352 415 2356
rect 419 2352 420 2356
rect 414 2351 420 2352
rect 574 2356 580 2357
rect 574 2352 575 2356
rect 579 2352 580 2356
rect 574 2351 580 2352
rect 734 2356 740 2357
rect 734 2352 735 2356
rect 739 2352 740 2356
rect 734 2351 740 2352
rect 886 2356 892 2357
rect 886 2352 887 2356
rect 891 2352 892 2356
rect 886 2351 892 2352
rect 1038 2356 1044 2357
rect 1038 2352 1039 2356
rect 1043 2352 1044 2356
rect 1038 2351 1044 2352
rect 1182 2356 1188 2357
rect 1182 2352 1183 2356
rect 1187 2352 1188 2356
rect 1182 2351 1188 2352
rect 1326 2356 1332 2357
rect 1326 2352 1327 2356
rect 1331 2352 1332 2356
rect 1326 2351 1332 2352
rect 1478 2356 1484 2357
rect 1478 2352 1479 2356
rect 1483 2352 1484 2356
rect 2006 2355 2007 2359
rect 2011 2355 2012 2359
rect 2006 2354 2012 2355
rect 1478 2351 1484 2352
rect 136 2327 138 2351
rect 256 2327 258 2351
rect 416 2327 418 2351
rect 576 2327 578 2351
rect 736 2327 738 2351
rect 888 2327 890 2351
rect 1040 2327 1042 2351
rect 1184 2327 1186 2351
rect 1328 2327 1330 2351
rect 1480 2327 1482 2351
rect 2008 2327 2010 2354
rect 2606 2349 2612 2350
rect 2046 2348 2052 2349
rect 2046 2344 2047 2348
rect 2051 2344 2052 2348
rect 2606 2345 2607 2349
rect 2611 2345 2612 2349
rect 2606 2344 2612 2345
rect 2814 2349 2820 2350
rect 2814 2345 2815 2349
rect 2819 2345 2820 2349
rect 2814 2344 2820 2345
rect 3006 2349 3012 2350
rect 3006 2345 3007 2349
rect 3011 2345 3012 2349
rect 3006 2344 3012 2345
rect 3190 2349 3196 2350
rect 3190 2345 3191 2349
rect 3195 2345 3196 2349
rect 3190 2344 3196 2345
rect 3358 2349 3364 2350
rect 3358 2345 3359 2349
rect 3363 2345 3364 2349
rect 3358 2344 3364 2345
rect 3518 2349 3524 2350
rect 3518 2345 3519 2349
rect 3523 2345 3524 2349
rect 3518 2344 3524 2345
rect 3678 2349 3684 2350
rect 3678 2345 3679 2349
rect 3683 2345 3684 2349
rect 3678 2344 3684 2345
rect 3838 2349 3844 2350
rect 3838 2345 3839 2349
rect 3843 2345 3844 2349
rect 3838 2344 3844 2345
rect 3942 2348 3948 2349
rect 3942 2344 3943 2348
rect 3947 2344 3948 2348
rect 2046 2343 2052 2344
rect 111 2326 115 2327
rect 111 2321 115 2322
rect 135 2326 139 2327
rect 135 2321 139 2322
rect 255 2326 259 2327
rect 255 2321 259 2322
rect 263 2326 267 2327
rect 263 2321 267 2322
rect 415 2326 419 2327
rect 415 2321 419 2322
rect 423 2326 427 2327
rect 423 2321 427 2322
rect 575 2326 579 2327
rect 575 2321 579 2322
rect 583 2326 587 2327
rect 583 2321 587 2322
rect 735 2326 739 2327
rect 735 2321 739 2322
rect 743 2326 747 2327
rect 743 2321 747 2322
rect 887 2326 891 2327
rect 887 2321 891 2322
rect 895 2326 899 2327
rect 895 2321 899 2322
rect 1039 2326 1043 2327
rect 1039 2321 1043 2322
rect 1047 2326 1051 2327
rect 1047 2321 1051 2322
rect 1183 2326 1187 2327
rect 1183 2321 1187 2322
rect 1199 2326 1203 2327
rect 1199 2321 1203 2322
rect 1327 2326 1331 2327
rect 1327 2321 1331 2322
rect 1351 2326 1355 2327
rect 1351 2321 1355 2322
rect 1479 2326 1483 2327
rect 1479 2321 1483 2322
rect 1503 2326 1507 2327
rect 1503 2321 1507 2322
rect 2007 2326 2011 2327
rect 2007 2321 2011 2322
rect 112 2294 114 2321
rect 136 2297 138 2321
rect 264 2297 266 2321
rect 424 2297 426 2321
rect 584 2297 586 2321
rect 744 2297 746 2321
rect 896 2297 898 2321
rect 1048 2297 1050 2321
rect 1200 2297 1202 2321
rect 1352 2297 1354 2321
rect 1504 2297 1506 2321
rect 134 2296 140 2297
rect 110 2293 116 2294
rect 110 2289 111 2293
rect 115 2289 116 2293
rect 134 2292 135 2296
rect 139 2292 140 2296
rect 134 2291 140 2292
rect 262 2296 268 2297
rect 262 2292 263 2296
rect 267 2292 268 2296
rect 262 2291 268 2292
rect 422 2296 428 2297
rect 422 2292 423 2296
rect 427 2292 428 2296
rect 422 2291 428 2292
rect 582 2296 588 2297
rect 582 2292 583 2296
rect 587 2292 588 2296
rect 582 2291 588 2292
rect 742 2296 748 2297
rect 742 2292 743 2296
rect 747 2292 748 2296
rect 742 2291 748 2292
rect 894 2296 900 2297
rect 894 2292 895 2296
rect 899 2292 900 2296
rect 894 2291 900 2292
rect 1046 2296 1052 2297
rect 1046 2292 1047 2296
rect 1051 2292 1052 2296
rect 1046 2291 1052 2292
rect 1198 2296 1204 2297
rect 1198 2292 1199 2296
rect 1203 2292 1204 2296
rect 1198 2291 1204 2292
rect 1350 2296 1356 2297
rect 1350 2292 1351 2296
rect 1355 2292 1356 2296
rect 1350 2291 1356 2292
rect 1502 2296 1508 2297
rect 1502 2292 1503 2296
rect 1507 2292 1508 2296
rect 2008 2294 2010 2321
rect 2048 2307 2050 2343
rect 2608 2307 2610 2344
rect 2816 2307 2818 2344
rect 3008 2307 3010 2344
rect 3192 2307 3194 2344
rect 3360 2307 3362 2344
rect 3520 2307 3522 2344
rect 3680 2307 3682 2344
rect 3840 2307 3842 2344
rect 3942 2343 3948 2344
rect 3944 2307 3946 2343
rect 2047 2306 2051 2307
rect 2047 2301 2051 2302
rect 2071 2306 2075 2307
rect 2071 2301 2075 2302
rect 2167 2306 2171 2307
rect 2167 2301 2171 2302
rect 2271 2306 2275 2307
rect 2271 2301 2275 2302
rect 2415 2306 2419 2307
rect 2415 2301 2419 2302
rect 2575 2306 2579 2307
rect 2575 2301 2579 2302
rect 2607 2306 2611 2307
rect 2607 2301 2611 2302
rect 2743 2306 2747 2307
rect 2743 2301 2747 2302
rect 2815 2306 2819 2307
rect 2815 2301 2819 2302
rect 2911 2306 2915 2307
rect 2911 2301 2915 2302
rect 3007 2306 3011 2307
rect 3007 2301 3011 2302
rect 3071 2306 3075 2307
rect 3071 2301 3075 2302
rect 3191 2306 3195 2307
rect 3191 2301 3195 2302
rect 3231 2306 3235 2307
rect 3231 2301 3235 2302
rect 3359 2306 3363 2307
rect 3359 2301 3363 2302
rect 3383 2306 3387 2307
rect 3383 2301 3387 2302
rect 3519 2306 3523 2307
rect 3519 2301 3523 2302
rect 3535 2306 3539 2307
rect 3535 2301 3539 2302
rect 3679 2306 3683 2307
rect 3679 2301 3683 2302
rect 3695 2306 3699 2307
rect 3695 2301 3699 2302
rect 3839 2306 3843 2307
rect 3839 2301 3843 2302
rect 3943 2306 3947 2307
rect 3943 2301 3947 2302
rect 1502 2291 1508 2292
rect 2006 2293 2012 2294
rect 110 2288 116 2289
rect 2006 2289 2007 2293
rect 2011 2289 2012 2293
rect 2006 2288 2012 2289
rect 2048 2281 2050 2301
rect 2046 2280 2052 2281
rect 2072 2280 2074 2301
rect 2168 2280 2170 2301
rect 2272 2280 2274 2301
rect 2416 2280 2418 2301
rect 2576 2280 2578 2301
rect 2744 2280 2746 2301
rect 2912 2280 2914 2301
rect 3072 2280 3074 2301
rect 3232 2280 3234 2301
rect 3384 2280 3386 2301
rect 3536 2280 3538 2301
rect 3696 2280 3698 2301
rect 3944 2281 3946 2301
rect 3942 2280 3948 2281
rect 134 2277 140 2278
rect 110 2276 116 2277
rect 110 2272 111 2276
rect 115 2272 116 2276
rect 134 2273 135 2277
rect 139 2273 140 2277
rect 134 2272 140 2273
rect 262 2277 268 2278
rect 262 2273 263 2277
rect 267 2273 268 2277
rect 262 2272 268 2273
rect 422 2277 428 2278
rect 422 2273 423 2277
rect 427 2273 428 2277
rect 422 2272 428 2273
rect 582 2277 588 2278
rect 582 2273 583 2277
rect 587 2273 588 2277
rect 582 2272 588 2273
rect 742 2277 748 2278
rect 742 2273 743 2277
rect 747 2273 748 2277
rect 742 2272 748 2273
rect 894 2277 900 2278
rect 894 2273 895 2277
rect 899 2273 900 2277
rect 894 2272 900 2273
rect 1046 2277 1052 2278
rect 1046 2273 1047 2277
rect 1051 2273 1052 2277
rect 1046 2272 1052 2273
rect 1198 2277 1204 2278
rect 1198 2273 1199 2277
rect 1203 2273 1204 2277
rect 1198 2272 1204 2273
rect 1350 2277 1356 2278
rect 1350 2273 1351 2277
rect 1355 2273 1356 2277
rect 1350 2272 1356 2273
rect 1502 2277 1508 2278
rect 1502 2273 1503 2277
rect 1507 2273 1508 2277
rect 1502 2272 1508 2273
rect 2006 2276 2012 2277
rect 2006 2272 2007 2276
rect 2011 2272 2012 2276
rect 2046 2276 2047 2280
rect 2051 2276 2052 2280
rect 2046 2275 2052 2276
rect 2070 2279 2076 2280
rect 2070 2275 2071 2279
rect 2075 2275 2076 2279
rect 2070 2274 2076 2275
rect 2166 2279 2172 2280
rect 2166 2275 2167 2279
rect 2171 2275 2172 2279
rect 2166 2274 2172 2275
rect 2270 2279 2276 2280
rect 2270 2275 2271 2279
rect 2275 2275 2276 2279
rect 2270 2274 2276 2275
rect 2414 2279 2420 2280
rect 2414 2275 2415 2279
rect 2419 2275 2420 2279
rect 2414 2274 2420 2275
rect 2574 2279 2580 2280
rect 2574 2275 2575 2279
rect 2579 2275 2580 2279
rect 2574 2274 2580 2275
rect 2742 2279 2748 2280
rect 2742 2275 2743 2279
rect 2747 2275 2748 2279
rect 2742 2274 2748 2275
rect 2910 2279 2916 2280
rect 2910 2275 2911 2279
rect 2915 2275 2916 2279
rect 2910 2274 2916 2275
rect 3070 2279 3076 2280
rect 3070 2275 3071 2279
rect 3075 2275 3076 2279
rect 3070 2274 3076 2275
rect 3230 2279 3236 2280
rect 3230 2275 3231 2279
rect 3235 2275 3236 2279
rect 3230 2274 3236 2275
rect 3382 2279 3388 2280
rect 3382 2275 3383 2279
rect 3387 2275 3388 2279
rect 3382 2274 3388 2275
rect 3534 2279 3540 2280
rect 3534 2275 3535 2279
rect 3539 2275 3540 2279
rect 3534 2274 3540 2275
rect 3694 2279 3700 2280
rect 3694 2275 3695 2279
rect 3699 2275 3700 2279
rect 3942 2276 3943 2280
rect 3947 2276 3948 2280
rect 3942 2275 3948 2276
rect 3694 2274 3700 2275
rect 110 2271 116 2272
rect 112 2247 114 2271
rect 136 2247 138 2272
rect 264 2247 266 2272
rect 424 2247 426 2272
rect 584 2247 586 2272
rect 744 2247 746 2272
rect 896 2247 898 2272
rect 1048 2247 1050 2272
rect 1200 2247 1202 2272
rect 1352 2247 1354 2272
rect 1504 2247 1506 2272
rect 2006 2271 2012 2272
rect 2008 2247 2010 2271
rect 2046 2263 2052 2264
rect 2046 2259 2047 2263
rect 2051 2259 2052 2263
rect 3942 2263 3948 2264
rect 2046 2258 2052 2259
rect 2070 2260 2076 2261
rect 111 2246 115 2247
rect 111 2241 115 2242
rect 135 2246 139 2247
rect 135 2241 139 2242
rect 223 2246 227 2247
rect 223 2241 227 2242
rect 263 2246 267 2247
rect 263 2241 267 2242
rect 351 2246 355 2247
rect 351 2241 355 2242
rect 423 2246 427 2247
rect 423 2241 427 2242
rect 495 2246 499 2247
rect 495 2241 499 2242
rect 583 2246 587 2247
rect 583 2241 587 2242
rect 647 2246 651 2247
rect 647 2241 651 2242
rect 743 2246 747 2247
rect 743 2241 747 2242
rect 799 2246 803 2247
rect 799 2241 803 2242
rect 895 2246 899 2247
rect 895 2241 899 2242
rect 959 2246 963 2247
rect 959 2241 963 2242
rect 1047 2246 1051 2247
rect 1047 2241 1051 2242
rect 1119 2246 1123 2247
rect 1119 2241 1123 2242
rect 1199 2246 1203 2247
rect 1199 2241 1203 2242
rect 1279 2246 1283 2247
rect 1279 2241 1283 2242
rect 1351 2246 1355 2247
rect 1351 2241 1355 2242
rect 1439 2246 1443 2247
rect 1439 2241 1443 2242
rect 1503 2246 1507 2247
rect 1503 2241 1507 2242
rect 1599 2246 1603 2247
rect 1599 2241 1603 2242
rect 2007 2246 2011 2247
rect 2007 2241 2011 2242
rect 112 2221 114 2241
rect 110 2220 116 2221
rect 224 2220 226 2241
rect 352 2220 354 2241
rect 496 2220 498 2241
rect 648 2220 650 2241
rect 800 2220 802 2241
rect 960 2220 962 2241
rect 1120 2220 1122 2241
rect 1280 2220 1282 2241
rect 1440 2220 1442 2241
rect 1600 2220 1602 2241
rect 2008 2221 2010 2241
rect 2048 2231 2050 2258
rect 2070 2256 2071 2260
rect 2075 2256 2076 2260
rect 2070 2255 2076 2256
rect 2166 2260 2172 2261
rect 2166 2256 2167 2260
rect 2171 2256 2172 2260
rect 2166 2255 2172 2256
rect 2270 2260 2276 2261
rect 2270 2256 2271 2260
rect 2275 2256 2276 2260
rect 2270 2255 2276 2256
rect 2414 2260 2420 2261
rect 2414 2256 2415 2260
rect 2419 2256 2420 2260
rect 2414 2255 2420 2256
rect 2574 2260 2580 2261
rect 2574 2256 2575 2260
rect 2579 2256 2580 2260
rect 2574 2255 2580 2256
rect 2742 2260 2748 2261
rect 2742 2256 2743 2260
rect 2747 2256 2748 2260
rect 2742 2255 2748 2256
rect 2910 2260 2916 2261
rect 2910 2256 2911 2260
rect 2915 2256 2916 2260
rect 2910 2255 2916 2256
rect 3070 2260 3076 2261
rect 3070 2256 3071 2260
rect 3075 2256 3076 2260
rect 3070 2255 3076 2256
rect 3230 2260 3236 2261
rect 3230 2256 3231 2260
rect 3235 2256 3236 2260
rect 3230 2255 3236 2256
rect 3382 2260 3388 2261
rect 3382 2256 3383 2260
rect 3387 2256 3388 2260
rect 3382 2255 3388 2256
rect 3534 2260 3540 2261
rect 3534 2256 3535 2260
rect 3539 2256 3540 2260
rect 3534 2255 3540 2256
rect 3694 2260 3700 2261
rect 3694 2256 3695 2260
rect 3699 2256 3700 2260
rect 3942 2259 3943 2263
rect 3947 2259 3948 2263
rect 3942 2258 3948 2259
rect 3694 2255 3700 2256
rect 2072 2231 2074 2255
rect 2168 2231 2170 2255
rect 2272 2231 2274 2255
rect 2416 2231 2418 2255
rect 2576 2231 2578 2255
rect 2744 2231 2746 2255
rect 2912 2231 2914 2255
rect 3072 2231 3074 2255
rect 3232 2231 3234 2255
rect 3384 2231 3386 2255
rect 3536 2231 3538 2255
rect 3696 2231 3698 2255
rect 3944 2231 3946 2258
rect 2047 2230 2051 2231
rect 2047 2225 2051 2226
rect 2071 2230 2075 2231
rect 2071 2225 2075 2226
rect 2167 2230 2171 2231
rect 2167 2225 2171 2226
rect 2175 2230 2179 2231
rect 2175 2225 2179 2226
rect 2271 2230 2275 2231
rect 2271 2225 2275 2226
rect 2319 2230 2323 2231
rect 2319 2225 2323 2226
rect 2415 2230 2419 2231
rect 2415 2225 2419 2226
rect 2471 2230 2475 2231
rect 2471 2225 2475 2226
rect 2575 2230 2579 2231
rect 2575 2225 2579 2226
rect 2623 2230 2627 2231
rect 2623 2225 2627 2226
rect 2743 2230 2747 2231
rect 2743 2225 2747 2226
rect 2783 2230 2787 2231
rect 2783 2225 2787 2226
rect 2911 2230 2915 2231
rect 2911 2225 2915 2226
rect 2935 2230 2939 2231
rect 2935 2225 2939 2226
rect 3071 2230 3075 2231
rect 3071 2225 3075 2226
rect 3079 2230 3083 2231
rect 3079 2225 3083 2226
rect 3223 2230 3227 2231
rect 3223 2225 3227 2226
rect 3231 2230 3235 2231
rect 3231 2225 3235 2226
rect 3367 2230 3371 2231
rect 3367 2225 3371 2226
rect 3383 2230 3387 2231
rect 3383 2225 3387 2226
rect 3519 2230 3523 2231
rect 3519 2225 3523 2226
rect 3535 2230 3539 2231
rect 3535 2225 3539 2226
rect 3695 2230 3699 2231
rect 3695 2225 3699 2226
rect 3943 2230 3947 2231
rect 3943 2225 3947 2226
rect 2006 2220 2012 2221
rect 110 2216 111 2220
rect 115 2216 116 2220
rect 110 2215 116 2216
rect 222 2219 228 2220
rect 222 2215 223 2219
rect 227 2215 228 2219
rect 222 2214 228 2215
rect 350 2219 356 2220
rect 350 2215 351 2219
rect 355 2215 356 2219
rect 350 2214 356 2215
rect 494 2219 500 2220
rect 494 2215 495 2219
rect 499 2215 500 2219
rect 494 2214 500 2215
rect 646 2219 652 2220
rect 646 2215 647 2219
rect 651 2215 652 2219
rect 646 2214 652 2215
rect 798 2219 804 2220
rect 798 2215 799 2219
rect 803 2215 804 2219
rect 798 2214 804 2215
rect 958 2219 964 2220
rect 958 2215 959 2219
rect 963 2215 964 2219
rect 958 2214 964 2215
rect 1118 2219 1124 2220
rect 1118 2215 1119 2219
rect 1123 2215 1124 2219
rect 1118 2214 1124 2215
rect 1278 2219 1284 2220
rect 1278 2215 1279 2219
rect 1283 2215 1284 2219
rect 1278 2214 1284 2215
rect 1438 2219 1444 2220
rect 1438 2215 1439 2219
rect 1443 2215 1444 2219
rect 1438 2214 1444 2215
rect 1598 2219 1604 2220
rect 1598 2215 1599 2219
rect 1603 2215 1604 2219
rect 2006 2216 2007 2220
rect 2011 2216 2012 2220
rect 2006 2215 2012 2216
rect 1598 2214 1604 2215
rect 110 2203 116 2204
rect 110 2199 111 2203
rect 115 2199 116 2203
rect 2006 2203 2012 2204
rect 110 2198 116 2199
rect 222 2200 228 2201
rect 112 2171 114 2198
rect 222 2196 223 2200
rect 227 2196 228 2200
rect 222 2195 228 2196
rect 350 2200 356 2201
rect 350 2196 351 2200
rect 355 2196 356 2200
rect 350 2195 356 2196
rect 494 2200 500 2201
rect 494 2196 495 2200
rect 499 2196 500 2200
rect 494 2195 500 2196
rect 646 2200 652 2201
rect 646 2196 647 2200
rect 651 2196 652 2200
rect 646 2195 652 2196
rect 798 2200 804 2201
rect 798 2196 799 2200
rect 803 2196 804 2200
rect 798 2195 804 2196
rect 958 2200 964 2201
rect 958 2196 959 2200
rect 963 2196 964 2200
rect 958 2195 964 2196
rect 1118 2200 1124 2201
rect 1118 2196 1119 2200
rect 1123 2196 1124 2200
rect 1118 2195 1124 2196
rect 1278 2200 1284 2201
rect 1278 2196 1279 2200
rect 1283 2196 1284 2200
rect 1278 2195 1284 2196
rect 1438 2200 1444 2201
rect 1438 2196 1439 2200
rect 1443 2196 1444 2200
rect 1438 2195 1444 2196
rect 1598 2200 1604 2201
rect 1598 2196 1599 2200
rect 1603 2196 1604 2200
rect 2006 2199 2007 2203
rect 2011 2199 2012 2203
rect 2006 2198 2012 2199
rect 2048 2198 2050 2225
rect 2072 2201 2074 2225
rect 2176 2201 2178 2225
rect 2320 2201 2322 2225
rect 2472 2201 2474 2225
rect 2624 2201 2626 2225
rect 2784 2201 2786 2225
rect 2936 2201 2938 2225
rect 3080 2201 3082 2225
rect 3224 2201 3226 2225
rect 3368 2201 3370 2225
rect 3520 2201 3522 2225
rect 2070 2200 2076 2201
rect 1598 2195 1604 2196
rect 224 2171 226 2195
rect 352 2171 354 2195
rect 496 2171 498 2195
rect 648 2171 650 2195
rect 800 2171 802 2195
rect 960 2171 962 2195
rect 1120 2171 1122 2195
rect 1280 2171 1282 2195
rect 1440 2171 1442 2195
rect 1600 2171 1602 2195
rect 2008 2171 2010 2198
rect 2046 2197 2052 2198
rect 2046 2193 2047 2197
rect 2051 2193 2052 2197
rect 2070 2196 2071 2200
rect 2075 2196 2076 2200
rect 2070 2195 2076 2196
rect 2174 2200 2180 2201
rect 2174 2196 2175 2200
rect 2179 2196 2180 2200
rect 2174 2195 2180 2196
rect 2318 2200 2324 2201
rect 2318 2196 2319 2200
rect 2323 2196 2324 2200
rect 2318 2195 2324 2196
rect 2470 2200 2476 2201
rect 2470 2196 2471 2200
rect 2475 2196 2476 2200
rect 2470 2195 2476 2196
rect 2622 2200 2628 2201
rect 2622 2196 2623 2200
rect 2627 2196 2628 2200
rect 2622 2195 2628 2196
rect 2782 2200 2788 2201
rect 2782 2196 2783 2200
rect 2787 2196 2788 2200
rect 2782 2195 2788 2196
rect 2934 2200 2940 2201
rect 2934 2196 2935 2200
rect 2939 2196 2940 2200
rect 2934 2195 2940 2196
rect 3078 2200 3084 2201
rect 3078 2196 3079 2200
rect 3083 2196 3084 2200
rect 3078 2195 3084 2196
rect 3222 2200 3228 2201
rect 3222 2196 3223 2200
rect 3227 2196 3228 2200
rect 3222 2195 3228 2196
rect 3366 2200 3372 2201
rect 3366 2196 3367 2200
rect 3371 2196 3372 2200
rect 3366 2195 3372 2196
rect 3518 2200 3524 2201
rect 3518 2196 3519 2200
rect 3523 2196 3524 2200
rect 3944 2198 3946 2225
rect 3518 2195 3524 2196
rect 3942 2197 3948 2198
rect 2046 2192 2052 2193
rect 3942 2193 3943 2197
rect 3947 2193 3948 2197
rect 3942 2192 3948 2193
rect 2070 2181 2076 2182
rect 2046 2180 2052 2181
rect 2046 2176 2047 2180
rect 2051 2176 2052 2180
rect 2070 2177 2071 2181
rect 2075 2177 2076 2181
rect 2070 2176 2076 2177
rect 2174 2181 2180 2182
rect 2174 2177 2175 2181
rect 2179 2177 2180 2181
rect 2174 2176 2180 2177
rect 2318 2181 2324 2182
rect 2318 2177 2319 2181
rect 2323 2177 2324 2181
rect 2318 2176 2324 2177
rect 2470 2181 2476 2182
rect 2470 2177 2471 2181
rect 2475 2177 2476 2181
rect 2470 2176 2476 2177
rect 2622 2181 2628 2182
rect 2622 2177 2623 2181
rect 2627 2177 2628 2181
rect 2622 2176 2628 2177
rect 2782 2181 2788 2182
rect 2782 2177 2783 2181
rect 2787 2177 2788 2181
rect 2782 2176 2788 2177
rect 2934 2181 2940 2182
rect 2934 2177 2935 2181
rect 2939 2177 2940 2181
rect 2934 2176 2940 2177
rect 3078 2181 3084 2182
rect 3078 2177 3079 2181
rect 3083 2177 3084 2181
rect 3078 2176 3084 2177
rect 3222 2181 3228 2182
rect 3222 2177 3223 2181
rect 3227 2177 3228 2181
rect 3222 2176 3228 2177
rect 3366 2181 3372 2182
rect 3366 2177 3367 2181
rect 3371 2177 3372 2181
rect 3366 2176 3372 2177
rect 3518 2181 3524 2182
rect 3518 2177 3519 2181
rect 3523 2177 3524 2181
rect 3518 2176 3524 2177
rect 3942 2180 3948 2181
rect 3942 2176 3943 2180
rect 3947 2176 3948 2180
rect 2046 2175 2052 2176
rect 111 2170 115 2171
rect 111 2165 115 2166
rect 223 2170 227 2171
rect 223 2165 227 2166
rect 351 2170 355 2171
rect 351 2165 355 2166
rect 471 2170 475 2171
rect 471 2165 475 2166
rect 495 2170 499 2171
rect 495 2165 499 2166
rect 567 2170 571 2171
rect 567 2165 571 2166
rect 647 2170 651 2171
rect 647 2165 651 2166
rect 679 2170 683 2171
rect 679 2165 683 2166
rect 799 2170 803 2171
rect 799 2165 803 2166
rect 807 2170 811 2171
rect 807 2165 811 2166
rect 943 2170 947 2171
rect 943 2165 947 2166
rect 959 2170 963 2171
rect 959 2165 963 2166
rect 1079 2170 1083 2171
rect 1079 2165 1083 2166
rect 1119 2170 1123 2171
rect 1119 2165 1123 2166
rect 1223 2170 1227 2171
rect 1223 2165 1227 2166
rect 1279 2170 1283 2171
rect 1279 2165 1283 2166
rect 1367 2170 1371 2171
rect 1367 2165 1371 2166
rect 1439 2170 1443 2171
rect 1439 2165 1443 2166
rect 1503 2170 1507 2171
rect 1503 2165 1507 2166
rect 1599 2170 1603 2171
rect 1599 2165 1603 2166
rect 1639 2170 1643 2171
rect 1639 2165 1643 2166
rect 1783 2170 1787 2171
rect 1783 2165 1787 2166
rect 1903 2170 1907 2171
rect 1903 2165 1907 2166
rect 2007 2170 2011 2171
rect 2007 2165 2011 2166
rect 112 2138 114 2165
rect 472 2141 474 2165
rect 568 2141 570 2165
rect 680 2141 682 2165
rect 808 2141 810 2165
rect 944 2141 946 2165
rect 1080 2141 1082 2165
rect 1224 2141 1226 2165
rect 1368 2141 1370 2165
rect 1504 2141 1506 2165
rect 1640 2141 1642 2165
rect 1784 2141 1786 2165
rect 1904 2141 1906 2165
rect 470 2140 476 2141
rect 110 2137 116 2138
rect 110 2133 111 2137
rect 115 2133 116 2137
rect 470 2136 471 2140
rect 475 2136 476 2140
rect 470 2135 476 2136
rect 566 2140 572 2141
rect 566 2136 567 2140
rect 571 2136 572 2140
rect 566 2135 572 2136
rect 678 2140 684 2141
rect 678 2136 679 2140
rect 683 2136 684 2140
rect 678 2135 684 2136
rect 806 2140 812 2141
rect 806 2136 807 2140
rect 811 2136 812 2140
rect 806 2135 812 2136
rect 942 2140 948 2141
rect 942 2136 943 2140
rect 947 2136 948 2140
rect 942 2135 948 2136
rect 1078 2140 1084 2141
rect 1078 2136 1079 2140
rect 1083 2136 1084 2140
rect 1078 2135 1084 2136
rect 1222 2140 1228 2141
rect 1222 2136 1223 2140
rect 1227 2136 1228 2140
rect 1222 2135 1228 2136
rect 1366 2140 1372 2141
rect 1366 2136 1367 2140
rect 1371 2136 1372 2140
rect 1366 2135 1372 2136
rect 1502 2140 1508 2141
rect 1502 2136 1503 2140
rect 1507 2136 1508 2140
rect 1502 2135 1508 2136
rect 1638 2140 1644 2141
rect 1638 2136 1639 2140
rect 1643 2136 1644 2140
rect 1638 2135 1644 2136
rect 1782 2140 1788 2141
rect 1782 2136 1783 2140
rect 1787 2136 1788 2140
rect 1782 2135 1788 2136
rect 1902 2140 1908 2141
rect 1902 2136 1903 2140
rect 1907 2136 1908 2140
rect 2008 2138 2010 2165
rect 1902 2135 1908 2136
rect 2006 2137 2012 2138
rect 110 2132 116 2133
rect 2006 2133 2007 2137
rect 2011 2133 2012 2137
rect 2048 2135 2050 2175
rect 2072 2135 2074 2176
rect 2176 2135 2178 2176
rect 2320 2135 2322 2176
rect 2472 2135 2474 2176
rect 2624 2135 2626 2176
rect 2784 2135 2786 2176
rect 2936 2135 2938 2176
rect 3080 2135 3082 2176
rect 3224 2135 3226 2176
rect 3368 2135 3370 2176
rect 3520 2135 3522 2176
rect 3942 2175 3948 2176
rect 3944 2135 3946 2175
rect 2006 2132 2012 2133
rect 2047 2134 2051 2135
rect 2047 2129 2051 2130
rect 2071 2134 2075 2135
rect 2071 2129 2075 2130
rect 2175 2134 2179 2135
rect 2175 2129 2179 2130
rect 2279 2134 2283 2135
rect 2279 2129 2283 2130
rect 2319 2134 2323 2135
rect 2319 2129 2323 2130
rect 2391 2134 2395 2135
rect 2391 2129 2395 2130
rect 2471 2134 2475 2135
rect 2471 2129 2475 2130
rect 2511 2134 2515 2135
rect 2511 2129 2515 2130
rect 2623 2134 2627 2135
rect 2623 2129 2627 2130
rect 2631 2134 2635 2135
rect 2631 2129 2635 2130
rect 2759 2134 2763 2135
rect 2759 2129 2763 2130
rect 2783 2134 2787 2135
rect 2783 2129 2787 2130
rect 2895 2134 2899 2135
rect 2895 2129 2899 2130
rect 2935 2134 2939 2135
rect 2935 2129 2939 2130
rect 3039 2134 3043 2135
rect 3039 2129 3043 2130
rect 3079 2134 3083 2135
rect 3079 2129 3083 2130
rect 3191 2134 3195 2135
rect 3191 2129 3195 2130
rect 3223 2134 3227 2135
rect 3223 2129 3227 2130
rect 3351 2134 3355 2135
rect 3351 2129 3355 2130
rect 3367 2134 3371 2135
rect 3367 2129 3371 2130
rect 3519 2134 3523 2135
rect 3519 2129 3523 2130
rect 3687 2134 3691 2135
rect 3687 2129 3691 2130
rect 3839 2134 3843 2135
rect 3839 2129 3843 2130
rect 3943 2134 3947 2135
rect 3943 2129 3947 2130
rect 470 2121 476 2122
rect 110 2120 116 2121
rect 110 2116 111 2120
rect 115 2116 116 2120
rect 470 2117 471 2121
rect 475 2117 476 2121
rect 470 2116 476 2117
rect 566 2121 572 2122
rect 566 2117 567 2121
rect 571 2117 572 2121
rect 566 2116 572 2117
rect 678 2121 684 2122
rect 678 2117 679 2121
rect 683 2117 684 2121
rect 678 2116 684 2117
rect 806 2121 812 2122
rect 806 2117 807 2121
rect 811 2117 812 2121
rect 806 2116 812 2117
rect 942 2121 948 2122
rect 942 2117 943 2121
rect 947 2117 948 2121
rect 942 2116 948 2117
rect 1078 2121 1084 2122
rect 1078 2117 1079 2121
rect 1083 2117 1084 2121
rect 1078 2116 1084 2117
rect 1222 2121 1228 2122
rect 1222 2117 1223 2121
rect 1227 2117 1228 2121
rect 1222 2116 1228 2117
rect 1366 2121 1372 2122
rect 1366 2117 1367 2121
rect 1371 2117 1372 2121
rect 1366 2116 1372 2117
rect 1502 2121 1508 2122
rect 1502 2117 1503 2121
rect 1507 2117 1508 2121
rect 1502 2116 1508 2117
rect 1638 2121 1644 2122
rect 1638 2117 1639 2121
rect 1643 2117 1644 2121
rect 1638 2116 1644 2117
rect 1782 2121 1788 2122
rect 1782 2117 1783 2121
rect 1787 2117 1788 2121
rect 1782 2116 1788 2117
rect 1902 2121 1908 2122
rect 1902 2117 1903 2121
rect 1907 2117 1908 2121
rect 1902 2116 1908 2117
rect 2006 2120 2012 2121
rect 2006 2116 2007 2120
rect 2011 2116 2012 2120
rect 110 2115 116 2116
rect 112 2095 114 2115
rect 472 2095 474 2116
rect 568 2095 570 2116
rect 680 2095 682 2116
rect 808 2095 810 2116
rect 944 2095 946 2116
rect 1080 2095 1082 2116
rect 1224 2095 1226 2116
rect 1368 2095 1370 2116
rect 1504 2095 1506 2116
rect 1640 2095 1642 2116
rect 1784 2095 1786 2116
rect 1904 2095 1906 2116
rect 2006 2115 2012 2116
rect 2008 2095 2010 2115
rect 2048 2109 2050 2129
rect 2046 2108 2052 2109
rect 2280 2108 2282 2129
rect 2392 2108 2394 2129
rect 2512 2108 2514 2129
rect 2632 2108 2634 2129
rect 2760 2108 2762 2129
rect 2896 2108 2898 2129
rect 3040 2108 3042 2129
rect 3192 2108 3194 2129
rect 3352 2108 3354 2129
rect 3520 2108 3522 2129
rect 3688 2108 3690 2129
rect 3840 2108 3842 2129
rect 3944 2109 3946 2129
rect 3942 2108 3948 2109
rect 2046 2104 2047 2108
rect 2051 2104 2052 2108
rect 2046 2103 2052 2104
rect 2278 2107 2284 2108
rect 2278 2103 2279 2107
rect 2283 2103 2284 2107
rect 2278 2102 2284 2103
rect 2390 2107 2396 2108
rect 2390 2103 2391 2107
rect 2395 2103 2396 2107
rect 2390 2102 2396 2103
rect 2510 2107 2516 2108
rect 2510 2103 2511 2107
rect 2515 2103 2516 2107
rect 2510 2102 2516 2103
rect 2630 2107 2636 2108
rect 2630 2103 2631 2107
rect 2635 2103 2636 2107
rect 2630 2102 2636 2103
rect 2758 2107 2764 2108
rect 2758 2103 2759 2107
rect 2763 2103 2764 2107
rect 2758 2102 2764 2103
rect 2894 2107 2900 2108
rect 2894 2103 2895 2107
rect 2899 2103 2900 2107
rect 2894 2102 2900 2103
rect 3038 2107 3044 2108
rect 3038 2103 3039 2107
rect 3043 2103 3044 2107
rect 3038 2102 3044 2103
rect 3190 2107 3196 2108
rect 3190 2103 3191 2107
rect 3195 2103 3196 2107
rect 3190 2102 3196 2103
rect 3350 2107 3356 2108
rect 3350 2103 3351 2107
rect 3355 2103 3356 2107
rect 3350 2102 3356 2103
rect 3518 2107 3524 2108
rect 3518 2103 3519 2107
rect 3523 2103 3524 2107
rect 3518 2102 3524 2103
rect 3686 2107 3692 2108
rect 3686 2103 3687 2107
rect 3691 2103 3692 2107
rect 3686 2102 3692 2103
rect 3838 2107 3844 2108
rect 3838 2103 3839 2107
rect 3843 2103 3844 2107
rect 3942 2104 3943 2108
rect 3947 2104 3948 2108
rect 3942 2103 3948 2104
rect 3838 2102 3844 2103
rect 111 2094 115 2095
rect 111 2089 115 2090
rect 471 2094 475 2095
rect 471 2089 475 2090
rect 567 2094 571 2095
rect 567 2089 571 2090
rect 623 2094 627 2095
rect 623 2089 627 2090
rect 679 2094 683 2095
rect 679 2089 683 2090
rect 735 2094 739 2095
rect 735 2089 739 2090
rect 807 2094 811 2095
rect 807 2089 811 2090
rect 855 2094 859 2095
rect 855 2089 859 2090
rect 943 2094 947 2095
rect 943 2089 947 2090
rect 983 2094 987 2095
rect 983 2089 987 2090
rect 1079 2094 1083 2095
rect 1079 2089 1083 2090
rect 1119 2094 1123 2095
rect 1119 2089 1123 2090
rect 1223 2094 1227 2095
rect 1223 2089 1227 2090
rect 1255 2094 1259 2095
rect 1255 2089 1259 2090
rect 1367 2094 1371 2095
rect 1367 2089 1371 2090
rect 1391 2094 1395 2095
rect 1391 2089 1395 2090
rect 1503 2094 1507 2095
rect 1503 2089 1507 2090
rect 1527 2094 1531 2095
rect 1527 2089 1531 2090
rect 1639 2094 1643 2095
rect 1639 2089 1643 2090
rect 1655 2094 1659 2095
rect 1655 2089 1659 2090
rect 1783 2094 1787 2095
rect 1783 2089 1787 2090
rect 1791 2094 1795 2095
rect 1791 2089 1795 2090
rect 1903 2094 1907 2095
rect 1903 2089 1907 2090
rect 2007 2094 2011 2095
rect 2007 2089 2011 2090
rect 2046 2091 2052 2092
rect 112 2069 114 2089
rect 110 2068 116 2069
rect 624 2068 626 2089
rect 736 2068 738 2089
rect 856 2068 858 2089
rect 984 2068 986 2089
rect 1120 2068 1122 2089
rect 1256 2068 1258 2089
rect 1392 2068 1394 2089
rect 1528 2068 1530 2089
rect 1656 2068 1658 2089
rect 1792 2068 1794 2089
rect 1904 2068 1906 2089
rect 2008 2069 2010 2089
rect 2046 2087 2047 2091
rect 2051 2087 2052 2091
rect 3942 2091 3948 2092
rect 2046 2086 2052 2087
rect 2278 2088 2284 2089
rect 2006 2068 2012 2069
rect 110 2064 111 2068
rect 115 2064 116 2068
rect 110 2063 116 2064
rect 622 2067 628 2068
rect 622 2063 623 2067
rect 627 2063 628 2067
rect 622 2062 628 2063
rect 734 2067 740 2068
rect 734 2063 735 2067
rect 739 2063 740 2067
rect 734 2062 740 2063
rect 854 2067 860 2068
rect 854 2063 855 2067
rect 859 2063 860 2067
rect 854 2062 860 2063
rect 982 2067 988 2068
rect 982 2063 983 2067
rect 987 2063 988 2067
rect 982 2062 988 2063
rect 1118 2067 1124 2068
rect 1118 2063 1119 2067
rect 1123 2063 1124 2067
rect 1118 2062 1124 2063
rect 1254 2067 1260 2068
rect 1254 2063 1255 2067
rect 1259 2063 1260 2067
rect 1254 2062 1260 2063
rect 1390 2067 1396 2068
rect 1390 2063 1391 2067
rect 1395 2063 1396 2067
rect 1390 2062 1396 2063
rect 1526 2067 1532 2068
rect 1526 2063 1527 2067
rect 1531 2063 1532 2067
rect 1526 2062 1532 2063
rect 1654 2067 1660 2068
rect 1654 2063 1655 2067
rect 1659 2063 1660 2067
rect 1654 2062 1660 2063
rect 1790 2067 1796 2068
rect 1790 2063 1791 2067
rect 1795 2063 1796 2067
rect 1790 2062 1796 2063
rect 1902 2067 1908 2068
rect 1902 2063 1903 2067
rect 1907 2063 1908 2067
rect 2006 2064 2007 2068
rect 2011 2064 2012 2068
rect 2006 2063 2012 2064
rect 1902 2062 1908 2063
rect 110 2051 116 2052
rect 110 2047 111 2051
rect 115 2047 116 2051
rect 2006 2051 2012 2052
rect 2048 2051 2050 2086
rect 2278 2084 2279 2088
rect 2283 2084 2284 2088
rect 2278 2083 2284 2084
rect 2390 2088 2396 2089
rect 2390 2084 2391 2088
rect 2395 2084 2396 2088
rect 2390 2083 2396 2084
rect 2510 2088 2516 2089
rect 2510 2084 2511 2088
rect 2515 2084 2516 2088
rect 2510 2083 2516 2084
rect 2630 2088 2636 2089
rect 2630 2084 2631 2088
rect 2635 2084 2636 2088
rect 2630 2083 2636 2084
rect 2758 2088 2764 2089
rect 2758 2084 2759 2088
rect 2763 2084 2764 2088
rect 2758 2083 2764 2084
rect 2894 2088 2900 2089
rect 2894 2084 2895 2088
rect 2899 2084 2900 2088
rect 2894 2083 2900 2084
rect 3038 2088 3044 2089
rect 3038 2084 3039 2088
rect 3043 2084 3044 2088
rect 3038 2083 3044 2084
rect 3190 2088 3196 2089
rect 3190 2084 3191 2088
rect 3195 2084 3196 2088
rect 3190 2083 3196 2084
rect 3350 2088 3356 2089
rect 3350 2084 3351 2088
rect 3355 2084 3356 2088
rect 3350 2083 3356 2084
rect 3518 2088 3524 2089
rect 3518 2084 3519 2088
rect 3523 2084 3524 2088
rect 3518 2083 3524 2084
rect 3686 2088 3692 2089
rect 3686 2084 3687 2088
rect 3691 2084 3692 2088
rect 3686 2083 3692 2084
rect 3838 2088 3844 2089
rect 3838 2084 3839 2088
rect 3843 2084 3844 2088
rect 3942 2087 3943 2091
rect 3947 2087 3948 2091
rect 3942 2086 3948 2087
rect 3838 2083 3844 2084
rect 2280 2051 2282 2083
rect 2392 2051 2394 2083
rect 2512 2051 2514 2083
rect 2632 2051 2634 2083
rect 2760 2051 2762 2083
rect 2896 2051 2898 2083
rect 3040 2051 3042 2083
rect 3192 2051 3194 2083
rect 3352 2051 3354 2083
rect 3520 2051 3522 2083
rect 3688 2051 3690 2083
rect 3840 2051 3842 2083
rect 3944 2051 3946 2086
rect 110 2046 116 2047
rect 622 2048 628 2049
rect 112 2015 114 2046
rect 622 2044 623 2048
rect 627 2044 628 2048
rect 622 2043 628 2044
rect 734 2048 740 2049
rect 734 2044 735 2048
rect 739 2044 740 2048
rect 734 2043 740 2044
rect 854 2048 860 2049
rect 854 2044 855 2048
rect 859 2044 860 2048
rect 854 2043 860 2044
rect 982 2048 988 2049
rect 982 2044 983 2048
rect 987 2044 988 2048
rect 982 2043 988 2044
rect 1118 2048 1124 2049
rect 1118 2044 1119 2048
rect 1123 2044 1124 2048
rect 1118 2043 1124 2044
rect 1254 2048 1260 2049
rect 1254 2044 1255 2048
rect 1259 2044 1260 2048
rect 1254 2043 1260 2044
rect 1390 2048 1396 2049
rect 1390 2044 1391 2048
rect 1395 2044 1396 2048
rect 1390 2043 1396 2044
rect 1526 2048 1532 2049
rect 1526 2044 1527 2048
rect 1531 2044 1532 2048
rect 1526 2043 1532 2044
rect 1654 2048 1660 2049
rect 1654 2044 1655 2048
rect 1659 2044 1660 2048
rect 1654 2043 1660 2044
rect 1790 2048 1796 2049
rect 1790 2044 1791 2048
rect 1795 2044 1796 2048
rect 1790 2043 1796 2044
rect 1902 2048 1908 2049
rect 1902 2044 1903 2048
rect 1907 2044 1908 2048
rect 2006 2047 2007 2051
rect 2011 2047 2012 2051
rect 2006 2046 2012 2047
rect 2047 2050 2051 2051
rect 1902 2043 1908 2044
rect 624 2015 626 2043
rect 736 2015 738 2043
rect 856 2015 858 2043
rect 984 2015 986 2043
rect 1120 2015 1122 2043
rect 1256 2015 1258 2043
rect 1392 2015 1394 2043
rect 1528 2015 1530 2043
rect 1656 2015 1658 2043
rect 1792 2015 1794 2043
rect 1904 2015 1906 2043
rect 2008 2015 2010 2046
rect 2047 2045 2051 2046
rect 2279 2050 2283 2051
rect 2279 2045 2283 2046
rect 2327 2050 2331 2051
rect 2327 2045 2331 2046
rect 2391 2050 2395 2051
rect 2391 2045 2395 2046
rect 2431 2050 2435 2051
rect 2431 2045 2435 2046
rect 2511 2050 2515 2051
rect 2511 2045 2515 2046
rect 2535 2050 2539 2051
rect 2535 2045 2539 2046
rect 2631 2050 2635 2051
rect 2631 2045 2635 2046
rect 2647 2050 2651 2051
rect 2647 2045 2651 2046
rect 2759 2050 2763 2051
rect 2759 2045 2763 2046
rect 2775 2050 2779 2051
rect 2775 2045 2779 2046
rect 2895 2050 2899 2051
rect 2895 2045 2899 2046
rect 2919 2050 2923 2051
rect 2919 2045 2923 2046
rect 3039 2050 3043 2051
rect 3039 2045 3043 2046
rect 3079 2050 3083 2051
rect 3079 2045 3083 2046
rect 3191 2050 3195 2051
rect 3191 2045 3195 2046
rect 3263 2050 3267 2051
rect 3263 2045 3267 2046
rect 3351 2050 3355 2051
rect 3351 2045 3355 2046
rect 3455 2050 3459 2051
rect 3455 2045 3459 2046
rect 3519 2050 3523 2051
rect 3519 2045 3523 2046
rect 3655 2050 3659 2051
rect 3655 2045 3659 2046
rect 3687 2050 3691 2051
rect 3687 2045 3691 2046
rect 3839 2050 3843 2051
rect 3839 2045 3843 2046
rect 3943 2050 3947 2051
rect 3943 2045 3947 2046
rect 2048 2018 2050 2045
rect 2328 2021 2330 2045
rect 2432 2021 2434 2045
rect 2536 2021 2538 2045
rect 2648 2021 2650 2045
rect 2776 2021 2778 2045
rect 2920 2021 2922 2045
rect 3080 2021 3082 2045
rect 3264 2021 3266 2045
rect 3456 2021 3458 2045
rect 3656 2021 3658 2045
rect 3840 2021 3842 2045
rect 2326 2020 2332 2021
rect 2046 2017 2052 2018
rect 111 2014 115 2015
rect 111 2009 115 2010
rect 447 2014 451 2015
rect 447 2009 451 2010
rect 575 2014 579 2015
rect 575 2009 579 2010
rect 623 2014 627 2015
rect 623 2009 627 2010
rect 727 2014 731 2015
rect 727 2009 731 2010
rect 735 2014 739 2015
rect 735 2009 739 2010
rect 855 2014 859 2015
rect 855 2009 859 2010
rect 887 2014 891 2015
rect 887 2009 891 2010
rect 983 2014 987 2015
rect 983 2009 987 2010
rect 1055 2014 1059 2015
rect 1055 2009 1059 2010
rect 1119 2014 1123 2015
rect 1119 2009 1123 2010
rect 1231 2014 1235 2015
rect 1231 2009 1235 2010
rect 1255 2014 1259 2015
rect 1255 2009 1259 2010
rect 1391 2014 1395 2015
rect 1391 2009 1395 2010
rect 1399 2014 1403 2015
rect 1399 2009 1403 2010
rect 1527 2014 1531 2015
rect 1527 2009 1531 2010
rect 1575 2014 1579 2015
rect 1575 2009 1579 2010
rect 1655 2014 1659 2015
rect 1655 2009 1659 2010
rect 1751 2014 1755 2015
rect 1751 2009 1755 2010
rect 1791 2014 1795 2015
rect 1791 2009 1795 2010
rect 1903 2014 1907 2015
rect 1903 2009 1907 2010
rect 2007 2014 2011 2015
rect 2046 2013 2047 2017
rect 2051 2013 2052 2017
rect 2326 2016 2327 2020
rect 2331 2016 2332 2020
rect 2326 2015 2332 2016
rect 2430 2020 2436 2021
rect 2430 2016 2431 2020
rect 2435 2016 2436 2020
rect 2430 2015 2436 2016
rect 2534 2020 2540 2021
rect 2534 2016 2535 2020
rect 2539 2016 2540 2020
rect 2534 2015 2540 2016
rect 2646 2020 2652 2021
rect 2646 2016 2647 2020
rect 2651 2016 2652 2020
rect 2646 2015 2652 2016
rect 2774 2020 2780 2021
rect 2774 2016 2775 2020
rect 2779 2016 2780 2020
rect 2774 2015 2780 2016
rect 2918 2020 2924 2021
rect 2918 2016 2919 2020
rect 2923 2016 2924 2020
rect 2918 2015 2924 2016
rect 3078 2020 3084 2021
rect 3078 2016 3079 2020
rect 3083 2016 3084 2020
rect 3078 2015 3084 2016
rect 3262 2020 3268 2021
rect 3262 2016 3263 2020
rect 3267 2016 3268 2020
rect 3262 2015 3268 2016
rect 3454 2020 3460 2021
rect 3454 2016 3455 2020
rect 3459 2016 3460 2020
rect 3454 2015 3460 2016
rect 3654 2020 3660 2021
rect 3654 2016 3655 2020
rect 3659 2016 3660 2020
rect 3654 2015 3660 2016
rect 3838 2020 3844 2021
rect 3838 2016 3839 2020
rect 3843 2016 3844 2020
rect 3944 2018 3946 2045
rect 3838 2015 3844 2016
rect 3942 2017 3948 2018
rect 2046 2012 2052 2013
rect 3942 2013 3943 2017
rect 3947 2013 3948 2017
rect 3942 2012 3948 2013
rect 2007 2009 2011 2010
rect 112 1982 114 2009
rect 448 1985 450 2009
rect 576 1985 578 2009
rect 728 1985 730 2009
rect 888 1985 890 2009
rect 1056 1985 1058 2009
rect 1232 1985 1234 2009
rect 1400 1985 1402 2009
rect 1576 1985 1578 2009
rect 1752 1985 1754 2009
rect 1904 1985 1906 2009
rect 446 1984 452 1985
rect 110 1981 116 1982
rect 110 1977 111 1981
rect 115 1977 116 1981
rect 446 1980 447 1984
rect 451 1980 452 1984
rect 446 1979 452 1980
rect 574 1984 580 1985
rect 574 1980 575 1984
rect 579 1980 580 1984
rect 574 1979 580 1980
rect 726 1984 732 1985
rect 726 1980 727 1984
rect 731 1980 732 1984
rect 726 1979 732 1980
rect 886 1984 892 1985
rect 886 1980 887 1984
rect 891 1980 892 1984
rect 886 1979 892 1980
rect 1054 1984 1060 1985
rect 1054 1980 1055 1984
rect 1059 1980 1060 1984
rect 1054 1979 1060 1980
rect 1230 1984 1236 1985
rect 1230 1980 1231 1984
rect 1235 1980 1236 1984
rect 1230 1979 1236 1980
rect 1398 1984 1404 1985
rect 1398 1980 1399 1984
rect 1403 1980 1404 1984
rect 1398 1979 1404 1980
rect 1574 1984 1580 1985
rect 1574 1980 1575 1984
rect 1579 1980 1580 1984
rect 1574 1979 1580 1980
rect 1750 1984 1756 1985
rect 1750 1980 1751 1984
rect 1755 1980 1756 1984
rect 1750 1979 1756 1980
rect 1902 1984 1908 1985
rect 1902 1980 1903 1984
rect 1907 1980 1908 1984
rect 2008 1982 2010 2009
rect 2326 2001 2332 2002
rect 2046 2000 2052 2001
rect 2046 1996 2047 2000
rect 2051 1996 2052 2000
rect 2326 1997 2327 2001
rect 2331 1997 2332 2001
rect 2326 1996 2332 1997
rect 2430 2001 2436 2002
rect 2430 1997 2431 2001
rect 2435 1997 2436 2001
rect 2430 1996 2436 1997
rect 2534 2001 2540 2002
rect 2534 1997 2535 2001
rect 2539 1997 2540 2001
rect 2534 1996 2540 1997
rect 2646 2001 2652 2002
rect 2646 1997 2647 2001
rect 2651 1997 2652 2001
rect 2646 1996 2652 1997
rect 2774 2001 2780 2002
rect 2774 1997 2775 2001
rect 2779 1997 2780 2001
rect 2774 1996 2780 1997
rect 2918 2001 2924 2002
rect 2918 1997 2919 2001
rect 2923 1997 2924 2001
rect 2918 1996 2924 1997
rect 3078 2001 3084 2002
rect 3078 1997 3079 2001
rect 3083 1997 3084 2001
rect 3078 1996 3084 1997
rect 3262 2001 3268 2002
rect 3262 1997 3263 2001
rect 3267 1997 3268 2001
rect 3262 1996 3268 1997
rect 3454 2001 3460 2002
rect 3454 1997 3455 2001
rect 3459 1997 3460 2001
rect 3454 1996 3460 1997
rect 3654 2001 3660 2002
rect 3654 1997 3655 2001
rect 3659 1997 3660 2001
rect 3654 1996 3660 1997
rect 3838 2001 3844 2002
rect 3838 1997 3839 2001
rect 3843 1997 3844 2001
rect 3838 1996 3844 1997
rect 3942 2000 3948 2001
rect 3942 1996 3943 2000
rect 3947 1996 3948 2000
rect 2046 1995 2052 1996
rect 1902 1979 1908 1980
rect 2006 1981 2012 1982
rect 110 1976 116 1977
rect 2006 1977 2007 1981
rect 2011 1977 2012 1981
rect 2006 1976 2012 1977
rect 2048 1971 2050 1995
rect 2328 1971 2330 1996
rect 2432 1971 2434 1996
rect 2536 1971 2538 1996
rect 2648 1971 2650 1996
rect 2776 1971 2778 1996
rect 2920 1971 2922 1996
rect 3080 1971 3082 1996
rect 3264 1971 3266 1996
rect 3456 1971 3458 1996
rect 3656 1971 3658 1996
rect 3840 1971 3842 1996
rect 3942 1995 3948 1996
rect 3944 1971 3946 1995
rect 2047 1970 2051 1971
rect 446 1965 452 1966
rect 110 1964 116 1965
rect 110 1960 111 1964
rect 115 1960 116 1964
rect 446 1961 447 1965
rect 451 1961 452 1965
rect 446 1960 452 1961
rect 574 1965 580 1966
rect 574 1961 575 1965
rect 579 1961 580 1965
rect 574 1960 580 1961
rect 726 1965 732 1966
rect 726 1961 727 1965
rect 731 1961 732 1965
rect 726 1960 732 1961
rect 886 1965 892 1966
rect 886 1961 887 1965
rect 891 1961 892 1965
rect 886 1960 892 1961
rect 1054 1965 1060 1966
rect 1054 1961 1055 1965
rect 1059 1961 1060 1965
rect 1054 1960 1060 1961
rect 1230 1965 1236 1966
rect 1230 1961 1231 1965
rect 1235 1961 1236 1965
rect 1230 1960 1236 1961
rect 1398 1965 1404 1966
rect 1398 1961 1399 1965
rect 1403 1961 1404 1965
rect 1398 1960 1404 1961
rect 1574 1965 1580 1966
rect 1574 1961 1575 1965
rect 1579 1961 1580 1965
rect 1574 1960 1580 1961
rect 1750 1965 1756 1966
rect 1750 1961 1751 1965
rect 1755 1961 1756 1965
rect 1750 1960 1756 1961
rect 1902 1965 1908 1966
rect 2047 1965 2051 1966
rect 2255 1970 2259 1971
rect 2255 1965 2259 1966
rect 2327 1970 2331 1971
rect 2327 1965 2331 1966
rect 2351 1970 2355 1971
rect 2351 1965 2355 1966
rect 2431 1970 2435 1971
rect 2431 1965 2435 1966
rect 2447 1970 2451 1971
rect 2447 1965 2451 1966
rect 2535 1970 2539 1971
rect 2535 1965 2539 1966
rect 2543 1970 2547 1971
rect 2543 1965 2547 1966
rect 2647 1970 2651 1971
rect 2647 1965 2651 1966
rect 2767 1970 2771 1971
rect 2767 1965 2771 1966
rect 2775 1970 2779 1971
rect 2775 1965 2779 1966
rect 2919 1970 2923 1971
rect 2919 1965 2923 1966
rect 3079 1970 3083 1971
rect 3079 1965 3083 1966
rect 3103 1970 3107 1971
rect 3103 1965 3107 1966
rect 3263 1970 3267 1971
rect 3263 1965 3267 1966
rect 3319 1970 3323 1971
rect 3319 1965 3323 1966
rect 3455 1970 3459 1971
rect 3455 1965 3459 1966
rect 3543 1970 3547 1971
rect 3543 1965 3547 1966
rect 3655 1970 3659 1971
rect 3655 1965 3659 1966
rect 3775 1970 3779 1971
rect 3775 1965 3779 1966
rect 3839 1970 3843 1971
rect 3839 1965 3843 1966
rect 3943 1970 3947 1971
rect 3943 1965 3947 1966
rect 1902 1961 1903 1965
rect 1907 1961 1908 1965
rect 1902 1960 1908 1961
rect 2006 1964 2012 1965
rect 2006 1960 2007 1964
rect 2011 1960 2012 1964
rect 110 1959 116 1960
rect 112 1939 114 1959
rect 448 1939 450 1960
rect 576 1939 578 1960
rect 728 1939 730 1960
rect 888 1939 890 1960
rect 1056 1939 1058 1960
rect 1232 1939 1234 1960
rect 1400 1939 1402 1960
rect 1576 1939 1578 1960
rect 1752 1939 1754 1960
rect 1904 1939 1906 1960
rect 2006 1959 2012 1960
rect 2008 1939 2010 1959
rect 2048 1945 2050 1965
rect 2046 1944 2052 1945
rect 2256 1944 2258 1965
rect 2352 1944 2354 1965
rect 2448 1944 2450 1965
rect 2544 1944 2546 1965
rect 2648 1944 2650 1965
rect 2768 1944 2770 1965
rect 2920 1944 2922 1965
rect 3104 1944 3106 1965
rect 3320 1944 3322 1965
rect 3544 1944 3546 1965
rect 3776 1944 3778 1965
rect 3944 1945 3946 1965
rect 3942 1944 3948 1945
rect 2046 1940 2047 1944
rect 2051 1940 2052 1944
rect 2046 1939 2052 1940
rect 2254 1943 2260 1944
rect 2254 1939 2255 1943
rect 2259 1939 2260 1943
rect 111 1938 115 1939
rect 111 1933 115 1934
rect 447 1938 451 1939
rect 447 1933 451 1934
rect 575 1938 579 1939
rect 575 1933 579 1934
rect 655 1938 659 1939
rect 655 1933 659 1934
rect 727 1938 731 1939
rect 727 1933 731 1934
rect 751 1938 755 1939
rect 751 1933 755 1934
rect 847 1938 851 1939
rect 847 1933 851 1934
rect 887 1938 891 1939
rect 887 1933 891 1934
rect 943 1938 947 1939
rect 943 1933 947 1934
rect 1039 1938 1043 1939
rect 1039 1933 1043 1934
rect 1055 1938 1059 1939
rect 1055 1933 1059 1934
rect 1135 1938 1139 1939
rect 1135 1933 1139 1934
rect 1231 1938 1235 1939
rect 1231 1933 1235 1934
rect 1327 1938 1331 1939
rect 1327 1933 1331 1934
rect 1399 1938 1403 1939
rect 1399 1933 1403 1934
rect 1423 1938 1427 1939
rect 1423 1933 1427 1934
rect 1575 1938 1579 1939
rect 1575 1933 1579 1934
rect 1751 1938 1755 1939
rect 1751 1933 1755 1934
rect 1903 1938 1907 1939
rect 1903 1933 1907 1934
rect 2007 1938 2011 1939
rect 2254 1938 2260 1939
rect 2350 1943 2356 1944
rect 2350 1939 2351 1943
rect 2355 1939 2356 1943
rect 2350 1938 2356 1939
rect 2446 1943 2452 1944
rect 2446 1939 2447 1943
rect 2451 1939 2452 1943
rect 2446 1938 2452 1939
rect 2542 1943 2548 1944
rect 2542 1939 2543 1943
rect 2547 1939 2548 1943
rect 2542 1938 2548 1939
rect 2646 1943 2652 1944
rect 2646 1939 2647 1943
rect 2651 1939 2652 1943
rect 2646 1938 2652 1939
rect 2766 1943 2772 1944
rect 2766 1939 2767 1943
rect 2771 1939 2772 1943
rect 2766 1938 2772 1939
rect 2918 1943 2924 1944
rect 2918 1939 2919 1943
rect 2923 1939 2924 1943
rect 2918 1938 2924 1939
rect 3102 1943 3108 1944
rect 3102 1939 3103 1943
rect 3107 1939 3108 1943
rect 3102 1938 3108 1939
rect 3318 1943 3324 1944
rect 3318 1939 3319 1943
rect 3323 1939 3324 1943
rect 3318 1938 3324 1939
rect 3542 1943 3548 1944
rect 3542 1939 3543 1943
rect 3547 1939 3548 1943
rect 3542 1938 3548 1939
rect 3774 1943 3780 1944
rect 3774 1939 3775 1943
rect 3779 1939 3780 1943
rect 3942 1940 3943 1944
rect 3947 1940 3948 1944
rect 3942 1939 3948 1940
rect 3774 1938 3780 1939
rect 2007 1933 2011 1934
rect 112 1913 114 1933
rect 110 1912 116 1913
rect 656 1912 658 1933
rect 752 1912 754 1933
rect 848 1912 850 1933
rect 944 1912 946 1933
rect 1040 1912 1042 1933
rect 1136 1912 1138 1933
rect 1232 1912 1234 1933
rect 1328 1912 1330 1933
rect 1424 1912 1426 1933
rect 2008 1913 2010 1933
rect 2046 1927 2052 1928
rect 2046 1923 2047 1927
rect 2051 1923 2052 1927
rect 3942 1927 3948 1928
rect 2046 1922 2052 1923
rect 2254 1924 2260 1925
rect 2006 1912 2012 1913
rect 110 1908 111 1912
rect 115 1908 116 1912
rect 110 1907 116 1908
rect 654 1911 660 1912
rect 654 1907 655 1911
rect 659 1907 660 1911
rect 654 1906 660 1907
rect 750 1911 756 1912
rect 750 1907 751 1911
rect 755 1907 756 1911
rect 750 1906 756 1907
rect 846 1911 852 1912
rect 846 1907 847 1911
rect 851 1907 852 1911
rect 846 1906 852 1907
rect 942 1911 948 1912
rect 942 1907 943 1911
rect 947 1907 948 1911
rect 942 1906 948 1907
rect 1038 1911 1044 1912
rect 1038 1907 1039 1911
rect 1043 1907 1044 1911
rect 1038 1906 1044 1907
rect 1134 1911 1140 1912
rect 1134 1907 1135 1911
rect 1139 1907 1140 1911
rect 1134 1906 1140 1907
rect 1230 1911 1236 1912
rect 1230 1907 1231 1911
rect 1235 1907 1236 1911
rect 1230 1906 1236 1907
rect 1326 1911 1332 1912
rect 1326 1907 1327 1911
rect 1331 1907 1332 1911
rect 1326 1906 1332 1907
rect 1422 1911 1428 1912
rect 1422 1907 1423 1911
rect 1427 1907 1428 1911
rect 2006 1908 2007 1912
rect 2011 1908 2012 1912
rect 2006 1907 2012 1908
rect 1422 1906 1428 1907
rect 110 1895 116 1896
rect 110 1891 111 1895
rect 115 1891 116 1895
rect 2006 1895 2012 1896
rect 110 1890 116 1891
rect 654 1892 660 1893
rect 112 1863 114 1890
rect 654 1888 655 1892
rect 659 1888 660 1892
rect 654 1887 660 1888
rect 750 1892 756 1893
rect 750 1888 751 1892
rect 755 1888 756 1892
rect 750 1887 756 1888
rect 846 1892 852 1893
rect 846 1888 847 1892
rect 851 1888 852 1892
rect 846 1887 852 1888
rect 942 1892 948 1893
rect 942 1888 943 1892
rect 947 1888 948 1892
rect 942 1887 948 1888
rect 1038 1892 1044 1893
rect 1038 1888 1039 1892
rect 1043 1888 1044 1892
rect 1038 1887 1044 1888
rect 1134 1892 1140 1893
rect 1134 1888 1135 1892
rect 1139 1888 1140 1892
rect 1134 1887 1140 1888
rect 1230 1892 1236 1893
rect 1230 1888 1231 1892
rect 1235 1888 1236 1892
rect 1230 1887 1236 1888
rect 1326 1892 1332 1893
rect 1326 1888 1327 1892
rect 1331 1888 1332 1892
rect 1326 1887 1332 1888
rect 1422 1892 1428 1893
rect 1422 1888 1423 1892
rect 1427 1888 1428 1892
rect 2006 1891 2007 1895
rect 2011 1891 2012 1895
rect 2006 1890 2012 1891
rect 1422 1887 1428 1888
rect 656 1863 658 1887
rect 752 1863 754 1887
rect 848 1863 850 1887
rect 944 1863 946 1887
rect 1040 1863 1042 1887
rect 1136 1863 1138 1887
rect 1232 1863 1234 1887
rect 1328 1863 1330 1887
rect 1424 1863 1426 1887
rect 2008 1863 2010 1890
rect 2048 1883 2050 1922
rect 2254 1920 2255 1924
rect 2259 1920 2260 1924
rect 2254 1919 2260 1920
rect 2350 1924 2356 1925
rect 2350 1920 2351 1924
rect 2355 1920 2356 1924
rect 2350 1919 2356 1920
rect 2446 1924 2452 1925
rect 2446 1920 2447 1924
rect 2451 1920 2452 1924
rect 2446 1919 2452 1920
rect 2542 1924 2548 1925
rect 2542 1920 2543 1924
rect 2547 1920 2548 1924
rect 2542 1919 2548 1920
rect 2646 1924 2652 1925
rect 2646 1920 2647 1924
rect 2651 1920 2652 1924
rect 2646 1919 2652 1920
rect 2766 1924 2772 1925
rect 2766 1920 2767 1924
rect 2771 1920 2772 1924
rect 2766 1919 2772 1920
rect 2918 1924 2924 1925
rect 2918 1920 2919 1924
rect 2923 1920 2924 1924
rect 2918 1919 2924 1920
rect 3102 1924 3108 1925
rect 3102 1920 3103 1924
rect 3107 1920 3108 1924
rect 3102 1919 3108 1920
rect 3318 1924 3324 1925
rect 3318 1920 3319 1924
rect 3323 1920 3324 1924
rect 3318 1919 3324 1920
rect 3542 1924 3548 1925
rect 3542 1920 3543 1924
rect 3547 1920 3548 1924
rect 3542 1919 3548 1920
rect 3774 1924 3780 1925
rect 3774 1920 3775 1924
rect 3779 1920 3780 1924
rect 3942 1923 3943 1927
rect 3947 1923 3948 1927
rect 3942 1922 3948 1923
rect 3774 1919 3780 1920
rect 2256 1883 2258 1919
rect 2352 1883 2354 1919
rect 2448 1883 2450 1919
rect 2544 1883 2546 1919
rect 2648 1883 2650 1919
rect 2768 1883 2770 1919
rect 2920 1883 2922 1919
rect 3104 1883 3106 1919
rect 3320 1883 3322 1919
rect 3544 1883 3546 1919
rect 3776 1883 3778 1919
rect 3944 1883 3946 1922
rect 2047 1882 2051 1883
rect 2047 1877 2051 1878
rect 2183 1882 2187 1883
rect 2183 1877 2187 1878
rect 2255 1882 2259 1883
rect 2255 1877 2259 1878
rect 2279 1882 2283 1883
rect 2279 1877 2283 1878
rect 2351 1882 2355 1883
rect 2351 1877 2355 1878
rect 2383 1882 2387 1883
rect 2383 1877 2387 1878
rect 2447 1882 2451 1883
rect 2447 1877 2451 1878
rect 2487 1882 2491 1883
rect 2487 1877 2491 1878
rect 2543 1882 2547 1883
rect 2543 1877 2547 1878
rect 2591 1882 2595 1883
rect 2591 1877 2595 1878
rect 2647 1882 2651 1883
rect 2647 1877 2651 1878
rect 2703 1882 2707 1883
rect 2703 1877 2707 1878
rect 2767 1882 2771 1883
rect 2767 1877 2771 1878
rect 2831 1882 2835 1883
rect 2831 1877 2835 1878
rect 2919 1882 2923 1883
rect 2919 1877 2923 1878
rect 2991 1882 2995 1883
rect 2991 1877 2995 1878
rect 3103 1882 3107 1883
rect 3103 1877 3107 1878
rect 3183 1882 3187 1883
rect 3183 1877 3187 1878
rect 3319 1882 3323 1883
rect 3319 1877 3323 1878
rect 3399 1882 3403 1883
rect 3399 1877 3403 1878
rect 3543 1882 3547 1883
rect 3543 1877 3547 1878
rect 3631 1882 3635 1883
rect 3631 1877 3635 1878
rect 3775 1882 3779 1883
rect 3775 1877 3779 1878
rect 3839 1882 3843 1883
rect 3839 1877 3843 1878
rect 3943 1882 3947 1883
rect 3943 1877 3947 1878
rect 111 1862 115 1863
rect 111 1857 115 1858
rect 319 1862 323 1863
rect 319 1857 323 1858
rect 447 1862 451 1863
rect 447 1857 451 1858
rect 583 1862 587 1863
rect 583 1857 587 1858
rect 655 1862 659 1863
rect 655 1857 659 1858
rect 719 1862 723 1863
rect 719 1857 723 1858
rect 751 1862 755 1863
rect 751 1857 755 1858
rect 847 1862 851 1863
rect 847 1857 851 1858
rect 855 1862 859 1863
rect 855 1857 859 1858
rect 943 1862 947 1863
rect 943 1857 947 1858
rect 991 1862 995 1863
rect 991 1857 995 1858
rect 1039 1862 1043 1863
rect 1039 1857 1043 1858
rect 1127 1862 1131 1863
rect 1127 1857 1131 1858
rect 1135 1862 1139 1863
rect 1135 1857 1139 1858
rect 1231 1862 1235 1863
rect 1231 1857 1235 1858
rect 1263 1862 1267 1863
rect 1263 1857 1267 1858
rect 1327 1862 1331 1863
rect 1327 1857 1331 1858
rect 1399 1862 1403 1863
rect 1399 1857 1403 1858
rect 1423 1862 1427 1863
rect 1423 1857 1427 1858
rect 1535 1862 1539 1863
rect 1535 1857 1539 1858
rect 2007 1862 2011 1863
rect 2007 1857 2011 1858
rect 112 1830 114 1857
rect 320 1833 322 1857
rect 448 1833 450 1857
rect 584 1833 586 1857
rect 720 1833 722 1857
rect 856 1833 858 1857
rect 992 1833 994 1857
rect 1128 1833 1130 1857
rect 1264 1833 1266 1857
rect 1400 1833 1402 1857
rect 1536 1833 1538 1857
rect 318 1832 324 1833
rect 110 1829 116 1830
rect 110 1825 111 1829
rect 115 1825 116 1829
rect 318 1828 319 1832
rect 323 1828 324 1832
rect 318 1827 324 1828
rect 446 1832 452 1833
rect 446 1828 447 1832
rect 451 1828 452 1832
rect 446 1827 452 1828
rect 582 1832 588 1833
rect 582 1828 583 1832
rect 587 1828 588 1832
rect 582 1827 588 1828
rect 718 1832 724 1833
rect 718 1828 719 1832
rect 723 1828 724 1832
rect 718 1827 724 1828
rect 854 1832 860 1833
rect 854 1828 855 1832
rect 859 1828 860 1832
rect 854 1827 860 1828
rect 990 1832 996 1833
rect 990 1828 991 1832
rect 995 1828 996 1832
rect 990 1827 996 1828
rect 1126 1832 1132 1833
rect 1126 1828 1127 1832
rect 1131 1828 1132 1832
rect 1126 1827 1132 1828
rect 1262 1832 1268 1833
rect 1262 1828 1263 1832
rect 1267 1828 1268 1832
rect 1262 1827 1268 1828
rect 1398 1832 1404 1833
rect 1398 1828 1399 1832
rect 1403 1828 1404 1832
rect 1398 1827 1404 1828
rect 1534 1832 1540 1833
rect 1534 1828 1535 1832
rect 1539 1828 1540 1832
rect 2008 1830 2010 1857
rect 2048 1850 2050 1877
rect 2184 1853 2186 1877
rect 2280 1853 2282 1877
rect 2384 1853 2386 1877
rect 2488 1853 2490 1877
rect 2592 1853 2594 1877
rect 2704 1853 2706 1877
rect 2832 1853 2834 1877
rect 2992 1853 2994 1877
rect 3184 1853 3186 1877
rect 3400 1853 3402 1877
rect 3632 1853 3634 1877
rect 3840 1853 3842 1877
rect 2182 1852 2188 1853
rect 2046 1849 2052 1850
rect 2046 1845 2047 1849
rect 2051 1845 2052 1849
rect 2182 1848 2183 1852
rect 2187 1848 2188 1852
rect 2182 1847 2188 1848
rect 2278 1852 2284 1853
rect 2278 1848 2279 1852
rect 2283 1848 2284 1852
rect 2278 1847 2284 1848
rect 2382 1852 2388 1853
rect 2382 1848 2383 1852
rect 2387 1848 2388 1852
rect 2382 1847 2388 1848
rect 2486 1852 2492 1853
rect 2486 1848 2487 1852
rect 2491 1848 2492 1852
rect 2486 1847 2492 1848
rect 2590 1852 2596 1853
rect 2590 1848 2591 1852
rect 2595 1848 2596 1852
rect 2590 1847 2596 1848
rect 2702 1852 2708 1853
rect 2702 1848 2703 1852
rect 2707 1848 2708 1852
rect 2702 1847 2708 1848
rect 2830 1852 2836 1853
rect 2830 1848 2831 1852
rect 2835 1848 2836 1852
rect 2830 1847 2836 1848
rect 2990 1852 2996 1853
rect 2990 1848 2991 1852
rect 2995 1848 2996 1852
rect 2990 1847 2996 1848
rect 3182 1852 3188 1853
rect 3182 1848 3183 1852
rect 3187 1848 3188 1852
rect 3182 1847 3188 1848
rect 3398 1852 3404 1853
rect 3398 1848 3399 1852
rect 3403 1848 3404 1852
rect 3398 1847 3404 1848
rect 3630 1852 3636 1853
rect 3630 1848 3631 1852
rect 3635 1848 3636 1852
rect 3630 1847 3636 1848
rect 3838 1852 3844 1853
rect 3838 1848 3839 1852
rect 3843 1848 3844 1852
rect 3944 1850 3946 1877
rect 3838 1847 3844 1848
rect 3942 1849 3948 1850
rect 2046 1844 2052 1845
rect 3942 1845 3943 1849
rect 3947 1845 3948 1849
rect 3942 1844 3948 1845
rect 2182 1833 2188 1834
rect 2046 1832 2052 1833
rect 1534 1827 1540 1828
rect 2006 1829 2012 1830
rect 110 1824 116 1825
rect 2006 1825 2007 1829
rect 2011 1825 2012 1829
rect 2046 1828 2047 1832
rect 2051 1828 2052 1832
rect 2182 1829 2183 1833
rect 2187 1829 2188 1833
rect 2182 1828 2188 1829
rect 2278 1833 2284 1834
rect 2278 1829 2279 1833
rect 2283 1829 2284 1833
rect 2278 1828 2284 1829
rect 2382 1833 2388 1834
rect 2382 1829 2383 1833
rect 2387 1829 2388 1833
rect 2382 1828 2388 1829
rect 2486 1833 2492 1834
rect 2486 1829 2487 1833
rect 2491 1829 2492 1833
rect 2486 1828 2492 1829
rect 2590 1833 2596 1834
rect 2590 1829 2591 1833
rect 2595 1829 2596 1833
rect 2590 1828 2596 1829
rect 2702 1833 2708 1834
rect 2702 1829 2703 1833
rect 2707 1829 2708 1833
rect 2702 1828 2708 1829
rect 2830 1833 2836 1834
rect 2830 1829 2831 1833
rect 2835 1829 2836 1833
rect 2830 1828 2836 1829
rect 2990 1833 2996 1834
rect 2990 1829 2991 1833
rect 2995 1829 2996 1833
rect 2990 1828 2996 1829
rect 3182 1833 3188 1834
rect 3182 1829 3183 1833
rect 3187 1829 3188 1833
rect 3182 1828 3188 1829
rect 3398 1833 3404 1834
rect 3398 1829 3399 1833
rect 3403 1829 3404 1833
rect 3398 1828 3404 1829
rect 3630 1833 3636 1834
rect 3630 1829 3631 1833
rect 3635 1829 3636 1833
rect 3630 1828 3636 1829
rect 3838 1833 3844 1834
rect 3838 1829 3839 1833
rect 3843 1829 3844 1833
rect 3838 1828 3844 1829
rect 3942 1832 3948 1833
rect 3942 1828 3943 1832
rect 3947 1828 3948 1832
rect 2046 1827 2052 1828
rect 2006 1824 2012 1825
rect 318 1813 324 1814
rect 110 1812 116 1813
rect 110 1808 111 1812
rect 115 1808 116 1812
rect 318 1809 319 1813
rect 323 1809 324 1813
rect 318 1808 324 1809
rect 446 1813 452 1814
rect 446 1809 447 1813
rect 451 1809 452 1813
rect 446 1808 452 1809
rect 582 1813 588 1814
rect 582 1809 583 1813
rect 587 1809 588 1813
rect 582 1808 588 1809
rect 718 1813 724 1814
rect 718 1809 719 1813
rect 723 1809 724 1813
rect 718 1808 724 1809
rect 854 1813 860 1814
rect 854 1809 855 1813
rect 859 1809 860 1813
rect 854 1808 860 1809
rect 990 1813 996 1814
rect 990 1809 991 1813
rect 995 1809 996 1813
rect 990 1808 996 1809
rect 1126 1813 1132 1814
rect 1126 1809 1127 1813
rect 1131 1809 1132 1813
rect 1126 1808 1132 1809
rect 1262 1813 1268 1814
rect 1262 1809 1263 1813
rect 1267 1809 1268 1813
rect 1262 1808 1268 1809
rect 1398 1813 1404 1814
rect 1398 1809 1399 1813
rect 1403 1809 1404 1813
rect 1398 1808 1404 1809
rect 1534 1813 1540 1814
rect 1534 1809 1535 1813
rect 1539 1809 1540 1813
rect 1534 1808 1540 1809
rect 2006 1812 2012 1813
rect 2006 1808 2007 1812
rect 2011 1808 2012 1812
rect 110 1807 116 1808
rect 112 1783 114 1807
rect 320 1783 322 1808
rect 448 1783 450 1808
rect 584 1783 586 1808
rect 720 1783 722 1808
rect 856 1783 858 1808
rect 992 1783 994 1808
rect 1128 1783 1130 1808
rect 1264 1783 1266 1808
rect 1400 1783 1402 1808
rect 1536 1783 1538 1808
rect 2006 1807 2012 1808
rect 2008 1783 2010 1807
rect 2048 1803 2050 1827
rect 2184 1803 2186 1828
rect 2280 1803 2282 1828
rect 2384 1803 2386 1828
rect 2488 1803 2490 1828
rect 2592 1803 2594 1828
rect 2704 1803 2706 1828
rect 2832 1803 2834 1828
rect 2992 1803 2994 1828
rect 3184 1803 3186 1828
rect 3400 1803 3402 1828
rect 3632 1803 3634 1828
rect 3840 1803 3842 1828
rect 3942 1827 3948 1828
rect 3944 1803 3946 1827
rect 2047 1802 2051 1803
rect 2047 1797 2051 1798
rect 2127 1802 2131 1803
rect 2127 1797 2131 1798
rect 2183 1802 2187 1803
rect 2183 1797 2187 1798
rect 2279 1802 2283 1803
rect 2279 1797 2283 1798
rect 2311 1802 2315 1803
rect 2311 1797 2315 1798
rect 2383 1802 2387 1803
rect 2383 1797 2387 1798
rect 2487 1802 2491 1803
rect 2487 1797 2491 1798
rect 2495 1802 2499 1803
rect 2495 1797 2499 1798
rect 2591 1802 2595 1803
rect 2591 1797 2595 1798
rect 2687 1802 2691 1803
rect 2687 1797 2691 1798
rect 2703 1802 2707 1803
rect 2703 1797 2707 1798
rect 2831 1802 2835 1803
rect 2831 1797 2835 1798
rect 2879 1802 2883 1803
rect 2879 1797 2883 1798
rect 2991 1802 2995 1803
rect 2991 1797 2995 1798
rect 3071 1802 3075 1803
rect 3071 1797 3075 1798
rect 3183 1802 3187 1803
rect 3183 1797 3187 1798
rect 3263 1802 3267 1803
rect 3263 1797 3267 1798
rect 3399 1802 3403 1803
rect 3399 1797 3403 1798
rect 3463 1802 3467 1803
rect 3463 1797 3467 1798
rect 3631 1802 3635 1803
rect 3631 1797 3635 1798
rect 3663 1802 3667 1803
rect 3663 1797 3667 1798
rect 3839 1802 3843 1803
rect 3839 1797 3843 1798
rect 3943 1802 3947 1803
rect 3943 1797 3947 1798
rect 111 1782 115 1783
rect 111 1777 115 1778
rect 255 1782 259 1783
rect 255 1777 259 1778
rect 319 1782 323 1783
rect 319 1777 323 1778
rect 391 1782 395 1783
rect 391 1777 395 1778
rect 447 1782 451 1783
rect 447 1777 451 1778
rect 535 1782 539 1783
rect 535 1777 539 1778
rect 583 1782 587 1783
rect 583 1777 587 1778
rect 695 1782 699 1783
rect 695 1777 699 1778
rect 719 1782 723 1783
rect 719 1777 723 1778
rect 855 1782 859 1783
rect 855 1777 859 1778
rect 863 1782 867 1783
rect 863 1777 867 1778
rect 991 1782 995 1783
rect 991 1777 995 1778
rect 1031 1782 1035 1783
rect 1031 1777 1035 1778
rect 1127 1782 1131 1783
rect 1127 1777 1131 1778
rect 1207 1782 1211 1783
rect 1207 1777 1211 1778
rect 1263 1782 1267 1783
rect 1263 1777 1267 1778
rect 1383 1782 1387 1783
rect 1383 1777 1387 1778
rect 1399 1782 1403 1783
rect 1399 1777 1403 1778
rect 1535 1782 1539 1783
rect 1535 1777 1539 1778
rect 1559 1782 1563 1783
rect 1559 1777 1563 1778
rect 1743 1782 1747 1783
rect 1743 1777 1747 1778
rect 2007 1782 2011 1783
rect 2007 1777 2011 1778
rect 2048 1777 2050 1797
rect 112 1757 114 1777
rect 110 1756 116 1757
rect 256 1756 258 1777
rect 392 1756 394 1777
rect 536 1756 538 1777
rect 696 1756 698 1777
rect 864 1756 866 1777
rect 1032 1756 1034 1777
rect 1208 1756 1210 1777
rect 1384 1756 1386 1777
rect 1560 1756 1562 1777
rect 1744 1756 1746 1777
rect 2008 1757 2010 1777
rect 2046 1776 2052 1777
rect 2128 1776 2130 1797
rect 2312 1776 2314 1797
rect 2496 1776 2498 1797
rect 2688 1776 2690 1797
rect 2880 1776 2882 1797
rect 3072 1776 3074 1797
rect 3264 1776 3266 1797
rect 3464 1776 3466 1797
rect 3664 1776 3666 1797
rect 3840 1776 3842 1797
rect 3944 1777 3946 1797
rect 3942 1776 3948 1777
rect 2046 1772 2047 1776
rect 2051 1772 2052 1776
rect 2046 1771 2052 1772
rect 2126 1775 2132 1776
rect 2126 1771 2127 1775
rect 2131 1771 2132 1775
rect 2126 1770 2132 1771
rect 2310 1775 2316 1776
rect 2310 1771 2311 1775
rect 2315 1771 2316 1775
rect 2310 1770 2316 1771
rect 2494 1775 2500 1776
rect 2494 1771 2495 1775
rect 2499 1771 2500 1775
rect 2494 1770 2500 1771
rect 2686 1775 2692 1776
rect 2686 1771 2687 1775
rect 2691 1771 2692 1775
rect 2686 1770 2692 1771
rect 2878 1775 2884 1776
rect 2878 1771 2879 1775
rect 2883 1771 2884 1775
rect 2878 1770 2884 1771
rect 3070 1775 3076 1776
rect 3070 1771 3071 1775
rect 3075 1771 3076 1775
rect 3070 1770 3076 1771
rect 3262 1775 3268 1776
rect 3262 1771 3263 1775
rect 3267 1771 3268 1775
rect 3262 1770 3268 1771
rect 3462 1775 3468 1776
rect 3462 1771 3463 1775
rect 3467 1771 3468 1775
rect 3462 1770 3468 1771
rect 3662 1775 3668 1776
rect 3662 1771 3663 1775
rect 3667 1771 3668 1775
rect 3662 1770 3668 1771
rect 3838 1775 3844 1776
rect 3838 1771 3839 1775
rect 3843 1771 3844 1775
rect 3942 1772 3943 1776
rect 3947 1772 3948 1776
rect 3942 1771 3948 1772
rect 3838 1770 3844 1771
rect 2046 1759 2052 1760
rect 2006 1756 2012 1757
rect 110 1752 111 1756
rect 115 1752 116 1756
rect 110 1751 116 1752
rect 254 1755 260 1756
rect 254 1751 255 1755
rect 259 1751 260 1755
rect 254 1750 260 1751
rect 390 1755 396 1756
rect 390 1751 391 1755
rect 395 1751 396 1755
rect 390 1750 396 1751
rect 534 1755 540 1756
rect 534 1751 535 1755
rect 539 1751 540 1755
rect 534 1750 540 1751
rect 694 1755 700 1756
rect 694 1751 695 1755
rect 699 1751 700 1755
rect 694 1750 700 1751
rect 862 1755 868 1756
rect 862 1751 863 1755
rect 867 1751 868 1755
rect 862 1750 868 1751
rect 1030 1755 1036 1756
rect 1030 1751 1031 1755
rect 1035 1751 1036 1755
rect 1030 1750 1036 1751
rect 1206 1755 1212 1756
rect 1206 1751 1207 1755
rect 1211 1751 1212 1755
rect 1206 1750 1212 1751
rect 1382 1755 1388 1756
rect 1382 1751 1383 1755
rect 1387 1751 1388 1755
rect 1382 1750 1388 1751
rect 1558 1755 1564 1756
rect 1558 1751 1559 1755
rect 1563 1751 1564 1755
rect 1558 1750 1564 1751
rect 1742 1755 1748 1756
rect 1742 1751 1743 1755
rect 1747 1751 1748 1755
rect 2006 1752 2007 1756
rect 2011 1752 2012 1756
rect 2046 1755 2047 1759
rect 2051 1755 2052 1759
rect 3942 1759 3948 1760
rect 2046 1754 2052 1755
rect 2126 1756 2132 1757
rect 2006 1751 2012 1752
rect 1742 1750 1748 1751
rect 110 1739 116 1740
rect 110 1735 111 1739
rect 115 1735 116 1739
rect 2006 1739 2012 1740
rect 110 1734 116 1735
rect 254 1736 260 1737
rect 112 1707 114 1734
rect 254 1732 255 1736
rect 259 1732 260 1736
rect 254 1731 260 1732
rect 390 1736 396 1737
rect 390 1732 391 1736
rect 395 1732 396 1736
rect 390 1731 396 1732
rect 534 1736 540 1737
rect 534 1732 535 1736
rect 539 1732 540 1736
rect 534 1731 540 1732
rect 694 1736 700 1737
rect 694 1732 695 1736
rect 699 1732 700 1736
rect 694 1731 700 1732
rect 862 1736 868 1737
rect 862 1732 863 1736
rect 867 1732 868 1736
rect 862 1731 868 1732
rect 1030 1736 1036 1737
rect 1030 1732 1031 1736
rect 1035 1732 1036 1736
rect 1030 1731 1036 1732
rect 1206 1736 1212 1737
rect 1206 1732 1207 1736
rect 1211 1732 1212 1736
rect 1206 1731 1212 1732
rect 1382 1736 1388 1737
rect 1382 1732 1383 1736
rect 1387 1732 1388 1736
rect 1382 1731 1388 1732
rect 1558 1736 1564 1737
rect 1558 1732 1559 1736
rect 1563 1732 1564 1736
rect 1558 1731 1564 1732
rect 1742 1736 1748 1737
rect 1742 1732 1743 1736
rect 1747 1732 1748 1736
rect 2006 1735 2007 1739
rect 2011 1735 2012 1739
rect 2006 1734 2012 1735
rect 1742 1731 1748 1732
rect 256 1707 258 1731
rect 392 1707 394 1731
rect 536 1707 538 1731
rect 696 1707 698 1731
rect 864 1707 866 1731
rect 1032 1707 1034 1731
rect 1208 1707 1210 1731
rect 1384 1707 1386 1731
rect 1560 1707 1562 1731
rect 1744 1707 1746 1731
rect 2008 1707 2010 1734
rect 2048 1723 2050 1754
rect 2126 1752 2127 1756
rect 2131 1752 2132 1756
rect 2126 1751 2132 1752
rect 2310 1756 2316 1757
rect 2310 1752 2311 1756
rect 2315 1752 2316 1756
rect 2310 1751 2316 1752
rect 2494 1756 2500 1757
rect 2494 1752 2495 1756
rect 2499 1752 2500 1756
rect 2494 1751 2500 1752
rect 2686 1756 2692 1757
rect 2686 1752 2687 1756
rect 2691 1752 2692 1756
rect 2686 1751 2692 1752
rect 2878 1756 2884 1757
rect 2878 1752 2879 1756
rect 2883 1752 2884 1756
rect 2878 1751 2884 1752
rect 3070 1756 3076 1757
rect 3070 1752 3071 1756
rect 3075 1752 3076 1756
rect 3070 1751 3076 1752
rect 3262 1756 3268 1757
rect 3262 1752 3263 1756
rect 3267 1752 3268 1756
rect 3262 1751 3268 1752
rect 3462 1756 3468 1757
rect 3462 1752 3463 1756
rect 3467 1752 3468 1756
rect 3462 1751 3468 1752
rect 3662 1756 3668 1757
rect 3662 1752 3663 1756
rect 3667 1752 3668 1756
rect 3662 1751 3668 1752
rect 3838 1756 3844 1757
rect 3838 1752 3839 1756
rect 3843 1752 3844 1756
rect 3942 1755 3943 1759
rect 3947 1755 3948 1759
rect 3942 1754 3948 1755
rect 3838 1751 3844 1752
rect 2128 1723 2130 1751
rect 2312 1723 2314 1751
rect 2496 1723 2498 1751
rect 2688 1723 2690 1751
rect 2880 1723 2882 1751
rect 3072 1723 3074 1751
rect 3264 1723 3266 1751
rect 3464 1723 3466 1751
rect 3664 1723 3666 1751
rect 3840 1723 3842 1751
rect 3944 1723 3946 1754
rect 2047 1722 2051 1723
rect 2047 1717 2051 1718
rect 2071 1722 2075 1723
rect 2071 1717 2075 1718
rect 2127 1722 2131 1723
rect 2127 1717 2131 1718
rect 2191 1722 2195 1723
rect 2191 1717 2195 1718
rect 2311 1722 2315 1723
rect 2311 1717 2315 1718
rect 2343 1722 2347 1723
rect 2343 1717 2347 1718
rect 2495 1722 2499 1723
rect 2495 1717 2499 1718
rect 2511 1722 2515 1723
rect 2511 1717 2515 1718
rect 2687 1722 2691 1723
rect 2687 1717 2691 1718
rect 2871 1722 2875 1723
rect 2871 1717 2875 1718
rect 2879 1722 2883 1723
rect 2879 1717 2883 1718
rect 3063 1722 3067 1723
rect 3063 1717 3067 1718
rect 3071 1722 3075 1723
rect 3071 1717 3075 1718
rect 3255 1722 3259 1723
rect 3255 1717 3259 1718
rect 3263 1722 3267 1723
rect 3263 1717 3267 1718
rect 3447 1722 3451 1723
rect 3447 1717 3451 1718
rect 3463 1722 3467 1723
rect 3463 1717 3467 1718
rect 3647 1722 3651 1723
rect 3647 1717 3651 1718
rect 3663 1722 3667 1723
rect 3663 1717 3667 1718
rect 3839 1722 3843 1723
rect 3839 1717 3843 1718
rect 3943 1722 3947 1723
rect 3943 1717 3947 1718
rect 111 1706 115 1707
rect 111 1701 115 1702
rect 135 1706 139 1707
rect 135 1701 139 1702
rect 255 1706 259 1707
rect 255 1701 259 1702
rect 263 1706 267 1707
rect 263 1701 267 1702
rect 391 1706 395 1707
rect 391 1701 395 1702
rect 431 1706 435 1707
rect 431 1701 435 1702
rect 535 1706 539 1707
rect 535 1701 539 1702
rect 607 1706 611 1707
rect 607 1701 611 1702
rect 695 1706 699 1707
rect 695 1701 699 1702
rect 799 1706 803 1707
rect 799 1701 803 1702
rect 863 1706 867 1707
rect 863 1701 867 1702
rect 999 1706 1003 1707
rect 999 1701 1003 1702
rect 1031 1706 1035 1707
rect 1031 1701 1035 1702
rect 1199 1706 1203 1707
rect 1199 1701 1203 1702
rect 1207 1706 1211 1707
rect 1207 1701 1211 1702
rect 1383 1706 1387 1707
rect 1383 1701 1387 1702
rect 1407 1706 1411 1707
rect 1407 1701 1411 1702
rect 1559 1706 1563 1707
rect 1559 1701 1563 1702
rect 1623 1706 1627 1707
rect 1623 1701 1627 1702
rect 1743 1706 1747 1707
rect 1743 1701 1747 1702
rect 1839 1706 1843 1707
rect 1839 1701 1843 1702
rect 2007 1706 2011 1707
rect 2007 1701 2011 1702
rect 112 1674 114 1701
rect 136 1677 138 1701
rect 264 1677 266 1701
rect 432 1677 434 1701
rect 608 1677 610 1701
rect 800 1677 802 1701
rect 1000 1677 1002 1701
rect 1200 1677 1202 1701
rect 1408 1677 1410 1701
rect 1624 1677 1626 1701
rect 1840 1677 1842 1701
rect 134 1676 140 1677
rect 110 1673 116 1674
rect 110 1669 111 1673
rect 115 1669 116 1673
rect 134 1672 135 1676
rect 139 1672 140 1676
rect 134 1671 140 1672
rect 262 1676 268 1677
rect 262 1672 263 1676
rect 267 1672 268 1676
rect 262 1671 268 1672
rect 430 1676 436 1677
rect 430 1672 431 1676
rect 435 1672 436 1676
rect 430 1671 436 1672
rect 606 1676 612 1677
rect 606 1672 607 1676
rect 611 1672 612 1676
rect 606 1671 612 1672
rect 798 1676 804 1677
rect 798 1672 799 1676
rect 803 1672 804 1676
rect 798 1671 804 1672
rect 998 1676 1004 1677
rect 998 1672 999 1676
rect 1003 1672 1004 1676
rect 998 1671 1004 1672
rect 1198 1676 1204 1677
rect 1198 1672 1199 1676
rect 1203 1672 1204 1676
rect 1198 1671 1204 1672
rect 1406 1676 1412 1677
rect 1406 1672 1407 1676
rect 1411 1672 1412 1676
rect 1406 1671 1412 1672
rect 1622 1676 1628 1677
rect 1622 1672 1623 1676
rect 1627 1672 1628 1676
rect 1622 1671 1628 1672
rect 1838 1676 1844 1677
rect 1838 1672 1839 1676
rect 1843 1672 1844 1676
rect 2008 1674 2010 1701
rect 2048 1690 2050 1717
rect 2072 1693 2074 1717
rect 2192 1693 2194 1717
rect 2344 1693 2346 1717
rect 2512 1693 2514 1717
rect 2688 1693 2690 1717
rect 2872 1693 2874 1717
rect 3064 1693 3066 1717
rect 3256 1693 3258 1717
rect 3448 1693 3450 1717
rect 3648 1693 3650 1717
rect 3840 1693 3842 1717
rect 2070 1692 2076 1693
rect 2046 1689 2052 1690
rect 2046 1685 2047 1689
rect 2051 1685 2052 1689
rect 2070 1688 2071 1692
rect 2075 1688 2076 1692
rect 2070 1687 2076 1688
rect 2190 1692 2196 1693
rect 2190 1688 2191 1692
rect 2195 1688 2196 1692
rect 2190 1687 2196 1688
rect 2342 1692 2348 1693
rect 2342 1688 2343 1692
rect 2347 1688 2348 1692
rect 2342 1687 2348 1688
rect 2510 1692 2516 1693
rect 2510 1688 2511 1692
rect 2515 1688 2516 1692
rect 2510 1687 2516 1688
rect 2686 1692 2692 1693
rect 2686 1688 2687 1692
rect 2691 1688 2692 1692
rect 2686 1687 2692 1688
rect 2870 1692 2876 1693
rect 2870 1688 2871 1692
rect 2875 1688 2876 1692
rect 2870 1687 2876 1688
rect 3062 1692 3068 1693
rect 3062 1688 3063 1692
rect 3067 1688 3068 1692
rect 3062 1687 3068 1688
rect 3254 1692 3260 1693
rect 3254 1688 3255 1692
rect 3259 1688 3260 1692
rect 3254 1687 3260 1688
rect 3446 1692 3452 1693
rect 3446 1688 3447 1692
rect 3451 1688 3452 1692
rect 3446 1687 3452 1688
rect 3646 1692 3652 1693
rect 3646 1688 3647 1692
rect 3651 1688 3652 1692
rect 3646 1687 3652 1688
rect 3838 1692 3844 1693
rect 3838 1688 3839 1692
rect 3843 1688 3844 1692
rect 3944 1690 3946 1717
rect 3838 1687 3844 1688
rect 3942 1689 3948 1690
rect 2046 1684 2052 1685
rect 3942 1685 3943 1689
rect 3947 1685 3948 1689
rect 3942 1684 3948 1685
rect 1838 1671 1844 1672
rect 2006 1673 2012 1674
rect 2070 1673 2076 1674
rect 110 1668 116 1669
rect 2006 1669 2007 1673
rect 2011 1669 2012 1673
rect 2006 1668 2012 1669
rect 2046 1672 2052 1673
rect 2046 1668 2047 1672
rect 2051 1668 2052 1672
rect 2070 1669 2071 1673
rect 2075 1669 2076 1673
rect 2070 1668 2076 1669
rect 2190 1673 2196 1674
rect 2190 1669 2191 1673
rect 2195 1669 2196 1673
rect 2190 1668 2196 1669
rect 2342 1673 2348 1674
rect 2342 1669 2343 1673
rect 2347 1669 2348 1673
rect 2342 1668 2348 1669
rect 2510 1673 2516 1674
rect 2510 1669 2511 1673
rect 2515 1669 2516 1673
rect 2510 1668 2516 1669
rect 2686 1673 2692 1674
rect 2686 1669 2687 1673
rect 2691 1669 2692 1673
rect 2686 1668 2692 1669
rect 2870 1673 2876 1674
rect 2870 1669 2871 1673
rect 2875 1669 2876 1673
rect 2870 1668 2876 1669
rect 3062 1673 3068 1674
rect 3062 1669 3063 1673
rect 3067 1669 3068 1673
rect 3062 1668 3068 1669
rect 3254 1673 3260 1674
rect 3254 1669 3255 1673
rect 3259 1669 3260 1673
rect 3254 1668 3260 1669
rect 3446 1673 3452 1674
rect 3446 1669 3447 1673
rect 3451 1669 3452 1673
rect 3446 1668 3452 1669
rect 3646 1673 3652 1674
rect 3646 1669 3647 1673
rect 3651 1669 3652 1673
rect 3646 1668 3652 1669
rect 3838 1673 3844 1674
rect 3838 1669 3839 1673
rect 3843 1669 3844 1673
rect 3838 1668 3844 1669
rect 3942 1672 3948 1673
rect 3942 1668 3943 1672
rect 3947 1668 3948 1672
rect 2046 1667 2052 1668
rect 134 1657 140 1658
rect 110 1656 116 1657
rect 110 1652 111 1656
rect 115 1652 116 1656
rect 134 1653 135 1657
rect 139 1653 140 1657
rect 134 1652 140 1653
rect 262 1657 268 1658
rect 262 1653 263 1657
rect 267 1653 268 1657
rect 262 1652 268 1653
rect 430 1657 436 1658
rect 430 1653 431 1657
rect 435 1653 436 1657
rect 430 1652 436 1653
rect 606 1657 612 1658
rect 606 1653 607 1657
rect 611 1653 612 1657
rect 606 1652 612 1653
rect 798 1657 804 1658
rect 798 1653 799 1657
rect 803 1653 804 1657
rect 798 1652 804 1653
rect 998 1657 1004 1658
rect 998 1653 999 1657
rect 1003 1653 1004 1657
rect 998 1652 1004 1653
rect 1198 1657 1204 1658
rect 1198 1653 1199 1657
rect 1203 1653 1204 1657
rect 1198 1652 1204 1653
rect 1406 1657 1412 1658
rect 1406 1653 1407 1657
rect 1411 1653 1412 1657
rect 1406 1652 1412 1653
rect 1622 1657 1628 1658
rect 1622 1653 1623 1657
rect 1627 1653 1628 1657
rect 1622 1652 1628 1653
rect 1838 1657 1844 1658
rect 1838 1653 1839 1657
rect 1843 1653 1844 1657
rect 1838 1652 1844 1653
rect 2006 1656 2012 1657
rect 2006 1652 2007 1656
rect 2011 1652 2012 1656
rect 110 1651 116 1652
rect 112 1631 114 1651
rect 136 1631 138 1652
rect 264 1631 266 1652
rect 432 1631 434 1652
rect 608 1631 610 1652
rect 800 1631 802 1652
rect 1000 1631 1002 1652
rect 1200 1631 1202 1652
rect 1408 1631 1410 1652
rect 1624 1631 1626 1652
rect 1840 1631 1842 1652
rect 2006 1651 2012 1652
rect 2008 1631 2010 1651
rect 2048 1647 2050 1667
rect 2072 1647 2074 1668
rect 2192 1647 2194 1668
rect 2344 1647 2346 1668
rect 2512 1647 2514 1668
rect 2688 1647 2690 1668
rect 2872 1647 2874 1668
rect 3064 1647 3066 1668
rect 3256 1647 3258 1668
rect 3448 1647 3450 1668
rect 3648 1647 3650 1668
rect 3840 1647 3842 1668
rect 3942 1667 3948 1668
rect 3944 1647 3946 1667
rect 2047 1646 2051 1647
rect 2047 1641 2051 1642
rect 2071 1646 2075 1647
rect 2071 1641 2075 1642
rect 2191 1646 2195 1647
rect 2191 1641 2195 1642
rect 2335 1646 2339 1647
rect 2335 1641 2339 1642
rect 2343 1646 2347 1647
rect 2343 1641 2347 1642
rect 2511 1646 2515 1647
rect 2511 1641 2515 1642
rect 2599 1646 2603 1647
rect 2599 1641 2603 1642
rect 2687 1646 2691 1647
rect 2687 1641 2691 1642
rect 2839 1646 2843 1647
rect 2839 1641 2843 1642
rect 2871 1646 2875 1647
rect 2871 1641 2875 1642
rect 3047 1646 3051 1647
rect 3047 1641 3051 1642
rect 3063 1646 3067 1647
rect 3063 1641 3067 1642
rect 3231 1646 3235 1647
rect 3231 1641 3235 1642
rect 3255 1646 3259 1647
rect 3255 1641 3259 1642
rect 3399 1646 3403 1647
rect 3399 1641 3403 1642
rect 3447 1646 3451 1647
rect 3447 1641 3451 1642
rect 3551 1646 3555 1647
rect 3551 1641 3555 1642
rect 3647 1646 3651 1647
rect 3647 1641 3651 1642
rect 3695 1646 3699 1647
rect 3695 1641 3699 1642
rect 3839 1646 3843 1647
rect 3839 1641 3843 1642
rect 3943 1646 3947 1647
rect 3943 1641 3947 1642
rect 111 1630 115 1631
rect 111 1625 115 1626
rect 135 1630 139 1631
rect 135 1625 139 1626
rect 263 1630 267 1631
rect 263 1625 267 1626
rect 287 1630 291 1631
rect 287 1625 291 1626
rect 431 1630 435 1631
rect 431 1625 435 1626
rect 471 1630 475 1631
rect 471 1625 475 1626
rect 607 1630 611 1631
rect 607 1625 611 1626
rect 655 1630 659 1631
rect 655 1625 659 1626
rect 799 1630 803 1631
rect 799 1625 803 1626
rect 839 1630 843 1631
rect 839 1625 843 1626
rect 999 1630 1003 1631
rect 999 1625 1003 1626
rect 1015 1630 1019 1631
rect 1015 1625 1019 1626
rect 1183 1630 1187 1631
rect 1183 1625 1187 1626
rect 1199 1630 1203 1631
rect 1199 1625 1203 1626
rect 1343 1630 1347 1631
rect 1343 1625 1347 1626
rect 1407 1630 1411 1631
rect 1407 1625 1411 1626
rect 1495 1630 1499 1631
rect 1495 1625 1499 1626
rect 1623 1630 1627 1631
rect 1623 1625 1627 1626
rect 1639 1630 1643 1631
rect 1639 1625 1643 1626
rect 1783 1630 1787 1631
rect 1783 1625 1787 1626
rect 1839 1630 1843 1631
rect 1839 1625 1843 1626
rect 1903 1630 1907 1631
rect 1903 1625 1907 1626
rect 2007 1630 2011 1631
rect 2007 1625 2011 1626
rect 112 1605 114 1625
rect 110 1604 116 1605
rect 136 1604 138 1625
rect 288 1604 290 1625
rect 472 1604 474 1625
rect 656 1604 658 1625
rect 840 1604 842 1625
rect 1016 1604 1018 1625
rect 1184 1604 1186 1625
rect 1344 1604 1346 1625
rect 1496 1604 1498 1625
rect 1640 1604 1642 1625
rect 1784 1604 1786 1625
rect 1904 1604 1906 1625
rect 2008 1605 2010 1625
rect 2048 1621 2050 1641
rect 2046 1620 2052 1621
rect 2072 1620 2074 1641
rect 2336 1620 2338 1641
rect 2600 1620 2602 1641
rect 2840 1620 2842 1641
rect 3048 1620 3050 1641
rect 3232 1620 3234 1641
rect 3400 1620 3402 1641
rect 3552 1620 3554 1641
rect 3696 1620 3698 1641
rect 3840 1620 3842 1641
rect 3944 1621 3946 1641
rect 3942 1620 3948 1621
rect 2046 1616 2047 1620
rect 2051 1616 2052 1620
rect 2046 1615 2052 1616
rect 2070 1619 2076 1620
rect 2070 1615 2071 1619
rect 2075 1615 2076 1619
rect 2070 1614 2076 1615
rect 2334 1619 2340 1620
rect 2334 1615 2335 1619
rect 2339 1615 2340 1619
rect 2334 1614 2340 1615
rect 2598 1619 2604 1620
rect 2598 1615 2599 1619
rect 2603 1615 2604 1619
rect 2598 1614 2604 1615
rect 2838 1619 2844 1620
rect 2838 1615 2839 1619
rect 2843 1615 2844 1619
rect 2838 1614 2844 1615
rect 3046 1619 3052 1620
rect 3046 1615 3047 1619
rect 3051 1615 3052 1619
rect 3046 1614 3052 1615
rect 3230 1619 3236 1620
rect 3230 1615 3231 1619
rect 3235 1615 3236 1619
rect 3230 1614 3236 1615
rect 3398 1619 3404 1620
rect 3398 1615 3399 1619
rect 3403 1615 3404 1619
rect 3398 1614 3404 1615
rect 3550 1619 3556 1620
rect 3550 1615 3551 1619
rect 3555 1615 3556 1619
rect 3550 1614 3556 1615
rect 3694 1619 3700 1620
rect 3694 1615 3695 1619
rect 3699 1615 3700 1619
rect 3694 1614 3700 1615
rect 3838 1619 3844 1620
rect 3838 1615 3839 1619
rect 3843 1615 3844 1619
rect 3942 1616 3943 1620
rect 3947 1616 3948 1620
rect 3942 1615 3948 1616
rect 3838 1614 3844 1615
rect 2006 1604 2012 1605
rect 110 1600 111 1604
rect 115 1600 116 1604
rect 110 1599 116 1600
rect 134 1603 140 1604
rect 134 1599 135 1603
rect 139 1599 140 1603
rect 134 1598 140 1599
rect 286 1603 292 1604
rect 286 1599 287 1603
rect 291 1599 292 1603
rect 286 1598 292 1599
rect 470 1603 476 1604
rect 470 1599 471 1603
rect 475 1599 476 1603
rect 470 1598 476 1599
rect 654 1603 660 1604
rect 654 1599 655 1603
rect 659 1599 660 1603
rect 654 1598 660 1599
rect 838 1603 844 1604
rect 838 1599 839 1603
rect 843 1599 844 1603
rect 838 1598 844 1599
rect 1014 1603 1020 1604
rect 1014 1599 1015 1603
rect 1019 1599 1020 1603
rect 1014 1598 1020 1599
rect 1182 1603 1188 1604
rect 1182 1599 1183 1603
rect 1187 1599 1188 1603
rect 1182 1598 1188 1599
rect 1342 1603 1348 1604
rect 1342 1599 1343 1603
rect 1347 1599 1348 1603
rect 1342 1598 1348 1599
rect 1494 1603 1500 1604
rect 1494 1599 1495 1603
rect 1499 1599 1500 1603
rect 1494 1598 1500 1599
rect 1638 1603 1644 1604
rect 1638 1599 1639 1603
rect 1643 1599 1644 1603
rect 1638 1598 1644 1599
rect 1782 1603 1788 1604
rect 1782 1599 1783 1603
rect 1787 1599 1788 1603
rect 1782 1598 1788 1599
rect 1902 1603 1908 1604
rect 1902 1599 1903 1603
rect 1907 1599 1908 1603
rect 2006 1600 2007 1604
rect 2011 1600 2012 1604
rect 2006 1599 2012 1600
rect 2046 1603 2052 1604
rect 2046 1599 2047 1603
rect 2051 1599 2052 1603
rect 3942 1603 3948 1604
rect 1902 1598 1908 1599
rect 2046 1598 2052 1599
rect 2070 1600 2076 1601
rect 110 1587 116 1588
rect 110 1583 111 1587
rect 115 1583 116 1587
rect 2006 1587 2012 1588
rect 110 1582 116 1583
rect 134 1584 140 1585
rect 112 1551 114 1582
rect 134 1580 135 1584
rect 139 1580 140 1584
rect 134 1579 140 1580
rect 286 1584 292 1585
rect 286 1580 287 1584
rect 291 1580 292 1584
rect 286 1579 292 1580
rect 470 1584 476 1585
rect 470 1580 471 1584
rect 475 1580 476 1584
rect 470 1579 476 1580
rect 654 1584 660 1585
rect 654 1580 655 1584
rect 659 1580 660 1584
rect 654 1579 660 1580
rect 838 1584 844 1585
rect 838 1580 839 1584
rect 843 1580 844 1584
rect 838 1579 844 1580
rect 1014 1584 1020 1585
rect 1014 1580 1015 1584
rect 1019 1580 1020 1584
rect 1014 1579 1020 1580
rect 1182 1584 1188 1585
rect 1182 1580 1183 1584
rect 1187 1580 1188 1584
rect 1182 1579 1188 1580
rect 1342 1584 1348 1585
rect 1342 1580 1343 1584
rect 1347 1580 1348 1584
rect 1342 1579 1348 1580
rect 1494 1584 1500 1585
rect 1494 1580 1495 1584
rect 1499 1580 1500 1584
rect 1494 1579 1500 1580
rect 1638 1584 1644 1585
rect 1638 1580 1639 1584
rect 1643 1580 1644 1584
rect 1638 1579 1644 1580
rect 1782 1584 1788 1585
rect 1782 1580 1783 1584
rect 1787 1580 1788 1584
rect 1782 1579 1788 1580
rect 1902 1584 1908 1585
rect 1902 1580 1903 1584
rect 1907 1580 1908 1584
rect 2006 1583 2007 1587
rect 2011 1583 2012 1587
rect 2006 1582 2012 1583
rect 1902 1579 1908 1580
rect 136 1551 138 1579
rect 288 1551 290 1579
rect 472 1551 474 1579
rect 656 1551 658 1579
rect 840 1551 842 1579
rect 1016 1551 1018 1579
rect 1184 1551 1186 1579
rect 1344 1551 1346 1579
rect 1496 1551 1498 1579
rect 1640 1551 1642 1579
rect 1784 1551 1786 1579
rect 1904 1551 1906 1579
rect 2008 1551 2010 1582
rect 2048 1567 2050 1598
rect 2070 1596 2071 1600
rect 2075 1596 2076 1600
rect 2070 1595 2076 1596
rect 2334 1600 2340 1601
rect 2334 1596 2335 1600
rect 2339 1596 2340 1600
rect 2334 1595 2340 1596
rect 2598 1600 2604 1601
rect 2598 1596 2599 1600
rect 2603 1596 2604 1600
rect 2598 1595 2604 1596
rect 2838 1600 2844 1601
rect 2838 1596 2839 1600
rect 2843 1596 2844 1600
rect 2838 1595 2844 1596
rect 3046 1600 3052 1601
rect 3046 1596 3047 1600
rect 3051 1596 3052 1600
rect 3046 1595 3052 1596
rect 3230 1600 3236 1601
rect 3230 1596 3231 1600
rect 3235 1596 3236 1600
rect 3230 1595 3236 1596
rect 3398 1600 3404 1601
rect 3398 1596 3399 1600
rect 3403 1596 3404 1600
rect 3398 1595 3404 1596
rect 3550 1600 3556 1601
rect 3550 1596 3551 1600
rect 3555 1596 3556 1600
rect 3550 1595 3556 1596
rect 3694 1600 3700 1601
rect 3694 1596 3695 1600
rect 3699 1596 3700 1600
rect 3694 1595 3700 1596
rect 3838 1600 3844 1601
rect 3838 1596 3839 1600
rect 3843 1596 3844 1600
rect 3942 1599 3943 1603
rect 3947 1599 3948 1603
rect 3942 1598 3948 1599
rect 3838 1595 3844 1596
rect 2072 1567 2074 1595
rect 2336 1567 2338 1595
rect 2600 1567 2602 1595
rect 2840 1567 2842 1595
rect 3048 1567 3050 1595
rect 3232 1567 3234 1595
rect 3400 1567 3402 1595
rect 3552 1567 3554 1595
rect 3696 1567 3698 1595
rect 3840 1567 3842 1595
rect 3944 1567 3946 1598
rect 2047 1566 2051 1567
rect 2047 1561 2051 1562
rect 2071 1566 2075 1567
rect 2071 1561 2075 1562
rect 2335 1566 2339 1567
rect 2335 1561 2339 1562
rect 2583 1566 2587 1567
rect 2583 1561 2587 1562
rect 2599 1566 2603 1567
rect 2599 1561 2603 1562
rect 2743 1566 2747 1567
rect 2743 1561 2747 1562
rect 2839 1566 2843 1567
rect 2839 1561 2843 1562
rect 2903 1566 2907 1567
rect 2903 1561 2907 1562
rect 3047 1566 3051 1567
rect 3047 1561 3051 1562
rect 3063 1566 3067 1567
rect 3063 1561 3067 1562
rect 3223 1566 3227 1567
rect 3223 1561 3227 1562
rect 3231 1566 3235 1567
rect 3231 1561 3235 1562
rect 3383 1566 3387 1567
rect 3383 1561 3387 1562
rect 3399 1566 3403 1567
rect 3399 1561 3403 1562
rect 3543 1566 3547 1567
rect 3543 1561 3547 1562
rect 3551 1566 3555 1567
rect 3551 1561 3555 1562
rect 3695 1566 3699 1567
rect 3695 1561 3699 1562
rect 3703 1566 3707 1567
rect 3703 1561 3707 1562
rect 3839 1566 3843 1567
rect 3839 1561 3843 1562
rect 3943 1566 3947 1567
rect 3943 1561 3947 1562
rect 111 1550 115 1551
rect 111 1545 115 1546
rect 135 1550 139 1551
rect 135 1545 139 1546
rect 287 1550 291 1551
rect 287 1545 291 1546
rect 295 1550 299 1551
rect 295 1545 299 1546
rect 471 1550 475 1551
rect 471 1545 475 1546
rect 487 1550 491 1551
rect 487 1545 491 1546
rect 655 1550 659 1551
rect 655 1545 659 1546
rect 687 1550 691 1551
rect 687 1545 691 1546
rect 839 1550 843 1551
rect 839 1545 843 1546
rect 887 1550 891 1551
rect 887 1545 891 1546
rect 1015 1550 1019 1551
rect 1015 1545 1019 1546
rect 1079 1550 1083 1551
rect 1079 1545 1083 1546
rect 1183 1550 1187 1551
rect 1183 1545 1187 1546
rect 1263 1550 1267 1551
rect 1263 1545 1267 1546
rect 1343 1550 1347 1551
rect 1343 1545 1347 1546
rect 1447 1550 1451 1551
rect 1447 1545 1451 1546
rect 1495 1550 1499 1551
rect 1495 1545 1499 1546
rect 1623 1550 1627 1551
rect 1623 1545 1627 1546
rect 1639 1550 1643 1551
rect 1639 1545 1643 1546
rect 1783 1550 1787 1551
rect 1783 1545 1787 1546
rect 1807 1550 1811 1551
rect 1807 1545 1811 1546
rect 1903 1550 1907 1551
rect 1903 1545 1907 1546
rect 2007 1550 2011 1551
rect 2007 1545 2011 1546
rect 112 1518 114 1545
rect 136 1521 138 1545
rect 296 1521 298 1545
rect 488 1521 490 1545
rect 688 1521 690 1545
rect 888 1521 890 1545
rect 1080 1521 1082 1545
rect 1264 1521 1266 1545
rect 1448 1521 1450 1545
rect 1624 1521 1626 1545
rect 1808 1521 1810 1545
rect 134 1520 140 1521
rect 110 1517 116 1518
rect 110 1513 111 1517
rect 115 1513 116 1517
rect 134 1516 135 1520
rect 139 1516 140 1520
rect 134 1515 140 1516
rect 294 1520 300 1521
rect 294 1516 295 1520
rect 299 1516 300 1520
rect 294 1515 300 1516
rect 486 1520 492 1521
rect 486 1516 487 1520
rect 491 1516 492 1520
rect 486 1515 492 1516
rect 686 1520 692 1521
rect 686 1516 687 1520
rect 691 1516 692 1520
rect 686 1515 692 1516
rect 886 1520 892 1521
rect 886 1516 887 1520
rect 891 1516 892 1520
rect 886 1515 892 1516
rect 1078 1520 1084 1521
rect 1078 1516 1079 1520
rect 1083 1516 1084 1520
rect 1078 1515 1084 1516
rect 1262 1520 1268 1521
rect 1262 1516 1263 1520
rect 1267 1516 1268 1520
rect 1262 1515 1268 1516
rect 1446 1520 1452 1521
rect 1446 1516 1447 1520
rect 1451 1516 1452 1520
rect 1446 1515 1452 1516
rect 1622 1520 1628 1521
rect 1622 1516 1623 1520
rect 1627 1516 1628 1520
rect 1622 1515 1628 1516
rect 1806 1520 1812 1521
rect 1806 1516 1807 1520
rect 1811 1516 1812 1520
rect 2008 1518 2010 1545
rect 2048 1534 2050 1561
rect 2584 1537 2586 1561
rect 2744 1537 2746 1561
rect 2904 1537 2906 1561
rect 3064 1537 3066 1561
rect 3224 1537 3226 1561
rect 3384 1537 3386 1561
rect 3544 1537 3546 1561
rect 3704 1537 3706 1561
rect 2582 1536 2588 1537
rect 2046 1533 2052 1534
rect 2046 1529 2047 1533
rect 2051 1529 2052 1533
rect 2582 1532 2583 1536
rect 2587 1532 2588 1536
rect 2582 1531 2588 1532
rect 2742 1536 2748 1537
rect 2742 1532 2743 1536
rect 2747 1532 2748 1536
rect 2742 1531 2748 1532
rect 2902 1536 2908 1537
rect 2902 1532 2903 1536
rect 2907 1532 2908 1536
rect 2902 1531 2908 1532
rect 3062 1536 3068 1537
rect 3062 1532 3063 1536
rect 3067 1532 3068 1536
rect 3062 1531 3068 1532
rect 3222 1536 3228 1537
rect 3222 1532 3223 1536
rect 3227 1532 3228 1536
rect 3222 1531 3228 1532
rect 3382 1536 3388 1537
rect 3382 1532 3383 1536
rect 3387 1532 3388 1536
rect 3382 1531 3388 1532
rect 3542 1536 3548 1537
rect 3542 1532 3543 1536
rect 3547 1532 3548 1536
rect 3542 1531 3548 1532
rect 3702 1536 3708 1537
rect 3702 1532 3703 1536
rect 3707 1532 3708 1536
rect 3944 1534 3946 1561
rect 3702 1531 3708 1532
rect 3942 1533 3948 1534
rect 2046 1528 2052 1529
rect 3942 1529 3943 1533
rect 3947 1529 3948 1533
rect 3942 1528 3948 1529
rect 1806 1515 1812 1516
rect 2006 1517 2012 1518
rect 2582 1517 2588 1518
rect 110 1512 116 1513
rect 2006 1513 2007 1517
rect 2011 1513 2012 1517
rect 2006 1512 2012 1513
rect 2046 1516 2052 1517
rect 2046 1512 2047 1516
rect 2051 1512 2052 1516
rect 2582 1513 2583 1517
rect 2587 1513 2588 1517
rect 2582 1512 2588 1513
rect 2742 1517 2748 1518
rect 2742 1513 2743 1517
rect 2747 1513 2748 1517
rect 2742 1512 2748 1513
rect 2902 1517 2908 1518
rect 2902 1513 2903 1517
rect 2907 1513 2908 1517
rect 2902 1512 2908 1513
rect 3062 1517 3068 1518
rect 3062 1513 3063 1517
rect 3067 1513 3068 1517
rect 3062 1512 3068 1513
rect 3222 1517 3228 1518
rect 3222 1513 3223 1517
rect 3227 1513 3228 1517
rect 3222 1512 3228 1513
rect 3382 1517 3388 1518
rect 3382 1513 3383 1517
rect 3387 1513 3388 1517
rect 3382 1512 3388 1513
rect 3542 1517 3548 1518
rect 3542 1513 3543 1517
rect 3547 1513 3548 1517
rect 3542 1512 3548 1513
rect 3702 1517 3708 1518
rect 3702 1513 3703 1517
rect 3707 1513 3708 1517
rect 3702 1512 3708 1513
rect 3942 1516 3948 1517
rect 3942 1512 3943 1516
rect 3947 1512 3948 1516
rect 2046 1511 2052 1512
rect 134 1501 140 1502
rect 110 1500 116 1501
rect 110 1496 111 1500
rect 115 1496 116 1500
rect 134 1497 135 1501
rect 139 1497 140 1501
rect 134 1496 140 1497
rect 294 1501 300 1502
rect 294 1497 295 1501
rect 299 1497 300 1501
rect 294 1496 300 1497
rect 486 1501 492 1502
rect 486 1497 487 1501
rect 491 1497 492 1501
rect 486 1496 492 1497
rect 686 1501 692 1502
rect 686 1497 687 1501
rect 691 1497 692 1501
rect 686 1496 692 1497
rect 886 1501 892 1502
rect 886 1497 887 1501
rect 891 1497 892 1501
rect 886 1496 892 1497
rect 1078 1501 1084 1502
rect 1078 1497 1079 1501
rect 1083 1497 1084 1501
rect 1078 1496 1084 1497
rect 1262 1501 1268 1502
rect 1262 1497 1263 1501
rect 1267 1497 1268 1501
rect 1262 1496 1268 1497
rect 1446 1501 1452 1502
rect 1446 1497 1447 1501
rect 1451 1497 1452 1501
rect 1446 1496 1452 1497
rect 1622 1501 1628 1502
rect 1622 1497 1623 1501
rect 1627 1497 1628 1501
rect 1622 1496 1628 1497
rect 1806 1501 1812 1502
rect 1806 1497 1807 1501
rect 1811 1497 1812 1501
rect 1806 1496 1812 1497
rect 2006 1500 2012 1501
rect 2006 1496 2007 1500
rect 2011 1496 2012 1500
rect 110 1495 116 1496
rect 112 1475 114 1495
rect 136 1475 138 1496
rect 296 1475 298 1496
rect 488 1475 490 1496
rect 688 1475 690 1496
rect 888 1475 890 1496
rect 1080 1475 1082 1496
rect 1264 1475 1266 1496
rect 1448 1475 1450 1496
rect 1624 1475 1626 1496
rect 1808 1475 1810 1496
rect 2006 1495 2012 1496
rect 2008 1475 2010 1495
rect 2048 1491 2050 1511
rect 2584 1491 2586 1512
rect 2744 1491 2746 1512
rect 2904 1491 2906 1512
rect 3064 1491 3066 1512
rect 3224 1491 3226 1512
rect 3384 1491 3386 1512
rect 3544 1491 3546 1512
rect 3704 1491 3706 1512
rect 3942 1511 3948 1512
rect 3944 1491 3946 1511
rect 2047 1490 2051 1491
rect 2047 1485 2051 1486
rect 2415 1490 2419 1491
rect 2415 1485 2419 1486
rect 2511 1490 2515 1491
rect 2511 1485 2515 1486
rect 2583 1490 2587 1491
rect 2583 1485 2587 1486
rect 2607 1490 2611 1491
rect 2607 1485 2611 1486
rect 2703 1490 2707 1491
rect 2703 1485 2707 1486
rect 2743 1490 2747 1491
rect 2743 1485 2747 1486
rect 2799 1490 2803 1491
rect 2799 1485 2803 1486
rect 2903 1490 2907 1491
rect 2903 1485 2907 1486
rect 2919 1490 2923 1491
rect 2919 1485 2923 1486
rect 3063 1490 3067 1491
rect 3063 1485 3067 1486
rect 3223 1490 3227 1491
rect 3223 1485 3227 1486
rect 3231 1490 3235 1491
rect 3231 1485 3235 1486
rect 3383 1490 3387 1491
rect 3383 1485 3387 1486
rect 3415 1490 3419 1491
rect 3415 1485 3419 1486
rect 3543 1490 3547 1491
rect 3543 1485 3547 1486
rect 3615 1490 3619 1491
rect 3615 1485 3619 1486
rect 3703 1490 3707 1491
rect 3703 1485 3707 1486
rect 3815 1490 3819 1491
rect 3815 1485 3819 1486
rect 3943 1490 3947 1491
rect 3943 1485 3947 1486
rect 111 1474 115 1475
rect 111 1469 115 1470
rect 135 1474 139 1475
rect 135 1469 139 1470
rect 175 1474 179 1475
rect 175 1469 179 1470
rect 295 1474 299 1475
rect 295 1469 299 1470
rect 359 1474 363 1475
rect 359 1469 363 1470
rect 487 1474 491 1475
rect 487 1469 491 1470
rect 567 1474 571 1475
rect 567 1469 571 1470
rect 687 1474 691 1475
rect 687 1469 691 1470
rect 783 1474 787 1475
rect 783 1469 787 1470
rect 887 1474 891 1475
rect 887 1469 891 1470
rect 1007 1474 1011 1475
rect 1007 1469 1011 1470
rect 1079 1474 1083 1475
rect 1079 1469 1083 1470
rect 1231 1474 1235 1475
rect 1231 1469 1235 1470
rect 1263 1474 1267 1475
rect 1263 1469 1267 1470
rect 1447 1474 1451 1475
rect 1447 1469 1451 1470
rect 1463 1474 1467 1475
rect 1463 1469 1467 1470
rect 1623 1474 1627 1475
rect 1623 1469 1627 1470
rect 1695 1474 1699 1475
rect 1695 1469 1699 1470
rect 1807 1474 1811 1475
rect 1807 1469 1811 1470
rect 1903 1474 1907 1475
rect 1903 1469 1907 1470
rect 2007 1474 2011 1475
rect 2007 1469 2011 1470
rect 112 1449 114 1469
rect 110 1448 116 1449
rect 176 1448 178 1469
rect 360 1448 362 1469
rect 568 1448 570 1469
rect 784 1448 786 1469
rect 1008 1448 1010 1469
rect 1232 1448 1234 1469
rect 1464 1448 1466 1469
rect 1696 1448 1698 1469
rect 1904 1448 1906 1469
rect 2008 1449 2010 1469
rect 2048 1465 2050 1485
rect 2046 1464 2052 1465
rect 2416 1464 2418 1485
rect 2512 1464 2514 1485
rect 2608 1464 2610 1485
rect 2704 1464 2706 1485
rect 2800 1464 2802 1485
rect 2920 1464 2922 1485
rect 3064 1464 3066 1485
rect 3232 1464 3234 1485
rect 3416 1464 3418 1485
rect 3616 1464 3618 1485
rect 3816 1464 3818 1485
rect 3944 1465 3946 1485
rect 3942 1464 3948 1465
rect 2046 1460 2047 1464
rect 2051 1460 2052 1464
rect 2046 1459 2052 1460
rect 2414 1463 2420 1464
rect 2414 1459 2415 1463
rect 2419 1459 2420 1463
rect 2414 1458 2420 1459
rect 2510 1463 2516 1464
rect 2510 1459 2511 1463
rect 2515 1459 2516 1463
rect 2510 1458 2516 1459
rect 2606 1463 2612 1464
rect 2606 1459 2607 1463
rect 2611 1459 2612 1463
rect 2606 1458 2612 1459
rect 2702 1463 2708 1464
rect 2702 1459 2703 1463
rect 2707 1459 2708 1463
rect 2702 1458 2708 1459
rect 2798 1463 2804 1464
rect 2798 1459 2799 1463
rect 2803 1459 2804 1463
rect 2798 1458 2804 1459
rect 2918 1463 2924 1464
rect 2918 1459 2919 1463
rect 2923 1459 2924 1463
rect 2918 1458 2924 1459
rect 3062 1463 3068 1464
rect 3062 1459 3063 1463
rect 3067 1459 3068 1463
rect 3062 1458 3068 1459
rect 3230 1463 3236 1464
rect 3230 1459 3231 1463
rect 3235 1459 3236 1463
rect 3230 1458 3236 1459
rect 3414 1463 3420 1464
rect 3414 1459 3415 1463
rect 3419 1459 3420 1463
rect 3414 1458 3420 1459
rect 3614 1463 3620 1464
rect 3614 1459 3615 1463
rect 3619 1459 3620 1463
rect 3614 1458 3620 1459
rect 3814 1463 3820 1464
rect 3814 1459 3815 1463
rect 3819 1459 3820 1463
rect 3942 1460 3943 1464
rect 3947 1460 3948 1464
rect 3942 1459 3948 1460
rect 3814 1458 3820 1459
rect 2006 1448 2012 1449
rect 110 1444 111 1448
rect 115 1444 116 1448
rect 110 1443 116 1444
rect 174 1447 180 1448
rect 174 1443 175 1447
rect 179 1443 180 1447
rect 174 1442 180 1443
rect 358 1447 364 1448
rect 358 1443 359 1447
rect 363 1443 364 1447
rect 358 1442 364 1443
rect 566 1447 572 1448
rect 566 1443 567 1447
rect 571 1443 572 1447
rect 566 1442 572 1443
rect 782 1447 788 1448
rect 782 1443 783 1447
rect 787 1443 788 1447
rect 782 1442 788 1443
rect 1006 1447 1012 1448
rect 1006 1443 1007 1447
rect 1011 1443 1012 1447
rect 1006 1442 1012 1443
rect 1230 1447 1236 1448
rect 1230 1443 1231 1447
rect 1235 1443 1236 1447
rect 1230 1442 1236 1443
rect 1462 1447 1468 1448
rect 1462 1443 1463 1447
rect 1467 1443 1468 1447
rect 1462 1442 1468 1443
rect 1694 1447 1700 1448
rect 1694 1443 1695 1447
rect 1699 1443 1700 1447
rect 1694 1442 1700 1443
rect 1902 1447 1908 1448
rect 1902 1443 1903 1447
rect 1907 1443 1908 1447
rect 2006 1444 2007 1448
rect 2011 1444 2012 1448
rect 2006 1443 2012 1444
rect 2046 1447 2052 1448
rect 2046 1443 2047 1447
rect 2051 1443 2052 1447
rect 3942 1447 3948 1448
rect 1902 1442 1908 1443
rect 2046 1442 2052 1443
rect 2414 1444 2420 1445
rect 110 1431 116 1432
rect 110 1427 111 1431
rect 115 1427 116 1431
rect 2006 1431 2012 1432
rect 110 1426 116 1427
rect 174 1428 180 1429
rect 112 1399 114 1426
rect 174 1424 175 1428
rect 179 1424 180 1428
rect 174 1423 180 1424
rect 358 1428 364 1429
rect 358 1424 359 1428
rect 363 1424 364 1428
rect 358 1423 364 1424
rect 566 1428 572 1429
rect 566 1424 567 1428
rect 571 1424 572 1428
rect 566 1423 572 1424
rect 782 1428 788 1429
rect 782 1424 783 1428
rect 787 1424 788 1428
rect 782 1423 788 1424
rect 1006 1428 1012 1429
rect 1006 1424 1007 1428
rect 1011 1424 1012 1428
rect 1006 1423 1012 1424
rect 1230 1428 1236 1429
rect 1230 1424 1231 1428
rect 1235 1424 1236 1428
rect 1230 1423 1236 1424
rect 1462 1428 1468 1429
rect 1462 1424 1463 1428
rect 1467 1424 1468 1428
rect 1462 1423 1468 1424
rect 1694 1428 1700 1429
rect 1694 1424 1695 1428
rect 1699 1424 1700 1428
rect 1694 1423 1700 1424
rect 1902 1428 1908 1429
rect 1902 1424 1903 1428
rect 1907 1424 1908 1428
rect 2006 1427 2007 1431
rect 2011 1427 2012 1431
rect 2006 1426 2012 1427
rect 1902 1423 1908 1424
rect 176 1399 178 1423
rect 360 1399 362 1423
rect 568 1399 570 1423
rect 784 1399 786 1423
rect 1008 1399 1010 1423
rect 1232 1399 1234 1423
rect 1464 1399 1466 1423
rect 1696 1399 1698 1423
rect 1904 1399 1906 1423
rect 2008 1399 2010 1426
rect 111 1398 115 1399
rect 111 1393 115 1394
rect 175 1398 179 1399
rect 175 1393 179 1394
rect 327 1398 331 1399
rect 327 1393 331 1394
rect 359 1398 363 1399
rect 359 1393 363 1394
rect 463 1398 467 1399
rect 463 1393 467 1394
rect 567 1398 571 1399
rect 567 1393 571 1394
rect 599 1398 603 1399
rect 599 1393 603 1394
rect 727 1398 731 1399
rect 727 1393 731 1394
rect 783 1398 787 1399
rect 783 1393 787 1394
rect 855 1398 859 1399
rect 855 1393 859 1394
rect 983 1398 987 1399
rect 983 1393 987 1394
rect 1007 1398 1011 1399
rect 1007 1393 1011 1394
rect 1119 1398 1123 1399
rect 1119 1393 1123 1394
rect 1231 1398 1235 1399
rect 1231 1393 1235 1394
rect 1263 1398 1267 1399
rect 1263 1393 1267 1394
rect 1423 1398 1427 1399
rect 1423 1393 1427 1394
rect 1463 1398 1467 1399
rect 1463 1393 1467 1394
rect 1583 1398 1587 1399
rect 1583 1393 1587 1394
rect 1695 1398 1699 1399
rect 1695 1393 1699 1394
rect 1751 1398 1755 1399
rect 1751 1393 1755 1394
rect 1903 1398 1907 1399
rect 1903 1393 1907 1394
rect 2007 1398 2011 1399
rect 2048 1395 2050 1442
rect 2414 1440 2415 1444
rect 2419 1440 2420 1444
rect 2414 1439 2420 1440
rect 2510 1444 2516 1445
rect 2510 1440 2511 1444
rect 2515 1440 2516 1444
rect 2510 1439 2516 1440
rect 2606 1444 2612 1445
rect 2606 1440 2607 1444
rect 2611 1440 2612 1444
rect 2606 1439 2612 1440
rect 2702 1444 2708 1445
rect 2702 1440 2703 1444
rect 2707 1440 2708 1444
rect 2702 1439 2708 1440
rect 2798 1444 2804 1445
rect 2798 1440 2799 1444
rect 2803 1440 2804 1444
rect 2798 1439 2804 1440
rect 2918 1444 2924 1445
rect 2918 1440 2919 1444
rect 2923 1440 2924 1444
rect 2918 1439 2924 1440
rect 3062 1444 3068 1445
rect 3062 1440 3063 1444
rect 3067 1440 3068 1444
rect 3062 1439 3068 1440
rect 3230 1444 3236 1445
rect 3230 1440 3231 1444
rect 3235 1440 3236 1444
rect 3230 1439 3236 1440
rect 3414 1444 3420 1445
rect 3414 1440 3415 1444
rect 3419 1440 3420 1444
rect 3414 1439 3420 1440
rect 3614 1444 3620 1445
rect 3614 1440 3615 1444
rect 3619 1440 3620 1444
rect 3614 1439 3620 1440
rect 3814 1444 3820 1445
rect 3814 1440 3815 1444
rect 3819 1440 3820 1444
rect 3942 1443 3943 1447
rect 3947 1443 3948 1447
rect 3942 1442 3948 1443
rect 3814 1439 3820 1440
rect 2416 1395 2418 1439
rect 2512 1395 2514 1439
rect 2608 1395 2610 1439
rect 2704 1395 2706 1439
rect 2800 1395 2802 1439
rect 2920 1395 2922 1439
rect 3064 1395 3066 1439
rect 3232 1395 3234 1439
rect 3416 1395 3418 1439
rect 3616 1395 3618 1439
rect 3816 1395 3818 1439
rect 3944 1395 3946 1442
rect 2007 1393 2011 1394
rect 2047 1394 2051 1395
rect 112 1366 114 1393
rect 328 1369 330 1393
rect 464 1369 466 1393
rect 600 1369 602 1393
rect 728 1369 730 1393
rect 856 1369 858 1393
rect 984 1369 986 1393
rect 1120 1369 1122 1393
rect 1264 1369 1266 1393
rect 1424 1369 1426 1393
rect 1584 1369 1586 1393
rect 1752 1369 1754 1393
rect 1904 1369 1906 1393
rect 326 1368 332 1369
rect 110 1365 116 1366
rect 110 1361 111 1365
rect 115 1361 116 1365
rect 326 1364 327 1368
rect 331 1364 332 1368
rect 326 1363 332 1364
rect 462 1368 468 1369
rect 462 1364 463 1368
rect 467 1364 468 1368
rect 462 1363 468 1364
rect 598 1368 604 1369
rect 598 1364 599 1368
rect 603 1364 604 1368
rect 598 1363 604 1364
rect 726 1368 732 1369
rect 726 1364 727 1368
rect 731 1364 732 1368
rect 726 1363 732 1364
rect 854 1368 860 1369
rect 854 1364 855 1368
rect 859 1364 860 1368
rect 854 1363 860 1364
rect 982 1368 988 1369
rect 982 1364 983 1368
rect 987 1364 988 1368
rect 982 1363 988 1364
rect 1118 1368 1124 1369
rect 1118 1364 1119 1368
rect 1123 1364 1124 1368
rect 1118 1363 1124 1364
rect 1262 1368 1268 1369
rect 1262 1364 1263 1368
rect 1267 1364 1268 1368
rect 1262 1363 1268 1364
rect 1422 1368 1428 1369
rect 1422 1364 1423 1368
rect 1427 1364 1428 1368
rect 1422 1363 1428 1364
rect 1582 1368 1588 1369
rect 1582 1364 1583 1368
rect 1587 1364 1588 1368
rect 1582 1363 1588 1364
rect 1750 1368 1756 1369
rect 1750 1364 1751 1368
rect 1755 1364 1756 1368
rect 1750 1363 1756 1364
rect 1902 1368 1908 1369
rect 1902 1364 1903 1368
rect 1907 1364 1908 1368
rect 2008 1366 2010 1393
rect 2047 1389 2051 1390
rect 2071 1394 2075 1395
rect 2071 1389 2075 1390
rect 2303 1394 2307 1395
rect 2303 1389 2307 1390
rect 2415 1394 2419 1395
rect 2415 1389 2419 1390
rect 2511 1394 2515 1395
rect 2511 1389 2515 1390
rect 2559 1394 2563 1395
rect 2559 1389 2563 1390
rect 2607 1394 2611 1395
rect 2607 1389 2611 1390
rect 2703 1394 2707 1395
rect 2703 1389 2707 1390
rect 2799 1394 2803 1395
rect 2799 1389 2803 1390
rect 2807 1394 2811 1395
rect 2807 1389 2811 1390
rect 2919 1394 2923 1395
rect 2919 1389 2923 1390
rect 3055 1394 3059 1395
rect 3055 1389 3059 1390
rect 3063 1394 3067 1395
rect 3063 1389 3067 1390
rect 3231 1394 3235 1395
rect 3231 1389 3235 1390
rect 3303 1394 3307 1395
rect 3303 1389 3307 1390
rect 3415 1394 3419 1395
rect 3415 1389 3419 1390
rect 3559 1394 3563 1395
rect 3559 1389 3563 1390
rect 3615 1394 3619 1395
rect 3615 1389 3619 1390
rect 3815 1394 3819 1395
rect 3815 1389 3819 1390
rect 3943 1394 3947 1395
rect 3943 1389 3947 1390
rect 1902 1363 1908 1364
rect 2006 1365 2012 1366
rect 110 1360 116 1361
rect 2006 1361 2007 1365
rect 2011 1361 2012 1365
rect 2048 1362 2050 1389
rect 2072 1365 2074 1389
rect 2304 1365 2306 1389
rect 2560 1365 2562 1389
rect 2808 1365 2810 1389
rect 3056 1365 3058 1389
rect 3304 1365 3306 1389
rect 3560 1365 3562 1389
rect 3816 1365 3818 1389
rect 2070 1364 2076 1365
rect 2006 1360 2012 1361
rect 2046 1361 2052 1362
rect 2046 1357 2047 1361
rect 2051 1357 2052 1361
rect 2070 1360 2071 1364
rect 2075 1360 2076 1364
rect 2070 1359 2076 1360
rect 2302 1364 2308 1365
rect 2302 1360 2303 1364
rect 2307 1360 2308 1364
rect 2302 1359 2308 1360
rect 2558 1364 2564 1365
rect 2558 1360 2559 1364
rect 2563 1360 2564 1364
rect 2558 1359 2564 1360
rect 2806 1364 2812 1365
rect 2806 1360 2807 1364
rect 2811 1360 2812 1364
rect 2806 1359 2812 1360
rect 3054 1364 3060 1365
rect 3054 1360 3055 1364
rect 3059 1360 3060 1364
rect 3054 1359 3060 1360
rect 3302 1364 3308 1365
rect 3302 1360 3303 1364
rect 3307 1360 3308 1364
rect 3302 1359 3308 1360
rect 3558 1364 3564 1365
rect 3558 1360 3559 1364
rect 3563 1360 3564 1364
rect 3558 1359 3564 1360
rect 3814 1364 3820 1365
rect 3814 1360 3815 1364
rect 3819 1360 3820 1364
rect 3944 1362 3946 1389
rect 3814 1359 3820 1360
rect 3942 1361 3948 1362
rect 2046 1356 2052 1357
rect 3942 1357 3943 1361
rect 3947 1357 3948 1361
rect 3942 1356 3948 1357
rect 326 1349 332 1350
rect 110 1348 116 1349
rect 110 1344 111 1348
rect 115 1344 116 1348
rect 326 1345 327 1349
rect 331 1345 332 1349
rect 326 1344 332 1345
rect 462 1349 468 1350
rect 462 1345 463 1349
rect 467 1345 468 1349
rect 462 1344 468 1345
rect 598 1349 604 1350
rect 598 1345 599 1349
rect 603 1345 604 1349
rect 598 1344 604 1345
rect 726 1349 732 1350
rect 726 1345 727 1349
rect 731 1345 732 1349
rect 726 1344 732 1345
rect 854 1349 860 1350
rect 854 1345 855 1349
rect 859 1345 860 1349
rect 854 1344 860 1345
rect 982 1349 988 1350
rect 982 1345 983 1349
rect 987 1345 988 1349
rect 982 1344 988 1345
rect 1118 1349 1124 1350
rect 1118 1345 1119 1349
rect 1123 1345 1124 1349
rect 1118 1344 1124 1345
rect 1262 1349 1268 1350
rect 1262 1345 1263 1349
rect 1267 1345 1268 1349
rect 1262 1344 1268 1345
rect 1422 1349 1428 1350
rect 1422 1345 1423 1349
rect 1427 1345 1428 1349
rect 1422 1344 1428 1345
rect 1582 1349 1588 1350
rect 1582 1345 1583 1349
rect 1587 1345 1588 1349
rect 1582 1344 1588 1345
rect 1750 1349 1756 1350
rect 1750 1345 1751 1349
rect 1755 1345 1756 1349
rect 1750 1344 1756 1345
rect 1902 1349 1908 1350
rect 1902 1345 1903 1349
rect 1907 1345 1908 1349
rect 1902 1344 1908 1345
rect 2006 1348 2012 1349
rect 2006 1344 2007 1348
rect 2011 1344 2012 1348
rect 2070 1345 2076 1346
rect 110 1343 116 1344
rect 112 1315 114 1343
rect 328 1315 330 1344
rect 464 1315 466 1344
rect 600 1315 602 1344
rect 728 1315 730 1344
rect 856 1315 858 1344
rect 984 1315 986 1344
rect 1120 1315 1122 1344
rect 1264 1315 1266 1344
rect 1424 1315 1426 1344
rect 1584 1315 1586 1344
rect 1752 1315 1754 1344
rect 1904 1315 1906 1344
rect 2006 1343 2012 1344
rect 2046 1344 2052 1345
rect 2008 1315 2010 1343
rect 2046 1340 2047 1344
rect 2051 1340 2052 1344
rect 2070 1341 2071 1345
rect 2075 1341 2076 1345
rect 2070 1340 2076 1341
rect 2302 1345 2308 1346
rect 2302 1341 2303 1345
rect 2307 1341 2308 1345
rect 2302 1340 2308 1341
rect 2558 1345 2564 1346
rect 2558 1341 2559 1345
rect 2563 1341 2564 1345
rect 2558 1340 2564 1341
rect 2806 1345 2812 1346
rect 2806 1341 2807 1345
rect 2811 1341 2812 1345
rect 2806 1340 2812 1341
rect 3054 1345 3060 1346
rect 3054 1341 3055 1345
rect 3059 1341 3060 1345
rect 3054 1340 3060 1341
rect 3302 1345 3308 1346
rect 3302 1341 3303 1345
rect 3307 1341 3308 1345
rect 3302 1340 3308 1341
rect 3558 1345 3564 1346
rect 3558 1341 3559 1345
rect 3563 1341 3564 1345
rect 3558 1340 3564 1341
rect 3814 1345 3820 1346
rect 3814 1341 3815 1345
rect 3819 1341 3820 1345
rect 3814 1340 3820 1341
rect 3942 1344 3948 1345
rect 3942 1340 3943 1344
rect 3947 1340 3948 1344
rect 2046 1339 2052 1340
rect 111 1314 115 1315
rect 111 1309 115 1310
rect 327 1314 331 1315
rect 327 1309 331 1310
rect 463 1314 467 1315
rect 463 1309 467 1310
rect 551 1314 555 1315
rect 551 1309 555 1310
rect 599 1314 603 1315
rect 599 1309 603 1310
rect 655 1314 659 1315
rect 655 1309 659 1310
rect 727 1314 731 1315
rect 727 1309 731 1310
rect 767 1314 771 1315
rect 767 1309 771 1310
rect 855 1314 859 1315
rect 855 1309 859 1310
rect 879 1314 883 1315
rect 879 1309 883 1310
rect 983 1314 987 1315
rect 983 1309 987 1310
rect 991 1314 995 1315
rect 991 1309 995 1310
rect 1103 1314 1107 1315
rect 1103 1309 1107 1310
rect 1119 1314 1123 1315
rect 1119 1309 1123 1310
rect 1215 1314 1219 1315
rect 1215 1309 1219 1310
rect 1263 1314 1267 1315
rect 1263 1309 1267 1310
rect 1327 1314 1331 1315
rect 1327 1309 1331 1310
rect 1423 1314 1427 1315
rect 1423 1309 1427 1310
rect 1439 1314 1443 1315
rect 1439 1309 1443 1310
rect 1559 1314 1563 1315
rect 1559 1309 1563 1310
rect 1583 1314 1587 1315
rect 1583 1309 1587 1310
rect 1751 1314 1755 1315
rect 1751 1309 1755 1310
rect 1903 1314 1907 1315
rect 1903 1309 1907 1310
rect 2007 1314 2011 1315
rect 2048 1311 2050 1339
rect 2072 1311 2074 1340
rect 2304 1311 2306 1340
rect 2560 1311 2562 1340
rect 2808 1311 2810 1340
rect 3056 1311 3058 1340
rect 3304 1311 3306 1340
rect 3560 1311 3562 1340
rect 3816 1311 3818 1340
rect 3942 1339 3948 1340
rect 3944 1311 3946 1339
rect 2007 1309 2011 1310
rect 2047 1310 2051 1311
rect 112 1289 114 1309
rect 110 1288 116 1289
rect 552 1288 554 1309
rect 656 1288 658 1309
rect 768 1288 770 1309
rect 880 1288 882 1309
rect 992 1288 994 1309
rect 1104 1288 1106 1309
rect 1216 1288 1218 1309
rect 1328 1288 1330 1309
rect 1440 1288 1442 1309
rect 1560 1288 1562 1309
rect 2008 1289 2010 1309
rect 2047 1305 2051 1306
rect 2071 1310 2075 1311
rect 2071 1305 2075 1306
rect 2223 1310 2227 1311
rect 2223 1305 2227 1306
rect 2303 1310 2307 1311
rect 2303 1305 2307 1306
rect 2415 1310 2419 1311
rect 2415 1305 2419 1306
rect 2559 1310 2563 1311
rect 2559 1305 2563 1306
rect 2615 1310 2619 1311
rect 2615 1305 2619 1306
rect 2807 1310 2811 1311
rect 2807 1305 2811 1306
rect 2815 1310 2819 1311
rect 2815 1305 2819 1306
rect 2999 1310 3003 1311
rect 2999 1305 3003 1306
rect 3055 1310 3059 1311
rect 3055 1305 3059 1306
rect 3175 1310 3179 1311
rect 3175 1305 3179 1306
rect 3303 1310 3307 1311
rect 3303 1305 3307 1306
rect 3343 1310 3347 1311
rect 3343 1305 3347 1306
rect 3503 1310 3507 1311
rect 3503 1305 3507 1306
rect 3559 1310 3563 1311
rect 3559 1305 3563 1306
rect 3663 1310 3667 1311
rect 3663 1305 3667 1306
rect 3815 1310 3819 1311
rect 3815 1305 3819 1306
rect 3831 1310 3835 1311
rect 3831 1305 3835 1306
rect 3943 1310 3947 1311
rect 3943 1305 3947 1306
rect 2006 1288 2012 1289
rect 110 1284 111 1288
rect 115 1284 116 1288
rect 110 1283 116 1284
rect 550 1287 556 1288
rect 550 1283 551 1287
rect 555 1283 556 1287
rect 550 1282 556 1283
rect 654 1287 660 1288
rect 654 1283 655 1287
rect 659 1283 660 1287
rect 654 1282 660 1283
rect 766 1287 772 1288
rect 766 1283 767 1287
rect 771 1283 772 1287
rect 766 1282 772 1283
rect 878 1287 884 1288
rect 878 1283 879 1287
rect 883 1283 884 1287
rect 878 1282 884 1283
rect 990 1287 996 1288
rect 990 1283 991 1287
rect 995 1283 996 1287
rect 990 1282 996 1283
rect 1102 1287 1108 1288
rect 1102 1283 1103 1287
rect 1107 1283 1108 1287
rect 1102 1282 1108 1283
rect 1214 1287 1220 1288
rect 1214 1283 1215 1287
rect 1219 1283 1220 1287
rect 1214 1282 1220 1283
rect 1326 1287 1332 1288
rect 1326 1283 1327 1287
rect 1331 1283 1332 1287
rect 1326 1282 1332 1283
rect 1438 1287 1444 1288
rect 1438 1283 1439 1287
rect 1443 1283 1444 1287
rect 1438 1282 1444 1283
rect 1558 1287 1564 1288
rect 1558 1283 1559 1287
rect 1563 1283 1564 1287
rect 2006 1284 2007 1288
rect 2011 1284 2012 1288
rect 2048 1285 2050 1305
rect 2006 1283 2012 1284
rect 2046 1284 2052 1285
rect 2072 1284 2074 1305
rect 2224 1284 2226 1305
rect 2416 1284 2418 1305
rect 2616 1284 2618 1305
rect 2816 1284 2818 1305
rect 3000 1284 3002 1305
rect 3176 1284 3178 1305
rect 3344 1284 3346 1305
rect 3504 1284 3506 1305
rect 3664 1284 3666 1305
rect 3832 1284 3834 1305
rect 3944 1285 3946 1305
rect 3942 1284 3948 1285
rect 1558 1282 1564 1283
rect 2046 1280 2047 1284
rect 2051 1280 2052 1284
rect 2046 1279 2052 1280
rect 2070 1283 2076 1284
rect 2070 1279 2071 1283
rect 2075 1279 2076 1283
rect 2070 1278 2076 1279
rect 2222 1283 2228 1284
rect 2222 1279 2223 1283
rect 2227 1279 2228 1283
rect 2222 1278 2228 1279
rect 2414 1283 2420 1284
rect 2414 1279 2415 1283
rect 2419 1279 2420 1283
rect 2414 1278 2420 1279
rect 2614 1283 2620 1284
rect 2614 1279 2615 1283
rect 2619 1279 2620 1283
rect 2614 1278 2620 1279
rect 2814 1283 2820 1284
rect 2814 1279 2815 1283
rect 2819 1279 2820 1283
rect 2814 1278 2820 1279
rect 2998 1283 3004 1284
rect 2998 1279 2999 1283
rect 3003 1279 3004 1283
rect 2998 1278 3004 1279
rect 3174 1283 3180 1284
rect 3174 1279 3175 1283
rect 3179 1279 3180 1283
rect 3174 1278 3180 1279
rect 3342 1283 3348 1284
rect 3342 1279 3343 1283
rect 3347 1279 3348 1283
rect 3342 1278 3348 1279
rect 3502 1283 3508 1284
rect 3502 1279 3503 1283
rect 3507 1279 3508 1283
rect 3502 1278 3508 1279
rect 3662 1283 3668 1284
rect 3662 1279 3663 1283
rect 3667 1279 3668 1283
rect 3662 1278 3668 1279
rect 3830 1283 3836 1284
rect 3830 1279 3831 1283
rect 3835 1279 3836 1283
rect 3942 1280 3943 1284
rect 3947 1280 3948 1284
rect 3942 1279 3948 1280
rect 3830 1278 3836 1279
rect 110 1271 116 1272
rect 110 1267 111 1271
rect 115 1267 116 1271
rect 2006 1271 2012 1272
rect 110 1266 116 1267
rect 550 1268 556 1269
rect 112 1239 114 1266
rect 550 1264 551 1268
rect 555 1264 556 1268
rect 550 1263 556 1264
rect 654 1268 660 1269
rect 654 1264 655 1268
rect 659 1264 660 1268
rect 654 1263 660 1264
rect 766 1268 772 1269
rect 766 1264 767 1268
rect 771 1264 772 1268
rect 766 1263 772 1264
rect 878 1268 884 1269
rect 878 1264 879 1268
rect 883 1264 884 1268
rect 878 1263 884 1264
rect 990 1268 996 1269
rect 990 1264 991 1268
rect 995 1264 996 1268
rect 990 1263 996 1264
rect 1102 1268 1108 1269
rect 1102 1264 1103 1268
rect 1107 1264 1108 1268
rect 1102 1263 1108 1264
rect 1214 1268 1220 1269
rect 1214 1264 1215 1268
rect 1219 1264 1220 1268
rect 1214 1263 1220 1264
rect 1326 1268 1332 1269
rect 1326 1264 1327 1268
rect 1331 1264 1332 1268
rect 1326 1263 1332 1264
rect 1438 1268 1444 1269
rect 1438 1264 1439 1268
rect 1443 1264 1444 1268
rect 1438 1263 1444 1264
rect 1558 1268 1564 1269
rect 1558 1264 1559 1268
rect 1563 1264 1564 1268
rect 2006 1267 2007 1271
rect 2011 1267 2012 1271
rect 2006 1266 2012 1267
rect 2046 1267 2052 1268
rect 1558 1263 1564 1264
rect 552 1239 554 1263
rect 656 1239 658 1263
rect 768 1239 770 1263
rect 880 1239 882 1263
rect 992 1239 994 1263
rect 1104 1239 1106 1263
rect 1216 1239 1218 1263
rect 1328 1239 1330 1263
rect 1440 1239 1442 1263
rect 1560 1239 1562 1263
rect 2008 1239 2010 1266
rect 2046 1263 2047 1267
rect 2051 1263 2052 1267
rect 3942 1267 3948 1268
rect 2046 1262 2052 1263
rect 2070 1264 2076 1265
rect 111 1238 115 1239
rect 111 1233 115 1234
rect 391 1238 395 1239
rect 391 1233 395 1234
rect 519 1238 523 1239
rect 519 1233 523 1234
rect 551 1238 555 1239
rect 551 1233 555 1234
rect 655 1238 659 1239
rect 655 1233 659 1234
rect 663 1238 667 1239
rect 663 1233 667 1234
rect 767 1238 771 1239
rect 767 1233 771 1234
rect 807 1238 811 1239
rect 807 1233 811 1234
rect 879 1238 883 1239
rect 879 1233 883 1234
rect 959 1238 963 1239
rect 959 1233 963 1234
rect 991 1238 995 1239
rect 991 1233 995 1234
rect 1103 1238 1107 1239
rect 1103 1233 1107 1234
rect 1111 1238 1115 1239
rect 1111 1233 1115 1234
rect 1215 1238 1219 1239
rect 1215 1233 1219 1234
rect 1255 1238 1259 1239
rect 1255 1233 1259 1234
rect 1327 1238 1331 1239
rect 1327 1233 1331 1234
rect 1407 1238 1411 1239
rect 1407 1233 1411 1234
rect 1439 1238 1443 1239
rect 1439 1233 1443 1234
rect 1559 1238 1563 1239
rect 1559 1233 1563 1234
rect 1711 1238 1715 1239
rect 1711 1233 1715 1234
rect 2007 1238 2011 1239
rect 2007 1233 2011 1234
rect 112 1206 114 1233
rect 392 1209 394 1233
rect 520 1209 522 1233
rect 664 1209 666 1233
rect 808 1209 810 1233
rect 960 1209 962 1233
rect 1112 1209 1114 1233
rect 1256 1209 1258 1233
rect 1408 1209 1410 1233
rect 1560 1209 1562 1233
rect 1712 1209 1714 1233
rect 390 1208 396 1209
rect 110 1205 116 1206
rect 110 1201 111 1205
rect 115 1201 116 1205
rect 390 1204 391 1208
rect 395 1204 396 1208
rect 390 1203 396 1204
rect 518 1208 524 1209
rect 518 1204 519 1208
rect 523 1204 524 1208
rect 518 1203 524 1204
rect 662 1208 668 1209
rect 662 1204 663 1208
rect 667 1204 668 1208
rect 662 1203 668 1204
rect 806 1208 812 1209
rect 806 1204 807 1208
rect 811 1204 812 1208
rect 806 1203 812 1204
rect 958 1208 964 1209
rect 958 1204 959 1208
rect 963 1204 964 1208
rect 958 1203 964 1204
rect 1110 1208 1116 1209
rect 1110 1204 1111 1208
rect 1115 1204 1116 1208
rect 1110 1203 1116 1204
rect 1254 1208 1260 1209
rect 1254 1204 1255 1208
rect 1259 1204 1260 1208
rect 1254 1203 1260 1204
rect 1406 1208 1412 1209
rect 1406 1204 1407 1208
rect 1411 1204 1412 1208
rect 1406 1203 1412 1204
rect 1558 1208 1564 1209
rect 1558 1204 1559 1208
rect 1563 1204 1564 1208
rect 1558 1203 1564 1204
rect 1710 1208 1716 1209
rect 1710 1204 1711 1208
rect 1715 1204 1716 1208
rect 2008 1206 2010 1233
rect 2048 1227 2050 1262
rect 2070 1260 2071 1264
rect 2075 1260 2076 1264
rect 2070 1259 2076 1260
rect 2222 1264 2228 1265
rect 2222 1260 2223 1264
rect 2227 1260 2228 1264
rect 2222 1259 2228 1260
rect 2414 1264 2420 1265
rect 2414 1260 2415 1264
rect 2419 1260 2420 1264
rect 2414 1259 2420 1260
rect 2614 1264 2620 1265
rect 2614 1260 2615 1264
rect 2619 1260 2620 1264
rect 2614 1259 2620 1260
rect 2814 1264 2820 1265
rect 2814 1260 2815 1264
rect 2819 1260 2820 1264
rect 2814 1259 2820 1260
rect 2998 1264 3004 1265
rect 2998 1260 2999 1264
rect 3003 1260 3004 1264
rect 2998 1259 3004 1260
rect 3174 1264 3180 1265
rect 3174 1260 3175 1264
rect 3179 1260 3180 1264
rect 3174 1259 3180 1260
rect 3342 1264 3348 1265
rect 3342 1260 3343 1264
rect 3347 1260 3348 1264
rect 3342 1259 3348 1260
rect 3502 1264 3508 1265
rect 3502 1260 3503 1264
rect 3507 1260 3508 1264
rect 3502 1259 3508 1260
rect 3662 1264 3668 1265
rect 3662 1260 3663 1264
rect 3667 1260 3668 1264
rect 3662 1259 3668 1260
rect 3830 1264 3836 1265
rect 3830 1260 3831 1264
rect 3835 1260 3836 1264
rect 3942 1263 3943 1267
rect 3947 1263 3948 1267
rect 3942 1262 3948 1263
rect 3830 1259 3836 1260
rect 2072 1227 2074 1259
rect 2224 1227 2226 1259
rect 2416 1227 2418 1259
rect 2616 1227 2618 1259
rect 2816 1227 2818 1259
rect 3000 1227 3002 1259
rect 3176 1227 3178 1259
rect 3344 1227 3346 1259
rect 3504 1227 3506 1259
rect 3664 1227 3666 1259
rect 3832 1227 3834 1259
rect 3944 1227 3946 1262
rect 2047 1226 2051 1227
rect 2047 1221 2051 1222
rect 2071 1226 2075 1227
rect 2071 1221 2075 1222
rect 2135 1226 2139 1227
rect 2135 1221 2139 1222
rect 2223 1226 2227 1227
rect 2223 1221 2227 1222
rect 2311 1226 2315 1227
rect 2311 1221 2315 1222
rect 2415 1226 2419 1227
rect 2415 1221 2419 1222
rect 2503 1226 2507 1227
rect 2503 1221 2507 1222
rect 2615 1226 2619 1227
rect 2615 1221 2619 1222
rect 2695 1226 2699 1227
rect 2695 1221 2699 1222
rect 2815 1226 2819 1227
rect 2815 1221 2819 1222
rect 2887 1226 2891 1227
rect 2887 1221 2891 1222
rect 2999 1226 3003 1227
rect 2999 1221 3003 1222
rect 3071 1226 3075 1227
rect 3071 1221 3075 1222
rect 3175 1226 3179 1227
rect 3175 1221 3179 1222
rect 3239 1226 3243 1227
rect 3239 1221 3243 1222
rect 3343 1226 3347 1227
rect 3343 1221 3347 1222
rect 3399 1226 3403 1227
rect 3399 1221 3403 1222
rect 3503 1226 3507 1227
rect 3503 1221 3507 1222
rect 3551 1226 3555 1227
rect 3551 1221 3555 1222
rect 3663 1226 3667 1227
rect 3663 1221 3667 1222
rect 3703 1226 3707 1227
rect 3703 1221 3707 1222
rect 3831 1226 3835 1227
rect 3831 1221 3835 1222
rect 3839 1226 3843 1227
rect 3839 1221 3843 1222
rect 3943 1226 3947 1227
rect 3943 1221 3947 1222
rect 1710 1203 1716 1204
rect 2006 1205 2012 1206
rect 110 1200 116 1201
rect 2006 1201 2007 1205
rect 2011 1201 2012 1205
rect 2006 1200 2012 1201
rect 2048 1194 2050 1221
rect 2136 1197 2138 1221
rect 2312 1197 2314 1221
rect 2504 1197 2506 1221
rect 2696 1197 2698 1221
rect 2888 1197 2890 1221
rect 3072 1197 3074 1221
rect 3240 1197 3242 1221
rect 3400 1197 3402 1221
rect 3552 1197 3554 1221
rect 3704 1197 3706 1221
rect 3840 1197 3842 1221
rect 2134 1196 2140 1197
rect 2046 1193 2052 1194
rect 390 1189 396 1190
rect 110 1188 116 1189
rect 110 1184 111 1188
rect 115 1184 116 1188
rect 390 1185 391 1189
rect 395 1185 396 1189
rect 390 1184 396 1185
rect 518 1189 524 1190
rect 518 1185 519 1189
rect 523 1185 524 1189
rect 518 1184 524 1185
rect 662 1189 668 1190
rect 662 1185 663 1189
rect 667 1185 668 1189
rect 662 1184 668 1185
rect 806 1189 812 1190
rect 806 1185 807 1189
rect 811 1185 812 1189
rect 806 1184 812 1185
rect 958 1189 964 1190
rect 958 1185 959 1189
rect 963 1185 964 1189
rect 958 1184 964 1185
rect 1110 1189 1116 1190
rect 1110 1185 1111 1189
rect 1115 1185 1116 1189
rect 1110 1184 1116 1185
rect 1254 1189 1260 1190
rect 1254 1185 1255 1189
rect 1259 1185 1260 1189
rect 1254 1184 1260 1185
rect 1406 1189 1412 1190
rect 1406 1185 1407 1189
rect 1411 1185 1412 1189
rect 1406 1184 1412 1185
rect 1558 1189 1564 1190
rect 1558 1185 1559 1189
rect 1563 1185 1564 1189
rect 1558 1184 1564 1185
rect 1710 1189 1716 1190
rect 2046 1189 2047 1193
rect 2051 1189 2052 1193
rect 2134 1192 2135 1196
rect 2139 1192 2140 1196
rect 2134 1191 2140 1192
rect 2310 1196 2316 1197
rect 2310 1192 2311 1196
rect 2315 1192 2316 1196
rect 2310 1191 2316 1192
rect 2502 1196 2508 1197
rect 2502 1192 2503 1196
rect 2507 1192 2508 1196
rect 2502 1191 2508 1192
rect 2694 1196 2700 1197
rect 2694 1192 2695 1196
rect 2699 1192 2700 1196
rect 2694 1191 2700 1192
rect 2886 1196 2892 1197
rect 2886 1192 2887 1196
rect 2891 1192 2892 1196
rect 2886 1191 2892 1192
rect 3070 1196 3076 1197
rect 3070 1192 3071 1196
rect 3075 1192 3076 1196
rect 3070 1191 3076 1192
rect 3238 1196 3244 1197
rect 3238 1192 3239 1196
rect 3243 1192 3244 1196
rect 3238 1191 3244 1192
rect 3398 1196 3404 1197
rect 3398 1192 3399 1196
rect 3403 1192 3404 1196
rect 3398 1191 3404 1192
rect 3550 1196 3556 1197
rect 3550 1192 3551 1196
rect 3555 1192 3556 1196
rect 3550 1191 3556 1192
rect 3702 1196 3708 1197
rect 3702 1192 3703 1196
rect 3707 1192 3708 1196
rect 3702 1191 3708 1192
rect 3838 1196 3844 1197
rect 3838 1192 3839 1196
rect 3843 1192 3844 1196
rect 3944 1194 3946 1221
rect 3838 1191 3844 1192
rect 3942 1193 3948 1194
rect 1710 1185 1711 1189
rect 1715 1185 1716 1189
rect 1710 1184 1716 1185
rect 2006 1188 2012 1189
rect 2046 1188 2052 1189
rect 3942 1189 3943 1193
rect 3947 1189 3948 1193
rect 3942 1188 3948 1189
rect 2006 1184 2007 1188
rect 2011 1184 2012 1188
rect 110 1183 116 1184
rect 112 1159 114 1183
rect 392 1159 394 1184
rect 520 1159 522 1184
rect 664 1159 666 1184
rect 808 1159 810 1184
rect 960 1159 962 1184
rect 1112 1159 1114 1184
rect 1256 1159 1258 1184
rect 1408 1159 1410 1184
rect 1560 1159 1562 1184
rect 1712 1159 1714 1184
rect 2006 1183 2012 1184
rect 2008 1159 2010 1183
rect 2134 1177 2140 1178
rect 2046 1176 2052 1177
rect 2046 1172 2047 1176
rect 2051 1172 2052 1176
rect 2134 1173 2135 1177
rect 2139 1173 2140 1177
rect 2134 1172 2140 1173
rect 2310 1177 2316 1178
rect 2310 1173 2311 1177
rect 2315 1173 2316 1177
rect 2310 1172 2316 1173
rect 2502 1177 2508 1178
rect 2502 1173 2503 1177
rect 2507 1173 2508 1177
rect 2502 1172 2508 1173
rect 2694 1177 2700 1178
rect 2694 1173 2695 1177
rect 2699 1173 2700 1177
rect 2694 1172 2700 1173
rect 2886 1177 2892 1178
rect 2886 1173 2887 1177
rect 2891 1173 2892 1177
rect 2886 1172 2892 1173
rect 3070 1177 3076 1178
rect 3070 1173 3071 1177
rect 3075 1173 3076 1177
rect 3070 1172 3076 1173
rect 3238 1177 3244 1178
rect 3238 1173 3239 1177
rect 3243 1173 3244 1177
rect 3238 1172 3244 1173
rect 3398 1177 3404 1178
rect 3398 1173 3399 1177
rect 3403 1173 3404 1177
rect 3398 1172 3404 1173
rect 3550 1177 3556 1178
rect 3550 1173 3551 1177
rect 3555 1173 3556 1177
rect 3550 1172 3556 1173
rect 3702 1177 3708 1178
rect 3702 1173 3703 1177
rect 3707 1173 3708 1177
rect 3702 1172 3708 1173
rect 3838 1177 3844 1178
rect 3838 1173 3839 1177
rect 3843 1173 3844 1177
rect 3838 1172 3844 1173
rect 3942 1176 3948 1177
rect 3942 1172 3943 1176
rect 3947 1172 3948 1176
rect 2046 1171 2052 1172
rect 111 1158 115 1159
rect 111 1153 115 1154
rect 175 1158 179 1159
rect 175 1153 179 1154
rect 327 1158 331 1159
rect 327 1153 331 1154
rect 391 1158 395 1159
rect 391 1153 395 1154
rect 495 1158 499 1159
rect 495 1153 499 1154
rect 519 1158 523 1159
rect 519 1153 523 1154
rect 663 1158 667 1159
rect 663 1153 667 1154
rect 671 1158 675 1159
rect 671 1153 675 1154
rect 807 1158 811 1159
rect 807 1153 811 1154
rect 847 1158 851 1159
rect 847 1153 851 1154
rect 959 1158 963 1159
rect 959 1153 963 1154
rect 1031 1158 1035 1159
rect 1031 1153 1035 1154
rect 1111 1158 1115 1159
rect 1111 1153 1115 1154
rect 1207 1158 1211 1159
rect 1207 1153 1211 1154
rect 1255 1158 1259 1159
rect 1255 1153 1259 1154
rect 1383 1158 1387 1159
rect 1383 1153 1387 1154
rect 1407 1158 1411 1159
rect 1407 1153 1411 1154
rect 1559 1158 1563 1159
rect 1559 1153 1563 1154
rect 1567 1158 1571 1159
rect 1567 1153 1571 1154
rect 1711 1158 1715 1159
rect 1711 1153 1715 1154
rect 1751 1158 1755 1159
rect 1751 1153 1755 1154
rect 2007 1158 2011 1159
rect 2007 1153 2011 1154
rect 112 1133 114 1153
rect 110 1132 116 1133
rect 176 1132 178 1153
rect 328 1132 330 1153
rect 496 1132 498 1153
rect 672 1132 674 1153
rect 848 1132 850 1153
rect 1032 1132 1034 1153
rect 1208 1132 1210 1153
rect 1384 1132 1386 1153
rect 1568 1132 1570 1153
rect 1752 1132 1754 1153
rect 2008 1133 2010 1153
rect 2048 1143 2050 1171
rect 2136 1143 2138 1172
rect 2312 1143 2314 1172
rect 2504 1143 2506 1172
rect 2696 1143 2698 1172
rect 2888 1143 2890 1172
rect 3072 1143 3074 1172
rect 3240 1143 3242 1172
rect 3400 1143 3402 1172
rect 3552 1143 3554 1172
rect 3704 1143 3706 1172
rect 3840 1143 3842 1172
rect 3942 1171 3948 1172
rect 3944 1143 3946 1171
rect 2047 1142 2051 1143
rect 2047 1137 2051 1138
rect 2135 1142 2139 1143
rect 2135 1137 2139 1138
rect 2295 1142 2299 1143
rect 2295 1137 2299 1138
rect 2311 1142 2315 1143
rect 2311 1137 2315 1138
rect 2423 1142 2427 1143
rect 2423 1137 2427 1138
rect 2503 1142 2507 1143
rect 2503 1137 2507 1138
rect 2559 1142 2563 1143
rect 2559 1137 2563 1138
rect 2695 1142 2699 1143
rect 2695 1137 2699 1138
rect 2839 1142 2843 1143
rect 2839 1137 2843 1138
rect 2887 1142 2891 1143
rect 2887 1137 2891 1138
rect 2991 1142 2995 1143
rect 2991 1137 2995 1138
rect 3071 1142 3075 1143
rect 3071 1137 3075 1138
rect 3151 1142 3155 1143
rect 3151 1137 3155 1138
rect 3239 1142 3243 1143
rect 3239 1137 3243 1138
rect 3319 1142 3323 1143
rect 3319 1137 3323 1138
rect 3399 1142 3403 1143
rect 3399 1137 3403 1138
rect 3495 1142 3499 1143
rect 3495 1137 3499 1138
rect 3551 1142 3555 1143
rect 3551 1137 3555 1138
rect 3679 1142 3683 1143
rect 3679 1137 3683 1138
rect 3703 1142 3707 1143
rect 3703 1137 3707 1138
rect 3839 1142 3843 1143
rect 3839 1137 3843 1138
rect 3943 1142 3947 1143
rect 3943 1137 3947 1138
rect 2006 1132 2012 1133
rect 110 1128 111 1132
rect 115 1128 116 1132
rect 110 1127 116 1128
rect 174 1131 180 1132
rect 174 1127 175 1131
rect 179 1127 180 1131
rect 174 1126 180 1127
rect 326 1131 332 1132
rect 326 1127 327 1131
rect 331 1127 332 1131
rect 326 1126 332 1127
rect 494 1131 500 1132
rect 494 1127 495 1131
rect 499 1127 500 1131
rect 494 1126 500 1127
rect 670 1131 676 1132
rect 670 1127 671 1131
rect 675 1127 676 1131
rect 670 1126 676 1127
rect 846 1131 852 1132
rect 846 1127 847 1131
rect 851 1127 852 1131
rect 846 1126 852 1127
rect 1030 1131 1036 1132
rect 1030 1127 1031 1131
rect 1035 1127 1036 1131
rect 1030 1126 1036 1127
rect 1206 1131 1212 1132
rect 1206 1127 1207 1131
rect 1211 1127 1212 1131
rect 1206 1126 1212 1127
rect 1382 1131 1388 1132
rect 1382 1127 1383 1131
rect 1387 1127 1388 1131
rect 1382 1126 1388 1127
rect 1566 1131 1572 1132
rect 1566 1127 1567 1131
rect 1571 1127 1572 1131
rect 1566 1126 1572 1127
rect 1750 1131 1756 1132
rect 1750 1127 1751 1131
rect 1755 1127 1756 1131
rect 2006 1128 2007 1132
rect 2011 1128 2012 1132
rect 2006 1127 2012 1128
rect 1750 1126 1756 1127
rect 2048 1117 2050 1137
rect 2046 1116 2052 1117
rect 2296 1116 2298 1137
rect 2424 1116 2426 1137
rect 2560 1116 2562 1137
rect 2696 1116 2698 1137
rect 2840 1116 2842 1137
rect 2992 1116 2994 1137
rect 3152 1116 3154 1137
rect 3320 1116 3322 1137
rect 3496 1116 3498 1137
rect 3680 1116 3682 1137
rect 3840 1116 3842 1137
rect 3944 1117 3946 1137
rect 3942 1116 3948 1117
rect 110 1115 116 1116
rect 110 1111 111 1115
rect 115 1111 116 1115
rect 2006 1115 2012 1116
rect 110 1110 116 1111
rect 174 1112 180 1113
rect 112 1075 114 1110
rect 174 1108 175 1112
rect 179 1108 180 1112
rect 174 1107 180 1108
rect 326 1112 332 1113
rect 326 1108 327 1112
rect 331 1108 332 1112
rect 326 1107 332 1108
rect 494 1112 500 1113
rect 494 1108 495 1112
rect 499 1108 500 1112
rect 494 1107 500 1108
rect 670 1112 676 1113
rect 670 1108 671 1112
rect 675 1108 676 1112
rect 670 1107 676 1108
rect 846 1112 852 1113
rect 846 1108 847 1112
rect 851 1108 852 1112
rect 846 1107 852 1108
rect 1030 1112 1036 1113
rect 1030 1108 1031 1112
rect 1035 1108 1036 1112
rect 1030 1107 1036 1108
rect 1206 1112 1212 1113
rect 1206 1108 1207 1112
rect 1211 1108 1212 1112
rect 1206 1107 1212 1108
rect 1382 1112 1388 1113
rect 1382 1108 1383 1112
rect 1387 1108 1388 1112
rect 1382 1107 1388 1108
rect 1566 1112 1572 1113
rect 1566 1108 1567 1112
rect 1571 1108 1572 1112
rect 1566 1107 1572 1108
rect 1750 1112 1756 1113
rect 1750 1108 1751 1112
rect 1755 1108 1756 1112
rect 2006 1111 2007 1115
rect 2011 1111 2012 1115
rect 2046 1112 2047 1116
rect 2051 1112 2052 1116
rect 2046 1111 2052 1112
rect 2294 1115 2300 1116
rect 2294 1111 2295 1115
rect 2299 1111 2300 1115
rect 2006 1110 2012 1111
rect 2294 1110 2300 1111
rect 2422 1115 2428 1116
rect 2422 1111 2423 1115
rect 2427 1111 2428 1115
rect 2422 1110 2428 1111
rect 2558 1115 2564 1116
rect 2558 1111 2559 1115
rect 2563 1111 2564 1115
rect 2558 1110 2564 1111
rect 2694 1115 2700 1116
rect 2694 1111 2695 1115
rect 2699 1111 2700 1115
rect 2694 1110 2700 1111
rect 2838 1115 2844 1116
rect 2838 1111 2839 1115
rect 2843 1111 2844 1115
rect 2838 1110 2844 1111
rect 2990 1115 2996 1116
rect 2990 1111 2991 1115
rect 2995 1111 2996 1115
rect 2990 1110 2996 1111
rect 3150 1115 3156 1116
rect 3150 1111 3151 1115
rect 3155 1111 3156 1115
rect 3150 1110 3156 1111
rect 3318 1115 3324 1116
rect 3318 1111 3319 1115
rect 3323 1111 3324 1115
rect 3318 1110 3324 1111
rect 3494 1115 3500 1116
rect 3494 1111 3495 1115
rect 3499 1111 3500 1115
rect 3494 1110 3500 1111
rect 3678 1115 3684 1116
rect 3678 1111 3679 1115
rect 3683 1111 3684 1115
rect 3678 1110 3684 1111
rect 3838 1115 3844 1116
rect 3838 1111 3839 1115
rect 3843 1111 3844 1115
rect 3942 1112 3943 1116
rect 3947 1112 3948 1116
rect 3942 1111 3948 1112
rect 3838 1110 3844 1111
rect 1750 1107 1756 1108
rect 176 1075 178 1107
rect 328 1075 330 1107
rect 496 1075 498 1107
rect 672 1075 674 1107
rect 848 1075 850 1107
rect 1032 1075 1034 1107
rect 1208 1075 1210 1107
rect 1384 1075 1386 1107
rect 1568 1075 1570 1107
rect 1752 1075 1754 1107
rect 2008 1075 2010 1110
rect 2046 1099 2052 1100
rect 2046 1095 2047 1099
rect 2051 1095 2052 1099
rect 3942 1099 3948 1100
rect 2046 1094 2052 1095
rect 2294 1096 2300 1097
rect 111 1074 115 1075
rect 111 1069 115 1070
rect 135 1074 139 1075
rect 135 1069 139 1070
rect 175 1074 179 1075
rect 175 1069 179 1070
rect 231 1074 235 1075
rect 231 1069 235 1070
rect 327 1074 331 1075
rect 327 1069 331 1070
rect 375 1074 379 1075
rect 375 1069 379 1070
rect 495 1074 499 1075
rect 495 1069 499 1070
rect 543 1074 547 1075
rect 543 1069 547 1070
rect 671 1074 675 1075
rect 671 1069 675 1070
rect 727 1074 731 1075
rect 727 1069 731 1070
rect 847 1074 851 1075
rect 847 1069 851 1070
rect 911 1074 915 1075
rect 911 1069 915 1070
rect 1031 1074 1035 1075
rect 1031 1069 1035 1070
rect 1095 1074 1099 1075
rect 1095 1069 1099 1070
rect 1207 1074 1211 1075
rect 1207 1069 1211 1070
rect 1279 1074 1283 1075
rect 1279 1069 1283 1070
rect 1383 1074 1387 1075
rect 1383 1069 1387 1070
rect 1463 1074 1467 1075
rect 1463 1069 1467 1070
rect 1567 1074 1571 1075
rect 1567 1069 1571 1070
rect 1647 1074 1651 1075
rect 1647 1069 1651 1070
rect 1751 1074 1755 1075
rect 1751 1069 1755 1070
rect 1831 1074 1835 1075
rect 1831 1069 1835 1070
rect 2007 1074 2011 1075
rect 2007 1069 2011 1070
rect 112 1042 114 1069
rect 136 1045 138 1069
rect 232 1045 234 1069
rect 376 1045 378 1069
rect 544 1045 546 1069
rect 728 1045 730 1069
rect 912 1045 914 1069
rect 1096 1045 1098 1069
rect 1280 1045 1282 1069
rect 1464 1045 1466 1069
rect 1648 1045 1650 1069
rect 1832 1045 1834 1069
rect 134 1044 140 1045
rect 110 1041 116 1042
rect 110 1037 111 1041
rect 115 1037 116 1041
rect 134 1040 135 1044
rect 139 1040 140 1044
rect 134 1039 140 1040
rect 230 1044 236 1045
rect 230 1040 231 1044
rect 235 1040 236 1044
rect 230 1039 236 1040
rect 374 1044 380 1045
rect 374 1040 375 1044
rect 379 1040 380 1044
rect 374 1039 380 1040
rect 542 1044 548 1045
rect 542 1040 543 1044
rect 547 1040 548 1044
rect 542 1039 548 1040
rect 726 1044 732 1045
rect 726 1040 727 1044
rect 731 1040 732 1044
rect 726 1039 732 1040
rect 910 1044 916 1045
rect 910 1040 911 1044
rect 915 1040 916 1044
rect 910 1039 916 1040
rect 1094 1044 1100 1045
rect 1094 1040 1095 1044
rect 1099 1040 1100 1044
rect 1094 1039 1100 1040
rect 1278 1044 1284 1045
rect 1278 1040 1279 1044
rect 1283 1040 1284 1044
rect 1278 1039 1284 1040
rect 1462 1044 1468 1045
rect 1462 1040 1463 1044
rect 1467 1040 1468 1044
rect 1462 1039 1468 1040
rect 1646 1044 1652 1045
rect 1646 1040 1647 1044
rect 1651 1040 1652 1044
rect 1646 1039 1652 1040
rect 1830 1044 1836 1045
rect 1830 1040 1831 1044
rect 1835 1040 1836 1044
rect 2008 1042 2010 1069
rect 2048 1063 2050 1094
rect 2294 1092 2295 1096
rect 2299 1092 2300 1096
rect 2294 1091 2300 1092
rect 2422 1096 2428 1097
rect 2422 1092 2423 1096
rect 2427 1092 2428 1096
rect 2422 1091 2428 1092
rect 2558 1096 2564 1097
rect 2558 1092 2559 1096
rect 2563 1092 2564 1096
rect 2558 1091 2564 1092
rect 2694 1096 2700 1097
rect 2694 1092 2695 1096
rect 2699 1092 2700 1096
rect 2694 1091 2700 1092
rect 2838 1096 2844 1097
rect 2838 1092 2839 1096
rect 2843 1092 2844 1096
rect 2838 1091 2844 1092
rect 2990 1096 2996 1097
rect 2990 1092 2991 1096
rect 2995 1092 2996 1096
rect 2990 1091 2996 1092
rect 3150 1096 3156 1097
rect 3150 1092 3151 1096
rect 3155 1092 3156 1096
rect 3150 1091 3156 1092
rect 3318 1096 3324 1097
rect 3318 1092 3319 1096
rect 3323 1092 3324 1096
rect 3318 1091 3324 1092
rect 3494 1096 3500 1097
rect 3494 1092 3495 1096
rect 3499 1092 3500 1096
rect 3494 1091 3500 1092
rect 3678 1096 3684 1097
rect 3678 1092 3679 1096
rect 3683 1092 3684 1096
rect 3678 1091 3684 1092
rect 3838 1096 3844 1097
rect 3838 1092 3839 1096
rect 3843 1092 3844 1096
rect 3942 1095 3943 1099
rect 3947 1095 3948 1099
rect 3942 1094 3948 1095
rect 3838 1091 3844 1092
rect 2296 1063 2298 1091
rect 2424 1063 2426 1091
rect 2560 1063 2562 1091
rect 2696 1063 2698 1091
rect 2840 1063 2842 1091
rect 2992 1063 2994 1091
rect 3152 1063 3154 1091
rect 3320 1063 3322 1091
rect 3496 1063 3498 1091
rect 3680 1063 3682 1091
rect 3840 1063 3842 1091
rect 3944 1063 3946 1094
rect 2047 1062 2051 1063
rect 2047 1057 2051 1058
rect 2295 1062 2299 1063
rect 2295 1057 2299 1058
rect 2423 1062 2427 1063
rect 2423 1057 2427 1058
rect 2495 1062 2499 1063
rect 2495 1057 2499 1058
rect 2559 1062 2563 1063
rect 2559 1057 2563 1058
rect 2599 1062 2603 1063
rect 2599 1057 2603 1058
rect 2695 1062 2699 1063
rect 2695 1057 2699 1058
rect 2711 1062 2715 1063
rect 2711 1057 2715 1058
rect 2839 1062 2843 1063
rect 2839 1057 2843 1058
rect 2847 1062 2851 1063
rect 2847 1057 2851 1058
rect 2991 1062 2995 1063
rect 2991 1057 2995 1058
rect 3007 1062 3011 1063
rect 3007 1057 3011 1058
rect 3151 1062 3155 1063
rect 3151 1057 3155 1058
rect 3199 1062 3203 1063
rect 3199 1057 3203 1058
rect 3319 1062 3323 1063
rect 3319 1057 3323 1058
rect 3407 1062 3411 1063
rect 3407 1057 3411 1058
rect 3495 1062 3499 1063
rect 3495 1057 3499 1058
rect 3631 1062 3635 1063
rect 3631 1057 3635 1058
rect 3679 1062 3683 1063
rect 3679 1057 3683 1058
rect 3839 1062 3843 1063
rect 3839 1057 3843 1058
rect 3943 1062 3947 1063
rect 3943 1057 3947 1058
rect 1830 1039 1836 1040
rect 2006 1041 2012 1042
rect 110 1036 116 1037
rect 2006 1037 2007 1041
rect 2011 1037 2012 1041
rect 2006 1036 2012 1037
rect 2048 1030 2050 1057
rect 2496 1033 2498 1057
rect 2600 1033 2602 1057
rect 2712 1033 2714 1057
rect 2848 1033 2850 1057
rect 3008 1033 3010 1057
rect 3200 1033 3202 1057
rect 3408 1033 3410 1057
rect 3632 1033 3634 1057
rect 3840 1033 3842 1057
rect 2494 1032 2500 1033
rect 2046 1029 2052 1030
rect 134 1025 140 1026
rect 110 1024 116 1025
rect 110 1020 111 1024
rect 115 1020 116 1024
rect 134 1021 135 1025
rect 139 1021 140 1025
rect 134 1020 140 1021
rect 230 1025 236 1026
rect 230 1021 231 1025
rect 235 1021 236 1025
rect 230 1020 236 1021
rect 374 1025 380 1026
rect 374 1021 375 1025
rect 379 1021 380 1025
rect 374 1020 380 1021
rect 542 1025 548 1026
rect 542 1021 543 1025
rect 547 1021 548 1025
rect 542 1020 548 1021
rect 726 1025 732 1026
rect 726 1021 727 1025
rect 731 1021 732 1025
rect 726 1020 732 1021
rect 910 1025 916 1026
rect 910 1021 911 1025
rect 915 1021 916 1025
rect 910 1020 916 1021
rect 1094 1025 1100 1026
rect 1094 1021 1095 1025
rect 1099 1021 1100 1025
rect 1094 1020 1100 1021
rect 1278 1025 1284 1026
rect 1278 1021 1279 1025
rect 1283 1021 1284 1025
rect 1278 1020 1284 1021
rect 1462 1025 1468 1026
rect 1462 1021 1463 1025
rect 1467 1021 1468 1025
rect 1462 1020 1468 1021
rect 1646 1025 1652 1026
rect 1646 1021 1647 1025
rect 1651 1021 1652 1025
rect 1646 1020 1652 1021
rect 1830 1025 1836 1026
rect 2046 1025 2047 1029
rect 2051 1025 2052 1029
rect 2494 1028 2495 1032
rect 2499 1028 2500 1032
rect 2494 1027 2500 1028
rect 2598 1032 2604 1033
rect 2598 1028 2599 1032
rect 2603 1028 2604 1032
rect 2598 1027 2604 1028
rect 2710 1032 2716 1033
rect 2710 1028 2711 1032
rect 2715 1028 2716 1032
rect 2710 1027 2716 1028
rect 2846 1032 2852 1033
rect 2846 1028 2847 1032
rect 2851 1028 2852 1032
rect 2846 1027 2852 1028
rect 3006 1032 3012 1033
rect 3006 1028 3007 1032
rect 3011 1028 3012 1032
rect 3006 1027 3012 1028
rect 3198 1032 3204 1033
rect 3198 1028 3199 1032
rect 3203 1028 3204 1032
rect 3198 1027 3204 1028
rect 3406 1032 3412 1033
rect 3406 1028 3407 1032
rect 3411 1028 3412 1032
rect 3406 1027 3412 1028
rect 3630 1032 3636 1033
rect 3630 1028 3631 1032
rect 3635 1028 3636 1032
rect 3630 1027 3636 1028
rect 3838 1032 3844 1033
rect 3838 1028 3839 1032
rect 3843 1028 3844 1032
rect 3944 1030 3946 1057
rect 3838 1027 3844 1028
rect 3942 1029 3948 1030
rect 1830 1021 1831 1025
rect 1835 1021 1836 1025
rect 1830 1020 1836 1021
rect 2006 1024 2012 1025
rect 2046 1024 2052 1025
rect 3942 1025 3943 1029
rect 3947 1025 3948 1029
rect 3942 1024 3948 1025
rect 2006 1020 2007 1024
rect 2011 1020 2012 1024
rect 110 1019 116 1020
rect 112 999 114 1019
rect 136 999 138 1020
rect 232 999 234 1020
rect 376 999 378 1020
rect 544 999 546 1020
rect 728 999 730 1020
rect 912 999 914 1020
rect 1096 999 1098 1020
rect 1280 999 1282 1020
rect 1464 999 1466 1020
rect 1648 999 1650 1020
rect 1832 999 1834 1020
rect 2006 1019 2012 1020
rect 2008 999 2010 1019
rect 2494 1013 2500 1014
rect 2046 1012 2052 1013
rect 2046 1008 2047 1012
rect 2051 1008 2052 1012
rect 2494 1009 2495 1013
rect 2499 1009 2500 1013
rect 2494 1008 2500 1009
rect 2598 1013 2604 1014
rect 2598 1009 2599 1013
rect 2603 1009 2604 1013
rect 2598 1008 2604 1009
rect 2710 1013 2716 1014
rect 2710 1009 2711 1013
rect 2715 1009 2716 1013
rect 2710 1008 2716 1009
rect 2846 1013 2852 1014
rect 2846 1009 2847 1013
rect 2851 1009 2852 1013
rect 2846 1008 2852 1009
rect 3006 1013 3012 1014
rect 3006 1009 3007 1013
rect 3011 1009 3012 1013
rect 3006 1008 3012 1009
rect 3198 1013 3204 1014
rect 3198 1009 3199 1013
rect 3203 1009 3204 1013
rect 3198 1008 3204 1009
rect 3406 1013 3412 1014
rect 3406 1009 3407 1013
rect 3411 1009 3412 1013
rect 3406 1008 3412 1009
rect 3630 1013 3636 1014
rect 3630 1009 3631 1013
rect 3635 1009 3636 1013
rect 3630 1008 3636 1009
rect 3838 1013 3844 1014
rect 3838 1009 3839 1013
rect 3843 1009 3844 1013
rect 3838 1008 3844 1009
rect 3942 1012 3948 1013
rect 3942 1008 3943 1012
rect 3947 1008 3948 1012
rect 2046 1007 2052 1008
rect 111 998 115 999
rect 111 993 115 994
rect 135 998 139 999
rect 135 993 139 994
rect 231 998 235 999
rect 231 993 235 994
rect 271 998 275 999
rect 271 993 275 994
rect 375 998 379 999
rect 375 993 379 994
rect 447 998 451 999
rect 447 993 451 994
rect 543 998 547 999
rect 543 993 547 994
rect 631 998 635 999
rect 631 993 635 994
rect 727 998 731 999
rect 727 993 731 994
rect 823 998 827 999
rect 823 993 827 994
rect 911 998 915 999
rect 911 993 915 994
rect 1007 998 1011 999
rect 1007 993 1011 994
rect 1095 998 1099 999
rect 1095 993 1099 994
rect 1175 998 1179 999
rect 1175 993 1179 994
rect 1279 998 1283 999
rect 1279 993 1283 994
rect 1335 998 1339 999
rect 1335 993 1339 994
rect 1463 998 1467 999
rect 1463 993 1467 994
rect 1487 998 1491 999
rect 1487 993 1491 994
rect 1631 998 1635 999
rect 1631 993 1635 994
rect 1647 998 1651 999
rect 1647 993 1651 994
rect 1775 998 1779 999
rect 1775 993 1779 994
rect 1831 998 1835 999
rect 1831 993 1835 994
rect 1903 998 1907 999
rect 1903 993 1907 994
rect 2007 998 2011 999
rect 2007 993 2011 994
rect 112 973 114 993
rect 110 972 116 973
rect 136 972 138 993
rect 272 972 274 993
rect 448 972 450 993
rect 632 972 634 993
rect 824 972 826 993
rect 1008 972 1010 993
rect 1176 972 1178 993
rect 1336 972 1338 993
rect 1488 972 1490 993
rect 1632 972 1634 993
rect 1776 972 1778 993
rect 1904 972 1906 993
rect 2008 973 2010 993
rect 2048 987 2050 1007
rect 2496 987 2498 1008
rect 2600 987 2602 1008
rect 2712 987 2714 1008
rect 2848 987 2850 1008
rect 3008 987 3010 1008
rect 3200 987 3202 1008
rect 3408 987 3410 1008
rect 3632 987 3634 1008
rect 3840 987 3842 1008
rect 3942 1007 3948 1008
rect 3944 987 3946 1007
rect 2047 986 2051 987
rect 2047 981 2051 982
rect 2495 986 2499 987
rect 2495 981 2499 982
rect 2599 986 2603 987
rect 2599 981 2603 982
rect 2647 986 2651 987
rect 2647 981 2651 982
rect 2711 986 2715 987
rect 2711 981 2715 982
rect 2743 986 2747 987
rect 2743 981 2747 982
rect 2847 986 2851 987
rect 2847 981 2851 982
rect 2967 986 2971 987
rect 2967 981 2971 982
rect 3007 986 3011 987
rect 3007 981 3011 982
rect 3111 986 3115 987
rect 3111 981 3115 982
rect 3199 986 3203 987
rect 3199 981 3203 982
rect 3279 986 3283 987
rect 3279 981 3283 982
rect 3407 986 3411 987
rect 3407 981 3411 982
rect 3463 986 3467 987
rect 3463 981 3467 982
rect 3631 986 3635 987
rect 3631 981 3635 982
rect 3663 986 3667 987
rect 3663 981 3667 982
rect 3839 986 3843 987
rect 3839 981 3843 982
rect 3943 986 3947 987
rect 3943 981 3947 982
rect 2006 972 2012 973
rect 110 968 111 972
rect 115 968 116 972
rect 110 967 116 968
rect 134 971 140 972
rect 134 967 135 971
rect 139 967 140 971
rect 134 966 140 967
rect 270 971 276 972
rect 270 967 271 971
rect 275 967 276 971
rect 270 966 276 967
rect 446 971 452 972
rect 446 967 447 971
rect 451 967 452 971
rect 446 966 452 967
rect 630 971 636 972
rect 630 967 631 971
rect 635 967 636 971
rect 630 966 636 967
rect 822 971 828 972
rect 822 967 823 971
rect 827 967 828 971
rect 822 966 828 967
rect 1006 971 1012 972
rect 1006 967 1007 971
rect 1011 967 1012 971
rect 1006 966 1012 967
rect 1174 971 1180 972
rect 1174 967 1175 971
rect 1179 967 1180 971
rect 1174 966 1180 967
rect 1334 971 1340 972
rect 1334 967 1335 971
rect 1339 967 1340 971
rect 1334 966 1340 967
rect 1486 971 1492 972
rect 1486 967 1487 971
rect 1491 967 1492 971
rect 1486 966 1492 967
rect 1630 971 1636 972
rect 1630 967 1631 971
rect 1635 967 1636 971
rect 1630 966 1636 967
rect 1774 971 1780 972
rect 1774 967 1775 971
rect 1779 967 1780 971
rect 1774 966 1780 967
rect 1902 971 1908 972
rect 1902 967 1903 971
rect 1907 967 1908 971
rect 2006 968 2007 972
rect 2011 968 2012 972
rect 2006 967 2012 968
rect 1902 966 1908 967
rect 2048 961 2050 981
rect 2046 960 2052 961
rect 2648 960 2650 981
rect 2744 960 2746 981
rect 2848 960 2850 981
rect 2968 960 2970 981
rect 3112 960 3114 981
rect 3280 960 3282 981
rect 3464 960 3466 981
rect 3664 960 3666 981
rect 3840 960 3842 981
rect 3944 961 3946 981
rect 3942 960 3948 961
rect 2046 956 2047 960
rect 2051 956 2052 960
rect 110 955 116 956
rect 110 951 111 955
rect 115 951 116 955
rect 2006 955 2012 956
rect 2046 955 2052 956
rect 2646 959 2652 960
rect 2646 955 2647 959
rect 2651 955 2652 959
rect 110 950 116 951
rect 134 952 140 953
rect 112 923 114 950
rect 134 948 135 952
rect 139 948 140 952
rect 134 947 140 948
rect 270 952 276 953
rect 270 948 271 952
rect 275 948 276 952
rect 270 947 276 948
rect 446 952 452 953
rect 446 948 447 952
rect 451 948 452 952
rect 446 947 452 948
rect 630 952 636 953
rect 630 948 631 952
rect 635 948 636 952
rect 630 947 636 948
rect 822 952 828 953
rect 822 948 823 952
rect 827 948 828 952
rect 822 947 828 948
rect 1006 952 1012 953
rect 1006 948 1007 952
rect 1011 948 1012 952
rect 1006 947 1012 948
rect 1174 952 1180 953
rect 1174 948 1175 952
rect 1179 948 1180 952
rect 1174 947 1180 948
rect 1334 952 1340 953
rect 1334 948 1335 952
rect 1339 948 1340 952
rect 1334 947 1340 948
rect 1486 952 1492 953
rect 1486 948 1487 952
rect 1491 948 1492 952
rect 1486 947 1492 948
rect 1630 952 1636 953
rect 1630 948 1631 952
rect 1635 948 1636 952
rect 1630 947 1636 948
rect 1774 952 1780 953
rect 1774 948 1775 952
rect 1779 948 1780 952
rect 1774 947 1780 948
rect 1902 952 1908 953
rect 1902 948 1903 952
rect 1907 948 1908 952
rect 2006 951 2007 955
rect 2011 951 2012 955
rect 2646 954 2652 955
rect 2742 959 2748 960
rect 2742 955 2743 959
rect 2747 955 2748 959
rect 2742 954 2748 955
rect 2846 959 2852 960
rect 2846 955 2847 959
rect 2851 955 2852 959
rect 2846 954 2852 955
rect 2966 959 2972 960
rect 2966 955 2967 959
rect 2971 955 2972 959
rect 2966 954 2972 955
rect 3110 959 3116 960
rect 3110 955 3111 959
rect 3115 955 3116 959
rect 3110 954 3116 955
rect 3278 959 3284 960
rect 3278 955 3279 959
rect 3283 955 3284 959
rect 3278 954 3284 955
rect 3462 959 3468 960
rect 3462 955 3463 959
rect 3467 955 3468 959
rect 3462 954 3468 955
rect 3662 959 3668 960
rect 3662 955 3663 959
rect 3667 955 3668 959
rect 3662 954 3668 955
rect 3838 959 3844 960
rect 3838 955 3839 959
rect 3843 955 3844 959
rect 3942 956 3943 960
rect 3947 956 3948 960
rect 3942 955 3948 956
rect 3838 954 3844 955
rect 2006 950 2012 951
rect 1902 947 1908 948
rect 136 923 138 947
rect 272 923 274 947
rect 448 923 450 947
rect 632 923 634 947
rect 824 923 826 947
rect 1008 923 1010 947
rect 1176 923 1178 947
rect 1336 923 1338 947
rect 1488 923 1490 947
rect 1632 923 1634 947
rect 1776 923 1778 947
rect 1904 923 1906 947
rect 2008 923 2010 950
rect 2046 943 2052 944
rect 2046 939 2047 943
rect 2051 939 2052 943
rect 3942 943 3948 944
rect 2046 938 2052 939
rect 2646 940 2652 941
rect 111 922 115 923
rect 111 917 115 918
rect 135 922 139 923
rect 135 917 139 918
rect 271 922 275 923
rect 271 917 275 918
rect 447 922 451 923
rect 447 917 451 918
rect 455 922 459 923
rect 455 917 459 918
rect 631 922 635 923
rect 631 917 635 918
rect 655 922 659 923
rect 655 917 659 918
rect 823 922 827 923
rect 823 917 827 918
rect 855 922 859 923
rect 855 917 859 918
rect 1007 922 1011 923
rect 1007 917 1011 918
rect 1055 922 1059 923
rect 1055 917 1059 918
rect 1175 922 1179 923
rect 1175 917 1179 918
rect 1239 922 1243 923
rect 1239 917 1243 918
rect 1335 922 1339 923
rect 1335 917 1339 918
rect 1415 922 1419 923
rect 1415 917 1419 918
rect 1487 922 1491 923
rect 1487 917 1491 918
rect 1583 922 1587 923
rect 1583 917 1587 918
rect 1631 922 1635 923
rect 1631 917 1635 918
rect 1751 922 1755 923
rect 1751 917 1755 918
rect 1775 922 1779 923
rect 1775 917 1779 918
rect 1903 922 1907 923
rect 1903 917 1907 918
rect 2007 922 2011 923
rect 2007 917 2011 918
rect 112 890 114 917
rect 136 893 138 917
rect 272 893 274 917
rect 456 893 458 917
rect 656 893 658 917
rect 856 893 858 917
rect 1056 893 1058 917
rect 1240 893 1242 917
rect 1416 893 1418 917
rect 1584 893 1586 917
rect 1752 893 1754 917
rect 1904 893 1906 917
rect 134 892 140 893
rect 110 889 116 890
rect 110 885 111 889
rect 115 885 116 889
rect 134 888 135 892
rect 139 888 140 892
rect 134 887 140 888
rect 270 892 276 893
rect 270 888 271 892
rect 275 888 276 892
rect 270 887 276 888
rect 454 892 460 893
rect 454 888 455 892
rect 459 888 460 892
rect 454 887 460 888
rect 654 892 660 893
rect 654 888 655 892
rect 659 888 660 892
rect 654 887 660 888
rect 854 892 860 893
rect 854 888 855 892
rect 859 888 860 892
rect 854 887 860 888
rect 1054 892 1060 893
rect 1054 888 1055 892
rect 1059 888 1060 892
rect 1054 887 1060 888
rect 1238 892 1244 893
rect 1238 888 1239 892
rect 1243 888 1244 892
rect 1238 887 1244 888
rect 1414 892 1420 893
rect 1414 888 1415 892
rect 1419 888 1420 892
rect 1414 887 1420 888
rect 1582 892 1588 893
rect 1582 888 1583 892
rect 1587 888 1588 892
rect 1582 887 1588 888
rect 1750 892 1756 893
rect 1750 888 1751 892
rect 1755 888 1756 892
rect 1750 887 1756 888
rect 1902 892 1908 893
rect 1902 888 1903 892
rect 1907 888 1908 892
rect 2008 890 2010 917
rect 2048 899 2050 938
rect 2646 936 2647 940
rect 2651 936 2652 940
rect 2646 935 2652 936
rect 2742 940 2748 941
rect 2742 936 2743 940
rect 2747 936 2748 940
rect 2742 935 2748 936
rect 2846 940 2852 941
rect 2846 936 2847 940
rect 2851 936 2852 940
rect 2846 935 2852 936
rect 2966 940 2972 941
rect 2966 936 2967 940
rect 2971 936 2972 940
rect 2966 935 2972 936
rect 3110 940 3116 941
rect 3110 936 3111 940
rect 3115 936 3116 940
rect 3110 935 3116 936
rect 3278 940 3284 941
rect 3278 936 3279 940
rect 3283 936 3284 940
rect 3278 935 3284 936
rect 3462 940 3468 941
rect 3462 936 3463 940
rect 3467 936 3468 940
rect 3462 935 3468 936
rect 3662 940 3668 941
rect 3662 936 3663 940
rect 3667 936 3668 940
rect 3662 935 3668 936
rect 3838 940 3844 941
rect 3838 936 3839 940
rect 3843 936 3844 940
rect 3942 939 3943 943
rect 3947 939 3948 943
rect 3942 938 3948 939
rect 3838 935 3844 936
rect 2648 899 2650 935
rect 2744 899 2746 935
rect 2848 899 2850 935
rect 2968 899 2970 935
rect 3112 899 3114 935
rect 3280 899 3282 935
rect 3464 899 3466 935
rect 3664 899 3666 935
rect 3840 899 3842 935
rect 3944 899 3946 938
rect 2047 898 2051 899
rect 2047 893 2051 894
rect 2071 898 2075 899
rect 2071 893 2075 894
rect 2255 898 2259 899
rect 2255 893 2259 894
rect 2463 898 2467 899
rect 2463 893 2467 894
rect 2647 898 2651 899
rect 2647 893 2651 894
rect 2679 898 2683 899
rect 2679 893 2683 894
rect 2743 898 2747 899
rect 2743 893 2747 894
rect 2847 898 2851 899
rect 2847 893 2851 894
rect 2895 898 2899 899
rect 2895 893 2899 894
rect 2967 898 2971 899
rect 2967 893 2971 894
rect 3111 898 3115 899
rect 3111 893 3115 894
rect 3127 898 3131 899
rect 3127 893 3131 894
rect 3279 898 3283 899
rect 3279 893 3283 894
rect 3367 898 3371 899
rect 3367 893 3371 894
rect 3463 898 3467 899
rect 3463 893 3467 894
rect 3615 898 3619 899
rect 3615 893 3619 894
rect 3663 898 3667 899
rect 3663 893 3667 894
rect 3839 898 3843 899
rect 3839 893 3843 894
rect 3943 898 3947 899
rect 3943 893 3947 894
rect 1902 887 1908 888
rect 2006 889 2012 890
rect 110 884 116 885
rect 2006 885 2007 889
rect 2011 885 2012 889
rect 2006 884 2012 885
rect 134 873 140 874
rect 110 872 116 873
rect 110 868 111 872
rect 115 868 116 872
rect 134 869 135 873
rect 139 869 140 873
rect 134 868 140 869
rect 270 873 276 874
rect 270 869 271 873
rect 275 869 276 873
rect 270 868 276 869
rect 454 873 460 874
rect 454 869 455 873
rect 459 869 460 873
rect 454 868 460 869
rect 654 873 660 874
rect 654 869 655 873
rect 659 869 660 873
rect 654 868 660 869
rect 854 873 860 874
rect 854 869 855 873
rect 859 869 860 873
rect 854 868 860 869
rect 1054 873 1060 874
rect 1054 869 1055 873
rect 1059 869 1060 873
rect 1054 868 1060 869
rect 1238 873 1244 874
rect 1238 869 1239 873
rect 1243 869 1244 873
rect 1238 868 1244 869
rect 1414 873 1420 874
rect 1414 869 1415 873
rect 1419 869 1420 873
rect 1414 868 1420 869
rect 1582 873 1588 874
rect 1582 869 1583 873
rect 1587 869 1588 873
rect 1582 868 1588 869
rect 1750 873 1756 874
rect 1750 869 1751 873
rect 1755 869 1756 873
rect 1750 868 1756 869
rect 1902 873 1908 874
rect 1902 869 1903 873
rect 1907 869 1908 873
rect 1902 868 1908 869
rect 2006 872 2012 873
rect 2006 868 2007 872
rect 2011 868 2012 872
rect 110 867 116 868
rect 112 847 114 867
rect 136 847 138 868
rect 272 847 274 868
rect 456 847 458 868
rect 656 847 658 868
rect 856 847 858 868
rect 1056 847 1058 868
rect 1240 847 1242 868
rect 1416 847 1418 868
rect 1584 847 1586 868
rect 1752 847 1754 868
rect 1904 847 1906 868
rect 2006 867 2012 868
rect 2008 847 2010 867
rect 2048 866 2050 893
rect 2072 869 2074 893
rect 2256 869 2258 893
rect 2464 869 2466 893
rect 2680 869 2682 893
rect 2896 869 2898 893
rect 3128 869 3130 893
rect 3368 869 3370 893
rect 3616 869 3618 893
rect 3840 869 3842 893
rect 2070 868 2076 869
rect 2046 865 2052 866
rect 2046 861 2047 865
rect 2051 861 2052 865
rect 2070 864 2071 868
rect 2075 864 2076 868
rect 2070 863 2076 864
rect 2254 868 2260 869
rect 2254 864 2255 868
rect 2259 864 2260 868
rect 2254 863 2260 864
rect 2462 868 2468 869
rect 2462 864 2463 868
rect 2467 864 2468 868
rect 2462 863 2468 864
rect 2678 868 2684 869
rect 2678 864 2679 868
rect 2683 864 2684 868
rect 2678 863 2684 864
rect 2894 868 2900 869
rect 2894 864 2895 868
rect 2899 864 2900 868
rect 2894 863 2900 864
rect 3126 868 3132 869
rect 3126 864 3127 868
rect 3131 864 3132 868
rect 3126 863 3132 864
rect 3366 868 3372 869
rect 3366 864 3367 868
rect 3371 864 3372 868
rect 3366 863 3372 864
rect 3614 868 3620 869
rect 3614 864 3615 868
rect 3619 864 3620 868
rect 3614 863 3620 864
rect 3838 868 3844 869
rect 3838 864 3839 868
rect 3843 864 3844 868
rect 3944 866 3946 893
rect 3838 863 3844 864
rect 3942 865 3948 866
rect 2046 860 2052 861
rect 3942 861 3943 865
rect 3947 861 3948 865
rect 3942 860 3948 861
rect 2070 849 2076 850
rect 2046 848 2052 849
rect 111 846 115 847
rect 111 841 115 842
rect 135 846 139 847
rect 135 841 139 842
rect 215 846 219 847
rect 215 841 219 842
rect 271 846 275 847
rect 271 841 275 842
rect 343 846 347 847
rect 343 841 347 842
rect 455 846 459 847
rect 455 841 459 842
rect 495 846 499 847
rect 495 841 499 842
rect 655 846 659 847
rect 655 841 659 842
rect 831 846 835 847
rect 831 841 835 842
rect 855 846 859 847
rect 855 841 859 842
rect 1007 846 1011 847
rect 1007 841 1011 842
rect 1055 846 1059 847
rect 1055 841 1059 842
rect 1183 846 1187 847
rect 1183 841 1187 842
rect 1239 846 1243 847
rect 1239 841 1243 842
rect 1359 846 1363 847
rect 1359 841 1363 842
rect 1415 846 1419 847
rect 1415 841 1419 842
rect 1535 846 1539 847
rect 1535 841 1539 842
rect 1583 846 1587 847
rect 1583 841 1587 842
rect 1719 846 1723 847
rect 1719 841 1723 842
rect 1751 846 1755 847
rect 1751 841 1755 842
rect 1903 846 1907 847
rect 1903 841 1907 842
rect 2007 846 2011 847
rect 2046 844 2047 848
rect 2051 844 2052 848
rect 2070 845 2071 849
rect 2075 845 2076 849
rect 2070 844 2076 845
rect 2254 849 2260 850
rect 2254 845 2255 849
rect 2259 845 2260 849
rect 2254 844 2260 845
rect 2462 849 2468 850
rect 2462 845 2463 849
rect 2467 845 2468 849
rect 2462 844 2468 845
rect 2678 849 2684 850
rect 2678 845 2679 849
rect 2683 845 2684 849
rect 2678 844 2684 845
rect 2894 849 2900 850
rect 2894 845 2895 849
rect 2899 845 2900 849
rect 2894 844 2900 845
rect 3126 849 3132 850
rect 3126 845 3127 849
rect 3131 845 3132 849
rect 3126 844 3132 845
rect 3366 849 3372 850
rect 3366 845 3367 849
rect 3371 845 3372 849
rect 3366 844 3372 845
rect 3614 849 3620 850
rect 3614 845 3615 849
rect 3619 845 3620 849
rect 3614 844 3620 845
rect 3838 849 3844 850
rect 3838 845 3839 849
rect 3843 845 3844 849
rect 3838 844 3844 845
rect 3942 848 3948 849
rect 3942 844 3943 848
rect 3947 844 3948 848
rect 2046 843 2052 844
rect 2007 841 2011 842
rect 112 821 114 841
rect 110 820 116 821
rect 216 820 218 841
rect 344 820 346 841
rect 496 820 498 841
rect 656 820 658 841
rect 832 820 834 841
rect 1008 820 1010 841
rect 1184 820 1186 841
rect 1360 820 1362 841
rect 1536 820 1538 841
rect 1720 820 1722 841
rect 2008 821 2010 841
rect 2048 823 2050 843
rect 2072 823 2074 844
rect 2256 823 2258 844
rect 2464 823 2466 844
rect 2680 823 2682 844
rect 2896 823 2898 844
rect 3128 823 3130 844
rect 3368 823 3370 844
rect 3616 823 3618 844
rect 3840 823 3842 844
rect 3942 843 3948 844
rect 3944 823 3946 843
rect 2047 822 2051 823
rect 2006 820 2012 821
rect 110 816 111 820
rect 115 816 116 820
rect 110 815 116 816
rect 214 819 220 820
rect 214 815 215 819
rect 219 815 220 819
rect 214 814 220 815
rect 342 819 348 820
rect 342 815 343 819
rect 347 815 348 819
rect 342 814 348 815
rect 494 819 500 820
rect 494 815 495 819
rect 499 815 500 819
rect 494 814 500 815
rect 654 819 660 820
rect 654 815 655 819
rect 659 815 660 819
rect 654 814 660 815
rect 830 819 836 820
rect 830 815 831 819
rect 835 815 836 819
rect 830 814 836 815
rect 1006 819 1012 820
rect 1006 815 1007 819
rect 1011 815 1012 819
rect 1006 814 1012 815
rect 1182 819 1188 820
rect 1182 815 1183 819
rect 1187 815 1188 819
rect 1182 814 1188 815
rect 1358 819 1364 820
rect 1358 815 1359 819
rect 1363 815 1364 819
rect 1358 814 1364 815
rect 1534 819 1540 820
rect 1534 815 1535 819
rect 1539 815 1540 819
rect 1534 814 1540 815
rect 1718 819 1724 820
rect 1718 815 1719 819
rect 1723 815 1724 819
rect 2006 816 2007 820
rect 2011 816 2012 820
rect 2047 817 2051 818
rect 2071 822 2075 823
rect 2071 817 2075 818
rect 2215 822 2219 823
rect 2215 817 2219 818
rect 2255 822 2259 823
rect 2255 817 2259 818
rect 2327 822 2331 823
rect 2327 817 2331 818
rect 2447 822 2451 823
rect 2447 817 2451 818
rect 2463 822 2467 823
rect 2463 817 2467 818
rect 2583 822 2587 823
rect 2583 817 2587 818
rect 2679 822 2683 823
rect 2679 817 2683 818
rect 2735 822 2739 823
rect 2735 817 2739 818
rect 2895 822 2899 823
rect 2895 817 2899 818
rect 3063 822 3067 823
rect 3063 817 3067 818
rect 3127 822 3131 823
rect 3127 817 3131 818
rect 3247 822 3251 823
rect 3247 817 3251 818
rect 3367 822 3371 823
rect 3367 817 3371 818
rect 3447 822 3451 823
rect 3447 817 3451 818
rect 3615 822 3619 823
rect 3615 817 3619 818
rect 3655 822 3659 823
rect 3655 817 3659 818
rect 3839 822 3843 823
rect 3839 817 3843 818
rect 3943 822 3947 823
rect 3943 817 3947 818
rect 2006 815 2012 816
rect 1718 814 1724 815
rect 110 803 116 804
rect 110 799 111 803
rect 115 799 116 803
rect 2006 803 2012 804
rect 110 798 116 799
rect 214 800 220 801
rect 112 771 114 798
rect 214 796 215 800
rect 219 796 220 800
rect 214 795 220 796
rect 342 800 348 801
rect 342 796 343 800
rect 347 796 348 800
rect 342 795 348 796
rect 494 800 500 801
rect 494 796 495 800
rect 499 796 500 800
rect 494 795 500 796
rect 654 800 660 801
rect 654 796 655 800
rect 659 796 660 800
rect 654 795 660 796
rect 830 800 836 801
rect 830 796 831 800
rect 835 796 836 800
rect 830 795 836 796
rect 1006 800 1012 801
rect 1006 796 1007 800
rect 1011 796 1012 800
rect 1006 795 1012 796
rect 1182 800 1188 801
rect 1182 796 1183 800
rect 1187 796 1188 800
rect 1182 795 1188 796
rect 1358 800 1364 801
rect 1358 796 1359 800
rect 1363 796 1364 800
rect 1358 795 1364 796
rect 1534 800 1540 801
rect 1534 796 1535 800
rect 1539 796 1540 800
rect 1534 795 1540 796
rect 1718 800 1724 801
rect 1718 796 1719 800
rect 1723 796 1724 800
rect 2006 799 2007 803
rect 2011 799 2012 803
rect 2006 798 2012 799
rect 1718 795 1724 796
rect 216 771 218 795
rect 344 771 346 795
rect 496 771 498 795
rect 656 771 658 795
rect 832 771 834 795
rect 1008 771 1010 795
rect 1184 771 1186 795
rect 1360 771 1362 795
rect 1536 771 1538 795
rect 1720 771 1722 795
rect 2008 771 2010 798
rect 2048 797 2050 817
rect 2046 796 2052 797
rect 2216 796 2218 817
rect 2328 796 2330 817
rect 2448 796 2450 817
rect 2584 796 2586 817
rect 2736 796 2738 817
rect 2896 796 2898 817
rect 3064 796 3066 817
rect 3248 796 3250 817
rect 3448 796 3450 817
rect 3656 796 3658 817
rect 3840 796 3842 817
rect 3944 797 3946 817
rect 3942 796 3948 797
rect 2046 792 2047 796
rect 2051 792 2052 796
rect 2046 791 2052 792
rect 2214 795 2220 796
rect 2214 791 2215 795
rect 2219 791 2220 795
rect 2214 790 2220 791
rect 2326 795 2332 796
rect 2326 791 2327 795
rect 2331 791 2332 795
rect 2326 790 2332 791
rect 2446 795 2452 796
rect 2446 791 2447 795
rect 2451 791 2452 795
rect 2446 790 2452 791
rect 2582 795 2588 796
rect 2582 791 2583 795
rect 2587 791 2588 795
rect 2582 790 2588 791
rect 2734 795 2740 796
rect 2734 791 2735 795
rect 2739 791 2740 795
rect 2734 790 2740 791
rect 2894 795 2900 796
rect 2894 791 2895 795
rect 2899 791 2900 795
rect 2894 790 2900 791
rect 3062 795 3068 796
rect 3062 791 3063 795
rect 3067 791 3068 795
rect 3062 790 3068 791
rect 3246 795 3252 796
rect 3246 791 3247 795
rect 3251 791 3252 795
rect 3246 790 3252 791
rect 3446 795 3452 796
rect 3446 791 3447 795
rect 3451 791 3452 795
rect 3446 790 3452 791
rect 3654 795 3660 796
rect 3654 791 3655 795
rect 3659 791 3660 795
rect 3654 790 3660 791
rect 3838 795 3844 796
rect 3838 791 3839 795
rect 3843 791 3844 795
rect 3942 792 3943 796
rect 3947 792 3948 796
rect 3942 791 3948 792
rect 3838 790 3844 791
rect 2046 779 2052 780
rect 2046 775 2047 779
rect 2051 775 2052 779
rect 3942 779 3948 780
rect 2046 774 2052 775
rect 2214 776 2220 777
rect 111 770 115 771
rect 111 765 115 766
rect 215 770 219 771
rect 215 765 219 766
rect 343 770 347 771
rect 343 765 347 766
rect 375 770 379 771
rect 375 765 379 766
rect 495 770 499 771
rect 495 765 499 766
rect 623 770 627 771
rect 623 765 627 766
rect 655 770 659 771
rect 655 765 659 766
rect 751 770 755 771
rect 751 765 755 766
rect 831 770 835 771
rect 831 765 835 766
rect 887 770 891 771
rect 887 765 891 766
rect 1007 770 1011 771
rect 1007 765 1011 766
rect 1023 770 1027 771
rect 1023 765 1027 766
rect 1167 770 1171 771
rect 1167 765 1171 766
rect 1183 770 1187 771
rect 1183 765 1187 766
rect 1311 770 1315 771
rect 1311 765 1315 766
rect 1359 770 1363 771
rect 1359 765 1363 766
rect 1455 770 1459 771
rect 1455 765 1459 766
rect 1535 770 1539 771
rect 1535 765 1539 766
rect 1599 770 1603 771
rect 1599 765 1603 766
rect 1719 770 1723 771
rect 1719 765 1723 766
rect 2007 770 2011 771
rect 2007 765 2011 766
rect 112 738 114 765
rect 376 741 378 765
rect 496 741 498 765
rect 624 741 626 765
rect 752 741 754 765
rect 888 741 890 765
rect 1024 741 1026 765
rect 1168 741 1170 765
rect 1312 741 1314 765
rect 1456 741 1458 765
rect 1600 741 1602 765
rect 374 740 380 741
rect 110 737 116 738
rect 110 733 111 737
rect 115 733 116 737
rect 374 736 375 740
rect 379 736 380 740
rect 374 735 380 736
rect 494 740 500 741
rect 494 736 495 740
rect 499 736 500 740
rect 494 735 500 736
rect 622 740 628 741
rect 622 736 623 740
rect 627 736 628 740
rect 622 735 628 736
rect 750 740 756 741
rect 750 736 751 740
rect 755 736 756 740
rect 750 735 756 736
rect 886 740 892 741
rect 886 736 887 740
rect 891 736 892 740
rect 886 735 892 736
rect 1022 740 1028 741
rect 1022 736 1023 740
rect 1027 736 1028 740
rect 1022 735 1028 736
rect 1166 740 1172 741
rect 1166 736 1167 740
rect 1171 736 1172 740
rect 1166 735 1172 736
rect 1310 740 1316 741
rect 1310 736 1311 740
rect 1315 736 1316 740
rect 1310 735 1316 736
rect 1454 740 1460 741
rect 1454 736 1455 740
rect 1459 736 1460 740
rect 1454 735 1460 736
rect 1598 740 1604 741
rect 1598 736 1599 740
rect 1603 736 1604 740
rect 2008 738 2010 765
rect 2048 743 2050 774
rect 2214 772 2215 776
rect 2219 772 2220 776
rect 2214 771 2220 772
rect 2326 776 2332 777
rect 2326 772 2327 776
rect 2331 772 2332 776
rect 2326 771 2332 772
rect 2446 776 2452 777
rect 2446 772 2447 776
rect 2451 772 2452 776
rect 2446 771 2452 772
rect 2582 776 2588 777
rect 2582 772 2583 776
rect 2587 772 2588 776
rect 2582 771 2588 772
rect 2734 776 2740 777
rect 2734 772 2735 776
rect 2739 772 2740 776
rect 2734 771 2740 772
rect 2894 776 2900 777
rect 2894 772 2895 776
rect 2899 772 2900 776
rect 2894 771 2900 772
rect 3062 776 3068 777
rect 3062 772 3063 776
rect 3067 772 3068 776
rect 3062 771 3068 772
rect 3246 776 3252 777
rect 3246 772 3247 776
rect 3251 772 3252 776
rect 3246 771 3252 772
rect 3446 776 3452 777
rect 3446 772 3447 776
rect 3451 772 3452 776
rect 3446 771 3452 772
rect 3654 776 3660 777
rect 3654 772 3655 776
rect 3659 772 3660 776
rect 3654 771 3660 772
rect 3838 776 3844 777
rect 3838 772 3839 776
rect 3843 772 3844 776
rect 3942 775 3943 779
rect 3947 775 3948 779
rect 3942 774 3948 775
rect 3838 771 3844 772
rect 2216 743 2218 771
rect 2328 743 2330 771
rect 2448 743 2450 771
rect 2584 743 2586 771
rect 2736 743 2738 771
rect 2896 743 2898 771
rect 3064 743 3066 771
rect 3248 743 3250 771
rect 3448 743 3450 771
rect 3656 743 3658 771
rect 3840 743 3842 771
rect 3944 743 3946 774
rect 2047 742 2051 743
rect 1598 735 1604 736
rect 2006 737 2012 738
rect 2047 737 2051 738
rect 2215 742 2219 743
rect 2215 737 2219 738
rect 2327 742 2331 743
rect 2327 737 2331 738
rect 2375 742 2379 743
rect 2375 737 2379 738
rect 2447 742 2451 743
rect 2447 737 2451 738
rect 2495 742 2499 743
rect 2495 737 2499 738
rect 2583 742 2587 743
rect 2583 737 2587 738
rect 2623 742 2627 743
rect 2623 737 2627 738
rect 2735 742 2739 743
rect 2735 737 2739 738
rect 2767 742 2771 743
rect 2767 737 2771 738
rect 2895 742 2899 743
rect 2895 737 2899 738
rect 2911 742 2915 743
rect 2911 737 2915 738
rect 3063 742 3067 743
rect 3063 737 3067 738
rect 3215 742 3219 743
rect 3215 737 3219 738
rect 3247 742 3251 743
rect 3247 737 3251 738
rect 3367 742 3371 743
rect 3367 737 3371 738
rect 3447 742 3451 743
rect 3447 737 3451 738
rect 3519 742 3523 743
rect 3519 737 3523 738
rect 3655 742 3659 743
rect 3655 737 3659 738
rect 3679 742 3683 743
rect 3679 737 3683 738
rect 3839 742 3843 743
rect 3839 737 3843 738
rect 3943 742 3947 743
rect 3943 737 3947 738
rect 110 732 116 733
rect 2006 733 2007 737
rect 2011 733 2012 737
rect 2006 732 2012 733
rect 374 721 380 722
rect 110 720 116 721
rect 110 716 111 720
rect 115 716 116 720
rect 374 717 375 721
rect 379 717 380 721
rect 374 716 380 717
rect 494 721 500 722
rect 494 717 495 721
rect 499 717 500 721
rect 494 716 500 717
rect 622 721 628 722
rect 622 717 623 721
rect 627 717 628 721
rect 622 716 628 717
rect 750 721 756 722
rect 750 717 751 721
rect 755 717 756 721
rect 750 716 756 717
rect 886 721 892 722
rect 886 717 887 721
rect 891 717 892 721
rect 886 716 892 717
rect 1022 721 1028 722
rect 1022 717 1023 721
rect 1027 717 1028 721
rect 1022 716 1028 717
rect 1166 721 1172 722
rect 1166 717 1167 721
rect 1171 717 1172 721
rect 1166 716 1172 717
rect 1310 721 1316 722
rect 1310 717 1311 721
rect 1315 717 1316 721
rect 1310 716 1316 717
rect 1454 721 1460 722
rect 1454 717 1455 721
rect 1459 717 1460 721
rect 1454 716 1460 717
rect 1598 721 1604 722
rect 1598 717 1599 721
rect 1603 717 1604 721
rect 1598 716 1604 717
rect 2006 720 2012 721
rect 2006 716 2007 720
rect 2011 716 2012 720
rect 110 715 116 716
rect 112 695 114 715
rect 376 695 378 716
rect 496 695 498 716
rect 624 695 626 716
rect 752 695 754 716
rect 888 695 890 716
rect 1024 695 1026 716
rect 1168 695 1170 716
rect 1312 695 1314 716
rect 1456 695 1458 716
rect 1600 695 1602 716
rect 2006 715 2012 716
rect 2008 695 2010 715
rect 2048 710 2050 737
rect 2376 713 2378 737
rect 2496 713 2498 737
rect 2624 713 2626 737
rect 2768 713 2770 737
rect 2912 713 2914 737
rect 3064 713 3066 737
rect 3216 713 3218 737
rect 3368 713 3370 737
rect 3520 713 3522 737
rect 3680 713 3682 737
rect 3840 713 3842 737
rect 2374 712 2380 713
rect 2046 709 2052 710
rect 2046 705 2047 709
rect 2051 705 2052 709
rect 2374 708 2375 712
rect 2379 708 2380 712
rect 2374 707 2380 708
rect 2494 712 2500 713
rect 2494 708 2495 712
rect 2499 708 2500 712
rect 2494 707 2500 708
rect 2622 712 2628 713
rect 2622 708 2623 712
rect 2627 708 2628 712
rect 2622 707 2628 708
rect 2766 712 2772 713
rect 2766 708 2767 712
rect 2771 708 2772 712
rect 2766 707 2772 708
rect 2910 712 2916 713
rect 2910 708 2911 712
rect 2915 708 2916 712
rect 2910 707 2916 708
rect 3062 712 3068 713
rect 3062 708 3063 712
rect 3067 708 3068 712
rect 3062 707 3068 708
rect 3214 712 3220 713
rect 3214 708 3215 712
rect 3219 708 3220 712
rect 3214 707 3220 708
rect 3366 712 3372 713
rect 3366 708 3367 712
rect 3371 708 3372 712
rect 3366 707 3372 708
rect 3518 712 3524 713
rect 3518 708 3519 712
rect 3523 708 3524 712
rect 3518 707 3524 708
rect 3678 712 3684 713
rect 3678 708 3679 712
rect 3683 708 3684 712
rect 3678 707 3684 708
rect 3838 712 3844 713
rect 3838 708 3839 712
rect 3843 708 3844 712
rect 3944 710 3946 737
rect 3838 707 3844 708
rect 3942 709 3948 710
rect 2046 704 2052 705
rect 3942 705 3943 709
rect 3947 705 3948 709
rect 3942 704 3948 705
rect 111 694 115 695
rect 111 689 115 690
rect 375 694 379 695
rect 375 689 379 690
rect 495 694 499 695
rect 495 689 499 690
rect 527 694 531 695
rect 527 689 531 690
rect 623 694 627 695
rect 623 689 627 690
rect 631 694 635 695
rect 631 689 635 690
rect 743 694 747 695
rect 743 689 747 690
rect 751 694 755 695
rect 751 689 755 690
rect 855 694 859 695
rect 855 689 859 690
rect 887 694 891 695
rect 887 689 891 690
rect 967 694 971 695
rect 967 689 971 690
rect 1023 694 1027 695
rect 1023 689 1027 690
rect 1071 694 1075 695
rect 1071 689 1075 690
rect 1167 694 1171 695
rect 1167 689 1171 690
rect 1183 694 1187 695
rect 1183 689 1187 690
rect 1295 694 1299 695
rect 1295 689 1299 690
rect 1311 694 1315 695
rect 1311 689 1315 690
rect 1407 694 1411 695
rect 1407 689 1411 690
rect 1455 694 1459 695
rect 1455 689 1459 690
rect 1519 694 1523 695
rect 1519 689 1523 690
rect 1599 694 1603 695
rect 1599 689 1603 690
rect 2007 694 2011 695
rect 2374 693 2380 694
rect 2007 689 2011 690
rect 2046 692 2052 693
rect 112 669 114 689
rect 110 668 116 669
rect 528 668 530 689
rect 632 668 634 689
rect 744 668 746 689
rect 856 668 858 689
rect 968 668 970 689
rect 1072 668 1074 689
rect 1184 668 1186 689
rect 1296 668 1298 689
rect 1408 668 1410 689
rect 1520 668 1522 689
rect 2008 669 2010 689
rect 2046 688 2047 692
rect 2051 688 2052 692
rect 2374 689 2375 693
rect 2379 689 2380 693
rect 2374 688 2380 689
rect 2494 693 2500 694
rect 2494 689 2495 693
rect 2499 689 2500 693
rect 2494 688 2500 689
rect 2622 693 2628 694
rect 2622 689 2623 693
rect 2627 689 2628 693
rect 2622 688 2628 689
rect 2766 693 2772 694
rect 2766 689 2767 693
rect 2771 689 2772 693
rect 2766 688 2772 689
rect 2910 693 2916 694
rect 2910 689 2911 693
rect 2915 689 2916 693
rect 2910 688 2916 689
rect 3062 693 3068 694
rect 3062 689 3063 693
rect 3067 689 3068 693
rect 3062 688 3068 689
rect 3214 693 3220 694
rect 3214 689 3215 693
rect 3219 689 3220 693
rect 3214 688 3220 689
rect 3366 693 3372 694
rect 3366 689 3367 693
rect 3371 689 3372 693
rect 3366 688 3372 689
rect 3518 693 3524 694
rect 3518 689 3519 693
rect 3523 689 3524 693
rect 3518 688 3524 689
rect 3678 693 3684 694
rect 3678 689 3679 693
rect 3683 689 3684 693
rect 3678 688 3684 689
rect 3838 693 3844 694
rect 3838 689 3839 693
rect 3843 689 3844 693
rect 3838 688 3844 689
rect 3942 692 3948 693
rect 3942 688 3943 692
rect 3947 688 3948 692
rect 2046 687 2052 688
rect 2006 668 2012 669
rect 110 664 111 668
rect 115 664 116 668
rect 110 663 116 664
rect 526 667 532 668
rect 526 663 527 667
rect 531 663 532 667
rect 526 662 532 663
rect 630 667 636 668
rect 630 663 631 667
rect 635 663 636 667
rect 630 662 636 663
rect 742 667 748 668
rect 742 663 743 667
rect 747 663 748 667
rect 742 662 748 663
rect 854 667 860 668
rect 854 663 855 667
rect 859 663 860 667
rect 854 662 860 663
rect 966 667 972 668
rect 966 663 967 667
rect 971 663 972 667
rect 966 662 972 663
rect 1070 667 1076 668
rect 1070 663 1071 667
rect 1075 663 1076 667
rect 1070 662 1076 663
rect 1182 667 1188 668
rect 1182 663 1183 667
rect 1187 663 1188 667
rect 1182 662 1188 663
rect 1294 667 1300 668
rect 1294 663 1295 667
rect 1299 663 1300 667
rect 1294 662 1300 663
rect 1406 667 1412 668
rect 1406 663 1407 667
rect 1411 663 1412 667
rect 1406 662 1412 663
rect 1518 667 1524 668
rect 1518 663 1519 667
rect 1523 663 1524 667
rect 2006 664 2007 668
rect 2011 664 2012 668
rect 2006 663 2012 664
rect 1518 662 1524 663
rect 2048 659 2050 687
rect 2376 659 2378 688
rect 2496 659 2498 688
rect 2624 659 2626 688
rect 2768 659 2770 688
rect 2912 659 2914 688
rect 3064 659 3066 688
rect 3216 659 3218 688
rect 3368 659 3370 688
rect 3520 659 3522 688
rect 3680 659 3682 688
rect 3840 659 3842 688
rect 3942 687 3948 688
rect 3944 659 3946 687
rect 2047 658 2051 659
rect 2047 653 2051 654
rect 2111 658 2115 659
rect 2111 653 2115 654
rect 2247 658 2251 659
rect 2247 653 2251 654
rect 2375 658 2379 659
rect 2375 653 2379 654
rect 2399 658 2403 659
rect 2399 653 2403 654
rect 2495 658 2499 659
rect 2495 653 2499 654
rect 2575 658 2579 659
rect 2575 653 2579 654
rect 2623 658 2627 659
rect 2623 653 2627 654
rect 2759 658 2763 659
rect 2759 653 2763 654
rect 2767 658 2771 659
rect 2767 653 2771 654
rect 2911 658 2915 659
rect 2911 653 2915 654
rect 2943 658 2947 659
rect 2943 653 2947 654
rect 3063 658 3067 659
rect 3063 653 3067 654
rect 3127 658 3131 659
rect 3127 653 3131 654
rect 3215 658 3219 659
rect 3215 653 3219 654
rect 3303 658 3307 659
rect 3303 653 3307 654
rect 3367 658 3371 659
rect 3367 653 3371 654
rect 3479 658 3483 659
rect 3479 653 3483 654
rect 3519 658 3523 659
rect 3519 653 3523 654
rect 3655 658 3659 659
rect 3655 653 3659 654
rect 3679 658 3683 659
rect 3679 653 3683 654
rect 3831 658 3835 659
rect 3831 653 3835 654
rect 3839 658 3843 659
rect 3839 653 3843 654
rect 3943 658 3947 659
rect 3943 653 3947 654
rect 110 651 116 652
rect 110 647 111 651
rect 115 647 116 651
rect 2006 651 2012 652
rect 110 646 116 647
rect 526 648 532 649
rect 112 619 114 646
rect 526 644 527 648
rect 531 644 532 648
rect 526 643 532 644
rect 630 648 636 649
rect 630 644 631 648
rect 635 644 636 648
rect 630 643 636 644
rect 742 648 748 649
rect 742 644 743 648
rect 747 644 748 648
rect 742 643 748 644
rect 854 648 860 649
rect 854 644 855 648
rect 859 644 860 648
rect 854 643 860 644
rect 966 648 972 649
rect 966 644 967 648
rect 971 644 972 648
rect 966 643 972 644
rect 1070 648 1076 649
rect 1070 644 1071 648
rect 1075 644 1076 648
rect 1070 643 1076 644
rect 1182 648 1188 649
rect 1182 644 1183 648
rect 1187 644 1188 648
rect 1182 643 1188 644
rect 1294 648 1300 649
rect 1294 644 1295 648
rect 1299 644 1300 648
rect 1294 643 1300 644
rect 1406 648 1412 649
rect 1406 644 1407 648
rect 1411 644 1412 648
rect 1406 643 1412 644
rect 1518 648 1524 649
rect 1518 644 1519 648
rect 1523 644 1524 648
rect 2006 647 2007 651
rect 2011 647 2012 651
rect 2006 646 2012 647
rect 1518 643 1524 644
rect 528 619 530 643
rect 632 619 634 643
rect 744 619 746 643
rect 856 619 858 643
rect 968 619 970 643
rect 1072 619 1074 643
rect 1184 619 1186 643
rect 1296 619 1298 643
rect 1408 619 1410 643
rect 1520 619 1522 643
rect 2008 619 2010 646
rect 2048 633 2050 653
rect 2046 632 2052 633
rect 2112 632 2114 653
rect 2248 632 2250 653
rect 2400 632 2402 653
rect 2576 632 2578 653
rect 2760 632 2762 653
rect 2944 632 2946 653
rect 3128 632 3130 653
rect 3304 632 3306 653
rect 3480 632 3482 653
rect 3656 632 3658 653
rect 3832 632 3834 653
rect 3944 633 3946 653
rect 3942 632 3948 633
rect 2046 628 2047 632
rect 2051 628 2052 632
rect 2046 627 2052 628
rect 2110 631 2116 632
rect 2110 627 2111 631
rect 2115 627 2116 631
rect 2110 626 2116 627
rect 2246 631 2252 632
rect 2246 627 2247 631
rect 2251 627 2252 631
rect 2246 626 2252 627
rect 2398 631 2404 632
rect 2398 627 2399 631
rect 2403 627 2404 631
rect 2398 626 2404 627
rect 2574 631 2580 632
rect 2574 627 2575 631
rect 2579 627 2580 631
rect 2574 626 2580 627
rect 2758 631 2764 632
rect 2758 627 2759 631
rect 2763 627 2764 631
rect 2758 626 2764 627
rect 2942 631 2948 632
rect 2942 627 2943 631
rect 2947 627 2948 631
rect 2942 626 2948 627
rect 3126 631 3132 632
rect 3126 627 3127 631
rect 3131 627 3132 631
rect 3126 626 3132 627
rect 3302 631 3308 632
rect 3302 627 3303 631
rect 3307 627 3308 631
rect 3302 626 3308 627
rect 3478 631 3484 632
rect 3478 627 3479 631
rect 3483 627 3484 631
rect 3478 626 3484 627
rect 3654 631 3660 632
rect 3654 627 3655 631
rect 3659 627 3660 631
rect 3654 626 3660 627
rect 3830 631 3836 632
rect 3830 627 3831 631
rect 3835 627 3836 631
rect 3942 628 3943 632
rect 3947 628 3948 632
rect 3942 627 3948 628
rect 3830 626 3836 627
rect 111 618 115 619
rect 111 613 115 614
rect 527 618 531 619
rect 527 613 531 614
rect 631 618 635 619
rect 631 613 635 614
rect 687 618 691 619
rect 687 613 691 614
rect 743 618 747 619
rect 743 613 747 614
rect 783 618 787 619
rect 783 613 787 614
rect 855 618 859 619
rect 855 613 859 614
rect 879 618 883 619
rect 879 613 883 614
rect 967 618 971 619
rect 967 613 971 614
rect 975 618 979 619
rect 975 613 979 614
rect 1071 618 1075 619
rect 1071 613 1075 614
rect 1167 618 1171 619
rect 1167 613 1171 614
rect 1183 618 1187 619
rect 1183 613 1187 614
rect 1263 618 1267 619
rect 1263 613 1267 614
rect 1295 618 1299 619
rect 1295 613 1299 614
rect 1359 618 1363 619
rect 1359 613 1363 614
rect 1407 618 1411 619
rect 1407 613 1411 614
rect 1455 618 1459 619
rect 1455 613 1459 614
rect 1519 618 1523 619
rect 1519 613 1523 614
rect 2007 618 2011 619
rect 2007 613 2011 614
rect 2046 615 2052 616
rect 112 586 114 613
rect 688 589 690 613
rect 784 589 786 613
rect 880 589 882 613
rect 976 589 978 613
rect 1072 589 1074 613
rect 1168 589 1170 613
rect 1264 589 1266 613
rect 1360 589 1362 613
rect 1456 589 1458 613
rect 686 588 692 589
rect 110 585 116 586
rect 110 581 111 585
rect 115 581 116 585
rect 686 584 687 588
rect 691 584 692 588
rect 686 583 692 584
rect 782 588 788 589
rect 782 584 783 588
rect 787 584 788 588
rect 782 583 788 584
rect 878 588 884 589
rect 878 584 879 588
rect 883 584 884 588
rect 878 583 884 584
rect 974 588 980 589
rect 974 584 975 588
rect 979 584 980 588
rect 974 583 980 584
rect 1070 588 1076 589
rect 1070 584 1071 588
rect 1075 584 1076 588
rect 1070 583 1076 584
rect 1166 588 1172 589
rect 1166 584 1167 588
rect 1171 584 1172 588
rect 1166 583 1172 584
rect 1262 588 1268 589
rect 1262 584 1263 588
rect 1267 584 1268 588
rect 1262 583 1268 584
rect 1358 588 1364 589
rect 1358 584 1359 588
rect 1363 584 1364 588
rect 1358 583 1364 584
rect 1454 588 1460 589
rect 1454 584 1455 588
rect 1459 584 1460 588
rect 2008 586 2010 613
rect 2046 611 2047 615
rect 2051 611 2052 615
rect 3942 615 3948 616
rect 2046 610 2052 611
rect 2110 612 2116 613
rect 1454 583 1460 584
rect 2006 585 2012 586
rect 110 580 116 581
rect 2006 581 2007 585
rect 2011 581 2012 585
rect 2006 580 2012 581
rect 2048 579 2050 610
rect 2110 608 2111 612
rect 2115 608 2116 612
rect 2110 607 2116 608
rect 2246 612 2252 613
rect 2246 608 2247 612
rect 2251 608 2252 612
rect 2246 607 2252 608
rect 2398 612 2404 613
rect 2398 608 2399 612
rect 2403 608 2404 612
rect 2398 607 2404 608
rect 2574 612 2580 613
rect 2574 608 2575 612
rect 2579 608 2580 612
rect 2574 607 2580 608
rect 2758 612 2764 613
rect 2758 608 2759 612
rect 2763 608 2764 612
rect 2758 607 2764 608
rect 2942 612 2948 613
rect 2942 608 2943 612
rect 2947 608 2948 612
rect 2942 607 2948 608
rect 3126 612 3132 613
rect 3126 608 3127 612
rect 3131 608 3132 612
rect 3126 607 3132 608
rect 3302 612 3308 613
rect 3302 608 3303 612
rect 3307 608 3308 612
rect 3302 607 3308 608
rect 3478 612 3484 613
rect 3478 608 3479 612
rect 3483 608 3484 612
rect 3478 607 3484 608
rect 3654 612 3660 613
rect 3654 608 3655 612
rect 3659 608 3660 612
rect 3654 607 3660 608
rect 3830 612 3836 613
rect 3830 608 3831 612
rect 3835 608 3836 612
rect 3942 611 3943 615
rect 3947 611 3948 615
rect 3942 610 3948 611
rect 3830 607 3836 608
rect 2112 579 2114 607
rect 2248 579 2250 607
rect 2400 579 2402 607
rect 2576 579 2578 607
rect 2760 579 2762 607
rect 2944 579 2946 607
rect 3128 579 3130 607
rect 3304 579 3306 607
rect 3480 579 3482 607
rect 3656 579 3658 607
rect 3832 579 3834 607
rect 3944 579 3946 610
rect 2047 578 2051 579
rect 2047 573 2051 574
rect 2071 578 2075 579
rect 2071 573 2075 574
rect 2111 578 2115 579
rect 2111 573 2115 574
rect 2183 578 2187 579
rect 2183 573 2187 574
rect 2247 578 2251 579
rect 2247 573 2251 574
rect 2335 578 2339 579
rect 2335 573 2339 574
rect 2399 578 2403 579
rect 2399 573 2403 574
rect 2503 578 2507 579
rect 2503 573 2507 574
rect 2575 578 2579 579
rect 2575 573 2579 574
rect 2687 578 2691 579
rect 2687 573 2691 574
rect 2759 578 2763 579
rect 2759 573 2763 574
rect 2879 578 2883 579
rect 2879 573 2883 574
rect 2943 578 2947 579
rect 2943 573 2947 574
rect 3071 578 3075 579
rect 3071 573 3075 574
rect 3127 578 3131 579
rect 3127 573 3131 574
rect 3263 578 3267 579
rect 3263 573 3267 574
rect 3303 578 3307 579
rect 3303 573 3307 574
rect 3455 578 3459 579
rect 3455 573 3459 574
rect 3479 578 3483 579
rect 3479 573 3483 574
rect 3647 578 3651 579
rect 3647 573 3651 574
rect 3655 578 3659 579
rect 3655 573 3659 574
rect 3831 578 3835 579
rect 3831 573 3835 574
rect 3839 578 3843 579
rect 3839 573 3843 574
rect 3943 578 3947 579
rect 3943 573 3947 574
rect 686 569 692 570
rect 110 568 116 569
rect 110 564 111 568
rect 115 564 116 568
rect 686 565 687 569
rect 691 565 692 569
rect 686 564 692 565
rect 782 569 788 570
rect 782 565 783 569
rect 787 565 788 569
rect 782 564 788 565
rect 878 569 884 570
rect 878 565 879 569
rect 883 565 884 569
rect 878 564 884 565
rect 974 569 980 570
rect 974 565 975 569
rect 979 565 980 569
rect 974 564 980 565
rect 1070 569 1076 570
rect 1070 565 1071 569
rect 1075 565 1076 569
rect 1070 564 1076 565
rect 1166 569 1172 570
rect 1166 565 1167 569
rect 1171 565 1172 569
rect 1166 564 1172 565
rect 1262 569 1268 570
rect 1262 565 1263 569
rect 1267 565 1268 569
rect 1262 564 1268 565
rect 1358 569 1364 570
rect 1358 565 1359 569
rect 1363 565 1364 569
rect 1358 564 1364 565
rect 1454 569 1460 570
rect 1454 565 1455 569
rect 1459 565 1460 569
rect 1454 564 1460 565
rect 2006 568 2012 569
rect 2006 564 2007 568
rect 2011 564 2012 568
rect 110 563 116 564
rect 112 523 114 563
rect 688 523 690 564
rect 784 523 786 564
rect 880 523 882 564
rect 976 523 978 564
rect 1072 523 1074 564
rect 1168 523 1170 564
rect 1264 523 1266 564
rect 1360 523 1362 564
rect 1456 523 1458 564
rect 2006 563 2012 564
rect 2008 523 2010 563
rect 2048 546 2050 573
rect 2072 549 2074 573
rect 2184 549 2186 573
rect 2336 549 2338 573
rect 2504 549 2506 573
rect 2688 549 2690 573
rect 2880 549 2882 573
rect 3072 549 3074 573
rect 3264 549 3266 573
rect 3456 549 3458 573
rect 3648 549 3650 573
rect 3840 549 3842 573
rect 2070 548 2076 549
rect 2046 545 2052 546
rect 2046 541 2047 545
rect 2051 541 2052 545
rect 2070 544 2071 548
rect 2075 544 2076 548
rect 2070 543 2076 544
rect 2182 548 2188 549
rect 2182 544 2183 548
rect 2187 544 2188 548
rect 2182 543 2188 544
rect 2334 548 2340 549
rect 2334 544 2335 548
rect 2339 544 2340 548
rect 2334 543 2340 544
rect 2502 548 2508 549
rect 2502 544 2503 548
rect 2507 544 2508 548
rect 2502 543 2508 544
rect 2686 548 2692 549
rect 2686 544 2687 548
rect 2691 544 2692 548
rect 2686 543 2692 544
rect 2878 548 2884 549
rect 2878 544 2879 548
rect 2883 544 2884 548
rect 2878 543 2884 544
rect 3070 548 3076 549
rect 3070 544 3071 548
rect 3075 544 3076 548
rect 3070 543 3076 544
rect 3262 548 3268 549
rect 3262 544 3263 548
rect 3267 544 3268 548
rect 3262 543 3268 544
rect 3454 548 3460 549
rect 3454 544 3455 548
rect 3459 544 3460 548
rect 3454 543 3460 544
rect 3646 548 3652 549
rect 3646 544 3647 548
rect 3651 544 3652 548
rect 3646 543 3652 544
rect 3838 548 3844 549
rect 3838 544 3839 548
rect 3843 544 3844 548
rect 3944 546 3946 573
rect 3838 543 3844 544
rect 3942 545 3948 546
rect 2046 540 2052 541
rect 3942 541 3943 545
rect 3947 541 3948 545
rect 3942 540 3948 541
rect 2070 529 2076 530
rect 2046 528 2052 529
rect 2046 524 2047 528
rect 2051 524 2052 528
rect 2070 525 2071 529
rect 2075 525 2076 529
rect 2070 524 2076 525
rect 2182 529 2188 530
rect 2182 525 2183 529
rect 2187 525 2188 529
rect 2182 524 2188 525
rect 2334 529 2340 530
rect 2334 525 2335 529
rect 2339 525 2340 529
rect 2334 524 2340 525
rect 2502 529 2508 530
rect 2502 525 2503 529
rect 2507 525 2508 529
rect 2502 524 2508 525
rect 2686 529 2692 530
rect 2686 525 2687 529
rect 2691 525 2692 529
rect 2686 524 2692 525
rect 2878 529 2884 530
rect 2878 525 2879 529
rect 2883 525 2884 529
rect 2878 524 2884 525
rect 3070 529 3076 530
rect 3070 525 3071 529
rect 3075 525 3076 529
rect 3070 524 3076 525
rect 3262 529 3268 530
rect 3262 525 3263 529
rect 3267 525 3268 529
rect 3262 524 3268 525
rect 3454 529 3460 530
rect 3454 525 3455 529
rect 3459 525 3460 529
rect 3454 524 3460 525
rect 3646 529 3652 530
rect 3646 525 3647 529
rect 3651 525 3652 529
rect 3646 524 3652 525
rect 3838 529 3844 530
rect 3838 525 3839 529
rect 3843 525 3844 529
rect 3838 524 3844 525
rect 3942 528 3948 529
rect 3942 524 3943 528
rect 3947 524 3948 528
rect 2046 523 2052 524
rect 111 522 115 523
rect 111 517 115 518
rect 383 522 387 523
rect 383 517 387 518
rect 479 522 483 523
rect 479 517 483 518
rect 575 522 579 523
rect 575 517 579 518
rect 671 522 675 523
rect 671 517 675 518
rect 687 522 691 523
rect 687 517 691 518
rect 767 522 771 523
rect 767 517 771 518
rect 783 522 787 523
rect 783 517 787 518
rect 863 522 867 523
rect 863 517 867 518
rect 879 522 883 523
rect 879 517 883 518
rect 959 522 963 523
rect 959 517 963 518
rect 975 522 979 523
rect 975 517 979 518
rect 1055 522 1059 523
rect 1055 517 1059 518
rect 1071 522 1075 523
rect 1071 517 1075 518
rect 1151 522 1155 523
rect 1151 517 1155 518
rect 1167 522 1171 523
rect 1167 517 1171 518
rect 1247 522 1251 523
rect 1247 517 1251 518
rect 1263 522 1267 523
rect 1263 517 1267 518
rect 1343 522 1347 523
rect 1343 517 1347 518
rect 1359 522 1363 523
rect 1359 517 1363 518
rect 1439 522 1443 523
rect 1439 517 1443 518
rect 1455 522 1459 523
rect 1455 517 1459 518
rect 1535 522 1539 523
rect 1535 517 1539 518
rect 2007 522 2011 523
rect 2007 517 2011 518
rect 112 497 114 517
rect 110 496 116 497
rect 384 496 386 517
rect 480 496 482 517
rect 576 496 578 517
rect 672 496 674 517
rect 768 496 770 517
rect 864 496 866 517
rect 960 496 962 517
rect 1056 496 1058 517
rect 1152 496 1154 517
rect 1248 496 1250 517
rect 1344 496 1346 517
rect 1440 496 1442 517
rect 1536 496 1538 517
rect 2008 497 2010 517
rect 2048 503 2050 523
rect 2072 503 2074 524
rect 2184 503 2186 524
rect 2336 503 2338 524
rect 2504 503 2506 524
rect 2688 503 2690 524
rect 2880 503 2882 524
rect 3072 503 3074 524
rect 3264 503 3266 524
rect 3456 503 3458 524
rect 3648 503 3650 524
rect 3840 503 3842 524
rect 3942 523 3948 524
rect 3944 503 3946 523
rect 2047 502 2051 503
rect 2047 497 2051 498
rect 2071 502 2075 503
rect 2071 497 2075 498
rect 2183 502 2187 503
rect 2183 497 2187 498
rect 2319 502 2323 503
rect 2319 497 2323 498
rect 2335 502 2339 503
rect 2335 497 2339 498
rect 2463 502 2467 503
rect 2463 497 2467 498
rect 2503 502 2507 503
rect 2503 497 2507 498
rect 2615 502 2619 503
rect 2615 497 2619 498
rect 2687 502 2691 503
rect 2687 497 2691 498
rect 2775 502 2779 503
rect 2775 497 2779 498
rect 2879 502 2883 503
rect 2879 497 2883 498
rect 2959 502 2963 503
rect 2959 497 2963 498
rect 3071 502 3075 503
rect 3071 497 3075 498
rect 3159 502 3163 503
rect 3159 497 3163 498
rect 3263 502 3267 503
rect 3263 497 3267 498
rect 3367 502 3371 503
rect 3367 497 3371 498
rect 3455 502 3459 503
rect 3455 497 3459 498
rect 3583 502 3587 503
rect 3583 497 3587 498
rect 3647 502 3651 503
rect 3647 497 3651 498
rect 3807 502 3811 503
rect 3807 497 3811 498
rect 3839 502 3843 503
rect 3839 497 3843 498
rect 3943 502 3947 503
rect 3943 497 3947 498
rect 2006 496 2012 497
rect 110 492 111 496
rect 115 492 116 496
rect 110 491 116 492
rect 382 495 388 496
rect 382 491 383 495
rect 387 491 388 495
rect 382 490 388 491
rect 478 495 484 496
rect 478 491 479 495
rect 483 491 484 495
rect 478 490 484 491
rect 574 495 580 496
rect 574 491 575 495
rect 579 491 580 495
rect 574 490 580 491
rect 670 495 676 496
rect 670 491 671 495
rect 675 491 676 495
rect 670 490 676 491
rect 766 495 772 496
rect 766 491 767 495
rect 771 491 772 495
rect 766 490 772 491
rect 862 495 868 496
rect 862 491 863 495
rect 867 491 868 495
rect 862 490 868 491
rect 958 495 964 496
rect 958 491 959 495
rect 963 491 964 495
rect 958 490 964 491
rect 1054 495 1060 496
rect 1054 491 1055 495
rect 1059 491 1060 495
rect 1054 490 1060 491
rect 1150 495 1156 496
rect 1150 491 1151 495
rect 1155 491 1156 495
rect 1150 490 1156 491
rect 1246 495 1252 496
rect 1246 491 1247 495
rect 1251 491 1252 495
rect 1246 490 1252 491
rect 1342 495 1348 496
rect 1342 491 1343 495
rect 1347 491 1348 495
rect 1342 490 1348 491
rect 1438 495 1444 496
rect 1438 491 1439 495
rect 1443 491 1444 495
rect 1438 490 1444 491
rect 1534 495 1540 496
rect 1534 491 1535 495
rect 1539 491 1540 495
rect 2006 492 2007 496
rect 2011 492 2012 496
rect 2006 491 2012 492
rect 1534 490 1540 491
rect 110 479 116 480
rect 110 475 111 479
rect 115 475 116 479
rect 2006 479 2012 480
rect 110 474 116 475
rect 382 476 388 477
rect 112 435 114 474
rect 382 472 383 476
rect 387 472 388 476
rect 382 471 388 472
rect 478 476 484 477
rect 478 472 479 476
rect 483 472 484 476
rect 478 471 484 472
rect 574 476 580 477
rect 574 472 575 476
rect 579 472 580 476
rect 574 471 580 472
rect 670 476 676 477
rect 670 472 671 476
rect 675 472 676 476
rect 670 471 676 472
rect 766 476 772 477
rect 766 472 767 476
rect 771 472 772 476
rect 766 471 772 472
rect 862 476 868 477
rect 862 472 863 476
rect 867 472 868 476
rect 862 471 868 472
rect 958 476 964 477
rect 958 472 959 476
rect 963 472 964 476
rect 958 471 964 472
rect 1054 476 1060 477
rect 1054 472 1055 476
rect 1059 472 1060 476
rect 1054 471 1060 472
rect 1150 476 1156 477
rect 1150 472 1151 476
rect 1155 472 1156 476
rect 1150 471 1156 472
rect 1246 476 1252 477
rect 1246 472 1247 476
rect 1251 472 1252 476
rect 1246 471 1252 472
rect 1342 476 1348 477
rect 1342 472 1343 476
rect 1347 472 1348 476
rect 1342 471 1348 472
rect 1438 476 1444 477
rect 1438 472 1439 476
rect 1443 472 1444 476
rect 1438 471 1444 472
rect 1534 476 1540 477
rect 1534 472 1535 476
rect 1539 472 1540 476
rect 2006 475 2007 479
rect 2011 475 2012 479
rect 2048 477 2050 497
rect 2006 474 2012 475
rect 2046 476 2052 477
rect 2184 476 2186 497
rect 2320 476 2322 497
rect 2464 476 2466 497
rect 2616 476 2618 497
rect 2776 476 2778 497
rect 2960 476 2962 497
rect 3160 476 3162 497
rect 3368 476 3370 497
rect 3584 476 3586 497
rect 3808 476 3810 497
rect 3944 477 3946 497
rect 3942 476 3948 477
rect 1534 471 1540 472
rect 384 435 386 471
rect 480 435 482 471
rect 576 435 578 471
rect 672 435 674 471
rect 768 435 770 471
rect 864 435 866 471
rect 960 435 962 471
rect 1056 435 1058 471
rect 1152 435 1154 471
rect 1248 435 1250 471
rect 1344 435 1346 471
rect 1440 435 1442 471
rect 1536 435 1538 471
rect 2008 435 2010 474
rect 2046 472 2047 476
rect 2051 472 2052 476
rect 2046 471 2052 472
rect 2182 475 2188 476
rect 2182 471 2183 475
rect 2187 471 2188 475
rect 2182 470 2188 471
rect 2318 475 2324 476
rect 2318 471 2319 475
rect 2323 471 2324 475
rect 2318 470 2324 471
rect 2462 475 2468 476
rect 2462 471 2463 475
rect 2467 471 2468 475
rect 2462 470 2468 471
rect 2614 475 2620 476
rect 2614 471 2615 475
rect 2619 471 2620 475
rect 2614 470 2620 471
rect 2774 475 2780 476
rect 2774 471 2775 475
rect 2779 471 2780 475
rect 2774 470 2780 471
rect 2958 475 2964 476
rect 2958 471 2959 475
rect 2963 471 2964 475
rect 2958 470 2964 471
rect 3158 475 3164 476
rect 3158 471 3159 475
rect 3163 471 3164 475
rect 3158 470 3164 471
rect 3366 475 3372 476
rect 3366 471 3367 475
rect 3371 471 3372 475
rect 3366 470 3372 471
rect 3582 475 3588 476
rect 3582 471 3583 475
rect 3587 471 3588 475
rect 3582 470 3588 471
rect 3806 475 3812 476
rect 3806 471 3807 475
rect 3811 471 3812 475
rect 3942 472 3943 476
rect 3947 472 3948 476
rect 3942 471 3948 472
rect 3806 470 3812 471
rect 2046 459 2052 460
rect 2046 455 2047 459
rect 2051 455 2052 459
rect 3942 459 3948 460
rect 2046 454 2052 455
rect 2182 456 2188 457
rect 111 434 115 435
rect 111 429 115 430
rect 383 434 387 435
rect 383 429 387 430
rect 479 434 483 435
rect 479 429 483 430
rect 487 434 491 435
rect 487 429 491 430
rect 575 434 579 435
rect 575 429 579 430
rect 583 434 587 435
rect 583 429 587 430
rect 671 434 675 435
rect 671 429 675 430
rect 687 434 691 435
rect 687 429 691 430
rect 767 434 771 435
rect 767 429 771 430
rect 791 434 795 435
rect 791 429 795 430
rect 863 434 867 435
rect 863 429 867 430
rect 895 434 899 435
rect 895 429 899 430
rect 959 434 963 435
rect 959 429 963 430
rect 999 434 1003 435
rect 999 429 1003 430
rect 1055 434 1059 435
rect 1055 429 1059 430
rect 1103 434 1107 435
rect 1103 429 1107 430
rect 1151 434 1155 435
rect 1151 429 1155 430
rect 1207 434 1211 435
rect 1207 429 1211 430
rect 1247 434 1251 435
rect 1247 429 1251 430
rect 1319 434 1323 435
rect 1319 429 1323 430
rect 1343 434 1347 435
rect 1343 429 1347 430
rect 1431 434 1435 435
rect 1431 429 1435 430
rect 1439 434 1443 435
rect 1439 429 1443 430
rect 1535 434 1539 435
rect 1535 429 1539 430
rect 2007 434 2011 435
rect 2007 429 2011 430
rect 112 402 114 429
rect 488 405 490 429
rect 584 405 586 429
rect 688 405 690 429
rect 792 405 794 429
rect 896 405 898 429
rect 1000 405 1002 429
rect 1104 405 1106 429
rect 1208 405 1210 429
rect 1320 405 1322 429
rect 1432 405 1434 429
rect 486 404 492 405
rect 110 401 116 402
rect 110 397 111 401
rect 115 397 116 401
rect 486 400 487 404
rect 491 400 492 404
rect 486 399 492 400
rect 582 404 588 405
rect 582 400 583 404
rect 587 400 588 404
rect 582 399 588 400
rect 686 404 692 405
rect 686 400 687 404
rect 691 400 692 404
rect 686 399 692 400
rect 790 404 796 405
rect 790 400 791 404
rect 795 400 796 404
rect 790 399 796 400
rect 894 404 900 405
rect 894 400 895 404
rect 899 400 900 404
rect 894 399 900 400
rect 998 404 1004 405
rect 998 400 999 404
rect 1003 400 1004 404
rect 998 399 1004 400
rect 1102 404 1108 405
rect 1102 400 1103 404
rect 1107 400 1108 404
rect 1102 399 1108 400
rect 1206 404 1212 405
rect 1206 400 1207 404
rect 1211 400 1212 404
rect 1206 399 1212 400
rect 1318 404 1324 405
rect 1318 400 1319 404
rect 1323 400 1324 404
rect 1318 399 1324 400
rect 1430 404 1436 405
rect 1430 400 1431 404
rect 1435 400 1436 404
rect 2008 402 2010 429
rect 2048 427 2050 454
rect 2182 452 2183 456
rect 2187 452 2188 456
rect 2182 451 2188 452
rect 2318 456 2324 457
rect 2318 452 2319 456
rect 2323 452 2324 456
rect 2318 451 2324 452
rect 2462 456 2468 457
rect 2462 452 2463 456
rect 2467 452 2468 456
rect 2462 451 2468 452
rect 2614 456 2620 457
rect 2614 452 2615 456
rect 2619 452 2620 456
rect 2614 451 2620 452
rect 2774 456 2780 457
rect 2774 452 2775 456
rect 2779 452 2780 456
rect 2774 451 2780 452
rect 2958 456 2964 457
rect 2958 452 2959 456
rect 2963 452 2964 456
rect 2958 451 2964 452
rect 3158 456 3164 457
rect 3158 452 3159 456
rect 3163 452 3164 456
rect 3158 451 3164 452
rect 3366 456 3372 457
rect 3366 452 3367 456
rect 3371 452 3372 456
rect 3366 451 3372 452
rect 3582 456 3588 457
rect 3582 452 3583 456
rect 3587 452 3588 456
rect 3582 451 3588 452
rect 3806 456 3812 457
rect 3806 452 3807 456
rect 3811 452 3812 456
rect 3942 455 3943 459
rect 3947 455 3948 459
rect 3942 454 3948 455
rect 3806 451 3812 452
rect 2184 427 2186 451
rect 2320 427 2322 451
rect 2464 427 2466 451
rect 2616 427 2618 451
rect 2776 427 2778 451
rect 2960 427 2962 451
rect 3160 427 3162 451
rect 3368 427 3370 451
rect 3584 427 3586 451
rect 3808 427 3810 451
rect 3944 427 3946 454
rect 2047 426 2051 427
rect 2047 421 2051 422
rect 2183 426 2187 427
rect 2183 421 2187 422
rect 2319 426 2323 427
rect 2319 421 2323 422
rect 2343 426 2347 427
rect 2343 421 2347 422
rect 2463 426 2467 427
rect 2463 421 2467 422
rect 2487 426 2491 427
rect 2487 421 2491 422
rect 2615 426 2619 427
rect 2615 421 2619 422
rect 2639 426 2643 427
rect 2639 421 2643 422
rect 2775 426 2779 427
rect 2775 421 2779 422
rect 2799 426 2803 427
rect 2799 421 2803 422
rect 2959 426 2963 427
rect 2959 421 2963 422
rect 3111 426 3115 427
rect 3111 421 3115 422
rect 3159 426 3163 427
rect 3159 421 3163 422
rect 3263 426 3267 427
rect 3263 421 3267 422
rect 3367 426 3371 427
rect 3367 421 3371 422
rect 3415 426 3419 427
rect 3415 421 3419 422
rect 3559 426 3563 427
rect 3559 421 3563 422
rect 3583 426 3587 427
rect 3583 421 3587 422
rect 3711 426 3715 427
rect 3711 421 3715 422
rect 3807 426 3811 427
rect 3807 421 3811 422
rect 3839 426 3843 427
rect 3839 421 3843 422
rect 3943 426 3947 427
rect 3943 421 3947 422
rect 1430 399 1436 400
rect 2006 401 2012 402
rect 110 396 116 397
rect 2006 397 2007 401
rect 2011 397 2012 401
rect 2006 396 2012 397
rect 2048 394 2050 421
rect 2344 397 2346 421
rect 2488 397 2490 421
rect 2640 397 2642 421
rect 2800 397 2802 421
rect 2960 397 2962 421
rect 3112 397 3114 421
rect 3264 397 3266 421
rect 3416 397 3418 421
rect 3560 397 3562 421
rect 3712 397 3714 421
rect 3840 397 3842 421
rect 2342 396 2348 397
rect 2046 393 2052 394
rect 2046 389 2047 393
rect 2051 389 2052 393
rect 2342 392 2343 396
rect 2347 392 2348 396
rect 2342 391 2348 392
rect 2486 396 2492 397
rect 2486 392 2487 396
rect 2491 392 2492 396
rect 2486 391 2492 392
rect 2638 396 2644 397
rect 2638 392 2639 396
rect 2643 392 2644 396
rect 2638 391 2644 392
rect 2798 396 2804 397
rect 2798 392 2799 396
rect 2803 392 2804 396
rect 2798 391 2804 392
rect 2958 396 2964 397
rect 2958 392 2959 396
rect 2963 392 2964 396
rect 2958 391 2964 392
rect 3110 396 3116 397
rect 3110 392 3111 396
rect 3115 392 3116 396
rect 3110 391 3116 392
rect 3262 396 3268 397
rect 3262 392 3263 396
rect 3267 392 3268 396
rect 3262 391 3268 392
rect 3414 396 3420 397
rect 3414 392 3415 396
rect 3419 392 3420 396
rect 3414 391 3420 392
rect 3558 396 3564 397
rect 3558 392 3559 396
rect 3563 392 3564 396
rect 3558 391 3564 392
rect 3710 396 3716 397
rect 3710 392 3711 396
rect 3715 392 3716 396
rect 3710 391 3716 392
rect 3838 396 3844 397
rect 3838 392 3839 396
rect 3843 392 3844 396
rect 3944 394 3946 421
rect 3838 391 3844 392
rect 3942 393 3948 394
rect 2046 388 2052 389
rect 3942 389 3943 393
rect 3947 389 3948 393
rect 3942 388 3948 389
rect 486 385 492 386
rect 110 384 116 385
rect 110 380 111 384
rect 115 380 116 384
rect 486 381 487 385
rect 491 381 492 385
rect 486 380 492 381
rect 582 385 588 386
rect 582 381 583 385
rect 587 381 588 385
rect 582 380 588 381
rect 686 385 692 386
rect 686 381 687 385
rect 691 381 692 385
rect 686 380 692 381
rect 790 385 796 386
rect 790 381 791 385
rect 795 381 796 385
rect 790 380 796 381
rect 894 385 900 386
rect 894 381 895 385
rect 899 381 900 385
rect 894 380 900 381
rect 998 385 1004 386
rect 998 381 999 385
rect 1003 381 1004 385
rect 998 380 1004 381
rect 1102 385 1108 386
rect 1102 381 1103 385
rect 1107 381 1108 385
rect 1102 380 1108 381
rect 1206 385 1212 386
rect 1206 381 1207 385
rect 1211 381 1212 385
rect 1206 380 1212 381
rect 1318 385 1324 386
rect 1318 381 1319 385
rect 1323 381 1324 385
rect 1318 380 1324 381
rect 1430 385 1436 386
rect 1430 381 1431 385
rect 1435 381 1436 385
rect 1430 380 1436 381
rect 2006 384 2012 385
rect 2006 380 2007 384
rect 2011 380 2012 384
rect 110 379 116 380
rect 112 355 114 379
rect 488 355 490 380
rect 584 355 586 380
rect 688 355 690 380
rect 792 355 794 380
rect 896 355 898 380
rect 1000 355 1002 380
rect 1104 355 1106 380
rect 1208 355 1210 380
rect 1320 355 1322 380
rect 1432 355 1434 380
rect 2006 379 2012 380
rect 2008 355 2010 379
rect 2342 377 2348 378
rect 2046 376 2052 377
rect 2046 372 2047 376
rect 2051 372 2052 376
rect 2342 373 2343 377
rect 2347 373 2348 377
rect 2342 372 2348 373
rect 2486 377 2492 378
rect 2486 373 2487 377
rect 2491 373 2492 377
rect 2486 372 2492 373
rect 2638 377 2644 378
rect 2638 373 2639 377
rect 2643 373 2644 377
rect 2638 372 2644 373
rect 2798 377 2804 378
rect 2798 373 2799 377
rect 2803 373 2804 377
rect 2798 372 2804 373
rect 2958 377 2964 378
rect 2958 373 2959 377
rect 2963 373 2964 377
rect 2958 372 2964 373
rect 3110 377 3116 378
rect 3110 373 3111 377
rect 3115 373 3116 377
rect 3110 372 3116 373
rect 3262 377 3268 378
rect 3262 373 3263 377
rect 3267 373 3268 377
rect 3262 372 3268 373
rect 3414 377 3420 378
rect 3414 373 3415 377
rect 3419 373 3420 377
rect 3414 372 3420 373
rect 3558 377 3564 378
rect 3558 373 3559 377
rect 3563 373 3564 377
rect 3558 372 3564 373
rect 3710 377 3716 378
rect 3710 373 3711 377
rect 3715 373 3716 377
rect 3710 372 3716 373
rect 3838 377 3844 378
rect 3838 373 3839 377
rect 3843 373 3844 377
rect 3838 372 3844 373
rect 3942 376 3948 377
rect 3942 372 3943 376
rect 3947 372 3948 376
rect 2046 371 2052 372
rect 111 354 115 355
rect 111 349 115 350
rect 327 354 331 355
rect 327 349 331 350
rect 463 354 467 355
rect 463 349 467 350
rect 487 354 491 355
rect 487 349 491 350
rect 583 354 587 355
rect 583 349 587 350
rect 615 354 619 355
rect 615 349 619 350
rect 687 354 691 355
rect 687 349 691 350
rect 767 354 771 355
rect 767 349 771 350
rect 791 354 795 355
rect 791 349 795 350
rect 895 354 899 355
rect 895 349 899 350
rect 919 354 923 355
rect 919 349 923 350
rect 999 354 1003 355
rect 999 349 1003 350
rect 1063 354 1067 355
rect 1063 349 1067 350
rect 1103 354 1107 355
rect 1103 349 1107 350
rect 1207 354 1211 355
rect 1207 349 1211 350
rect 1319 354 1323 355
rect 1319 349 1323 350
rect 1351 354 1355 355
rect 1351 349 1355 350
rect 1431 354 1435 355
rect 1431 349 1435 350
rect 1495 354 1499 355
rect 1495 349 1499 350
rect 1639 354 1643 355
rect 1639 349 1643 350
rect 2007 354 2011 355
rect 2007 349 2011 350
rect 112 329 114 349
rect 110 328 116 329
rect 328 328 330 349
rect 464 328 466 349
rect 616 328 618 349
rect 768 328 770 349
rect 920 328 922 349
rect 1064 328 1066 349
rect 1208 328 1210 349
rect 1352 328 1354 349
rect 1496 328 1498 349
rect 1640 328 1642 349
rect 2008 329 2010 349
rect 2048 347 2050 371
rect 2344 347 2346 372
rect 2488 347 2490 372
rect 2640 347 2642 372
rect 2800 347 2802 372
rect 2960 347 2962 372
rect 3112 347 3114 372
rect 3264 347 3266 372
rect 3416 347 3418 372
rect 3560 347 3562 372
rect 3712 347 3714 372
rect 3840 347 3842 372
rect 3942 371 3948 372
rect 3944 347 3946 371
rect 2047 346 2051 347
rect 2047 341 2051 342
rect 2343 346 2347 347
rect 2343 341 2347 342
rect 2487 346 2491 347
rect 2487 341 2491 342
rect 2495 346 2499 347
rect 2495 341 2499 342
rect 2639 346 2643 347
rect 2639 341 2643 342
rect 2799 346 2803 347
rect 2799 341 2803 342
rect 2959 346 2963 347
rect 2959 341 2963 342
rect 3111 346 3115 347
rect 3111 341 3115 342
rect 3119 346 3123 347
rect 3119 341 3123 342
rect 3263 346 3267 347
rect 3263 341 3267 342
rect 3271 346 3275 347
rect 3271 341 3275 342
rect 3415 346 3419 347
rect 3415 341 3419 342
rect 3423 346 3427 347
rect 3423 341 3427 342
rect 3559 346 3563 347
rect 3559 341 3563 342
rect 3567 346 3571 347
rect 3567 341 3571 342
rect 3711 346 3715 347
rect 3711 341 3715 342
rect 3839 346 3843 347
rect 3839 341 3843 342
rect 3943 346 3947 347
rect 3943 341 3947 342
rect 2006 328 2012 329
rect 110 324 111 328
rect 115 324 116 328
rect 110 323 116 324
rect 326 327 332 328
rect 326 323 327 327
rect 331 323 332 327
rect 326 322 332 323
rect 462 327 468 328
rect 462 323 463 327
rect 467 323 468 327
rect 462 322 468 323
rect 614 327 620 328
rect 614 323 615 327
rect 619 323 620 327
rect 614 322 620 323
rect 766 327 772 328
rect 766 323 767 327
rect 771 323 772 327
rect 766 322 772 323
rect 918 327 924 328
rect 918 323 919 327
rect 923 323 924 327
rect 918 322 924 323
rect 1062 327 1068 328
rect 1062 323 1063 327
rect 1067 323 1068 327
rect 1062 322 1068 323
rect 1206 327 1212 328
rect 1206 323 1207 327
rect 1211 323 1212 327
rect 1206 322 1212 323
rect 1350 327 1356 328
rect 1350 323 1351 327
rect 1355 323 1356 327
rect 1350 322 1356 323
rect 1494 327 1500 328
rect 1494 323 1495 327
rect 1499 323 1500 327
rect 1494 322 1500 323
rect 1638 327 1644 328
rect 1638 323 1639 327
rect 1643 323 1644 327
rect 2006 324 2007 328
rect 2011 324 2012 328
rect 2006 323 2012 324
rect 1638 322 1644 323
rect 2048 321 2050 341
rect 2046 320 2052 321
rect 2496 320 2498 341
rect 2640 320 2642 341
rect 2800 320 2802 341
rect 2960 320 2962 341
rect 3120 320 3122 341
rect 3272 320 3274 341
rect 3424 320 3426 341
rect 3568 320 3570 341
rect 3712 320 3714 341
rect 3840 320 3842 341
rect 3944 321 3946 341
rect 3942 320 3948 321
rect 2046 316 2047 320
rect 2051 316 2052 320
rect 2046 315 2052 316
rect 2494 319 2500 320
rect 2494 315 2495 319
rect 2499 315 2500 319
rect 2494 314 2500 315
rect 2638 319 2644 320
rect 2638 315 2639 319
rect 2643 315 2644 319
rect 2638 314 2644 315
rect 2798 319 2804 320
rect 2798 315 2799 319
rect 2803 315 2804 319
rect 2798 314 2804 315
rect 2958 319 2964 320
rect 2958 315 2959 319
rect 2963 315 2964 319
rect 2958 314 2964 315
rect 3118 319 3124 320
rect 3118 315 3119 319
rect 3123 315 3124 319
rect 3118 314 3124 315
rect 3270 319 3276 320
rect 3270 315 3271 319
rect 3275 315 3276 319
rect 3270 314 3276 315
rect 3422 319 3428 320
rect 3422 315 3423 319
rect 3427 315 3428 319
rect 3422 314 3428 315
rect 3566 319 3572 320
rect 3566 315 3567 319
rect 3571 315 3572 319
rect 3566 314 3572 315
rect 3710 319 3716 320
rect 3710 315 3711 319
rect 3715 315 3716 319
rect 3710 314 3716 315
rect 3838 319 3844 320
rect 3838 315 3839 319
rect 3843 315 3844 319
rect 3942 316 3943 320
rect 3947 316 3948 320
rect 3942 315 3948 316
rect 3838 314 3844 315
rect 110 311 116 312
rect 110 307 111 311
rect 115 307 116 311
rect 2006 311 2012 312
rect 110 306 116 307
rect 326 308 332 309
rect 112 271 114 306
rect 326 304 327 308
rect 331 304 332 308
rect 326 303 332 304
rect 462 308 468 309
rect 462 304 463 308
rect 467 304 468 308
rect 462 303 468 304
rect 614 308 620 309
rect 614 304 615 308
rect 619 304 620 308
rect 614 303 620 304
rect 766 308 772 309
rect 766 304 767 308
rect 771 304 772 308
rect 766 303 772 304
rect 918 308 924 309
rect 918 304 919 308
rect 923 304 924 308
rect 918 303 924 304
rect 1062 308 1068 309
rect 1062 304 1063 308
rect 1067 304 1068 308
rect 1062 303 1068 304
rect 1206 308 1212 309
rect 1206 304 1207 308
rect 1211 304 1212 308
rect 1206 303 1212 304
rect 1350 308 1356 309
rect 1350 304 1351 308
rect 1355 304 1356 308
rect 1350 303 1356 304
rect 1494 308 1500 309
rect 1494 304 1495 308
rect 1499 304 1500 308
rect 1494 303 1500 304
rect 1638 308 1644 309
rect 1638 304 1639 308
rect 1643 304 1644 308
rect 2006 307 2007 311
rect 2011 307 2012 311
rect 2006 306 2012 307
rect 1638 303 1644 304
rect 328 271 330 303
rect 464 271 466 303
rect 616 271 618 303
rect 768 271 770 303
rect 920 271 922 303
rect 1064 271 1066 303
rect 1208 271 1210 303
rect 1352 271 1354 303
rect 1496 271 1498 303
rect 1640 271 1642 303
rect 2008 271 2010 306
rect 2046 303 2052 304
rect 2046 299 2047 303
rect 2051 299 2052 303
rect 3942 303 3948 304
rect 2046 298 2052 299
rect 2494 300 2500 301
rect 2048 271 2050 298
rect 2494 296 2495 300
rect 2499 296 2500 300
rect 2494 295 2500 296
rect 2638 300 2644 301
rect 2638 296 2639 300
rect 2643 296 2644 300
rect 2638 295 2644 296
rect 2798 300 2804 301
rect 2798 296 2799 300
rect 2803 296 2804 300
rect 2798 295 2804 296
rect 2958 300 2964 301
rect 2958 296 2959 300
rect 2963 296 2964 300
rect 2958 295 2964 296
rect 3118 300 3124 301
rect 3118 296 3119 300
rect 3123 296 3124 300
rect 3118 295 3124 296
rect 3270 300 3276 301
rect 3270 296 3271 300
rect 3275 296 3276 300
rect 3270 295 3276 296
rect 3422 300 3428 301
rect 3422 296 3423 300
rect 3427 296 3428 300
rect 3422 295 3428 296
rect 3566 300 3572 301
rect 3566 296 3567 300
rect 3571 296 3572 300
rect 3566 295 3572 296
rect 3710 300 3716 301
rect 3710 296 3711 300
rect 3715 296 3716 300
rect 3710 295 3716 296
rect 3838 300 3844 301
rect 3838 296 3839 300
rect 3843 296 3844 300
rect 3942 299 3943 303
rect 3947 299 3948 303
rect 3942 298 3948 299
rect 3838 295 3844 296
rect 2496 271 2498 295
rect 2640 271 2642 295
rect 2800 271 2802 295
rect 2960 271 2962 295
rect 3120 271 3122 295
rect 3272 271 3274 295
rect 3424 271 3426 295
rect 3568 271 3570 295
rect 3712 271 3714 295
rect 3840 271 3842 295
rect 3944 271 3946 298
rect 111 270 115 271
rect 111 265 115 266
rect 167 270 171 271
rect 167 265 171 266
rect 327 270 331 271
rect 327 265 331 266
rect 463 270 467 271
rect 463 265 467 266
rect 503 270 507 271
rect 503 265 507 266
rect 615 270 619 271
rect 615 265 619 266
rect 687 270 691 271
rect 687 265 691 266
rect 767 270 771 271
rect 767 265 771 266
rect 871 270 875 271
rect 871 265 875 266
rect 919 270 923 271
rect 919 265 923 266
rect 1047 270 1051 271
rect 1047 265 1051 266
rect 1063 270 1067 271
rect 1063 265 1067 266
rect 1207 270 1211 271
rect 1207 265 1211 266
rect 1215 270 1219 271
rect 1215 265 1219 266
rect 1351 270 1355 271
rect 1351 265 1355 266
rect 1367 270 1371 271
rect 1367 265 1371 266
rect 1495 270 1499 271
rect 1495 265 1499 266
rect 1511 270 1515 271
rect 1511 265 1515 266
rect 1639 270 1643 271
rect 1639 265 1643 266
rect 1647 270 1651 271
rect 1647 265 1651 266
rect 1783 270 1787 271
rect 1783 265 1787 266
rect 1903 270 1907 271
rect 1903 265 1907 266
rect 2007 270 2011 271
rect 2007 265 2011 266
rect 2047 270 2051 271
rect 2047 265 2051 266
rect 2071 270 2075 271
rect 2071 265 2075 266
rect 2271 270 2275 271
rect 2271 265 2275 266
rect 2495 270 2499 271
rect 2495 265 2499 266
rect 2639 270 2643 271
rect 2639 265 2643 266
rect 2703 270 2707 271
rect 2703 265 2707 266
rect 2799 270 2803 271
rect 2799 265 2803 266
rect 2903 270 2907 271
rect 2903 265 2907 266
rect 2959 270 2963 271
rect 2959 265 2963 266
rect 3095 270 3099 271
rect 3095 265 3099 266
rect 3119 270 3123 271
rect 3119 265 3123 266
rect 3271 270 3275 271
rect 3271 265 3275 266
rect 3287 270 3291 271
rect 3287 265 3291 266
rect 3423 270 3427 271
rect 3423 265 3427 266
rect 3479 270 3483 271
rect 3479 265 3483 266
rect 3567 270 3571 271
rect 3567 265 3571 266
rect 3671 270 3675 271
rect 3671 265 3675 266
rect 3711 270 3715 271
rect 3711 265 3715 266
rect 3839 270 3843 271
rect 3839 265 3843 266
rect 3943 270 3947 271
rect 3943 265 3947 266
rect 112 238 114 265
rect 168 241 170 265
rect 328 241 330 265
rect 504 241 506 265
rect 688 241 690 265
rect 872 241 874 265
rect 1048 241 1050 265
rect 1216 241 1218 265
rect 1368 241 1370 265
rect 1512 241 1514 265
rect 1648 241 1650 265
rect 1784 241 1786 265
rect 1904 241 1906 265
rect 166 240 172 241
rect 110 237 116 238
rect 110 233 111 237
rect 115 233 116 237
rect 166 236 167 240
rect 171 236 172 240
rect 166 235 172 236
rect 326 240 332 241
rect 326 236 327 240
rect 331 236 332 240
rect 326 235 332 236
rect 502 240 508 241
rect 502 236 503 240
rect 507 236 508 240
rect 502 235 508 236
rect 686 240 692 241
rect 686 236 687 240
rect 691 236 692 240
rect 686 235 692 236
rect 870 240 876 241
rect 870 236 871 240
rect 875 236 876 240
rect 870 235 876 236
rect 1046 240 1052 241
rect 1046 236 1047 240
rect 1051 236 1052 240
rect 1046 235 1052 236
rect 1214 240 1220 241
rect 1214 236 1215 240
rect 1219 236 1220 240
rect 1214 235 1220 236
rect 1366 240 1372 241
rect 1366 236 1367 240
rect 1371 236 1372 240
rect 1366 235 1372 236
rect 1510 240 1516 241
rect 1510 236 1511 240
rect 1515 236 1516 240
rect 1510 235 1516 236
rect 1646 240 1652 241
rect 1646 236 1647 240
rect 1651 236 1652 240
rect 1646 235 1652 236
rect 1782 240 1788 241
rect 1782 236 1783 240
rect 1787 236 1788 240
rect 1782 235 1788 236
rect 1902 240 1908 241
rect 1902 236 1903 240
rect 1907 236 1908 240
rect 2008 238 2010 265
rect 2048 238 2050 265
rect 2072 241 2074 265
rect 2272 241 2274 265
rect 2496 241 2498 265
rect 2704 241 2706 265
rect 2904 241 2906 265
rect 3096 241 3098 265
rect 3288 241 3290 265
rect 3480 241 3482 265
rect 3672 241 3674 265
rect 3840 241 3842 265
rect 2070 240 2076 241
rect 1902 235 1908 236
rect 2006 237 2012 238
rect 110 232 116 233
rect 2006 233 2007 237
rect 2011 233 2012 237
rect 2006 232 2012 233
rect 2046 237 2052 238
rect 2046 233 2047 237
rect 2051 233 2052 237
rect 2070 236 2071 240
rect 2075 236 2076 240
rect 2070 235 2076 236
rect 2270 240 2276 241
rect 2270 236 2271 240
rect 2275 236 2276 240
rect 2270 235 2276 236
rect 2494 240 2500 241
rect 2494 236 2495 240
rect 2499 236 2500 240
rect 2494 235 2500 236
rect 2702 240 2708 241
rect 2702 236 2703 240
rect 2707 236 2708 240
rect 2702 235 2708 236
rect 2902 240 2908 241
rect 2902 236 2903 240
rect 2907 236 2908 240
rect 2902 235 2908 236
rect 3094 240 3100 241
rect 3094 236 3095 240
rect 3099 236 3100 240
rect 3094 235 3100 236
rect 3286 240 3292 241
rect 3286 236 3287 240
rect 3291 236 3292 240
rect 3286 235 3292 236
rect 3478 240 3484 241
rect 3478 236 3479 240
rect 3483 236 3484 240
rect 3478 235 3484 236
rect 3670 240 3676 241
rect 3670 236 3671 240
rect 3675 236 3676 240
rect 3670 235 3676 236
rect 3838 240 3844 241
rect 3838 236 3839 240
rect 3843 236 3844 240
rect 3944 238 3946 265
rect 3838 235 3844 236
rect 3942 237 3948 238
rect 2046 232 2052 233
rect 3942 233 3943 237
rect 3947 233 3948 237
rect 3942 232 3948 233
rect 166 221 172 222
rect 110 220 116 221
rect 110 216 111 220
rect 115 216 116 220
rect 166 217 167 221
rect 171 217 172 221
rect 166 216 172 217
rect 326 221 332 222
rect 326 217 327 221
rect 331 217 332 221
rect 326 216 332 217
rect 502 221 508 222
rect 502 217 503 221
rect 507 217 508 221
rect 502 216 508 217
rect 686 221 692 222
rect 686 217 687 221
rect 691 217 692 221
rect 686 216 692 217
rect 870 221 876 222
rect 870 217 871 221
rect 875 217 876 221
rect 870 216 876 217
rect 1046 221 1052 222
rect 1046 217 1047 221
rect 1051 217 1052 221
rect 1046 216 1052 217
rect 1214 221 1220 222
rect 1214 217 1215 221
rect 1219 217 1220 221
rect 1214 216 1220 217
rect 1366 221 1372 222
rect 1366 217 1367 221
rect 1371 217 1372 221
rect 1366 216 1372 217
rect 1510 221 1516 222
rect 1510 217 1511 221
rect 1515 217 1516 221
rect 1510 216 1516 217
rect 1646 221 1652 222
rect 1646 217 1647 221
rect 1651 217 1652 221
rect 1646 216 1652 217
rect 1782 221 1788 222
rect 1782 217 1783 221
rect 1787 217 1788 221
rect 1782 216 1788 217
rect 1902 221 1908 222
rect 2070 221 2076 222
rect 1902 217 1903 221
rect 1907 217 1908 221
rect 1902 216 1908 217
rect 2006 220 2012 221
rect 2006 216 2007 220
rect 2011 216 2012 220
rect 110 215 116 216
rect 112 167 114 215
rect 168 167 170 216
rect 328 167 330 216
rect 504 167 506 216
rect 688 167 690 216
rect 872 167 874 216
rect 1048 167 1050 216
rect 1216 167 1218 216
rect 1368 167 1370 216
rect 1512 167 1514 216
rect 1648 167 1650 216
rect 1784 167 1786 216
rect 1904 167 1906 216
rect 2006 215 2012 216
rect 2046 220 2052 221
rect 2046 216 2047 220
rect 2051 216 2052 220
rect 2070 217 2071 221
rect 2075 217 2076 221
rect 2070 216 2076 217
rect 2270 221 2276 222
rect 2270 217 2271 221
rect 2275 217 2276 221
rect 2270 216 2276 217
rect 2494 221 2500 222
rect 2494 217 2495 221
rect 2499 217 2500 221
rect 2494 216 2500 217
rect 2702 221 2708 222
rect 2702 217 2703 221
rect 2707 217 2708 221
rect 2702 216 2708 217
rect 2902 221 2908 222
rect 2902 217 2903 221
rect 2907 217 2908 221
rect 2902 216 2908 217
rect 3094 221 3100 222
rect 3094 217 3095 221
rect 3099 217 3100 221
rect 3094 216 3100 217
rect 3286 221 3292 222
rect 3286 217 3287 221
rect 3291 217 3292 221
rect 3286 216 3292 217
rect 3478 221 3484 222
rect 3478 217 3479 221
rect 3483 217 3484 221
rect 3478 216 3484 217
rect 3670 221 3676 222
rect 3670 217 3671 221
rect 3675 217 3676 221
rect 3670 216 3676 217
rect 3838 221 3844 222
rect 3838 217 3839 221
rect 3843 217 3844 221
rect 3838 216 3844 217
rect 3942 220 3948 221
rect 3942 216 3943 220
rect 3947 216 3948 220
rect 2046 215 2052 216
rect 2008 167 2010 215
rect 2048 171 2050 215
rect 2072 171 2074 216
rect 2272 171 2274 216
rect 2496 171 2498 216
rect 2704 171 2706 216
rect 2904 171 2906 216
rect 3096 171 3098 216
rect 3288 171 3290 216
rect 3480 171 3482 216
rect 3672 171 3674 216
rect 3840 171 3842 216
rect 3942 215 3948 216
rect 3944 171 3946 215
rect 2047 170 2051 171
rect 111 166 115 167
rect 111 161 115 162
rect 135 166 139 167
rect 135 161 139 162
rect 167 166 171 167
rect 167 161 171 162
rect 231 166 235 167
rect 231 161 235 162
rect 327 166 331 167
rect 327 161 331 162
rect 423 166 427 167
rect 423 161 427 162
rect 503 166 507 167
rect 503 161 507 162
rect 527 166 531 167
rect 527 161 531 162
rect 647 166 651 167
rect 647 161 651 162
rect 687 166 691 167
rect 687 161 691 162
rect 775 166 779 167
rect 775 161 779 162
rect 871 166 875 167
rect 871 161 875 162
rect 903 166 907 167
rect 903 161 907 162
rect 1031 166 1035 167
rect 1031 161 1035 162
rect 1047 166 1051 167
rect 1047 161 1051 162
rect 1151 166 1155 167
rect 1151 161 1155 162
rect 1215 166 1219 167
rect 1215 161 1219 162
rect 1271 166 1275 167
rect 1271 161 1275 162
rect 1367 166 1371 167
rect 1367 161 1371 162
rect 1383 166 1387 167
rect 1383 161 1387 162
rect 1487 166 1491 167
rect 1487 161 1491 162
rect 1511 166 1515 167
rect 1511 161 1515 162
rect 1591 166 1595 167
rect 1591 161 1595 162
rect 1647 166 1651 167
rect 1647 161 1651 162
rect 1703 166 1707 167
rect 1703 161 1707 162
rect 1783 166 1787 167
rect 1783 161 1787 162
rect 1807 166 1811 167
rect 1807 161 1811 162
rect 1903 166 1907 167
rect 1903 161 1907 162
rect 2007 166 2011 167
rect 2047 165 2051 166
rect 2071 170 2075 171
rect 2071 165 2075 166
rect 2167 170 2171 171
rect 2167 165 2171 166
rect 2263 170 2267 171
rect 2263 165 2267 166
rect 2271 170 2275 171
rect 2271 165 2275 166
rect 2359 170 2363 171
rect 2359 165 2363 166
rect 2455 170 2459 171
rect 2455 165 2459 166
rect 2495 170 2499 171
rect 2495 165 2499 166
rect 2551 170 2555 171
rect 2551 165 2555 166
rect 2655 170 2659 171
rect 2655 165 2659 166
rect 2703 170 2707 171
rect 2703 165 2707 166
rect 2759 170 2763 171
rect 2759 165 2763 166
rect 2863 170 2867 171
rect 2863 165 2867 166
rect 2903 170 2907 171
rect 2903 165 2907 166
rect 2975 170 2979 171
rect 2975 165 2979 166
rect 3095 170 3099 171
rect 3095 165 3099 166
rect 3103 170 3107 171
rect 3103 165 3107 166
rect 3239 170 3243 171
rect 3239 165 3243 166
rect 3287 170 3291 171
rect 3287 165 3291 166
rect 3383 170 3387 171
rect 3383 165 3387 166
rect 3479 170 3483 171
rect 3479 165 3483 166
rect 3535 170 3539 171
rect 3535 165 3539 166
rect 3671 170 3675 171
rect 3671 165 3675 166
rect 3695 170 3699 171
rect 3695 165 3699 166
rect 3839 170 3843 171
rect 3839 165 3843 166
rect 3943 170 3947 171
rect 3943 165 3947 166
rect 2007 161 2011 162
rect 112 141 114 161
rect 110 140 116 141
rect 136 140 138 161
rect 232 140 234 161
rect 328 140 330 161
rect 424 140 426 161
rect 528 140 530 161
rect 648 140 650 161
rect 776 140 778 161
rect 904 140 906 161
rect 1032 140 1034 161
rect 1152 140 1154 161
rect 1272 140 1274 161
rect 1384 140 1386 161
rect 1488 140 1490 161
rect 1592 140 1594 161
rect 1704 140 1706 161
rect 1808 140 1810 161
rect 1904 140 1906 161
rect 2008 141 2010 161
rect 2048 145 2050 165
rect 2046 144 2052 145
rect 2072 144 2074 165
rect 2168 144 2170 165
rect 2264 144 2266 165
rect 2360 144 2362 165
rect 2456 144 2458 165
rect 2552 144 2554 165
rect 2656 144 2658 165
rect 2760 144 2762 165
rect 2864 144 2866 165
rect 2976 144 2978 165
rect 3104 144 3106 165
rect 3240 144 3242 165
rect 3384 144 3386 165
rect 3536 144 3538 165
rect 3696 144 3698 165
rect 3840 144 3842 165
rect 3944 145 3946 165
rect 3942 144 3948 145
rect 2006 140 2012 141
rect 110 136 111 140
rect 115 136 116 140
rect 110 135 116 136
rect 134 139 140 140
rect 134 135 135 139
rect 139 135 140 139
rect 134 134 140 135
rect 230 139 236 140
rect 230 135 231 139
rect 235 135 236 139
rect 230 134 236 135
rect 326 139 332 140
rect 326 135 327 139
rect 331 135 332 139
rect 326 134 332 135
rect 422 139 428 140
rect 422 135 423 139
rect 427 135 428 139
rect 422 134 428 135
rect 526 139 532 140
rect 526 135 527 139
rect 531 135 532 139
rect 526 134 532 135
rect 646 139 652 140
rect 646 135 647 139
rect 651 135 652 139
rect 646 134 652 135
rect 774 139 780 140
rect 774 135 775 139
rect 779 135 780 139
rect 774 134 780 135
rect 902 139 908 140
rect 902 135 903 139
rect 907 135 908 139
rect 902 134 908 135
rect 1030 139 1036 140
rect 1030 135 1031 139
rect 1035 135 1036 139
rect 1030 134 1036 135
rect 1150 139 1156 140
rect 1150 135 1151 139
rect 1155 135 1156 139
rect 1150 134 1156 135
rect 1270 139 1276 140
rect 1270 135 1271 139
rect 1275 135 1276 139
rect 1270 134 1276 135
rect 1382 139 1388 140
rect 1382 135 1383 139
rect 1387 135 1388 139
rect 1382 134 1388 135
rect 1486 139 1492 140
rect 1486 135 1487 139
rect 1491 135 1492 139
rect 1486 134 1492 135
rect 1590 139 1596 140
rect 1590 135 1591 139
rect 1595 135 1596 139
rect 1590 134 1596 135
rect 1702 139 1708 140
rect 1702 135 1703 139
rect 1707 135 1708 139
rect 1702 134 1708 135
rect 1806 139 1812 140
rect 1806 135 1807 139
rect 1811 135 1812 139
rect 1806 134 1812 135
rect 1902 139 1908 140
rect 1902 135 1903 139
rect 1907 135 1908 139
rect 2006 136 2007 140
rect 2011 136 2012 140
rect 2046 140 2047 144
rect 2051 140 2052 144
rect 2046 139 2052 140
rect 2070 143 2076 144
rect 2070 139 2071 143
rect 2075 139 2076 143
rect 2070 138 2076 139
rect 2166 143 2172 144
rect 2166 139 2167 143
rect 2171 139 2172 143
rect 2166 138 2172 139
rect 2262 143 2268 144
rect 2262 139 2263 143
rect 2267 139 2268 143
rect 2262 138 2268 139
rect 2358 143 2364 144
rect 2358 139 2359 143
rect 2363 139 2364 143
rect 2358 138 2364 139
rect 2454 143 2460 144
rect 2454 139 2455 143
rect 2459 139 2460 143
rect 2454 138 2460 139
rect 2550 143 2556 144
rect 2550 139 2551 143
rect 2555 139 2556 143
rect 2550 138 2556 139
rect 2654 143 2660 144
rect 2654 139 2655 143
rect 2659 139 2660 143
rect 2654 138 2660 139
rect 2758 143 2764 144
rect 2758 139 2759 143
rect 2763 139 2764 143
rect 2758 138 2764 139
rect 2862 143 2868 144
rect 2862 139 2863 143
rect 2867 139 2868 143
rect 2862 138 2868 139
rect 2974 143 2980 144
rect 2974 139 2975 143
rect 2979 139 2980 143
rect 2974 138 2980 139
rect 3102 143 3108 144
rect 3102 139 3103 143
rect 3107 139 3108 143
rect 3102 138 3108 139
rect 3238 143 3244 144
rect 3238 139 3239 143
rect 3243 139 3244 143
rect 3238 138 3244 139
rect 3382 143 3388 144
rect 3382 139 3383 143
rect 3387 139 3388 143
rect 3382 138 3388 139
rect 3534 143 3540 144
rect 3534 139 3535 143
rect 3539 139 3540 143
rect 3534 138 3540 139
rect 3694 143 3700 144
rect 3694 139 3695 143
rect 3699 139 3700 143
rect 3694 138 3700 139
rect 3838 143 3844 144
rect 3838 139 3839 143
rect 3843 139 3844 143
rect 3942 140 3943 144
rect 3947 140 3948 144
rect 3942 139 3948 140
rect 3838 138 3844 139
rect 2006 135 2012 136
rect 1902 134 1908 135
rect 2046 127 2052 128
rect 110 123 116 124
rect 110 119 111 123
rect 115 119 116 123
rect 2006 123 2012 124
rect 110 118 116 119
rect 134 120 140 121
rect 112 91 114 118
rect 134 116 135 120
rect 139 116 140 120
rect 134 115 140 116
rect 230 120 236 121
rect 230 116 231 120
rect 235 116 236 120
rect 230 115 236 116
rect 326 120 332 121
rect 326 116 327 120
rect 331 116 332 120
rect 326 115 332 116
rect 422 120 428 121
rect 422 116 423 120
rect 427 116 428 120
rect 422 115 428 116
rect 526 120 532 121
rect 526 116 527 120
rect 531 116 532 120
rect 526 115 532 116
rect 646 120 652 121
rect 646 116 647 120
rect 651 116 652 120
rect 646 115 652 116
rect 774 120 780 121
rect 774 116 775 120
rect 779 116 780 120
rect 774 115 780 116
rect 902 120 908 121
rect 902 116 903 120
rect 907 116 908 120
rect 902 115 908 116
rect 1030 120 1036 121
rect 1030 116 1031 120
rect 1035 116 1036 120
rect 1030 115 1036 116
rect 1150 120 1156 121
rect 1150 116 1151 120
rect 1155 116 1156 120
rect 1150 115 1156 116
rect 1270 120 1276 121
rect 1270 116 1271 120
rect 1275 116 1276 120
rect 1270 115 1276 116
rect 1382 120 1388 121
rect 1382 116 1383 120
rect 1387 116 1388 120
rect 1382 115 1388 116
rect 1486 120 1492 121
rect 1486 116 1487 120
rect 1491 116 1492 120
rect 1486 115 1492 116
rect 1590 120 1596 121
rect 1590 116 1591 120
rect 1595 116 1596 120
rect 1590 115 1596 116
rect 1702 120 1708 121
rect 1702 116 1703 120
rect 1707 116 1708 120
rect 1702 115 1708 116
rect 1806 120 1812 121
rect 1806 116 1807 120
rect 1811 116 1812 120
rect 1806 115 1812 116
rect 1902 120 1908 121
rect 1902 116 1903 120
rect 1907 116 1908 120
rect 2006 119 2007 123
rect 2011 119 2012 123
rect 2046 123 2047 127
rect 2051 123 2052 127
rect 3942 127 3948 128
rect 2046 122 2052 123
rect 2070 124 2076 125
rect 2006 118 2012 119
rect 1902 115 1908 116
rect 136 91 138 115
rect 232 91 234 115
rect 328 91 330 115
rect 424 91 426 115
rect 528 91 530 115
rect 648 91 650 115
rect 776 91 778 115
rect 904 91 906 115
rect 1032 91 1034 115
rect 1152 91 1154 115
rect 1272 91 1274 115
rect 1384 91 1386 115
rect 1488 91 1490 115
rect 1592 91 1594 115
rect 1704 91 1706 115
rect 1808 91 1810 115
rect 1904 91 1906 115
rect 2008 91 2010 118
rect 2048 95 2050 122
rect 2070 120 2071 124
rect 2075 120 2076 124
rect 2070 119 2076 120
rect 2166 124 2172 125
rect 2166 120 2167 124
rect 2171 120 2172 124
rect 2166 119 2172 120
rect 2262 124 2268 125
rect 2262 120 2263 124
rect 2267 120 2268 124
rect 2262 119 2268 120
rect 2358 124 2364 125
rect 2358 120 2359 124
rect 2363 120 2364 124
rect 2358 119 2364 120
rect 2454 124 2460 125
rect 2454 120 2455 124
rect 2459 120 2460 124
rect 2454 119 2460 120
rect 2550 124 2556 125
rect 2550 120 2551 124
rect 2555 120 2556 124
rect 2550 119 2556 120
rect 2654 124 2660 125
rect 2654 120 2655 124
rect 2659 120 2660 124
rect 2654 119 2660 120
rect 2758 124 2764 125
rect 2758 120 2759 124
rect 2763 120 2764 124
rect 2758 119 2764 120
rect 2862 124 2868 125
rect 2862 120 2863 124
rect 2867 120 2868 124
rect 2862 119 2868 120
rect 2974 124 2980 125
rect 2974 120 2975 124
rect 2979 120 2980 124
rect 2974 119 2980 120
rect 3102 124 3108 125
rect 3102 120 3103 124
rect 3107 120 3108 124
rect 3102 119 3108 120
rect 3238 124 3244 125
rect 3238 120 3239 124
rect 3243 120 3244 124
rect 3238 119 3244 120
rect 3382 124 3388 125
rect 3382 120 3383 124
rect 3387 120 3388 124
rect 3382 119 3388 120
rect 3534 124 3540 125
rect 3534 120 3535 124
rect 3539 120 3540 124
rect 3534 119 3540 120
rect 3694 124 3700 125
rect 3694 120 3695 124
rect 3699 120 3700 124
rect 3694 119 3700 120
rect 3838 124 3844 125
rect 3838 120 3839 124
rect 3843 120 3844 124
rect 3942 123 3943 127
rect 3947 123 3948 127
rect 3942 122 3948 123
rect 3838 119 3844 120
rect 2072 95 2074 119
rect 2168 95 2170 119
rect 2264 95 2266 119
rect 2360 95 2362 119
rect 2456 95 2458 119
rect 2552 95 2554 119
rect 2656 95 2658 119
rect 2760 95 2762 119
rect 2864 95 2866 119
rect 2976 95 2978 119
rect 3104 95 3106 119
rect 3240 95 3242 119
rect 3384 95 3386 119
rect 3536 95 3538 119
rect 3696 95 3698 119
rect 3840 95 3842 119
rect 3944 95 3946 122
rect 2047 94 2051 95
rect 111 90 115 91
rect 111 85 115 86
rect 135 90 139 91
rect 135 85 139 86
rect 231 90 235 91
rect 231 85 235 86
rect 327 90 331 91
rect 327 85 331 86
rect 423 90 427 91
rect 423 85 427 86
rect 527 90 531 91
rect 527 85 531 86
rect 647 90 651 91
rect 647 85 651 86
rect 775 90 779 91
rect 775 85 779 86
rect 903 90 907 91
rect 903 85 907 86
rect 1031 90 1035 91
rect 1031 85 1035 86
rect 1151 90 1155 91
rect 1151 85 1155 86
rect 1271 90 1275 91
rect 1271 85 1275 86
rect 1383 90 1387 91
rect 1383 85 1387 86
rect 1487 90 1491 91
rect 1487 85 1491 86
rect 1591 90 1595 91
rect 1591 85 1595 86
rect 1703 90 1707 91
rect 1703 85 1707 86
rect 1807 90 1811 91
rect 1807 85 1811 86
rect 1903 90 1907 91
rect 1903 85 1907 86
rect 2007 90 2011 91
rect 2047 89 2051 90
rect 2071 94 2075 95
rect 2071 89 2075 90
rect 2167 94 2171 95
rect 2167 89 2171 90
rect 2263 94 2267 95
rect 2263 89 2267 90
rect 2359 94 2363 95
rect 2359 89 2363 90
rect 2455 94 2459 95
rect 2455 89 2459 90
rect 2551 94 2555 95
rect 2551 89 2555 90
rect 2655 94 2659 95
rect 2655 89 2659 90
rect 2759 94 2763 95
rect 2759 89 2763 90
rect 2863 94 2867 95
rect 2863 89 2867 90
rect 2975 94 2979 95
rect 2975 89 2979 90
rect 3103 94 3107 95
rect 3103 89 3107 90
rect 3239 94 3243 95
rect 3239 89 3243 90
rect 3383 94 3387 95
rect 3383 89 3387 90
rect 3535 94 3539 95
rect 3535 89 3539 90
rect 3695 94 3699 95
rect 3695 89 3699 90
rect 3839 94 3843 95
rect 3839 89 3843 90
rect 3943 94 3947 95
rect 3943 89 3947 90
rect 2007 85 2011 86
<< m4c >>
rect 111 4026 115 4030
rect 1519 4026 1523 4030
rect 1615 4026 1619 4030
rect 1711 4026 1715 4030
rect 1807 4026 1811 4030
rect 1903 4026 1907 4030
rect 2007 4026 2011 4030
rect 2047 4014 2051 4018
rect 2071 4014 2075 4018
rect 2167 4014 2171 4018
rect 2263 4014 2267 4018
rect 3943 4014 3947 4018
rect 111 3950 115 3954
rect 199 3950 203 3954
rect 295 3950 299 3954
rect 391 3950 395 3954
rect 495 3950 499 3954
rect 615 3950 619 3954
rect 743 3950 747 3954
rect 871 3950 875 3954
rect 999 3950 1003 3954
rect 1127 3950 1131 3954
rect 1255 3950 1259 3954
rect 1383 3950 1387 3954
rect 1511 3950 1515 3954
rect 1519 3950 1523 3954
rect 1615 3950 1619 3954
rect 1647 3950 1651 3954
rect 1711 3950 1715 3954
rect 1807 3950 1811 3954
rect 1903 3950 1907 3954
rect 2007 3950 2011 3954
rect 2047 3938 2051 3942
rect 2071 3938 2075 3942
rect 2159 3938 2163 3942
rect 2167 3938 2171 3942
rect 2263 3938 2267 3942
rect 2287 3938 2291 3942
rect 2415 3938 2419 3942
rect 2551 3938 2555 3942
rect 2687 3938 2691 3942
rect 2823 3938 2827 3942
rect 2951 3938 2955 3942
rect 3071 3938 3075 3942
rect 3191 3938 3195 3942
rect 3303 3938 3307 3942
rect 3407 3938 3411 3942
rect 3519 3938 3523 3942
rect 3631 3938 3635 3942
rect 3743 3938 3747 3942
rect 3943 3938 3947 3942
rect 111 3874 115 3878
rect 199 3874 203 3878
rect 295 3874 299 3878
rect 335 3874 339 3878
rect 391 3874 395 3878
rect 455 3874 459 3878
rect 495 3874 499 3878
rect 583 3874 587 3878
rect 615 3874 619 3878
rect 719 3874 723 3878
rect 743 3874 747 3878
rect 847 3874 851 3878
rect 871 3874 875 3878
rect 975 3874 979 3878
rect 999 3874 1003 3878
rect 1103 3874 1107 3878
rect 1127 3874 1131 3878
rect 1231 3874 1235 3878
rect 1255 3874 1259 3878
rect 1359 3874 1363 3878
rect 1383 3874 1387 3878
rect 1487 3874 1491 3878
rect 1511 3874 1515 3878
rect 1647 3874 1651 3878
rect 2007 3874 2011 3878
rect 2047 3854 2051 3858
rect 2159 3854 2163 3858
rect 2207 3854 2211 3858
rect 2287 3854 2291 3858
rect 2343 3854 2347 3858
rect 2415 3854 2419 3858
rect 2487 3854 2491 3858
rect 2551 3854 2555 3858
rect 2647 3854 2651 3858
rect 2687 3854 2691 3858
rect 2823 3854 2827 3858
rect 2951 3854 2955 3858
rect 3015 3854 3019 3858
rect 3071 3854 3075 3858
rect 3191 3854 3195 3858
rect 3223 3854 3227 3858
rect 3303 3854 3307 3858
rect 3407 3854 3411 3858
rect 3439 3854 3443 3858
rect 3519 3854 3523 3858
rect 3631 3854 3635 3858
rect 3655 3854 3659 3858
rect 3743 3854 3747 3858
rect 3943 3854 3947 3858
rect 111 3794 115 3798
rect 335 3794 339 3798
rect 455 3794 459 3798
rect 503 3794 507 3798
rect 583 3794 587 3798
rect 615 3794 619 3798
rect 719 3794 723 3798
rect 735 3794 739 3798
rect 847 3794 851 3798
rect 863 3794 867 3798
rect 975 3794 979 3798
rect 999 3794 1003 3798
rect 1103 3794 1107 3798
rect 1143 3794 1147 3798
rect 1231 3794 1235 3798
rect 1287 3794 1291 3798
rect 1359 3794 1363 3798
rect 1431 3794 1435 3798
rect 1487 3794 1491 3798
rect 1583 3794 1587 3798
rect 2007 3794 2011 3798
rect 2047 3778 2051 3782
rect 2191 3778 2195 3782
rect 2207 3778 2211 3782
rect 2343 3778 2347 3782
rect 2375 3778 2379 3782
rect 2487 3778 2491 3782
rect 2559 3778 2563 3782
rect 2647 3778 2651 3782
rect 2743 3778 2747 3782
rect 2823 3778 2827 3782
rect 2935 3778 2939 3782
rect 3015 3778 3019 3782
rect 3127 3778 3131 3782
rect 3223 3778 3227 3782
rect 3319 3778 3323 3782
rect 3439 3778 3443 3782
rect 3511 3778 3515 3782
rect 3655 3778 3659 3782
rect 3711 3778 3715 3782
rect 3943 3778 3947 3782
rect 111 3710 115 3714
rect 495 3710 499 3714
rect 503 3710 507 3714
rect 591 3710 595 3714
rect 615 3710 619 3714
rect 687 3710 691 3714
rect 735 3710 739 3714
rect 791 3710 795 3714
rect 863 3710 867 3714
rect 911 3710 915 3714
rect 999 3710 1003 3714
rect 1039 3710 1043 3714
rect 1143 3710 1147 3714
rect 1183 3710 1187 3714
rect 1287 3710 1291 3714
rect 1335 3710 1339 3714
rect 1431 3710 1435 3714
rect 1495 3710 1499 3714
rect 1583 3710 1587 3714
rect 1655 3710 1659 3714
rect 2007 3710 2011 3714
rect 2047 3698 2051 3702
rect 2127 3698 2131 3702
rect 2191 3698 2195 3702
rect 2351 3698 2355 3702
rect 2375 3698 2379 3702
rect 2559 3698 2563 3702
rect 2583 3698 2587 3702
rect 2743 3698 2747 3702
rect 2815 3698 2819 3702
rect 2935 3698 2939 3702
rect 3047 3698 3051 3702
rect 3127 3698 3131 3702
rect 3279 3698 3283 3702
rect 3319 3698 3323 3702
rect 3511 3698 3515 3702
rect 3711 3698 3715 3702
rect 3751 3698 3755 3702
rect 3943 3698 3947 3702
rect 111 3626 115 3630
rect 335 3626 339 3630
rect 463 3626 467 3630
rect 495 3626 499 3630
rect 591 3626 595 3630
rect 607 3626 611 3630
rect 687 3626 691 3630
rect 759 3626 763 3630
rect 791 3626 795 3630
rect 911 3626 915 3630
rect 927 3626 931 3630
rect 1039 3626 1043 3630
rect 1095 3626 1099 3630
rect 1183 3626 1187 3630
rect 1263 3626 1267 3630
rect 1335 3626 1339 3630
rect 1439 3626 1443 3630
rect 1495 3626 1499 3630
rect 1615 3626 1619 3630
rect 1655 3626 1659 3630
rect 1791 3626 1795 3630
rect 2007 3626 2011 3630
rect 2047 3614 2051 3618
rect 2127 3614 2131 3618
rect 2191 3614 2195 3618
rect 2327 3614 2331 3618
rect 2351 3614 2355 3618
rect 2455 3614 2459 3618
rect 2583 3614 2587 3618
rect 2719 3614 2723 3618
rect 2815 3614 2819 3618
rect 2855 3614 2859 3618
rect 2999 3614 3003 3618
rect 3047 3614 3051 3618
rect 3143 3614 3147 3618
rect 3279 3614 3283 3618
rect 3295 3614 3299 3618
rect 3455 3614 3459 3618
rect 3511 3614 3515 3618
rect 3623 3614 3627 3618
rect 3751 3614 3755 3618
rect 3943 3614 3947 3618
rect 111 3538 115 3542
rect 159 3538 163 3542
rect 303 3538 307 3542
rect 335 3538 339 3542
rect 463 3538 467 3542
rect 607 3538 611 3542
rect 639 3538 643 3542
rect 759 3538 763 3542
rect 815 3538 819 3542
rect 927 3538 931 3542
rect 999 3538 1003 3542
rect 1095 3538 1099 3542
rect 1175 3538 1179 3542
rect 1263 3538 1267 3542
rect 1351 3538 1355 3542
rect 1439 3538 1443 3542
rect 1527 3538 1531 3542
rect 1615 3538 1619 3542
rect 1703 3538 1707 3542
rect 1791 3538 1795 3542
rect 1879 3538 1883 3542
rect 2007 3538 2011 3542
rect 2047 3538 2051 3542
rect 2103 3538 2107 3542
rect 2191 3538 2195 3542
rect 2271 3538 2275 3542
rect 2327 3538 2331 3542
rect 2447 3538 2451 3542
rect 2455 3538 2459 3542
rect 2583 3538 2587 3542
rect 2631 3538 2635 3542
rect 2719 3538 2723 3542
rect 2815 3538 2819 3542
rect 2855 3538 2859 3542
rect 2999 3538 3003 3542
rect 3143 3538 3147 3542
rect 3175 3538 3179 3542
rect 3295 3538 3299 3542
rect 3351 3538 3355 3542
rect 3455 3538 3459 3542
rect 3519 3538 3523 3542
rect 3623 3538 3627 3542
rect 3687 3538 3691 3542
rect 3839 3538 3843 3542
rect 3943 3538 3947 3542
rect 111 3454 115 3458
rect 135 3454 139 3458
rect 159 3454 163 3458
rect 303 3454 307 3458
rect 319 3454 323 3458
rect 463 3454 467 3458
rect 535 3454 539 3458
rect 639 3454 643 3458
rect 751 3454 755 3458
rect 815 3454 819 3458
rect 959 3454 963 3458
rect 999 3454 1003 3458
rect 1159 3454 1163 3458
rect 1175 3454 1179 3458
rect 1351 3454 1355 3458
rect 1527 3454 1531 3458
rect 1535 3454 1539 3458
rect 1703 3454 1707 3458
rect 1719 3454 1723 3458
rect 1879 3454 1883 3458
rect 1903 3454 1907 3458
rect 2007 3454 2011 3458
rect 2047 3458 2051 3462
rect 2103 3458 2107 3462
rect 2127 3458 2131 3462
rect 2271 3458 2275 3462
rect 2311 3458 2315 3462
rect 2447 3458 2451 3462
rect 2495 3458 2499 3462
rect 2631 3458 2635 3462
rect 2679 3458 2683 3462
rect 2815 3458 2819 3462
rect 2863 3458 2867 3462
rect 2999 3458 3003 3462
rect 3047 3458 3051 3462
rect 3175 3458 3179 3462
rect 3223 3458 3227 3462
rect 3351 3458 3355 3462
rect 3407 3458 3411 3462
rect 3519 3458 3523 3462
rect 3591 3458 3595 3462
rect 3687 3458 3691 3462
rect 3775 3458 3779 3462
rect 3839 3458 3843 3462
rect 3943 3458 3947 3462
rect 111 3378 115 3382
rect 135 3378 139 3382
rect 231 3378 235 3382
rect 319 3378 323 3382
rect 375 3378 379 3382
rect 535 3378 539 3382
rect 703 3378 707 3382
rect 751 3378 755 3382
rect 871 3378 875 3382
rect 959 3378 963 3382
rect 1047 3378 1051 3382
rect 1159 3378 1163 3382
rect 1215 3378 1219 3382
rect 1351 3378 1355 3382
rect 1383 3378 1387 3382
rect 1535 3378 1539 3382
rect 1543 3378 1547 3382
rect 1703 3378 1707 3382
rect 1719 3378 1723 3382
rect 1871 3378 1875 3382
rect 1903 3378 1907 3382
rect 2007 3378 2011 3382
rect 2047 3366 2051 3370
rect 2071 3366 2075 3370
rect 2127 3366 2131 3370
rect 2215 3366 2219 3370
rect 2311 3366 2315 3370
rect 2359 3366 2363 3370
rect 2495 3366 2499 3370
rect 2511 3366 2515 3370
rect 2655 3366 2659 3370
rect 2679 3366 2683 3370
rect 2799 3366 2803 3370
rect 2863 3366 2867 3370
rect 2935 3366 2939 3370
rect 3047 3366 3051 3370
rect 3079 3366 3083 3370
rect 3223 3366 3227 3370
rect 3375 3366 3379 3370
rect 3407 3366 3411 3370
rect 3535 3366 3539 3370
rect 3591 3366 3595 3370
rect 3695 3366 3699 3370
rect 3775 3366 3779 3370
rect 3839 3366 3843 3370
rect 3943 3366 3947 3370
rect 111 3302 115 3306
rect 135 3302 139 3306
rect 231 3302 235 3306
rect 279 3302 283 3306
rect 375 3302 379 3306
rect 463 3302 467 3306
rect 535 3302 539 3306
rect 663 3302 667 3306
rect 703 3302 707 3306
rect 871 3302 875 3306
rect 1047 3302 1051 3306
rect 1079 3302 1083 3306
rect 1215 3302 1219 3306
rect 1295 3302 1299 3306
rect 1383 3302 1387 3306
rect 1519 3302 1523 3306
rect 1543 3302 1547 3306
rect 1703 3302 1707 3306
rect 1743 3302 1747 3306
rect 1871 3302 1875 3306
rect 2007 3302 2011 3306
rect 2047 3282 2051 3286
rect 2071 3282 2075 3286
rect 2111 3282 2115 3286
rect 2215 3282 2219 3286
rect 2247 3282 2251 3286
rect 2359 3282 2363 3286
rect 2399 3282 2403 3286
rect 2511 3282 2515 3286
rect 2575 3282 2579 3286
rect 2655 3282 2659 3286
rect 2783 3282 2787 3286
rect 2799 3282 2803 3286
rect 2935 3282 2939 3286
rect 3015 3282 3019 3286
rect 3079 3282 3083 3286
rect 3223 3282 3227 3286
rect 3263 3282 3267 3286
rect 3375 3282 3379 3286
rect 3527 3282 3531 3286
rect 3535 3282 3539 3286
rect 3695 3282 3699 3286
rect 3791 3282 3795 3286
rect 3839 3282 3843 3286
rect 3943 3282 3947 3286
rect 111 3226 115 3230
rect 135 3226 139 3230
rect 279 3226 283 3230
rect 287 3226 291 3230
rect 447 3226 451 3230
rect 463 3226 467 3230
rect 615 3226 619 3230
rect 663 3226 667 3230
rect 791 3226 795 3230
rect 871 3226 875 3230
rect 967 3226 971 3230
rect 1079 3226 1083 3230
rect 1143 3226 1147 3230
rect 1295 3226 1299 3230
rect 1327 3226 1331 3230
rect 1511 3226 1515 3230
rect 1519 3226 1523 3230
rect 1695 3226 1699 3230
rect 1743 3226 1747 3230
rect 2007 3226 2011 3230
rect 2047 3206 2051 3210
rect 2071 3206 2075 3210
rect 2111 3206 2115 3210
rect 2167 3206 2171 3210
rect 2247 3206 2251 3210
rect 2263 3206 2267 3210
rect 2359 3206 2363 3210
rect 2399 3206 2403 3210
rect 2455 3206 2459 3210
rect 2551 3206 2555 3210
rect 2575 3206 2579 3210
rect 2647 3206 2651 3210
rect 2743 3206 2747 3210
rect 2783 3206 2787 3210
rect 2839 3206 2843 3210
rect 2935 3206 2939 3210
rect 3015 3206 3019 3210
rect 3031 3206 3035 3210
rect 3127 3206 3131 3210
rect 3223 3206 3227 3210
rect 3263 3206 3267 3210
rect 3319 3206 3323 3210
rect 3439 3206 3443 3210
rect 3527 3206 3531 3210
rect 3575 3206 3579 3210
rect 3719 3206 3723 3210
rect 3791 3206 3795 3210
rect 3839 3206 3843 3210
rect 3943 3206 3947 3210
rect 111 3146 115 3150
rect 135 3146 139 3150
rect 287 3146 291 3150
rect 311 3146 315 3150
rect 439 3146 443 3150
rect 447 3146 451 3150
rect 583 3146 587 3150
rect 615 3146 619 3150
rect 743 3146 747 3150
rect 791 3146 795 3150
rect 903 3146 907 3150
rect 967 3146 971 3150
rect 1063 3146 1067 3150
rect 1143 3146 1147 3150
rect 1223 3146 1227 3150
rect 1327 3146 1331 3150
rect 1391 3146 1395 3150
rect 1511 3146 1515 3150
rect 1559 3146 1563 3150
rect 1695 3146 1699 3150
rect 1727 3146 1731 3150
rect 2007 3146 2011 3150
rect 2047 3118 2051 3122
rect 2071 3118 2075 3122
rect 2167 3118 2171 3122
rect 2263 3118 2267 3122
rect 2335 3118 2339 3122
rect 2359 3118 2363 3122
rect 2455 3118 2459 3122
rect 2551 3118 2555 3122
rect 2623 3118 2627 3122
rect 2647 3118 2651 3122
rect 2743 3118 2747 3122
rect 2839 3118 2843 3122
rect 2911 3118 2915 3122
rect 2935 3118 2939 3122
rect 3031 3118 3035 3122
rect 3127 3118 3131 3122
rect 3207 3118 3211 3122
rect 3223 3118 3227 3122
rect 3319 3118 3323 3122
rect 3439 3118 3443 3122
rect 3503 3118 3507 3122
rect 3575 3118 3579 3122
rect 3719 3118 3723 3122
rect 3799 3118 3803 3122
rect 3839 3118 3843 3122
rect 3943 3118 3947 3122
rect 111 3062 115 3066
rect 311 3062 315 3066
rect 439 3062 443 3066
rect 503 3062 507 3066
rect 583 3062 587 3066
rect 599 3062 603 3066
rect 703 3062 707 3066
rect 743 3062 747 3066
rect 815 3062 819 3066
rect 903 3062 907 3066
rect 935 3062 939 3066
rect 1063 3062 1067 3066
rect 1071 3062 1075 3066
rect 1223 3062 1227 3066
rect 1383 3062 1387 3066
rect 1391 3062 1395 3066
rect 1551 3062 1555 3066
rect 1559 3062 1563 3066
rect 1719 3062 1723 3066
rect 1727 3062 1731 3066
rect 2007 3062 2011 3066
rect 2047 3042 2051 3046
rect 2071 3042 2075 3046
rect 2335 3042 2339 3046
rect 2383 3042 2387 3046
rect 2623 3042 2627 3046
rect 2703 3042 2707 3046
rect 2911 3042 2915 3046
rect 2999 3042 3003 3046
rect 3207 3042 3211 3046
rect 3287 3042 3291 3046
rect 3503 3042 3507 3046
rect 3575 3042 3579 3046
rect 3799 3042 3803 3046
rect 3839 3042 3843 3046
rect 3943 3042 3947 3046
rect 111 2982 115 2986
rect 503 2982 507 2986
rect 551 2982 555 2986
rect 599 2982 603 2986
rect 647 2982 651 2986
rect 703 2982 707 2986
rect 759 2982 763 2986
rect 815 2982 819 2986
rect 887 2982 891 2986
rect 935 2982 939 2986
rect 1023 2982 1027 2986
rect 1071 2982 1075 2986
rect 1175 2982 1179 2986
rect 1223 2982 1227 2986
rect 1327 2982 1331 2986
rect 1383 2982 1387 2986
rect 1487 2982 1491 2986
rect 1551 2982 1555 2986
rect 1655 2982 1659 2986
rect 1719 2982 1723 2986
rect 1823 2982 1827 2986
rect 2007 2982 2011 2986
rect 2047 2962 2051 2966
rect 2071 2962 2075 2966
rect 2383 2962 2387 2966
rect 2391 2962 2395 2966
rect 2703 2962 2707 2966
rect 2975 2962 2979 2966
rect 2999 2962 3003 2966
rect 3215 2962 3219 2966
rect 3287 2962 3291 2966
rect 3439 2962 3443 2966
rect 3575 2962 3579 2966
rect 3647 2962 3651 2966
rect 3839 2962 3843 2966
rect 3943 2962 3947 2966
rect 111 2898 115 2902
rect 471 2898 475 2902
rect 551 2898 555 2902
rect 575 2898 579 2902
rect 647 2898 651 2902
rect 695 2898 699 2902
rect 759 2898 763 2902
rect 839 2898 843 2902
rect 887 2898 891 2902
rect 991 2898 995 2902
rect 1023 2898 1027 2902
rect 1151 2898 1155 2902
rect 1175 2898 1179 2902
rect 1319 2898 1323 2902
rect 1327 2898 1331 2902
rect 1487 2898 1491 2902
rect 1495 2898 1499 2902
rect 1655 2898 1659 2902
rect 1671 2898 1675 2902
rect 1823 2898 1827 2902
rect 1847 2898 1851 2902
rect 2007 2898 2011 2902
rect 2047 2886 2051 2890
rect 2071 2886 2075 2890
rect 2295 2886 2299 2890
rect 2391 2886 2395 2890
rect 2535 2886 2539 2890
rect 2703 2886 2707 2890
rect 2767 2886 2771 2890
rect 2975 2886 2979 2890
rect 2991 2886 2995 2890
rect 3215 2886 3219 2890
rect 3431 2886 3435 2890
rect 3439 2886 3443 2890
rect 3647 2886 3651 2890
rect 3839 2886 3843 2890
rect 3943 2886 3947 2890
rect 111 2818 115 2822
rect 471 2818 475 2822
rect 479 2818 483 2822
rect 575 2818 579 2822
rect 679 2818 683 2822
rect 695 2818 699 2822
rect 799 2818 803 2822
rect 839 2818 843 2822
rect 935 2818 939 2822
rect 991 2818 995 2822
rect 1079 2818 1083 2822
rect 1151 2818 1155 2822
rect 1239 2818 1243 2822
rect 1319 2818 1323 2822
rect 1415 2818 1419 2822
rect 1495 2818 1499 2822
rect 1599 2818 1603 2822
rect 1671 2818 1675 2822
rect 1783 2818 1787 2822
rect 1847 2818 1851 2822
rect 2007 2818 2011 2822
rect 2047 2806 2051 2810
rect 2071 2806 2075 2810
rect 2199 2806 2203 2810
rect 2295 2806 2299 2810
rect 2367 2806 2371 2810
rect 2535 2806 2539 2810
rect 2551 2806 2555 2810
rect 2735 2806 2739 2810
rect 2767 2806 2771 2810
rect 2927 2806 2931 2810
rect 2991 2806 2995 2810
rect 3111 2806 3115 2810
rect 3215 2806 3219 2810
rect 3295 2806 3299 2810
rect 3431 2806 3435 2810
rect 3479 2806 3483 2810
rect 3647 2806 3651 2810
rect 3671 2806 3675 2810
rect 3839 2806 3843 2810
rect 3943 2806 3947 2810
rect 111 2738 115 2742
rect 479 2738 483 2742
rect 511 2738 515 2742
rect 575 2738 579 2742
rect 623 2738 627 2742
rect 679 2738 683 2742
rect 743 2738 747 2742
rect 799 2738 803 2742
rect 879 2738 883 2742
rect 935 2738 939 2742
rect 1015 2738 1019 2742
rect 1079 2738 1083 2742
rect 1159 2738 1163 2742
rect 1239 2738 1243 2742
rect 1311 2738 1315 2742
rect 1415 2738 1419 2742
rect 1463 2738 1467 2742
rect 1599 2738 1603 2742
rect 1623 2738 1627 2742
rect 1783 2738 1787 2742
rect 2007 2738 2011 2742
rect 2047 2726 2051 2730
rect 2071 2726 2075 2730
rect 2191 2726 2195 2730
rect 2199 2726 2203 2730
rect 2319 2726 2323 2730
rect 2367 2726 2371 2730
rect 2447 2726 2451 2730
rect 2551 2726 2555 2730
rect 2583 2726 2587 2730
rect 2727 2726 2731 2730
rect 2735 2726 2739 2730
rect 2887 2726 2891 2730
rect 2927 2726 2931 2730
rect 3063 2726 3067 2730
rect 3111 2726 3115 2730
rect 3255 2726 3259 2730
rect 3295 2726 3299 2730
rect 3455 2726 3459 2730
rect 3479 2726 3483 2730
rect 3655 2726 3659 2730
rect 3671 2726 3675 2730
rect 3839 2726 3843 2730
rect 3943 2726 3947 2730
rect 111 2658 115 2662
rect 367 2658 371 2662
rect 487 2658 491 2662
rect 511 2658 515 2662
rect 615 2658 619 2662
rect 623 2658 627 2662
rect 743 2658 747 2662
rect 751 2658 755 2662
rect 879 2658 883 2662
rect 895 2658 899 2662
rect 1015 2658 1019 2662
rect 1031 2658 1035 2662
rect 1159 2658 1163 2662
rect 1167 2658 1171 2662
rect 1303 2658 1307 2662
rect 1311 2658 1315 2662
rect 1431 2658 1435 2662
rect 1463 2658 1467 2662
rect 1567 2658 1571 2662
rect 1623 2658 1627 2662
rect 1703 2658 1707 2662
rect 1783 2658 1787 2662
rect 2007 2658 2011 2662
rect 2047 2642 2051 2646
rect 2071 2642 2075 2646
rect 2191 2642 2195 2646
rect 2231 2642 2235 2646
rect 2319 2642 2323 2646
rect 2335 2642 2339 2646
rect 2447 2642 2451 2646
rect 2559 2642 2563 2646
rect 2583 2642 2587 2646
rect 2671 2642 2675 2646
rect 2727 2642 2731 2646
rect 2791 2642 2795 2646
rect 2887 2642 2891 2646
rect 2911 2642 2915 2646
rect 3031 2642 3035 2646
rect 3063 2642 3067 2646
rect 3151 2642 3155 2646
rect 3255 2642 3259 2646
rect 3455 2642 3459 2646
rect 3655 2642 3659 2646
rect 3839 2642 3843 2646
rect 3943 2642 3947 2646
rect 111 2582 115 2586
rect 135 2582 139 2586
rect 287 2582 291 2586
rect 367 2582 371 2586
rect 447 2582 451 2586
rect 487 2582 491 2586
rect 607 2582 611 2586
rect 615 2582 619 2586
rect 751 2582 755 2586
rect 767 2582 771 2586
rect 895 2582 899 2586
rect 919 2582 923 2586
rect 1031 2582 1035 2586
rect 1063 2582 1067 2586
rect 1167 2582 1171 2586
rect 1199 2582 1203 2586
rect 1303 2582 1307 2586
rect 1335 2582 1339 2586
rect 1431 2582 1435 2586
rect 1463 2582 1467 2586
rect 1567 2582 1571 2586
rect 1591 2582 1595 2586
rect 1703 2582 1707 2586
rect 1727 2582 1731 2586
rect 2007 2582 2011 2586
rect 2047 2562 2051 2566
rect 2231 2562 2235 2566
rect 2335 2562 2339 2566
rect 2383 2562 2387 2566
rect 2447 2562 2451 2566
rect 2495 2562 2499 2566
rect 2559 2562 2563 2566
rect 2615 2562 2619 2566
rect 2671 2562 2675 2566
rect 2743 2562 2747 2566
rect 2791 2562 2795 2566
rect 2871 2562 2875 2566
rect 2911 2562 2915 2566
rect 2991 2562 2995 2566
rect 3031 2562 3035 2566
rect 3111 2562 3115 2566
rect 3151 2562 3155 2566
rect 3231 2562 3235 2566
rect 3359 2562 3363 2566
rect 3487 2562 3491 2566
rect 3943 2562 3947 2566
rect 111 2490 115 2494
rect 135 2490 139 2494
rect 231 2490 235 2494
rect 287 2490 291 2494
rect 327 2490 331 2494
rect 423 2490 427 2494
rect 447 2490 451 2494
rect 519 2490 523 2494
rect 607 2490 611 2494
rect 767 2490 771 2494
rect 919 2490 923 2494
rect 1063 2490 1067 2494
rect 1199 2490 1203 2494
rect 1335 2490 1339 2494
rect 1463 2490 1467 2494
rect 1591 2490 1595 2494
rect 1727 2490 1731 2494
rect 2007 2490 2011 2494
rect 2047 2482 2051 2486
rect 2383 2482 2387 2486
rect 2495 2482 2499 2486
rect 2535 2482 2539 2486
rect 2615 2482 2619 2486
rect 2711 2482 2715 2486
rect 2743 2482 2747 2486
rect 2871 2482 2875 2486
rect 2879 2482 2883 2486
rect 2991 2482 2995 2486
rect 3047 2482 3051 2486
rect 3111 2482 3115 2486
rect 3207 2482 3211 2486
rect 3231 2482 3235 2486
rect 3359 2482 3363 2486
rect 3487 2482 3491 2486
rect 3503 2482 3507 2486
rect 3655 2482 3659 2486
rect 3807 2482 3811 2486
rect 3943 2482 3947 2486
rect 111 2398 115 2402
rect 135 2398 139 2402
rect 231 2398 235 2402
rect 255 2398 259 2402
rect 327 2398 331 2402
rect 415 2398 419 2402
rect 423 2398 427 2402
rect 519 2398 523 2402
rect 575 2398 579 2402
rect 735 2398 739 2402
rect 887 2398 891 2402
rect 1039 2398 1043 2402
rect 1183 2398 1187 2402
rect 1327 2398 1331 2402
rect 1479 2398 1483 2402
rect 2007 2398 2011 2402
rect 2047 2394 2051 2398
rect 2535 2394 2539 2398
rect 2607 2394 2611 2398
rect 2711 2394 2715 2398
rect 2815 2394 2819 2398
rect 2879 2394 2883 2398
rect 3007 2394 3011 2398
rect 3047 2394 3051 2398
rect 3191 2394 3195 2398
rect 3207 2394 3211 2398
rect 3359 2394 3363 2398
rect 3503 2394 3507 2398
rect 3519 2394 3523 2398
rect 3655 2394 3659 2398
rect 3679 2394 3683 2398
rect 3807 2394 3811 2398
rect 3839 2394 3843 2398
rect 3943 2394 3947 2398
rect 111 2322 115 2326
rect 135 2322 139 2326
rect 255 2322 259 2326
rect 263 2322 267 2326
rect 415 2322 419 2326
rect 423 2322 427 2326
rect 575 2322 579 2326
rect 583 2322 587 2326
rect 735 2322 739 2326
rect 743 2322 747 2326
rect 887 2322 891 2326
rect 895 2322 899 2326
rect 1039 2322 1043 2326
rect 1047 2322 1051 2326
rect 1183 2322 1187 2326
rect 1199 2322 1203 2326
rect 1327 2322 1331 2326
rect 1351 2322 1355 2326
rect 1479 2322 1483 2326
rect 1503 2322 1507 2326
rect 2007 2322 2011 2326
rect 2047 2302 2051 2306
rect 2071 2302 2075 2306
rect 2167 2302 2171 2306
rect 2271 2302 2275 2306
rect 2415 2302 2419 2306
rect 2575 2302 2579 2306
rect 2607 2302 2611 2306
rect 2743 2302 2747 2306
rect 2815 2302 2819 2306
rect 2911 2302 2915 2306
rect 3007 2302 3011 2306
rect 3071 2302 3075 2306
rect 3191 2302 3195 2306
rect 3231 2302 3235 2306
rect 3359 2302 3363 2306
rect 3383 2302 3387 2306
rect 3519 2302 3523 2306
rect 3535 2302 3539 2306
rect 3679 2302 3683 2306
rect 3695 2302 3699 2306
rect 3839 2302 3843 2306
rect 3943 2302 3947 2306
rect 111 2242 115 2246
rect 135 2242 139 2246
rect 223 2242 227 2246
rect 263 2242 267 2246
rect 351 2242 355 2246
rect 423 2242 427 2246
rect 495 2242 499 2246
rect 583 2242 587 2246
rect 647 2242 651 2246
rect 743 2242 747 2246
rect 799 2242 803 2246
rect 895 2242 899 2246
rect 959 2242 963 2246
rect 1047 2242 1051 2246
rect 1119 2242 1123 2246
rect 1199 2242 1203 2246
rect 1279 2242 1283 2246
rect 1351 2242 1355 2246
rect 1439 2242 1443 2246
rect 1503 2242 1507 2246
rect 1599 2242 1603 2246
rect 2007 2242 2011 2246
rect 2047 2226 2051 2230
rect 2071 2226 2075 2230
rect 2167 2226 2171 2230
rect 2175 2226 2179 2230
rect 2271 2226 2275 2230
rect 2319 2226 2323 2230
rect 2415 2226 2419 2230
rect 2471 2226 2475 2230
rect 2575 2226 2579 2230
rect 2623 2226 2627 2230
rect 2743 2226 2747 2230
rect 2783 2226 2787 2230
rect 2911 2226 2915 2230
rect 2935 2226 2939 2230
rect 3071 2226 3075 2230
rect 3079 2226 3083 2230
rect 3223 2226 3227 2230
rect 3231 2226 3235 2230
rect 3367 2226 3371 2230
rect 3383 2226 3387 2230
rect 3519 2226 3523 2230
rect 3535 2226 3539 2230
rect 3695 2226 3699 2230
rect 3943 2226 3947 2230
rect 111 2166 115 2170
rect 223 2166 227 2170
rect 351 2166 355 2170
rect 471 2166 475 2170
rect 495 2166 499 2170
rect 567 2166 571 2170
rect 647 2166 651 2170
rect 679 2166 683 2170
rect 799 2166 803 2170
rect 807 2166 811 2170
rect 943 2166 947 2170
rect 959 2166 963 2170
rect 1079 2166 1083 2170
rect 1119 2166 1123 2170
rect 1223 2166 1227 2170
rect 1279 2166 1283 2170
rect 1367 2166 1371 2170
rect 1439 2166 1443 2170
rect 1503 2166 1507 2170
rect 1599 2166 1603 2170
rect 1639 2166 1643 2170
rect 1783 2166 1787 2170
rect 1903 2166 1907 2170
rect 2007 2166 2011 2170
rect 2047 2130 2051 2134
rect 2071 2130 2075 2134
rect 2175 2130 2179 2134
rect 2279 2130 2283 2134
rect 2319 2130 2323 2134
rect 2391 2130 2395 2134
rect 2471 2130 2475 2134
rect 2511 2130 2515 2134
rect 2623 2130 2627 2134
rect 2631 2130 2635 2134
rect 2759 2130 2763 2134
rect 2783 2130 2787 2134
rect 2895 2130 2899 2134
rect 2935 2130 2939 2134
rect 3039 2130 3043 2134
rect 3079 2130 3083 2134
rect 3191 2130 3195 2134
rect 3223 2130 3227 2134
rect 3351 2130 3355 2134
rect 3367 2130 3371 2134
rect 3519 2130 3523 2134
rect 3687 2130 3691 2134
rect 3839 2130 3843 2134
rect 3943 2130 3947 2134
rect 111 2090 115 2094
rect 471 2090 475 2094
rect 567 2090 571 2094
rect 623 2090 627 2094
rect 679 2090 683 2094
rect 735 2090 739 2094
rect 807 2090 811 2094
rect 855 2090 859 2094
rect 943 2090 947 2094
rect 983 2090 987 2094
rect 1079 2090 1083 2094
rect 1119 2090 1123 2094
rect 1223 2090 1227 2094
rect 1255 2090 1259 2094
rect 1367 2090 1371 2094
rect 1391 2090 1395 2094
rect 1503 2090 1507 2094
rect 1527 2090 1531 2094
rect 1639 2090 1643 2094
rect 1655 2090 1659 2094
rect 1783 2090 1787 2094
rect 1791 2090 1795 2094
rect 1903 2090 1907 2094
rect 2007 2090 2011 2094
rect 2047 2046 2051 2050
rect 2279 2046 2283 2050
rect 2327 2046 2331 2050
rect 2391 2046 2395 2050
rect 2431 2046 2435 2050
rect 2511 2046 2515 2050
rect 2535 2046 2539 2050
rect 2631 2046 2635 2050
rect 2647 2046 2651 2050
rect 2759 2046 2763 2050
rect 2775 2046 2779 2050
rect 2895 2046 2899 2050
rect 2919 2046 2923 2050
rect 3039 2046 3043 2050
rect 3079 2046 3083 2050
rect 3191 2046 3195 2050
rect 3263 2046 3267 2050
rect 3351 2046 3355 2050
rect 3455 2046 3459 2050
rect 3519 2046 3523 2050
rect 3655 2046 3659 2050
rect 3687 2046 3691 2050
rect 3839 2046 3843 2050
rect 3943 2046 3947 2050
rect 111 2010 115 2014
rect 447 2010 451 2014
rect 575 2010 579 2014
rect 623 2010 627 2014
rect 727 2010 731 2014
rect 735 2010 739 2014
rect 855 2010 859 2014
rect 887 2010 891 2014
rect 983 2010 987 2014
rect 1055 2010 1059 2014
rect 1119 2010 1123 2014
rect 1231 2010 1235 2014
rect 1255 2010 1259 2014
rect 1391 2010 1395 2014
rect 1399 2010 1403 2014
rect 1527 2010 1531 2014
rect 1575 2010 1579 2014
rect 1655 2010 1659 2014
rect 1751 2010 1755 2014
rect 1791 2010 1795 2014
rect 1903 2010 1907 2014
rect 2007 2010 2011 2014
rect 2047 1966 2051 1970
rect 2255 1966 2259 1970
rect 2327 1966 2331 1970
rect 2351 1966 2355 1970
rect 2431 1966 2435 1970
rect 2447 1966 2451 1970
rect 2535 1966 2539 1970
rect 2543 1966 2547 1970
rect 2647 1966 2651 1970
rect 2767 1966 2771 1970
rect 2775 1966 2779 1970
rect 2919 1966 2923 1970
rect 3079 1966 3083 1970
rect 3103 1966 3107 1970
rect 3263 1966 3267 1970
rect 3319 1966 3323 1970
rect 3455 1966 3459 1970
rect 3543 1966 3547 1970
rect 3655 1966 3659 1970
rect 3775 1966 3779 1970
rect 3839 1966 3843 1970
rect 3943 1966 3947 1970
rect 111 1934 115 1938
rect 447 1934 451 1938
rect 575 1934 579 1938
rect 655 1934 659 1938
rect 727 1934 731 1938
rect 751 1934 755 1938
rect 847 1934 851 1938
rect 887 1934 891 1938
rect 943 1934 947 1938
rect 1039 1934 1043 1938
rect 1055 1934 1059 1938
rect 1135 1934 1139 1938
rect 1231 1934 1235 1938
rect 1327 1934 1331 1938
rect 1399 1934 1403 1938
rect 1423 1934 1427 1938
rect 1575 1934 1579 1938
rect 1751 1934 1755 1938
rect 1903 1934 1907 1938
rect 2007 1934 2011 1938
rect 2047 1878 2051 1882
rect 2183 1878 2187 1882
rect 2255 1878 2259 1882
rect 2279 1878 2283 1882
rect 2351 1878 2355 1882
rect 2383 1878 2387 1882
rect 2447 1878 2451 1882
rect 2487 1878 2491 1882
rect 2543 1878 2547 1882
rect 2591 1878 2595 1882
rect 2647 1878 2651 1882
rect 2703 1878 2707 1882
rect 2767 1878 2771 1882
rect 2831 1878 2835 1882
rect 2919 1878 2923 1882
rect 2991 1878 2995 1882
rect 3103 1878 3107 1882
rect 3183 1878 3187 1882
rect 3319 1878 3323 1882
rect 3399 1878 3403 1882
rect 3543 1878 3547 1882
rect 3631 1878 3635 1882
rect 3775 1878 3779 1882
rect 3839 1878 3843 1882
rect 3943 1878 3947 1882
rect 111 1858 115 1862
rect 319 1858 323 1862
rect 447 1858 451 1862
rect 583 1858 587 1862
rect 655 1858 659 1862
rect 719 1858 723 1862
rect 751 1858 755 1862
rect 847 1858 851 1862
rect 855 1858 859 1862
rect 943 1858 947 1862
rect 991 1858 995 1862
rect 1039 1858 1043 1862
rect 1127 1858 1131 1862
rect 1135 1858 1139 1862
rect 1231 1858 1235 1862
rect 1263 1858 1267 1862
rect 1327 1858 1331 1862
rect 1399 1858 1403 1862
rect 1423 1858 1427 1862
rect 1535 1858 1539 1862
rect 2007 1858 2011 1862
rect 2047 1798 2051 1802
rect 2127 1798 2131 1802
rect 2183 1798 2187 1802
rect 2279 1798 2283 1802
rect 2311 1798 2315 1802
rect 2383 1798 2387 1802
rect 2487 1798 2491 1802
rect 2495 1798 2499 1802
rect 2591 1798 2595 1802
rect 2687 1798 2691 1802
rect 2703 1798 2707 1802
rect 2831 1798 2835 1802
rect 2879 1798 2883 1802
rect 2991 1798 2995 1802
rect 3071 1798 3075 1802
rect 3183 1798 3187 1802
rect 3263 1798 3267 1802
rect 3399 1798 3403 1802
rect 3463 1798 3467 1802
rect 3631 1798 3635 1802
rect 3663 1798 3667 1802
rect 3839 1798 3843 1802
rect 3943 1798 3947 1802
rect 111 1778 115 1782
rect 255 1778 259 1782
rect 319 1778 323 1782
rect 391 1778 395 1782
rect 447 1778 451 1782
rect 535 1778 539 1782
rect 583 1778 587 1782
rect 695 1778 699 1782
rect 719 1778 723 1782
rect 855 1778 859 1782
rect 863 1778 867 1782
rect 991 1778 995 1782
rect 1031 1778 1035 1782
rect 1127 1778 1131 1782
rect 1207 1778 1211 1782
rect 1263 1778 1267 1782
rect 1383 1778 1387 1782
rect 1399 1778 1403 1782
rect 1535 1778 1539 1782
rect 1559 1778 1563 1782
rect 1743 1778 1747 1782
rect 2007 1778 2011 1782
rect 2047 1718 2051 1722
rect 2071 1718 2075 1722
rect 2127 1718 2131 1722
rect 2191 1718 2195 1722
rect 2311 1718 2315 1722
rect 2343 1718 2347 1722
rect 2495 1718 2499 1722
rect 2511 1718 2515 1722
rect 2687 1718 2691 1722
rect 2871 1718 2875 1722
rect 2879 1718 2883 1722
rect 3063 1718 3067 1722
rect 3071 1718 3075 1722
rect 3255 1718 3259 1722
rect 3263 1718 3267 1722
rect 3447 1718 3451 1722
rect 3463 1718 3467 1722
rect 3647 1718 3651 1722
rect 3663 1718 3667 1722
rect 3839 1718 3843 1722
rect 3943 1718 3947 1722
rect 111 1702 115 1706
rect 135 1702 139 1706
rect 255 1702 259 1706
rect 263 1702 267 1706
rect 391 1702 395 1706
rect 431 1702 435 1706
rect 535 1702 539 1706
rect 607 1702 611 1706
rect 695 1702 699 1706
rect 799 1702 803 1706
rect 863 1702 867 1706
rect 999 1702 1003 1706
rect 1031 1702 1035 1706
rect 1199 1702 1203 1706
rect 1207 1702 1211 1706
rect 1383 1702 1387 1706
rect 1407 1702 1411 1706
rect 1559 1702 1563 1706
rect 1623 1702 1627 1706
rect 1743 1702 1747 1706
rect 1839 1702 1843 1706
rect 2007 1702 2011 1706
rect 2047 1642 2051 1646
rect 2071 1642 2075 1646
rect 2191 1642 2195 1646
rect 2335 1642 2339 1646
rect 2343 1642 2347 1646
rect 2511 1642 2515 1646
rect 2599 1642 2603 1646
rect 2687 1642 2691 1646
rect 2839 1642 2843 1646
rect 2871 1642 2875 1646
rect 3047 1642 3051 1646
rect 3063 1642 3067 1646
rect 3231 1642 3235 1646
rect 3255 1642 3259 1646
rect 3399 1642 3403 1646
rect 3447 1642 3451 1646
rect 3551 1642 3555 1646
rect 3647 1642 3651 1646
rect 3695 1642 3699 1646
rect 3839 1642 3843 1646
rect 3943 1642 3947 1646
rect 111 1626 115 1630
rect 135 1626 139 1630
rect 263 1626 267 1630
rect 287 1626 291 1630
rect 431 1626 435 1630
rect 471 1626 475 1630
rect 607 1626 611 1630
rect 655 1626 659 1630
rect 799 1626 803 1630
rect 839 1626 843 1630
rect 999 1626 1003 1630
rect 1015 1626 1019 1630
rect 1183 1626 1187 1630
rect 1199 1626 1203 1630
rect 1343 1626 1347 1630
rect 1407 1626 1411 1630
rect 1495 1626 1499 1630
rect 1623 1626 1627 1630
rect 1639 1626 1643 1630
rect 1783 1626 1787 1630
rect 1839 1626 1843 1630
rect 1903 1626 1907 1630
rect 2007 1626 2011 1630
rect 2047 1562 2051 1566
rect 2071 1562 2075 1566
rect 2335 1562 2339 1566
rect 2583 1562 2587 1566
rect 2599 1562 2603 1566
rect 2743 1562 2747 1566
rect 2839 1562 2843 1566
rect 2903 1562 2907 1566
rect 3047 1562 3051 1566
rect 3063 1562 3067 1566
rect 3223 1562 3227 1566
rect 3231 1562 3235 1566
rect 3383 1562 3387 1566
rect 3399 1562 3403 1566
rect 3543 1562 3547 1566
rect 3551 1562 3555 1566
rect 3695 1562 3699 1566
rect 3703 1562 3707 1566
rect 3839 1562 3843 1566
rect 3943 1562 3947 1566
rect 111 1546 115 1550
rect 135 1546 139 1550
rect 287 1546 291 1550
rect 295 1546 299 1550
rect 471 1546 475 1550
rect 487 1546 491 1550
rect 655 1546 659 1550
rect 687 1546 691 1550
rect 839 1546 843 1550
rect 887 1546 891 1550
rect 1015 1546 1019 1550
rect 1079 1546 1083 1550
rect 1183 1546 1187 1550
rect 1263 1546 1267 1550
rect 1343 1546 1347 1550
rect 1447 1546 1451 1550
rect 1495 1546 1499 1550
rect 1623 1546 1627 1550
rect 1639 1546 1643 1550
rect 1783 1546 1787 1550
rect 1807 1546 1811 1550
rect 1903 1546 1907 1550
rect 2007 1546 2011 1550
rect 2047 1486 2051 1490
rect 2415 1486 2419 1490
rect 2511 1486 2515 1490
rect 2583 1486 2587 1490
rect 2607 1486 2611 1490
rect 2703 1486 2707 1490
rect 2743 1486 2747 1490
rect 2799 1486 2803 1490
rect 2903 1486 2907 1490
rect 2919 1486 2923 1490
rect 3063 1486 3067 1490
rect 3223 1486 3227 1490
rect 3231 1486 3235 1490
rect 3383 1486 3387 1490
rect 3415 1486 3419 1490
rect 3543 1486 3547 1490
rect 3615 1486 3619 1490
rect 3703 1486 3707 1490
rect 3815 1486 3819 1490
rect 3943 1486 3947 1490
rect 111 1470 115 1474
rect 135 1470 139 1474
rect 175 1470 179 1474
rect 295 1470 299 1474
rect 359 1470 363 1474
rect 487 1470 491 1474
rect 567 1470 571 1474
rect 687 1470 691 1474
rect 783 1470 787 1474
rect 887 1470 891 1474
rect 1007 1470 1011 1474
rect 1079 1470 1083 1474
rect 1231 1470 1235 1474
rect 1263 1470 1267 1474
rect 1447 1470 1451 1474
rect 1463 1470 1467 1474
rect 1623 1470 1627 1474
rect 1695 1470 1699 1474
rect 1807 1470 1811 1474
rect 1903 1470 1907 1474
rect 2007 1470 2011 1474
rect 111 1394 115 1398
rect 175 1394 179 1398
rect 327 1394 331 1398
rect 359 1394 363 1398
rect 463 1394 467 1398
rect 567 1394 571 1398
rect 599 1394 603 1398
rect 727 1394 731 1398
rect 783 1394 787 1398
rect 855 1394 859 1398
rect 983 1394 987 1398
rect 1007 1394 1011 1398
rect 1119 1394 1123 1398
rect 1231 1394 1235 1398
rect 1263 1394 1267 1398
rect 1423 1394 1427 1398
rect 1463 1394 1467 1398
rect 1583 1394 1587 1398
rect 1695 1394 1699 1398
rect 1751 1394 1755 1398
rect 1903 1394 1907 1398
rect 2007 1394 2011 1398
rect 2047 1390 2051 1394
rect 2071 1390 2075 1394
rect 2303 1390 2307 1394
rect 2415 1390 2419 1394
rect 2511 1390 2515 1394
rect 2559 1390 2563 1394
rect 2607 1390 2611 1394
rect 2703 1390 2707 1394
rect 2799 1390 2803 1394
rect 2807 1390 2811 1394
rect 2919 1390 2923 1394
rect 3055 1390 3059 1394
rect 3063 1390 3067 1394
rect 3231 1390 3235 1394
rect 3303 1390 3307 1394
rect 3415 1390 3419 1394
rect 3559 1390 3563 1394
rect 3615 1390 3619 1394
rect 3815 1390 3819 1394
rect 3943 1390 3947 1394
rect 111 1310 115 1314
rect 327 1310 331 1314
rect 463 1310 467 1314
rect 551 1310 555 1314
rect 599 1310 603 1314
rect 655 1310 659 1314
rect 727 1310 731 1314
rect 767 1310 771 1314
rect 855 1310 859 1314
rect 879 1310 883 1314
rect 983 1310 987 1314
rect 991 1310 995 1314
rect 1103 1310 1107 1314
rect 1119 1310 1123 1314
rect 1215 1310 1219 1314
rect 1263 1310 1267 1314
rect 1327 1310 1331 1314
rect 1423 1310 1427 1314
rect 1439 1310 1443 1314
rect 1559 1310 1563 1314
rect 1583 1310 1587 1314
rect 1751 1310 1755 1314
rect 1903 1310 1907 1314
rect 2007 1310 2011 1314
rect 2047 1306 2051 1310
rect 2071 1306 2075 1310
rect 2223 1306 2227 1310
rect 2303 1306 2307 1310
rect 2415 1306 2419 1310
rect 2559 1306 2563 1310
rect 2615 1306 2619 1310
rect 2807 1306 2811 1310
rect 2815 1306 2819 1310
rect 2999 1306 3003 1310
rect 3055 1306 3059 1310
rect 3175 1306 3179 1310
rect 3303 1306 3307 1310
rect 3343 1306 3347 1310
rect 3503 1306 3507 1310
rect 3559 1306 3563 1310
rect 3663 1306 3667 1310
rect 3815 1306 3819 1310
rect 3831 1306 3835 1310
rect 3943 1306 3947 1310
rect 111 1234 115 1238
rect 391 1234 395 1238
rect 519 1234 523 1238
rect 551 1234 555 1238
rect 655 1234 659 1238
rect 663 1234 667 1238
rect 767 1234 771 1238
rect 807 1234 811 1238
rect 879 1234 883 1238
rect 959 1234 963 1238
rect 991 1234 995 1238
rect 1103 1234 1107 1238
rect 1111 1234 1115 1238
rect 1215 1234 1219 1238
rect 1255 1234 1259 1238
rect 1327 1234 1331 1238
rect 1407 1234 1411 1238
rect 1439 1234 1443 1238
rect 1559 1234 1563 1238
rect 1711 1234 1715 1238
rect 2007 1234 2011 1238
rect 2047 1222 2051 1226
rect 2071 1222 2075 1226
rect 2135 1222 2139 1226
rect 2223 1222 2227 1226
rect 2311 1222 2315 1226
rect 2415 1222 2419 1226
rect 2503 1222 2507 1226
rect 2615 1222 2619 1226
rect 2695 1222 2699 1226
rect 2815 1222 2819 1226
rect 2887 1222 2891 1226
rect 2999 1222 3003 1226
rect 3071 1222 3075 1226
rect 3175 1222 3179 1226
rect 3239 1222 3243 1226
rect 3343 1222 3347 1226
rect 3399 1222 3403 1226
rect 3503 1222 3507 1226
rect 3551 1222 3555 1226
rect 3663 1222 3667 1226
rect 3703 1222 3707 1226
rect 3831 1222 3835 1226
rect 3839 1222 3843 1226
rect 3943 1222 3947 1226
rect 111 1154 115 1158
rect 175 1154 179 1158
rect 327 1154 331 1158
rect 391 1154 395 1158
rect 495 1154 499 1158
rect 519 1154 523 1158
rect 663 1154 667 1158
rect 671 1154 675 1158
rect 807 1154 811 1158
rect 847 1154 851 1158
rect 959 1154 963 1158
rect 1031 1154 1035 1158
rect 1111 1154 1115 1158
rect 1207 1154 1211 1158
rect 1255 1154 1259 1158
rect 1383 1154 1387 1158
rect 1407 1154 1411 1158
rect 1559 1154 1563 1158
rect 1567 1154 1571 1158
rect 1711 1154 1715 1158
rect 1751 1154 1755 1158
rect 2007 1154 2011 1158
rect 2047 1138 2051 1142
rect 2135 1138 2139 1142
rect 2295 1138 2299 1142
rect 2311 1138 2315 1142
rect 2423 1138 2427 1142
rect 2503 1138 2507 1142
rect 2559 1138 2563 1142
rect 2695 1138 2699 1142
rect 2839 1138 2843 1142
rect 2887 1138 2891 1142
rect 2991 1138 2995 1142
rect 3071 1138 3075 1142
rect 3151 1138 3155 1142
rect 3239 1138 3243 1142
rect 3319 1138 3323 1142
rect 3399 1138 3403 1142
rect 3495 1138 3499 1142
rect 3551 1138 3555 1142
rect 3679 1138 3683 1142
rect 3703 1138 3707 1142
rect 3839 1138 3843 1142
rect 3943 1138 3947 1142
rect 111 1070 115 1074
rect 135 1070 139 1074
rect 175 1070 179 1074
rect 231 1070 235 1074
rect 327 1070 331 1074
rect 375 1070 379 1074
rect 495 1070 499 1074
rect 543 1070 547 1074
rect 671 1070 675 1074
rect 727 1070 731 1074
rect 847 1070 851 1074
rect 911 1070 915 1074
rect 1031 1070 1035 1074
rect 1095 1070 1099 1074
rect 1207 1070 1211 1074
rect 1279 1070 1283 1074
rect 1383 1070 1387 1074
rect 1463 1070 1467 1074
rect 1567 1070 1571 1074
rect 1647 1070 1651 1074
rect 1751 1070 1755 1074
rect 1831 1070 1835 1074
rect 2007 1070 2011 1074
rect 2047 1058 2051 1062
rect 2295 1058 2299 1062
rect 2423 1058 2427 1062
rect 2495 1058 2499 1062
rect 2559 1058 2563 1062
rect 2599 1058 2603 1062
rect 2695 1058 2699 1062
rect 2711 1058 2715 1062
rect 2839 1058 2843 1062
rect 2847 1058 2851 1062
rect 2991 1058 2995 1062
rect 3007 1058 3011 1062
rect 3151 1058 3155 1062
rect 3199 1058 3203 1062
rect 3319 1058 3323 1062
rect 3407 1058 3411 1062
rect 3495 1058 3499 1062
rect 3631 1058 3635 1062
rect 3679 1058 3683 1062
rect 3839 1058 3843 1062
rect 3943 1058 3947 1062
rect 111 994 115 998
rect 135 994 139 998
rect 231 994 235 998
rect 271 994 275 998
rect 375 994 379 998
rect 447 994 451 998
rect 543 994 547 998
rect 631 994 635 998
rect 727 994 731 998
rect 823 994 827 998
rect 911 994 915 998
rect 1007 994 1011 998
rect 1095 994 1099 998
rect 1175 994 1179 998
rect 1279 994 1283 998
rect 1335 994 1339 998
rect 1463 994 1467 998
rect 1487 994 1491 998
rect 1631 994 1635 998
rect 1647 994 1651 998
rect 1775 994 1779 998
rect 1831 994 1835 998
rect 1903 994 1907 998
rect 2007 994 2011 998
rect 2047 982 2051 986
rect 2495 982 2499 986
rect 2599 982 2603 986
rect 2647 982 2651 986
rect 2711 982 2715 986
rect 2743 982 2747 986
rect 2847 982 2851 986
rect 2967 982 2971 986
rect 3007 982 3011 986
rect 3111 982 3115 986
rect 3199 982 3203 986
rect 3279 982 3283 986
rect 3407 982 3411 986
rect 3463 982 3467 986
rect 3631 982 3635 986
rect 3663 982 3667 986
rect 3839 982 3843 986
rect 3943 982 3947 986
rect 111 918 115 922
rect 135 918 139 922
rect 271 918 275 922
rect 447 918 451 922
rect 455 918 459 922
rect 631 918 635 922
rect 655 918 659 922
rect 823 918 827 922
rect 855 918 859 922
rect 1007 918 1011 922
rect 1055 918 1059 922
rect 1175 918 1179 922
rect 1239 918 1243 922
rect 1335 918 1339 922
rect 1415 918 1419 922
rect 1487 918 1491 922
rect 1583 918 1587 922
rect 1631 918 1635 922
rect 1751 918 1755 922
rect 1775 918 1779 922
rect 1903 918 1907 922
rect 2007 918 2011 922
rect 2047 894 2051 898
rect 2071 894 2075 898
rect 2255 894 2259 898
rect 2463 894 2467 898
rect 2647 894 2651 898
rect 2679 894 2683 898
rect 2743 894 2747 898
rect 2847 894 2851 898
rect 2895 894 2899 898
rect 2967 894 2971 898
rect 3111 894 3115 898
rect 3127 894 3131 898
rect 3279 894 3283 898
rect 3367 894 3371 898
rect 3463 894 3467 898
rect 3615 894 3619 898
rect 3663 894 3667 898
rect 3839 894 3843 898
rect 3943 894 3947 898
rect 111 842 115 846
rect 135 842 139 846
rect 215 842 219 846
rect 271 842 275 846
rect 343 842 347 846
rect 455 842 459 846
rect 495 842 499 846
rect 655 842 659 846
rect 831 842 835 846
rect 855 842 859 846
rect 1007 842 1011 846
rect 1055 842 1059 846
rect 1183 842 1187 846
rect 1239 842 1243 846
rect 1359 842 1363 846
rect 1415 842 1419 846
rect 1535 842 1539 846
rect 1583 842 1587 846
rect 1719 842 1723 846
rect 1751 842 1755 846
rect 1903 842 1907 846
rect 2007 842 2011 846
rect 2047 818 2051 822
rect 2071 818 2075 822
rect 2215 818 2219 822
rect 2255 818 2259 822
rect 2327 818 2331 822
rect 2447 818 2451 822
rect 2463 818 2467 822
rect 2583 818 2587 822
rect 2679 818 2683 822
rect 2735 818 2739 822
rect 2895 818 2899 822
rect 3063 818 3067 822
rect 3127 818 3131 822
rect 3247 818 3251 822
rect 3367 818 3371 822
rect 3447 818 3451 822
rect 3615 818 3619 822
rect 3655 818 3659 822
rect 3839 818 3843 822
rect 3943 818 3947 822
rect 111 766 115 770
rect 215 766 219 770
rect 343 766 347 770
rect 375 766 379 770
rect 495 766 499 770
rect 623 766 627 770
rect 655 766 659 770
rect 751 766 755 770
rect 831 766 835 770
rect 887 766 891 770
rect 1007 766 1011 770
rect 1023 766 1027 770
rect 1167 766 1171 770
rect 1183 766 1187 770
rect 1311 766 1315 770
rect 1359 766 1363 770
rect 1455 766 1459 770
rect 1535 766 1539 770
rect 1599 766 1603 770
rect 1719 766 1723 770
rect 2007 766 2011 770
rect 2047 738 2051 742
rect 2215 738 2219 742
rect 2327 738 2331 742
rect 2375 738 2379 742
rect 2447 738 2451 742
rect 2495 738 2499 742
rect 2583 738 2587 742
rect 2623 738 2627 742
rect 2735 738 2739 742
rect 2767 738 2771 742
rect 2895 738 2899 742
rect 2911 738 2915 742
rect 3063 738 3067 742
rect 3215 738 3219 742
rect 3247 738 3251 742
rect 3367 738 3371 742
rect 3447 738 3451 742
rect 3519 738 3523 742
rect 3655 738 3659 742
rect 3679 738 3683 742
rect 3839 738 3843 742
rect 3943 738 3947 742
rect 111 690 115 694
rect 375 690 379 694
rect 495 690 499 694
rect 527 690 531 694
rect 623 690 627 694
rect 631 690 635 694
rect 743 690 747 694
rect 751 690 755 694
rect 855 690 859 694
rect 887 690 891 694
rect 967 690 971 694
rect 1023 690 1027 694
rect 1071 690 1075 694
rect 1167 690 1171 694
rect 1183 690 1187 694
rect 1295 690 1299 694
rect 1311 690 1315 694
rect 1407 690 1411 694
rect 1455 690 1459 694
rect 1519 690 1523 694
rect 1599 690 1603 694
rect 2007 690 2011 694
rect 2047 654 2051 658
rect 2111 654 2115 658
rect 2247 654 2251 658
rect 2375 654 2379 658
rect 2399 654 2403 658
rect 2495 654 2499 658
rect 2575 654 2579 658
rect 2623 654 2627 658
rect 2759 654 2763 658
rect 2767 654 2771 658
rect 2911 654 2915 658
rect 2943 654 2947 658
rect 3063 654 3067 658
rect 3127 654 3131 658
rect 3215 654 3219 658
rect 3303 654 3307 658
rect 3367 654 3371 658
rect 3479 654 3483 658
rect 3519 654 3523 658
rect 3655 654 3659 658
rect 3679 654 3683 658
rect 3831 654 3835 658
rect 3839 654 3843 658
rect 3943 654 3947 658
rect 111 614 115 618
rect 527 614 531 618
rect 631 614 635 618
rect 687 614 691 618
rect 743 614 747 618
rect 783 614 787 618
rect 855 614 859 618
rect 879 614 883 618
rect 967 614 971 618
rect 975 614 979 618
rect 1071 614 1075 618
rect 1167 614 1171 618
rect 1183 614 1187 618
rect 1263 614 1267 618
rect 1295 614 1299 618
rect 1359 614 1363 618
rect 1407 614 1411 618
rect 1455 614 1459 618
rect 1519 614 1523 618
rect 2007 614 2011 618
rect 2047 574 2051 578
rect 2071 574 2075 578
rect 2111 574 2115 578
rect 2183 574 2187 578
rect 2247 574 2251 578
rect 2335 574 2339 578
rect 2399 574 2403 578
rect 2503 574 2507 578
rect 2575 574 2579 578
rect 2687 574 2691 578
rect 2759 574 2763 578
rect 2879 574 2883 578
rect 2943 574 2947 578
rect 3071 574 3075 578
rect 3127 574 3131 578
rect 3263 574 3267 578
rect 3303 574 3307 578
rect 3455 574 3459 578
rect 3479 574 3483 578
rect 3647 574 3651 578
rect 3655 574 3659 578
rect 3831 574 3835 578
rect 3839 574 3843 578
rect 3943 574 3947 578
rect 111 518 115 522
rect 383 518 387 522
rect 479 518 483 522
rect 575 518 579 522
rect 671 518 675 522
rect 687 518 691 522
rect 767 518 771 522
rect 783 518 787 522
rect 863 518 867 522
rect 879 518 883 522
rect 959 518 963 522
rect 975 518 979 522
rect 1055 518 1059 522
rect 1071 518 1075 522
rect 1151 518 1155 522
rect 1167 518 1171 522
rect 1247 518 1251 522
rect 1263 518 1267 522
rect 1343 518 1347 522
rect 1359 518 1363 522
rect 1439 518 1443 522
rect 1455 518 1459 522
rect 1535 518 1539 522
rect 2007 518 2011 522
rect 2047 498 2051 502
rect 2071 498 2075 502
rect 2183 498 2187 502
rect 2319 498 2323 502
rect 2335 498 2339 502
rect 2463 498 2467 502
rect 2503 498 2507 502
rect 2615 498 2619 502
rect 2687 498 2691 502
rect 2775 498 2779 502
rect 2879 498 2883 502
rect 2959 498 2963 502
rect 3071 498 3075 502
rect 3159 498 3163 502
rect 3263 498 3267 502
rect 3367 498 3371 502
rect 3455 498 3459 502
rect 3583 498 3587 502
rect 3647 498 3651 502
rect 3807 498 3811 502
rect 3839 498 3843 502
rect 3943 498 3947 502
rect 111 430 115 434
rect 383 430 387 434
rect 479 430 483 434
rect 487 430 491 434
rect 575 430 579 434
rect 583 430 587 434
rect 671 430 675 434
rect 687 430 691 434
rect 767 430 771 434
rect 791 430 795 434
rect 863 430 867 434
rect 895 430 899 434
rect 959 430 963 434
rect 999 430 1003 434
rect 1055 430 1059 434
rect 1103 430 1107 434
rect 1151 430 1155 434
rect 1207 430 1211 434
rect 1247 430 1251 434
rect 1319 430 1323 434
rect 1343 430 1347 434
rect 1431 430 1435 434
rect 1439 430 1443 434
rect 1535 430 1539 434
rect 2007 430 2011 434
rect 2047 422 2051 426
rect 2183 422 2187 426
rect 2319 422 2323 426
rect 2343 422 2347 426
rect 2463 422 2467 426
rect 2487 422 2491 426
rect 2615 422 2619 426
rect 2639 422 2643 426
rect 2775 422 2779 426
rect 2799 422 2803 426
rect 2959 422 2963 426
rect 3111 422 3115 426
rect 3159 422 3163 426
rect 3263 422 3267 426
rect 3367 422 3371 426
rect 3415 422 3419 426
rect 3559 422 3563 426
rect 3583 422 3587 426
rect 3711 422 3715 426
rect 3807 422 3811 426
rect 3839 422 3843 426
rect 3943 422 3947 426
rect 111 350 115 354
rect 327 350 331 354
rect 463 350 467 354
rect 487 350 491 354
rect 583 350 587 354
rect 615 350 619 354
rect 687 350 691 354
rect 767 350 771 354
rect 791 350 795 354
rect 895 350 899 354
rect 919 350 923 354
rect 999 350 1003 354
rect 1063 350 1067 354
rect 1103 350 1107 354
rect 1207 350 1211 354
rect 1319 350 1323 354
rect 1351 350 1355 354
rect 1431 350 1435 354
rect 1495 350 1499 354
rect 1639 350 1643 354
rect 2007 350 2011 354
rect 2047 342 2051 346
rect 2343 342 2347 346
rect 2487 342 2491 346
rect 2495 342 2499 346
rect 2639 342 2643 346
rect 2799 342 2803 346
rect 2959 342 2963 346
rect 3111 342 3115 346
rect 3119 342 3123 346
rect 3263 342 3267 346
rect 3271 342 3275 346
rect 3415 342 3419 346
rect 3423 342 3427 346
rect 3559 342 3563 346
rect 3567 342 3571 346
rect 3711 342 3715 346
rect 3839 342 3843 346
rect 3943 342 3947 346
rect 111 266 115 270
rect 167 266 171 270
rect 327 266 331 270
rect 463 266 467 270
rect 503 266 507 270
rect 615 266 619 270
rect 687 266 691 270
rect 767 266 771 270
rect 871 266 875 270
rect 919 266 923 270
rect 1047 266 1051 270
rect 1063 266 1067 270
rect 1207 266 1211 270
rect 1215 266 1219 270
rect 1351 266 1355 270
rect 1367 266 1371 270
rect 1495 266 1499 270
rect 1511 266 1515 270
rect 1639 266 1643 270
rect 1647 266 1651 270
rect 1783 266 1787 270
rect 1903 266 1907 270
rect 2007 266 2011 270
rect 2047 266 2051 270
rect 2071 266 2075 270
rect 2271 266 2275 270
rect 2495 266 2499 270
rect 2639 266 2643 270
rect 2703 266 2707 270
rect 2799 266 2803 270
rect 2903 266 2907 270
rect 2959 266 2963 270
rect 3095 266 3099 270
rect 3119 266 3123 270
rect 3271 266 3275 270
rect 3287 266 3291 270
rect 3423 266 3427 270
rect 3479 266 3483 270
rect 3567 266 3571 270
rect 3671 266 3675 270
rect 3711 266 3715 270
rect 3839 266 3843 270
rect 3943 266 3947 270
rect 111 162 115 166
rect 135 162 139 166
rect 167 162 171 166
rect 231 162 235 166
rect 327 162 331 166
rect 423 162 427 166
rect 503 162 507 166
rect 527 162 531 166
rect 647 162 651 166
rect 687 162 691 166
rect 775 162 779 166
rect 871 162 875 166
rect 903 162 907 166
rect 1031 162 1035 166
rect 1047 162 1051 166
rect 1151 162 1155 166
rect 1215 162 1219 166
rect 1271 162 1275 166
rect 1367 162 1371 166
rect 1383 162 1387 166
rect 1487 162 1491 166
rect 1511 162 1515 166
rect 1591 162 1595 166
rect 1647 162 1651 166
rect 1703 162 1707 166
rect 1783 162 1787 166
rect 1807 162 1811 166
rect 1903 162 1907 166
rect 2007 162 2011 166
rect 2047 166 2051 170
rect 2071 166 2075 170
rect 2167 166 2171 170
rect 2263 166 2267 170
rect 2271 166 2275 170
rect 2359 166 2363 170
rect 2455 166 2459 170
rect 2495 166 2499 170
rect 2551 166 2555 170
rect 2655 166 2659 170
rect 2703 166 2707 170
rect 2759 166 2763 170
rect 2863 166 2867 170
rect 2903 166 2907 170
rect 2975 166 2979 170
rect 3095 166 3099 170
rect 3103 166 3107 170
rect 3239 166 3243 170
rect 3287 166 3291 170
rect 3383 166 3387 170
rect 3479 166 3483 170
rect 3535 166 3539 170
rect 3671 166 3675 170
rect 3695 166 3699 170
rect 3839 166 3843 170
rect 3943 166 3947 170
rect 111 86 115 90
rect 135 86 139 90
rect 231 86 235 90
rect 327 86 331 90
rect 423 86 427 90
rect 527 86 531 90
rect 647 86 651 90
rect 775 86 779 90
rect 903 86 907 90
rect 1031 86 1035 90
rect 1151 86 1155 90
rect 1271 86 1275 90
rect 1383 86 1387 90
rect 1487 86 1491 90
rect 1591 86 1595 90
rect 1703 86 1707 90
rect 1807 86 1811 90
rect 1903 86 1907 90
rect 2007 86 2011 90
rect 2047 90 2051 94
rect 2071 90 2075 94
rect 2167 90 2171 94
rect 2263 90 2267 94
rect 2359 90 2363 94
rect 2455 90 2459 94
rect 2551 90 2555 94
rect 2655 90 2659 94
rect 2759 90 2763 94
rect 2863 90 2867 94
rect 2975 90 2979 94
rect 3103 90 3107 94
rect 3239 90 3243 94
rect 3383 90 3387 94
rect 3535 90 3539 94
rect 3695 90 3699 94
rect 3839 90 3843 94
rect 3943 90 3947 94
<< m4 >>
rect 96 4025 97 4031
rect 103 4030 2031 4031
rect 103 4026 111 4030
rect 115 4026 1519 4030
rect 1523 4026 1615 4030
rect 1619 4026 1711 4030
rect 1715 4026 1807 4030
rect 1811 4026 1903 4030
rect 1907 4026 2007 4030
rect 2011 4026 2031 4030
rect 103 4025 2031 4026
rect 2037 4025 2038 4031
rect 2018 4013 2019 4019
rect 2025 4018 3967 4019
rect 2025 4014 2047 4018
rect 2051 4014 2071 4018
rect 2075 4014 2167 4018
rect 2171 4014 2263 4018
rect 2267 4014 3943 4018
rect 3947 4014 3967 4018
rect 2025 4013 3967 4014
rect 3973 4013 3974 4019
rect 84 3949 85 3955
rect 91 3954 2019 3955
rect 91 3950 111 3954
rect 115 3950 199 3954
rect 203 3950 295 3954
rect 299 3950 391 3954
rect 395 3950 495 3954
rect 499 3950 615 3954
rect 619 3950 743 3954
rect 747 3950 871 3954
rect 875 3950 999 3954
rect 1003 3950 1127 3954
rect 1131 3950 1255 3954
rect 1259 3950 1383 3954
rect 1387 3950 1511 3954
rect 1515 3950 1519 3954
rect 1523 3950 1615 3954
rect 1619 3950 1647 3954
rect 1651 3950 1711 3954
rect 1715 3950 1807 3954
rect 1811 3950 1903 3954
rect 1907 3950 2007 3954
rect 2011 3950 2019 3954
rect 91 3949 2019 3950
rect 2025 3949 2026 3955
rect 2030 3937 2031 3943
rect 2037 3942 3979 3943
rect 2037 3938 2047 3942
rect 2051 3938 2071 3942
rect 2075 3938 2159 3942
rect 2163 3938 2167 3942
rect 2171 3938 2263 3942
rect 2267 3938 2287 3942
rect 2291 3938 2415 3942
rect 2419 3938 2551 3942
rect 2555 3938 2687 3942
rect 2691 3938 2823 3942
rect 2827 3938 2951 3942
rect 2955 3938 3071 3942
rect 3075 3938 3191 3942
rect 3195 3938 3303 3942
rect 3307 3938 3407 3942
rect 3411 3938 3519 3942
rect 3523 3938 3631 3942
rect 3635 3938 3743 3942
rect 3747 3938 3943 3942
rect 3947 3938 3979 3942
rect 2037 3937 3979 3938
rect 3985 3937 3986 3943
rect 96 3873 97 3879
rect 103 3878 2031 3879
rect 103 3874 111 3878
rect 115 3874 199 3878
rect 203 3874 295 3878
rect 299 3874 335 3878
rect 339 3874 391 3878
rect 395 3874 455 3878
rect 459 3874 495 3878
rect 499 3874 583 3878
rect 587 3874 615 3878
rect 619 3874 719 3878
rect 723 3874 743 3878
rect 747 3874 847 3878
rect 851 3874 871 3878
rect 875 3874 975 3878
rect 979 3874 999 3878
rect 1003 3874 1103 3878
rect 1107 3874 1127 3878
rect 1131 3874 1231 3878
rect 1235 3874 1255 3878
rect 1259 3874 1359 3878
rect 1363 3874 1383 3878
rect 1387 3874 1487 3878
rect 1491 3874 1511 3878
rect 1515 3874 1647 3878
rect 1651 3874 2007 3878
rect 2011 3874 2031 3878
rect 103 3873 2031 3874
rect 2037 3873 2038 3879
rect 2018 3853 2019 3859
rect 2025 3858 3967 3859
rect 2025 3854 2047 3858
rect 2051 3854 2159 3858
rect 2163 3854 2207 3858
rect 2211 3854 2287 3858
rect 2291 3854 2343 3858
rect 2347 3854 2415 3858
rect 2419 3854 2487 3858
rect 2491 3854 2551 3858
rect 2555 3854 2647 3858
rect 2651 3854 2687 3858
rect 2691 3854 2823 3858
rect 2827 3854 2951 3858
rect 2955 3854 3015 3858
rect 3019 3854 3071 3858
rect 3075 3854 3191 3858
rect 3195 3854 3223 3858
rect 3227 3854 3303 3858
rect 3307 3854 3407 3858
rect 3411 3854 3439 3858
rect 3443 3854 3519 3858
rect 3523 3854 3631 3858
rect 3635 3854 3655 3858
rect 3659 3854 3743 3858
rect 3747 3854 3943 3858
rect 3947 3854 3967 3858
rect 2025 3853 3967 3854
rect 3973 3853 3974 3859
rect 84 3793 85 3799
rect 91 3798 2019 3799
rect 91 3794 111 3798
rect 115 3794 335 3798
rect 339 3794 455 3798
rect 459 3794 503 3798
rect 507 3794 583 3798
rect 587 3794 615 3798
rect 619 3794 719 3798
rect 723 3794 735 3798
rect 739 3794 847 3798
rect 851 3794 863 3798
rect 867 3794 975 3798
rect 979 3794 999 3798
rect 1003 3794 1103 3798
rect 1107 3794 1143 3798
rect 1147 3794 1231 3798
rect 1235 3794 1287 3798
rect 1291 3794 1359 3798
rect 1363 3794 1431 3798
rect 1435 3794 1487 3798
rect 1491 3794 1583 3798
rect 1587 3794 2007 3798
rect 2011 3794 2019 3798
rect 91 3793 2019 3794
rect 2025 3793 2026 3799
rect 2030 3777 2031 3783
rect 2037 3782 3979 3783
rect 2037 3778 2047 3782
rect 2051 3778 2191 3782
rect 2195 3778 2207 3782
rect 2211 3778 2343 3782
rect 2347 3778 2375 3782
rect 2379 3778 2487 3782
rect 2491 3778 2559 3782
rect 2563 3778 2647 3782
rect 2651 3778 2743 3782
rect 2747 3778 2823 3782
rect 2827 3778 2935 3782
rect 2939 3778 3015 3782
rect 3019 3778 3127 3782
rect 3131 3778 3223 3782
rect 3227 3778 3319 3782
rect 3323 3778 3439 3782
rect 3443 3778 3511 3782
rect 3515 3778 3655 3782
rect 3659 3778 3711 3782
rect 3715 3778 3943 3782
rect 3947 3778 3979 3782
rect 2037 3777 3979 3778
rect 3985 3777 3986 3783
rect 96 3709 97 3715
rect 103 3714 2031 3715
rect 103 3710 111 3714
rect 115 3710 495 3714
rect 499 3710 503 3714
rect 507 3710 591 3714
rect 595 3710 615 3714
rect 619 3710 687 3714
rect 691 3710 735 3714
rect 739 3710 791 3714
rect 795 3710 863 3714
rect 867 3710 911 3714
rect 915 3710 999 3714
rect 1003 3710 1039 3714
rect 1043 3710 1143 3714
rect 1147 3710 1183 3714
rect 1187 3710 1287 3714
rect 1291 3710 1335 3714
rect 1339 3710 1431 3714
rect 1435 3710 1495 3714
rect 1499 3710 1583 3714
rect 1587 3710 1655 3714
rect 1659 3710 2007 3714
rect 2011 3710 2031 3714
rect 103 3709 2031 3710
rect 2037 3709 2038 3715
rect 2018 3697 2019 3703
rect 2025 3702 3967 3703
rect 2025 3698 2047 3702
rect 2051 3698 2127 3702
rect 2131 3698 2191 3702
rect 2195 3698 2351 3702
rect 2355 3698 2375 3702
rect 2379 3698 2559 3702
rect 2563 3698 2583 3702
rect 2587 3698 2743 3702
rect 2747 3698 2815 3702
rect 2819 3698 2935 3702
rect 2939 3698 3047 3702
rect 3051 3698 3127 3702
rect 3131 3698 3279 3702
rect 3283 3698 3319 3702
rect 3323 3698 3511 3702
rect 3515 3698 3711 3702
rect 3715 3698 3751 3702
rect 3755 3698 3943 3702
rect 3947 3698 3967 3702
rect 2025 3697 3967 3698
rect 3973 3697 3974 3703
rect 84 3625 85 3631
rect 91 3630 2019 3631
rect 91 3626 111 3630
rect 115 3626 335 3630
rect 339 3626 463 3630
rect 467 3626 495 3630
rect 499 3626 591 3630
rect 595 3626 607 3630
rect 611 3626 687 3630
rect 691 3626 759 3630
rect 763 3626 791 3630
rect 795 3626 911 3630
rect 915 3626 927 3630
rect 931 3626 1039 3630
rect 1043 3626 1095 3630
rect 1099 3626 1183 3630
rect 1187 3626 1263 3630
rect 1267 3626 1335 3630
rect 1339 3626 1439 3630
rect 1443 3626 1495 3630
rect 1499 3626 1615 3630
rect 1619 3626 1655 3630
rect 1659 3626 1791 3630
rect 1795 3626 2007 3630
rect 2011 3626 2019 3630
rect 91 3625 2019 3626
rect 2025 3625 2026 3631
rect 2030 3613 2031 3619
rect 2037 3618 3979 3619
rect 2037 3614 2047 3618
rect 2051 3614 2127 3618
rect 2131 3614 2191 3618
rect 2195 3614 2327 3618
rect 2331 3614 2351 3618
rect 2355 3614 2455 3618
rect 2459 3614 2583 3618
rect 2587 3614 2719 3618
rect 2723 3614 2815 3618
rect 2819 3614 2855 3618
rect 2859 3614 2999 3618
rect 3003 3614 3047 3618
rect 3051 3614 3143 3618
rect 3147 3614 3279 3618
rect 3283 3614 3295 3618
rect 3299 3614 3455 3618
rect 3459 3614 3511 3618
rect 3515 3614 3623 3618
rect 3627 3614 3751 3618
rect 3755 3614 3943 3618
rect 3947 3614 3979 3618
rect 2037 3613 3979 3614
rect 3985 3613 3986 3619
rect 2018 3547 2019 3553
rect 2025 3547 2050 3553
rect 2044 3543 2050 3547
rect 96 3537 97 3543
rect 103 3542 2031 3543
rect 103 3538 111 3542
rect 115 3538 159 3542
rect 163 3538 303 3542
rect 307 3538 335 3542
rect 339 3538 463 3542
rect 467 3538 607 3542
rect 611 3538 639 3542
rect 643 3538 759 3542
rect 763 3538 815 3542
rect 819 3538 927 3542
rect 931 3538 999 3542
rect 1003 3538 1095 3542
rect 1099 3538 1175 3542
rect 1179 3538 1263 3542
rect 1267 3538 1351 3542
rect 1355 3538 1439 3542
rect 1443 3538 1527 3542
rect 1531 3538 1615 3542
rect 1619 3538 1703 3542
rect 1707 3538 1791 3542
rect 1795 3538 1879 3542
rect 1883 3538 2007 3542
rect 2011 3538 2031 3542
rect 103 3537 2031 3538
rect 2037 3537 2038 3543
rect 2044 3542 3967 3543
rect 2044 3538 2047 3542
rect 2051 3538 2103 3542
rect 2107 3538 2191 3542
rect 2195 3538 2271 3542
rect 2275 3538 2327 3542
rect 2331 3538 2447 3542
rect 2451 3538 2455 3542
rect 2459 3538 2583 3542
rect 2587 3538 2631 3542
rect 2635 3538 2719 3542
rect 2723 3538 2815 3542
rect 2819 3538 2855 3542
rect 2859 3538 2999 3542
rect 3003 3538 3143 3542
rect 3147 3538 3175 3542
rect 3179 3538 3295 3542
rect 3299 3538 3351 3542
rect 3355 3538 3455 3542
rect 3459 3538 3519 3542
rect 3523 3538 3623 3542
rect 3627 3538 3687 3542
rect 3691 3538 3839 3542
rect 3843 3538 3943 3542
rect 3947 3538 3967 3542
rect 2044 3537 3967 3538
rect 3973 3537 3974 3543
rect 84 3453 85 3459
rect 91 3458 2019 3459
rect 91 3454 111 3458
rect 115 3454 135 3458
rect 139 3454 159 3458
rect 163 3454 303 3458
rect 307 3454 319 3458
rect 323 3454 463 3458
rect 467 3454 535 3458
rect 539 3454 639 3458
rect 643 3454 751 3458
rect 755 3454 815 3458
rect 819 3454 959 3458
rect 963 3454 999 3458
rect 1003 3454 1159 3458
rect 1163 3454 1175 3458
rect 1179 3454 1351 3458
rect 1355 3454 1527 3458
rect 1531 3454 1535 3458
rect 1539 3454 1703 3458
rect 1707 3454 1719 3458
rect 1723 3454 1879 3458
rect 1883 3454 1903 3458
rect 1907 3454 2007 3458
rect 2011 3454 2019 3458
rect 91 3453 2019 3454
rect 2025 3453 2026 3459
rect 2030 3457 2031 3463
rect 2037 3462 3979 3463
rect 2037 3458 2047 3462
rect 2051 3458 2103 3462
rect 2107 3458 2127 3462
rect 2131 3458 2271 3462
rect 2275 3458 2311 3462
rect 2315 3458 2447 3462
rect 2451 3458 2495 3462
rect 2499 3458 2631 3462
rect 2635 3458 2679 3462
rect 2683 3458 2815 3462
rect 2819 3458 2863 3462
rect 2867 3458 2999 3462
rect 3003 3458 3047 3462
rect 3051 3458 3175 3462
rect 3179 3458 3223 3462
rect 3227 3458 3351 3462
rect 3355 3458 3407 3462
rect 3411 3458 3519 3462
rect 3523 3458 3591 3462
rect 3595 3458 3687 3462
rect 3691 3458 3775 3462
rect 3779 3458 3839 3462
rect 3843 3458 3943 3462
rect 3947 3458 3979 3462
rect 2037 3457 3979 3458
rect 3985 3457 3986 3463
rect 96 3377 97 3383
rect 103 3382 2031 3383
rect 103 3378 111 3382
rect 115 3378 135 3382
rect 139 3378 231 3382
rect 235 3378 319 3382
rect 323 3378 375 3382
rect 379 3378 535 3382
rect 539 3378 703 3382
rect 707 3378 751 3382
rect 755 3378 871 3382
rect 875 3378 959 3382
rect 963 3378 1047 3382
rect 1051 3378 1159 3382
rect 1163 3378 1215 3382
rect 1219 3378 1351 3382
rect 1355 3378 1383 3382
rect 1387 3378 1535 3382
rect 1539 3378 1543 3382
rect 1547 3378 1703 3382
rect 1707 3378 1719 3382
rect 1723 3378 1871 3382
rect 1875 3378 1903 3382
rect 1907 3378 2007 3382
rect 2011 3378 2031 3382
rect 103 3377 2031 3378
rect 2037 3377 2038 3383
rect 2018 3365 2019 3371
rect 2025 3370 3967 3371
rect 2025 3366 2047 3370
rect 2051 3366 2071 3370
rect 2075 3366 2127 3370
rect 2131 3366 2215 3370
rect 2219 3366 2311 3370
rect 2315 3366 2359 3370
rect 2363 3366 2495 3370
rect 2499 3366 2511 3370
rect 2515 3366 2655 3370
rect 2659 3366 2679 3370
rect 2683 3366 2799 3370
rect 2803 3366 2863 3370
rect 2867 3366 2935 3370
rect 2939 3366 3047 3370
rect 3051 3366 3079 3370
rect 3083 3366 3223 3370
rect 3227 3366 3375 3370
rect 3379 3366 3407 3370
rect 3411 3366 3535 3370
rect 3539 3366 3591 3370
rect 3595 3366 3695 3370
rect 3699 3366 3775 3370
rect 3779 3366 3839 3370
rect 3843 3366 3943 3370
rect 3947 3366 3967 3370
rect 2025 3365 3967 3366
rect 3973 3365 3974 3371
rect 84 3301 85 3307
rect 91 3306 2019 3307
rect 91 3302 111 3306
rect 115 3302 135 3306
rect 139 3302 231 3306
rect 235 3302 279 3306
rect 283 3302 375 3306
rect 379 3302 463 3306
rect 467 3302 535 3306
rect 539 3302 663 3306
rect 667 3302 703 3306
rect 707 3302 871 3306
rect 875 3302 1047 3306
rect 1051 3302 1079 3306
rect 1083 3302 1215 3306
rect 1219 3302 1295 3306
rect 1299 3302 1383 3306
rect 1387 3302 1519 3306
rect 1523 3302 1543 3306
rect 1547 3302 1703 3306
rect 1707 3302 1743 3306
rect 1747 3302 1871 3306
rect 1875 3302 2007 3306
rect 2011 3302 2019 3306
rect 91 3301 2019 3302
rect 2025 3301 2026 3307
rect 2030 3281 2031 3287
rect 2037 3286 3979 3287
rect 2037 3282 2047 3286
rect 2051 3282 2071 3286
rect 2075 3282 2111 3286
rect 2115 3282 2215 3286
rect 2219 3282 2247 3286
rect 2251 3282 2359 3286
rect 2363 3282 2399 3286
rect 2403 3282 2511 3286
rect 2515 3282 2575 3286
rect 2579 3282 2655 3286
rect 2659 3282 2783 3286
rect 2787 3282 2799 3286
rect 2803 3282 2935 3286
rect 2939 3282 3015 3286
rect 3019 3282 3079 3286
rect 3083 3282 3223 3286
rect 3227 3282 3263 3286
rect 3267 3282 3375 3286
rect 3379 3282 3527 3286
rect 3531 3282 3535 3286
rect 3539 3282 3695 3286
rect 3699 3282 3791 3286
rect 3795 3282 3839 3286
rect 3843 3282 3943 3286
rect 3947 3282 3979 3286
rect 2037 3281 3979 3282
rect 3985 3281 3986 3287
rect 96 3225 97 3231
rect 103 3230 2031 3231
rect 103 3226 111 3230
rect 115 3226 135 3230
rect 139 3226 279 3230
rect 283 3226 287 3230
rect 291 3226 447 3230
rect 451 3226 463 3230
rect 467 3226 615 3230
rect 619 3226 663 3230
rect 667 3226 791 3230
rect 795 3226 871 3230
rect 875 3226 967 3230
rect 971 3226 1079 3230
rect 1083 3226 1143 3230
rect 1147 3226 1295 3230
rect 1299 3226 1327 3230
rect 1331 3226 1511 3230
rect 1515 3226 1519 3230
rect 1523 3226 1695 3230
rect 1699 3226 1743 3230
rect 1747 3226 2007 3230
rect 2011 3226 2031 3230
rect 103 3225 2031 3226
rect 2037 3225 2038 3231
rect 2018 3205 2019 3211
rect 2025 3210 3967 3211
rect 2025 3206 2047 3210
rect 2051 3206 2071 3210
rect 2075 3206 2111 3210
rect 2115 3206 2167 3210
rect 2171 3206 2247 3210
rect 2251 3206 2263 3210
rect 2267 3206 2359 3210
rect 2363 3206 2399 3210
rect 2403 3206 2455 3210
rect 2459 3206 2551 3210
rect 2555 3206 2575 3210
rect 2579 3206 2647 3210
rect 2651 3206 2743 3210
rect 2747 3206 2783 3210
rect 2787 3206 2839 3210
rect 2843 3206 2935 3210
rect 2939 3206 3015 3210
rect 3019 3206 3031 3210
rect 3035 3206 3127 3210
rect 3131 3206 3223 3210
rect 3227 3206 3263 3210
rect 3267 3206 3319 3210
rect 3323 3206 3439 3210
rect 3443 3206 3527 3210
rect 3531 3206 3575 3210
rect 3579 3206 3719 3210
rect 3723 3206 3791 3210
rect 3795 3206 3839 3210
rect 3843 3206 3943 3210
rect 3947 3206 3967 3210
rect 2025 3205 3967 3206
rect 3973 3205 3974 3211
rect 84 3145 85 3151
rect 91 3150 2019 3151
rect 91 3146 111 3150
rect 115 3146 135 3150
rect 139 3146 287 3150
rect 291 3146 311 3150
rect 315 3146 439 3150
rect 443 3146 447 3150
rect 451 3146 583 3150
rect 587 3146 615 3150
rect 619 3146 743 3150
rect 747 3146 791 3150
rect 795 3146 903 3150
rect 907 3146 967 3150
rect 971 3146 1063 3150
rect 1067 3146 1143 3150
rect 1147 3146 1223 3150
rect 1227 3146 1327 3150
rect 1331 3146 1391 3150
rect 1395 3146 1511 3150
rect 1515 3146 1559 3150
rect 1563 3146 1695 3150
rect 1699 3146 1727 3150
rect 1731 3146 2007 3150
rect 2011 3146 2019 3150
rect 91 3145 2019 3146
rect 2025 3145 2026 3151
rect 2030 3117 2031 3123
rect 2037 3122 3979 3123
rect 2037 3118 2047 3122
rect 2051 3118 2071 3122
rect 2075 3118 2167 3122
rect 2171 3118 2263 3122
rect 2267 3118 2335 3122
rect 2339 3118 2359 3122
rect 2363 3118 2455 3122
rect 2459 3118 2551 3122
rect 2555 3118 2623 3122
rect 2627 3118 2647 3122
rect 2651 3118 2743 3122
rect 2747 3118 2839 3122
rect 2843 3118 2911 3122
rect 2915 3118 2935 3122
rect 2939 3118 3031 3122
rect 3035 3118 3127 3122
rect 3131 3118 3207 3122
rect 3211 3118 3223 3122
rect 3227 3118 3319 3122
rect 3323 3118 3439 3122
rect 3443 3118 3503 3122
rect 3507 3118 3575 3122
rect 3579 3118 3719 3122
rect 3723 3118 3799 3122
rect 3803 3118 3839 3122
rect 3843 3118 3943 3122
rect 3947 3118 3979 3122
rect 2037 3117 3979 3118
rect 3985 3117 3986 3123
rect 96 3061 97 3067
rect 103 3066 2031 3067
rect 103 3062 111 3066
rect 115 3062 311 3066
rect 315 3062 439 3066
rect 443 3062 503 3066
rect 507 3062 583 3066
rect 587 3062 599 3066
rect 603 3062 703 3066
rect 707 3062 743 3066
rect 747 3062 815 3066
rect 819 3062 903 3066
rect 907 3062 935 3066
rect 939 3062 1063 3066
rect 1067 3062 1071 3066
rect 1075 3062 1223 3066
rect 1227 3062 1383 3066
rect 1387 3062 1391 3066
rect 1395 3062 1551 3066
rect 1555 3062 1559 3066
rect 1563 3062 1719 3066
rect 1723 3062 1727 3066
rect 1731 3062 2007 3066
rect 2011 3062 2031 3066
rect 103 3061 2031 3062
rect 2037 3061 2038 3067
rect 2018 3041 2019 3047
rect 2025 3046 3967 3047
rect 2025 3042 2047 3046
rect 2051 3042 2071 3046
rect 2075 3042 2335 3046
rect 2339 3042 2383 3046
rect 2387 3042 2623 3046
rect 2627 3042 2703 3046
rect 2707 3042 2911 3046
rect 2915 3042 2999 3046
rect 3003 3042 3207 3046
rect 3211 3042 3287 3046
rect 3291 3042 3503 3046
rect 3507 3042 3575 3046
rect 3579 3042 3799 3046
rect 3803 3042 3839 3046
rect 3843 3042 3943 3046
rect 3947 3042 3967 3046
rect 2025 3041 3967 3042
rect 3973 3041 3974 3047
rect 84 2981 85 2987
rect 91 2986 2019 2987
rect 91 2982 111 2986
rect 115 2982 503 2986
rect 507 2982 551 2986
rect 555 2982 599 2986
rect 603 2982 647 2986
rect 651 2982 703 2986
rect 707 2982 759 2986
rect 763 2982 815 2986
rect 819 2982 887 2986
rect 891 2982 935 2986
rect 939 2982 1023 2986
rect 1027 2982 1071 2986
rect 1075 2982 1175 2986
rect 1179 2982 1223 2986
rect 1227 2982 1327 2986
rect 1331 2982 1383 2986
rect 1387 2982 1487 2986
rect 1491 2982 1551 2986
rect 1555 2982 1655 2986
rect 1659 2982 1719 2986
rect 1723 2982 1823 2986
rect 1827 2982 2007 2986
rect 2011 2982 2019 2986
rect 91 2981 2019 2982
rect 2025 2981 2026 2987
rect 2030 2961 2031 2967
rect 2037 2966 3979 2967
rect 2037 2962 2047 2966
rect 2051 2962 2071 2966
rect 2075 2962 2383 2966
rect 2387 2962 2391 2966
rect 2395 2962 2703 2966
rect 2707 2962 2975 2966
rect 2979 2962 2999 2966
rect 3003 2962 3215 2966
rect 3219 2962 3287 2966
rect 3291 2962 3439 2966
rect 3443 2962 3575 2966
rect 3579 2962 3647 2966
rect 3651 2962 3839 2966
rect 3843 2962 3943 2966
rect 3947 2962 3979 2966
rect 2037 2961 3979 2962
rect 3985 2961 3986 2967
rect 96 2897 97 2903
rect 103 2902 2031 2903
rect 103 2898 111 2902
rect 115 2898 471 2902
rect 475 2898 551 2902
rect 555 2898 575 2902
rect 579 2898 647 2902
rect 651 2898 695 2902
rect 699 2898 759 2902
rect 763 2898 839 2902
rect 843 2898 887 2902
rect 891 2898 991 2902
rect 995 2898 1023 2902
rect 1027 2898 1151 2902
rect 1155 2898 1175 2902
rect 1179 2898 1319 2902
rect 1323 2898 1327 2902
rect 1331 2898 1487 2902
rect 1491 2898 1495 2902
rect 1499 2898 1655 2902
rect 1659 2898 1671 2902
rect 1675 2898 1823 2902
rect 1827 2898 1847 2902
rect 1851 2898 2007 2902
rect 2011 2898 2031 2902
rect 103 2897 2031 2898
rect 2037 2897 2038 2903
rect 2018 2885 2019 2891
rect 2025 2890 3967 2891
rect 2025 2886 2047 2890
rect 2051 2886 2071 2890
rect 2075 2886 2295 2890
rect 2299 2886 2391 2890
rect 2395 2886 2535 2890
rect 2539 2886 2703 2890
rect 2707 2886 2767 2890
rect 2771 2886 2975 2890
rect 2979 2886 2991 2890
rect 2995 2886 3215 2890
rect 3219 2886 3431 2890
rect 3435 2886 3439 2890
rect 3443 2886 3647 2890
rect 3651 2886 3839 2890
rect 3843 2886 3943 2890
rect 3947 2886 3967 2890
rect 2025 2885 3967 2886
rect 3973 2885 3974 2891
rect 84 2817 85 2823
rect 91 2822 2019 2823
rect 91 2818 111 2822
rect 115 2818 471 2822
rect 475 2818 479 2822
rect 483 2818 575 2822
rect 579 2818 679 2822
rect 683 2818 695 2822
rect 699 2818 799 2822
rect 803 2818 839 2822
rect 843 2818 935 2822
rect 939 2818 991 2822
rect 995 2818 1079 2822
rect 1083 2818 1151 2822
rect 1155 2818 1239 2822
rect 1243 2818 1319 2822
rect 1323 2818 1415 2822
rect 1419 2818 1495 2822
rect 1499 2818 1599 2822
rect 1603 2818 1671 2822
rect 1675 2818 1783 2822
rect 1787 2818 1847 2822
rect 1851 2818 2007 2822
rect 2011 2818 2019 2822
rect 91 2817 2019 2818
rect 2025 2817 2026 2823
rect 2030 2805 2031 2811
rect 2037 2810 3979 2811
rect 2037 2806 2047 2810
rect 2051 2806 2071 2810
rect 2075 2806 2199 2810
rect 2203 2806 2295 2810
rect 2299 2806 2367 2810
rect 2371 2806 2535 2810
rect 2539 2806 2551 2810
rect 2555 2806 2735 2810
rect 2739 2806 2767 2810
rect 2771 2806 2927 2810
rect 2931 2806 2991 2810
rect 2995 2806 3111 2810
rect 3115 2806 3215 2810
rect 3219 2806 3295 2810
rect 3299 2806 3431 2810
rect 3435 2806 3479 2810
rect 3483 2806 3647 2810
rect 3651 2806 3671 2810
rect 3675 2806 3839 2810
rect 3843 2806 3943 2810
rect 3947 2806 3979 2810
rect 2037 2805 3979 2806
rect 3985 2805 3986 2811
rect 96 2737 97 2743
rect 103 2742 2031 2743
rect 103 2738 111 2742
rect 115 2738 479 2742
rect 483 2738 511 2742
rect 515 2738 575 2742
rect 579 2738 623 2742
rect 627 2738 679 2742
rect 683 2738 743 2742
rect 747 2738 799 2742
rect 803 2738 879 2742
rect 883 2738 935 2742
rect 939 2738 1015 2742
rect 1019 2738 1079 2742
rect 1083 2738 1159 2742
rect 1163 2738 1239 2742
rect 1243 2738 1311 2742
rect 1315 2738 1415 2742
rect 1419 2738 1463 2742
rect 1467 2738 1599 2742
rect 1603 2738 1623 2742
rect 1627 2738 1783 2742
rect 1787 2738 2007 2742
rect 2011 2738 2031 2742
rect 103 2737 2031 2738
rect 2037 2737 2038 2743
rect 2018 2725 2019 2731
rect 2025 2730 3967 2731
rect 2025 2726 2047 2730
rect 2051 2726 2071 2730
rect 2075 2726 2191 2730
rect 2195 2726 2199 2730
rect 2203 2726 2319 2730
rect 2323 2726 2367 2730
rect 2371 2726 2447 2730
rect 2451 2726 2551 2730
rect 2555 2726 2583 2730
rect 2587 2726 2727 2730
rect 2731 2726 2735 2730
rect 2739 2726 2887 2730
rect 2891 2726 2927 2730
rect 2931 2726 3063 2730
rect 3067 2726 3111 2730
rect 3115 2726 3255 2730
rect 3259 2726 3295 2730
rect 3299 2726 3455 2730
rect 3459 2726 3479 2730
rect 3483 2726 3655 2730
rect 3659 2726 3671 2730
rect 3675 2726 3839 2730
rect 3843 2726 3943 2730
rect 3947 2726 3967 2730
rect 2025 2725 3967 2726
rect 3973 2725 3974 2731
rect 84 2657 85 2663
rect 91 2662 2019 2663
rect 91 2658 111 2662
rect 115 2658 367 2662
rect 371 2658 487 2662
rect 491 2658 511 2662
rect 515 2658 615 2662
rect 619 2658 623 2662
rect 627 2658 743 2662
rect 747 2658 751 2662
rect 755 2658 879 2662
rect 883 2658 895 2662
rect 899 2658 1015 2662
rect 1019 2658 1031 2662
rect 1035 2658 1159 2662
rect 1163 2658 1167 2662
rect 1171 2658 1303 2662
rect 1307 2658 1311 2662
rect 1315 2658 1431 2662
rect 1435 2658 1463 2662
rect 1467 2658 1567 2662
rect 1571 2658 1623 2662
rect 1627 2658 1703 2662
rect 1707 2658 1783 2662
rect 1787 2658 2007 2662
rect 2011 2658 2019 2662
rect 91 2657 2019 2658
rect 2025 2657 2026 2663
rect 2030 2641 2031 2647
rect 2037 2646 3979 2647
rect 2037 2642 2047 2646
rect 2051 2642 2071 2646
rect 2075 2642 2191 2646
rect 2195 2642 2231 2646
rect 2235 2642 2319 2646
rect 2323 2642 2335 2646
rect 2339 2642 2447 2646
rect 2451 2642 2559 2646
rect 2563 2642 2583 2646
rect 2587 2642 2671 2646
rect 2675 2642 2727 2646
rect 2731 2642 2791 2646
rect 2795 2642 2887 2646
rect 2891 2642 2911 2646
rect 2915 2642 3031 2646
rect 3035 2642 3063 2646
rect 3067 2642 3151 2646
rect 3155 2642 3255 2646
rect 3259 2642 3455 2646
rect 3459 2642 3655 2646
rect 3659 2642 3839 2646
rect 3843 2642 3943 2646
rect 3947 2642 3979 2646
rect 2037 2641 3979 2642
rect 3985 2641 3986 2647
rect 96 2581 97 2587
rect 103 2586 2031 2587
rect 103 2582 111 2586
rect 115 2582 135 2586
rect 139 2582 287 2586
rect 291 2582 367 2586
rect 371 2582 447 2586
rect 451 2582 487 2586
rect 491 2582 607 2586
rect 611 2582 615 2586
rect 619 2582 751 2586
rect 755 2582 767 2586
rect 771 2582 895 2586
rect 899 2582 919 2586
rect 923 2582 1031 2586
rect 1035 2582 1063 2586
rect 1067 2582 1167 2586
rect 1171 2582 1199 2586
rect 1203 2582 1303 2586
rect 1307 2582 1335 2586
rect 1339 2582 1431 2586
rect 1435 2582 1463 2586
rect 1467 2582 1567 2586
rect 1571 2582 1591 2586
rect 1595 2582 1703 2586
rect 1707 2582 1727 2586
rect 1731 2582 2007 2586
rect 2011 2582 2031 2586
rect 103 2581 2031 2582
rect 2037 2581 2038 2587
rect 2018 2561 2019 2567
rect 2025 2566 3967 2567
rect 2025 2562 2047 2566
rect 2051 2562 2231 2566
rect 2235 2562 2335 2566
rect 2339 2562 2383 2566
rect 2387 2562 2447 2566
rect 2451 2562 2495 2566
rect 2499 2562 2559 2566
rect 2563 2562 2615 2566
rect 2619 2562 2671 2566
rect 2675 2562 2743 2566
rect 2747 2562 2791 2566
rect 2795 2562 2871 2566
rect 2875 2562 2911 2566
rect 2915 2562 2991 2566
rect 2995 2562 3031 2566
rect 3035 2562 3111 2566
rect 3115 2562 3151 2566
rect 3155 2562 3231 2566
rect 3235 2562 3359 2566
rect 3363 2562 3487 2566
rect 3491 2562 3943 2566
rect 3947 2562 3967 2566
rect 2025 2561 3967 2562
rect 3973 2561 3974 2567
rect 84 2489 85 2495
rect 91 2494 2019 2495
rect 91 2490 111 2494
rect 115 2490 135 2494
rect 139 2490 231 2494
rect 235 2490 287 2494
rect 291 2490 327 2494
rect 331 2490 423 2494
rect 427 2490 447 2494
rect 451 2490 519 2494
rect 523 2490 607 2494
rect 611 2490 767 2494
rect 771 2490 919 2494
rect 923 2490 1063 2494
rect 1067 2490 1199 2494
rect 1203 2490 1335 2494
rect 1339 2490 1463 2494
rect 1467 2490 1591 2494
rect 1595 2490 1727 2494
rect 1731 2490 2007 2494
rect 2011 2490 2019 2494
rect 91 2489 2019 2490
rect 2025 2489 2026 2495
rect 2030 2481 2031 2487
rect 2037 2486 3979 2487
rect 2037 2482 2047 2486
rect 2051 2482 2383 2486
rect 2387 2482 2495 2486
rect 2499 2482 2535 2486
rect 2539 2482 2615 2486
rect 2619 2482 2711 2486
rect 2715 2482 2743 2486
rect 2747 2482 2871 2486
rect 2875 2482 2879 2486
rect 2883 2482 2991 2486
rect 2995 2482 3047 2486
rect 3051 2482 3111 2486
rect 3115 2482 3207 2486
rect 3211 2482 3231 2486
rect 3235 2482 3359 2486
rect 3363 2482 3487 2486
rect 3491 2482 3503 2486
rect 3507 2482 3655 2486
rect 3659 2482 3807 2486
rect 3811 2482 3943 2486
rect 3947 2482 3979 2486
rect 2037 2481 3979 2482
rect 3985 2481 3986 2487
rect 2018 2407 2019 2413
rect 2025 2407 2050 2413
rect 96 2397 97 2403
rect 103 2402 2031 2403
rect 103 2398 111 2402
rect 115 2398 135 2402
rect 139 2398 231 2402
rect 235 2398 255 2402
rect 259 2398 327 2402
rect 331 2398 415 2402
rect 419 2398 423 2402
rect 427 2398 519 2402
rect 523 2398 575 2402
rect 579 2398 735 2402
rect 739 2398 887 2402
rect 891 2398 1039 2402
rect 1043 2398 1183 2402
rect 1187 2398 1327 2402
rect 1331 2398 1479 2402
rect 1483 2398 2007 2402
rect 2011 2398 2031 2402
rect 103 2397 2031 2398
rect 2037 2397 2038 2403
rect 2044 2399 2050 2407
rect 2044 2398 3967 2399
rect 2044 2394 2047 2398
rect 2051 2394 2535 2398
rect 2539 2394 2607 2398
rect 2611 2394 2711 2398
rect 2715 2394 2815 2398
rect 2819 2394 2879 2398
rect 2883 2394 3007 2398
rect 3011 2394 3047 2398
rect 3051 2394 3191 2398
rect 3195 2394 3207 2398
rect 3211 2394 3359 2398
rect 3363 2394 3503 2398
rect 3507 2394 3519 2398
rect 3523 2394 3655 2398
rect 3659 2394 3679 2398
rect 3683 2394 3807 2398
rect 3811 2394 3839 2398
rect 3843 2394 3943 2398
rect 3947 2394 3967 2398
rect 2044 2393 3967 2394
rect 3973 2393 3974 2399
rect 84 2321 85 2327
rect 91 2326 2019 2327
rect 91 2322 111 2326
rect 115 2322 135 2326
rect 139 2322 255 2326
rect 259 2322 263 2326
rect 267 2322 415 2326
rect 419 2322 423 2326
rect 427 2322 575 2326
rect 579 2322 583 2326
rect 587 2322 735 2326
rect 739 2322 743 2326
rect 747 2322 887 2326
rect 891 2322 895 2326
rect 899 2322 1039 2326
rect 1043 2322 1047 2326
rect 1051 2322 1183 2326
rect 1187 2322 1199 2326
rect 1203 2322 1327 2326
rect 1331 2322 1351 2326
rect 1355 2322 1479 2326
rect 1483 2322 1503 2326
rect 1507 2322 2007 2326
rect 2011 2322 2019 2326
rect 91 2321 2019 2322
rect 2025 2321 2026 2327
rect 2030 2301 2031 2307
rect 2037 2306 3979 2307
rect 2037 2302 2047 2306
rect 2051 2302 2071 2306
rect 2075 2302 2167 2306
rect 2171 2302 2271 2306
rect 2275 2302 2415 2306
rect 2419 2302 2575 2306
rect 2579 2302 2607 2306
rect 2611 2302 2743 2306
rect 2747 2302 2815 2306
rect 2819 2302 2911 2306
rect 2915 2302 3007 2306
rect 3011 2302 3071 2306
rect 3075 2302 3191 2306
rect 3195 2302 3231 2306
rect 3235 2302 3359 2306
rect 3363 2302 3383 2306
rect 3387 2302 3519 2306
rect 3523 2302 3535 2306
rect 3539 2302 3679 2306
rect 3683 2302 3695 2306
rect 3699 2302 3839 2306
rect 3843 2302 3943 2306
rect 3947 2302 3979 2306
rect 2037 2301 3979 2302
rect 3985 2301 3986 2307
rect 96 2241 97 2247
rect 103 2246 2031 2247
rect 103 2242 111 2246
rect 115 2242 135 2246
rect 139 2242 223 2246
rect 227 2242 263 2246
rect 267 2242 351 2246
rect 355 2242 423 2246
rect 427 2242 495 2246
rect 499 2242 583 2246
rect 587 2242 647 2246
rect 651 2242 743 2246
rect 747 2242 799 2246
rect 803 2242 895 2246
rect 899 2242 959 2246
rect 963 2242 1047 2246
rect 1051 2242 1119 2246
rect 1123 2242 1199 2246
rect 1203 2242 1279 2246
rect 1283 2242 1351 2246
rect 1355 2242 1439 2246
rect 1443 2242 1503 2246
rect 1507 2242 1599 2246
rect 1603 2242 2007 2246
rect 2011 2242 2031 2246
rect 103 2241 2031 2242
rect 2037 2241 2038 2247
rect 2018 2225 2019 2231
rect 2025 2230 3967 2231
rect 2025 2226 2047 2230
rect 2051 2226 2071 2230
rect 2075 2226 2167 2230
rect 2171 2226 2175 2230
rect 2179 2226 2271 2230
rect 2275 2226 2319 2230
rect 2323 2226 2415 2230
rect 2419 2226 2471 2230
rect 2475 2226 2575 2230
rect 2579 2226 2623 2230
rect 2627 2226 2743 2230
rect 2747 2226 2783 2230
rect 2787 2226 2911 2230
rect 2915 2226 2935 2230
rect 2939 2226 3071 2230
rect 3075 2226 3079 2230
rect 3083 2226 3223 2230
rect 3227 2226 3231 2230
rect 3235 2226 3367 2230
rect 3371 2226 3383 2230
rect 3387 2226 3519 2230
rect 3523 2226 3535 2230
rect 3539 2226 3695 2230
rect 3699 2226 3943 2230
rect 3947 2226 3967 2230
rect 2025 2225 3967 2226
rect 3973 2225 3974 2231
rect 84 2165 85 2171
rect 91 2170 2019 2171
rect 91 2166 111 2170
rect 115 2166 223 2170
rect 227 2166 351 2170
rect 355 2166 471 2170
rect 475 2166 495 2170
rect 499 2166 567 2170
rect 571 2166 647 2170
rect 651 2166 679 2170
rect 683 2166 799 2170
rect 803 2166 807 2170
rect 811 2166 943 2170
rect 947 2166 959 2170
rect 963 2166 1079 2170
rect 1083 2166 1119 2170
rect 1123 2166 1223 2170
rect 1227 2166 1279 2170
rect 1283 2166 1367 2170
rect 1371 2166 1439 2170
rect 1443 2166 1503 2170
rect 1507 2166 1599 2170
rect 1603 2166 1639 2170
rect 1643 2166 1783 2170
rect 1787 2166 1903 2170
rect 1907 2166 2007 2170
rect 2011 2166 2019 2170
rect 91 2165 2019 2166
rect 2025 2165 2026 2171
rect 2030 2129 2031 2135
rect 2037 2134 3979 2135
rect 2037 2130 2047 2134
rect 2051 2130 2071 2134
rect 2075 2130 2175 2134
rect 2179 2130 2279 2134
rect 2283 2130 2319 2134
rect 2323 2130 2391 2134
rect 2395 2130 2471 2134
rect 2475 2130 2511 2134
rect 2515 2130 2623 2134
rect 2627 2130 2631 2134
rect 2635 2130 2759 2134
rect 2763 2130 2783 2134
rect 2787 2130 2895 2134
rect 2899 2130 2935 2134
rect 2939 2130 3039 2134
rect 3043 2130 3079 2134
rect 3083 2130 3191 2134
rect 3195 2130 3223 2134
rect 3227 2130 3351 2134
rect 3355 2130 3367 2134
rect 3371 2130 3519 2134
rect 3523 2130 3687 2134
rect 3691 2130 3839 2134
rect 3843 2130 3943 2134
rect 3947 2130 3979 2134
rect 2037 2129 3979 2130
rect 3985 2129 3986 2135
rect 96 2089 97 2095
rect 103 2094 2031 2095
rect 103 2090 111 2094
rect 115 2090 471 2094
rect 475 2090 567 2094
rect 571 2090 623 2094
rect 627 2090 679 2094
rect 683 2090 735 2094
rect 739 2090 807 2094
rect 811 2090 855 2094
rect 859 2090 943 2094
rect 947 2090 983 2094
rect 987 2090 1079 2094
rect 1083 2090 1119 2094
rect 1123 2090 1223 2094
rect 1227 2090 1255 2094
rect 1259 2090 1367 2094
rect 1371 2090 1391 2094
rect 1395 2090 1503 2094
rect 1507 2090 1527 2094
rect 1531 2090 1639 2094
rect 1643 2090 1655 2094
rect 1659 2090 1783 2094
rect 1787 2090 1791 2094
rect 1795 2090 1903 2094
rect 1907 2090 2007 2094
rect 2011 2090 2031 2094
rect 103 2089 2031 2090
rect 2037 2089 2038 2095
rect 2018 2045 2019 2051
rect 2025 2050 3967 2051
rect 2025 2046 2047 2050
rect 2051 2046 2279 2050
rect 2283 2046 2327 2050
rect 2331 2046 2391 2050
rect 2395 2046 2431 2050
rect 2435 2046 2511 2050
rect 2515 2046 2535 2050
rect 2539 2046 2631 2050
rect 2635 2046 2647 2050
rect 2651 2046 2759 2050
rect 2763 2046 2775 2050
rect 2779 2046 2895 2050
rect 2899 2046 2919 2050
rect 2923 2046 3039 2050
rect 3043 2046 3079 2050
rect 3083 2046 3191 2050
rect 3195 2046 3263 2050
rect 3267 2046 3351 2050
rect 3355 2046 3455 2050
rect 3459 2046 3519 2050
rect 3523 2046 3655 2050
rect 3659 2046 3687 2050
rect 3691 2046 3839 2050
rect 3843 2046 3943 2050
rect 3947 2046 3967 2050
rect 2025 2045 3967 2046
rect 3973 2045 3974 2051
rect 84 2009 85 2015
rect 91 2014 2019 2015
rect 91 2010 111 2014
rect 115 2010 447 2014
rect 451 2010 575 2014
rect 579 2010 623 2014
rect 627 2010 727 2014
rect 731 2010 735 2014
rect 739 2010 855 2014
rect 859 2010 887 2014
rect 891 2010 983 2014
rect 987 2010 1055 2014
rect 1059 2010 1119 2014
rect 1123 2010 1231 2014
rect 1235 2010 1255 2014
rect 1259 2010 1391 2014
rect 1395 2010 1399 2014
rect 1403 2010 1527 2014
rect 1531 2010 1575 2014
rect 1579 2010 1655 2014
rect 1659 2010 1751 2014
rect 1755 2010 1791 2014
rect 1795 2010 1903 2014
rect 1907 2010 2007 2014
rect 2011 2010 2019 2014
rect 91 2009 2019 2010
rect 2025 2009 2026 2015
rect 2030 1965 2031 1971
rect 2037 1970 3979 1971
rect 2037 1966 2047 1970
rect 2051 1966 2255 1970
rect 2259 1966 2327 1970
rect 2331 1966 2351 1970
rect 2355 1966 2431 1970
rect 2435 1966 2447 1970
rect 2451 1966 2535 1970
rect 2539 1966 2543 1970
rect 2547 1966 2647 1970
rect 2651 1966 2767 1970
rect 2771 1966 2775 1970
rect 2779 1966 2919 1970
rect 2923 1966 3079 1970
rect 3083 1966 3103 1970
rect 3107 1966 3263 1970
rect 3267 1966 3319 1970
rect 3323 1966 3455 1970
rect 3459 1966 3543 1970
rect 3547 1966 3655 1970
rect 3659 1966 3775 1970
rect 3779 1966 3839 1970
rect 3843 1966 3943 1970
rect 3947 1966 3979 1970
rect 2037 1965 3979 1966
rect 3985 1965 3986 1971
rect 96 1933 97 1939
rect 103 1938 2031 1939
rect 103 1934 111 1938
rect 115 1934 447 1938
rect 451 1934 575 1938
rect 579 1934 655 1938
rect 659 1934 727 1938
rect 731 1934 751 1938
rect 755 1934 847 1938
rect 851 1934 887 1938
rect 891 1934 943 1938
rect 947 1934 1039 1938
rect 1043 1934 1055 1938
rect 1059 1934 1135 1938
rect 1139 1934 1231 1938
rect 1235 1934 1327 1938
rect 1331 1934 1399 1938
rect 1403 1934 1423 1938
rect 1427 1934 1575 1938
rect 1579 1934 1751 1938
rect 1755 1934 1903 1938
rect 1907 1934 2007 1938
rect 2011 1934 2031 1938
rect 103 1933 2031 1934
rect 2037 1933 2038 1939
rect 2018 1877 2019 1883
rect 2025 1882 3967 1883
rect 2025 1878 2047 1882
rect 2051 1878 2183 1882
rect 2187 1878 2255 1882
rect 2259 1878 2279 1882
rect 2283 1878 2351 1882
rect 2355 1878 2383 1882
rect 2387 1878 2447 1882
rect 2451 1878 2487 1882
rect 2491 1878 2543 1882
rect 2547 1878 2591 1882
rect 2595 1878 2647 1882
rect 2651 1878 2703 1882
rect 2707 1878 2767 1882
rect 2771 1878 2831 1882
rect 2835 1878 2919 1882
rect 2923 1878 2991 1882
rect 2995 1878 3103 1882
rect 3107 1878 3183 1882
rect 3187 1878 3319 1882
rect 3323 1878 3399 1882
rect 3403 1878 3543 1882
rect 3547 1878 3631 1882
rect 3635 1878 3775 1882
rect 3779 1878 3839 1882
rect 3843 1878 3943 1882
rect 3947 1878 3967 1882
rect 2025 1877 3967 1878
rect 3973 1877 3974 1883
rect 84 1857 85 1863
rect 91 1862 2019 1863
rect 91 1858 111 1862
rect 115 1858 319 1862
rect 323 1858 447 1862
rect 451 1858 583 1862
rect 587 1858 655 1862
rect 659 1858 719 1862
rect 723 1858 751 1862
rect 755 1858 847 1862
rect 851 1858 855 1862
rect 859 1858 943 1862
rect 947 1858 991 1862
rect 995 1858 1039 1862
rect 1043 1858 1127 1862
rect 1131 1858 1135 1862
rect 1139 1858 1231 1862
rect 1235 1858 1263 1862
rect 1267 1858 1327 1862
rect 1331 1858 1399 1862
rect 1403 1858 1423 1862
rect 1427 1858 1535 1862
rect 1539 1858 2007 1862
rect 2011 1858 2019 1862
rect 91 1857 2019 1858
rect 2025 1857 2026 1863
rect 2030 1797 2031 1803
rect 2037 1802 3979 1803
rect 2037 1798 2047 1802
rect 2051 1798 2127 1802
rect 2131 1798 2183 1802
rect 2187 1798 2279 1802
rect 2283 1798 2311 1802
rect 2315 1798 2383 1802
rect 2387 1798 2487 1802
rect 2491 1798 2495 1802
rect 2499 1798 2591 1802
rect 2595 1798 2687 1802
rect 2691 1798 2703 1802
rect 2707 1798 2831 1802
rect 2835 1798 2879 1802
rect 2883 1798 2991 1802
rect 2995 1798 3071 1802
rect 3075 1798 3183 1802
rect 3187 1798 3263 1802
rect 3267 1798 3399 1802
rect 3403 1798 3463 1802
rect 3467 1798 3631 1802
rect 3635 1798 3663 1802
rect 3667 1798 3839 1802
rect 3843 1798 3943 1802
rect 3947 1798 3979 1802
rect 2037 1797 3979 1798
rect 3985 1797 3986 1803
rect 96 1777 97 1783
rect 103 1782 2031 1783
rect 103 1778 111 1782
rect 115 1778 255 1782
rect 259 1778 319 1782
rect 323 1778 391 1782
rect 395 1778 447 1782
rect 451 1778 535 1782
rect 539 1778 583 1782
rect 587 1778 695 1782
rect 699 1778 719 1782
rect 723 1778 855 1782
rect 859 1778 863 1782
rect 867 1778 991 1782
rect 995 1778 1031 1782
rect 1035 1778 1127 1782
rect 1131 1778 1207 1782
rect 1211 1778 1263 1782
rect 1267 1778 1383 1782
rect 1387 1778 1399 1782
rect 1403 1778 1535 1782
rect 1539 1778 1559 1782
rect 1563 1778 1743 1782
rect 1747 1778 2007 1782
rect 2011 1778 2031 1782
rect 103 1777 2031 1778
rect 2037 1777 2038 1783
rect 2018 1717 2019 1723
rect 2025 1722 3967 1723
rect 2025 1718 2047 1722
rect 2051 1718 2071 1722
rect 2075 1718 2127 1722
rect 2131 1718 2191 1722
rect 2195 1718 2311 1722
rect 2315 1718 2343 1722
rect 2347 1718 2495 1722
rect 2499 1718 2511 1722
rect 2515 1718 2687 1722
rect 2691 1718 2871 1722
rect 2875 1718 2879 1722
rect 2883 1718 3063 1722
rect 3067 1718 3071 1722
rect 3075 1718 3255 1722
rect 3259 1718 3263 1722
rect 3267 1718 3447 1722
rect 3451 1718 3463 1722
rect 3467 1718 3647 1722
rect 3651 1718 3663 1722
rect 3667 1718 3839 1722
rect 3843 1718 3943 1722
rect 3947 1718 3967 1722
rect 2025 1717 3967 1718
rect 3973 1717 3974 1723
rect 84 1701 85 1707
rect 91 1706 2019 1707
rect 91 1702 111 1706
rect 115 1702 135 1706
rect 139 1702 255 1706
rect 259 1702 263 1706
rect 267 1702 391 1706
rect 395 1702 431 1706
rect 435 1702 535 1706
rect 539 1702 607 1706
rect 611 1702 695 1706
rect 699 1702 799 1706
rect 803 1702 863 1706
rect 867 1702 999 1706
rect 1003 1702 1031 1706
rect 1035 1702 1199 1706
rect 1203 1702 1207 1706
rect 1211 1702 1383 1706
rect 1387 1702 1407 1706
rect 1411 1702 1559 1706
rect 1563 1702 1623 1706
rect 1627 1702 1743 1706
rect 1747 1702 1839 1706
rect 1843 1702 2007 1706
rect 2011 1702 2019 1706
rect 91 1701 2019 1702
rect 2025 1701 2026 1707
rect 2030 1641 2031 1647
rect 2037 1646 3979 1647
rect 2037 1642 2047 1646
rect 2051 1642 2071 1646
rect 2075 1642 2191 1646
rect 2195 1642 2335 1646
rect 2339 1642 2343 1646
rect 2347 1642 2511 1646
rect 2515 1642 2599 1646
rect 2603 1642 2687 1646
rect 2691 1642 2839 1646
rect 2843 1642 2871 1646
rect 2875 1642 3047 1646
rect 3051 1642 3063 1646
rect 3067 1642 3231 1646
rect 3235 1642 3255 1646
rect 3259 1642 3399 1646
rect 3403 1642 3447 1646
rect 3451 1642 3551 1646
rect 3555 1642 3647 1646
rect 3651 1642 3695 1646
rect 3699 1642 3839 1646
rect 3843 1642 3943 1646
rect 3947 1642 3979 1646
rect 2037 1641 3979 1642
rect 3985 1641 3986 1647
rect 96 1625 97 1631
rect 103 1630 2031 1631
rect 103 1626 111 1630
rect 115 1626 135 1630
rect 139 1626 263 1630
rect 267 1626 287 1630
rect 291 1626 431 1630
rect 435 1626 471 1630
rect 475 1626 607 1630
rect 611 1626 655 1630
rect 659 1626 799 1630
rect 803 1626 839 1630
rect 843 1626 999 1630
rect 1003 1626 1015 1630
rect 1019 1626 1183 1630
rect 1187 1626 1199 1630
rect 1203 1626 1343 1630
rect 1347 1626 1407 1630
rect 1411 1626 1495 1630
rect 1499 1626 1623 1630
rect 1627 1626 1639 1630
rect 1643 1626 1783 1630
rect 1787 1626 1839 1630
rect 1843 1626 1903 1630
rect 1907 1626 2007 1630
rect 2011 1626 2031 1630
rect 103 1625 2031 1626
rect 2037 1625 2038 1631
rect 2018 1561 2019 1567
rect 2025 1566 3967 1567
rect 2025 1562 2047 1566
rect 2051 1562 2071 1566
rect 2075 1562 2335 1566
rect 2339 1562 2583 1566
rect 2587 1562 2599 1566
rect 2603 1562 2743 1566
rect 2747 1562 2839 1566
rect 2843 1562 2903 1566
rect 2907 1562 3047 1566
rect 3051 1562 3063 1566
rect 3067 1562 3223 1566
rect 3227 1562 3231 1566
rect 3235 1562 3383 1566
rect 3387 1562 3399 1566
rect 3403 1562 3543 1566
rect 3547 1562 3551 1566
rect 3555 1562 3695 1566
rect 3699 1562 3703 1566
rect 3707 1562 3839 1566
rect 3843 1562 3943 1566
rect 3947 1562 3967 1566
rect 2025 1561 3967 1562
rect 3973 1561 3974 1567
rect 84 1545 85 1551
rect 91 1550 2019 1551
rect 91 1546 111 1550
rect 115 1546 135 1550
rect 139 1546 287 1550
rect 291 1546 295 1550
rect 299 1546 471 1550
rect 475 1546 487 1550
rect 491 1546 655 1550
rect 659 1546 687 1550
rect 691 1546 839 1550
rect 843 1546 887 1550
rect 891 1546 1015 1550
rect 1019 1546 1079 1550
rect 1083 1546 1183 1550
rect 1187 1546 1263 1550
rect 1267 1546 1343 1550
rect 1347 1546 1447 1550
rect 1451 1546 1495 1550
rect 1499 1546 1623 1550
rect 1627 1546 1639 1550
rect 1643 1546 1783 1550
rect 1787 1546 1807 1550
rect 1811 1546 1903 1550
rect 1907 1546 2007 1550
rect 2011 1546 2019 1550
rect 91 1545 2019 1546
rect 2025 1545 2026 1551
rect 2030 1485 2031 1491
rect 2037 1490 3979 1491
rect 2037 1486 2047 1490
rect 2051 1486 2415 1490
rect 2419 1486 2511 1490
rect 2515 1486 2583 1490
rect 2587 1486 2607 1490
rect 2611 1486 2703 1490
rect 2707 1486 2743 1490
rect 2747 1486 2799 1490
rect 2803 1486 2903 1490
rect 2907 1486 2919 1490
rect 2923 1486 3063 1490
rect 3067 1486 3223 1490
rect 3227 1486 3231 1490
rect 3235 1486 3383 1490
rect 3387 1486 3415 1490
rect 3419 1486 3543 1490
rect 3547 1486 3615 1490
rect 3619 1486 3703 1490
rect 3707 1486 3815 1490
rect 3819 1486 3943 1490
rect 3947 1486 3979 1490
rect 2037 1485 3979 1486
rect 3985 1485 3986 1491
rect 96 1469 97 1475
rect 103 1474 2031 1475
rect 103 1470 111 1474
rect 115 1470 135 1474
rect 139 1470 175 1474
rect 179 1470 295 1474
rect 299 1470 359 1474
rect 363 1470 487 1474
rect 491 1470 567 1474
rect 571 1470 687 1474
rect 691 1470 783 1474
rect 787 1470 887 1474
rect 891 1470 1007 1474
rect 1011 1470 1079 1474
rect 1083 1470 1231 1474
rect 1235 1470 1263 1474
rect 1267 1470 1447 1474
rect 1451 1470 1463 1474
rect 1467 1470 1623 1474
rect 1627 1470 1695 1474
rect 1699 1470 1807 1474
rect 1811 1470 1903 1474
rect 1907 1470 2007 1474
rect 2011 1470 2031 1474
rect 103 1469 2031 1470
rect 2037 1469 2038 1475
rect 84 1393 85 1399
rect 91 1398 2019 1399
rect 91 1394 111 1398
rect 115 1394 175 1398
rect 179 1394 327 1398
rect 331 1394 359 1398
rect 363 1394 463 1398
rect 467 1394 567 1398
rect 571 1394 599 1398
rect 603 1394 727 1398
rect 731 1394 783 1398
rect 787 1394 855 1398
rect 859 1394 983 1398
rect 987 1394 1007 1398
rect 1011 1394 1119 1398
rect 1123 1394 1231 1398
rect 1235 1394 1263 1398
rect 1267 1394 1423 1398
rect 1427 1394 1463 1398
rect 1467 1394 1583 1398
rect 1587 1394 1695 1398
rect 1699 1394 1751 1398
rect 1755 1394 1903 1398
rect 1907 1394 2007 1398
rect 2011 1394 2019 1398
rect 91 1393 2019 1394
rect 2025 1395 2026 1399
rect 2025 1394 3974 1395
rect 2025 1393 2047 1394
rect 2018 1390 2047 1393
rect 2051 1390 2071 1394
rect 2075 1390 2303 1394
rect 2307 1390 2415 1394
rect 2419 1390 2511 1394
rect 2515 1390 2559 1394
rect 2563 1390 2607 1394
rect 2611 1390 2703 1394
rect 2707 1390 2799 1394
rect 2803 1390 2807 1394
rect 2811 1390 2919 1394
rect 2923 1390 3055 1394
rect 3059 1390 3063 1394
rect 3067 1390 3231 1394
rect 3235 1390 3303 1394
rect 3307 1390 3415 1394
rect 3419 1390 3559 1394
rect 3563 1390 3615 1394
rect 3619 1390 3815 1394
rect 3819 1390 3943 1394
rect 3947 1390 3974 1394
rect 2018 1389 3974 1390
rect 96 1309 97 1315
rect 103 1314 2031 1315
rect 103 1310 111 1314
rect 115 1310 327 1314
rect 331 1310 463 1314
rect 467 1310 551 1314
rect 555 1310 599 1314
rect 603 1310 655 1314
rect 659 1310 727 1314
rect 731 1310 767 1314
rect 771 1310 855 1314
rect 859 1310 879 1314
rect 883 1310 983 1314
rect 987 1310 991 1314
rect 995 1310 1103 1314
rect 1107 1310 1119 1314
rect 1123 1310 1215 1314
rect 1219 1310 1263 1314
rect 1267 1310 1327 1314
rect 1331 1310 1423 1314
rect 1427 1310 1439 1314
rect 1443 1310 1559 1314
rect 1563 1310 1583 1314
rect 1587 1310 1751 1314
rect 1755 1310 1903 1314
rect 1907 1310 2007 1314
rect 2011 1310 2031 1314
rect 103 1309 2031 1310
rect 2037 1311 2038 1315
rect 2037 1310 3986 1311
rect 2037 1309 2047 1310
rect 2030 1306 2047 1309
rect 2051 1306 2071 1310
rect 2075 1306 2223 1310
rect 2227 1306 2303 1310
rect 2307 1306 2415 1310
rect 2419 1306 2559 1310
rect 2563 1306 2615 1310
rect 2619 1306 2807 1310
rect 2811 1306 2815 1310
rect 2819 1306 2999 1310
rect 3003 1306 3055 1310
rect 3059 1306 3175 1310
rect 3179 1306 3303 1310
rect 3307 1306 3343 1310
rect 3347 1306 3503 1310
rect 3507 1306 3559 1310
rect 3563 1306 3663 1310
rect 3667 1306 3815 1310
rect 3819 1306 3831 1310
rect 3835 1306 3943 1310
rect 3947 1306 3986 1310
rect 2030 1305 3986 1306
rect 84 1233 85 1239
rect 91 1238 2019 1239
rect 91 1234 111 1238
rect 115 1234 391 1238
rect 395 1234 519 1238
rect 523 1234 551 1238
rect 555 1234 655 1238
rect 659 1234 663 1238
rect 667 1234 767 1238
rect 771 1234 807 1238
rect 811 1234 879 1238
rect 883 1234 959 1238
rect 963 1234 991 1238
rect 995 1234 1103 1238
rect 1107 1234 1111 1238
rect 1115 1234 1215 1238
rect 1219 1234 1255 1238
rect 1259 1234 1327 1238
rect 1331 1234 1407 1238
rect 1411 1234 1439 1238
rect 1443 1234 1559 1238
rect 1563 1234 1711 1238
rect 1715 1234 2007 1238
rect 2011 1234 2019 1238
rect 91 1233 2019 1234
rect 2025 1233 2026 1239
rect 2018 1221 2019 1227
rect 2025 1226 3967 1227
rect 2025 1222 2047 1226
rect 2051 1222 2071 1226
rect 2075 1222 2135 1226
rect 2139 1222 2223 1226
rect 2227 1222 2311 1226
rect 2315 1222 2415 1226
rect 2419 1222 2503 1226
rect 2507 1222 2615 1226
rect 2619 1222 2695 1226
rect 2699 1222 2815 1226
rect 2819 1222 2887 1226
rect 2891 1222 2999 1226
rect 3003 1222 3071 1226
rect 3075 1222 3175 1226
rect 3179 1222 3239 1226
rect 3243 1222 3343 1226
rect 3347 1222 3399 1226
rect 3403 1222 3503 1226
rect 3507 1222 3551 1226
rect 3555 1222 3663 1226
rect 3667 1222 3703 1226
rect 3707 1222 3831 1226
rect 3835 1222 3839 1226
rect 3843 1222 3943 1226
rect 3947 1222 3967 1226
rect 2025 1221 3967 1222
rect 3973 1221 3974 1227
rect 96 1153 97 1159
rect 103 1158 2031 1159
rect 103 1154 111 1158
rect 115 1154 175 1158
rect 179 1154 327 1158
rect 331 1154 391 1158
rect 395 1154 495 1158
rect 499 1154 519 1158
rect 523 1154 663 1158
rect 667 1154 671 1158
rect 675 1154 807 1158
rect 811 1154 847 1158
rect 851 1154 959 1158
rect 963 1154 1031 1158
rect 1035 1154 1111 1158
rect 1115 1154 1207 1158
rect 1211 1154 1255 1158
rect 1259 1154 1383 1158
rect 1387 1154 1407 1158
rect 1411 1154 1559 1158
rect 1563 1154 1567 1158
rect 1571 1154 1711 1158
rect 1715 1154 1751 1158
rect 1755 1154 2007 1158
rect 2011 1154 2031 1158
rect 103 1153 2031 1154
rect 2037 1153 2038 1159
rect 2030 1137 2031 1143
rect 2037 1142 3979 1143
rect 2037 1138 2047 1142
rect 2051 1138 2135 1142
rect 2139 1138 2295 1142
rect 2299 1138 2311 1142
rect 2315 1138 2423 1142
rect 2427 1138 2503 1142
rect 2507 1138 2559 1142
rect 2563 1138 2695 1142
rect 2699 1138 2839 1142
rect 2843 1138 2887 1142
rect 2891 1138 2991 1142
rect 2995 1138 3071 1142
rect 3075 1138 3151 1142
rect 3155 1138 3239 1142
rect 3243 1138 3319 1142
rect 3323 1138 3399 1142
rect 3403 1138 3495 1142
rect 3499 1138 3551 1142
rect 3555 1138 3679 1142
rect 3683 1138 3703 1142
rect 3707 1138 3839 1142
rect 3843 1138 3943 1142
rect 3947 1138 3979 1142
rect 2037 1137 3979 1138
rect 3985 1137 3986 1143
rect 84 1069 85 1075
rect 91 1074 2019 1075
rect 91 1070 111 1074
rect 115 1070 135 1074
rect 139 1070 175 1074
rect 179 1070 231 1074
rect 235 1070 327 1074
rect 331 1070 375 1074
rect 379 1070 495 1074
rect 499 1070 543 1074
rect 547 1070 671 1074
rect 675 1070 727 1074
rect 731 1070 847 1074
rect 851 1070 911 1074
rect 915 1070 1031 1074
rect 1035 1070 1095 1074
rect 1099 1070 1207 1074
rect 1211 1070 1279 1074
rect 1283 1070 1383 1074
rect 1387 1070 1463 1074
rect 1467 1070 1567 1074
rect 1571 1070 1647 1074
rect 1651 1070 1751 1074
rect 1755 1070 1831 1074
rect 1835 1070 2007 1074
rect 2011 1070 2019 1074
rect 91 1069 2019 1070
rect 2025 1069 2026 1075
rect 2018 1057 2019 1063
rect 2025 1062 3967 1063
rect 2025 1058 2047 1062
rect 2051 1058 2295 1062
rect 2299 1058 2423 1062
rect 2427 1058 2495 1062
rect 2499 1058 2559 1062
rect 2563 1058 2599 1062
rect 2603 1058 2695 1062
rect 2699 1058 2711 1062
rect 2715 1058 2839 1062
rect 2843 1058 2847 1062
rect 2851 1058 2991 1062
rect 2995 1058 3007 1062
rect 3011 1058 3151 1062
rect 3155 1058 3199 1062
rect 3203 1058 3319 1062
rect 3323 1058 3407 1062
rect 3411 1058 3495 1062
rect 3499 1058 3631 1062
rect 3635 1058 3679 1062
rect 3683 1058 3839 1062
rect 3843 1058 3943 1062
rect 3947 1058 3967 1062
rect 2025 1057 3967 1058
rect 3973 1057 3974 1063
rect 96 993 97 999
rect 103 998 2031 999
rect 103 994 111 998
rect 115 994 135 998
rect 139 994 231 998
rect 235 994 271 998
rect 275 994 375 998
rect 379 994 447 998
rect 451 994 543 998
rect 547 994 631 998
rect 635 994 727 998
rect 731 994 823 998
rect 827 994 911 998
rect 915 994 1007 998
rect 1011 994 1095 998
rect 1099 994 1175 998
rect 1179 994 1279 998
rect 1283 994 1335 998
rect 1339 994 1463 998
rect 1467 994 1487 998
rect 1491 994 1631 998
rect 1635 994 1647 998
rect 1651 994 1775 998
rect 1779 994 1831 998
rect 1835 994 1903 998
rect 1907 994 2007 998
rect 2011 994 2031 998
rect 103 993 2031 994
rect 2037 993 2038 999
rect 2030 981 2031 987
rect 2037 986 3979 987
rect 2037 982 2047 986
rect 2051 982 2495 986
rect 2499 982 2599 986
rect 2603 982 2647 986
rect 2651 982 2711 986
rect 2715 982 2743 986
rect 2747 982 2847 986
rect 2851 982 2967 986
rect 2971 982 3007 986
rect 3011 982 3111 986
rect 3115 982 3199 986
rect 3203 982 3279 986
rect 3283 982 3407 986
rect 3411 982 3463 986
rect 3467 982 3631 986
rect 3635 982 3663 986
rect 3667 982 3839 986
rect 3843 982 3943 986
rect 3947 982 3979 986
rect 2037 981 3979 982
rect 3985 981 3986 987
rect 84 917 85 923
rect 91 922 2019 923
rect 91 918 111 922
rect 115 918 135 922
rect 139 918 271 922
rect 275 918 447 922
rect 451 918 455 922
rect 459 918 631 922
rect 635 918 655 922
rect 659 918 823 922
rect 827 918 855 922
rect 859 918 1007 922
rect 1011 918 1055 922
rect 1059 918 1175 922
rect 1179 918 1239 922
rect 1243 918 1335 922
rect 1339 918 1415 922
rect 1419 918 1487 922
rect 1491 918 1583 922
rect 1587 918 1631 922
rect 1635 918 1751 922
rect 1755 918 1775 922
rect 1779 918 1903 922
rect 1907 918 2007 922
rect 2011 918 2019 922
rect 91 917 2019 918
rect 2025 917 2026 923
rect 2018 893 2019 899
rect 2025 898 3967 899
rect 2025 894 2047 898
rect 2051 894 2071 898
rect 2075 894 2255 898
rect 2259 894 2463 898
rect 2467 894 2647 898
rect 2651 894 2679 898
rect 2683 894 2743 898
rect 2747 894 2847 898
rect 2851 894 2895 898
rect 2899 894 2967 898
rect 2971 894 3111 898
rect 3115 894 3127 898
rect 3131 894 3279 898
rect 3283 894 3367 898
rect 3371 894 3463 898
rect 3467 894 3615 898
rect 3619 894 3663 898
rect 3667 894 3839 898
rect 3843 894 3943 898
rect 3947 894 3967 898
rect 2025 893 3967 894
rect 3973 893 3974 899
rect 96 841 97 847
rect 103 846 2031 847
rect 103 842 111 846
rect 115 842 135 846
rect 139 842 215 846
rect 219 842 271 846
rect 275 842 343 846
rect 347 842 455 846
rect 459 842 495 846
rect 499 842 655 846
rect 659 842 831 846
rect 835 842 855 846
rect 859 842 1007 846
rect 1011 842 1055 846
rect 1059 842 1183 846
rect 1187 842 1239 846
rect 1243 842 1359 846
rect 1363 842 1415 846
rect 1419 842 1535 846
rect 1539 842 1583 846
rect 1587 842 1719 846
rect 1723 842 1751 846
rect 1755 842 1903 846
rect 1907 842 2007 846
rect 2011 842 2031 846
rect 103 841 2031 842
rect 2037 841 2038 847
rect 2030 817 2031 823
rect 2037 822 3979 823
rect 2037 818 2047 822
rect 2051 818 2071 822
rect 2075 818 2215 822
rect 2219 818 2255 822
rect 2259 818 2327 822
rect 2331 818 2447 822
rect 2451 818 2463 822
rect 2467 818 2583 822
rect 2587 818 2679 822
rect 2683 818 2735 822
rect 2739 818 2895 822
rect 2899 818 3063 822
rect 3067 818 3127 822
rect 3131 818 3247 822
rect 3251 818 3367 822
rect 3371 818 3447 822
rect 3451 818 3615 822
rect 3619 818 3655 822
rect 3659 818 3839 822
rect 3843 818 3943 822
rect 3947 818 3979 822
rect 2037 817 3979 818
rect 3985 817 3986 823
rect 84 765 85 771
rect 91 770 2019 771
rect 91 766 111 770
rect 115 766 215 770
rect 219 766 343 770
rect 347 766 375 770
rect 379 766 495 770
rect 499 766 623 770
rect 627 766 655 770
rect 659 766 751 770
rect 755 766 831 770
rect 835 766 887 770
rect 891 766 1007 770
rect 1011 766 1023 770
rect 1027 766 1167 770
rect 1171 766 1183 770
rect 1187 766 1311 770
rect 1315 766 1359 770
rect 1363 766 1455 770
rect 1459 766 1535 770
rect 1539 766 1599 770
rect 1603 766 1719 770
rect 1723 766 2007 770
rect 2011 766 2019 770
rect 91 765 2019 766
rect 2025 765 2026 771
rect 2018 737 2019 743
rect 2025 742 3967 743
rect 2025 738 2047 742
rect 2051 738 2215 742
rect 2219 738 2327 742
rect 2331 738 2375 742
rect 2379 738 2447 742
rect 2451 738 2495 742
rect 2499 738 2583 742
rect 2587 738 2623 742
rect 2627 738 2735 742
rect 2739 738 2767 742
rect 2771 738 2895 742
rect 2899 738 2911 742
rect 2915 738 3063 742
rect 3067 738 3215 742
rect 3219 738 3247 742
rect 3251 738 3367 742
rect 3371 738 3447 742
rect 3451 738 3519 742
rect 3523 738 3655 742
rect 3659 738 3679 742
rect 3683 738 3839 742
rect 3843 738 3943 742
rect 3947 738 3967 742
rect 2025 737 3967 738
rect 3973 737 3974 743
rect 96 689 97 695
rect 103 694 2031 695
rect 103 690 111 694
rect 115 690 375 694
rect 379 690 495 694
rect 499 690 527 694
rect 531 690 623 694
rect 627 690 631 694
rect 635 690 743 694
rect 747 690 751 694
rect 755 690 855 694
rect 859 690 887 694
rect 891 690 967 694
rect 971 690 1023 694
rect 1027 690 1071 694
rect 1075 690 1167 694
rect 1171 690 1183 694
rect 1187 690 1295 694
rect 1299 690 1311 694
rect 1315 690 1407 694
rect 1411 690 1455 694
rect 1459 690 1519 694
rect 1523 690 1599 694
rect 1603 690 2007 694
rect 2011 690 2031 694
rect 103 689 2031 690
rect 2037 689 2038 695
rect 2030 653 2031 659
rect 2037 658 3979 659
rect 2037 654 2047 658
rect 2051 654 2111 658
rect 2115 654 2247 658
rect 2251 654 2375 658
rect 2379 654 2399 658
rect 2403 654 2495 658
rect 2499 654 2575 658
rect 2579 654 2623 658
rect 2627 654 2759 658
rect 2763 654 2767 658
rect 2771 654 2911 658
rect 2915 654 2943 658
rect 2947 654 3063 658
rect 3067 654 3127 658
rect 3131 654 3215 658
rect 3219 654 3303 658
rect 3307 654 3367 658
rect 3371 654 3479 658
rect 3483 654 3519 658
rect 3523 654 3655 658
rect 3659 654 3679 658
rect 3683 654 3831 658
rect 3835 654 3839 658
rect 3843 654 3943 658
rect 3947 654 3979 658
rect 2037 653 3979 654
rect 3985 653 3986 659
rect 84 613 85 619
rect 91 618 2019 619
rect 91 614 111 618
rect 115 614 527 618
rect 531 614 631 618
rect 635 614 687 618
rect 691 614 743 618
rect 747 614 783 618
rect 787 614 855 618
rect 859 614 879 618
rect 883 614 967 618
rect 971 614 975 618
rect 979 614 1071 618
rect 1075 614 1167 618
rect 1171 614 1183 618
rect 1187 614 1263 618
rect 1267 614 1295 618
rect 1299 614 1359 618
rect 1363 614 1407 618
rect 1411 614 1455 618
rect 1459 614 1519 618
rect 1523 614 2007 618
rect 2011 614 2019 618
rect 91 613 2019 614
rect 2025 613 2026 619
rect 2018 573 2019 579
rect 2025 578 3967 579
rect 2025 574 2047 578
rect 2051 574 2071 578
rect 2075 574 2111 578
rect 2115 574 2183 578
rect 2187 574 2247 578
rect 2251 574 2335 578
rect 2339 574 2399 578
rect 2403 574 2503 578
rect 2507 574 2575 578
rect 2579 574 2687 578
rect 2691 574 2759 578
rect 2763 574 2879 578
rect 2883 574 2943 578
rect 2947 574 3071 578
rect 3075 574 3127 578
rect 3131 574 3263 578
rect 3267 574 3303 578
rect 3307 574 3455 578
rect 3459 574 3479 578
rect 3483 574 3647 578
rect 3651 574 3655 578
rect 3659 574 3831 578
rect 3835 574 3839 578
rect 3843 574 3943 578
rect 3947 574 3967 578
rect 2025 573 3967 574
rect 3973 573 3974 579
rect 96 517 97 523
rect 103 522 2031 523
rect 103 518 111 522
rect 115 518 383 522
rect 387 518 479 522
rect 483 518 575 522
rect 579 518 671 522
rect 675 518 687 522
rect 691 518 767 522
rect 771 518 783 522
rect 787 518 863 522
rect 867 518 879 522
rect 883 518 959 522
rect 963 518 975 522
rect 979 518 1055 522
rect 1059 518 1071 522
rect 1075 518 1151 522
rect 1155 518 1167 522
rect 1171 518 1247 522
rect 1251 518 1263 522
rect 1267 518 1343 522
rect 1347 518 1359 522
rect 1363 518 1439 522
rect 1443 518 1455 522
rect 1459 518 1535 522
rect 1539 518 2007 522
rect 2011 518 2031 522
rect 103 517 2031 518
rect 2037 517 2038 523
rect 2030 497 2031 503
rect 2037 502 3979 503
rect 2037 498 2047 502
rect 2051 498 2071 502
rect 2075 498 2183 502
rect 2187 498 2319 502
rect 2323 498 2335 502
rect 2339 498 2463 502
rect 2467 498 2503 502
rect 2507 498 2615 502
rect 2619 498 2687 502
rect 2691 498 2775 502
rect 2779 498 2879 502
rect 2883 498 2959 502
rect 2963 498 3071 502
rect 3075 498 3159 502
rect 3163 498 3263 502
rect 3267 498 3367 502
rect 3371 498 3455 502
rect 3459 498 3583 502
rect 3587 498 3647 502
rect 3651 498 3807 502
rect 3811 498 3839 502
rect 3843 498 3943 502
rect 3947 498 3979 502
rect 2037 497 3979 498
rect 3985 497 3986 503
rect 84 429 85 435
rect 91 434 2019 435
rect 91 430 111 434
rect 115 430 383 434
rect 387 430 479 434
rect 483 430 487 434
rect 491 430 575 434
rect 579 430 583 434
rect 587 430 671 434
rect 675 430 687 434
rect 691 430 767 434
rect 771 430 791 434
rect 795 430 863 434
rect 867 430 895 434
rect 899 430 959 434
rect 963 430 999 434
rect 1003 430 1055 434
rect 1059 430 1103 434
rect 1107 430 1151 434
rect 1155 430 1207 434
rect 1211 430 1247 434
rect 1251 430 1319 434
rect 1323 430 1343 434
rect 1347 430 1431 434
rect 1435 430 1439 434
rect 1443 430 1535 434
rect 1539 430 2007 434
rect 2011 430 2019 434
rect 91 429 2019 430
rect 2025 429 2026 435
rect 2018 427 2026 429
rect 2018 421 2019 427
rect 2025 426 3967 427
rect 2025 422 2047 426
rect 2051 422 2183 426
rect 2187 422 2319 426
rect 2323 422 2343 426
rect 2347 422 2463 426
rect 2467 422 2487 426
rect 2491 422 2615 426
rect 2619 422 2639 426
rect 2643 422 2775 426
rect 2779 422 2799 426
rect 2803 422 2959 426
rect 2963 422 3111 426
rect 3115 422 3159 426
rect 3163 422 3263 426
rect 3267 422 3367 426
rect 3371 422 3415 426
rect 3419 422 3559 426
rect 3563 422 3583 426
rect 3587 422 3711 426
rect 3715 422 3807 426
rect 3811 422 3839 426
rect 3843 422 3943 426
rect 3947 422 3967 426
rect 2025 421 3967 422
rect 3973 421 3974 427
rect 96 349 97 355
rect 103 354 2031 355
rect 103 350 111 354
rect 115 350 327 354
rect 331 350 463 354
rect 467 350 487 354
rect 491 350 583 354
rect 587 350 615 354
rect 619 350 687 354
rect 691 350 767 354
rect 771 350 791 354
rect 795 350 895 354
rect 899 350 919 354
rect 923 350 999 354
rect 1003 350 1063 354
rect 1067 350 1103 354
rect 1107 350 1207 354
rect 1211 350 1319 354
rect 1323 350 1351 354
rect 1355 350 1431 354
rect 1435 350 1495 354
rect 1499 350 1639 354
rect 1643 350 2007 354
rect 2011 350 2031 354
rect 103 349 2031 350
rect 2037 349 2038 355
rect 2030 347 2038 349
rect 2030 341 2031 347
rect 2037 346 3979 347
rect 2037 342 2047 346
rect 2051 342 2343 346
rect 2347 342 2487 346
rect 2491 342 2495 346
rect 2499 342 2639 346
rect 2643 342 2799 346
rect 2803 342 2959 346
rect 2963 342 3111 346
rect 3115 342 3119 346
rect 3123 342 3263 346
rect 3267 342 3271 346
rect 3275 342 3415 346
rect 3419 342 3423 346
rect 3427 342 3559 346
rect 3563 342 3567 346
rect 3571 342 3711 346
rect 3715 342 3839 346
rect 3843 342 3943 346
rect 3947 342 3979 346
rect 2037 341 3979 342
rect 3985 341 3986 347
rect 84 265 85 271
rect 91 270 2019 271
rect 91 266 111 270
rect 115 266 167 270
rect 171 266 327 270
rect 331 266 463 270
rect 467 266 503 270
rect 507 266 615 270
rect 619 266 687 270
rect 691 266 767 270
rect 771 266 871 270
rect 875 266 919 270
rect 923 266 1047 270
rect 1051 266 1063 270
rect 1067 266 1207 270
rect 1211 266 1215 270
rect 1219 266 1351 270
rect 1355 266 1367 270
rect 1371 266 1495 270
rect 1499 266 1511 270
rect 1515 266 1639 270
rect 1643 266 1647 270
rect 1651 266 1783 270
rect 1787 266 1903 270
rect 1907 266 2007 270
rect 2011 266 2019 270
rect 91 265 2019 266
rect 2025 270 3974 271
rect 2025 266 2047 270
rect 2051 266 2071 270
rect 2075 266 2271 270
rect 2275 266 2495 270
rect 2499 266 2639 270
rect 2643 266 2703 270
rect 2707 266 2799 270
rect 2803 266 2903 270
rect 2907 266 2959 270
rect 2963 266 3095 270
rect 3099 266 3119 270
rect 3123 266 3271 270
rect 3275 266 3287 270
rect 3291 266 3423 270
rect 3427 266 3479 270
rect 3483 266 3567 270
rect 3571 266 3671 270
rect 3675 266 3711 270
rect 3715 266 3839 270
rect 3843 266 3943 270
rect 3947 266 3974 270
rect 2025 265 3974 266
rect 2030 170 3986 171
rect 2030 167 2047 170
rect 96 161 97 167
rect 103 166 2031 167
rect 103 162 111 166
rect 115 162 135 166
rect 139 162 167 166
rect 171 162 231 166
rect 235 162 327 166
rect 331 162 423 166
rect 427 162 503 166
rect 507 162 527 166
rect 531 162 647 166
rect 651 162 687 166
rect 691 162 775 166
rect 779 162 871 166
rect 875 162 903 166
rect 907 162 1031 166
rect 1035 162 1047 166
rect 1051 162 1151 166
rect 1155 162 1215 166
rect 1219 162 1271 166
rect 1275 162 1367 166
rect 1371 162 1383 166
rect 1387 162 1487 166
rect 1491 162 1511 166
rect 1515 162 1591 166
rect 1595 162 1647 166
rect 1651 162 1703 166
rect 1707 162 1783 166
rect 1787 162 1807 166
rect 1811 162 1903 166
rect 1907 162 2007 166
rect 2011 162 2031 166
rect 103 161 2031 162
rect 2037 166 2047 167
rect 2051 166 2071 170
rect 2075 166 2167 170
rect 2171 166 2263 170
rect 2267 166 2271 170
rect 2275 166 2359 170
rect 2363 166 2455 170
rect 2459 166 2495 170
rect 2499 166 2551 170
rect 2555 166 2655 170
rect 2659 166 2703 170
rect 2707 166 2759 170
rect 2763 166 2863 170
rect 2867 166 2903 170
rect 2907 166 2975 170
rect 2979 166 3095 170
rect 3099 166 3103 170
rect 3107 166 3239 170
rect 3243 166 3287 170
rect 3291 166 3383 170
rect 3387 166 3479 170
rect 3483 166 3535 170
rect 3539 166 3671 170
rect 3675 166 3695 170
rect 3699 166 3839 170
rect 3843 166 3943 170
rect 3947 166 3986 170
rect 2037 165 3986 166
rect 2037 161 2038 165
rect 2018 94 3974 95
rect 2018 91 2047 94
rect 84 85 85 91
rect 91 90 2019 91
rect 91 86 111 90
rect 115 86 135 90
rect 139 86 231 90
rect 235 86 327 90
rect 331 86 423 90
rect 427 86 527 90
rect 531 86 647 90
rect 651 86 775 90
rect 779 86 903 90
rect 907 86 1031 90
rect 1035 86 1151 90
rect 1155 86 1271 90
rect 1275 86 1383 90
rect 1387 86 1487 90
rect 1491 86 1591 90
rect 1595 86 1703 90
rect 1707 86 1807 90
rect 1811 86 1903 90
rect 1907 86 2007 90
rect 2011 86 2019 90
rect 91 85 2019 86
rect 2025 90 2047 91
rect 2051 90 2071 94
rect 2075 90 2167 94
rect 2171 90 2263 94
rect 2267 90 2359 94
rect 2363 90 2455 94
rect 2459 90 2551 94
rect 2555 90 2655 94
rect 2659 90 2759 94
rect 2763 90 2863 94
rect 2867 90 2975 94
rect 2979 90 3103 94
rect 3107 90 3239 94
rect 3243 90 3383 94
rect 3387 90 3535 94
rect 3539 90 3695 94
rect 3699 90 3839 94
rect 3843 90 3943 94
rect 3947 90 3974 94
rect 2025 89 3974 90
rect 2025 85 2026 89
<< m5c >>
rect 97 4025 103 4031
rect 2031 4025 2037 4031
rect 2019 4013 2025 4019
rect 3967 4013 3973 4019
rect 85 3949 91 3955
rect 2019 3949 2025 3955
rect 2031 3937 2037 3943
rect 3979 3937 3985 3943
rect 97 3873 103 3879
rect 2031 3873 2037 3879
rect 2019 3853 2025 3859
rect 3967 3853 3973 3859
rect 85 3793 91 3799
rect 2019 3793 2025 3799
rect 2031 3777 2037 3783
rect 3979 3777 3985 3783
rect 97 3709 103 3715
rect 2031 3709 2037 3715
rect 2019 3697 2025 3703
rect 3967 3697 3973 3703
rect 85 3625 91 3631
rect 2019 3625 2025 3631
rect 2031 3613 2037 3619
rect 3979 3613 3985 3619
rect 2019 3547 2025 3553
rect 97 3537 103 3543
rect 2031 3537 2037 3543
rect 3967 3537 3973 3543
rect 85 3453 91 3459
rect 2019 3453 2025 3459
rect 2031 3457 2037 3463
rect 3979 3457 3985 3463
rect 97 3377 103 3383
rect 2031 3377 2037 3383
rect 2019 3365 2025 3371
rect 3967 3365 3973 3371
rect 85 3301 91 3307
rect 2019 3301 2025 3307
rect 2031 3281 2037 3287
rect 3979 3281 3985 3287
rect 97 3225 103 3231
rect 2031 3225 2037 3231
rect 2019 3205 2025 3211
rect 3967 3205 3973 3211
rect 85 3145 91 3151
rect 2019 3145 2025 3151
rect 2031 3117 2037 3123
rect 3979 3117 3985 3123
rect 97 3061 103 3067
rect 2031 3061 2037 3067
rect 2019 3041 2025 3047
rect 3967 3041 3973 3047
rect 85 2981 91 2987
rect 2019 2981 2025 2987
rect 2031 2961 2037 2967
rect 3979 2961 3985 2967
rect 97 2897 103 2903
rect 2031 2897 2037 2903
rect 2019 2885 2025 2891
rect 3967 2885 3973 2891
rect 85 2817 91 2823
rect 2019 2817 2025 2823
rect 2031 2805 2037 2811
rect 3979 2805 3985 2811
rect 97 2737 103 2743
rect 2031 2737 2037 2743
rect 2019 2725 2025 2731
rect 3967 2725 3973 2731
rect 85 2657 91 2663
rect 2019 2657 2025 2663
rect 2031 2641 2037 2647
rect 3979 2641 3985 2647
rect 97 2581 103 2587
rect 2031 2581 2037 2587
rect 2019 2561 2025 2567
rect 3967 2561 3973 2567
rect 85 2489 91 2495
rect 2019 2489 2025 2495
rect 2031 2481 2037 2487
rect 3979 2481 3985 2487
rect 2019 2407 2025 2413
rect 97 2397 103 2403
rect 2031 2397 2037 2403
rect 3967 2393 3973 2399
rect 85 2321 91 2327
rect 2019 2321 2025 2327
rect 2031 2301 2037 2307
rect 3979 2301 3985 2307
rect 97 2241 103 2247
rect 2031 2241 2037 2247
rect 2019 2225 2025 2231
rect 3967 2225 3973 2231
rect 85 2165 91 2171
rect 2019 2165 2025 2171
rect 2031 2129 2037 2135
rect 3979 2129 3985 2135
rect 97 2089 103 2095
rect 2031 2089 2037 2095
rect 2019 2045 2025 2051
rect 3967 2045 3973 2051
rect 85 2009 91 2015
rect 2019 2009 2025 2015
rect 2031 1965 2037 1971
rect 3979 1965 3985 1971
rect 97 1933 103 1939
rect 2031 1933 2037 1939
rect 2019 1877 2025 1883
rect 3967 1877 3973 1883
rect 85 1857 91 1863
rect 2019 1857 2025 1863
rect 2031 1797 2037 1803
rect 3979 1797 3985 1803
rect 97 1777 103 1783
rect 2031 1777 2037 1783
rect 2019 1717 2025 1723
rect 3967 1717 3973 1723
rect 85 1701 91 1707
rect 2019 1701 2025 1707
rect 2031 1641 2037 1647
rect 3979 1641 3985 1647
rect 97 1625 103 1631
rect 2031 1625 2037 1631
rect 2019 1561 2025 1567
rect 3967 1561 3973 1567
rect 85 1545 91 1551
rect 2019 1545 2025 1551
rect 2031 1485 2037 1491
rect 3979 1485 3985 1491
rect 97 1469 103 1475
rect 2031 1469 2037 1475
rect 85 1393 91 1399
rect 2019 1393 2025 1399
rect 97 1309 103 1315
rect 2031 1309 2037 1315
rect 85 1233 91 1239
rect 2019 1233 2025 1239
rect 2019 1221 2025 1227
rect 3967 1221 3973 1227
rect 97 1153 103 1159
rect 2031 1153 2037 1159
rect 2031 1137 2037 1143
rect 3979 1137 3985 1143
rect 85 1069 91 1075
rect 2019 1069 2025 1075
rect 2019 1057 2025 1063
rect 3967 1057 3973 1063
rect 97 993 103 999
rect 2031 993 2037 999
rect 2031 981 2037 987
rect 3979 981 3985 987
rect 85 917 91 923
rect 2019 917 2025 923
rect 2019 893 2025 899
rect 3967 893 3973 899
rect 97 841 103 847
rect 2031 841 2037 847
rect 2031 817 2037 823
rect 3979 817 3985 823
rect 85 765 91 771
rect 2019 765 2025 771
rect 2019 737 2025 743
rect 3967 737 3973 743
rect 97 689 103 695
rect 2031 689 2037 695
rect 2031 653 2037 659
rect 3979 653 3985 659
rect 85 613 91 619
rect 2019 613 2025 619
rect 2019 573 2025 579
rect 3967 573 3973 579
rect 97 517 103 523
rect 2031 517 2037 523
rect 2031 497 2037 503
rect 3979 497 3985 503
rect 85 429 91 435
rect 2019 429 2025 435
rect 2019 421 2025 427
rect 3967 421 3973 427
rect 97 349 103 355
rect 2031 349 2037 355
rect 2031 341 2037 347
rect 3979 341 3985 347
rect 85 265 91 271
rect 2019 265 2025 271
rect 97 161 103 167
rect 2031 161 2037 167
rect 85 85 91 91
rect 2019 85 2025 91
<< m5 >>
rect 84 3955 92 4032
rect 84 3949 85 3955
rect 91 3949 92 3955
rect 84 3799 92 3949
rect 84 3793 85 3799
rect 91 3793 92 3799
rect 84 3631 92 3793
rect 84 3625 85 3631
rect 91 3625 92 3631
rect 84 3459 92 3625
rect 84 3453 85 3459
rect 91 3453 92 3459
rect 84 3307 92 3453
rect 84 3301 85 3307
rect 91 3301 92 3307
rect 84 3151 92 3301
rect 84 3145 85 3151
rect 91 3145 92 3151
rect 84 2987 92 3145
rect 84 2981 85 2987
rect 91 2981 92 2987
rect 84 2823 92 2981
rect 84 2817 85 2823
rect 91 2817 92 2823
rect 84 2663 92 2817
rect 84 2657 85 2663
rect 91 2657 92 2663
rect 84 2495 92 2657
rect 84 2489 85 2495
rect 91 2489 92 2495
rect 84 2327 92 2489
rect 84 2321 85 2327
rect 91 2321 92 2327
rect 84 2171 92 2321
rect 84 2165 85 2171
rect 91 2165 92 2171
rect 84 2015 92 2165
rect 84 2009 85 2015
rect 91 2009 92 2015
rect 84 1863 92 2009
rect 84 1857 85 1863
rect 91 1857 92 1863
rect 84 1707 92 1857
rect 84 1701 85 1707
rect 91 1701 92 1707
rect 84 1551 92 1701
rect 84 1545 85 1551
rect 91 1545 92 1551
rect 84 1399 92 1545
rect 84 1393 85 1399
rect 91 1393 92 1399
rect 84 1239 92 1393
rect 84 1233 85 1239
rect 91 1233 92 1239
rect 84 1075 92 1233
rect 84 1069 85 1075
rect 91 1069 92 1075
rect 84 923 92 1069
rect 84 917 85 923
rect 91 917 92 923
rect 84 771 92 917
rect 84 765 85 771
rect 91 765 92 771
rect 84 619 92 765
rect 84 613 85 619
rect 91 613 92 619
rect 84 435 92 613
rect 84 429 85 435
rect 91 429 92 435
rect 84 271 92 429
rect 84 265 85 271
rect 91 265 92 271
rect 84 91 92 265
rect 84 85 85 91
rect 91 85 92 91
rect 84 72 92 85
rect 96 4031 104 4032
rect 96 4025 97 4031
rect 103 4025 104 4031
rect 96 3879 104 4025
rect 96 3873 97 3879
rect 103 3873 104 3879
rect 96 3715 104 3873
rect 96 3709 97 3715
rect 103 3709 104 3715
rect 96 3543 104 3709
rect 96 3537 97 3543
rect 103 3537 104 3543
rect 96 3383 104 3537
rect 96 3377 97 3383
rect 103 3377 104 3383
rect 96 3231 104 3377
rect 96 3225 97 3231
rect 103 3225 104 3231
rect 96 3067 104 3225
rect 96 3061 97 3067
rect 103 3061 104 3067
rect 96 2903 104 3061
rect 96 2897 97 2903
rect 103 2897 104 2903
rect 96 2743 104 2897
rect 96 2737 97 2743
rect 103 2737 104 2743
rect 96 2587 104 2737
rect 96 2581 97 2587
rect 103 2581 104 2587
rect 96 2403 104 2581
rect 96 2397 97 2403
rect 103 2397 104 2403
rect 96 2247 104 2397
rect 96 2241 97 2247
rect 103 2241 104 2247
rect 96 2095 104 2241
rect 96 2089 97 2095
rect 103 2089 104 2095
rect 96 1939 104 2089
rect 96 1933 97 1939
rect 103 1933 104 1939
rect 96 1783 104 1933
rect 96 1777 97 1783
rect 103 1777 104 1783
rect 96 1631 104 1777
rect 96 1625 97 1631
rect 103 1625 104 1631
rect 96 1475 104 1625
rect 96 1469 97 1475
rect 103 1469 104 1475
rect 96 1315 104 1469
rect 96 1309 97 1315
rect 103 1309 104 1315
rect 96 1159 104 1309
rect 96 1153 97 1159
rect 103 1153 104 1159
rect 96 999 104 1153
rect 96 993 97 999
rect 103 993 104 999
rect 96 847 104 993
rect 96 841 97 847
rect 103 841 104 847
rect 96 695 104 841
rect 96 689 97 695
rect 103 689 104 695
rect 96 523 104 689
rect 96 517 97 523
rect 103 517 104 523
rect 96 355 104 517
rect 96 349 97 355
rect 103 349 104 355
rect 96 167 104 349
rect 96 161 97 167
rect 103 161 104 167
rect 96 72 104 161
rect 2018 4019 2026 4032
rect 2018 4013 2019 4019
rect 2025 4013 2026 4019
rect 2018 3955 2026 4013
rect 2018 3949 2019 3955
rect 2025 3949 2026 3955
rect 2018 3859 2026 3949
rect 2018 3853 2019 3859
rect 2025 3853 2026 3859
rect 2018 3799 2026 3853
rect 2018 3793 2019 3799
rect 2025 3793 2026 3799
rect 2018 3703 2026 3793
rect 2018 3697 2019 3703
rect 2025 3697 2026 3703
rect 2018 3631 2026 3697
rect 2018 3625 2019 3631
rect 2025 3625 2026 3631
rect 2018 3553 2026 3625
rect 2018 3547 2019 3553
rect 2025 3547 2026 3553
rect 2018 3459 2026 3547
rect 2018 3453 2019 3459
rect 2025 3453 2026 3459
rect 2018 3371 2026 3453
rect 2018 3365 2019 3371
rect 2025 3365 2026 3371
rect 2018 3307 2026 3365
rect 2018 3301 2019 3307
rect 2025 3301 2026 3307
rect 2018 3211 2026 3301
rect 2018 3205 2019 3211
rect 2025 3205 2026 3211
rect 2018 3151 2026 3205
rect 2018 3145 2019 3151
rect 2025 3145 2026 3151
rect 2018 3047 2026 3145
rect 2018 3041 2019 3047
rect 2025 3041 2026 3047
rect 2018 2987 2026 3041
rect 2018 2981 2019 2987
rect 2025 2981 2026 2987
rect 2018 2891 2026 2981
rect 2018 2885 2019 2891
rect 2025 2885 2026 2891
rect 2018 2823 2026 2885
rect 2018 2817 2019 2823
rect 2025 2817 2026 2823
rect 2018 2731 2026 2817
rect 2018 2725 2019 2731
rect 2025 2725 2026 2731
rect 2018 2663 2026 2725
rect 2018 2657 2019 2663
rect 2025 2657 2026 2663
rect 2018 2567 2026 2657
rect 2018 2561 2019 2567
rect 2025 2561 2026 2567
rect 2018 2495 2026 2561
rect 2018 2489 2019 2495
rect 2025 2489 2026 2495
rect 2018 2413 2026 2489
rect 2018 2407 2019 2413
rect 2025 2407 2026 2413
rect 2018 2327 2026 2407
rect 2018 2321 2019 2327
rect 2025 2321 2026 2327
rect 2018 2231 2026 2321
rect 2018 2225 2019 2231
rect 2025 2225 2026 2231
rect 2018 2171 2026 2225
rect 2018 2165 2019 2171
rect 2025 2165 2026 2171
rect 2018 2051 2026 2165
rect 2018 2045 2019 2051
rect 2025 2045 2026 2051
rect 2018 2015 2026 2045
rect 2018 2009 2019 2015
rect 2025 2009 2026 2015
rect 2018 1883 2026 2009
rect 2018 1877 2019 1883
rect 2025 1877 2026 1883
rect 2018 1863 2026 1877
rect 2018 1857 2019 1863
rect 2025 1857 2026 1863
rect 2018 1723 2026 1857
rect 2018 1717 2019 1723
rect 2025 1717 2026 1723
rect 2018 1707 2026 1717
rect 2018 1701 2019 1707
rect 2025 1701 2026 1707
rect 2018 1567 2026 1701
rect 2018 1561 2019 1567
rect 2025 1561 2026 1567
rect 2018 1551 2026 1561
rect 2018 1545 2019 1551
rect 2025 1545 2026 1551
rect 2018 1399 2026 1545
rect 2018 1393 2019 1399
rect 2025 1393 2026 1399
rect 2018 1239 2026 1393
rect 2018 1233 2019 1239
rect 2025 1233 2026 1239
rect 2018 1227 2026 1233
rect 2018 1221 2019 1227
rect 2025 1221 2026 1227
rect 2018 1075 2026 1221
rect 2018 1069 2019 1075
rect 2025 1069 2026 1075
rect 2018 1063 2026 1069
rect 2018 1057 2019 1063
rect 2025 1057 2026 1063
rect 2018 923 2026 1057
rect 2018 917 2019 923
rect 2025 917 2026 923
rect 2018 899 2026 917
rect 2018 893 2019 899
rect 2025 893 2026 899
rect 2018 771 2026 893
rect 2018 765 2019 771
rect 2025 765 2026 771
rect 2018 743 2026 765
rect 2018 737 2019 743
rect 2025 737 2026 743
rect 2018 619 2026 737
rect 2018 613 2019 619
rect 2025 613 2026 619
rect 2018 579 2026 613
rect 2018 573 2019 579
rect 2025 573 2026 579
rect 2018 435 2026 573
rect 2018 429 2019 435
rect 2025 429 2026 435
rect 2018 427 2026 429
rect 2018 421 2019 427
rect 2025 421 2026 427
rect 2018 271 2026 421
rect 2018 265 2019 271
rect 2025 265 2026 271
rect 2018 91 2026 265
rect 2018 85 2019 91
rect 2025 85 2026 91
rect 2018 72 2026 85
rect 2030 4031 2038 4032
rect 2030 4025 2031 4031
rect 2037 4025 2038 4031
rect 2030 3943 2038 4025
rect 2030 3937 2031 3943
rect 2037 3937 2038 3943
rect 2030 3879 2038 3937
rect 2030 3873 2031 3879
rect 2037 3873 2038 3879
rect 2030 3783 2038 3873
rect 2030 3777 2031 3783
rect 2037 3777 2038 3783
rect 2030 3715 2038 3777
rect 2030 3709 2031 3715
rect 2037 3709 2038 3715
rect 2030 3619 2038 3709
rect 2030 3613 2031 3619
rect 2037 3613 2038 3619
rect 2030 3543 2038 3613
rect 2030 3537 2031 3543
rect 2037 3537 2038 3543
rect 2030 3463 2038 3537
rect 2030 3457 2031 3463
rect 2037 3457 2038 3463
rect 2030 3383 2038 3457
rect 2030 3377 2031 3383
rect 2037 3377 2038 3383
rect 2030 3287 2038 3377
rect 2030 3281 2031 3287
rect 2037 3281 2038 3287
rect 2030 3231 2038 3281
rect 2030 3225 2031 3231
rect 2037 3225 2038 3231
rect 2030 3123 2038 3225
rect 2030 3117 2031 3123
rect 2037 3117 2038 3123
rect 2030 3067 2038 3117
rect 2030 3061 2031 3067
rect 2037 3061 2038 3067
rect 2030 2967 2038 3061
rect 2030 2961 2031 2967
rect 2037 2961 2038 2967
rect 2030 2903 2038 2961
rect 2030 2897 2031 2903
rect 2037 2897 2038 2903
rect 2030 2811 2038 2897
rect 2030 2805 2031 2811
rect 2037 2805 2038 2811
rect 2030 2743 2038 2805
rect 2030 2737 2031 2743
rect 2037 2737 2038 2743
rect 2030 2647 2038 2737
rect 2030 2641 2031 2647
rect 2037 2641 2038 2647
rect 2030 2587 2038 2641
rect 2030 2581 2031 2587
rect 2037 2581 2038 2587
rect 2030 2487 2038 2581
rect 2030 2481 2031 2487
rect 2037 2481 2038 2487
rect 2030 2403 2038 2481
rect 2030 2397 2031 2403
rect 2037 2397 2038 2403
rect 2030 2307 2038 2397
rect 2030 2301 2031 2307
rect 2037 2301 2038 2307
rect 2030 2247 2038 2301
rect 2030 2241 2031 2247
rect 2037 2241 2038 2247
rect 2030 2135 2038 2241
rect 2030 2129 2031 2135
rect 2037 2129 2038 2135
rect 2030 2095 2038 2129
rect 2030 2089 2031 2095
rect 2037 2089 2038 2095
rect 2030 1971 2038 2089
rect 2030 1965 2031 1971
rect 2037 1965 2038 1971
rect 2030 1939 2038 1965
rect 2030 1933 2031 1939
rect 2037 1933 2038 1939
rect 2030 1803 2038 1933
rect 2030 1797 2031 1803
rect 2037 1797 2038 1803
rect 2030 1783 2038 1797
rect 2030 1777 2031 1783
rect 2037 1777 2038 1783
rect 2030 1647 2038 1777
rect 2030 1641 2031 1647
rect 2037 1641 2038 1647
rect 2030 1631 2038 1641
rect 2030 1625 2031 1631
rect 2037 1625 2038 1631
rect 2030 1491 2038 1625
rect 2030 1485 2031 1491
rect 2037 1485 2038 1491
rect 2030 1475 2038 1485
rect 2030 1469 2031 1475
rect 2037 1469 2038 1475
rect 2030 1315 2038 1469
rect 2030 1309 2031 1315
rect 2037 1309 2038 1315
rect 2030 1159 2038 1309
rect 2030 1153 2031 1159
rect 2037 1153 2038 1159
rect 2030 1143 2038 1153
rect 2030 1137 2031 1143
rect 2037 1137 2038 1143
rect 2030 999 2038 1137
rect 2030 993 2031 999
rect 2037 993 2038 999
rect 2030 987 2038 993
rect 2030 981 2031 987
rect 2037 981 2038 987
rect 2030 847 2038 981
rect 2030 841 2031 847
rect 2037 841 2038 847
rect 2030 823 2038 841
rect 2030 817 2031 823
rect 2037 817 2038 823
rect 2030 695 2038 817
rect 2030 689 2031 695
rect 2037 689 2038 695
rect 2030 659 2038 689
rect 2030 653 2031 659
rect 2037 653 2038 659
rect 2030 523 2038 653
rect 2030 517 2031 523
rect 2037 517 2038 523
rect 2030 503 2038 517
rect 2030 497 2031 503
rect 2037 497 2038 503
rect 2030 355 2038 497
rect 2030 349 2031 355
rect 2037 349 2038 355
rect 2030 347 2038 349
rect 2030 341 2031 347
rect 2037 341 2038 347
rect 2030 167 2038 341
rect 2030 161 2031 167
rect 2037 161 2038 167
rect 2030 72 2038 161
rect 3966 4019 3974 4032
rect 3966 4013 3967 4019
rect 3973 4013 3974 4019
rect 3966 3859 3974 4013
rect 3966 3853 3967 3859
rect 3973 3853 3974 3859
rect 3966 3703 3974 3853
rect 3966 3697 3967 3703
rect 3973 3697 3974 3703
rect 3966 3543 3974 3697
rect 3966 3537 3967 3543
rect 3973 3537 3974 3543
rect 3966 3371 3974 3537
rect 3966 3365 3967 3371
rect 3973 3365 3974 3371
rect 3966 3211 3974 3365
rect 3966 3205 3967 3211
rect 3973 3205 3974 3211
rect 3966 3047 3974 3205
rect 3966 3041 3967 3047
rect 3973 3041 3974 3047
rect 3966 2891 3974 3041
rect 3966 2885 3967 2891
rect 3973 2885 3974 2891
rect 3966 2731 3974 2885
rect 3966 2725 3967 2731
rect 3973 2725 3974 2731
rect 3966 2567 3974 2725
rect 3966 2561 3967 2567
rect 3973 2561 3974 2567
rect 3966 2399 3974 2561
rect 3966 2393 3967 2399
rect 3973 2393 3974 2399
rect 3966 2231 3974 2393
rect 3966 2225 3967 2231
rect 3973 2225 3974 2231
rect 3966 2051 3974 2225
rect 3966 2045 3967 2051
rect 3973 2045 3974 2051
rect 3966 1883 3974 2045
rect 3966 1877 3967 1883
rect 3973 1877 3974 1883
rect 3966 1723 3974 1877
rect 3966 1717 3967 1723
rect 3973 1717 3974 1723
rect 3966 1567 3974 1717
rect 3966 1561 3967 1567
rect 3973 1561 3974 1567
rect 3966 1227 3974 1561
rect 3966 1221 3967 1227
rect 3973 1221 3974 1227
rect 3966 1063 3974 1221
rect 3966 1057 3967 1063
rect 3973 1057 3974 1063
rect 3966 899 3974 1057
rect 3966 893 3967 899
rect 3973 893 3974 899
rect 3966 743 3974 893
rect 3966 737 3967 743
rect 3973 737 3974 743
rect 3966 579 3974 737
rect 3966 573 3967 579
rect 3973 573 3974 579
rect 3966 427 3974 573
rect 3966 421 3967 427
rect 3973 421 3974 427
rect 3966 72 3974 421
rect 3978 3943 3986 4032
rect 3978 3937 3979 3943
rect 3985 3937 3986 3943
rect 3978 3783 3986 3937
rect 3978 3777 3979 3783
rect 3985 3777 3986 3783
rect 3978 3619 3986 3777
rect 3978 3613 3979 3619
rect 3985 3613 3986 3619
rect 3978 3463 3986 3613
rect 3978 3457 3979 3463
rect 3985 3457 3986 3463
rect 3978 3287 3986 3457
rect 3978 3281 3979 3287
rect 3985 3281 3986 3287
rect 3978 3123 3986 3281
rect 3978 3117 3979 3123
rect 3985 3117 3986 3123
rect 3978 2967 3986 3117
rect 3978 2961 3979 2967
rect 3985 2961 3986 2967
rect 3978 2811 3986 2961
rect 3978 2805 3979 2811
rect 3985 2805 3986 2811
rect 3978 2647 3986 2805
rect 3978 2641 3979 2647
rect 3985 2641 3986 2647
rect 3978 2487 3986 2641
rect 3978 2481 3979 2487
rect 3985 2481 3986 2487
rect 3978 2307 3986 2481
rect 3978 2301 3979 2307
rect 3985 2301 3986 2307
rect 3978 2135 3986 2301
rect 3978 2129 3979 2135
rect 3985 2129 3986 2135
rect 3978 1971 3986 2129
rect 3978 1965 3979 1971
rect 3985 1965 3986 1971
rect 3978 1803 3986 1965
rect 3978 1797 3979 1803
rect 3985 1797 3986 1803
rect 3978 1647 3986 1797
rect 3978 1641 3979 1647
rect 3985 1641 3986 1647
rect 3978 1491 3986 1641
rect 3978 1485 3979 1491
rect 3985 1485 3986 1491
rect 3978 1143 3986 1485
rect 3978 1137 3979 1143
rect 3985 1137 3986 1143
rect 3978 987 3986 1137
rect 3978 981 3979 987
rect 3985 981 3986 987
rect 3978 823 3986 981
rect 3978 817 3979 823
rect 3985 817 3986 823
rect 3978 659 3986 817
rect 3978 653 3979 659
rect 3985 653 3986 659
rect 3978 503 3986 653
rect 3978 497 3979 503
rect 3985 497 3986 503
rect 3978 347 3986 497
rect 3978 341 3979 347
rect 3985 341 3986 347
rect 3978 72 3986 341
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__193
timestamp 1731220340
transform 1 0 3936 0 -1 3988
box 7 3 12 24
use welltap_svt  __well_tap__192
timestamp 1731220340
transform 1 0 2040 0 -1 3988
box 7 3 12 24
use welltap_svt  __well_tap__191
timestamp 1731220340
transform 1 0 3936 0 1 3892
box 7 3 12 24
use welltap_svt  __well_tap__190
timestamp 1731220340
transform 1 0 2040 0 1 3892
box 7 3 12 24
use welltap_svt  __well_tap__189
timestamp 1731220340
transform 1 0 3936 0 -1 3828
box 7 3 12 24
use welltap_svt  __well_tap__188
timestamp 1731220340
transform 1 0 2040 0 -1 3828
box 7 3 12 24
use welltap_svt  __well_tap__187
timestamp 1731220340
transform 1 0 3936 0 1 3732
box 7 3 12 24
use welltap_svt  __well_tap__186
timestamp 1731220340
transform 1 0 2040 0 1 3732
box 7 3 12 24
use welltap_svt  __well_tap__185
timestamp 1731220340
transform 1 0 3936 0 -1 3672
box 7 3 12 24
use welltap_svt  __well_tap__184
timestamp 1731220340
transform 1 0 2040 0 -1 3672
box 7 3 12 24
use welltap_svt  __well_tap__183
timestamp 1731220340
transform 1 0 3936 0 1 3568
box 7 3 12 24
use welltap_svt  __well_tap__182
timestamp 1731220340
transform 1 0 2040 0 1 3568
box 7 3 12 24
use welltap_svt  __well_tap__181
timestamp 1731220340
transform 1 0 3936 0 -1 3512
box 7 3 12 24
use welltap_svt  __well_tap__180
timestamp 1731220340
transform 1 0 2040 0 -1 3512
box 7 3 12 24
use welltap_svt  __well_tap__179
timestamp 1731220340
transform 1 0 3936 0 1 3412
box 7 3 12 24
use welltap_svt  __well_tap__178
timestamp 1731220340
transform 1 0 2040 0 1 3412
box 7 3 12 24
use welltap_svt  __well_tap__177
timestamp 1731220340
transform 1 0 3936 0 -1 3340
box 7 3 12 24
use welltap_svt  __well_tap__176
timestamp 1731220340
transform 1 0 2040 0 -1 3340
box 7 3 12 24
use welltap_svt  __well_tap__175
timestamp 1731220340
transform 1 0 3936 0 1 3236
box 7 3 12 24
use welltap_svt  __well_tap__174
timestamp 1731220340
transform 1 0 2040 0 1 3236
box 7 3 12 24
use welltap_svt  __well_tap__173
timestamp 1731220340
transform 1 0 3936 0 -1 3180
box 7 3 12 24
use welltap_svt  __well_tap__172
timestamp 1731220340
transform 1 0 2040 0 -1 3180
box 7 3 12 24
use welltap_svt  __well_tap__171
timestamp 1731220340
transform 1 0 3936 0 1 3072
box 7 3 12 24
use welltap_svt  __well_tap__170
timestamp 1731220340
transform 1 0 2040 0 1 3072
box 7 3 12 24
use welltap_svt  __well_tap__169
timestamp 1731220340
transform 1 0 3936 0 -1 3016
box 7 3 12 24
use welltap_svt  __well_tap__168
timestamp 1731220340
transform 1 0 2040 0 -1 3016
box 7 3 12 24
use welltap_svt  __well_tap__167
timestamp 1731220340
transform 1 0 3936 0 1 2916
box 7 3 12 24
use welltap_svt  __well_tap__166
timestamp 1731220340
transform 1 0 2040 0 1 2916
box 7 3 12 24
use welltap_svt  __well_tap__165
timestamp 1731220340
transform 1 0 3936 0 -1 2860
box 7 3 12 24
use welltap_svt  __well_tap__164
timestamp 1731220340
transform 1 0 2040 0 -1 2860
box 7 3 12 24
use welltap_svt  __well_tap__163
timestamp 1731220340
transform 1 0 3936 0 1 2760
box 7 3 12 24
use welltap_svt  __well_tap__162
timestamp 1731220340
transform 1 0 2040 0 1 2760
box 7 3 12 24
use welltap_svt  __well_tap__161
timestamp 1731220340
transform 1 0 3936 0 -1 2700
box 7 3 12 24
use welltap_svt  __well_tap__160
timestamp 1731220340
transform 1 0 2040 0 -1 2700
box 7 3 12 24
use welltap_svt  __well_tap__159
timestamp 1731220340
transform 1 0 3936 0 1 2596
box 7 3 12 24
use welltap_svt  __well_tap__158
timestamp 1731220340
transform 1 0 2040 0 1 2596
box 7 3 12 24
use welltap_svt  __well_tap__157
timestamp 1731220340
transform 1 0 3936 0 -1 2536
box 7 3 12 24
use welltap_svt  __well_tap__156
timestamp 1731220340
transform 1 0 2040 0 -1 2536
box 7 3 12 24
use welltap_svt  __well_tap__155
timestamp 1731220340
transform 1 0 3936 0 1 2436
box 7 3 12 24
use welltap_svt  __well_tap__154
timestamp 1731220340
transform 1 0 2040 0 1 2436
box 7 3 12 24
use welltap_svt  __well_tap__153
timestamp 1731220340
transform 1 0 3936 0 -1 2368
box 7 3 12 24
use welltap_svt  __well_tap__152
timestamp 1731220340
transform 1 0 2040 0 -1 2368
box 7 3 12 24
use welltap_svt  __well_tap__151
timestamp 1731220340
transform 1 0 3936 0 1 2256
box 7 3 12 24
use welltap_svt  __well_tap__150
timestamp 1731220340
transform 1 0 2040 0 1 2256
box 7 3 12 24
use welltap_svt  __well_tap__149
timestamp 1731220340
transform 1 0 3936 0 -1 2200
box 7 3 12 24
use welltap_svt  __well_tap__148
timestamp 1731220340
transform 1 0 2040 0 -1 2200
box 7 3 12 24
use welltap_svt  __well_tap__147
timestamp 1731220340
transform 1 0 3936 0 1 2084
box 7 3 12 24
use welltap_svt  __well_tap__146
timestamp 1731220340
transform 1 0 2040 0 1 2084
box 7 3 12 24
use welltap_svt  __well_tap__145
timestamp 1731220340
transform 1 0 3936 0 -1 2020
box 7 3 12 24
use welltap_svt  __well_tap__144
timestamp 1731220340
transform 1 0 2040 0 -1 2020
box 7 3 12 24
use welltap_svt  __well_tap__143
timestamp 1731220340
transform 1 0 3936 0 1 1920
box 7 3 12 24
use welltap_svt  __well_tap__142
timestamp 1731220340
transform 1 0 2040 0 1 1920
box 7 3 12 24
use welltap_svt  __well_tap__141
timestamp 1731220340
transform 1 0 3936 0 -1 1852
box 7 3 12 24
use welltap_svt  __well_tap__140
timestamp 1731220340
transform 1 0 2040 0 -1 1852
box 7 3 12 24
use welltap_svt  __well_tap__139
timestamp 1731220340
transform 1 0 3936 0 1 1752
box 7 3 12 24
use welltap_svt  __well_tap__138
timestamp 1731220340
transform 1 0 2040 0 1 1752
box 7 3 12 24
use welltap_svt  __well_tap__137
timestamp 1731220340
transform 1 0 3936 0 -1 1692
box 7 3 12 24
use welltap_svt  __well_tap__136
timestamp 1731220340
transform 1 0 2040 0 -1 1692
box 7 3 12 24
use welltap_svt  __well_tap__135
timestamp 1731220340
transform 1 0 3936 0 1 1596
box 7 3 12 24
use welltap_svt  __well_tap__134
timestamp 1731220340
transform 1 0 2040 0 1 1596
box 7 3 12 24
use welltap_svt  __well_tap__133
timestamp 1731220340
transform 1 0 3936 0 -1 1536
box 7 3 12 24
use welltap_svt  __well_tap__132
timestamp 1731220340
transform 1 0 2040 0 -1 1536
box 7 3 12 24
use welltap_svt  __well_tap__131
timestamp 1731220340
transform 1 0 3936 0 1 1440
box 7 3 12 24
use welltap_svt  __well_tap__130
timestamp 1731220340
transform 1 0 2040 0 1 1440
box 7 3 12 24
use welltap_svt  __well_tap__129
timestamp 1731220340
transform 1 0 3936 0 -1 1364
box 7 3 12 24
use welltap_svt  __well_tap__128
timestamp 1731220340
transform 1 0 2040 0 -1 1364
box 7 3 12 24
use welltap_svt  __well_tap__127
timestamp 1731220340
transform 1 0 3936 0 1 1260
box 7 3 12 24
use welltap_svt  __well_tap__126
timestamp 1731220340
transform 1 0 2040 0 1 1260
box 7 3 12 24
use welltap_svt  __well_tap__125
timestamp 1731220340
transform 1 0 3936 0 -1 1196
box 7 3 12 24
use welltap_svt  __well_tap__124
timestamp 1731220340
transform 1 0 2040 0 -1 1196
box 7 3 12 24
use welltap_svt  __well_tap__123
timestamp 1731220340
transform 1 0 3936 0 1 1092
box 7 3 12 24
use welltap_svt  __well_tap__122
timestamp 1731220340
transform 1 0 2040 0 1 1092
box 7 3 12 24
use welltap_svt  __well_tap__121
timestamp 1731220340
transform 1 0 3936 0 -1 1032
box 7 3 12 24
use welltap_svt  __well_tap__120
timestamp 1731220340
transform 1 0 2040 0 -1 1032
box 7 3 12 24
use welltap_svt  __well_tap__119
timestamp 1731220340
transform 1 0 3936 0 1 936
box 7 3 12 24
use welltap_svt  __well_tap__118
timestamp 1731220340
transform 1 0 2040 0 1 936
box 7 3 12 24
use welltap_svt  __well_tap__117
timestamp 1731220340
transform 1 0 3936 0 -1 868
box 7 3 12 24
use welltap_svt  __well_tap__116
timestamp 1731220340
transform 1 0 2040 0 -1 868
box 7 3 12 24
use welltap_svt  __well_tap__115
timestamp 1731220340
transform 1 0 3936 0 1 772
box 7 3 12 24
use welltap_svt  __well_tap__114
timestamp 1731220340
transform 1 0 2040 0 1 772
box 7 3 12 24
use welltap_svt  __well_tap__113
timestamp 1731220340
transform 1 0 3936 0 -1 712
box 7 3 12 24
use welltap_svt  __well_tap__112
timestamp 1731220340
transform 1 0 2040 0 -1 712
box 7 3 12 24
use welltap_svt  __well_tap__111
timestamp 1731220340
transform 1 0 3936 0 1 608
box 7 3 12 24
use welltap_svt  __well_tap__110
timestamp 1731220340
transform 1 0 2040 0 1 608
box 7 3 12 24
use welltap_svt  __well_tap__109
timestamp 1731220340
transform 1 0 3936 0 -1 548
box 7 3 12 24
use welltap_svt  __well_tap__108
timestamp 1731220340
transform 1 0 2040 0 -1 548
box 7 3 12 24
use welltap_svt  __well_tap__107
timestamp 1731220340
transform 1 0 3936 0 1 452
box 7 3 12 24
use welltap_svt  __well_tap__106
timestamp 1731220340
transform 1 0 2040 0 1 452
box 7 3 12 24
use welltap_svt  __well_tap__105
timestamp 1731220340
transform 1 0 3936 0 -1 396
box 7 3 12 24
use welltap_svt  __well_tap__104
timestamp 1731220340
transform 1 0 2040 0 -1 396
box 7 3 12 24
use welltap_svt  __well_tap__103
timestamp 1731220340
transform 1 0 3936 0 1 296
box 7 3 12 24
use welltap_svt  __well_tap__102
timestamp 1731220340
transform 1 0 2040 0 1 296
box 7 3 12 24
use welltap_svt  __well_tap__101
timestamp 1731220340
transform 1 0 3936 0 -1 240
box 7 3 12 24
use welltap_svt  __well_tap__100
timestamp 1731220340
transform 1 0 2040 0 -1 240
box 7 3 12 24
use welltap_svt  __well_tap__99
timestamp 1731220340
transform 1 0 3936 0 1 120
box 7 3 12 24
use welltap_svt  __well_tap__98
timestamp 1731220340
transform 1 0 2040 0 1 120
box 7 3 12 24
use welltap_svt  __well_tap__97
timestamp 1731220340
transform 1 0 2000 0 1 3980
box 7 3 12 24
use welltap_svt  __well_tap__96
timestamp 1731220340
transform 1 0 104 0 1 3980
box 7 3 12 24
use welltap_svt  __well_tap__95
timestamp 1731220340
transform 1 0 2000 0 -1 3924
box 7 3 12 24
use welltap_svt  __well_tap__94
timestamp 1731220340
transform 1 0 104 0 -1 3924
box 7 3 12 24
use welltap_svt  __well_tap__93
timestamp 1731220340
transform 1 0 2000 0 1 3828
box 7 3 12 24
use welltap_svt  __well_tap__92
timestamp 1731220340
transform 1 0 104 0 1 3828
box 7 3 12 24
use welltap_svt  __well_tap__91
timestamp 1731220340
transform 1 0 2000 0 -1 3768
box 7 3 12 24
use welltap_svt  __well_tap__90
timestamp 1731220340
transform 1 0 104 0 -1 3768
box 7 3 12 24
use welltap_svt  __well_tap__89
timestamp 1731220340
transform 1 0 2000 0 1 3664
box 7 3 12 24
use welltap_svt  __well_tap__88
timestamp 1731220340
transform 1 0 104 0 1 3664
box 7 3 12 24
use welltap_svt  __well_tap__87
timestamp 1731220340
transform 1 0 2000 0 -1 3600
box 7 3 12 24
use welltap_svt  __well_tap__86
timestamp 1731220340
transform 1 0 104 0 -1 3600
box 7 3 12 24
use welltap_svt  __well_tap__85
timestamp 1731220340
transform 1 0 2000 0 1 3492
box 7 3 12 24
use welltap_svt  __well_tap__84
timestamp 1731220340
transform 1 0 104 0 1 3492
box 7 3 12 24
use welltap_svt  __well_tap__83
timestamp 1731220340
transform 1 0 2000 0 -1 3428
box 7 3 12 24
use welltap_svt  __well_tap__82
timestamp 1731220340
transform 1 0 104 0 -1 3428
box 7 3 12 24
use welltap_svt  __well_tap__81
timestamp 1731220340
transform 1 0 2000 0 1 3332
box 7 3 12 24
use welltap_svt  __well_tap__80
timestamp 1731220340
transform 1 0 104 0 1 3332
box 7 3 12 24
use welltap_svt  __well_tap__79
timestamp 1731220340
transform 1 0 2000 0 -1 3276
box 7 3 12 24
use welltap_svt  __well_tap__78
timestamp 1731220340
transform 1 0 104 0 -1 3276
box 7 3 12 24
use welltap_svt  __well_tap__77
timestamp 1731220340
transform 1 0 2000 0 1 3180
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220340
transform 1 0 104 0 1 3180
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220340
transform 1 0 2000 0 -1 3120
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220340
transform 1 0 104 0 -1 3120
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220340
transform 1 0 2000 0 1 3016
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220340
transform 1 0 104 0 1 3016
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220340
transform 1 0 2000 0 -1 2956
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220340
transform 1 0 104 0 -1 2956
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220340
transform 1 0 2000 0 1 2852
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220340
transform 1 0 104 0 1 2852
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220340
transform 1 0 2000 0 -1 2792
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220340
transform 1 0 104 0 -1 2792
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220340
transform 1 0 2000 0 1 2692
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220340
transform 1 0 104 0 1 2692
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220340
transform 1 0 2000 0 -1 2632
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220340
transform 1 0 104 0 -1 2632
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220340
transform 1 0 2000 0 1 2536
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220340
transform 1 0 104 0 1 2536
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220340
transform 1 0 2000 0 -1 2464
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220340
transform 1 0 104 0 -1 2464
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220340
transform 1 0 2000 0 1 2352
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220340
transform 1 0 104 0 1 2352
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220340
transform 1 0 2000 0 -1 2296
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220340
transform 1 0 104 0 -1 2296
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220340
transform 1 0 2000 0 1 2196
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220340
transform 1 0 104 0 1 2196
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220340
transform 1 0 2000 0 -1 2140
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220340
transform 1 0 104 0 -1 2140
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220340
transform 1 0 2000 0 1 2044
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220340
transform 1 0 104 0 1 2044
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220340
transform 1 0 2000 0 -1 1984
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220340
transform 1 0 104 0 -1 1984
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220340
transform 1 0 2000 0 1 1888
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220340
transform 1 0 104 0 1 1888
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220340
transform 1 0 2000 0 -1 1832
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220340
transform 1 0 104 0 -1 1832
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220340
transform 1 0 2000 0 1 1732
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220340
transform 1 0 104 0 1 1732
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220340
transform 1 0 2000 0 -1 1676
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220340
transform 1 0 104 0 -1 1676
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220340
transform 1 0 2000 0 1 1580
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220340
transform 1 0 104 0 1 1580
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220340
transform 1 0 2000 0 -1 1520
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220340
transform 1 0 104 0 -1 1520
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220340
transform 1 0 2000 0 1 1424
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220340
transform 1 0 104 0 1 1424
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220340
transform 1 0 2000 0 -1 1368
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220340
transform 1 0 104 0 -1 1368
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220340
transform 1 0 2000 0 1 1264
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220340
transform 1 0 104 0 1 1264
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220340
transform 1 0 2000 0 -1 1208
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220340
transform 1 0 104 0 -1 1208
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220340
transform 1 0 2000 0 1 1108
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220340
transform 1 0 104 0 1 1108
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220340
transform 1 0 2000 0 -1 1044
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220340
transform 1 0 104 0 -1 1044
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220340
transform 1 0 2000 0 1 948
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220340
transform 1 0 104 0 1 948
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220340
transform 1 0 2000 0 -1 892
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220340
transform 1 0 104 0 -1 892
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220340
transform 1 0 2000 0 1 796
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220340
transform 1 0 104 0 1 796
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220340
transform 1 0 2000 0 -1 740
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220340
transform 1 0 104 0 -1 740
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220340
transform 1 0 2000 0 1 644
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220340
transform 1 0 104 0 1 644
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220340
transform 1 0 2000 0 -1 588
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220340
transform 1 0 104 0 -1 588
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220340
transform 1 0 2000 0 1 472
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220340
transform 1 0 104 0 1 472
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220340
transform 1 0 2000 0 -1 404
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220340
transform 1 0 104 0 -1 404
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220340
transform 1 0 2000 0 1 304
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220340
transform 1 0 104 0 1 304
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220340
transform 1 0 2000 0 -1 240
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220340
transform 1 0 104 0 -1 240
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220340
transform 1 0 2000 0 1 116
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220340
transform 1 0 104 0 1 116
box 7 3 12 24
use _0_0cell_0_0gcelem3x0  tst_5999_6
timestamp 1731220340
transform 1 0 3680 0 -1 3540
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5998_6
timestamp 1731220340
transform 1 0 3832 0 -1 3540
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5997_6
timestamp 1731220340
transform 1 0 3832 0 -1 3368
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5996_6
timestamp 1731220340
transform 1 0 3832 0 -1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5995_6
timestamp 1731220340
transform 1 0 3832 0 -1 3044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5994_6
timestamp 1731220340
transform 1 0 3832 0 -1 2888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5993_6
timestamp 1731220340
transform 1 0 3832 0 1 2732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5992_6
timestamp 1731220340
transform 1 0 3832 0 -1 2728
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5991_6
timestamp 1731220340
transform 1 0 3648 0 -1 2728
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5990_6
timestamp 1731220340
transform 1 0 3664 0 1 2732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5989_6
timestamp 1731220340
transform 1 0 3792 0 1 3044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5988_6
timestamp 1731220340
transform 1 0 3784 0 1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5987_6
timestamp 1731220340
transform 1 0 3768 0 1 3384
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5986_6
timestamp 1731220340
transform 1 0 3744 0 -1 3700
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5985_6
timestamp 1731220340
transform 1 0 3704 0 1 3704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5984_6
timestamp 1731220340
transform 1 0 3648 0 -1 3856
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5983_6
timestamp 1731220340
transform 1 0 3736 0 1 3864
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5982_6
timestamp 1731220340
transform 1 0 3624 0 1 3864
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5981_6
timestamp 1731220340
transform 1 0 3512 0 1 3864
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5980_6
timestamp 1731220340
transform 1 0 3400 0 1 3864
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5979_6
timestamp 1731220340
transform 1 0 3296 0 1 3864
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5978_6
timestamp 1731220340
transform 1 0 3184 0 1 3864
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5977_6
timestamp 1731220340
transform 1 0 3064 0 1 3864
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5976_6
timestamp 1731220340
transform 1 0 2944 0 1 3864
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5975_6
timestamp 1731220340
transform 1 0 2816 0 1 3864
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5974_6
timestamp 1731220340
transform 1 0 3008 0 -1 3856
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5973_6
timestamp 1731220340
transform 1 0 3216 0 -1 3856
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5972_6
timestamp 1731220340
transform 1 0 3432 0 -1 3856
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5971_6
timestamp 1731220340
transform 1 0 3312 0 1 3704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5970_6
timestamp 1731220340
transform 1 0 3120 0 1 3704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5969_6
timestamp 1731220340
transform 1 0 2928 0 1 3704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5968_6
timestamp 1731220340
transform 1 0 3504 0 1 3704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5967_6
timestamp 1731220340
transform 1 0 3504 0 -1 3700
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5966_6
timestamp 1731220340
transform 1 0 3272 0 -1 3700
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5965_6
timestamp 1731220340
transform 1 0 3040 0 -1 3700
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5964_6
timestamp 1731220340
transform 1 0 3448 0 1 3540
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5963_6
timestamp 1731220340
transform 1 0 3616 0 1 3540
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5962_6
timestamp 1731220340
transform 1 0 3512 0 -1 3540
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5961_6
timestamp 1731220340
transform 1 0 3344 0 -1 3540
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5960_6
timestamp 1731220340
transform 1 0 3400 0 1 3384
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5959_6
timestamp 1731220340
transform 1 0 3584 0 1 3384
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5958_6
timestamp 1731220340
transform 1 0 3688 0 -1 3368
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5957_6
timestamp 1731220340
transform 1 0 3528 0 -1 3368
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5956_6
timestamp 1731220340
transform 1 0 3368 0 -1 3368
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5955_6
timestamp 1731220340
transform 1 0 3520 0 1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5954_6
timestamp 1731220340
transform 1 0 3216 0 -1 3368
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5953_6
timestamp 1731220340
transform 1 0 3072 0 -1 3368
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5952_6
timestamp 1731220340
transform 1 0 2928 0 -1 3368
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5951_6
timestamp 1731220340
transform 1 0 2856 0 1 3384
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5950_6
timestamp 1731220340
transform 1 0 3040 0 1 3384
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5949_6
timestamp 1731220340
transform 1 0 3216 0 1 3384
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5948_6
timestamp 1731220340
transform 1 0 3168 0 -1 3540
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5947_6
timestamp 1731220340
transform 1 0 2992 0 -1 3540
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5946_6
timestamp 1731220340
transform 1 0 3288 0 1 3540
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5945_6
timestamp 1731220340
transform 1 0 3136 0 1 3540
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5944_6
timestamp 1731220340
transform 1 0 2992 0 1 3540
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5943_6
timestamp 1731220340
transform 1 0 2848 0 1 3540
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5942_6
timestamp 1731220340
transform 1 0 2712 0 1 3540
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5941_6
timestamp 1731220340
transform 1 0 2576 0 1 3540
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5940_6
timestamp 1731220340
transform 1 0 2448 0 1 3540
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5939_6
timestamp 1731220340
transform 1 0 2320 0 1 3540
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5938_6
timestamp 1731220340
transform 1 0 2440 0 -1 3540
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5937_6
timestamp 1731220340
transform 1 0 2624 0 -1 3540
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5936_6
timestamp 1731220340
transform 1 0 2808 0 -1 3540
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5935_6
timestamp 1731220340
transform 1 0 2672 0 1 3384
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5934_6
timestamp 1731220340
transform 1 0 2488 0 1 3384
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5933_6
timestamp 1731220340
transform 1 0 2304 0 1 3384
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5932_6
timestamp 1731220340
transform 1 0 2352 0 -1 3368
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5931_6
timestamp 1731220340
transform 1 0 2504 0 -1 3368
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5930_6
timestamp 1731220340
transform 1 0 2648 0 -1 3368
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5929_6
timestamp 1731220340
transform 1 0 2792 0 -1 3368
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5928_6
timestamp 1731220340
transform 1 0 3008 0 1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5927_6
timestamp 1731220340
transform 1 0 2776 0 1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5926_6
timestamp 1731220340
transform 1 0 2568 0 1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5925_6
timestamp 1731220340
transform 1 0 2392 0 1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5924_6
timestamp 1731220340
transform 1 0 2240 0 1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5923_6
timestamp 1731220340
transform 1 0 2256 0 -1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5922_6
timestamp 1731220340
transform 1 0 2352 0 -1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5921_6
timestamp 1731220340
transform 1 0 2448 0 -1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5920_6
timestamp 1731220340
transform 1 0 2544 0 -1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5919_6
timestamp 1731220340
transform 1 0 2640 0 -1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5918_6
timestamp 1731220340
transform 1 0 2736 0 -1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5917_6
timestamp 1731220340
transform 1 0 2832 0 -1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5916_6
timestamp 1731220340
transform 1 0 2928 0 -1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5915_6
timestamp 1731220340
transform 1 0 3024 0 -1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5914_6
timestamp 1731220340
transform 1 0 3120 0 -1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5913_6
timestamp 1731220340
transform 1 0 3216 0 -1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5912_6
timestamp 1731220340
transform 1 0 3256 0 1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5911_6
timestamp 1731220340
transform 1 0 3312 0 -1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5910_6
timestamp 1731220340
transform 1 0 3432 0 -1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5909_6
timestamp 1731220340
transform 1 0 3712 0 -1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5908_6
timestamp 1731220340
transform 1 0 3568 0 -1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5907_6
timestamp 1731220340
transform 1 0 3496 0 1 3044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5906_6
timestamp 1731220340
transform 1 0 3200 0 1 3044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5905_6
timestamp 1731220340
transform 1 0 2904 0 1 3044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5904_6
timestamp 1731220340
transform 1 0 2616 0 1 3044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5903_6
timestamp 1731220340
transform 1 0 2696 0 -1 3044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5902_6
timestamp 1731220340
transform 1 0 2992 0 -1 3044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5901_6
timestamp 1731220340
transform 1 0 3280 0 -1 3044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5900_6
timestamp 1731220340
transform 1 0 3568 0 -1 3044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5899_6
timestamp 1731220340
transform 1 0 3832 0 1 2888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5898_6
timestamp 1731220340
transform 1 0 3640 0 1 2888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5897_6
timestamp 1731220340
transform 1 0 3432 0 1 2888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5896_6
timestamp 1731220340
transform 1 0 3208 0 1 2888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5895_6
timestamp 1731220340
transform 1 0 2968 0 1 2888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5894_6
timestamp 1731220340
transform 1 0 2696 0 1 2888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5893_6
timestamp 1731220340
transform 1 0 3640 0 -1 2888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5892_6
timestamp 1731220340
transform 1 0 3424 0 -1 2888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5891_6
timestamp 1731220340
transform 1 0 3208 0 -1 2888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5890_6
timestamp 1731220340
transform 1 0 2984 0 -1 2888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5889_6
timestamp 1731220340
transform 1 0 3472 0 1 2732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5888_6
timestamp 1731220340
transform 1 0 3288 0 1 2732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5887_6
timestamp 1731220340
transform 1 0 3104 0 1 2732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5886_6
timestamp 1731220340
transform 1 0 2920 0 1 2732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5885_6
timestamp 1731220340
transform 1 0 3448 0 -1 2728
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5884_6
timestamp 1731220340
transform 1 0 3248 0 -1 2728
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5883_6
timestamp 1731220340
transform 1 0 3056 0 -1 2728
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5882_6
timestamp 1731220340
transform 1 0 2880 0 -1 2728
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5881_6
timestamp 1731220340
transform 1 0 2720 0 -1 2728
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5880_6
timestamp 1731220340
transform 1 0 2784 0 1 2568
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5879_6
timestamp 1731220340
transform 1 0 2904 0 1 2568
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5878_6
timestamp 1731220340
transform 1 0 3144 0 1 2568
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5877_6
timestamp 1731220340
transform 1 0 3024 0 1 2568
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5876_6
timestamp 1731220340
transform 1 0 2984 0 -1 2564
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5875_6
timestamp 1731220340
transform 1 0 3104 0 -1 2564
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5874_6
timestamp 1731220340
transform 1 0 3224 0 -1 2564
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5873_6
timestamp 1731220340
transform 1 0 3352 0 -1 2564
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5872_6
timestamp 1731220340
transform 1 0 3480 0 -1 2564
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5871_6
timestamp 1731220340
transform 1 0 3352 0 1 2408
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5870_6
timestamp 1731220340
transform 1 0 3200 0 1 2408
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5869_6
timestamp 1731220340
transform 1 0 3496 0 1 2408
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5868_6
timestamp 1731220340
transform 1 0 3648 0 1 2408
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5867_6
timestamp 1731220340
transform 1 0 3800 0 1 2408
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5866_6
timestamp 1731220340
transform 1 0 3832 0 -1 2396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5865_6
timestamp 1731220340
transform 1 0 3672 0 -1 2396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5864_6
timestamp 1731220340
transform 1 0 3512 0 -1 2396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5863_6
timestamp 1731220340
transform 1 0 3352 0 -1 2396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5862_6
timestamp 1731220340
transform 1 0 3184 0 -1 2396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5861_6
timestamp 1731220340
transform 1 0 3688 0 1 2228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5860_6
timestamp 1731220340
transform 1 0 3528 0 1 2228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5859_6
timestamp 1731220340
transform 1 0 3376 0 1 2228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5858_6
timestamp 1731220340
transform 1 0 3224 0 1 2228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5857_6
timestamp 1731220340
transform 1 0 3064 0 1 2228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5856_6
timestamp 1731220340
transform 1 0 3512 0 -1 2228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5855_6
timestamp 1731220340
transform 1 0 3360 0 -1 2228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5854_6
timestamp 1731220340
transform 1 0 3216 0 -1 2228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5853_6
timestamp 1731220340
transform 1 0 3072 0 -1 2228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5852_6
timestamp 1731220340
transform 1 0 2928 0 -1 2228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5851_6
timestamp 1731220340
transform 1 0 3512 0 1 2056
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5850_6
timestamp 1731220340
transform 1 0 3344 0 1 2056
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5849_6
timestamp 1731220340
transform 1 0 3184 0 1 2056
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5848_6
timestamp 1731220340
transform 1 0 3032 0 1 2056
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5847_6
timestamp 1731220340
transform 1 0 2888 0 1 2056
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5846_6
timestamp 1731220340
transform 1 0 3448 0 -1 2048
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5845_6
timestamp 1731220340
transform 1 0 3256 0 -1 2048
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5844_6
timestamp 1731220340
transform 1 0 3072 0 -1 2048
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5843_6
timestamp 1731220340
transform 1 0 2912 0 -1 2048
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5842_6
timestamp 1731220340
transform 1 0 2768 0 -1 2048
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5841_6
timestamp 1731220340
transform 1 0 2760 0 1 1892
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5840_6
timestamp 1731220340
transform 1 0 2912 0 1 1892
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5839_6
timestamp 1731220340
transform 1 0 3096 0 1 1892
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5838_6
timestamp 1731220340
transform 1 0 3312 0 1 1892
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5837_6
timestamp 1731220340
transform 1 0 3536 0 1 1892
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5836_6
timestamp 1731220340
transform 1 0 3624 0 -1 1880
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5835_6
timestamp 1731220340
transform 1 0 3392 0 -1 1880
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5834_6
timestamp 1731220340
transform 1 0 3176 0 -1 1880
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5833_6
timestamp 1731220340
transform 1 0 2984 0 -1 1880
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5832_6
timestamp 1731220340
transform 1 0 2824 0 -1 1880
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5831_6
timestamp 1731220340
transform 1 0 2872 0 1 1724
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5830_6
timestamp 1731220340
transform 1 0 3064 0 1 1724
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5829_6
timestamp 1731220340
transform 1 0 3256 0 1 1724
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5828_6
timestamp 1731220340
transform 1 0 3456 0 1 1724
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5827_6
timestamp 1731220340
transform 1 0 3440 0 -1 1720
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5826_6
timestamp 1731220340
transform 1 0 3248 0 -1 1720
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5825_6
timestamp 1731220340
transform 1 0 3056 0 -1 1720
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5824_6
timestamp 1731220340
transform 1 0 3040 0 1 1568
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5823_6
timestamp 1731220340
transform 1 0 2832 0 1 1568
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5822_6
timestamp 1731220340
transform 1 0 3224 0 1 1568
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5821_6
timestamp 1731220340
transform 1 0 3392 0 1 1568
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5820_6
timestamp 1731220340
transform 1 0 3376 0 -1 1564
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5819_6
timestamp 1731220340
transform 1 0 3216 0 -1 1564
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5818_6
timestamp 1731220340
transform 1 0 3536 0 -1 1564
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5817_6
timestamp 1731220340
transform 1 0 3696 0 -1 1564
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5816_6
timestamp 1731220340
transform 1 0 3688 0 1 1568
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5815_6
timestamp 1731220340
transform 1 0 3544 0 1 1568
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5814_6
timestamp 1731220340
transform 1 0 3640 0 -1 1720
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5813_6
timestamp 1731220340
transform 1 0 3656 0 1 1724
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5812_6
timestamp 1731220340
transform 1 0 3768 0 1 1892
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5811_6
timestamp 1731220340
transform 1 0 3832 0 1 2056
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5810_6
timestamp 1731220340
transform 1 0 3680 0 1 2056
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5809_6
timestamp 1731220340
transform 1 0 3648 0 -1 2048
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5808_6
timestamp 1731220340
transform 1 0 3832 0 -1 2048
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5807_6
timestamp 1731220340
transform 1 0 3832 0 -1 1880
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5806_6
timestamp 1731220340
transform 1 0 3832 0 1 1724
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5805_6
timestamp 1731220340
transform 1 0 3832 0 -1 1720
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5804_6
timestamp 1731220340
transform 1 0 3832 0 1 1568
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5803_6
timestamp 1731220340
transform 1 0 3808 0 1 1412
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5802_6
timestamp 1731220340
transform 1 0 3808 0 -1 1392
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5801_6
timestamp 1731220340
transform 1 0 3824 0 1 1232
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5800_6
timestamp 1731220340
transform 1 0 3832 0 -1 1224
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5799_6
timestamp 1731220340
transform 1 0 3832 0 1 1064
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5798_6
timestamp 1731220340
transform 1 0 3832 0 -1 1060
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5797_6
timestamp 1731220340
transform 1 0 3832 0 1 908
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5796_6
timestamp 1731220340
transform 1 0 3832 0 -1 896
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5795_6
timestamp 1731220340
transform 1 0 3832 0 1 744
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5794_6
timestamp 1731220340
transform 1 0 3832 0 -1 740
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5793_6
timestamp 1731220340
transform 1 0 3824 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5792_6
timestamp 1731220340
transform 1 0 3832 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5791_6
timestamp 1731220340
transform 1 0 3640 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5790_6
timestamp 1731220340
transform 1 0 3448 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5789_6
timestamp 1731220340
transform 1 0 3296 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5788_6
timestamp 1731220340
transform 1 0 3472 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5787_6
timestamp 1731220340
transform 1 0 3648 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5786_6
timestamp 1731220340
transform 1 0 3672 0 -1 740
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5785_6
timestamp 1731220340
transform 1 0 3512 0 -1 740
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5784_6
timestamp 1731220340
transform 1 0 3360 0 -1 740
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5783_6
timestamp 1731220340
transform 1 0 3208 0 -1 740
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5782_6
timestamp 1731220340
transform 1 0 3240 0 1 744
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5781_6
timestamp 1731220340
transform 1 0 3440 0 1 744
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5780_6
timestamp 1731220340
transform 1 0 3648 0 1 744
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5779_6
timestamp 1731220340
transform 1 0 3608 0 -1 896
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5778_6
timestamp 1731220340
transform 1 0 3360 0 -1 896
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5777_6
timestamp 1731220340
transform 1 0 3120 0 -1 896
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5776_6
timestamp 1731220340
transform 1 0 3656 0 1 908
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5775_6
timestamp 1731220340
transform 1 0 3456 0 1 908
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5774_6
timestamp 1731220340
transform 1 0 3272 0 1 908
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5773_6
timestamp 1731220340
transform 1 0 3104 0 1 908
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5772_6
timestamp 1731220340
transform 1 0 2960 0 1 908
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5771_6
timestamp 1731220340
transform 1 0 3000 0 -1 1060
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5770_6
timestamp 1731220340
transform 1 0 3624 0 -1 1060
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5769_6
timestamp 1731220340
transform 1 0 3400 0 -1 1060
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5768_6
timestamp 1731220340
transform 1 0 3192 0 -1 1060
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5767_6
timestamp 1731220340
transform 1 0 3144 0 1 1064
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5766_6
timestamp 1731220340
transform 1 0 2984 0 1 1064
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5765_6
timestamp 1731220340
transform 1 0 3312 0 1 1064
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5764_6
timestamp 1731220340
transform 1 0 3672 0 1 1064
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5763_6
timestamp 1731220340
transform 1 0 3488 0 1 1064
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5762_6
timestamp 1731220340
transform 1 0 3392 0 -1 1224
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5761_6
timestamp 1731220340
transform 1 0 3232 0 -1 1224
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5760_6
timestamp 1731220340
transform 1 0 3064 0 -1 1224
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5759_6
timestamp 1731220340
transform 1 0 3544 0 -1 1224
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5758_6
timestamp 1731220340
transform 1 0 3696 0 -1 1224
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5757_6
timestamp 1731220340
transform 1 0 3656 0 1 1232
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5756_6
timestamp 1731220340
transform 1 0 3496 0 1 1232
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5755_6
timestamp 1731220340
transform 1 0 3336 0 1 1232
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5754_6
timestamp 1731220340
transform 1 0 3168 0 1 1232
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5753_6
timestamp 1731220340
transform 1 0 2992 0 1 1232
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5752_6
timestamp 1731220340
transform 1 0 3552 0 -1 1392
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5751_6
timestamp 1731220340
transform 1 0 3296 0 -1 1392
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5750_6
timestamp 1731220340
transform 1 0 3048 0 -1 1392
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5749_6
timestamp 1731220340
transform 1 0 2800 0 -1 1392
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5748_6
timestamp 1731220340
transform 1 0 2552 0 -1 1392
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5747_6
timestamp 1731220340
transform 1 0 3608 0 1 1412
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5746_6
timestamp 1731220340
transform 1 0 3408 0 1 1412
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5745_6
timestamp 1731220340
transform 1 0 3224 0 1 1412
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5744_6
timestamp 1731220340
transform 1 0 3056 0 1 1412
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5743_6
timestamp 1731220340
transform 1 0 2912 0 1 1412
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5742_6
timestamp 1731220340
transform 1 0 2792 0 1 1412
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5741_6
timestamp 1731220340
transform 1 0 2696 0 1 1412
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5740_6
timestamp 1731220340
transform 1 0 2600 0 1 1412
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5739_6
timestamp 1731220340
transform 1 0 2504 0 1 1412
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5738_6
timestamp 1731220340
transform 1 0 2408 0 1 1412
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5737_6
timestamp 1731220340
transform 1 0 3056 0 -1 1564
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5736_6
timestamp 1731220340
transform 1 0 2896 0 -1 1564
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5735_6
timestamp 1731220340
transform 1 0 2736 0 -1 1564
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5734_6
timestamp 1731220340
transform 1 0 2576 0 -1 1564
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5733_6
timestamp 1731220340
transform 1 0 2592 0 1 1568
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5732_6
timestamp 1731220340
transform 1 0 2680 0 -1 1720
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5731_6
timestamp 1731220340
transform 1 0 2864 0 -1 1720
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5730_6
timestamp 1731220340
transform 1 0 2680 0 1 1724
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5729_6
timestamp 1731220340
transform 1 0 2696 0 -1 1880
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5728_6
timestamp 1731220340
transform 1 0 2584 0 -1 1880
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5727_6
timestamp 1731220340
transform 1 0 2640 0 1 1892
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5726_6
timestamp 1731220340
transform 1 0 2640 0 -1 2048
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5725_6
timestamp 1731220340
transform 1 0 2624 0 1 2056
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5724_6
timestamp 1731220340
transform 1 0 2752 0 1 2056
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5723_6
timestamp 1731220340
transform 1 0 2776 0 -1 2228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5722_6
timestamp 1731220340
transform 1 0 2904 0 1 2228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5721_6
timestamp 1731220340
transform 1 0 2808 0 -1 2396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5720_6
timestamp 1731220340
transform 1 0 2600 0 -1 2396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5719_6
timestamp 1731220340
transform 1 0 3000 0 -1 2396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5718_6
timestamp 1731220340
transform 1 0 3040 0 1 2408
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5717_6
timestamp 1731220340
transform 1 0 2872 0 1 2408
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5716_6
timestamp 1731220340
transform 1 0 2704 0 1 2408
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5715_6
timestamp 1731220340
transform 1 0 2528 0 1 2408
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5714_6
timestamp 1731220340
transform 1 0 2864 0 -1 2564
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5713_6
timestamp 1731220340
transform 1 0 2736 0 -1 2564
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5712_6
timestamp 1731220340
transform 1 0 2608 0 -1 2564
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5711_6
timestamp 1731220340
transform 1 0 2488 0 -1 2564
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5710_6
timestamp 1731220340
transform 1 0 2376 0 -1 2564
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5709_6
timestamp 1731220340
transform 1 0 2664 0 1 2568
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5708_6
timestamp 1731220340
transform 1 0 2552 0 1 2568
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5707_6
timestamp 1731220340
transform 1 0 2440 0 1 2568
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5706_6
timestamp 1731220340
transform 1 0 2328 0 1 2568
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5705_6
timestamp 1731220340
transform 1 0 2224 0 1 2568
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5704_6
timestamp 1731220340
transform 1 0 2576 0 -1 2728
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5703_6
timestamp 1731220340
transform 1 0 2440 0 -1 2728
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5702_6
timestamp 1731220340
transform 1 0 2312 0 -1 2728
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5701_6
timestamp 1731220340
transform 1 0 2184 0 -1 2728
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5700_6
timestamp 1731220340
transform 1 0 2064 0 -1 2728
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5699_6
timestamp 1731220340
transform 1 0 2728 0 1 2732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5698_6
timestamp 1731220340
transform 1 0 2544 0 1 2732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5697_6
timestamp 1731220340
transform 1 0 2360 0 1 2732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5696_6
timestamp 1731220340
transform 1 0 2192 0 1 2732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5695_6
timestamp 1731220340
transform 1 0 2064 0 1 2732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5694_6
timestamp 1731220340
transform 1 0 2760 0 -1 2888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5693_6
timestamp 1731220340
transform 1 0 2528 0 -1 2888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5692_6
timestamp 1731220340
transform 1 0 2288 0 -1 2888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5691_6
timestamp 1731220340
transform 1 0 2064 0 -1 2888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5690_6
timestamp 1731220340
transform 1 0 2064 0 1 2888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5689_6
timestamp 1731220340
transform 1 0 2384 0 1 2888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5688_6
timestamp 1731220340
transform 1 0 2376 0 -1 3044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5687_6
timestamp 1731220340
transform 1 0 2064 0 -1 3044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5686_6
timestamp 1731220340
transform 1 0 2064 0 1 3044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5685_6
timestamp 1731220340
transform 1 0 2328 0 1 3044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5684_6
timestamp 1731220340
transform 1 0 2160 0 -1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5683_6
timestamp 1731220340
transform 1 0 2064 0 -1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5682_6
timestamp 1731220340
transform 1 0 2104 0 1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5681_6
timestamp 1731220340
transform 1 0 2064 0 -1 3368
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5680_6
timestamp 1731220340
transform 1 0 2208 0 -1 3368
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5679_6
timestamp 1731220340
transform 1 0 2120 0 1 3384
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5678_6
timestamp 1731220340
transform 1 0 2096 0 -1 3540
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5677_6
timestamp 1731220340
transform 1 0 2264 0 -1 3540
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5676_6
timestamp 1731220340
transform 1 0 2184 0 1 3540
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5675_6
timestamp 1731220340
transform 1 0 2120 0 -1 3700
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5674_6
timestamp 1731220340
transform 1 0 2344 0 -1 3700
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5673_6
timestamp 1731220340
transform 1 0 2576 0 -1 3700
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5672_6
timestamp 1731220340
transform 1 0 2808 0 -1 3700
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5671_6
timestamp 1731220340
transform 1 0 2736 0 1 3704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5670_6
timestamp 1731220340
transform 1 0 2552 0 1 3704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5669_6
timestamp 1731220340
transform 1 0 2368 0 1 3704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5668_6
timestamp 1731220340
transform 1 0 2184 0 1 3704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5667_6
timestamp 1731220340
transform 1 0 2200 0 -1 3856
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5666_6
timestamp 1731220340
transform 1 0 2336 0 -1 3856
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5665_6
timestamp 1731220340
transform 1 0 2480 0 -1 3856
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5664_6
timestamp 1731220340
transform 1 0 2640 0 -1 3856
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5663_6
timestamp 1731220340
transform 1 0 2816 0 -1 3856
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5662_6
timestamp 1731220340
transform 1 0 2680 0 1 3864
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5661_6
timestamp 1731220340
transform 1 0 2544 0 1 3864
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5660_6
timestamp 1731220340
transform 1 0 2408 0 1 3864
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5659_6
timestamp 1731220340
transform 1 0 2280 0 1 3864
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5658_6
timestamp 1731220340
transform 1 0 2152 0 1 3864
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5657_6
timestamp 1731220340
transform 1 0 2256 0 -1 4016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5656_6
timestamp 1731220340
transform 1 0 2160 0 -1 4016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5655_6
timestamp 1731220340
transform 1 0 2064 0 -1 4016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5654_6
timestamp 1731220340
transform 1 0 1896 0 1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5653_6
timestamp 1731220340
transform 1 0 1800 0 1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5652_6
timestamp 1731220340
transform 1 0 1704 0 1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5651_6
timestamp 1731220340
transform 1 0 1608 0 1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5650_6
timestamp 1731220340
transform 1 0 1512 0 1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5649_6
timestamp 1731220340
transform 1 0 1640 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5648_6
timestamp 1731220340
transform 1 0 1504 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5647_6
timestamp 1731220340
transform 1 0 1376 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5646_6
timestamp 1731220340
transform 1 0 1248 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5645_6
timestamp 1731220340
transform 1 0 1120 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5644_6
timestamp 1731220340
transform 1 0 1096 0 1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5643_6
timestamp 1731220340
transform 1 0 1224 0 1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5642_6
timestamp 1731220340
transform 1 0 1352 0 1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5641_6
timestamp 1731220340
transform 1 0 1480 0 1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5640_6
timestamp 1731220340
transform 1 0 1424 0 -1 3796
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5639_6
timestamp 1731220340
transform 1 0 1280 0 -1 3796
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5638_6
timestamp 1731220340
transform 1 0 1576 0 -1 3796
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5637_6
timestamp 1731220340
transform 1 0 1488 0 1 3636
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5636_6
timestamp 1731220340
transform 1 0 1648 0 1 3636
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5635_6
timestamp 1731220340
transform 1 0 1608 0 -1 3628
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5634_6
timestamp 1731220340
transform 1 0 1432 0 -1 3628
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5633_6
timestamp 1731220340
transform 1 0 1784 0 -1 3628
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5632_6
timestamp 1731220340
transform 1 0 1872 0 1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5631_6
timestamp 1731220340
transform 1 0 1696 0 1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5630_6
timestamp 1731220340
transform 1 0 1520 0 1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5629_6
timestamp 1731220340
transform 1 0 1528 0 -1 3456
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5628_6
timestamp 1731220340
transform 1 0 1712 0 -1 3456
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5627_6
timestamp 1731220340
transform 1 0 1896 0 -1 3456
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5626_6
timestamp 1731220340
transform 1 0 1864 0 1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5625_6
timestamp 1731220340
transform 1 0 1696 0 1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5624_6
timestamp 1731220340
transform 1 0 1536 0 1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5623_6
timestamp 1731220340
transform 1 0 1512 0 -1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5622_6
timestamp 1731220340
transform 1 0 1736 0 -1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5621_6
timestamp 1731220340
transform 1 0 1688 0 1 3152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5620_6
timestamp 1731220340
transform 1 0 1504 0 1 3152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5619_6
timestamp 1731220340
transform 1 0 1384 0 -1 3148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5618_6
timestamp 1731220340
transform 1 0 1552 0 -1 3148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5617_6
timestamp 1731220340
transform 1 0 1720 0 -1 3148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5616_6
timestamp 1731220340
transform 1 0 1712 0 1 2988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5615_6
timestamp 1731220340
transform 1 0 1544 0 1 2988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5614_6
timestamp 1731220340
transform 1 0 1480 0 -1 2984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5613_6
timestamp 1731220340
transform 1 0 1648 0 -1 2984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5612_6
timestamp 1731220340
transform 1 0 1816 0 -1 2984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5611_6
timestamp 1731220340
transform 1 0 1840 0 1 2824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5610_6
timestamp 1731220340
transform 1 0 1664 0 1 2824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5609_6
timestamp 1731220340
transform 1 0 1488 0 1 2824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5608_6
timestamp 1731220340
transform 1 0 1592 0 -1 2820
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5607_6
timestamp 1731220340
transform 1 0 1776 0 -1 2820
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5606_6
timestamp 1731220340
transform 1 0 1776 0 1 2664
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5605_6
timestamp 1731220340
transform 1 0 1616 0 1 2664
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5604_6
timestamp 1731220340
transform 1 0 1456 0 1 2664
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5603_6
timestamp 1731220340
transform 1 0 1424 0 -1 2660
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5602_6
timestamp 1731220340
transform 1 0 1560 0 -1 2660
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5601_6
timestamp 1731220340
transform 1 0 1696 0 -1 2660
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5600_6
timestamp 1731220340
transform 1 0 1720 0 1 2508
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5599_6
timestamp 1731220340
transform 1 0 1584 0 1 2508
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5598_6
timestamp 1731220340
transform 1 0 1456 0 1 2508
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5597_6
timestamp 1731220340
transform 1 0 1328 0 1 2508
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5596_6
timestamp 1731220340
transform 1 0 1192 0 1 2508
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5595_6
timestamp 1731220340
transform 1 0 1056 0 1 2508
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5594_6
timestamp 1731220340
transform 1 0 912 0 1 2508
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5593_6
timestamp 1731220340
transform 1 0 1024 0 -1 2660
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5592_6
timestamp 1731220340
transform 1 0 1160 0 -1 2660
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5591_6
timestamp 1731220340
transform 1 0 1296 0 -1 2660
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5590_6
timestamp 1731220340
transform 1 0 1304 0 1 2664
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5589_6
timestamp 1731220340
transform 1 0 1152 0 1 2664
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5588_6
timestamp 1731220340
transform 1 0 1072 0 -1 2820
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5587_6
timestamp 1731220340
transform 1 0 1232 0 -1 2820
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5586_6
timestamp 1731220340
transform 1 0 1408 0 -1 2820
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5585_6
timestamp 1731220340
transform 1 0 1312 0 1 2824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5584_6
timestamp 1731220340
transform 1 0 1144 0 1 2824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5583_6
timestamp 1731220340
transform 1 0 1320 0 -1 2984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5582_6
timestamp 1731220340
transform 1 0 1168 0 -1 2984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5581_6
timestamp 1731220340
transform 1 0 1064 0 1 2988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5580_6
timestamp 1731220340
transform 1 0 1216 0 1 2988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5579_6
timestamp 1731220340
transform 1 0 1376 0 1 2988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5578_6
timestamp 1731220340
transform 1 0 1216 0 -1 3148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5577_6
timestamp 1731220340
transform 1 0 1056 0 -1 3148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5576_6
timestamp 1731220340
transform 1 0 960 0 1 3152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5575_6
timestamp 1731220340
transform 1 0 1136 0 1 3152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5574_6
timestamp 1731220340
transform 1 0 1320 0 1 3152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5573_6
timestamp 1731220340
transform 1 0 1288 0 -1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5572_6
timestamp 1731220340
transform 1 0 1072 0 -1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5571_6
timestamp 1731220340
transform 1 0 1040 0 1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5570_6
timestamp 1731220340
transform 1 0 1208 0 1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5569_6
timestamp 1731220340
transform 1 0 1376 0 1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5568_6
timestamp 1731220340
transform 1 0 1344 0 -1 3456
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5567_6
timestamp 1731220340
transform 1 0 1152 0 -1 3456
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5566_6
timestamp 1731220340
transform 1 0 952 0 -1 3456
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5565_6
timestamp 1731220340
transform 1 0 992 0 1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5564_6
timestamp 1731220340
transform 1 0 1168 0 1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5563_6
timestamp 1731220340
transform 1 0 1344 0 1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5562_6
timestamp 1731220340
transform 1 0 1256 0 -1 3628
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5561_6
timestamp 1731220340
transform 1 0 1088 0 -1 3628
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5560_6
timestamp 1731220340
transform 1 0 1032 0 1 3636
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5559_6
timestamp 1731220340
transform 1 0 1328 0 1 3636
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5558_6
timestamp 1731220340
transform 1 0 1176 0 1 3636
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5557_6
timestamp 1731220340
transform 1 0 1136 0 -1 3796
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5556_6
timestamp 1731220340
transform 1 0 992 0 -1 3796
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5555_6
timestamp 1731220340
transform 1 0 968 0 1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5554_6
timestamp 1731220340
transform 1 0 840 0 1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5553_6
timestamp 1731220340
transform 1 0 712 0 1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5552_6
timestamp 1731220340
transform 1 0 992 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5551_6
timestamp 1731220340
transform 1 0 864 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5550_6
timestamp 1731220340
transform 1 0 736 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5549_6
timestamp 1731220340
transform 1 0 608 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5548_6
timestamp 1731220340
transform 1 0 488 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5547_6
timestamp 1731220340
transform 1 0 384 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5546_6
timestamp 1731220340
transform 1 0 288 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5545_6
timestamp 1731220340
transform 1 0 192 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5544_6
timestamp 1731220340
transform 1 0 328 0 1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5543_6
timestamp 1731220340
transform 1 0 448 0 1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5542_6
timestamp 1731220340
transform 1 0 576 0 1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5541_6
timestamp 1731220340
transform 1 0 496 0 -1 3796
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5540_6
timestamp 1731220340
transform 1 0 608 0 -1 3796
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5539_6
timestamp 1731220340
transform 1 0 728 0 -1 3796
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5538_6
timestamp 1731220340
transform 1 0 856 0 -1 3796
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5537_6
timestamp 1731220340
transform 1 0 904 0 1 3636
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5536_6
timestamp 1731220340
transform 1 0 784 0 1 3636
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5535_6
timestamp 1731220340
transform 1 0 680 0 1 3636
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5534_6
timestamp 1731220340
transform 1 0 584 0 1 3636
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5533_6
timestamp 1731220340
transform 1 0 488 0 1 3636
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5532_6
timestamp 1731220340
transform 1 0 920 0 -1 3628
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5531_6
timestamp 1731220340
transform 1 0 752 0 -1 3628
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5530_6
timestamp 1731220340
transform 1 0 600 0 -1 3628
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5529_6
timestamp 1731220340
transform 1 0 456 0 -1 3628
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5528_6
timestamp 1731220340
transform 1 0 328 0 -1 3628
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5527_6
timestamp 1731220340
transform 1 0 808 0 1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5526_6
timestamp 1731220340
transform 1 0 632 0 1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5525_6
timestamp 1731220340
transform 1 0 456 0 1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5524_6
timestamp 1731220340
transform 1 0 296 0 1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5523_6
timestamp 1731220340
transform 1 0 152 0 1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5522_6
timestamp 1731220340
transform 1 0 744 0 -1 3456
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5521_6
timestamp 1731220340
transform 1 0 528 0 -1 3456
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5520_6
timestamp 1731220340
transform 1 0 312 0 -1 3456
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5519_6
timestamp 1731220340
transform 1 0 128 0 -1 3456
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5518_6
timestamp 1731220340
transform 1 0 864 0 1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5517_6
timestamp 1731220340
transform 1 0 696 0 1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5516_6
timestamp 1731220340
transform 1 0 528 0 1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5515_6
timestamp 1731220340
transform 1 0 368 0 1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5514_6
timestamp 1731220340
transform 1 0 224 0 1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5513_6
timestamp 1731220340
transform 1 0 128 0 1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5512_6
timestamp 1731220340
transform 1 0 128 0 -1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5511_6
timestamp 1731220340
transform 1 0 272 0 -1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5510_6
timestamp 1731220340
transform 1 0 864 0 -1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5509_6
timestamp 1731220340
transform 1 0 656 0 -1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5508_6
timestamp 1731220340
transform 1 0 456 0 -1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5507_6
timestamp 1731220340
transform 1 0 440 0 1 3152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5506_6
timestamp 1731220340
transform 1 0 280 0 1 3152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5505_6
timestamp 1731220340
transform 1 0 128 0 1 3152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5504_6
timestamp 1731220340
transform 1 0 608 0 1 3152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5503_6
timestamp 1731220340
transform 1 0 784 0 1 3152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5502_6
timestamp 1731220340
transform 1 0 896 0 -1 3148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5501_6
timestamp 1731220340
transform 1 0 736 0 -1 3148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5500_6
timestamp 1731220340
transform 1 0 576 0 -1 3148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5499_6
timestamp 1731220340
transform 1 0 432 0 -1 3148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5498_6
timestamp 1731220340
transform 1 0 304 0 -1 3148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5497_6
timestamp 1731220340
transform 1 0 496 0 1 2988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5496_6
timestamp 1731220340
transform 1 0 592 0 1 2988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5495_6
timestamp 1731220340
transform 1 0 696 0 1 2988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5494_6
timestamp 1731220340
transform 1 0 808 0 1 2988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5493_6
timestamp 1731220340
transform 1 0 928 0 1 2988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5492_6
timestamp 1731220340
transform 1 0 1016 0 -1 2984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5491_6
timestamp 1731220340
transform 1 0 880 0 -1 2984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5490_6
timestamp 1731220340
transform 1 0 752 0 -1 2984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5489_6
timestamp 1731220340
transform 1 0 640 0 -1 2984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5488_6
timestamp 1731220340
transform 1 0 544 0 -1 2984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5487_6
timestamp 1731220340
transform 1 0 984 0 1 2824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5486_6
timestamp 1731220340
transform 1 0 832 0 1 2824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5485_6
timestamp 1731220340
transform 1 0 688 0 1 2824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5484_6
timestamp 1731220340
transform 1 0 568 0 1 2824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5483_6
timestamp 1731220340
transform 1 0 464 0 1 2824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5482_6
timestamp 1731220340
transform 1 0 472 0 -1 2820
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5481_6
timestamp 1731220340
transform 1 0 568 0 -1 2820
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5480_6
timestamp 1731220340
transform 1 0 672 0 -1 2820
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5479_6
timestamp 1731220340
transform 1 0 792 0 -1 2820
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5478_6
timestamp 1731220340
transform 1 0 928 0 -1 2820
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5477_6
timestamp 1731220340
transform 1 0 1008 0 1 2664
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5476_6
timestamp 1731220340
transform 1 0 872 0 1 2664
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5475_6
timestamp 1731220340
transform 1 0 736 0 1 2664
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5474_6
timestamp 1731220340
transform 1 0 616 0 1 2664
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5473_6
timestamp 1731220340
transform 1 0 504 0 1 2664
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5472_6
timestamp 1731220340
transform 1 0 888 0 -1 2660
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5471_6
timestamp 1731220340
transform 1 0 744 0 -1 2660
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5470_6
timestamp 1731220340
transform 1 0 608 0 -1 2660
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5469_6
timestamp 1731220340
transform 1 0 480 0 -1 2660
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5468_6
timestamp 1731220340
transform 1 0 360 0 -1 2660
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5467_6
timestamp 1731220340
transform 1 0 760 0 1 2508
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5466_6
timestamp 1731220340
transform 1 0 600 0 1 2508
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5465_6
timestamp 1731220340
transform 1 0 440 0 1 2508
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5464_6
timestamp 1731220340
transform 1 0 280 0 1 2508
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5463_6
timestamp 1731220340
transform 1 0 128 0 1 2508
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5462_6
timestamp 1731220340
transform 1 0 512 0 -1 2492
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5461_6
timestamp 1731220340
transform 1 0 416 0 -1 2492
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5460_6
timestamp 1731220340
transform 1 0 320 0 -1 2492
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5459_6
timestamp 1731220340
transform 1 0 224 0 -1 2492
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5458_6
timestamp 1731220340
transform 1 0 128 0 -1 2492
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5457_6
timestamp 1731220340
transform 1 0 128 0 1 2324
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5456_6
timestamp 1731220340
transform 1 0 248 0 1 2324
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5455_6
timestamp 1731220340
transform 1 0 408 0 1 2324
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5454_6
timestamp 1731220340
transform 1 0 568 0 1 2324
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5453_6
timestamp 1731220340
transform 1 0 728 0 1 2324
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5452_6
timestamp 1731220340
transform 1 0 736 0 -1 2324
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5451_6
timestamp 1731220340
transform 1 0 576 0 -1 2324
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5450_6
timestamp 1731220340
transform 1 0 416 0 -1 2324
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5449_6
timestamp 1731220340
transform 1 0 256 0 -1 2324
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5448_6
timestamp 1731220340
transform 1 0 128 0 -1 2324
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5447_6
timestamp 1731220340
transform 1 0 216 0 1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5446_6
timestamp 1731220340
transform 1 0 344 0 1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5445_6
timestamp 1731220340
transform 1 0 488 0 1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5444_6
timestamp 1731220340
transform 1 0 640 0 1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5443_6
timestamp 1731220340
transform 1 0 792 0 1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5442_6
timestamp 1731220340
transform 1 0 672 0 -1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5441_6
timestamp 1731220340
transform 1 0 560 0 -1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5440_6
timestamp 1731220340
transform 1 0 464 0 -1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5439_6
timestamp 1731220340
transform 1 0 800 0 -1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5438_6
timestamp 1731220340
transform 1 0 936 0 -1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5437_6
timestamp 1731220340
transform 1 0 1112 0 1 2016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5436_6
timestamp 1731220340
transform 1 0 976 0 1 2016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5435_6
timestamp 1731220340
transform 1 0 848 0 1 2016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5434_6
timestamp 1731220340
transform 1 0 728 0 1 2016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5433_6
timestamp 1731220340
transform 1 0 616 0 1 2016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5432_6
timestamp 1731220340
transform 1 0 880 0 -1 2012
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5431_6
timestamp 1731220340
transform 1 0 720 0 -1 2012
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5430_6
timestamp 1731220340
transform 1 0 568 0 -1 2012
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5429_6
timestamp 1731220340
transform 1 0 440 0 -1 2012
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5428_6
timestamp 1731220340
transform 1 0 440 0 -1 1860
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5427_6
timestamp 1731220340
transform 1 0 312 0 -1 1860
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5426_6
timestamp 1731220340
transform 1 0 248 0 1 1704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5425_6
timestamp 1731220340
transform 1 0 384 0 1 1704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5424_6
timestamp 1731220340
transform 1 0 424 0 -1 1704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5423_6
timestamp 1731220340
transform 1 0 256 0 -1 1704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5422_6
timestamp 1731220340
transform 1 0 128 0 -1 1704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5421_6
timestamp 1731220340
transform 1 0 128 0 1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5420_6
timestamp 1731220340
transform 1 0 280 0 1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5419_6
timestamp 1731220340
transform 1 0 480 0 -1 1548
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5418_6
timestamp 1731220340
transform 1 0 288 0 -1 1548
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5417_6
timestamp 1731220340
transform 1 0 128 0 -1 1548
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5416_6
timestamp 1731220340
transform 1 0 168 0 1 1396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5415_6
timestamp 1731220340
transform 1 0 352 0 1 1396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5414_6
timestamp 1731220340
transform 1 0 320 0 -1 1396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5413_6
timestamp 1731220340
transform 1 0 560 0 1 1396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5412_6
timestamp 1731220340
transform 1 0 776 0 1 1396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5411_6
timestamp 1731220340
transform 1 0 880 0 -1 1548
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5410_6
timestamp 1731220340
transform 1 0 680 0 -1 1548
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5409_6
timestamp 1731220340
transform 1 0 648 0 1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5408_6
timestamp 1731220340
transform 1 0 464 0 1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5407_6
timestamp 1731220340
transform 1 0 832 0 1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5406_6
timestamp 1731220340
transform 1 0 792 0 -1 1704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5405_6
timestamp 1731220340
transform 1 0 600 0 -1 1704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5404_6
timestamp 1731220340
transform 1 0 528 0 1 1704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5403_6
timestamp 1731220340
transform 1 0 688 0 1 1704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5402_6
timestamp 1731220340
transform 1 0 856 0 1 1704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5401_6
timestamp 1731220340
transform 1 0 848 0 -1 1860
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5400_6
timestamp 1731220340
transform 1 0 712 0 -1 1860
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5399_6
timestamp 1731220340
transform 1 0 576 0 -1 1860
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5398_6
timestamp 1731220340
transform 1 0 648 0 1 1860
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5397_6
timestamp 1731220340
transform 1 0 744 0 1 1860
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5396_6
timestamp 1731220340
transform 1 0 840 0 1 1860
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5395_6
timestamp 1731220340
transform 1 0 936 0 1 1860
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5394_6
timestamp 1731220340
transform 1 0 1032 0 1 1860
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5393_6
timestamp 1731220340
transform 1 0 1048 0 -1 2012
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5392_6
timestamp 1731220340
transform 1 0 1128 0 1 1860
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5391_6
timestamp 1731220340
transform 1 0 1224 0 -1 2012
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5390_6
timestamp 1731220340
transform 1 0 1248 0 1 2016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5389_6
timestamp 1731220340
transform 1 0 1216 0 -1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5388_6
timestamp 1731220340
transform 1 0 1072 0 -1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5387_6
timestamp 1731220340
transform 1 0 1112 0 1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5386_6
timestamp 1731220340
transform 1 0 952 0 1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5385_6
timestamp 1731220340
transform 1 0 1040 0 -1 2324
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5384_6
timestamp 1731220340
transform 1 0 888 0 -1 2324
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5383_6
timestamp 1731220340
transform 1 0 880 0 1 2324
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5382_6
timestamp 1731220340
transform 1 0 1032 0 1 2324
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5381_6
timestamp 1731220340
transform 1 0 1176 0 1 2324
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5380_6
timestamp 1731220340
transform 1 0 1320 0 1 2324
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5379_6
timestamp 1731220340
transform 1 0 1472 0 1 2324
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5378_6
timestamp 1731220340
transform 1 0 1496 0 -1 2324
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5377_6
timestamp 1731220340
transform 1 0 1344 0 -1 2324
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5376_6
timestamp 1731220340
transform 1 0 1192 0 -1 2324
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5375_6
timestamp 1731220340
transform 1 0 1272 0 1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5374_6
timestamp 1731220340
transform 1 0 1432 0 1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5373_6
timestamp 1731220340
transform 1 0 1592 0 1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5372_6
timestamp 1731220340
transform 1 0 1496 0 -1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5371_6
timestamp 1731220340
transform 1 0 1360 0 -1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5370_6
timestamp 1731220340
transform 1 0 1632 0 -1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5369_6
timestamp 1731220340
transform 1 0 1648 0 1 2016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5368_6
timestamp 1731220340
transform 1 0 1520 0 1 2016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5367_6
timestamp 1731220340
transform 1 0 1384 0 1 2016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5366_6
timestamp 1731220340
transform 1 0 1392 0 -1 2012
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5365_6
timestamp 1731220340
transform 1 0 1568 0 -1 2012
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5364_6
timestamp 1731220340
transform 1 0 1744 0 -1 2012
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5363_6
timestamp 1731220340
transform 1 0 1896 0 -1 2012
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5362_6
timestamp 1731220340
transform 1 0 1896 0 1 2016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5361_6
timestamp 1731220340
transform 1 0 1784 0 1 2016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5360_6
timestamp 1731220340
transform 1 0 1776 0 -1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5359_6
timestamp 1731220340
transform 1 0 1896 0 -1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5358_6
timestamp 1731220340
transform 1 0 2064 0 -1 2228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5357_6
timestamp 1731220340
transform 1 0 2168 0 -1 2228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5356_6
timestamp 1731220340
transform 1 0 2160 0 1 2228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5355_6
timestamp 1731220340
transform 1 0 2064 0 1 2228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5354_6
timestamp 1731220340
transform 1 0 2264 0 1 2228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5353_6
timestamp 1731220340
transform 1 0 2408 0 1 2228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5352_6
timestamp 1731220340
transform 1 0 2568 0 1 2228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5351_6
timestamp 1731220340
transform 1 0 2736 0 1 2228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5350_6
timestamp 1731220340
transform 1 0 2616 0 -1 2228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5349_6
timestamp 1731220340
transform 1 0 2464 0 -1 2228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5348_6
timestamp 1731220340
transform 1 0 2312 0 -1 2228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5347_6
timestamp 1731220340
transform 1 0 2272 0 1 2056
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5346_6
timestamp 1731220340
transform 1 0 2384 0 1 2056
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5345_6
timestamp 1731220340
transform 1 0 2504 0 1 2056
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5344_6
timestamp 1731220340
transform 1 0 2424 0 -1 2048
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5343_6
timestamp 1731220340
transform 1 0 2320 0 -1 2048
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5342_6
timestamp 1731220340
transform 1 0 2528 0 -1 2048
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5341_6
timestamp 1731220340
transform 1 0 2536 0 1 1892
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5340_6
timestamp 1731220340
transform 1 0 2440 0 1 1892
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5339_6
timestamp 1731220340
transform 1 0 2344 0 1 1892
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5338_6
timestamp 1731220340
transform 1 0 2248 0 1 1892
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5337_6
timestamp 1731220340
transform 1 0 2480 0 -1 1880
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5336_6
timestamp 1731220340
transform 1 0 2376 0 -1 1880
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5335_6
timestamp 1731220340
transform 1 0 2272 0 -1 1880
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5334_6
timestamp 1731220340
transform 1 0 2176 0 -1 1880
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5333_6
timestamp 1731220340
transform 1 0 2120 0 1 1724
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5332_6
timestamp 1731220340
transform 1 0 2304 0 1 1724
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5331_6
timestamp 1731220340
transform 1 0 2488 0 1 1724
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5330_6
timestamp 1731220340
transform 1 0 2504 0 -1 1720
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5329_6
timestamp 1731220340
transform 1 0 2336 0 -1 1720
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5328_6
timestamp 1731220340
transform 1 0 2184 0 -1 1720
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5327_6
timestamp 1731220340
transform 1 0 2064 0 -1 1720
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5326_6
timestamp 1731220340
transform 1 0 2328 0 1 1568
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5325_6
timestamp 1731220340
transform 1 0 2064 0 1 1568
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5324_6
timestamp 1731220340
transform 1 0 1896 0 1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5323_6
timestamp 1731220340
transform 1 0 1776 0 1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5322_6
timestamp 1731220340
transform 1 0 1632 0 1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5321_6
timestamp 1731220340
transform 1 0 1488 0 1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5320_6
timestamp 1731220340
transform 1 0 1616 0 -1 1704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5319_6
timestamp 1731220340
transform 1 0 1832 0 -1 1704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5318_6
timestamp 1731220340
transform 1 0 1736 0 1 1704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5317_6
timestamp 1731220340
transform 1 0 1552 0 1 1704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5316_6
timestamp 1731220340
transform 1 0 1376 0 1 1704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5315_6
timestamp 1731220340
transform 1 0 1392 0 -1 1860
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5314_6
timestamp 1731220340
transform 1 0 1528 0 -1 1860
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5313_6
timestamp 1731220340
transform 1 0 1416 0 1 1860
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5312_6
timestamp 1731220340
transform 1 0 1320 0 1 1860
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5311_6
timestamp 1731220340
transform 1 0 1224 0 1 1860
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5310_6
timestamp 1731220340
transform 1 0 1256 0 -1 1860
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5309_6
timestamp 1731220340
transform 1 0 1120 0 -1 1860
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5308_6
timestamp 1731220340
transform 1 0 984 0 -1 1860
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5307_6
timestamp 1731220340
transform 1 0 1200 0 1 1704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5306_6
timestamp 1731220340
transform 1 0 1024 0 1 1704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5305_6
timestamp 1731220340
transform 1 0 992 0 -1 1704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5304_6
timestamp 1731220340
transform 1 0 1400 0 -1 1704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5303_6
timestamp 1731220340
transform 1 0 1192 0 -1 1704
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5302_6
timestamp 1731220340
transform 1 0 1176 0 1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5301_6
timestamp 1731220340
transform 1 0 1008 0 1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5300_6
timestamp 1731220340
transform 1 0 1336 0 1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5299_6
timestamp 1731220340
transform 1 0 1256 0 -1 1548
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5298_6
timestamp 1731220340
transform 1 0 1072 0 -1 1548
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5297_6
timestamp 1731220340
transform 1 0 1440 0 -1 1548
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5296_6
timestamp 1731220340
transform 1 0 1616 0 -1 1548
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5295_6
timestamp 1731220340
transform 1 0 1800 0 -1 1548
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5294_6
timestamp 1731220340
transform 1 0 1896 0 1 1396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5293_6
timestamp 1731220340
transform 1 0 1688 0 1 1396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5292_6
timestamp 1731220340
transform 1 0 1456 0 1 1396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5291_6
timestamp 1731220340
transform 1 0 1744 0 -1 1396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5290_6
timestamp 1731220340
transform 1 0 1896 0 -1 1396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5289_6
timestamp 1731220340
transform 1 0 2064 0 -1 1392
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5288_6
timestamp 1731220340
transform 1 0 2296 0 -1 1392
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5287_6
timestamp 1731220340
transform 1 0 2216 0 1 1232
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5286_6
timestamp 1731220340
transform 1 0 2064 0 1 1232
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5285_6
timestamp 1731220340
transform 1 0 2408 0 1 1232
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5284_6
timestamp 1731220340
transform 1 0 2808 0 1 1232
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5283_6
timestamp 1731220340
transform 1 0 2608 0 1 1232
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5282_6
timestamp 1731220340
transform 1 0 2496 0 -1 1224
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5281_6
timestamp 1731220340
transform 1 0 2304 0 -1 1224
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5280_6
timestamp 1731220340
transform 1 0 2128 0 -1 1224
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5279_6
timestamp 1731220340
transform 1 0 2688 0 -1 1224
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5278_6
timestamp 1731220340
transform 1 0 2880 0 -1 1224
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5277_6
timestamp 1731220340
transform 1 0 2832 0 1 1064
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5276_6
timestamp 1731220340
transform 1 0 2688 0 1 1064
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5275_6
timestamp 1731220340
transform 1 0 2552 0 1 1064
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5274_6
timestamp 1731220340
transform 1 0 2416 0 1 1064
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5273_6
timestamp 1731220340
transform 1 0 2288 0 1 1064
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5272_6
timestamp 1731220340
transform 1 0 2488 0 -1 1060
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5271_6
timestamp 1731220340
transform 1 0 2592 0 -1 1060
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5270_6
timestamp 1731220340
transform 1 0 2704 0 -1 1060
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5269_6
timestamp 1731220340
transform 1 0 2840 0 -1 1060
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5268_6
timestamp 1731220340
transform 1 0 2840 0 1 908
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5267_6
timestamp 1731220340
transform 1 0 2736 0 1 908
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5266_6
timestamp 1731220340
transform 1 0 2640 0 1 908
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5265_6
timestamp 1731220340
transform 1 0 2672 0 -1 896
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5264_6
timestamp 1731220340
transform 1 0 2888 0 -1 896
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5263_6
timestamp 1731220340
transform 1 0 2888 0 1 744
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5262_6
timestamp 1731220340
transform 1 0 3056 0 1 744
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5261_6
timestamp 1731220340
transform 1 0 3056 0 -1 740
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5260_6
timestamp 1731220340
transform 1 0 3120 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5259_6
timestamp 1731220340
transform 1 0 2936 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5258_6
timestamp 1731220340
transform 1 0 2872 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5257_6
timestamp 1731220340
transform 1 0 3064 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5256_6
timestamp 1731220340
transform 1 0 3256 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5255_6
timestamp 1731220340
transform 1 0 3152 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5254_6
timestamp 1731220340
transform 1 0 2952 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5253_6
timestamp 1731220340
transform 1 0 3360 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5252_6
timestamp 1731220340
transform 1 0 3576 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5251_6
timestamp 1731220340
transform 1 0 3408 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5250_6
timestamp 1731220340
transform 1 0 3256 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5249_6
timestamp 1731220340
transform 1 0 3104 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5248_6
timestamp 1731220340
transform 1 0 3552 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5247_6
timestamp 1731220340
transform 1 0 3704 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5246_6
timestamp 1731220340
transform 1 0 3704 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5245_6
timestamp 1731220340
transform 1 0 3800 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5244_6
timestamp 1731220340
transform 1 0 3832 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5243_6
timestamp 1731220340
transform 1 0 3832 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5242_6
timestamp 1731220340
transform 1 0 3832 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5241_6
timestamp 1731220340
transform 1 0 3832 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5240_6
timestamp 1731220340
transform 1 0 3688 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5239_6
timestamp 1731220340
transform 1 0 3560 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5238_6
timestamp 1731220340
transform 1 0 3416 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5237_6
timestamp 1731220340
transform 1 0 3264 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5236_6
timestamp 1731220340
transform 1 0 3664 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5235_6
timestamp 1731220340
transform 1 0 3472 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5234_6
timestamp 1731220340
transform 1 0 3280 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5233_6
timestamp 1731220340
transform 1 0 3088 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5232_6
timestamp 1731220340
transform 1 0 3528 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5231_6
timestamp 1731220340
transform 1 0 3376 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5230_6
timestamp 1731220340
transform 1 0 3232 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5229_6
timestamp 1731220340
transform 1 0 3096 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5228_6
timestamp 1731220340
transform 1 0 2968 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5227_6
timestamp 1731220340
transform 1 0 2856 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5226_6
timestamp 1731220340
transform 1 0 2752 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5225_6
timestamp 1731220340
transform 1 0 2648 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5224_6
timestamp 1731220340
transform 1 0 2488 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5223_6
timestamp 1731220340
transform 1 0 2696 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5222_6
timestamp 1731220340
transform 1 0 2896 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5221_6
timestamp 1731220340
transform 1 0 3112 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5220_6
timestamp 1731220340
transform 1 0 2952 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5219_6
timestamp 1731220340
transform 1 0 2792 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5218_6
timestamp 1731220340
transform 1 0 2632 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5217_6
timestamp 1731220340
transform 1 0 2488 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5216_6
timestamp 1731220340
transform 1 0 2952 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5215_6
timestamp 1731220340
transform 1 0 2792 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5214_6
timestamp 1731220340
transform 1 0 2632 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5213_6
timestamp 1731220340
transform 1 0 2480 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5212_6
timestamp 1731220340
transform 1 0 2336 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5211_6
timestamp 1731220340
transform 1 0 2768 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5210_6
timestamp 1731220340
transform 1 0 2608 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5209_6
timestamp 1731220340
transform 1 0 2456 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5208_6
timestamp 1731220340
transform 1 0 2312 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5207_6
timestamp 1731220340
transform 1 0 2176 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5206_6
timestamp 1731220340
transform 1 0 2680 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5205_6
timestamp 1731220340
transform 1 0 2496 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5204_6
timestamp 1731220340
transform 1 0 2328 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5203_6
timestamp 1731220340
transform 1 0 2176 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5202_6
timestamp 1731220340
transform 1 0 2064 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5201_6
timestamp 1731220340
transform 1 0 2104 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5200_6
timestamp 1731220340
transform 1 0 2240 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5199_6
timestamp 1731220340
transform 1 0 2392 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5198_6
timestamp 1731220340
transform 1 0 2752 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5197_6
timestamp 1731220340
transform 1 0 2568 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5196_6
timestamp 1731220340
transform 1 0 2488 0 -1 740
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5195_6
timestamp 1731220340
transform 1 0 2368 0 -1 740
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5194_6
timestamp 1731220340
transform 1 0 2616 0 -1 740
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5193_6
timestamp 1731220340
transform 1 0 2904 0 -1 740
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5192_6
timestamp 1731220340
transform 1 0 2760 0 -1 740
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5191_6
timestamp 1731220340
transform 1 0 2728 0 1 744
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5190_6
timestamp 1731220340
transform 1 0 2576 0 1 744
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5189_6
timestamp 1731220340
transform 1 0 2440 0 1 744
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5188_6
timestamp 1731220340
transform 1 0 2320 0 1 744
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5187_6
timestamp 1731220340
transform 1 0 2208 0 1 744
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5186_6
timestamp 1731220340
transform 1 0 2456 0 -1 896
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5185_6
timestamp 1731220340
transform 1 0 2248 0 -1 896
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5184_6
timestamp 1731220340
transform 1 0 2064 0 -1 896
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5183_6
timestamp 1731220340
transform 1 0 1896 0 -1 920
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5182_6
timestamp 1731220340
transform 1 0 1744 0 -1 920
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5181_6
timestamp 1731220340
transform 1 0 1896 0 1 920
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5180_6
timestamp 1731220340
transform 1 0 1768 0 1 920
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5179_6
timestamp 1731220340
transform 1 0 1624 0 1 920
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5178_6
timestamp 1731220340
transform 1 0 1480 0 1 920
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5177_6
timestamp 1731220340
transform 1 0 1640 0 -1 1072
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5176_6
timestamp 1731220340
transform 1 0 1824 0 -1 1072
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5175_6
timestamp 1731220340
transform 1 0 1744 0 1 1080
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5174_6
timestamp 1731220340
transform 1 0 1560 0 1 1080
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5173_6
timestamp 1731220340
transform 1 0 1704 0 -1 1236
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5172_6
timestamp 1731220340
transform 1 0 1552 0 -1 1236
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5171_6
timestamp 1731220340
transform 1 0 1400 0 -1 1236
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5170_6
timestamp 1731220340
transform 1 0 1432 0 1 1236
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5169_6
timestamp 1731220340
transform 1 0 1552 0 1 1236
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5168_6
timestamp 1731220340
transform 1 0 1576 0 -1 1396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5167_6
timestamp 1731220340
transform 1 0 1320 0 1 1236
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5166_6
timestamp 1731220340
transform 1 0 1208 0 1 1236
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5165_6
timestamp 1731220340
transform 1 0 1104 0 -1 1236
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5164_6
timestamp 1731220340
transform 1 0 1248 0 -1 1236
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5163_6
timestamp 1731220340
transform 1 0 1200 0 1 1080
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5162_6
timestamp 1731220340
transform 1 0 1376 0 1 1080
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5161_6
timestamp 1731220340
transform 1 0 1456 0 -1 1072
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5160_6
timestamp 1731220340
transform 1 0 1272 0 -1 1072
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5159_6
timestamp 1731220340
transform 1 0 1328 0 1 920
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5158_6
timestamp 1731220340
transform 1 0 1168 0 1 920
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5157_6
timestamp 1731220340
transform 1 0 1232 0 -1 920
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5156_6
timestamp 1731220340
transform 1 0 1408 0 -1 920
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5155_6
timestamp 1731220340
transform 1 0 1576 0 -1 920
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5154_6
timestamp 1731220340
transform 1 0 1528 0 1 768
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5153_6
timestamp 1731220340
transform 1 0 1352 0 1 768
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5152_6
timestamp 1731220340
transform 1 0 1712 0 1 768
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5151_6
timestamp 1731220340
transform 1 0 1592 0 -1 768
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5150_6
timestamp 1731220340
transform 1 0 1448 0 -1 768
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5149_6
timestamp 1731220340
transform 1 0 1304 0 -1 768
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5148_6
timestamp 1731220340
transform 1 0 1288 0 1 616
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5147_6
timestamp 1731220340
transform 1 0 1400 0 1 616
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5146_6
timestamp 1731220340
transform 1 0 1512 0 1 616
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5145_6
timestamp 1731220340
transform 1 0 1448 0 -1 616
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5144_6
timestamp 1731220340
transform 1 0 1352 0 -1 616
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5143_6
timestamp 1731220340
transform 1 0 1256 0 -1 616
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5142_6
timestamp 1731220340
transform 1 0 1160 0 -1 616
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5141_6
timestamp 1731220340
transform 1 0 1064 0 1 616
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5140_6
timestamp 1731220340
transform 1 0 1176 0 1 616
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5139_6
timestamp 1731220340
transform 1 0 1160 0 -1 768
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5138_6
timestamp 1731220340
transform 1 0 1016 0 -1 768
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5137_6
timestamp 1731220340
transform 1 0 1000 0 1 768
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5136_6
timestamp 1731220340
transform 1 0 1176 0 1 768
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5135_6
timestamp 1731220340
transform 1 0 1048 0 -1 920
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5134_6
timestamp 1731220340
transform 1 0 1000 0 1 920
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5133_6
timestamp 1731220340
transform 1 0 1088 0 -1 1072
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5132_6
timestamp 1731220340
transform 1 0 1024 0 1 1080
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5131_6
timestamp 1731220340
transform 1 0 1096 0 1 1236
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5130_6
timestamp 1731220340
transform 1 0 1416 0 -1 1396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5129_6
timestamp 1731220340
transform 1 0 1256 0 -1 1396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5128_6
timestamp 1731220340
transform 1 0 1112 0 -1 1396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5127_6
timestamp 1731220340
transform 1 0 976 0 -1 1396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5126_6
timestamp 1731220340
transform 1 0 1224 0 1 1396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5125_6
timestamp 1731220340
transform 1 0 1000 0 1 1396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5124_6
timestamp 1731220340
transform 1 0 848 0 -1 1396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5123_6
timestamp 1731220340
transform 1 0 720 0 -1 1396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5122_6
timestamp 1731220340
transform 1 0 592 0 -1 1396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5121_6
timestamp 1731220340
transform 1 0 456 0 -1 1396
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5120_6
timestamp 1731220340
transform 1 0 984 0 1 1236
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5119_6
timestamp 1731220340
transform 1 0 872 0 1 1236
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5118_6
timestamp 1731220340
transform 1 0 760 0 1 1236
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5117_6
timestamp 1731220340
transform 1 0 648 0 1 1236
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5116_6
timestamp 1731220340
transform 1 0 544 0 1 1236
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5115_6
timestamp 1731220340
transform 1 0 952 0 -1 1236
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5114_6
timestamp 1731220340
transform 1 0 800 0 -1 1236
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5113_6
timestamp 1731220340
transform 1 0 656 0 -1 1236
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5112_6
timestamp 1731220340
transform 1 0 512 0 -1 1236
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5111_6
timestamp 1731220340
transform 1 0 384 0 -1 1236
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5110_6
timestamp 1731220340
transform 1 0 840 0 1 1080
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5109_6
timestamp 1731220340
transform 1 0 664 0 1 1080
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5108_6
timestamp 1731220340
transform 1 0 488 0 1 1080
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5107_6
timestamp 1731220340
transform 1 0 320 0 1 1080
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5106_6
timestamp 1731220340
transform 1 0 168 0 1 1080
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5105_6
timestamp 1731220340
transform 1 0 904 0 -1 1072
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5104_6
timestamp 1731220340
transform 1 0 720 0 -1 1072
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5103_6
timestamp 1731220340
transform 1 0 536 0 -1 1072
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5102_6
timestamp 1731220340
transform 1 0 368 0 -1 1072
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5101_6
timestamp 1731220340
transform 1 0 224 0 -1 1072
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5100_6
timestamp 1731220340
transform 1 0 128 0 -1 1072
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_599_6
timestamp 1731220340
transform 1 0 128 0 1 920
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_598_6
timestamp 1731220340
transform 1 0 264 0 1 920
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_597_6
timestamp 1731220340
transform 1 0 440 0 1 920
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_596_6
timestamp 1731220340
transform 1 0 624 0 1 920
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_595_6
timestamp 1731220340
transform 1 0 816 0 1 920
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_594_6
timestamp 1731220340
transform 1 0 848 0 -1 920
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_593_6
timestamp 1731220340
transform 1 0 648 0 -1 920
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_592_6
timestamp 1731220340
transform 1 0 448 0 -1 920
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_591_6
timestamp 1731220340
transform 1 0 264 0 -1 920
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_590_6
timestamp 1731220340
transform 1 0 128 0 -1 920
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_589_6
timestamp 1731220340
transform 1 0 208 0 1 768
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_588_6
timestamp 1731220340
transform 1 0 336 0 1 768
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_587_6
timestamp 1731220340
transform 1 0 488 0 1 768
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_586_6
timestamp 1731220340
transform 1 0 648 0 1 768
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_585_6
timestamp 1731220340
transform 1 0 824 0 1 768
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_584_6
timestamp 1731220340
transform 1 0 880 0 -1 768
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_583_6
timestamp 1731220340
transform 1 0 616 0 -1 768
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_582_6
timestamp 1731220340
transform 1 0 488 0 -1 768
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_581_6
timestamp 1731220340
transform 1 0 368 0 -1 768
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_580_6
timestamp 1731220340
transform 1 0 744 0 -1 768
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_579_6
timestamp 1731220340
transform 1 0 736 0 1 616
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_578_6
timestamp 1731220340
transform 1 0 624 0 1 616
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_577_6
timestamp 1731220340
transform 1 0 520 0 1 616
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_576_6
timestamp 1731220340
transform 1 0 848 0 1 616
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_575_6
timestamp 1731220340
transform 1 0 960 0 1 616
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_574_6
timestamp 1731220340
transform 1 0 872 0 -1 616
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_573_6
timestamp 1731220340
transform 1 0 776 0 -1 616
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_572_6
timestamp 1731220340
transform 1 0 680 0 -1 616
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_571_6
timestamp 1731220340
transform 1 0 968 0 -1 616
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_570_6
timestamp 1731220340
transform 1 0 1064 0 -1 616
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_569_6
timestamp 1731220340
transform 1 0 1336 0 1 444
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_568_6
timestamp 1731220340
transform 1 0 1528 0 1 444
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_567_6
timestamp 1731220340
transform 1 0 1432 0 1 444
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_566_6
timestamp 1731220340
transform 1 0 1424 0 -1 432
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_565_6
timestamp 1731220340
transform 1 0 1312 0 -1 432
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_564_6
timestamp 1731220340
transform 1 0 1344 0 1 276
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_563_6
timestamp 1731220340
transform 1 0 1488 0 1 276
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_562_6
timestamp 1731220340
transform 1 0 1632 0 1 276
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_561_6
timestamp 1731220340
transform 1 0 1504 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_560_6
timestamp 1731220340
transform 1 0 1640 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_559_6
timestamp 1731220340
transform 1 0 1776 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_558_6
timestamp 1731220340
transform 1 0 1896 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_557_6
timestamp 1731220340
transform 1 0 2064 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_556_6
timestamp 1731220340
transform 1 0 2264 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_555_6
timestamp 1731220340
transform 1 0 2544 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_554_6
timestamp 1731220340
transform 1 0 2448 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_553_6
timestamp 1731220340
transform 1 0 2352 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_552_6
timestamp 1731220340
transform 1 0 2256 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_551_6
timestamp 1731220340
transform 1 0 2160 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_550_6
timestamp 1731220340
transform 1 0 2064 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_549_6
timestamp 1731220340
transform 1 0 1896 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_548_6
timestamp 1731220340
transform 1 0 1800 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_547_6
timestamp 1731220340
transform 1 0 1696 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_546_6
timestamp 1731220340
transform 1 0 1584 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_545_6
timestamp 1731220340
transform 1 0 1480 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_544_6
timestamp 1731220340
transform 1 0 1376 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_543_6
timestamp 1731220340
transform 1 0 1264 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_542_6
timestamp 1731220340
transform 1 0 1144 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_541_6
timestamp 1731220340
transform 1 0 1024 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_540_6
timestamp 1731220340
transform 1 0 1040 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_539_6
timestamp 1731220340
transform 1 0 1360 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_538_6
timestamp 1731220340
transform 1 0 1208 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_537_6
timestamp 1731220340
transform 1 0 1200 0 1 276
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_536_6
timestamp 1731220340
transform 1 0 1056 0 1 276
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_535_6
timestamp 1731220340
transform 1 0 992 0 -1 432
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_534_6
timestamp 1731220340
transform 1 0 1096 0 -1 432
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_533_6
timestamp 1731220340
transform 1 0 1200 0 -1 432
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_532_6
timestamp 1731220340
transform 1 0 1240 0 1 444
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_531_6
timestamp 1731220340
transform 1 0 1144 0 1 444
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_530_6
timestamp 1731220340
transform 1 0 1048 0 1 444
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_529_6
timestamp 1731220340
transform 1 0 952 0 1 444
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_528_6
timestamp 1731220340
transform 1 0 856 0 1 444
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_527_6
timestamp 1731220340
transform 1 0 760 0 1 444
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_526_6
timestamp 1731220340
transform 1 0 664 0 1 444
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_525_6
timestamp 1731220340
transform 1 0 568 0 1 444
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_524_6
timestamp 1731220340
transform 1 0 472 0 1 444
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_523_6
timestamp 1731220340
transform 1 0 376 0 1 444
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_522_6
timestamp 1731220340
transform 1 0 888 0 -1 432
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_521_6
timestamp 1731220340
transform 1 0 784 0 -1 432
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_520_6
timestamp 1731220340
transform 1 0 680 0 -1 432
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_519_6
timestamp 1731220340
transform 1 0 576 0 -1 432
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_518_6
timestamp 1731220340
transform 1 0 480 0 -1 432
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_517_6
timestamp 1731220340
transform 1 0 912 0 1 276
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_516_6
timestamp 1731220340
transform 1 0 760 0 1 276
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_515_6
timestamp 1731220340
transform 1 0 608 0 1 276
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_514_6
timestamp 1731220340
transform 1 0 456 0 1 276
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_513_6
timestamp 1731220340
transform 1 0 320 0 1 276
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_512_6
timestamp 1731220340
transform 1 0 864 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_511_6
timestamp 1731220340
transform 1 0 680 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_510_6
timestamp 1731220340
transform 1 0 496 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_59_6
timestamp 1731220340
transform 1 0 320 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_58_6
timestamp 1731220340
transform 1 0 160 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_57_6
timestamp 1731220340
transform 1 0 896 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_56_6
timestamp 1731220340
transform 1 0 768 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_55_6
timestamp 1731220340
transform 1 0 640 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_54_6
timestamp 1731220340
transform 1 0 520 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_53_6
timestamp 1731220340
transform 1 0 416 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_52_6
timestamp 1731220340
transform 1 0 320 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_51_6
timestamp 1731220340
transform 1 0 224 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_50_6
timestamp 1731220340
transform 1 0 128 0 1 88
box 8 5 92 72
<< end >>
