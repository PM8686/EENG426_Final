magic
tech sky130l
timestamp 1731220306
<< checkpaint >>
rect -24 32 132 100
rect -24 21 131 32
rect -24 20 121 21
rect -16 -18 121 20
rect -16 -20 116 -18
rect -16 -27 87 -20
<< ndiffusion >>
rect 16 23 21 24
rect 16 20 17 23
rect 20 20 21 23
rect 16 14 21 20
rect 23 18 28 24
rect 23 15 24 18
rect 27 15 28 18
rect 23 14 28 15
rect 30 23 35 24
rect 30 20 31 23
rect 34 20 35 23
rect 30 14 35 20
rect 41 23 46 24
rect 41 20 42 23
rect 45 20 46 23
rect 41 14 46 20
rect 48 18 55 24
rect 48 15 51 18
rect 54 15 55 18
rect 48 14 55 15
rect 57 23 62 24
rect 57 20 58 23
rect 61 20 62 23
rect 57 14 62 20
rect 68 23 73 24
rect 68 20 69 23
rect 72 20 73 23
rect 68 14 73 20
rect 75 18 82 24
rect 75 15 76 18
rect 79 15 82 18
rect 75 14 82 15
rect 84 23 89 24
rect 84 20 85 23
rect 88 20 89 23
rect 84 14 89 20
<< ndc >>
rect 17 20 20 23
rect 24 15 27 18
rect 31 20 34 23
rect 42 20 45 23
rect 51 15 54 18
rect 58 20 61 23
rect 69 20 72 23
rect 76 15 79 18
rect 85 20 88 23
<< ntransistor >>
rect 21 14 23 24
rect 28 14 30 24
rect 46 14 48 24
rect 55 14 57 24
rect 73 14 75 24
rect 82 14 84 24
<< pdiffusion >>
rect 16 45 21 46
rect 16 42 17 45
rect 20 42 21 45
rect 16 31 21 42
rect 23 45 28 46
rect 23 42 24 45
rect 27 42 28 45
rect 23 31 28 42
rect 30 45 35 46
rect 30 42 31 45
rect 34 42 35 45
rect 30 31 35 42
rect 51 41 55 51
rect 41 35 46 41
rect 41 32 42 35
rect 45 32 46 35
rect 41 31 46 32
rect 48 35 55 41
rect 48 32 51 35
rect 54 32 55 35
rect 48 31 55 32
rect 57 42 62 51
rect 57 39 58 42
rect 61 39 62 42
rect 78 41 82 51
rect 57 31 62 39
rect 68 35 73 41
rect 68 32 69 35
rect 72 32 73 35
rect 68 31 73 32
rect 75 40 82 41
rect 75 37 78 40
rect 81 37 82 40
rect 75 31 82 37
rect 84 42 89 51
rect 84 39 85 42
rect 88 39 89 42
rect 84 31 89 39
<< pdc >>
rect 17 42 20 45
rect 24 42 27 45
rect 31 42 34 45
rect 42 32 45 35
rect 51 32 54 35
rect 58 39 61 42
rect 69 32 72 35
rect 78 37 81 40
rect 85 39 88 42
<< ptransistor >>
rect 21 31 23 46
rect 28 31 30 46
rect 46 31 48 41
rect 55 31 57 51
rect 73 31 75 41
rect 82 31 84 51
<< polysilicon >>
rect 52 58 57 59
rect 52 55 53 58
rect 56 55 57 58
rect 52 54 57 55
rect 55 51 57 54
rect 82 58 88 59
rect 82 55 84 58
rect 87 55 88 58
rect 82 54 88 55
rect 82 51 84 54
rect 21 46 23 48
rect 28 46 30 48
rect 46 41 48 43
rect 70 49 75 50
rect 70 46 71 49
rect 74 46 75 49
rect 70 45 75 46
rect 73 41 75 45
rect 21 24 23 31
rect 28 24 30 31
rect 46 24 48 31
rect 55 24 57 31
rect 73 24 75 31
rect 82 24 84 31
rect 21 10 23 14
rect 18 9 23 10
rect 18 6 19 9
rect 22 6 23 9
rect 28 12 30 14
rect 46 12 48 14
rect 55 12 57 14
rect 73 12 75 14
rect 82 12 84 14
rect 28 11 34 12
rect 28 8 30 11
rect 33 8 34 11
rect 28 7 34 8
rect 43 11 48 12
rect 43 8 44 11
rect 47 8 48 11
rect 43 7 48 8
rect 18 5 23 6
<< pc >>
rect 53 55 56 58
rect 84 55 87 58
rect 71 46 74 49
rect 19 6 22 9
rect 30 8 33 11
rect 44 8 47 11
<< m1 >>
rect 8 55 12 68
rect 40 64 44 68
rect 96 64 100 68
rect 40 58 43 64
rect 84 58 87 59
rect 8 52 20 55
rect 17 49 20 52
rect 17 45 20 46
rect 17 23 20 42
rect 24 53 25 56
rect 24 45 28 53
rect 27 42 28 45
rect 24 41 28 42
rect 31 55 53 58
rect 56 55 57 58
rect 78 56 81 57
rect 31 45 34 55
rect 96 56 99 64
rect 87 55 99 56
rect 84 53 99 55
rect 70 46 71 49
rect 74 46 75 49
rect 17 19 20 20
rect 31 23 34 42
rect 57 39 58 42
rect 61 39 62 42
rect 78 40 81 53
rect 84 39 85 42
rect 88 39 89 42
rect 78 36 81 37
rect 51 35 54 36
rect 41 32 42 35
rect 45 32 46 35
rect 68 32 69 35
rect 72 32 73 35
rect 41 20 42 23
rect 45 20 46 23
rect 31 19 34 20
rect 24 18 27 19
rect 51 18 54 32
rect 57 20 58 23
rect 61 20 69 23
rect 72 20 73 23
rect 84 20 85 23
rect 88 20 89 23
rect 24 14 27 15
rect 30 12 36 16
rect 76 18 79 19
rect 30 11 48 12
rect 18 6 19 9
rect 22 6 23 9
rect 33 8 44 11
rect 47 8 48 11
rect 51 9 54 15
rect 71 13 72 16
rect 75 15 76 16
rect 75 13 79 15
rect 71 12 79 13
rect 30 7 33 8
rect 51 5 54 6
<< m2c >>
rect 17 46 20 49
rect 25 53 28 56
rect 78 53 81 56
rect 71 46 74 49
rect 58 39 61 42
rect 85 39 88 42
rect 42 32 45 35
rect 69 32 72 35
rect 42 20 45 23
rect 24 15 27 18
rect 85 20 88 23
rect 19 6 22 9
rect 72 13 75 16
rect 51 6 54 9
<< m2 >>
rect 24 56 82 57
rect 24 53 25 56
rect 28 53 78 56
rect 81 53 82 56
rect 24 52 82 53
rect 16 49 75 50
rect 16 46 17 49
rect 20 46 71 49
rect 74 46 75 49
rect 16 45 75 46
rect 57 42 89 43
rect 57 39 58 42
rect 61 39 85 42
rect 88 39 89 42
rect 57 38 89 39
rect 41 35 73 36
rect 41 32 42 35
rect 45 32 69 35
rect 72 32 73 35
rect 41 31 73 32
rect 41 23 89 24
rect 41 20 42 23
rect 45 20 85 23
rect 88 20 89 23
rect 41 19 89 20
rect 23 18 28 19
rect 23 15 24 18
rect 27 17 28 18
rect 27 16 76 17
rect 27 15 72 16
rect 23 13 72 15
rect 75 13 76 16
rect 23 12 76 13
rect 16 9 55 10
rect 16 6 19 9
rect 22 6 51 9
rect 54 6 55 9
rect 16 5 55 6
<< labels >>
rlabel space 0 0 104 72 6 prboundary
rlabel polysilicon 83 25 83 25 3 D
rlabel polysilicon 83 52 83 52 3 D
rlabel polysilicon 83 55 83 55 3 D
rlabel polysilicon 83 56 83 56 3 D
rlabel polysilicon 83 59 83 59 3 D
rlabel ndiffusion 85 15 85 15 3 #5
rlabel ndiffusion 85 24 85 24 3 #5
rlabel ndiffusion 80 16 80 16 3 GND
rlabel pdiffusion 85 32 85 32 3 #7
rlabel pdiffusion 85 43 85 43 3 #7
rlabel pdiffusion 82 38 82 38 3 Vdd
rlabel pdiffusion 79 42 79 42 3 Vdd
rlabel ntransistor 83 15 83 15 3 D
rlabel ptransistor 83 32 83 32 3 D
rlabel ndiffusion 76 15 76 15 3 GND
rlabel ndiffusion 76 19 76 19 3 GND
rlabel ndiffusion 69 21 69 21 3 #10
rlabel pdiffusion 76 32 76 32 3 Vdd
rlabel pdiffusion 76 38 76 38 3 Vdd
rlabel pdiffusion 76 41 76 41 3 Vdd
rlabel polysilicon 74 42 74 42 3 Q
rlabel ntransistor 74 15 74 15 3 Q
rlabel polysilicon 74 25 74 25 3 Q
rlabel ptransistor 74 32 74 32 3 Q
rlabel polysilicon 71 46 71 46 3 Q
rlabel polysilicon 71 50 71 50 3 Q
rlabel polysilicon 83 13 83 13 3 D
rlabel ndiffusion 69 15 69 15 3 #10
rlabel ndiffusion 69 24 69 24 3 #10
rlabel pdiffusion 69 32 69 32 3 #8
rlabel pdiffusion 69 36 69 36 3 #8
rlabel polysilicon 56 25 56 25 3 _clk
rlabel polysilicon 56 52 56 52 3 _clk
rlabel polysilicon 74 13 74 13 3 Q
rlabel ndiffusion 58 15 58 15 3 #10
rlabel ndiffusion 58 24 58 24 3 #10
rlabel ndiffusion 55 16 55 16 3 _q
rlabel pdiffusion 58 32 58 32 3 #7
rlabel pdiffusion 55 33 55 33 3 _q
rlabel polysilicon 53 55 53 55 3 _clk
rlabel polysilicon 53 56 53 56 3 _clk
rlabel polysilicon 53 59 53 59 3 _clk
rlabel polysilicon 44 9 44 9 3 CLK
rlabel ntransistor 56 15 56 15 3 _clk
rlabel ptransistor 56 32 56 32 3 _clk
rlabel pdiffusion 52 42 52 42 3 _q
rlabel polysilicon 56 13 56 13 3 _clk
rlabel ndiffusion 49 15 49 15 3 _q
rlabel ndiffusion 49 16 49 16 3 _q
rlabel ndiffusion 49 19 49 19 3 _q
rlabel pdiffusion 49 32 49 32 3 _q
rlabel pdiffusion 49 33 49 33 3 _q
rlabel pdiffusion 49 36 49 36 3 _q
rlabel polysilicon 44 8 44 8 3 CLK
rlabel ntransistor 47 15 47 15 3 CLK
rlabel polysilicon 47 25 47 25 3 CLK
rlabel ptransistor 47 32 47 32 3 CLK
rlabel polysilicon 47 42 47 42 3 CLK
rlabel polysilicon 44 12 44 12 3 CLK
rlabel polysilicon 47 13 47 13 3 CLK
rlabel ndiffusion 42 15 42 15 3 #5
rlabel ndiffusion 35 21 35 21 3 _clk
rlabel pdiffusion 35 43 35 43 3 _clk
rlabel polysilicon 29 8 29 8 3 CLK
rlabel polysilicon 29 9 29 9 3 CLK
rlabel polysilicon 29 12 29 12 3 CLK
rlabel polysilicon 29 13 29 13 3 CLK
rlabel ndiffusion 31 15 31 15 3 _clk
rlabel ndiffusion 31 21 31 21 3 _clk
rlabel ndiffusion 31 24 31 24 3 _clk
rlabel pdiffusion 31 32 31 32 3 _clk
rlabel pdiffusion 31 43 31 43 3 _clk
rlabel pdiffusion 31 46 31 46 3 _clk
rlabel ntransistor 29 15 29 15 3 CLK
rlabel polysilicon 29 25 29 25 3 CLK
rlabel ptransistor 29 32 29 32 3 CLK
rlabel polysilicon 29 47 29 47 3 CLK
rlabel polysilicon 22 11 22 11 3 _q
rlabel ndiffusion 24 15 24 15 3 GND
rlabel ndiffusion 21 21 21 21 3 Q
rlabel pdiffusion 24 32 24 32 3 Vdd
rlabel pdiffusion 24 43 24 43 3 Vdd
rlabel pdiffusion 24 46 24 46 3 Vdd
rlabel pdiffusion 21 43 21 43 3 Q
rlabel polysilicon 19 6 19 6 3 _q
rlabel polysilicon 19 10 19 10 3 _q
rlabel ntransistor 22 15 22 15 3 _q
rlabel polysilicon 22 25 22 25 3 _q
rlabel ptransistor 22 32 22 32 3 _q
rlabel polysilicon 22 47 22 47 3 _q
rlabel ndiffusion 17 15 17 15 3 Q
rlabel ndiffusion 17 21 17 21 3 Q
rlabel ndiffusion 17 24 17 24 3 Q
rlabel pdiffusion 17 32 17 32 3 Q
rlabel pdiffusion 17 43 17 43 3 Q
rlabel m1 97 57 97 57 3 D
port 1 e
rlabel m1 97 65 97 65 3 D
port 1 e
rlabel m1 88 56 88 56 3 D
port 1 e
rlabel m1 85 40 85 40 3 #7
rlabel m1 85 54 85 54 3 D
port 1 e
rlabel pc 85 56 85 56 3 D
port 1 e
rlabel m1 85 59 85 59 3 D
port 1 e
rlabel m1 79 57 79 57 3 Vdd
rlabel m1 85 21 85 21 3 #5
rlabel m1 79 37 79 37 3 Vdd
rlabel pdc 79 38 79 38 3 Vdd
rlabel m1 79 41 79 41 3 Vdd
rlabel ndc 77 16 77 16 3 GND
rlabel m1 76 16 76 16 3 GND
rlabel m1 71 47 71 47 3 Q
port 2 e
rlabel m1 73 21 73 21 3 #10
rlabel m1 72 13 72 13 3 GND
rlabel m1 72 14 72 14 3 GND
rlabel m1 77 19 77 19 3 GND
rlabel ndc 70 21 70 21 3 #10
rlabel m1 69 33 69 33 3 #8
rlabel m1 62 21 62 21 3 #10
rlabel pdc 52 33 52 33 3 _q
rlabel m1 52 36 52 36 3 _q
rlabel m1 52 10 52 10 3 _q
rlabel ndc 59 21 59 21 3 #10
rlabel m1 58 21 58 21 3 #10
rlabel m1 32 20 32 20 3 _clk
rlabel m1 48 9 48 9 3 CLK
port 3 e
rlabel pc 45 9 45 9 3 CLK
port 3 e
rlabel ndc 52 16 52 16 3 _q
rlabel m1 52 19 52 19 3 _q
rlabel m1 57 56 57 56 3 _clk
rlabel m1 41 59 41 59 3 CLK
port 3 e
rlabel m1 41 65 41 65 3 CLK
port 3 e
rlabel m1 52 6 52 6 3 _q
rlabel m1 34 9 34 9 3 CLK
port 3 e
rlabel m1 25 15 25 15 3 GND
rlabel m1 25 19 25 19 3 GND
rlabel pdc 32 43 32 43 3 _clk
rlabel pc 54 56 54 56 3 _clk
rlabel m1 31 8 31 8 3 CLK
port 3 e
rlabel pc 31 9 31 9 3 CLK
port 3 e
rlabel m1 31 12 31 12 3 CLK
port 3 e
rlabel m1 31 13 31 13 3 CLK
port 3 e
rlabel m1 32 46 32 46 3 _clk
rlabel m1 32 56 32 56 3 _clk
rlabel ndc 32 21 32 21 3 _clk
rlabel m1 32 24 32 24 3 _clk
rlabel m1 28 43 28 43 3 Vdd
rlabel m1 25 42 25 42 3 Vdd
rlabel pdc 25 43 25 43 3 Vdd
rlabel m1 25 46 25 46 3 Vdd
rlabel m1 19 7 19 7 3 _q
rlabel m1 18 20 18 20 3 Q
port 2 e
rlabel ndc 18 21 18 21 3 Q
port 2 e
rlabel m1 18 24 18 24 3 Q
port 2 e
rlabel pdc 18 43 18 43 3 Q
port 2 e
rlabel m1 18 46 18 46 3 Q
port 2 e
rlabel m1 18 50 18 50 3 Q
port 2 e
rlabel m1 9 53 9 53 3 Q
port 2 e
rlabel m1 9 56 9 56 3 Q
port 2 e
rlabel m2 89 40 89 40 3 #7
rlabel m2c 86 40 86 40 3 #7
rlabel m2 62 40 62 40 3 #7
rlabel m2 89 21 89 21 3 #5
rlabel m2 73 33 73 33 3 #8
rlabel m2c 59 40 59 40 3 #7
rlabel m2c 86 21 86 21 3 #5
rlabel m2c 70 33 70 33 3 #8
rlabel m2 58 39 58 39 3 #7
rlabel m2 58 40 58 40 3 #7
rlabel m2 58 43 58 43 3 #7
rlabel m2 46 21 46 21 3 #5
rlabel m2 46 33 46 33 3 #8
rlabel m2c 43 21 43 21 3 #5
rlabel m2c 43 33 43 33 3 #8
rlabel m2 82 54 82 54 3 Vdd
rlabel m2 76 14 76 14 3 GND
rlabel m2 28 16 28 16 3 GND
rlabel m2 28 17 28 17 3 GND
rlabel m2 28 18 28 18 3 GND
rlabel m2 42 20 42 20 3 #5
rlabel m2 42 21 42 21 3 #5
rlabel m2 42 24 42 24 3 #5
rlabel m2 42 32 42 32 3 #8
rlabel m2 42 33 42 33 3 #8
rlabel m2 42 36 42 36 3 #8
rlabel m2c 79 54 79 54 3 Vdd
rlabel m2c 73 14 73 14 3 GND
rlabel m2c 25 16 25 16 3 GND
rlabel m2 29 54 29 54 3 Vdd
rlabel m2 55 7 55 7 3 _q
rlabel m2 24 13 24 13 3 GND
rlabel m2 24 14 24 14 3 GND
rlabel m2 24 16 24 16 3 GND
rlabel m2 24 19 24 19 3 GND
rlabel m2 75 47 75 47 3 Q
port 2 e
rlabel m2c 26 54 26 54 3 Vdd
rlabel m2c 52 7 52 7 3 _q
rlabel m2c 72 47 72 47 3 Q
port 2 e
rlabel m2 25 53 25 53 3 Vdd
rlabel m2 25 54 25 54 3 Vdd
rlabel m2 25 57 25 57 3 Vdd
rlabel m2 23 7 23 7 3 _q
rlabel m2 21 47 21 47 3 Q
port 2 e
rlabel m2c 20 7 20 7 3 _q
rlabel m2c 18 47 18 47 3 Q
port 2 e
rlabel m2 17 6 17 6 3 _q
rlabel m2 17 7 17 7 3 _q
rlabel m2 17 10 17 10 3 _q
rlabel m2 17 46 17 46 3 Q
port 2 e
rlabel m2 17 47 17 47 3 Q
port 2 e
rlabel m2 17 50 17 50 3 Q
port 2 e
<< end >>
