magic
tech sky130l
timestamp 1730254909
<< ndiffusion >>
rect 8 11 13 16
rect 8 8 9 11
rect 12 8 13 11
rect 8 6 13 8
rect 15 6 20 16
rect 22 14 27 16
rect 22 11 23 14
rect 26 11 27 14
rect 22 6 27 11
rect 33 15 38 16
rect 33 12 34 15
rect 37 12 38 15
rect 33 10 38 12
rect 40 14 47 16
rect 40 11 41 14
rect 44 11 47 14
rect 40 10 47 11
rect 43 6 47 10
rect 49 11 54 16
rect 49 8 50 11
rect 53 8 54 11
rect 49 6 54 8
rect 60 14 65 16
rect 60 11 61 14
rect 64 11 65 14
rect 60 6 65 11
rect 67 11 72 16
rect 67 8 68 11
rect 71 8 72 11
rect 67 6 72 8
<< ndc >>
rect 9 8 12 11
rect 23 11 26 14
rect 34 12 37 15
rect 41 11 44 14
rect 50 8 53 11
rect 61 11 64 14
rect 68 8 71 11
<< ntransistor >>
rect 13 6 15 16
rect 20 6 22 16
rect 38 10 40 16
rect 47 6 49 16
rect 65 6 67 16
<< pdiffusion >>
rect 8 35 13 38
rect 8 32 9 35
rect 12 32 13 35
rect 8 23 13 32
rect 15 31 19 38
rect 15 30 20 31
rect 15 27 16 30
rect 19 27 20 30
rect 15 23 20 27
rect 22 27 27 31
rect 22 24 23 27
rect 26 24 27 27
rect 22 23 27 24
rect 33 28 38 38
rect 33 25 34 28
rect 37 25 38 28
rect 33 23 38 25
rect 40 23 47 38
rect 49 37 54 38
rect 49 34 50 37
rect 53 34 54 37
rect 49 23 54 34
rect 60 35 65 38
rect 60 32 61 35
rect 64 32 65 35
rect 60 23 65 32
rect 67 28 72 38
rect 67 25 68 28
rect 71 25 72 28
rect 67 23 72 25
<< pdc >>
rect 9 32 12 35
rect 16 27 19 30
rect 23 24 26 27
rect 34 25 37 28
rect 50 34 53 37
rect 61 32 64 35
rect 68 25 71 28
<< ptransistor >>
rect 13 23 15 38
rect 20 23 22 31
rect 38 23 40 38
rect 47 23 49 38
rect 65 23 67 38
<< polysilicon >>
rect 9 45 15 46
rect 9 42 10 45
rect 13 42 15 45
rect 9 41 15 42
rect 32 45 40 46
rect 32 42 33 45
rect 36 42 40 45
rect 32 41 40 42
rect 43 45 49 46
rect 43 42 44 45
rect 47 42 49 45
rect 43 41 49 42
rect 13 38 15 41
rect 20 38 28 39
rect 38 38 40 41
rect 47 38 49 41
rect 65 38 67 40
rect 20 35 24 38
rect 27 35 28 38
rect 20 34 28 35
rect 20 31 22 34
rect 13 16 15 23
rect 20 16 22 23
rect 38 16 40 23
rect 47 16 49 23
rect 65 22 67 23
rect 65 21 80 22
rect 65 20 76 21
rect 65 16 67 20
rect 75 18 76 20
rect 79 18 80 21
rect 75 17 80 18
rect 38 8 40 10
rect 13 4 15 6
rect 20 4 22 6
rect 47 4 49 6
rect 65 4 67 6
<< pc >>
rect 10 42 13 45
rect 33 42 36 45
rect 44 42 47 45
rect 24 35 27 38
rect 76 18 79 21
<< m1 >>
rect 8 45 13 46
rect 8 42 10 45
rect 8 40 13 42
rect 16 42 20 44
rect 19 40 20 42
rect 24 42 33 45
rect 36 42 37 45
rect 24 41 37 42
rect 8 32 9 35
rect 12 32 13 35
rect 16 30 19 39
rect 24 38 28 41
rect 40 40 44 45
rect 47 42 48 45
rect 51 42 54 43
rect 27 35 28 38
rect 51 37 54 39
rect 24 34 28 35
rect 49 34 50 37
rect 53 34 54 37
rect 60 32 61 35
rect 64 32 65 35
rect 56 28 60 29
rect 16 26 19 27
rect 23 27 26 28
rect 33 25 34 28
rect 37 25 38 28
rect 59 25 60 28
rect 67 25 68 28
rect 71 25 72 28
rect 23 21 26 24
rect 23 17 26 18
rect 34 21 37 22
rect 34 15 37 18
rect 56 15 60 25
rect 75 18 76 21
rect 79 18 80 21
rect 8 11 12 12
rect 22 11 23 14
rect 26 11 27 14
rect 34 11 37 12
rect 41 14 44 15
rect 56 14 64 15
rect 8 8 9 11
rect 8 7 12 8
rect 8 4 9 7
rect 8 3 12 4
rect 41 7 44 11
rect 41 3 44 4
rect 50 11 53 12
rect 50 7 53 8
rect 56 11 61 14
rect 56 10 64 11
rect 68 11 71 12
rect 56 4 60 10
rect 68 7 71 8
rect 50 3 53 4
rect 68 3 71 4
<< m2c >>
rect 16 39 19 42
rect 9 32 12 35
rect 51 39 54 42
rect 61 32 64 35
rect 34 25 37 28
rect 56 25 59 28
rect 68 25 71 28
rect 23 18 26 21
rect 34 18 37 21
rect 76 18 79 21
rect 23 11 26 14
rect 9 4 12 7
rect 41 4 44 7
rect 50 4 53 7
rect 61 11 64 14
rect 68 4 71 7
<< m2 >>
rect 15 42 55 43
rect 15 39 16 42
rect 19 39 51 42
rect 54 39 55 42
rect 15 38 55 39
rect 8 35 65 36
rect 8 32 9 35
rect 12 32 61 35
rect 64 32 65 35
rect 8 31 65 32
rect 33 28 72 29
rect 33 25 34 28
rect 37 25 56 28
rect 59 25 68 28
rect 71 25 72 28
rect 33 24 72 25
rect 22 21 80 22
rect 22 18 23 21
rect 26 18 34 21
rect 37 18 76 21
rect 79 18 80 21
rect 22 17 80 18
rect 22 14 65 15
rect 22 11 23 14
rect 26 11 61 14
rect 64 11 65 14
rect 22 10 65 11
rect 8 7 46 8
rect 8 4 9 7
rect 12 4 41 7
rect 44 4 46 7
rect 8 3 46 4
rect 49 7 72 8
rect 49 4 50 7
rect 53 4 68 7
rect 71 4 72 7
rect 49 3 72 4
<< labels >>
rlabel m1 s 10 42 13 45 6 A
port 1 nsew signal input
rlabel m1 s 8 40 13 42 6 A
port 1 nsew signal input
rlabel m1 s 8 42 10 45 6 A
port 1 nsew signal input
rlabel m1 s 8 45 13 46 6 A
port 1 nsew signal input
rlabel m1 s 47 42 48 45 6 B
port 2 nsew signal input
rlabel m1 s 44 42 47 45 6 B
port 2 nsew signal input
rlabel m1 s 40 40 44 45 6 B
port 2 nsew signal input
rlabel m1 s 36 42 37 45 6 S
port 3 nsew signal input
rlabel m1 s 27 35 28 38 6 S
port 3 nsew signal input
rlabel m1 s 33 42 36 45 6 S
port 3 nsew signal input
rlabel m1 s 24 34 28 35 6 S
port 3 nsew signal input
rlabel m1 s 24 35 27 38 6 S
port 3 nsew signal input
rlabel m1 s 24 38 28 41 6 S
port 3 nsew signal input
rlabel m1 s 24 41 37 42 6 S
port 3 nsew signal input
rlabel m1 s 24 42 33 45 6 S
port 3 nsew signal input
rlabel m2 s 71 25 72 28 6 Y
port 4 nsew signal output
rlabel m2 s 68 25 71 28 6 Y
port 4 nsew signal output
rlabel m2 s 59 25 68 28 6 Y
port 4 nsew signal output
rlabel m2 s 56 25 59 28 6 Y
port 4 nsew signal output
rlabel m2 s 37 25 56 28 6 Y
port 4 nsew signal output
rlabel m2 s 64 11 65 14 6 Y
port 4 nsew signal output
rlabel m2 s 34 25 37 28 6 Y
port 4 nsew signal output
rlabel m2 s 61 11 64 14 6 Y
port 4 nsew signal output
rlabel m2 s 33 24 72 25 6 Y
port 4 nsew signal output
rlabel m2 s 33 25 34 28 6 Y
port 4 nsew signal output
rlabel m2 s 33 28 72 29 6 Y
port 4 nsew signal output
rlabel m2 s 26 11 61 14 6 Y
port 4 nsew signal output
rlabel m2 s 23 11 26 14 6 Y
port 4 nsew signal output
rlabel m2 s 22 10 65 11 6 Y
port 4 nsew signal output
rlabel m2 s 22 11 23 14 6 Y
port 4 nsew signal output
rlabel m2 s 22 14 65 15 6 Y
port 4 nsew signal output
rlabel m2c s 68 25 71 28 6 Y
port 4 nsew signal output
rlabel m2c s 61 11 64 14 6 Y
port 4 nsew signal output
rlabel m2c s 56 25 59 28 6 Y
port 4 nsew signal output
rlabel m2c s 34 25 37 28 6 Y
port 4 nsew signal output
rlabel m2c s 23 11 26 14 6 Y
port 4 nsew signal output
rlabel m1 s 71 25 72 28 6 Y
port 4 nsew signal output
rlabel m1 s 68 25 71 28 6 Y
port 4 nsew signal output
rlabel m1 s 67 25 68 28 6 Y
port 4 nsew signal output
rlabel m1 s 61 11 64 14 6 Y
port 4 nsew signal output
rlabel m1 s 59 25 60 28 6 Y
port 4 nsew signal output
rlabel m1 s 56 11 61 14 6 Y
port 4 nsew signal output
rlabel m1 s 56 14 64 15 6 Y
port 4 nsew signal output
rlabel m1 s 56 15 60 25 6 Y
port 4 nsew signal output
rlabel m1 s 56 25 59 28 6 Y
port 4 nsew signal output
rlabel m1 s 56 28 60 29 6 Y
port 4 nsew signal output
rlabel m1 s 37 25 38 28 6 Y
port 4 nsew signal output
rlabel m1 s 34 25 37 28 6 Y
port 4 nsew signal output
rlabel m1 s 33 25 34 28 6 Y
port 4 nsew signal output
rlabel m1 s 56 4 60 10 6 Y
port 4 nsew signal output
rlabel m1 s 56 10 64 11 6 Y
port 4 nsew signal output
rlabel m1 s 26 11 27 14 6 Y
port 4 nsew signal output
rlabel m1 s 23 11 26 14 6 Y
port 4 nsew signal output
rlabel m1 s 22 11 23 14 6 Y
port 4 nsew signal output
rlabel m2 s 54 39 55 42 6 Vdd
port 5 nsew power input
rlabel m2 s 51 39 54 42 6 Vdd
port 5 nsew power input
rlabel m2 s 19 39 51 42 6 Vdd
port 5 nsew power input
rlabel m2 s 16 39 19 42 6 Vdd
port 5 nsew power input
rlabel m2 s 15 38 55 39 6 Vdd
port 5 nsew power input
rlabel m2 s 15 39 16 42 6 Vdd
port 5 nsew power input
rlabel m2 s 15 42 55 43 6 Vdd
port 5 nsew power input
rlabel m2c s 51 39 54 42 6 Vdd
port 5 nsew power input
rlabel m2c s 16 39 19 42 6 Vdd
port 5 nsew power input
rlabel m1 s 53 34 54 37 6 Vdd
port 5 nsew power input
rlabel m1 s 51 37 54 39 6 Vdd
port 5 nsew power input
rlabel m1 s 51 39 54 42 6 Vdd
port 5 nsew power input
rlabel m1 s 51 42 54 43 6 Vdd
port 5 nsew power input
rlabel m1 s 50 34 53 37 6 Vdd
port 5 nsew power input
rlabel m1 s 49 34 50 37 6 Vdd
port 5 nsew power input
rlabel m1 s 19 40 20 42 6 Vdd
port 5 nsew power input
rlabel m1 s 16 39 19 42 6 Vdd
port 5 nsew power input
rlabel m1 s 16 26 19 27 6 Vdd
port 5 nsew power input
rlabel m1 s 16 27 19 30 6 Vdd
port 5 nsew power input
rlabel m1 s 16 30 19 39 6 Vdd
port 5 nsew power input
rlabel m1 s 16 42 20 44 6 Vdd
port 5 nsew power input
rlabel m2 s 44 4 46 7 6 GND
port 6 nsew ground input
rlabel m2 s 41 4 44 7 6 GND
port 6 nsew ground input
rlabel m2 s 12 4 41 7 6 GND
port 6 nsew ground input
rlabel m2 s 9 4 12 7 6 GND
port 6 nsew ground input
rlabel m2 s 8 3 46 4 6 GND
port 6 nsew ground input
rlabel m2 s 8 4 9 7 6 GND
port 6 nsew ground input
rlabel m2 s 8 7 46 8 6 GND
port 6 nsew ground input
rlabel m2c s 41 4 44 7 6 GND
port 6 nsew ground input
rlabel m2c s 9 4 12 7 6 GND
port 6 nsew ground input
rlabel m1 s 41 14 44 15 6 GND
port 6 nsew ground input
rlabel m1 s 41 11 44 14 6 GND
port 6 nsew ground input
rlabel m1 s 41 3 44 4 6 GND
port 6 nsew ground input
rlabel m1 s 41 4 44 7 6 GND
port 6 nsew ground input
rlabel m1 s 41 7 44 11 6 GND
port 6 nsew ground input
rlabel m1 s 9 4 12 7 6 GND
port 6 nsew ground input
rlabel m1 s 9 8 12 11 6 GND
port 6 nsew ground input
rlabel m1 s 8 3 12 4 6 GND
port 6 nsew ground input
rlabel m1 s 8 4 9 7 6 GND
port 6 nsew ground input
rlabel m1 s 8 7 12 8 6 GND
port 6 nsew ground input
rlabel m1 s 8 8 9 11 6 GND
port 6 nsew ground input
rlabel m1 s 8 11 12 12 6 GND
port 6 nsew ground input
rlabel space 0 0 88 48 1 prboundary
rlabel ndiffusion 72 9 72 9 3 #10
rlabel polysilicon 76 18 76 18 3 _S
rlabel ndiffusion 68 7 68 7 3 #10
rlabel ndiffusion 68 9 68 9 3 #10
rlabel ndiffusion 68 12 68 12 3 #10
rlabel pdiffusion 68 24 68 24 3 Y
rlabel pdiffusion 68 29 68 29 3 Y
rlabel polysilicon 48 39 48 39 3 B
rlabel ntransistor 66 7 66 7 3 _S
rlabel polysilicon 66 17 66 17 3 _S
rlabel polysilicon 66 21 66 21 3 _S
rlabel polysilicon 66 22 66 22 3 _S
rlabel polysilicon 66 23 66 23 3 _S
rlabel ptransistor 66 24 66 24 3 _S
rlabel polysilicon 66 39 66 39 3 _S
rlabel pdiffusion 50 24 50 24 3 Vdd
rlabel pdiffusion 50 38 50 38 3 Vdd
rlabel polysilicon 44 42 44 42 3 B
rlabel polysilicon 44 43 44 43 3 B
rlabel polysilicon 44 46 44 46 3 B
rlabel ndiffusion 61 7 61 7 3 Y
rlabel ndiffusion 54 9 54 9 3 #10
rlabel ndiffusion 61 12 61 12 3 Y
rlabel ndiffusion 61 15 61 15 3 Y
rlabel pdiffusion 61 24 61 24 3 #5
rlabel pdiffusion 61 36 61 36 3 #5
rlabel ndiffusion 45 12 45 12 3 GND
rlabel ndiffusion 38 13 38 13 3 _S
rlabel polysilicon 48 17 48 17 3 B
rlabel ptransistor 48 24 48 24 3 B
rlabel polysilicon 39 39 39 39 3 S
rlabel ndiffusion 50 7 50 7 3 #10
rlabel ndiffusion 50 9 50 9 3 #10
rlabel ndiffusion 50 12 50 12 3 #10
rlabel ndiffusion 41 11 41 11 3 GND
rlabel ndiffusion 41 12 41 12 3 GND
rlabel ndiffusion 41 15 41 15 3 GND
rlabel ndiffusion 34 13 34 13 3 _S
rlabel polysilicon 39 17 39 17 3 S
rlabel ptransistor 39 24 39 24 3 S
rlabel polysilicon 66 5 66 5 3 _S
rlabel ntransistor 48 7 48 7 3 B
rlabel polysilicon 39 9 39 9 3 S
rlabel ntransistor 39 11 39 11 3 S
rlabel ndiffusion 34 16 34 16 3 _S
rlabel pdiffusion 34 24 34 24 3 Y
rlabel ndiffusion 44 7 44 7 3 GND
rlabel ndiffusion 34 11 34 11 3 _S
rlabel pdiffusion 27 25 27 25 3 _S
rlabel polysilicon 33 42 33 42 3 S
rlabel polysilicon 33 43 33 43 3 S
rlabel polysilicon 33 46 33 46 3 S
rlabel polysilicon 48 5 48 5 3 B
rlabel ndiffusion 23 7 23 7 3 Y
rlabel pdiffusion 23 24 23 24 3 _S
rlabel pdiffusion 23 25 23 25 3 _S
rlabel pdiffusion 23 28 23 28 3 _S
rlabel pdiffusion 20 28 20 28 3 Vdd
rlabel polysilicon 21 32 21 32 3 S
rlabel polysilicon 21 35 21 35 3 S
rlabel polysilicon 21 36 21 36 3 S
rlabel polysilicon 21 39 21 39 3 S
rlabel polysilicon 21 5 21 5 3 S
rlabel ntransistor 21 7 21 7 3 S
rlabel polysilicon 21 17 21 17 3 S
rlabel ptransistor 21 24 21 24 3 S
rlabel polysilicon 14 43 14 43 3 A
rlabel ndiffusion 13 9 13 9 3 GND
rlabel pdiffusion 16 24 16 24 3 Vdd
rlabel pdiffusion 16 28 16 28 3 Vdd
rlabel pdiffusion 16 31 16 31 3 Vdd
rlabel pdiffusion 16 32 16 32 3 Vdd
rlabel polysilicon 14 39 14 39 3 A
rlabel polysilicon 14 5 14 5 3 A
rlabel ntransistor 14 7 14 7 3 A
rlabel polysilicon 14 17 14 17 3 A
rlabel ptransistor 14 24 14 24 3 A
rlabel polysilicon 10 42 10 42 3 A
rlabel polysilicon 10 43 10 43 3 A
rlabel polysilicon 10 46 10 46 3 A
rlabel ndiffusion 9 7 9 7 3 GND
rlabel pdiffusion 9 24 9 24 3 #5
rlabel m1 76 19 76 19 3 _S
rlabel m1 69 12 69 12 3 #10
rlabel m1 68 26 68 26 3 Y
port 4 e default output
rlabel m1 61 33 61 33 3 #5
rlabel m1 57 12 57 12 3 Y
port 4 e default output
rlabel m1 57 15 57 15 3 Y
port 4 e default output
rlabel m1 57 16 57 16 3 Y
port 4 e default output
rlabel m1 57 29 57 29 3 Y
port 4 e default output
rlabel m1 54 35 54 35 3 Vdd
rlabel m1 52 38 52 38 3 Vdd
rlabel m1 52 43 52 43 3 Vdd
rlabel pdc 51 35 51 35 3 Vdd
rlabel m1 48 43 48 43 3 B
port 2 e default input
rlabel m1 51 12 51 12 3 #10
rlabel m1 50 35 50 35 3 Vdd
rlabel pc 45 43 45 43 3 B
port 2 e
rlabel m1 42 15 42 15 3 GND
rlabel m1 41 41 41 41 3 B
port 2 e
rlabel ndc 42 12 42 12 3 GND
rlabel m1 35 12 35 12 3 _S
rlabel ndc 35 13 35 13 3 _S
rlabel m1 35 16 35 16 3 _S
rlabel m1 35 22 35 22 3 _S
rlabel m1 69 8 69 8 3 #10
rlabel ndc 69 9 69 9 3 #10
rlabel m1 37 43 37 43 3 S
port 3 e default input
rlabel m1 69 4 69 4 3 #10
rlabel m1 28 36 28 36 3 S
port 3 e default input
rlabel pc 34 43 34 43 3 S
port 3 e default input
rlabel m1 57 5 57 5 3 Y
port 4 e default output
rlabel m1 57 11 57 11 3 Y
port 4 e default output
rlabel m1 25 35 25 35 3 S
port 3 e default input
rlabel pc 25 36 25 36 3 S
port 3 e default input
rlabel m1 25 39 25 39 3 S
port 3 e default input
rlabel m1 25 42 25 42 3 S
port 3 e default input
rlabel m1 25 43 25 43 3 S
port 3 e
rlabel m1 24 18 24 18 3 _S
rlabel m1 24 22 24 22 3 _S
rlabel pdc 24 25 24 25 3 _S
rlabel m1 24 28 24 28 3 _S
rlabel m1 20 41 20 41 3 Vdd
rlabel m1 51 4 51 4 3 #10
rlabel m1 51 8 51 8 3 #10
rlabel ndc 51 9 51 9 3 #10
rlabel m1 17 27 17 27 3 Vdd
rlabel pdc 17 28 17 28 3 Vdd
rlabel m1 17 31 17 31 3 Vdd
rlabel m1 17 43 17 43 3 Vdd
rlabel m1 42 4 42 4 3 GND
rlabel m1 42 8 42 8 3 GND
rlabel ndc 10 9 10 9 3 GND
rlabel pc 11 43 11 43 3 A
port 1 e default input
rlabel m1 9 9 9 9 3 GND
rlabel m1 9 12 9 12 3 GND
rlabel m1 9 41 9 41 3 A
port 1 e default input
rlabel m1 9 43 9 43 3 A
port 1 e
rlabel m1 9 46 9 46 3 A
port 1 e
rlabel m2 72 26 72 26 3 Y
port 4 e default output
rlabel m2c 69 26 69 26 3 Y
port 4 e default output
rlabel m2 60 26 60 26 3 Y
port 4 e default output
rlabel m2 72 5 72 5 3 #10
rlabel m2 80 19 80 19 3 _S
rlabel m2c 57 26 57 26 3 Y
port 4 e default output
rlabel m2c 69 5 69 5 3 #10
rlabel m2c 77 19 77 19 3 _S
rlabel m2 38 26 38 26 3 Y
port 4 e default output
rlabel m2 54 5 54 5 3 #10
rlabel m2 65 12 65 12 3 Y
port 4 e default output
rlabel m2 38 19 38 19 3 _S
rlabel m2c 35 26 35 26 3 Y
port 4 e default output
rlabel m2c 51 5 51 5 3 #10
rlabel m2c 62 12 62 12 3 Y
port 4 e default output
rlabel m2c 35 19 35 19 3 _S
rlabel m2 34 25 34 25 3 Y
port 4 e default output
rlabel m2 34 26 34 26 3 Y
port 4 e default output
rlabel m2 34 29 34 29 3 Y
port 4 e default output
rlabel m2 55 40 55 40 3 Vdd
rlabel m2 50 5 50 5 3 #10
rlabel m2 27 12 27 12 3 Y
port 4 e
rlabel m2 27 19 27 19 3 _S
rlabel m2c 52 40 52 40 3 Vdd
rlabel m2c 24 12 24 12 3 Y
port 4 e
rlabel m2c 24 19 24 19 3 _S
rlabel m2 20 40 20 40 3 Vdd
rlabel m2 45 5 45 5 3 GND
rlabel m2 23 11 23 11 3 Y
port 4 e
rlabel m2 23 12 23 12 3 Y
port 4 e
rlabel m2 23 15 23 15 3 Y
port 4 e
rlabel m2 23 18 23 18 3 _S
rlabel m2 23 19 23 19 3 _S
rlabel m2 23 22 23 22 3 _S
rlabel m2 65 33 65 33 3 #5
rlabel m2c 17 40 17 40 3 Vdd
rlabel m2c 42 5 42 5 3 GND
rlabel m2c 62 33 62 33 3 #5
rlabel m2 16 39 16 39 3 Vdd
rlabel m2 16 40 16 40 3 Vdd
rlabel m2 16 43 16 43 3 Vdd
rlabel m2 50 4 50 4 3 #10
rlabel m2 13 5 13 5 3 GND
rlabel m2 50 8 50 8 3 #10
rlabel m2 13 33 13 33 3 #5
rlabel m2c 10 5 10 5 3 GND
rlabel m2c 10 33 10 33 3 #5
rlabel m2 9 4 9 4 3 GND
rlabel m2 9 5 9 5 3 GND
rlabel m2 9 8 9 8 3 GND
rlabel m2 9 32 9 32 3 #5
rlabel m2 9 33 9 33 3 #5
rlabel m2 9 36 9 36 3 #5
<< properties >>
string LEFsite CoreSite
string LEFclass CORE
string FIXED_BBOX 0 0 88 48
string LEFsymmetry X Y
string LEFview TRUE
<< end >>
