magic
tech sky130l
timestamp 1731220556
<< m2 >>
rect 142 3642 148 3643
rect 142 3638 143 3642
rect 147 3638 148 3642
rect 142 3637 148 3638
rect 222 3642 228 3643
rect 222 3638 223 3642
rect 227 3638 228 3642
rect 222 3637 228 3638
rect 350 3642 356 3643
rect 350 3638 351 3642
rect 355 3638 356 3642
rect 350 3637 356 3638
rect 494 3642 500 3643
rect 494 3638 495 3642
rect 499 3638 500 3642
rect 494 3637 500 3638
rect 646 3642 652 3643
rect 646 3638 647 3642
rect 651 3638 652 3642
rect 646 3637 652 3638
rect 806 3642 812 3643
rect 806 3638 807 3642
rect 811 3638 812 3642
rect 806 3637 812 3638
rect 974 3642 980 3643
rect 974 3638 975 3642
rect 979 3638 980 3642
rect 974 3637 980 3638
rect 1150 3642 1156 3643
rect 1150 3638 1151 3642
rect 1155 3638 1156 3642
rect 1150 3637 1156 3638
rect 1334 3642 1340 3643
rect 1334 3638 1335 3642
rect 1339 3638 1340 3642
rect 1334 3637 1340 3638
rect 110 3624 116 3625
rect 110 3620 111 3624
rect 115 3620 116 3624
rect 110 3619 116 3620
rect 1830 3624 1836 3625
rect 1830 3620 1831 3624
rect 1835 3620 1836 3624
rect 1830 3619 1836 3620
rect 1926 3614 1932 3615
rect 1926 3610 1927 3614
rect 1931 3610 1932 3614
rect 1926 3609 1932 3610
rect 2006 3614 2012 3615
rect 2006 3610 2007 3614
rect 2011 3610 2012 3614
rect 2006 3609 2012 3610
rect 2102 3614 2108 3615
rect 2102 3610 2103 3614
rect 2107 3610 2108 3614
rect 2102 3609 2108 3610
rect 2206 3614 2212 3615
rect 2206 3610 2207 3614
rect 2211 3610 2212 3614
rect 2206 3609 2212 3610
rect 2318 3614 2324 3615
rect 2318 3610 2319 3614
rect 2323 3610 2324 3614
rect 2318 3609 2324 3610
rect 2430 3614 2436 3615
rect 2430 3610 2431 3614
rect 2435 3610 2436 3614
rect 2430 3609 2436 3610
rect 2550 3614 2556 3615
rect 2550 3610 2551 3614
rect 2555 3610 2556 3614
rect 2550 3609 2556 3610
rect 2662 3614 2668 3615
rect 2662 3610 2663 3614
rect 2667 3610 2668 3614
rect 2662 3609 2668 3610
rect 2774 3614 2780 3615
rect 2774 3610 2775 3614
rect 2779 3610 2780 3614
rect 2774 3609 2780 3610
rect 2878 3614 2884 3615
rect 2878 3610 2879 3614
rect 2883 3610 2884 3614
rect 2878 3609 2884 3610
rect 2982 3614 2988 3615
rect 2982 3610 2983 3614
rect 2987 3610 2988 3614
rect 2982 3609 2988 3610
rect 3094 3614 3100 3615
rect 3094 3610 3095 3614
rect 3099 3610 3100 3614
rect 3094 3609 3100 3610
rect 3206 3614 3212 3615
rect 3206 3610 3207 3614
rect 3211 3610 3212 3614
rect 3206 3609 3212 3610
rect 110 3607 116 3608
rect 110 3603 111 3607
rect 115 3603 116 3607
rect 1830 3607 1836 3608
rect 110 3602 116 3603
rect 134 3604 140 3605
rect 134 3600 135 3604
rect 139 3600 140 3604
rect 134 3599 140 3600
rect 214 3604 220 3605
rect 214 3600 215 3604
rect 219 3600 220 3604
rect 214 3599 220 3600
rect 342 3604 348 3605
rect 342 3600 343 3604
rect 347 3600 348 3604
rect 342 3599 348 3600
rect 486 3604 492 3605
rect 486 3600 487 3604
rect 491 3600 492 3604
rect 486 3599 492 3600
rect 638 3604 644 3605
rect 638 3600 639 3604
rect 643 3600 644 3604
rect 638 3599 644 3600
rect 798 3604 804 3605
rect 798 3600 799 3604
rect 803 3600 804 3604
rect 798 3599 804 3600
rect 966 3604 972 3605
rect 966 3600 967 3604
rect 971 3600 972 3604
rect 966 3599 972 3600
rect 1142 3604 1148 3605
rect 1142 3600 1143 3604
rect 1147 3600 1148 3604
rect 1142 3599 1148 3600
rect 1326 3604 1332 3605
rect 1326 3600 1327 3604
rect 1331 3600 1332 3604
rect 1830 3603 1831 3607
rect 1835 3603 1836 3607
rect 1830 3602 1836 3603
rect 1326 3599 1332 3600
rect 1870 3596 1876 3597
rect 1870 3592 1871 3596
rect 1875 3592 1876 3596
rect 1870 3591 1876 3592
rect 3590 3596 3596 3597
rect 3590 3592 3591 3596
rect 3595 3592 3596 3596
rect 3590 3591 3596 3592
rect 1870 3579 1876 3580
rect 1870 3575 1871 3579
rect 1875 3575 1876 3579
rect 3590 3579 3596 3580
rect 1870 3574 1876 3575
rect 1918 3576 1924 3577
rect 1918 3572 1919 3576
rect 1923 3572 1924 3576
rect 1918 3571 1924 3572
rect 1998 3576 2004 3577
rect 1998 3572 1999 3576
rect 2003 3572 2004 3576
rect 1998 3571 2004 3572
rect 2094 3576 2100 3577
rect 2094 3572 2095 3576
rect 2099 3572 2100 3576
rect 2094 3571 2100 3572
rect 2198 3576 2204 3577
rect 2198 3572 2199 3576
rect 2203 3572 2204 3576
rect 2198 3571 2204 3572
rect 2310 3576 2316 3577
rect 2310 3572 2311 3576
rect 2315 3572 2316 3576
rect 2310 3571 2316 3572
rect 2422 3576 2428 3577
rect 2422 3572 2423 3576
rect 2427 3572 2428 3576
rect 2422 3571 2428 3572
rect 2542 3576 2548 3577
rect 2542 3572 2543 3576
rect 2547 3572 2548 3576
rect 2542 3571 2548 3572
rect 2654 3576 2660 3577
rect 2654 3572 2655 3576
rect 2659 3572 2660 3576
rect 2654 3571 2660 3572
rect 2766 3576 2772 3577
rect 2766 3572 2767 3576
rect 2771 3572 2772 3576
rect 2766 3571 2772 3572
rect 2870 3576 2876 3577
rect 2870 3572 2871 3576
rect 2875 3572 2876 3576
rect 2870 3571 2876 3572
rect 2974 3576 2980 3577
rect 2974 3572 2975 3576
rect 2979 3572 2980 3576
rect 2974 3571 2980 3572
rect 3086 3576 3092 3577
rect 3086 3572 3087 3576
rect 3091 3572 3092 3576
rect 3086 3571 3092 3572
rect 3198 3576 3204 3577
rect 3198 3572 3199 3576
rect 3203 3572 3204 3576
rect 3590 3575 3591 3579
rect 3595 3575 3596 3579
rect 3590 3574 3596 3575
rect 3198 3571 3204 3572
rect 238 3560 244 3561
rect 110 3557 116 3558
rect 110 3553 111 3557
rect 115 3553 116 3557
rect 238 3556 239 3560
rect 243 3556 244 3560
rect 238 3555 244 3556
rect 358 3560 364 3561
rect 358 3556 359 3560
rect 363 3556 364 3560
rect 358 3555 364 3556
rect 478 3560 484 3561
rect 478 3556 479 3560
rect 483 3556 484 3560
rect 478 3555 484 3556
rect 606 3560 612 3561
rect 606 3556 607 3560
rect 611 3556 612 3560
rect 606 3555 612 3556
rect 734 3560 740 3561
rect 734 3556 735 3560
rect 739 3556 740 3560
rect 734 3555 740 3556
rect 862 3560 868 3561
rect 862 3556 863 3560
rect 867 3556 868 3560
rect 862 3555 868 3556
rect 982 3560 988 3561
rect 982 3556 983 3560
rect 987 3556 988 3560
rect 982 3555 988 3556
rect 1094 3560 1100 3561
rect 1094 3556 1095 3560
rect 1099 3556 1100 3560
rect 1094 3555 1100 3556
rect 1206 3560 1212 3561
rect 1206 3556 1207 3560
rect 1211 3556 1212 3560
rect 1206 3555 1212 3556
rect 1318 3560 1324 3561
rect 1318 3556 1319 3560
rect 1323 3556 1324 3560
rect 1318 3555 1324 3556
rect 1438 3560 1444 3561
rect 1438 3556 1439 3560
rect 1443 3556 1444 3560
rect 1438 3555 1444 3556
rect 1830 3557 1836 3558
rect 110 3552 116 3553
rect 1830 3553 1831 3557
rect 1835 3553 1836 3557
rect 1830 3552 1836 3553
rect 110 3540 116 3541
rect 110 3536 111 3540
rect 115 3536 116 3540
rect 110 3535 116 3536
rect 1830 3540 1836 3541
rect 1830 3536 1831 3540
rect 1835 3536 1836 3540
rect 1830 3535 1836 3536
rect 1942 3532 1948 3533
rect 1870 3529 1876 3530
rect 1870 3525 1871 3529
rect 1875 3525 1876 3529
rect 1942 3528 1943 3532
rect 1947 3528 1948 3532
rect 1942 3527 1948 3528
rect 2126 3532 2132 3533
rect 2126 3528 2127 3532
rect 2131 3528 2132 3532
rect 2126 3527 2132 3528
rect 2302 3532 2308 3533
rect 2302 3528 2303 3532
rect 2307 3528 2308 3532
rect 2302 3527 2308 3528
rect 2478 3532 2484 3533
rect 2478 3528 2479 3532
rect 2483 3528 2484 3532
rect 2478 3527 2484 3528
rect 2646 3532 2652 3533
rect 2646 3528 2647 3532
rect 2651 3528 2652 3532
rect 2646 3527 2652 3528
rect 2814 3532 2820 3533
rect 2814 3528 2815 3532
rect 2819 3528 2820 3532
rect 2814 3527 2820 3528
rect 2974 3532 2980 3533
rect 2974 3528 2975 3532
rect 2979 3528 2980 3532
rect 2974 3527 2980 3528
rect 3134 3532 3140 3533
rect 3134 3528 3135 3532
rect 3139 3528 3140 3532
rect 3134 3527 3140 3528
rect 3302 3532 3308 3533
rect 3302 3528 3303 3532
rect 3307 3528 3308 3532
rect 3302 3527 3308 3528
rect 3590 3529 3596 3530
rect 1870 3524 1876 3525
rect 3590 3525 3591 3529
rect 3595 3525 3596 3529
rect 3590 3524 3596 3525
rect 246 3522 252 3523
rect 246 3518 247 3522
rect 251 3518 252 3522
rect 246 3517 252 3518
rect 366 3522 372 3523
rect 366 3518 367 3522
rect 371 3518 372 3522
rect 366 3517 372 3518
rect 486 3522 492 3523
rect 486 3518 487 3522
rect 491 3518 492 3522
rect 486 3517 492 3518
rect 614 3522 620 3523
rect 614 3518 615 3522
rect 619 3518 620 3522
rect 614 3517 620 3518
rect 742 3522 748 3523
rect 742 3518 743 3522
rect 747 3518 748 3522
rect 742 3517 748 3518
rect 870 3522 876 3523
rect 870 3518 871 3522
rect 875 3518 876 3522
rect 870 3517 876 3518
rect 990 3522 996 3523
rect 990 3518 991 3522
rect 995 3518 996 3522
rect 990 3517 996 3518
rect 1102 3522 1108 3523
rect 1102 3518 1103 3522
rect 1107 3518 1108 3522
rect 1102 3517 1108 3518
rect 1214 3522 1220 3523
rect 1214 3518 1215 3522
rect 1219 3518 1220 3522
rect 1214 3517 1220 3518
rect 1326 3522 1332 3523
rect 1326 3518 1327 3522
rect 1331 3518 1332 3522
rect 1326 3517 1332 3518
rect 1446 3522 1452 3523
rect 1446 3518 1447 3522
rect 1451 3518 1452 3522
rect 1446 3517 1452 3518
rect 1870 3512 1876 3513
rect 1870 3508 1871 3512
rect 1875 3508 1876 3512
rect 1870 3507 1876 3508
rect 3590 3512 3596 3513
rect 3590 3508 3591 3512
rect 3595 3508 3596 3512
rect 3590 3507 3596 3508
rect 1950 3494 1956 3495
rect 166 3490 172 3491
rect 166 3486 167 3490
rect 171 3486 172 3490
rect 166 3485 172 3486
rect 286 3490 292 3491
rect 286 3486 287 3490
rect 291 3486 292 3490
rect 286 3485 292 3486
rect 414 3490 420 3491
rect 414 3486 415 3490
rect 419 3486 420 3490
rect 414 3485 420 3486
rect 550 3490 556 3491
rect 550 3486 551 3490
rect 555 3486 556 3490
rect 550 3485 556 3486
rect 686 3490 692 3491
rect 686 3486 687 3490
rect 691 3486 692 3490
rect 686 3485 692 3486
rect 822 3490 828 3491
rect 822 3486 823 3490
rect 827 3486 828 3490
rect 822 3485 828 3486
rect 950 3490 956 3491
rect 950 3486 951 3490
rect 955 3486 956 3490
rect 950 3485 956 3486
rect 1070 3490 1076 3491
rect 1070 3486 1071 3490
rect 1075 3486 1076 3490
rect 1070 3485 1076 3486
rect 1182 3490 1188 3491
rect 1182 3486 1183 3490
rect 1187 3486 1188 3490
rect 1182 3485 1188 3486
rect 1302 3490 1308 3491
rect 1302 3486 1303 3490
rect 1307 3486 1308 3490
rect 1302 3485 1308 3486
rect 1422 3490 1428 3491
rect 1422 3486 1423 3490
rect 1427 3486 1428 3490
rect 1950 3490 1951 3494
rect 1955 3490 1956 3494
rect 1950 3489 1956 3490
rect 2134 3494 2140 3495
rect 2134 3490 2135 3494
rect 2139 3490 2140 3494
rect 2134 3489 2140 3490
rect 2310 3494 2316 3495
rect 2310 3490 2311 3494
rect 2315 3490 2316 3494
rect 2310 3489 2316 3490
rect 2486 3494 2492 3495
rect 2486 3490 2487 3494
rect 2491 3490 2492 3494
rect 2486 3489 2492 3490
rect 2654 3494 2660 3495
rect 2654 3490 2655 3494
rect 2659 3490 2660 3494
rect 2654 3489 2660 3490
rect 2822 3494 2828 3495
rect 2822 3490 2823 3494
rect 2827 3490 2828 3494
rect 2822 3489 2828 3490
rect 2982 3494 2988 3495
rect 2982 3490 2983 3494
rect 2987 3490 2988 3494
rect 2982 3489 2988 3490
rect 3142 3494 3148 3495
rect 3142 3490 3143 3494
rect 3147 3490 3148 3494
rect 3142 3489 3148 3490
rect 3310 3494 3316 3495
rect 3310 3490 3311 3494
rect 3315 3490 3316 3494
rect 3310 3489 3316 3490
rect 1422 3485 1428 3486
rect 110 3472 116 3473
rect 110 3468 111 3472
rect 115 3468 116 3472
rect 110 3467 116 3468
rect 1830 3472 1836 3473
rect 1830 3468 1831 3472
rect 1835 3468 1836 3472
rect 1830 3467 1836 3468
rect 1958 3462 1964 3463
rect 1958 3458 1959 3462
rect 1963 3458 1964 3462
rect 1958 3457 1964 3458
rect 2078 3462 2084 3463
rect 2078 3458 2079 3462
rect 2083 3458 2084 3462
rect 2078 3457 2084 3458
rect 2198 3462 2204 3463
rect 2198 3458 2199 3462
rect 2203 3458 2204 3462
rect 2198 3457 2204 3458
rect 2334 3462 2340 3463
rect 2334 3458 2335 3462
rect 2339 3458 2340 3462
rect 2334 3457 2340 3458
rect 2478 3462 2484 3463
rect 2478 3458 2479 3462
rect 2483 3458 2484 3462
rect 2478 3457 2484 3458
rect 2630 3462 2636 3463
rect 2630 3458 2631 3462
rect 2635 3458 2636 3462
rect 2630 3457 2636 3458
rect 2790 3462 2796 3463
rect 2790 3458 2791 3462
rect 2795 3458 2796 3462
rect 2790 3457 2796 3458
rect 2958 3462 2964 3463
rect 2958 3458 2959 3462
rect 2963 3458 2964 3462
rect 2958 3457 2964 3458
rect 3126 3462 3132 3463
rect 3126 3458 3127 3462
rect 3131 3458 3132 3462
rect 3126 3457 3132 3458
rect 3302 3462 3308 3463
rect 3302 3458 3303 3462
rect 3307 3458 3308 3462
rect 3302 3457 3308 3458
rect 110 3455 116 3456
rect 110 3451 111 3455
rect 115 3451 116 3455
rect 1830 3455 1836 3456
rect 110 3450 116 3451
rect 158 3452 164 3453
rect 158 3448 159 3452
rect 163 3448 164 3452
rect 158 3447 164 3448
rect 278 3452 284 3453
rect 278 3448 279 3452
rect 283 3448 284 3452
rect 278 3447 284 3448
rect 406 3452 412 3453
rect 406 3448 407 3452
rect 411 3448 412 3452
rect 406 3447 412 3448
rect 542 3452 548 3453
rect 542 3448 543 3452
rect 547 3448 548 3452
rect 542 3447 548 3448
rect 678 3452 684 3453
rect 678 3448 679 3452
rect 683 3448 684 3452
rect 678 3447 684 3448
rect 814 3452 820 3453
rect 814 3448 815 3452
rect 819 3448 820 3452
rect 814 3447 820 3448
rect 942 3452 948 3453
rect 942 3448 943 3452
rect 947 3448 948 3452
rect 942 3447 948 3448
rect 1062 3452 1068 3453
rect 1062 3448 1063 3452
rect 1067 3448 1068 3452
rect 1062 3447 1068 3448
rect 1174 3452 1180 3453
rect 1174 3448 1175 3452
rect 1179 3448 1180 3452
rect 1174 3447 1180 3448
rect 1294 3452 1300 3453
rect 1294 3448 1295 3452
rect 1299 3448 1300 3452
rect 1294 3447 1300 3448
rect 1414 3452 1420 3453
rect 1414 3448 1415 3452
rect 1419 3448 1420 3452
rect 1830 3451 1831 3455
rect 1835 3451 1836 3455
rect 1830 3450 1836 3451
rect 1414 3447 1420 3448
rect 1870 3444 1876 3445
rect 1870 3440 1871 3444
rect 1875 3440 1876 3444
rect 1870 3439 1876 3440
rect 3590 3444 3596 3445
rect 3590 3440 3591 3444
rect 3595 3440 3596 3444
rect 3590 3439 3596 3440
rect 1870 3427 1876 3428
rect 1870 3423 1871 3427
rect 1875 3423 1876 3427
rect 3590 3427 3596 3428
rect 1870 3422 1876 3423
rect 1950 3424 1956 3425
rect 1950 3420 1951 3424
rect 1955 3420 1956 3424
rect 1950 3419 1956 3420
rect 2070 3424 2076 3425
rect 2070 3420 2071 3424
rect 2075 3420 2076 3424
rect 2070 3419 2076 3420
rect 2190 3424 2196 3425
rect 2190 3420 2191 3424
rect 2195 3420 2196 3424
rect 2190 3419 2196 3420
rect 2326 3424 2332 3425
rect 2326 3420 2327 3424
rect 2331 3420 2332 3424
rect 2326 3419 2332 3420
rect 2470 3424 2476 3425
rect 2470 3420 2471 3424
rect 2475 3420 2476 3424
rect 2470 3419 2476 3420
rect 2622 3424 2628 3425
rect 2622 3420 2623 3424
rect 2627 3420 2628 3424
rect 2622 3419 2628 3420
rect 2782 3424 2788 3425
rect 2782 3420 2783 3424
rect 2787 3420 2788 3424
rect 2782 3419 2788 3420
rect 2950 3424 2956 3425
rect 2950 3420 2951 3424
rect 2955 3420 2956 3424
rect 2950 3419 2956 3420
rect 3118 3424 3124 3425
rect 3118 3420 3119 3424
rect 3123 3420 3124 3424
rect 3118 3419 3124 3420
rect 3294 3424 3300 3425
rect 3294 3420 3295 3424
rect 3299 3420 3300 3424
rect 3590 3423 3591 3427
rect 3595 3423 3596 3427
rect 3590 3422 3596 3423
rect 3294 3419 3300 3420
rect 134 3400 140 3401
rect 110 3397 116 3398
rect 110 3393 111 3397
rect 115 3393 116 3397
rect 134 3396 135 3400
rect 139 3396 140 3400
rect 134 3395 140 3396
rect 246 3400 252 3401
rect 246 3396 247 3400
rect 251 3396 252 3400
rect 246 3395 252 3396
rect 374 3400 380 3401
rect 374 3396 375 3400
rect 379 3396 380 3400
rect 374 3395 380 3396
rect 502 3400 508 3401
rect 502 3396 503 3400
rect 507 3396 508 3400
rect 502 3395 508 3396
rect 638 3400 644 3401
rect 638 3396 639 3400
rect 643 3396 644 3400
rect 638 3395 644 3396
rect 774 3400 780 3401
rect 774 3396 775 3400
rect 779 3396 780 3400
rect 774 3395 780 3396
rect 902 3400 908 3401
rect 902 3396 903 3400
rect 907 3396 908 3400
rect 902 3395 908 3396
rect 1030 3400 1036 3401
rect 1030 3396 1031 3400
rect 1035 3396 1036 3400
rect 1030 3395 1036 3396
rect 1158 3400 1164 3401
rect 1158 3396 1159 3400
rect 1163 3396 1164 3400
rect 1158 3395 1164 3396
rect 1286 3400 1292 3401
rect 1286 3396 1287 3400
rect 1291 3396 1292 3400
rect 1286 3395 1292 3396
rect 1414 3400 1420 3401
rect 1414 3396 1415 3400
rect 1419 3396 1420 3400
rect 1414 3395 1420 3396
rect 1830 3397 1836 3398
rect 110 3392 116 3393
rect 1830 3393 1831 3397
rect 1835 3393 1836 3397
rect 1830 3392 1836 3393
rect 110 3380 116 3381
rect 110 3376 111 3380
rect 115 3376 116 3380
rect 110 3375 116 3376
rect 1830 3380 1836 3381
rect 1830 3376 1831 3380
rect 1835 3376 1836 3380
rect 1830 3375 1836 3376
rect 1974 3372 1980 3373
rect 1870 3369 1876 3370
rect 1870 3365 1871 3369
rect 1875 3365 1876 3369
rect 1974 3368 1975 3372
rect 1979 3368 1980 3372
rect 1974 3367 1980 3368
rect 2134 3372 2140 3373
rect 2134 3368 2135 3372
rect 2139 3368 2140 3372
rect 2134 3367 2140 3368
rect 2286 3372 2292 3373
rect 2286 3368 2287 3372
rect 2291 3368 2292 3372
rect 2286 3367 2292 3368
rect 2430 3372 2436 3373
rect 2430 3368 2431 3372
rect 2435 3368 2436 3372
rect 2430 3367 2436 3368
rect 2558 3372 2564 3373
rect 2558 3368 2559 3372
rect 2563 3368 2564 3372
rect 2558 3367 2564 3368
rect 2678 3372 2684 3373
rect 2678 3368 2679 3372
rect 2683 3368 2684 3372
rect 2678 3367 2684 3368
rect 2790 3372 2796 3373
rect 2790 3368 2791 3372
rect 2795 3368 2796 3372
rect 2790 3367 2796 3368
rect 2894 3372 2900 3373
rect 2894 3368 2895 3372
rect 2899 3368 2900 3372
rect 2894 3367 2900 3368
rect 2990 3372 2996 3373
rect 2990 3368 2991 3372
rect 2995 3368 2996 3372
rect 2990 3367 2996 3368
rect 3078 3372 3084 3373
rect 3078 3368 3079 3372
rect 3083 3368 3084 3372
rect 3078 3367 3084 3368
rect 3166 3372 3172 3373
rect 3166 3368 3167 3372
rect 3171 3368 3172 3372
rect 3166 3367 3172 3368
rect 3254 3372 3260 3373
rect 3254 3368 3255 3372
rect 3259 3368 3260 3372
rect 3254 3367 3260 3368
rect 3342 3372 3348 3373
rect 3342 3368 3343 3372
rect 3347 3368 3348 3372
rect 3342 3367 3348 3368
rect 3422 3372 3428 3373
rect 3422 3368 3423 3372
rect 3427 3368 3428 3372
rect 3422 3367 3428 3368
rect 3502 3372 3508 3373
rect 3502 3368 3503 3372
rect 3507 3368 3508 3372
rect 3502 3367 3508 3368
rect 3590 3369 3596 3370
rect 1870 3364 1876 3365
rect 3590 3365 3591 3369
rect 3595 3365 3596 3369
rect 3590 3364 3596 3365
rect 142 3362 148 3363
rect 142 3358 143 3362
rect 147 3358 148 3362
rect 142 3357 148 3358
rect 254 3362 260 3363
rect 254 3358 255 3362
rect 259 3358 260 3362
rect 254 3357 260 3358
rect 382 3362 388 3363
rect 382 3358 383 3362
rect 387 3358 388 3362
rect 382 3357 388 3358
rect 510 3362 516 3363
rect 510 3358 511 3362
rect 515 3358 516 3362
rect 510 3357 516 3358
rect 646 3362 652 3363
rect 646 3358 647 3362
rect 651 3358 652 3362
rect 646 3357 652 3358
rect 782 3362 788 3363
rect 782 3358 783 3362
rect 787 3358 788 3362
rect 782 3357 788 3358
rect 910 3362 916 3363
rect 910 3358 911 3362
rect 915 3358 916 3362
rect 910 3357 916 3358
rect 1038 3362 1044 3363
rect 1038 3358 1039 3362
rect 1043 3358 1044 3362
rect 1038 3357 1044 3358
rect 1166 3362 1172 3363
rect 1166 3358 1167 3362
rect 1171 3358 1172 3362
rect 1166 3357 1172 3358
rect 1294 3362 1300 3363
rect 1294 3358 1295 3362
rect 1299 3358 1300 3362
rect 1294 3357 1300 3358
rect 1422 3362 1428 3363
rect 1422 3358 1423 3362
rect 1427 3358 1428 3362
rect 1422 3357 1428 3358
rect 1870 3352 1876 3353
rect 1870 3348 1871 3352
rect 1875 3348 1876 3352
rect 1870 3347 1876 3348
rect 3590 3352 3596 3353
rect 3590 3348 3591 3352
rect 3595 3348 3596 3352
rect 3590 3347 3596 3348
rect 1982 3334 1988 3335
rect 1982 3330 1983 3334
rect 1987 3330 1988 3334
rect 1982 3329 1988 3330
rect 2142 3334 2148 3335
rect 2142 3330 2143 3334
rect 2147 3330 2148 3334
rect 2142 3329 2148 3330
rect 2294 3334 2300 3335
rect 2294 3330 2295 3334
rect 2299 3330 2300 3334
rect 2294 3329 2300 3330
rect 2438 3334 2444 3335
rect 2438 3330 2439 3334
rect 2443 3330 2444 3334
rect 2438 3329 2444 3330
rect 2566 3334 2572 3335
rect 2566 3330 2567 3334
rect 2571 3330 2572 3334
rect 2566 3329 2572 3330
rect 2686 3334 2692 3335
rect 2686 3330 2687 3334
rect 2691 3330 2692 3334
rect 2686 3329 2692 3330
rect 2798 3334 2804 3335
rect 2798 3330 2799 3334
rect 2803 3330 2804 3334
rect 2798 3329 2804 3330
rect 2902 3334 2908 3335
rect 2902 3330 2903 3334
rect 2907 3330 2908 3334
rect 2902 3329 2908 3330
rect 2998 3334 3004 3335
rect 2998 3330 2999 3334
rect 3003 3330 3004 3334
rect 2998 3329 3004 3330
rect 3086 3334 3092 3335
rect 3086 3330 3087 3334
rect 3091 3330 3092 3334
rect 3086 3329 3092 3330
rect 3174 3334 3180 3335
rect 3174 3330 3175 3334
rect 3179 3330 3180 3334
rect 3174 3329 3180 3330
rect 3262 3334 3268 3335
rect 3262 3330 3263 3334
rect 3267 3330 3268 3334
rect 3262 3329 3268 3330
rect 3350 3334 3356 3335
rect 3350 3330 3351 3334
rect 3355 3330 3356 3334
rect 3350 3329 3356 3330
rect 3430 3334 3436 3335
rect 3430 3330 3431 3334
rect 3435 3330 3436 3334
rect 3430 3329 3436 3330
rect 3510 3334 3516 3335
rect 3510 3330 3511 3334
rect 3515 3330 3516 3334
rect 3510 3329 3516 3330
rect 270 3326 276 3327
rect 270 3322 271 3326
rect 275 3322 276 3326
rect 270 3321 276 3322
rect 390 3326 396 3327
rect 390 3322 391 3326
rect 395 3322 396 3326
rect 390 3321 396 3322
rect 518 3326 524 3327
rect 518 3322 519 3326
rect 523 3322 524 3326
rect 518 3321 524 3322
rect 654 3326 660 3327
rect 654 3322 655 3326
rect 659 3322 660 3326
rect 654 3321 660 3322
rect 790 3326 796 3327
rect 790 3322 791 3326
rect 795 3322 796 3326
rect 790 3321 796 3322
rect 918 3326 924 3327
rect 918 3322 919 3326
rect 923 3322 924 3326
rect 918 3321 924 3322
rect 1054 3326 1060 3327
rect 1054 3322 1055 3326
rect 1059 3322 1060 3326
rect 1054 3321 1060 3322
rect 1190 3326 1196 3327
rect 1190 3322 1191 3326
rect 1195 3322 1196 3326
rect 1190 3321 1196 3322
rect 1326 3326 1332 3327
rect 1326 3322 1327 3326
rect 1331 3322 1332 3326
rect 1326 3321 1332 3322
rect 1462 3326 1468 3327
rect 1462 3322 1463 3326
rect 1467 3322 1468 3326
rect 1462 3321 1468 3322
rect 110 3308 116 3309
rect 110 3304 111 3308
rect 115 3304 116 3308
rect 110 3303 116 3304
rect 1830 3308 1836 3309
rect 1830 3304 1831 3308
rect 1835 3304 1836 3308
rect 1830 3303 1836 3304
rect 1934 3298 1940 3299
rect 1934 3294 1935 3298
rect 1939 3294 1940 3298
rect 1934 3293 1940 3294
rect 2070 3298 2076 3299
rect 2070 3294 2071 3298
rect 2075 3294 2076 3298
rect 2070 3293 2076 3294
rect 2206 3298 2212 3299
rect 2206 3294 2207 3298
rect 2211 3294 2212 3298
rect 2206 3293 2212 3294
rect 2366 3298 2372 3299
rect 2366 3294 2367 3298
rect 2371 3294 2372 3298
rect 2366 3293 2372 3294
rect 2550 3298 2556 3299
rect 2550 3294 2551 3298
rect 2555 3294 2556 3298
rect 2550 3293 2556 3294
rect 2766 3298 2772 3299
rect 2766 3294 2767 3298
rect 2771 3294 2772 3298
rect 2766 3293 2772 3294
rect 3006 3298 3012 3299
rect 3006 3294 3007 3298
rect 3011 3294 3012 3298
rect 3006 3293 3012 3294
rect 3254 3298 3260 3299
rect 3254 3294 3255 3298
rect 3259 3294 3260 3298
rect 3254 3293 3260 3294
rect 3510 3298 3516 3299
rect 3510 3294 3511 3298
rect 3515 3294 3516 3298
rect 3510 3293 3516 3294
rect 110 3291 116 3292
rect 110 3287 111 3291
rect 115 3287 116 3291
rect 1830 3291 1836 3292
rect 110 3286 116 3287
rect 262 3288 268 3289
rect 262 3284 263 3288
rect 267 3284 268 3288
rect 262 3283 268 3284
rect 382 3288 388 3289
rect 382 3284 383 3288
rect 387 3284 388 3288
rect 382 3283 388 3284
rect 510 3288 516 3289
rect 510 3284 511 3288
rect 515 3284 516 3288
rect 510 3283 516 3284
rect 646 3288 652 3289
rect 646 3284 647 3288
rect 651 3284 652 3288
rect 646 3283 652 3284
rect 782 3288 788 3289
rect 782 3284 783 3288
rect 787 3284 788 3288
rect 782 3283 788 3284
rect 910 3288 916 3289
rect 910 3284 911 3288
rect 915 3284 916 3288
rect 910 3283 916 3284
rect 1046 3288 1052 3289
rect 1046 3284 1047 3288
rect 1051 3284 1052 3288
rect 1046 3283 1052 3284
rect 1182 3288 1188 3289
rect 1182 3284 1183 3288
rect 1187 3284 1188 3288
rect 1182 3283 1188 3284
rect 1318 3288 1324 3289
rect 1318 3284 1319 3288
rect 1323 3284 1324 3288
rect 1318 3283 1324 3284
rect 1454 3288 1460 3289
rect 1454 3284 1455 3288
rect 1459 3284 1460 3288
rect 1830 3287 1831 3291
rect 1835 3287 1836 3291
rect 1830 3286 1836 3287
rect 1454 3283 1460 3284
rect 1870 3280 1876 3281
rect 1870 3276 1871 3280
rect 1875 3276 1876 3280
rect 1870 3275 1876 3276
rect 3590 3280 3596 3281
rect 3590 3276 3591 3280
rect 3595 3276 3596 3280
rect 3590 3275 3596 3276
rect 1870 3263 1876 3264
rect 1870 3259 1871 3263
rect 1875 3259 1876 3263
rect 3590 3263 3596 3264
rect 1870 3258 1876 3259
rect 1926 3260 1932 3261
rect 1926 3256 1927 3260
rect 1931 3256 1932 3260
rect 1926 3255 1932 3256
rect 2062 3260 2068 3261
rect 2062 3256 2063 3260
rect 2067 3256 2068 3260
rect 2062 3255 2068 3256
rect 2198 3260 2204 3261
rect 2198 3256 2199 3260
rect 2203 3256 2204 3260
rect 2198 3255 2204 3256
rect 2358 3260 2364 3261
rect 2358 3256 2359 3260
rect 2363 3256 2364 3260
rect 2358 3255 2364 3256
rect 2542 3260 2548 3261
rect 2542 3256 2543 3260
rect 2547 3256 2548 3260
rect 2542 3255 2548 3256
rect 2758 3260 2764 3261
rect 2758 3256 2759 3260
rect 2763 3256 2764 3260
rect 2758 3255 2764 3256
rect 2998 3260 3004 3261
rect 2998 3256 2999 3260
rect 3003 3256 3004 3260
rect 2998 3255 3004 3256
rect 3246 3260 3252 3261
rect 3246 3256 3247 3260
rect 3251 3256 3252 3260
rect 3246 3255 3252 3256
rect 3502 3260 3508 3261
rect 3502 3256 3503 3260
rect 3507 3256 3508 3260
rect 3590 3259 3591 3263
rect 3595 3259 3596 3263
rect 3590 3258 3596 3259
rect 3502 3255 3508 3256
rect 382 3240 388 3241
rect 110 3237 116 3238
rect 110 3233 111 3237
rect 115 3233 116 3237
rect 382 3236 383 3240
rect 387 3236 388 3240
rect 382 3235 388 3236
rect 470 3240 476 3241
rect 470 3236 471 3240
rect 475 3236 476 3240
rect 470 3235 476 3236
rect 574 3240 580 3241
rect 574 3236 575 3240
rect 579 3236 580 3240
rect 574 3235 580 3236
rect 686 3240 692 3241
rect 686 3236 687 3240
rect 691 3236 692 3240
rect 686 3235 692 3236
rect 806 3240 812 3241
rect 806 3236 807 3240
rect 811 3236 812 3240
rect 806 3235 812 3236
rect 934 3240 940 3241
rect 934 3236 935 3240
rect 939 3236 940 3240
rect 934 3235 940 3236
rect 1062 3240 1068 3241
rect 1062 3236 1063 3240
rect 1067 3236 1068 3240
rect 1062 3235 1068 3236
rect 1190 3240 1196 3241
rect 1190 3236 1191 3240
rect 1195 3236 1196 3240
rect 1190 3235 1196 3236
rect 1318 3240 1324 3241
rect 1318 3236 1319 3240
rect 1323 3236 1324 3240
rect 1318 3235 1324 3236
rect 1446 3240 1452 3241
rect 1446 3236 1447 3240
rect 1451 3236 1452 3240
rect 1446 3235 1452 3236
rect 1574 3240 1580 3241
rect 1574 3236 1575 3240
rect 1579 3236 1580 3240
rect 1574 3235 1580 3236
rect 1830 3237 1836 3238
rect 110 3232 116 3233
rect 1830 3233 1831 3237
rect 1835 3233 1836 3237
rect 1830 3232 1836 3233
rect 110 3220 116 3221
rect 110 3216 111 3220
rect 115 3216 116 3220
rect 110 3215 116 3216
rect 1830 3220 1836 3221
rect 1830 3216 1831 3220
rect 1835 3216 1836 3220
rect 1830 3215 1836 3216
rect 1894 3212 1900 3213
rect 1870 3209 1876 3210
rect 1870 3205 1871 3209
rect 1875 3205 1876 3209
rect 1894 3208 1895 3212
rect 1899 3208 1900 3212
rect 1894 3207 1900 3208
rect 2006 3212 2012 3213
rect 2006 3208 2007 3212
rect 2011 3208 2012 3212
rect 2006 3207 2012 3208
rect 2142 3212 2148 3213
rect 2142 3208 2143 3212
rect 2147 3208 2148 3212
rect 2142 3207 2148 3208
rect 2278 3212 2284 3213
rect 2278 3208 2279 3212
rect 2283 3208 2284 3212
rect 2278 3207 2284 3208
rect 2414 3212 2420 3213
rect 2414 3208 2415 3212
rect 2419 3208 2420 3212
rect 2414 3207 2420 3208
rect 2566 3212 2572 3213
rect 2566 3208 2567 3212
rect 2571 3208 2572 3212
rect 2566 3207 2572 3208
rect 2726 3212 2732 3213
rect 2726 3208 2727 3212
rect 2731 3208 2732 3212
rect 2726 3207 2732 3208
rect 2910 3212 2916 3213
rect 2910 3208 2911 3212
rect 2915 3208 2916 3212
rect 2910 3207 2916 3208
rect 3102 3212 3108 3213
rect 3102 3208 3103 3212
rect 3107 3208 3108 3212
rect 3102 3207 3108 3208
rect 3310 3212 3316 3213
rect 3310 3208 3311 3212
rect 3315 3208 3316 3212
rect 3310 3207 3316 3208
rect 3502 3212 3508 3213
rect 3502 3208 3503 3212
rect 3507 3208 3508 3212
rect 3502 3207 3508 3208
rect 3590 3209 3596 3210
rect 1870 3204 1876 3205
rect 3590 3205 3591 3209
rect 3595 3205 3596 3209
rect 3590 3204 3596 3205
rect 390 3202 396 3203
rect 390 3198 391 3202
rect 395 3198 396 3202
rect 390 3197 396 3198
rect 478 3202 484 3203
rect 478 3198 479 3202
rect 483 3198 484 3202
rect 478 3197 484 3198
rect 582 3202 588 3203
rect 582 3198 583 3202
rect 587 3198 588 3202
rect 582 3197 588 3198
rect 694 3202 700 3203
rect 694 3198 695 3202
rect 699 3198 700 3202
rect 694 3197 700 3198
rect 814 3202 820 3203
rect 814 3198 815 3202
rect 819 3198 820 3202
rect 814 3197 820 3198
rect 942 3202 948 3203
rect 942 3198 943 3202
rect 947 3198 948 3202
rect 942 3197 948 3198
rect 1070 3202 1076 3203
rect 1070 3198 1071 3202
rect 1075 3198 1076 3202
rect 1070 3197 1076 3198
rect 1198 3202 1204 3203
rect 1198 3198 1199 3202
rect 1203 3198 1204 3202
rect 1198 3197 1204 3198
rect 1326 3202 1332 3203
rect 1326 3198 1327 3202
rect 1331 3198 1332 3202
rect 1326 3197 1332 3198
rect 1454 3202 1460 3203
rect 1454 3198 1455 3202
rect 1459 3198 1460 3202
rect 1454 3197 1460 3198
rect 1582 3202 1588 3203
rect 1582 3198 1583 3202
rect 1587 3198 1588 3202
rect 1582 3197 1588 3198
rect 1870 3192 1876 3193
rect 1870 3188 1871 3192
rect 1875 3188 1876 3192
rect 1870 3187 1876 3188
rect 3590 3192 3596 3193
rect 3590 3188 3591 3192
rect 3595 3188 3596 3192
rect 3590 3187 3596 3188
rect 1902 3174 1908 3175
rect 1902 3170 1903 3174
rect 1907 3170 1908 3174
rect 1902 3169 1908 3170
rect 2014 3174 2020 3175
rect 2014 3170 2015 3174
rect 2019 3170 2020 3174
rect 2014 3169 2020 3170
rect 2150 3174 2156 3175
rect 2150 3170 2151 3174
rect 2155 3170 2156 3174
rect 2150 3169 2156 3170
rect 2286 3174 2292 3175
rect 2286 3170 2287 3174
rect 2291 3170 2292 3174
rect 2286 3169 2292 3170
rect 2422 3174 2428 3175
rect 2422 3170 2423 3174
rect 2427 3170 2428 3174
rect 2422 3169 2428 3170
rect 2574 3174 2580 3175
rect 2574 3170 2575 3174
rect 2579 3170 2580 3174
rect 2574 3169 2580 3170
rect 2734 3174 2740 3175
rect 2734 3170 2735 3174
rect 2739 3170 2740 3174
rect 2734 3169 2740 3170
rect 2918 3174 2924 3175
rect 2918 3170 2919 3174
rect 2923 3170 2924 3174
rect 2918 3169 2924 3170
rect 3110 3174 3116 3175
rect 3110 3170 3111 3174
rect 3115 3170 3116 3174
rect 3110 3169 3116 3170
rect 3318 3174 3324 3175
rect 3318 3170 3319 3174
rect 3323 3170 3324 3174
rect 3318 3169 3324 3170
rect 3510 3174 3516 3175
rect 3510 3170 3511 3174
rect 3515 3170 3516 3174
rect 3510 3169 3516 3170
rect 382 3162 388 3163
rect 382 3158 383 3162
rect 387 3158 388 3162
rect 382 3157 388 3158
rect 462 3162 468 3163
rect 462 3158 463 3162
rect 467 3158 468 3162
rect 462 3157 468 3158
rect 542 3162 548 3163
rect 542 3158 543 3162
rect 547 3158 548 3162
rect 542 3157 548 3158
rect 622 3162 628 3163
rect 622 3158 623 3162
rect 627 3158 628 3162
rect 622 3157 628 3158
rect 710 3162 716 3163
rect 710 3158 711 3162
rect 715 3158 716 3162
rect 710 3157 716 3158
rect 814 3162 820 3163
rect 814 3158 815 3162
rect 819 3158 820 3162
rect 814 3157 820 3158
rect 926 3162 932 3163
rect 926 3158 927 3162
rect 931 3158 932 3162
rect 926 3157 932 3158
rect 1038 3162 1044 3163
rect 1038 3158 1039 3162
rect 1043 3158 1044 3162
rect 1038 3157 1044 3158
rect 1158 3162 1164 3163
rect 1158 3158 1159 3162
rect 1163 3158 1164 3162
rect 1158 3157 1164 3158
rect 1270 3162 1276 3163
rect 1270 3158 1271 3162
rect 1275 3158 1276 3162
rect 1270 3157 1276 3158
rect 1382 3162 1388 3163
rect 1382 3158 1383 3162
rect 1387 3158 1388 3162
rect 1382 3157 1388 3158
rect 1494 3162 1500 3163
rect 1494 3158 1495 3162
rect 1499 3158 1500 3162
rect 1494 3157 1500 3158
rect 1614 3162 1620 3163
rect 1614 3158 1615 3162
rect 1619 3158 1620 3162
rect 1614 3157 1620 3158
rect 1734 3162 1740 3163
rect 1734 3158 1735 3162
rect 1739 3158 1740 3162
rect 1734 3157 1740 3158
rect 110 3144 116 3145
rect 110 3140 111 3144
rect 115 3140 116 3144
rect 110 3139 116 3140
rect 1830 3144 1836 3145
rect 1830 3140 1831 3144
rect 1835 3140 1836 3144
rect 1830 3139 1836 3140
rect 1902 3142 1908 3143
rect 1902 3138 1903 3142
rect 1907 3138 1908 3142
rect 1902 3137 1908 3138
rect 2078 3142 2084 3143
rect 2078 3138 2079 3142
rect 2083 3138 2084 3142
rect 2078 3137 2084 3138
rect 2270 3142 2276 3143
rect 2270 3138 2271 3142
rect 2275 3138 2276 3142
rect 2270 3137 2276 3138
rect 2454 3142 2460 3143
rect 2454 3138 2455 3142
rect 2459 3138 2460 3142
rect 2454 3137 2460 3138
rect 2622 3142 2628 3143
rect 2622 3138 2623 3142
rect 2627 3138 2628 3142
rect 2622 3137 2628 3138
rect 2782 3142 2788 3143
rect 2782 3138 2783 3142
rect 2787 3138 2788 3142
rect 2782 3137 2788 3138
rect 2934 3142 2940 3143
rect 2934 3138 2935 3142
rect 2939 3138 2940 3142
rect 2934 3137 2940 3138
rect 3078 3142 3084 3143
rect 3078 3138 3079 3142
rect 3083 3138 3084 3142
rect 3078 3137 3084 3138
rect 3230 3142 3236 3143
rect 3230 3138 3231 3142
rect 3235 3138 3236 3142
rect 3230 3137 3236 3138
rect 110 3127 116 3128
rect 110 3123 111 3127
rect 115 3123 116 3127
rect 1830 3127 1836 3128
rect 110 3122 116 3123
rect 374 3124 380 3125
rect 374 3120 375 3124
rect 379 3120 380 3124
rect 374 3119 380 3120
rect 454 3124 460 3125
rect 454 3120 455 3124
rect 459 3120 460 3124
rect 454 3119 460 3120
rect 534 3124 540 3125
rect 534 3120 535 3124
rect 539 3120 540 3124
rect 534 3119 540 3120
rect 614 3124 620 3125
rect 614 3120 615 3124
rect 619 3120 620 3124
rect 614 3119 620 3120
rect 702 3124 708 3125
rect 702 3120 703 3124
rect 707 3120 708 3124
rect 702 3119 708 3120
rect 806 3124 812 3125
rect 806 3120 807 3124
rect 811 3120 812 3124
rect 806 3119 812 3120
rect 918 3124 924 3125
rect 918 3120 919 3124
rect 923 3120 924 3124
rect 918 3119 924 3120
rect 1030 3124 1036 3125
rect 1030 3120 1031 3124
rect 1035 3120 1036 3124
rect 1030 3119 1036 3120
rect 1150 3124 1156 3125
rect 1150 3120 1151 3124
rect 1155 3120 1156 3124
rect 1150 3119 1156 3120
rect 1262 3124 1268 3125
rect 1262 3120 1263 3124
rect 1267 3120 1268 3124
rect 1262 3119 1268 3120
rect 1374 3124 1380 3125
rect 1374 3120 1375 3124
rect 1379 3120 1380 3124
rect 1374 3119 1380 3120
rect 1486 3124 1492 3125
rect 1486 3120 1487 3124
rect 1491 3120 1492 3124
rect 1486 3119 1492 3120
rect 1606 3124 1612 3125
rect 1606 3120 1607 3124
rect 1611 3120 1612 3124
rect 1606 3119 1612 3120
rect 1726 3124 1732 3125
rect 1726 3120 1727 3124
rect 1731 3120 1732 3124
rect 1830 3123 1831 3127
rect 1835 3123 1836 3127
rect 1830 3122 1836 3123
rect 1870 3124 1876 3125
rect 1726 3119 1732 3120
rect 1870 3120 1871 3124
rect 1875 3120 1876 3124
rect 1870 3119 1876 3120
rect 3590 3124 3596 3125
rect 3590 3120 3591 3124
rect 3595 3120 3596 3124
rect 3590 3119 3596 3120
rect 1870 3107 1876 3108
rect 1870 3103 1871 3107
rect 1875 3103 1876 3107
rect 3590 3107 3596 3108
rect 1870 3102 1876 3103
rect 1894 3104 1900 3105
rect 1894 3100 1895 3104
rect 1899 3100 1900 3104
rect 1894 3099 1900 3100
rect 2070 3104 2076 3105
rect 2070 3100 2071 3104
rect 2075 3100 2076 3104
rect 2070 3099 2076 3100
rect 2262 3104 2268 3105
rect 2262 3100 2263 3104
rect 2267 3100 2268 3104
rect 2262 3099 2268 3100
rect 2446 3104 2452 3105
rect 2446 3100 2447 3104
rect 2451 3100 2452 3104
rect 2446 3099 2452 3100
rect 2614 3104 2620 3105
rect 2614 3100 2615 3104
rect 2619 3100 2620 3104
rect 2614 3099 2620 3100
rect 2774 3104 2780 3105
rect 2774 3100 2775 3104
rect 2779 3100 2780 3104
rect 2774 3099 2780 3100
rect 2926 3104 2932 3105
rect 2926 3100 2927 3104
rect 2931 3100 2932 3104
rect 2926 3099 2932 3100
rect 3070 3104 3076 3105
rect 3070 3100 3071 3104
rect 3075 3100 3076 3104
rect 3070 3099 3076 3100
rect 3222 3104 3228 3105
rect 3222 3100 3223 3104
rect 3227 3100 3228 3104
rect 3590 3103 3591 3107
rect 3595 3103 3596 3107
rect 3590 3102 3596 3103
rect 3222 3099 3228 3100
rect 942 3080 948 3081
rect 110 3077 116 3078
rect 110 3073 111 3077
rect 115 3073 116 3077
rect 942 3076 943 3080
rect 947 3076 948 3080
rect 942 3075 948 3076
rect 1022 3080 1028 3081
rect 1022 3076 1023 3080
rect 1027 3076 1028 3080
rect 1022 3075 1028 3076
rect 1102 3080 1108 3081
rect 1102 3076 1103 3080
rect 1107 3076 1108 3080
rect 1102 3075 1108 3076
rect 1182 3080 1188 3081
rect 1182 3076 1183 3080
rect 1187 3076 1188 3080
rect 1182 3075 1188 3076
rect 1262 3080 1268 3081
rect 1262 3076 1263 3080
rect 1267 3076 1268 3080
rect 1262 3075 1268 3076
rect 1342 3080 1348 3081
rect 1342 3076 1343 3080
rect 1347 3076 1348 3080
rect 1342 3075 1348 3076
rect 1422 3080 1428 3081
rect 1422 3076 1423 3080
rect 1427 3076 1428 3080
rect 1422 3075 1428 3076
rect 1502 3080 1508 3081
rect 1502 3076 1503 3080
rect 1507 3076 1508 3080
rect 1502 3075 1508 3076
rect 1582 3080 1588 3081
rect 1582 3076 1583 3080
rect 1587 3076 1588 3080
rect 1582 3075 1588 3076
rect 1662 3080 1668 3081
rect 1662 3076 1663 3080
rect 1667 3076 1668 3080
rect 1662 3075 1668 3076
rect 1742 3080 1748 3081
rect 1742 3076 1743 3080
rect 1747 3076 1748 3080
rect 1742 3075 1748 3076
rect 1830 3077 1836 3078
rect 110 3072 116 3073
rect 1830 3073 1831 3077
rect 1835 3073 1836 3077
rect 1830 3072 1836 3073
rect 110 3060 116 3061
rect 110 3056 111 3060
rect 115 3056 116 3060
rect 110 3055 116 3056
rect 1830 3060 1836 3061
rect 1830 3056 1831 3060
rect 1835 3056 1836 3060
rect 1830 3055 1836 3056
rect 1990 3052 1996 3053
rect 1870 3049 1876 3050
rect 1870 3045 1871 3049
rect 1875 3045 1876 3049
rect 1990 3048 1991 3052
rect 1995 3048 1996 3052
rect 1990 3047 1996 3048
rect 2246 3052 2252 3053
rect 2246 3048 2247 3052
rect 2251 3048 2252 3052
rect 2246 3047 2252 3048
rect 2486 3052 2492 3053
rect 2486 3048 2487 3052
rect 2491 3048 2492 3052
rect 2486 3047 2492 3048
rect 2702 3052 2708 3053
rect 2702 3048 2703 3052
rect 2707 3048 2708 3052
rect 2702 3047 2708 3048
rect 2894 3052 2900 3053
rect 2894 3048 2895 3052
rect 2899 3048 2900 3052
rect 2894 3047 2900 3048
rect 3062 3052 3068 3053
rect 3062 3048 3063 3052
rect 3067 3048 3068 3052
rect 3062 3047 3068 3048
rect 3222 3052 3228 3053
rect 3222 3048 3223 3052
rect 3227 3048 3228 3052
rect 3222 3047 3228 3048
rect 3374 3052 3380 3053
rect 3374 3048 3375 3052
rect 3379 3048 3380 3052
rect 3374 3047 3380 3048
rect 3502 3052 3508 3053
rect 3502 3048 3503 3052
rect 3507 3048 3508 3052
rect 3502 3047 3508 3048
rect 3590 3049 3596 3050
rect 1870 3044 1876 3045
rect 3590 3045 3591 3049
rect 3595 3045 3596 3049
rect 3590 3044 3596 3045
rect 950 3042 956 3043
rect 950 3038 951 3042
rect 955 3038 956 3042
rect 950 3037 956 3038
rect 1030 3042 1036 3043
rect 1030 3038 1031 3042
rect 1035 3038 1036 3042
rect 1030 3037 1036 3038
rect 1110 3042 1116 3043
rect 1110 3038 1111 3042
rect 1115 3038 1116 3042
rect 1110 3037 1116 3038
rect 1190 3042 1196 3043
rect 1190 3038 1191 3042
rect 1195 3038 1196 3042
rect 1190 3037 1196 3038
rect 1270 3042 1276 3043
rect 1270 3038 1271 3042
rect 1275 3038 1276 3042
rect 1270 3037 1276 3038
rect 1350 3042 1356 3043
rect 1350 3038 1351 3042
rect 1355 3038 1356 3042
rect 1350 3037 1356 3038
rect 1430 3042 1436 3043
rect 1430 3038 1431 3042
rect 1435 3038 1436 3042
rect 1430 3037 1436 3038
rect 1510 3042 1516 3043
rect 1510 3038 1511 3042
rect 1515 3038 1516 3042
rect 1510 3037 1516 3038
rect 1590 3042 1596 3043
rect 1590 3038 1591 3042
rect 1595 3038 1596 3042
rect 1590 3037 1596 3038
rect 1670 3042 1676 3043
rect 1670 3038 1671 3042
rect 1675 3038 1676 3042
rect 1670 3037 1676 3038
rect 1750 3042 1756 3043
rect 1750 3038 1751 3042
rect 1755 3038 1756 3042
rect 1750 3037 1756 3038
rect 1870 3032 1876 3033
rect 1870 3028 1871 3032
rect 1875 3028 1876 3032
rect 1870 3027 1876 3028
rect 3590 3032 3596 3033
rect 3590 3028 3591 3032
rect 3595 3028 3596 3032
rect 3590 3027 3596 3028
rect 1998 3014 2004 3015
rect 1998 3010 1999 3014
rect 2003 3010 2004 3014
rect 1998 3009 2004 3010
rect 2254 3014 2260 3015
rect 2254 3010 2255 3014
rect 2259 3010 2260 3014
rect 2254 3009 2260 3010
rect 2494 3014 2500 3015
rect 2494 3010 2495 3014
rect 2499 3010 2500 3014
rect 2494 3009 2500 3010
rect 2710 3014 2716 3015
rect 2710 3010 2711 3014
rect 2715 3010 2716 3014
rect 2710 3009 2716 3010
rect 2902 3014 2908 3015
rect 2902 3010 2903 3014
rect 2907 3010 2908 3014
rect 2902 3009 2908 3010
rect 3070 3014 3076 3015
rect 3070 3010 3071 3014
rect 3075 3010 3076 3014
rect 3070 3009 3076 3010
rect 3230 3014 3236 3015
rect 3230 3010 3231 3014
rect 3235 3010 3236 3014
rect 3230 3009 3236 3010
rect 3382 3014 3388 3015
rect 3382 3010 3383 3014
rect 3387 3010 3388 3014
rect 3382 3009 3388 3010
rect 3510 3014 3516 3015
rect 3510 3010 3511 3014
rect 3515 3010 3516 3014
rect 3510 3009 3516 3010
rect 206 2994 212 2995
rect 206 2990 207 2994
rect 211 2990 212 2994
rect 206 2989 212 2990
rect 326 2994 332 2995
rect 326 2990 327 2994
rect 331 2990 332 2994
rect 326 2989 332 2990
rect 470 2994 476 2995
rect 470 2990 471 2994
rect 475 2990 476 2994
rect 470 2989 476 2990
rect 630 2994 636 2995
rect 630 2990 631 2994
rect 635 2990 636 2994
rect 630 2989 636 2990
rect 806 2994 812 2995
rect 806 2990 807 2994
rect 811 2990 812 2994
rect 806 2989 812 2990
rect 982 2994 988 2995
rect 982 2990 983 2994
rect 987 2990 988 2994
rect 982 2989 988 2990
rect 1150 2994 1156 2995
rect 1150 2990 1151 2994
rect 1155 2990 1156 2994
rect 1150 2989 1156 2990
rect 1310 2994 1316 2995
rect 1310 2990 1311 2994
rect 1315 2990 1316 2994
rect 1310 2989 1316 2990
rect 1462 2994 1468 2995
rect 1462 2990 1463 2994
rect 1467 2990 1468 2994
rect 1462 2989 1468 2990
rect 1614 2994 1620 2995
rect 1614 2990 1615 2994
rect 1619 2990 1620 2994
rect 1614 2989 1620 2990
rect 1750 2994 1756 2995
rect 1750 2990 1751 2994
rect 1755 2990 1756 2994
rect 1750 2989 1756 2990
rect 1902 2978 1908 2979
rect 110 2976 116 2977
rect 110 2972 111 2976
rect 115 2972 116 2976
rect 110 2971 116 2972
rect 1830 2976 1836 2977
rect 1830 2972 1831 2976
rect 1835 2972 1836 2976
rect 1902 2974 1903 2978
rect 1907 2974 1908 2978
rect 1902 2973 1908 2974
rect 2142 2978 2148 2979
rect 2142 2974 2143 2978
rect 2147 2974 2148 2978
rect 2142 2973 2148 2974
rect 2390 2978 2396 2979
rect 2390 2974 2391 2978
rect 2395 2974 2396 2978
rect 2390 2973 2396 2974
rect 2606 2978 2612 2979
rect 2606 2974 2607 2978
rect 2611 2974 2612 2978
rect 2606 2973 2612 2974
rect 2798 2978 2804 2979
rect 2798 2974 2799 2978
rect 2803 2974 2804 2978
rect 2798 2973 2804 2974
rect 2966 2978 2972 2979
rect 2966 2974 2967 2978
rect 2971 2974 2972 2978
rect 2966 2973 2972 2974
rect 3118 2978 3124 2979
rect 3118 2974 3119 2978
rect 3123 2974 3124 2978
rect 3118 2973 3124 2974
rect 3262 2978 3268 2979
rect 3262 2974 3263 2978
rect 3267 2974 3268 2978
rect 3262 2973 3268 2974
rect 3398 2978 3404 2979
rect 3398 2974 3399 2978
rect 3403 2974 3404 2978
rect 3398 2973 3404 2974
rect 3510 2978 3516 2979
rect 3510 2974 3511 2978
rect 3515 2974 3516 2978
rect 3510 2973 3516 2974
rect 1830 2971 1836 2972
rect 1870 2960 1876 2961
rect 110 2959 116 2960
rect 110 2955 111 2959
rect 115 2955 116 2959
rect 1830 2959 1836 2960
rect 110 2954 116 2955
rect 198 2956 204 2957
rect 198 2952 199 2956
rect 203 2952 204 2956
rect 198 2951 204 2952
rect 318 2956 324 2957
rect 318 2952 319 2956
rect 323 2952 324 2956
rect 318 2951 324 2952
rect 462 2956 468 2957
rect 462 2952 463 2956
rect 467 2952 468 2956
rect 462 2951 468 2952
rect 622 2956 628 2957
rect 622 2952 623 2956
rect 627 2952 628 2956
rect 622 2951 628 2952
rect 798 2956 804 2957
rect 798 2952 799 2956
rect 803 2952 804 2956
rect 798 2951 804 2952
rect 974 2956 980 2957
rect 974 2952 975 2956
rect 979 2952 980 2956
rect 974 2951 980 2952
rect 1142 2956 1148 2957
rect 1142 2952 1143 2956
rect 1147 2952 1148 2956
rect 1142 2951 1148 2952
rect 1302 2956 1308 2957
rect 1302 2952 1303 2956
rect 1307 2952 1308 2956
rect 1302 2951 1308 2952
rect 1454 2956 1460 2957
rect 1454 2952 1455 2956
rect 1459 2952 1460 2956
rect 1454 2951 1460 2952
rect 1606 2956 1612 2957
rect 1606 2952 1607 2956
rect 1611 2952 1612 2956
rect 1606 2951 1612 2952
rect 1742 2956 1748 2957
rect 1742 2952 1743 2956
rect 1747 2952 1748 2956
rect 1830 2955 1831 2959
rect 1835 2955 1836 2959
rect 1870 2956 1871 2960
rect 1875 2956 1876 2960
rect 1870 2955 1876 2956
rect 3590 2960 3596 2961
rect 3590 2956 3591 2960
rect 3595 2956 3596 2960
rect 3590 2955 3596 2956
rect 1830 2954 1836 2955
rect 1742 2951 1748 2952
rect 1870 2943 1876 2944
rect 1870 2939 1871 2943
rect 1875 2939 1876 2943
rect 3590 2943 3596 2944
rect 1870 2938 1876 2939
rect 1894 2940 1900 2941
rect 1894 2936 1895 2940
rect 1899 2936 1900 2940
rect 1894 2935 1900 2936
rect 2134 2940 2140 2941
rect 2134 2936 2135 2940
rect 2139 2936 2140 2940
rect 2134 2935 2140 2936
rect 2382 2940 2388 2941
rect 2382 2936 2383 2940
rect 2387 2936 2388 2940
rect 2382 2935 2388 2936
rect 2598 2940 2604 2941
rect 2598 2936 2599 2940
rect 2603 2936 2604 2940
rect 2598 2935 2604 2936
rect 2790 2940 2796 2941
rect 2790 2936 2791 2940
rect 2795 2936 2796 2940
rect 2790 2935 2796 2936
rect 2958 2940 2964 2941
rect 2958 2936 2959 2940
rect 2963 2936 2964 2940
rect 2958 2935 2964 2936
rect 3110 2940 3116 2941
rect 3110 2936 3111 2940
rect 3115 2936 3116 2940
rect 3110 2935 3116 2936
rect 3254 2940 3260 2941
rect 3254 2936 3255 2940
rect 3259 2936 3260 2940
rect 3254 2935 3260 2936
rect 3390 2940 3396 2941
rect 3390 2936 3391 2940
rect 3395 2936 3396 2940
rect 3390 2935 3396 2936
rect 3502 2940 3508 2941
rect 3502 2936 3503 2940
rect 3507 2936 3508 2940
rect 3590 2939 3591 2943
rect 3595 2939 3596 2943
rect 3590 2938 3596 2939
rect 3502 2935 3508 2936
rect 246 2912 252 2913
rect 110 2909 116 2910
rect 110 2905 111 2909
rect 115 2905 116 2909
rect 246 2908 247 2912
rect 251 2908 252 2912
rect 246 2907 252 2908
rect 350 2912 356 2913
rect 350 2908 351 2912
rect 355 2908 356 2912
rect 350 2907 356 2908
rect 470 2912 476 2913
rect 470 2908 471 2912
rect 475 2908 476 2912
rect 470 2907 476 2908
rect 606 2912 612 2913
rect 606 2908 607 2912
rect 611 2908 612 2912
rect 606 2907 612 2908
rect 750 2912 756 2913
rect 750 2908 751 2912
rect 755 2908 756 2912
rect 750 2907 756 2908
rect 894 2912 900 2913
rect 894 2908 895 2912
rect 899 2908 900 2912
rect 894 2907 900 2908
rect 1030 2912 1036 2913
rect 1030 2908 1031 2912
rect 1035 2908 1036 2912
rect 1030 2907 1036 2908
rect 1158 2912 1164 2913
rect 1158 2908 1159 2912
rect 1163 2908 1164 2912
rect 1158 2907 1164 2908
rect 1278 2912 1284 2913
rect 1278 2908 1279 2912
rect 1283 2908 1284 2912
rect 1278 2907 1284 2908
rect 1398 2912 1404 2913
rect 1398 2908 1399 2912
rect 1403 2908 1404 2912
rect 1398 2907 1404 2908
rect 1518 2912 1524 2913
rect 1518 2908 1519 2912
rect 1523 2908 1524 2912
rect 1518 2907 1524 2908
rect 1638 2912 1644 2913
rect 1638 2908 1639 2912
rect 1643 2908 1644 2912
rect 1638 2907 1644 2908
rect 1830 2909 1836 2910
rect 110 2904 116 2905
rect 1830 2905 1831 2909
rect 1835 2905 1836 2909
rect 1830 2904 1836 2905
rect 110 2892 116 2893
rect 110 2888 111 2892
rect 115 2888 116 2892
rect 110 2887 116 2888
rect 1830 2892 1836 2893
rect 1830 2888 1831 2892
rect 1835 2888 1836 2892
rect 1830 2887 1836 2888
rect 2350 2884 2356 2885
rect 1870 2881 1876 2882
rect 1870 2877 1871 2881
rect 1875 2877 1876 2881
rect 2350 2880 2351 2884
rect 2355 2880 2356 2884
rect 2350 2879 2356 2880
rect 2446 2884 2452 2885
rect 2446 2880 2447 2884
rect 2451 2880 2452 2884
rect 2446 2879 2452 2880
rect 2550 2884 2556 2885
rect 2550 2880 2551 2884
rect 2555 2880 2556 2884
rect 2550 2879 2556 2880
rect 2654 2884 2660 2885
rect 2654 2880 2655 2884
rect 2659 2880 2660 2884
rect 2654 2879 2660 2880
rect 2758 2884 2764 2885
rect 2758 2880 2759 2884
rect 2763 2880 2764 2884
rect 2758 2879 2764 2880
rect 2870 2884 2876 2885
rect 2870 2880 2871 2884
rect 2875 2880 2876 2884
rect 2870 2879 2876 2880
rect 2982 2884 2988 2885
rect 2982 2880 2983 2884
rect 2987 2880 2988 2884
rect 2982 2879 2988 2880
rect 3094 2884 3100 2885
rect 3094 2880 3095 2884
rect 3099 2880 3100 2884
rect 3094 2879 3100 2880
rect 3206 2884 3212 2885
rect 3206 2880 3207 2884
rect 3211 2880 3212 2884
rect 3206 2879 3212 2880
rect 3590 2881 3596 2882
rect 1870 2876 1876 2877
rect 3590 2877 3591 2881
rect 3595 2877 3596 2881
rect 3590 2876 3596 2877
rect 254 2874 260 2875
rect 254 2870 255 2874
rect 259 2870 260 2874
rect 254 2869 260 2870
rect 358 2874 364 2875
rect 358 2870 359 2874
rect 363 2870 364 2874
rect 358 2869 364 2870
rect 478 2874 484 2875
rect 478 2870 479 2874
rect 483 2870 484 2874
rect 478 2869 484 2870
rect 614 2874 620 2875
rect 614 2870 615 2874
rect 619 2870 620 2874
rect 614 2869 620 2870
rect 758 2874 764 2875
rect 758 2870 759 2874
rect 763 2870 764 2874
rect 758 2869 764 2870
rect 902 2874 908 2875
rect 902 2870 903 2874
rect 907 2870 908 2874
rect 902 2869 908 2870
rect 1038 2874 1044 2875
rect 1038 2870 1039 2874
rect 1043 2870 1044 2874
rect 1038 2869 1044 2870
rect 1166 2874 1172 2875
rect 1166 2870 1167 2874
rect 1171 2870 1172 2874
rect 1166 2869 1172 2870
rect 1286 2874 1292 2875
rect 1286 2870 1287 2874
rect 1291 2870 1292 2874
rect 1286 2869 1292 2870
rect 1406 2874 1412 2875
rect 1406 2870 1407 2874
rect 1411 2870 1412 2874
rect 1406 2869 1412 2870
rect 1526 2874 1532 2875
rect 1526 2870 1527 2874
rect 1531 2870 1532 2874
rect 1526 2869 1532 2870
rect 1646 2874 1652 2875
rect 1646 2870 1647 2874
rect 1651 2870 1652 2874
rect 1646 2869 1652 2870
rect 1870 2864 1876 2865
rect 1870 2860 1871 2864
rect 1875 2860 1876 2864
rect 1870 2859 1876 2860
rect 3590 2864 3596 2865
rect 3590 2860 3591 2864
rect 3595 2860 3596 2864
rect 3590 2859 3596 2860
rect 2358 2846 2364 2847
rect 150 2842 156 2843
rect 150 2838 151 2842
rect 155 2838 156 2842
rect 150 2837 156 2838
rect 278 2842 284 2843
rect 278 2838 279 2842
rect 283 2838 284 2842
rect 278 2837 284 2838
rect 406 2842 412 2843
rect 406 2838 407 2842
rect 411 2838 412 2842
rect 406 2837 412 2838
rect 542 2842 548 2843
rect 542 2838 543 2842
rect 547 2838 548 2842
rect 542 2837 548 2838
rect 670 2842 676 2843
rect 670 2838 671 2842
rect 675 2838 676 2842
rect 670 2837 676 2838
rect 798 2842 804 2843
rect 798 2838 799 2842
rect 803 2838 804 2842
rect 798 2837 804 2838
rect 918 2842 924 2843
rect 918 2838 919 2842
rect 923 2838 924 2842
rect 918 2837 924 2838
rect 1038 2842 1044 2843
rect 1038 2838 1039 2842
rect 1043 2838 1044 2842
rect 1038 2837 1044 2838
rect 1150 2842 1156 2843
rect 1150 2838 1151 2842
rect 1155 2838 1156 2842
rect 1150 2837 1156 2838
rect 1270 2842 1276 2843
rect 1270 2838 1271 2842
rect 1275 2838 1276 2842
rect 1270 2837 1276 2838
rect 1390 2842 1396 2843
rect 1390 2838 1391 2842
rect 1395 2838 1396 2842
rect 2358 2842 2359 2846
rect 2363 2842 2364 2846
rect 2358 2841 2364 2842
rect 2454 2846 2460 2847
rect 2454 2842 2455 2846
rect 2459 2842 2460 2846
rect 2454 2841 2460 2842
rect 2558 2846 2564 2847
rect 2558 2842 2559 2846
rect 2563 2842 2564 2846
rect 2558 2841 2564 2842
rect 2662 2846 2668 2847
rect 2662 2842 2663 2846
rect 2667 2842 2668 2846
rect 2662 2841 2668 2842
rect 2766 2846 2772 2847
rect 2766 2842 2767 2846
rect 2771 2842 2772 2846
rect 2766 2841 2772 2842
rect 2878 2846 2884 2847
rect 2878 2842 2879 2846
rect 2883 2842 2884 2846
rect 2878 2841 2884 2842
rect 2990 2846 2996 2847
rect 2990 2842 2991 2846
rect 2995 2842 2996 2846
rect 2990 2841 2996 2842
rect 3102 2846 3108 2847
rect 3102 2842 3103 2846
rect 3107 2842 3108 2846
rect 3102 2841 3108 2842
rect 3214 2846 3220 2847
rect 3214 2842 3215 2846
rect 3219 2842 3220 2846
rect 3214 2841 3220 2842
rect 1390 2837 1396 2838
rect 110 2824 116 2825
rect 110 2820 111 2824
rect 115 2820 116 2824
rect 110 2819 116 2820
rect 1830 2824 1836 2825
rect 1830 2820 1831 2824
rect 1835 2820 1836 2824
rect 1830 2819 1836 2820
rect 2238 2814 2244 2815
rect 2238 2810 2239 2814
rect 2243 2810 2244 2814
rect 2238 2809 2244 2810
rect 2318 2814 2324 2815
rect 2318 2810 2319 2814
rect 2323 2810 2324 2814
rect 2318 2809 2324 2810
rect 2398 2814 2404 2815
rect 2398 2810 2399 2814
rect 2403 2810 2404 2814
rect 2398 2809 2404 2810
rect 2478 2814 2484 2815
rect 2478 2810 2479 2814
rect 2483 2810 2484 2814
rect 2478 2809 2484 2810
rect 2566 2814 2572 2815
rect 2566 2810 2567 2814
rect 2571 2810 2572 2814
rect 2566 2809 2572 2810
rect 2670 2814 2676 2815
rect 2670 2810 2671 2814
rect 2675 2810 2676 2814
rect 2670 2809 2676 2810
rect 2806 2814 2812 2815
rect 2806 2810 2807 2814
rect 2811 2810 2812 2814
rect 2806 2809 2812 2810
rect 2966 2814 2972 2815
rect 2966 2810 2967 2814
rect 2971 2810 2972 2814
rect 2966 2809 2972 2810
rect 3142 2814 3148 2815
rect 3142 2810 3143 2814
rect 3147 2810 3148 2814
rect 3142 2809 3148 2810
rect 3334 2814 3340 2815
rect 3334 2810 3335 2814
rect 3339 2810 3340 2814
rect 3334 2809 3340 2810
rect 3510 2814 3516 2815
rect 3510 2810 3511 2814
rect 3515 2810 3516 2814
rect 3510 2809 3516 2810
rect 110 2807 116 2808
rect 110 2803 111 2807
rect 115 2803 116 2807
rect 1830 2807 1836 2808
rect 110 2802 116 2803
rect 142 2804 148 2805
rect 142 2800 143 2804
rect 147 2800 148 2804
rect 142 2799 148 2800
rect 270 2804 276 2805
rect 270 2800 271 2804
rect 275 2800 276 2804
rect 270 2799 276 2800
rect 398 2804 404 2805
rect 398 2800 399 2804
rect 403 2800 404 2804
rect 398 2799 404 2800
rect 534 2804 540 2805
rect 534 2800 535 2804
rect 539 2800 540 2804
rect 534 2799 540 2800
rect 662 2804 668 2805
rect 662 2800 663 2804
rect 667 2800 668 2804
rect 662 2799 668 2800
rect 790 2804 796 2805
rect 790 2800 791 2804
rect 795 2800 796 2804
rect 790 2799 796 2800
rect 910 2804 916 2805
rect 910 2800 911 2804
rect 915 2800 916 2804
rect 910 2799 916 2800
rect 1030 2804 1036 2805
rect 1030 2800 1031 2804
rect 1035 2800 1036 2804
rect 1030 2799 1036 2800
rect 1142 2804 1148 2805
rect 1142 2800 1143 2804
rect 1147 2800 1148 2804
rect 1142 2799 1148 2800
rect 1262 2804 1268 2805
rect 1262 2800 1263 2804
rect 1267 2800 1268 2804
rect 1262 2799 1268 2800
rect 1382 2804 1388 2805
rect 1382 2800 1383 2804
rect 1387 2800 1388 2804
rect 1830 2803 1831 2807
rect 1835 2803 1836 2807
rect 1830 2802 1836 2803
rect 1382 2799 1388 2800
rect 1870 2796 1876 2797
rect 1870 2792 1871 2796
rect 1875 2792 1876 2796
rect 1870 2791 1876 2792
rect 3590 2796 3596 2797
rect 3590 2792 3591 2796
rect 3595 2792 3596 2796
rect 3590 2791 3596 2792
rect 1870 2779 1876 2780
rect 1870 2775 1871 2779
rect 1875 2775 1876 2779
rect 3590 2779 3596 2780
rect 1870 2774 1876 2775
rect 2230 2776 2236 2777
rect 2230 2772 2231 2776
rect 2235 2772 2236 2776
rect 2230 2771 2236 2772
rect 2310 2776 2316 2777
rect 2310 2772 2311 2776
rect 2315 2772 2316 2776
rect 2310 2771 2316 2772
rect 2390 2776 2396 2777
rect 2390 2772 2391 2776
rect 2395 2772 2396 2776
rect 2390 2771 2396 2772
rect 2470 2776 2476 2777
rect 2470 2772 2471 2776
rect 2475 2772 2476 2776
rect 2470 2771 2476 2772
rect 2558 2776 2564 2777
rect 2558 2772 2559 2776
rect 2563 2772 2564 2776
rect 2558 2771 2564 2772
rect 2662 2776 2668 2777
rect 2662 2772 2663 2776
rect 2667 2772 2668 2776
rect 2662 2771 2668 2772
rect 2798 2776 2804 2777
rect 2798 2772 2799 2776
rect 2803 2772 2804 2776
rect 2798 2771 2804 2772
rect 2958 2776 2964 2777
rect 2958 2772 2959 2776
rect 2963 2772 2964 2776
rect 2958 2771 2964 2772
rect 3134 2776 3140 2777
rect 3134 2772 3135 2776
rect 3139 2772 3140 2776
rect 3134 2771 3140 2772
rect 3326 2776 3332 2777
rect 3326 2772 3327 2776
rect 3331 2772 3332 2776
rect 3326 2771 3332 2772
rect 3502 2776 3508 2777
rect 3502 2772 3503 2776
rect 3507 2772 3508 2776
rect 3590 2775 3591 2779
rect 3595 2775 3596 2779
rect 3590 2774 3596 2775
rect 3502 2771 3508 2772
rect 142 2752 148 2753
rect 110 2749 116 2750
rect 110 2745 111 2749
rect 115 2745 116 2749
rect 142 2748 143 2752
rect 147 2748 148 2752
rect 142 2747 148 2748
rect 294 2752 300 2753
rect 294 2748 295 2752
rect 299 2748 300 2752
rect 294 2747 300 2748
rect 438 2752 444 2753
rect 438 2748 439 2752
rect 443 2748 444 2752
rect 438 2747 444 2748
rect 566 2752 572 2753
rect 566 2748 567 2752
rect 571 2748 572 2752
rect 566 2747 572 2748
rect 686 2752 692 2753
rect 686 2748 687 2752
rect 691 2748 692 2752
rect 686 2747 692 2748
rect 798 2752 804 2753
rect 798 2748 799 2752
rect 803 2748 804 2752
rect 798 2747 804 2748
rect 902 2752 908 2753
rect 902 2748 903 2752
rect 907 2748 908 2752
rect 902 2747 908 2748
rect 1006 2752 1012 2753
rect 1006 2748 1007 2752
rect 1011 2748 1012 2752
rect 1006 2747 1012 2748
rect 1102 2752 1108 2753
rect 1102 2748 1103 2752
rect 1107 2748 1108 2752
rect 1102 2747 1108 2748
rect 1198 2752 1204 2753
rect 1198 2748 1199 2752
rect 1203 2748 1204 2752
rect 1198 2747 1204 2748
rect 1302 2752 1308 2753
rect 1302 2748 1303 2752
rect 1307 2748 1308 2752
rect 1302 2747 1308 2748
rect 1830 2749 1836 2750
rect 110 2744 116 2745
rect 1830 2745 1831 2749
rect 1835 2745 1836 2749
rect 1830 2744 1836 2745
rect 110 2732 116 2733
rect 110 2728 111 2732
rect 115 2728 116 2732
rect 110 2727 116 2728
rect 1830 2732 1836 2733
rect 1830 2728 1831 2732
rect 1835 2728 1836 2732
rect 1830 2727 1836 2728
rect 2046 2720 2052 2721
rect 1870 2717 1876 2718
rect 150 2714 156 2715
rect 150 2710 151 2714
rect 155 2710 156 2714
rect 150 2709 156 2710
rect 302 2714 308 2715
rect 302 2710 303 2714
rect 307 2710 308 2714
rect 302 2709 308 2710
rect 446 2714 452 2715
rect 446 2710 447 2714
rect 451 2710 452 2714
rect 446 2709 452 2710
rect 574 2714 580 2715
rect 574 2710 575 2714
rect 579 2710 580 2714
rect 574 2709 580 2710
rect 694 2714 700 2715
rect 694 2710 695 2714
rect 699 2710 700 2714
rect 694 2709 700 2710
rect 806 2714 812 2715
rect 806 2710 807 2714
rect 811 2710 812 2714
rect 806 2709 812 2710
rect 910 2714 916 2715
rect 910 2710 911 2714
rect 915 2710 916 2714
rect 910 2709 916 2710
rect 1014 2714 1020 2715
rect 1014 2710 1015 2714
rect 1019 2710 1020 2714
rect 1014 2709 1020 2710
rect 1110 2714 1116 2715
rect 1110 2710 1111 2714
rect 1115 2710 1116 2714
rect 1110 2709 1116 2710
rect 1206 2714 1212 2715
rect 1206 2710 1207 2714
rect 1211 2710 1212 2714
rect 1206 2709 1212 2710
rect 1310 2714 1316 2715
rect 1310 2710 1311 2714
rect 1315 2710 1316 2714
rect 1870 2713 1871 2717
rect 1875 2713 1876 2717
rect 2046 2716 2047 2720
rect 2051 2716 2052 2720
rect 2046 2715 2052 2716
rect 2134 2720 2140 2721
rect 2134 2716 2135 2720
rect 2139 2716 2140 2720
rect 2134 2715 2140 2716
rect 2230 2720 2236 2721
rect 2230 2716 2231 2720
rect 2235 2716 2236 2720
rect 2230 2715 2236 2716
rect 2326 2720 2332 2721
rect 2326 2716 2327 2720
rect 2331 2716 2332 2720
rect 2326 2715 2332 2716
rect 2422 2720 2428 2721
rect 2422 2716 2423 2720
rect 2427 2716 2428 2720
rect 2422 2715 2428 2716
rect 2518 2720 2524 2721
rect 2518 2716 2519 2720
rect 2523 2716 2524 2720
rect 2518 2715 2524 2716
rect 2614 2720 2620 2721
rect 2614 2716 2615 2720
rect 2619 2716 2620 2720
rect 2614 2715 2620 2716
rect 2726 2720 2732 2721
rect 2726 2716 2727 2720
rect 2731 2716 2732 2720
rect 2726 2715 2732 2716
rect 2854 2720 2860 2721
rect 2854 2716 2855 2720
rect 2859 2716 2860 2720
rect 2854 2715 2860 2716
rect 3006 2720 3012 2721
rect 3006 2716 3007 2720
rect 3011 2716 3012 2720
rect 3006 2715 3012 2716
rect 3174 2720 3180 2721
rect 3174 2716 3175 2720
rect 3179 2716 3180 2720
rect 3174 2715 3180 2716
rect 3350 2720 3356 2721
rect 3350 2716 3351 2720
rect 3355 2716 3356 2720
rect 3350 2715 3356 2716
rect 3502 2720 3508 2721
rect 3502 2716 3503 2720
rect 3507 2716 3508 2720
rect 3502 2715 3508 2716
rect 3590 2717 3596 2718
rect 1870 2712 1876 2713
rect 3590 2713 3591 2717
rect 3595 2713 3596 2717
rect 3590 2712 3596 2713
rect 1310 2709 1316 2710
rect 1870 2700 1876 2701
rect 1870 2696 1871 2700
rect 1875 2696 1876 2700
rect 1870 2695 1876 2696
rect 3590 2700 3596 2701
rect 3590 2696 3591 2700
rect 3595 2696 3596 2700
rect 3590 2695 3596 2696
rect 2054 2682 2060 2683
rect 142 2678 148 2679
rect 142 2674 143 2678
rect 147 2674 148 2678
rect 142 2673 148 2674
rect 262 2678 268 2679
rect 262 2674 263 2678
rect 267 2674 268 2678
rect 262 2673 268 2674
rect 406 2678 412 2679
rect 406 2674 407 2678
rect 411 2674 412 2678
rect 406 2673 412 2674
rect 542 2678 548 2679
rect 542 2674 543 2678
rect 547 2674 548 2678
rect 542 2673 548 2674
rect 670 2678 676 2679
rect 670 2674 671 2678
rect 675 2674 676 2678
rect 670 2673 676 2674
rect 790 2678 796 2679
rect 790 2674 791 2678
rect 795 2674 796 2678
rect 790 2673 796 2674
rect 902 2678 908 2679
rect 902 2674 903 2678
rect 907 2674 908 2678
rect 902 2673 908 2674
rect 1014 2678 1020 2679
rect 1014 2674 1015 2678
rect 1019 2674 1020 2678
rect 1014 2673 1020 2674
rect 1118 2678 1124 2679
rect 1118 2674 1119 2678
rect 1123 2674 1124 2678
rect 1118 2673 1124 2674
rect 1214 2678 1220 2679
rect 1214 2674 1215 2678
rect 1219 2674 1220 2678
rect 1214 2673 1220 2674
rect 1318 2678 1324 2679
rect 1318 2674 1319 2678
rect 1323 2674 1324 2678
rect 1318 2673 1324 2674
rect 1422 2678 1428 2679
rect 1422 2674 1423 2678
rect 1427 2674 1428 2678
rect 2054 2678 2055 2682
rect 2059 2678 2060 2682
rect 2054 2677 2060 2678
rect 2142 2682 2148 2683
rect 2142 2678 2143 2682
rect 2147 2678 2148 2682
rect 2142 2677 2148 2678
rect 2238 2682 2244 2683
rect 2238 2678 2239 2682
rect 2243 2678 2244 2682
rect 2238 2677 2244 2678
rect 2334 2682 2340 2683
rect 2334 2678 2335 2682
rect 2339 2678 2340 2682
rect 2334 2677 2340 2678
rect 2430 2682 2436 2683
rect 2430 2678 2431 2682
rect 2435 2678 2436 2682
rect 2430 2677 2436 2678
rect 2526 2682 2532 2683
rect 2526 2678 2527 2682
rect 2531 2678 2532 2682
rect 2526 2677 2532 2678
rect 2622 2682 2628 2683
rect 2622 2678 2623 2682
rect 2627 2678 2628 2682
rect 2622 2677 2628 2678
rect 2734 2682 2740 2683
rect 2734 2678 2735 2682
rect 2739 2678 2740 2682
rect 2734 2677 2740 2678
rect 2862 2682 2868 2683
rect 2862 2678 2863 2682
rect 2867 2678 2868 2682
rect 2862 2677 2868 2678
rect 3014 2682 3020 2683
rect 3014 2678 3015 2682
rect 3019 2678 3020 2682
rect 3014 2677 3020 2678
rect 3182 2682 3188 2683
rect 3182 2678 3183 2682
rect 3187 2678 3188 2682
rect 3182 2677 3188 2678
rect 3358 2682 3364 2683
rect 3358 2678 3359 2682
rect 3363 2678 3364 2682
rect 3358 2677 3364 2678
rect 3510 2682 3516 2683
rect 3510 2678 3511 2682
rect 3515 2678 3516 2682
rect 3510 2677 3516 2678
rect 1422 2673 1428 2674
rect 110 2660 116 2661
rect 110 2656 111 2660
rect 115 2656 116 2660
rect 110 2655 116 2656
rect 1830 2660 1836 2661
rect 1830 2656 1831 2660
rect 1835 2656 1836 2660
rect 1830 2655 1836 2656
rect 2070 2650 2076 2651
rect 2070 2646 2071 2650
rect 2075 2646 2076 2650
rect 2070 2645 2076 2646
rect 2294 2650 2300 2651
rect 2294 2646 2295 2650
rect 2299 2646 2300 2650
rect 2294 2645 2300 2646
rect 2566 2650 2572 2651
rect 2566 2646 2567 2650
rect 2571 2646 2572 2650
rect 2566 2645 2572 2646
rect 2870 2650 2876 2651
rect 2870 2646 2871 2650
rect 2875 2646 2876 2650
rect 2870 2645 2876 2646
rect 3198 2650 3204 2651
rect 3198 2646 3199 2650
rect 3203 2646 3204 2650
rect 3198 2645 3204 2646
rect 3510 2650 3516 2651
rect 3510 2646 3511 2650
rect 3515 2646 3516 2650
rect 3510 2645 3516 2646
rect 110 2643 116 2644
rect 110 2639 111 2643
rect 115 2639 116 2643
rect 1830 2643 1836 2644
rect 110 2638 116 2639
rect 134 2640 140 2641
rect 134 2636 135 2640
rect 139 2636 140 2640
rect 134 2635 140 2636
rect 254 2640 260 2641
rect 254 2636 255 2640
rect 259 2636 260 2640
rect 254 2635 260 2636
rect 398 2640 404 2641
rect 398 2636 399 2640
rect 403 2636 404 2640
rect 398 2635 404 2636
rect 534 2640 540 2641
rect 534 2636 535 2640
rect 539 2636 540 2640
rect 534 2635 540 2636
rect 662 2640 668 2641
rect 662 2636 663 2640
rect 667 2636 668 2640
rect 662 2635 668 2636
rect 782 2640 788 2641
rect 782 2636 783 2640
rect 787 2636 788 2640
rect 782 2635 788 2636
rect 894 2640 900 2641
rect 894 2636 895 2640
rect 899 2636 900 2640
rect 894 2635 900 2636
rect 1006 2640 1012 2641
rect 1006 2636 1007 2640
rect 1011 2636 1012 2640
rect 1006 2635 1012 2636
rect 1110 2640 1116 2641
rect 1110 2636 1111 2640
rect 1115 2636 1116 2640
rect 1110 2635 1116 2636
rect 1206 2640 1212 2641
rect 1206 2636 1207 2640
rect 1211 2636 1212 2640
rect 1206 2635 1212 2636
rect 1310 2640 1316 2641
rect 1310 2636 1311 2640
rect 1315 2636 1316 2640
rect 1310 2635 1316 2636
rect 1414 2640 1420 2641
rect 1414 2636 1415 2640
rect 1419 2636 1420 2640
rect 1830 2639 1831 2643
rect 1835 2639 1836 2643
rect 1830 2638 1836 2639
rect 1414 2635 1420 2636
rect 1870 2632 1876 2633
rect 1870 2628 1871 2632
rect 1875 2628 1876 2632
rect 1870 2627 1876 2628
rect 3590 2632 3596 2633
rect 3590 2628 3591 2632
rect 3595 2628 3596 2632
rect 3590 2627 3596 2628
rect 1870 2615 1876 2616
rect 1870 2611 1871 2615
rect 1875 2611 1876 2615
rect 3590 2615 3596 2616
rect 1870 2610 1876 2611
rect 2062 2612 2068 2613
rect 2062 2608 2063 2612
rect 2067 2608 2068 2612
rect 2062 2607 2068 2608
rect 2286 2612 2292 2613
rect 2286 2608 2287 2612
rect 2291 2608 2292 2612
rect 2286 2607 2292 2608
rect 2558 2612 2564 2613
rect 2558 2608 2559 2612
rect 2563 2608 2564 2612
rect 2558 2607 2564 2608
rect 2862 2612 2868 2613
rect 2862 2608 2863 2612
rect 2867 2608 2868 2612
rect 2862 2607 2868 2608
rect 3190 2612 3196 2613
rect 3190 2608 3191 2612
rect 3195 2608 3196 2612
rect 3190 2607 3196 2608
rect 3502 2612 3508 2613
rect 3502 2608 3503 2612
rect 3507 2608 3508 2612
rect 3590 2611 3591 2615
rect 3595 2611 3596 2615
rect 3590 2610 3596 2611
rect 3502 2607 3508 2608
rect 142 2588 148 2589
rect 110 2585 116 2586
rect 110 2581 111 2585
rect 115 2581 116 2585
rect 142 2584 143 2588
rect 147 2584 148 2588
rect 142 2583 148 2584
rect 310 2588 316 2589
rect 310 2584 311 2588
rect 315 2584 316 2588
rect 310 2583 316 2584
rect 478 2588 484 2589
rect 478 2584 479 2588
rect 483 2584 484 2588
rect 478 2583 484 2584
rect 638 2588 644 2589
rect 638 2584 639 2588
rect 643 2584 644 2588
rect 638 2583 644 2584
rect 790 2588 796 2589
rect 790 2584 791 2588
rect 795 2584 796 2588
rect 790 2583 796 2584
rect 926 2588 932 2589
rect 926 2584 927 2588
rect 931 2584 932 2588
rect 926 2583 932 2584
rect 1054 2588 1060 2589
rect 1054 2584 1055 2588
rect 1059 2584 1060 2588
rect 1054 2583 1060 2584
rect 1174 2588 1180 2589
rect 1174 2584 1175 2588
rect 1179 2584 1180 2588
rect 1174 2583 1180 2584
rect 1294 2588 1300 2589
rect 1294 2584 1295 2588
rect 1299 2584 1300 2588
rect 1294 2583 1300 2584
rect 1406 2588 1412 2589
rect 1406 2584 1407 2588
rect 1411 2584 1412 2588
rect 1406 2583 1412 2584
rect 1526 2588 1532 2589
rect 1526 2584 1527 2588
rect 1531 2584 1532 2588
rect 1526 2583 1532 2584
rect 1830 2585 1836 2586
rect 110 2580 116 2581
rect 1830 2581 1831 2585
rect 1835 2581 1836 2585
rect 1830 2580 1836 2581
rect 110 2568 116 2569
rect 110 2564 111 2568
rect 115 2564 116 2568
rect 110 2563 116 2564
rect 1830 2568 1836 2569
rect 1830 2564 1831 2568
rect 1835 2564 1836 2568
rect 1830 2563 1836 2564
rect 2166 2564 2172 2565
rect 1870 2561 1876 2562
rect 1870 2557 1871 2561
rect 1875 2557 1876 2561
rect 2166 2560 2167 2564
rect 2171 2560 2172 2564
rect 2166 2559 2172 2560
rect 2262 2564 2268 2565
rect 2262 2560 2263 2564
rect 2267 2560 2268 2564
rect 2262 2559 2268 2560
rect 2366 2564 2372 2565
rect 2366 2560 2367 2564
rect 2371 2560 2372 2564
rect 2366 2559 2372 2560
rect 2478 2564 2484 2565
rect 2478 2560 2479 2564
rect 2483 2560 2484 2564
rect 2478 2559 2484 2560
rect 2590 2564 2596 2565
rect 2590 2560 2591 2564
rect 2595 2560 2596 2564
rect 2590 2559 2596 2560
rect 2694 2564 2700 2565
rect 2694 2560 2695 2564
rect 2699 2560 2700 2564
rect 2694 2559 2700 2560
rect 2798 2564 2804 2565
rect 2798 2560 2799 2564
rect 2803 2560 2804 2564
rect 2798 2559 2804 2560
rect 2902 2564 2908 2565
rect 2902 2560 2903 2564
rect 2907 2560 2908 2564
rect 2902 2559 2908 2560
rect 3014 2564 3020 2565
rect 3014 2560 3015 2564
rect 3019 2560 3020 2564
rect 3014 2559 3020 2560
rect 3134 2564 3140 2565
rect 3134 2560 3135 2564
rect 3139 2560 3140 2564
rect 3134 2559 3140 2560
rect 3262 2564 3268 2565
rect 3262 2560 3263 2564
rect 3267 2560 3268 2564
rect 3262 2559 3268 2560
rect 3390 2564 3396 2565
rect 3390 2560 3391 2564
rect 3395 2560 3396 2564
rect 3390 2559 3396 2560
rect 3502 2564 3508 2565
rect 3502 2560 3503 2564
rect 3507 2560 3508 2564
rect 3502 2559 3508 2560
rect 3590 2561 3596 2562
rect 1870 2556 1876 2557
rect 3590 2557 3591 2561
rect 3595 2557 3596 2561
rect 3590 2556 3596 2557
rect 150 2550 156 2551
rect 150 2546 151 2550
rect 155 2546 156 2550
rect 150 2545 156 2546
rect 318 2550 324 2551
rect 318 2546 319 2550
rect 323 2546 324 2550
rect 318 2545 324 2546
rect 486 2550 492 2551
rect 486 2546 487 2550
rect 491 2546 492 2550
rect 486 2545 492 2546
rect 646 2550 652 2551
rect 646 2546 647 2550
rect 651 2546 652 2550
rect 646 2545 652 2546
rect 798 2550 804 2551
rect 798 2546 799 2550
rect 803 2546 804 2550
rect 798 2545 804 2546
rect 934 2550 940 2551
rect 934 2546 935 2550
rect 939 2546 940 2550
rect 934 2545 940 2546
rect 1062 2550 1068 2551
rect 1062 2546 1063 2550
rect 1067 2546 1068 2550
rect 1062 2545 1068 2546
rect 1182 2550 1188 2551
rect 1182 2546 1183 2550
rect 1187 2546 1188 2550
rect 1182 2545 1188 2546
rect 1302 2550 1308 2551
rect 1302 2546 1303 2550
rect 1307 2546 1308 2550
rect 1302 2545 1308 2546
rect 1414 2550 1420 2551
rect 1414 2546 1415 2550
rect 1419 2546 1420 2550
rect 1414 2545 1420 2546
rect 1534 2550 1540 2551
rect 1534 2546 1535 2550
rect 1539 2546 1540 2550
rect 1534 2545 1540 2546
rect 1870 2544 1876 2545
rect 1870 2540 1871 2544
rect 1875 2540 1876 2544
rect 1870 2539 1876 2540
rect 3590 2544 3596 2545
rect 3590 2540 3591 2544
rect 3595 2540 3596 2544
rect 3590 2539 3596 2540
rect 2174 2526 2180 2527
rect 2174 2522 2175 2526
rect 2179 2522 2180 2526
rect 2174 2521 2180 2522
rect 2270 2526 2276 2527
rect 2270 2522 2271 2526
rect 2275 2522 2276 2526
rect 2270 2521 2276 2522
rect 2374 2526 2380 2527
rect 2374 2522 2375 2526
rect 2379 2522 2380 2526
rect 2374 2521 2380 2522
rect 2486 2526 2492 2527
rect 2486 2522 2487 2526
rect 2491 2522 2492 2526
rect 2486 2521 2492 2522
rect 2598 2526 2604 2527
rect 2598 2522 2599 2526
rect 2603 2522 2604 2526
rect 2598 2521 2604 2522
rect 2702 2526 2708 2527
rect 2702 2522 2703 2526
rect 2707 2522 2708 2526
rect 2702 2521 2708 2522
rect 2806 2526 2812 2527
rect 2806 2522 2807 2526
rect 2811 2522 2812 2526
rect 2806 2521 2812 2522
rect 2910 2526 2916 2527
rect 2910 2522 2911 2526
rect 2915 2522 2916 2526
rect 2910 2521 2916 2522
rect 3022 2526 3028 2527
rect 3022 2522 3023 2526
rect 3027 2522 3028 2526
rect 3022 2521 3028 2522
rect 3142 2526 3148 2527
rect 3142 2522 3143 2526
rect 3147 2522 3148 2526
rect 3142 2521 3148 2522
rect 3270 2526 3276 2527
rect 3270 2522 3271 2526
rect 3275 2522 3276 2526
rect 3270 2521 3276 2522
rect 3398 2526 3404 2527
rect 3398 2522 3399 2526
rect 3403 2522 3404 2526
rect 3398 2521 3404 2522
rect 3510 2526 3516 2527
rect 3510 2522 3511 2526
rect 3515 2522 3516 2526
rect 3510 2521 3516 2522
rect 142 2510 148 2511
rect 142 2506 143 2510
rect 147 2506 148 2510
rect 142 2505 148 2506
rect 294 2510 300 2511
rect 294 2506 295 2510
rect 299 2506 300 2510
rect 294 2505 300 2506
rect 446 2510 452 2511
rect 446 2506 447 2510
rect 451 2506 452 2510
rect 446 2505 452 2506
rect 590 2510 596 2511
rect 590 2506 591 2510
rect 595 2506 596 2510
rect 590 2505 596 2506
rect 734 2510 740 2511
rect 734 2506 735 2510
rect 739 2506 740 2510
rect 734 2505 740 2506
rect 878 2510 884 2511
rect 878 2506 879 2510
rect 883 2506 884 2510
rect 878 2505 884 2506
rect 1014 2510 1020 2511
rect 1014 2506 1015 2510
rect 1019 2506 1020 2510
rect 1014 2505 1020 2506
rect 1142 2510 1148 2511
rect 1142 2506 1143 2510
rect 1147 2506 1148 2510
rect 1142 2505 1148 2506
rect 1270 2510 1276 2511
rect 1270 2506 1271 2510
rect 1275 2506 1276 2510
rect 1270 2505 1276 2506
rect 1398 2510 1404 2511
rect 1398 2506 1399 2510
rect 1403 2506 1404 2510
rect 1398 2505 1404 2506
rect 1534 2510 1540 2511
rect 1534 2506 1535 2510
rect 1539 2506 1540 2510
rect 1534 2505 1540 2506
rect 2134 2494 2140 2495
rect 110 2492 116 2493
rect 110 2488 111 2492
rect 115 2488 116 2492
rect 110 2487 116 2488
rect 1830 2492 1836 2493
rect 1830 2488 1831 2492
rect 1835 2488 1836 2492
rect 2134 2490 2135 2494
rect 2139 2490 2140 2494
rect 2134 2489 2140 2490
rect 2222 2494 2228 2495
rect 2222 2490 2223 2494
rect 2227 2490 2228 2494
rect 2222 2489 2228 2490
rect 2318 2494 2324 2495
rect 2318 2490 2319 2494
rect 2323 2490 2324 2494
rect 2318 2489 2324 2490
rect 2422 2494 2428 2495
rect 2422 2490 2423 2494
rect 2427 2490 2428 2494
rect 2422 2489 2428 2490
rect 2534 2494 2540 2495
rect 2534 2490 2535 2494
rect 2539 2490 2540 2494
rect 2534 2489 2540 2490
rect 2654 2494 2660 2495
rect 2654 2490 2655 2494
rect 2659 2490 2660 2494
rect 2654 2489 2660 2490
rect 2782 2494 2788 2495
rect 2782 2490 2783 2494
rect 2787 2490 2788 2494
rect 2782 2489 2788 2490
rect 2918 2494 2924 2495
rect 2918 2490 2919 2494
rect 2923 2490 2924 2494
rect 2918 2489 2924 2490
rect 3062 2494 3068 2495
rect 3062 2490 3063 2494
rect 3067 2490 3068 2494
rect 3062 2489 3068 2490
rect 3214 2494 3220 2495
rect 3214 2490 3215 2494
rect 3219 2490 3220 2494
rect 3214 2489 3220 2490
rect 3374 2494 3380 2495
rect 3374 2490 3375 2494
rect 3379 2490 3380 2494
rect 3374 2489 3380 2490
rect 3510 2494 3516 2495
rect 3510 2490 3511 2494
rect 3515 2490 3516 2494
rect 3510 2489 3516 2490
rect 1830 2487 1836 2488
rect 1870 2476 1876 2477
rect 110 2475 116 2476
rect 110 2471 111 2475
rect 115 2471 116 2475
rect 1830 2475 1836 2476
rect 110 2470 116 2471
rect 134 2472 140 2473
rect 134 2468 135 2472
rect 139 2468 140 2472
rect 134 2467 140 2468
rect 286 2472 292 2473
rect 286 2468 287 2472
rect 291 2468 292 2472
rect 286 2467 292 2468
rect 438 2472 444 2473
rect 438 2468 439 2472
rect 443 2468 444 2472
rect 438 2467 444 2468
rect 582 2472 588 2473
rect 582 2468 583 2472
rect 587 2468 588 2472
rect 582 2467 588 2468
rect 726 2472 732 2473
rect 726 2468 727 2472
rect 731 2468 732 2472
rect 726 2467 732 2468
rect 870 2472 876 2473
rect 870 2468 871 2472
rect 875 2468 876 2472
rect 870 2467 876 2468
rect 1006 2472 1012 2473
rect 1006 2468 1007 2472
rect 1011 2468 1012 2472
rect 1006 2467 1012 2468
rect 1134 2472 1140 2473
rect 1134 2468 1135 2472
rect 1139 2468 1140 2472
rect 1134 2467 1140 2468
rect 1262 2472 1268 2473
rect 1262 2468 1263 2472
rect 1267 2468 1268 2472
rect 1262 2467 1268 2468
rect 1390 2472 1396 2473
rect 1390 2468 1391 2472
rect 1395 2468 1396 2472
rect 1390 2467 1396 2468
rect 1526 2472 1532 2473
rect 1526 2468 1527 2472
rect 1531 2468 1532 2472
rect 1830 2471 1831 2475
rect 1835 2471 1836 2475
rect 1870 2472 1871 2476
rect 1875 2472 1876 2476
rect 1870 2471 1876 2472
rect 3590 2476 3596 2477
rect 3590 2472 3591 2476
rect 3595 2472 3596 2476
rect 3590 2471 3596 2472
rect 1830 2470 1836 2471
rect 1526 2467 1532 2468
rect 1870 2459 1876 2460
rect 1870 2455 1871 2459
rect 1875 2455 1876 2459
rect 3590 2459 3596 2460
rect 1870 2454 1876 2455
rect 2126 2456 2132 2457
rect 2126 2452 2127 2456
rect 2131 2452 2132 2456
rect 2126 2451 2132 2452
rect 2214 2456 2220 2457
rect 2214 2452 2215 2456
rect 2219 2452 2220 2456
rect 2214 2451 2220 2452
rect 2310 2456 2316 2457
rect 2310 2452 2311 2456
rect 2315 2452 2316 2456
rect 2310 2451 2316 2452
rect 2414 2456 2420 2457
rect 2414 2452 2415 2456
rect 2419 2452 2420 2456
rect 2414 2451 2420 2452
rect 2526 2456 2532 2457
rect 2526 2452 2527 2456
rect 2531 2452 2532 2456
rect 2526 2451 2532 2452
rect 2646 2456 2652 2457
rect 2646 2452 2647 2456
rect 2651 2452 2652 2456
rect 2646 2451 2652 2452
rect 2774 2456 2780 2457
rect 2774 2452 2775 2456
rect 2779 2452 2780 2456
rect 2774 2451 2780 2452
rect 2910 2456 2916 2457
rect 2910 2452 2911 2456
rect 2915 2452 2916 2456
rect 2910 2451 2916 2452
rect 3054 2456 3060 2457
rect 3054 2452 3055 2456
rect 3059 2452 3060 2456
rect 3054 2451 3060 2452
rect 3206 2456 3212 2457
rect 3206 2452 3207 2456
rect 3211 2452 3212 2456
rect 3206 2451 3212 2452
rect 3366 2456 3372 2457
rect 3366 2452 3367 2456
rect 3371 2452 3372 2456
rect 3366 2451 3372 2452
rect 3502 2456 3508 2457
rect 3502 2452 3503 2456
rect 3507 2452 3508 2456
rect 3590 2455 3591 2459
rect 3595 2455 3596 2459
rect 3590 2454 3596 2455
rect 3502 2451 3508 2452
rect 198 2424 204 2425
rect 110 2421 116 2422
rect 110 2417 111 2421
rect 115 2417 116 2421
rect 198 2420 199 2424
rect 203 2420 204 2424
rect 198 2419 204 2420
rect 350 2424 356 2425
rect 350 2420 351 2424
rect 355 2420 356 2424
rect 350 2419 356 2420
rect 494 2424 500 2425
rect 494 2420 495 2424
rect 499 2420 500 2424
rect 494 2419 500 2420
rect 638 2424 644 2425
rect 638 2420 639 2424
rect 643 2420 644 2424
rect 638 2419 644 2420
rect 782 2424 788 2425
rect 782 2420 783 2424
rect 787 2420 788 2424
rect 782 2419 788 2420
rect 918 2424 924 2425
rect 918 2420 919 2424
rect 923 2420 924 2424
rect 918 2419 924 2420
rect 1046 2424 1052 2425
rect 1046 2420 1047 2424
rect 1051 2420 1052 2424
rect 1046 2419 1052 2420
rect 1174 2424 1180 2425
rect 1174 2420 1175 2424
rect 1179 2420 1180 2424
rect 1174 2419 1180 2420
rect 1310 2424 1316 2425
rect 1310 2420 1311 2424
rect 1315 2420 1316 2424
rect 1310 2419 1316 2420
rect 1446 2424 1452 2425
rect 1446 2420 1447 2424
rect 1451 2420 1452 2424
rect 1446 2419 1452 2420
rect 1830 2421 1836 2422
rect 110 2416 116 2417
rect 1830 2417 1831 2421
rect 1835 2417 1836 2421
rect 1830 2416 1836 2417
rect 110 2404 116 2405
rect 110 2400 111 2404
rect 115 2400 116 2404
rect 110 2399 116 2400
rect 1830 2404 1836 2405
rect 1830 2400 1831 2404
rect 1835 2400 1836 2404
rect 1974 2404 1980 2405
rect 1830 2399 1836 2400
rect 1870 2401 1876 2402
rect 1870 2397 1871 2401
rect 1875 2397 1876 2401
rect 1974 2400 1975 2404
rect 1979 2400 1980 2404
rect 1974 2399 1980 2400
rect 2086 2404 2092 2405
rect 2086 2400 2087 2404
rect 2091 2400 2092 2404
rect 2086 2399 2092 2400
rect 2206 2404 2212 2405
rect 2206 2400 2207 2404
rect 2211 2400 2212 2404
rect 2206 2399 2212 2400
rect 2334 2404 2340 2405
rect 2334 2400 2335 2404
rect 2339 2400 2340 2404
rect 2334 2399 2340 2400
rect 2478 2404 2484 2405
rect 2478 2400 2479 2404
rect 2483 2400 2484 2404
rect 2478 2399 2484 2400
rect 2630 2404 2636 2405
rect 2630 2400 2631 2404
rect 2635 2400 2636 2404
rect 2630 2399 2636 2400
rect 2790 2404 2796 2405
rect 2790 2400 2791 2404
rect 2795 2400 2796 2404
rect 2790 2399 2796 2400
rect 2966 2404 2972 2405
rect 2966 2400 2967 2404
rect 2971 2400 2972 2404
rect 2966 2399 2972 2400
rect 3150 2404 3156 2405
rect 3150 2400 3151 2404
rect 3155 2400 3156 2404
rect 3150 2399 3156 2400
rect 3334 2404 3340 2405
rect 3334 2400 3335 2404
rect 3339 2400 3340 2404
rect 3334 2399 3340 2400
rect 3502 2404 3508 2405
rect 3502 2400 3503 2404
rect 3507 2400 3508 2404
rect 3502 2399 3508 2400
rect 3590 2401 3596 2402
rect 1870 2396 1876 2397
rect 3590 2397 3591 2401
rect 3595 2397 3596 2401
rect 3590 2396 3596 2397
rect 206 2386 212 2387
rect 206 2382 207 2386
rect 211 2382 212 2386
rect 206 2381 212 2382
rect 358 2386 364 2387
rect 358 2382 359 2386
rect 363 2382 364 2386
rect 358 2381 364 2382
rect 502 2386 508 2387
rect 502 2382 503 2386
rect 507 2382 508 2386
rect 502 2381 508 2382
rect 646 2386 652 2387
rect 646 2382 647 2386
rect 651 2382 652 2386
rect 646 2381 652 2382
rect 790 2386 796 2387
rect 790 2382 791 2386
rect 795 2382 796 2386
rect 790 2381 796 2382
rect 926 2386 932 2387
rect 926 2382 927 2386
rect 931 2382 932 2386
rect 926 2381 932 2382
rect 1054 2386 1060 2387
rect 1054 2382 1055 2386
rect 1059 2382 1060 2386
rect 1054 2381 1060 2382
rect 1182 2386 1188 2387
rect 1182 2382 1183 2386
rect 1187 2382 1188 2386
rect 1182 2381 1188 2382
rect 1318 2386 1324 2387
rect 1318 2382 1319 2386
rect 1323 2382 1324 2386
rect 1318 2381 1324 2382
rect 1454 2386 1460 2387
rect 1454 2382 1455 2386
rect 1459 2382 1460 2386
rect 1454 2381 1460 2382
rect 1870 2384 1876 2385
rect 1870 2380 1871 2384
rect 1875 2380 1876 2384
rect 1870 2379 1876 2380
rect 3590 2384 3596 2385
rect 3590 2380 3591 2384
rect 3595 2380 3596 2384
rect 3590 2379 3596 2380
rect 1982 2366 1988 2367
rect 1982 2362 1983 2366
rect 1987 2362 1988 2366
rect 1982 2361 1988 2362
rect 2094 2366 2100 2367
rect 2094 2362 2095 2366
rect 2099 2362 2100 2366
rect 2094 2361 2100 2362
rect 2214 2366 2220 2367
rect 2214 2362 2215 2366
rect 2219 2362 2220 2366
rect 2214 2361 2220 2362
rect 2342 2366 2348 2367
rect 2342 2362 2343 2366
rect 2347 2362 2348 2366
rect 2342 2361 2348 2362
rect 2486 2366 2492 2367
rect 2486 2362 2487 2366
rect 2491 2362 2492 2366
rect 2486 2361 2492 2362
rect 2638 2366 2644 2367
rect 2638 2362 2639 2366
rect 2643 2362 2644 2366
rect 2638 2361 2644 2362
rect 2798 2366 2804 2367
rect 2798 2362 2799 2366
rect 2803 2362 2804 2366
rect 2798 2361 2804 2362
rect 2974 2366 2980 2367
rect 2974 2362 2975 2366
rect 2979 2362 2980 2366
rect 2974 2361 2980 2362
rect 3158 2366 3164 2367
rect 3158 2362 3159 2366
rect 3163 2362 3164 2366
rect 3158 2361 3164 2362
rect 3342 2366 3348 2367
rect 3342 2362 3343 2366
rect 3347 2362 3348 2366
rect 3342 2361 3348 2362
rect 3510 2366 3516 2367
rect 3510 2362 3511 2366
rect 3515 2362 3516 2366
rect 3510 2361 3516 2362
rect 222 2346 228 2347
rect 222 2342 223 2346
rect 227 2342 228 2346
rect 222 2341 228 2342
rect 326 2346 332 2347
rect 326 2342 327 2346
rect 331 2342 332 2346
rect 326 2341 332 2342
rect 438 2346 444 2347
rect 438 2342 439 2346
rect 443 2342 444 2346
rect 438 2341 444 2342
rect 558 2346 564 2347
rect 558 2342 559 2346
rect 563 2342 564 2346
rect 558 2341 564 2342
rect 678 2346 684 2347
rect 678 2342 679 2346
rect 683 2342 684 2346
rect 678 2341 684 2342
rect 798 2346 804 2347
rect 798 2342 799 2346
rect 803 2342 804 2346
rect 798 2341 804 2342
rect 910 2346 916 2347
rect 910 2342 911 2346
rect 915 2342 916 2346
rect 910 2341 916 2342
rect 1022 2346 1028 2347
rect 1022 2342 1023 2346
rect 1027 2342 1028 2346
rect 1022 2341 1028 2342
rect 1134 2346 1140 2347
rect 1134 2342 1135 2346
rect 1139 2342 1140 2346
rect 1134 2341 1140 2342
rect 1246 2346 1252 2347
rect 1246 2342 1247 2346
rect 1251 2342 1252 2346
rect 1246 2341 1252 2342
rect 1366 2346 1372 2347
rect 1366 2342 1367 2346
rect 1371 2342 1372 2346
rect 1366 2341 1372 2342
rect 1902 2330 1908 2331
rect 110 2328 116 2329
rect 110 2324 111 2328
rect 115 2324 116 2328
rect 110 2323 116 2324
rect 1830 2328 1836 2329
rect 1830 2324 1831 2328
rect 1835 2324 1836 2328
rect 1902 2326 1903 2330
rect 1907 2326 1908 2330
rect 1902 2325 1908 2326
rect 2014 2330 2020 2331
rect 2014 2326 2015 2330
rect 2019 2326 2020 2330
rect 2014 2325 2020 2326
rect 2166 2330 2172 2331
rect 2166 2326 2167 2330
rect 2171 2326 2172 2330
rect 2166 2325 2172 2326
rect 2318 2330 2324 2331
rect 2318 2326 2319 2330
rect 2323 2326 2324 2330
rect 2318 2325 2324 2326
rect 2470 2330 2476 2331
rect 2470 2326 2471 2330
rect 2475 2326 2476 2330
rect 2470 2325 2476 2326
rect 2622 2330 2628 2331
rect 2622 2326 2623 2330
rect 2627 2326 2628 2330
rect 2622 2325 2628 2326
rect 2774 2330 2780 2331
rect 2774 2326 2775 2330
rect 2779 2326 2780 2330
rect 2774 2325 2780 2326
rect 2926 2330 2932 2331
rect 2926 2326 2927 2330
rect 2931 2326 2932 2330
rect 2926 2325 2932 2326
rect 3086 2330 3092 2331
rect 3086 2326 3087 2330
rect 3091 2326 3092 2330
rect 3086 2325 3092 2326
rect 3246 2330 3252 2331
rect 3246 2326 3247 2330
rect 3251 2326 3252 2330
rect 3246 2325 3252 2326
rect 3414 2330 3420 2331
rect 3414 2326 3415 2330
rect 3419 2326 3420 2330
rect 3414 2325 3420 2326
rect 1830 2323 1836 2324
rect 1870 2312 1876 2313
rect 110 2311 116 2312
rect 110 2307 111 2311
rect 115 2307 116 2311
rect 1830 2311 1836 2312
rect 110 2306 116 2307
rect 214 2308 220 2309
rect 214 2304 215 2308
rect 219 2304 220 2308
rect 214 2303 220 2304
rect 318 2308 324 2309
rect 318 2304 319 2308
rect 323 2304 324 2308
rect 318 2303 324 2304
rect 430 2308 436 2309
rect 430 2304 431 2308
rect 435 2304 436 2308
rect 430 2303 436 2304
rect 550 2308 556 2309
rect 550 2304 551 2308
rect 555 2304 556 2308
rect 550 2303 556 2304
rect 670 2308 676 2309
rect 670 2304 671 2308
rect 675 2304 676 2308
rect 670 2303 676 2304
rect 790 2308 796 2309
rect 790 2304 791 2308
rect 795 2304 796 2308
rect 790 2303 796 2304
rect 902 2308 908 2309
rect 902 2304 903 2308
rect 907 2304 908 2308
rect 902 2303 908 2304
rect 1014 2308 1020 2309
rect 1014 2304 1015 2308
rect 1019 2304 1020 2308
rect 1014 2303 1020 2304
rect 1126 2308 1132 2309
rect 1126 2304 1127 2308
rect 1131 2304 1132 2308
rect 1126 2303 1132 2304
rect 1238 2308 1244 2309
rect 1238 2304 1239 2308
rect 1243 2304 1244 2308
rect 1238 2303 1244 2304
rect 1358 2308 1364 2309
rect 1358 2304 1359 2308
rect 1363 2304 1364 2308
rect 1830 2307 1831 2311
rect 1835 2307 1836 2311
rect 1870 2308 1871 2312
rect 1875 2308 1876 2312
rect 1870 2307 1876 2308
rect 3590 2312 3596 2313
rect 3590 2308 3591 2312
rect 3595 2308 3596 2312
rect 3590 2307 3596 2308
rect 1830 2306 1836 2307
rect 1358 2303 1364 2304
rect 1870 2295 1876 2296
rect 1870 2291 1871 2295
rect 1875 2291 1876 2295
rect 3590 2295 3596 2296
rect 1870 2290 1876 2291
rect 1894 2292 1900 2293
rect 1894 2288 1895 2292
rect 1899 2288 1900 2292
rect 1894 2287 1900 2288
rect 2006 2292 2012 2293
rect 2006 2288 2007 2292
rect 2011 2288 2012 2292
rect 2006 2287 2012 2288
rect 2158 2292 2164 2293
rect 2158 2288 2159 2292
rect 2163 2288 2164 2292
rect 2158 2287 2164 2288
rect 2310 2292 2316 2293
rect 2310 2288 2311 2292
rect 2315 2288 2316 2292
rect 2310 2287 2316 2288
rect 2462 2292 2468 2293
rect 2462 2288 2463 2292
rect 2467 2288 2468 2292
rect 2462 2287 2468 2288
rect 2614 2292 2620 2293
rect 2614 2288 2615 2292
rect 2619 2288 2620 2292
rect 2614 2287 2620 2288
rect 2766 2292 2772 2293
rect 2766 2288 2767 2292
rect 2771 2288 2772 2292
rect 2766 2287 2772 2288
rect 2918 2292 2924 2293
rect 2918 2288 2919 2292
rect 2923 2288 2924 2292
rect 2918 2287 2924 2288
rect 3078 2292 3084 2293
rect 3078 2288 3079 2292
rect 3083 2288 3084 2292
rect 3078 2287 3084 2288
rect 3238 2292 3244 2293
rect 3238 2288 3239 2292
rect 3243 2288 3244 2292
rect 3238 2287 3244 2288
rect 3406 2292 3412 2293
rect 3406 2288 3407 2292
rect 3411 2288 3412 2292
rect 3590 2291 3591 2295
rect 3595 2291 3596 2295
rect 3590 2290 3596 2291
rect 3406 2287 3412 2288
rect 310 2252 316 2253
rect 110 2249 116 2250
rect 110 2245 111 2249
rect 115 2245 116 2249
rect 310 2248 311 2252
rect 315 2248 316 2252
rect 310 2247 316 2248
rect 406 2252 412 2253
rect 406 2248 407 2252
rect 411 2248 412 2252
rect 406 2247 412 2248
rect 502 2252 508 2253
rect 502 2248 503 2252
rect 507 2248 508 2252
rect 502 2247 508 2248
rect 606 2252 612 2253
rect 606 2248 607 2252
rect 611 2248 612 2252
rect 606 2247 612 2248
rect 710 2252 716 2253
rect 710 2248 711 2252
rect 715 2248 716 2252
rect 710 2247 716 2248
rect 814 2252 820 2253
rect 814 2248 815 2252
rect 819 2248 820 2252
rect 814 2247 820 2248
rect 910 2252 916 2253
rect 910 2248 911 2252
rect 915 2248 916 2252
rect 910 2247 916 2248
rect 1006 2252 1012 2253
rect 1006 2248 1007 2252
rect 1011 2248 1012 2252
rect 1006 2247 1012 2248
rect 1102 2252 1108 2253
rect 1102 2248 1103 2252
rect 1107 2248 1108 2252
rect 1102 2247 1108 2248
rect 1198 2252 1204 2253
rect 1198 2248 1199 2252
rect 1203 2248 1204 2252
rect 1198 2247 1204 2248
rect 1302 2252 1308 2253
rect 1302 2248 1303 2252
rect 1307 2248 1308 2252
rect 1302 2247 1308 2248
rect 1830 2249 1836 2250
rect 110 2244 116 2245
rect 1830 2245 1831 2249
rect 1835 2245 1836 2249
rect 1894 2248 1900 2249
rect 1830 2244 1836 2245
rect 1870 2245 1876 2246
rect 1870 2241 1871 2245
rect 1875 2241 1876 2245
rect 1894 2244 1895 2248
rect 1899 2244 1900 2248
rect 1894 2243 1900 2244
rect 2030 2248 2036 2249
rect 2030 2244 2031 2248
rect 2035 2244 2036 2248
rect 2030 2243 2036 2244
rect 2206 2248 2212 2249
rect 2206 2244 2207 2248
rect 2211 2244 2212 2248
rect 2206 2243 2212 2244
rect 2390 2248 2396 2249
rect 2390 2244 2391 2248
rect 2395 2244 2396 2248
rect 2390 2243 2396 2244
rect 2574 2248 2580 2249
rect 2574 2244 2575 2248
rect 2579 2244 2580 2248
rect 2574 2243 2580 2244
rect 2766 2248 2772 2249
rect 2766 2244 2767 2248
rect 2771 2244 2772 2248
rect 2766 2243 2772 2244
rect 2950 2248 2956 2249
rect 2950 2244 2951 2248
rect 2955 2244 2956 2248
rect 2950 2243 2956 2244
rect 3142 2248 3148 2249
rect 3142 2244 3143 2248
rect 3147 2244 3148 2248
rect 3142 2243 3148 2244
rect 3334 2248 3340 2249
rect 3334 2244 3335 2248
rect 3339 2244 3340 2248
rect 3334 2243 3340 2244
rect 3502 2248 3508 2249
rect 3502 2244 3503 2248
rect 3507 2244 3508 2248
rect 3502 2243 3508 2244
rect 3590 2245 3596 2246
rect 1870 2240 1876 2241
rect 3590 2241 3591 2245
rect 3595 2241 3596 2245
rect 3590 2240 3596 2241
rect 110 2232 116 2233
rect 110 2228 111 2232
rect 115 2228 116 2232
rect 110 2227 116 2228
rect 1830 2232 1836 2233
rect 1830 2228 1831 2232
rect 1835 2228 1836 2232
rect 1830 2227 1836 2228
rect 1870 2228 1876 2229
rect 1870 2224 1871 2228
rect 1875 2224 1876 2228
rect 1870 2223 1876 2224
rect 3590 2228 3596 2229
rect 3590 2224 3591 2228
rect 3595 2224 3596 2228
rect 3590 2223 3596 2224
rect 318 2214 324 2215
rect 318 2210 319 2214
rect 323 2210 324 2214
rect 318 2209 324 2210
rect 414 2214 420 2215
rect 414 2210 415 2214
rect 419 2210 420 2214
rect 414 2209 420 2210
rect 510 2214 516 2215
rect 510 2210 511 2214
rect 515 2210 516 2214
rect 510 2209 516 2210
rect 614 2214 620 2215
rect 614 2210 615 2214
rect 619 2210 620 2214
rect 614 2209 620 2210
rect 718 2214 724 2215
rect 718 2210 719 2214
rect 723 2210 724 2214
rect 718 2209 724 2210
rect 822 2214 828 2215
rect 822 2210 823 2214
rect 827 2210 828 2214
rect 822 2209 828 2210
rect 918 2214 924 2215
rect 918 2210 919 2214
rect 923 2210 924 2214
rect 918 2209 924 2210
rect 1014 2214 1020 2215
rect 1014 2210 1015 2214
rect 1019 2210 1020 2214
rect 1014 2209 1020 2210
rect 1110 2214 1116 2215
rect 1110 2210 1111 2214
rect 1115 2210 1116 2214
rect 1110 2209 1116 2210
rect 1206 2214 1212 2215
rect 1206 2210 1207 2214
rect 1211 2210 1212 2214
rect 1206 2209 1212 2210
rect 1310 2214 1316 2215
rect 1310 2210 1311 2214
rect 1315 2210 1316 2214
rect 1310 2209 1316 2210
rect 1902 2210 1908 2211
rect 1902 2206 1903 2210
rect 1907 2206 1908 2210
rect 1902 2205 1908 2206
rect 2038 2210 2044 2211
rect 2038 2206 2039 2210
rect 2043 2206 2044 2210
rect 2038 2205 2044 2206
rect 2214 2210 2220 2211
rect 2214 2206 2215 2210
rect 2219 2206 2220 2210
rect 2214 2205 2220 2206
rect 2398 2210 2404 2211
rect 2398 2206 2399 2210
rect 2403 2206 2404 2210
rect 2398 2205 2404 2206
rect 2582 2210 2588 2211
rect 2582 2206 2583 2210
rect 2587 2206 2588 2210
rect 2582 2205 2588 2206
rect 2774 2210 2780 2211
rect 2774 2206 2775 2210
rect 2779 2206 2780 2210
rect 2774 2205 2780 2206
rect 2958 2210 2964 2211
rect 2958 2206 2959 2210
rect 2963 2206 2964 2210
rect 2958 2205 2964 2206
rect 3150 2210 3156 2211
rect 3150 2206 3151 2210
rect 3155 2206 3156 2210
rect 3150 2205 3156 2206
rect 3342 2210 3348 2211
rect 3342 2206 3343 2210
rect 3347 2206 3348 2210
rect 3342 2205 3348 2206
rect 3510 2210 3516 2211
rect 3510 2206 3511 2210
rect 3515 2206 3516 2210
rect 3510 2205 3516 2206
rect 318 2178 324 2179
rect 318 2174 319 2178
rect 323 2174 324 2178
rect 318 2173 324 2174
rect 414 2178 420 2179
rect 414 2174 415 2178
rect 419 2174 420 2178
rect 414 2173 420 2174
rect 518 2178 524 2179
rect 518 2174 519 2178
rect 523 2174 524 2178
rect 518 2173 524 2174
rect 622 2178 628 2179
rect 622 2174 623 2178
rect 627 2174 628 2178
rect 622 2173 628 2174
rect 726 2178 732 2179
rect 726 2174 727 2178
rect 731 2174 732 2178
rect 726 2173 732 2174
rect 830 2178 836 2179
rect 830 2174 831 2178
rect 835 2174 836 2178
rect 830 2173 836 2174
rect 934 2178 940 2179
rect 934 2174 935 2178
rect 939 2174 940 2178
rect 934 2173 940 2174
rect 1038 2178 1044 2179
rect 1038 2174 1039 2178
rect 1043 2174 1044 2178
rect 1038 2173 1044 2174
rect 1150 2178 1156 2179
rect 1150 2174 1151 2178
rect 1155 2174 1156 2178
rect 1150 2173 1156 2174
rect 1262 2178 1268 2179
rect 1262 2174 1263 2178
rect 1267 2174 1268 2178
rect 1262 2173 1268 2174
rect 1966 2170 1972 2171
rect 1966 2166 1967 2170
rect 1971 2166 1972 2170
rect 1966 2165 1972 2166
rect 2078 2170 2084 2171
rect 2078 2166 2079 2170
rect 2083 2166 2084 2170
rect 2078 2165 2084 2166
rect 2214 2170 2220 2171
rect 2214 2166 2215 2170
rect 2219 2166 2220 2170
rect 2214 2165 2220 2166
rect 2366 2170 2372 2171
rect 2366 2166 2367 2170
rect 2371 2166 2372 2170
rect 2366 2165 2372 2166
rect 2526 2170 2532 2171
rect 2526 2166 2527 2170
rect 2531 2166 2532 2170
rect 2526 2165 2532 2166
rect 2686 2170 2692 2171
rect 2686 2166 2687 2170
rect 2691 2166 2692 2170
rect 2686 2165 2692 2166
rect 2846 2170 2852 2171
rect 2846 2166 2847 2170
rect 2851 2166 2852 2170
rect 2846 2165 2852 2166
rect 2990 2170 2996 2171
rect 2990 2166 2991 2170
rect 2995 2166 2996 2170
rect 2990 2165 2996 2166
rect 3126 2170 3132 2171
rect 3126 2166 3127 2170
rect 3131 2166 3132 2170
rect 3126 2165 3132 2166
rect 3262 2170 3268 2171
rect 3262 2166 3263 2170
rect 3267 2166 3268 2170
rect 3262 2165 3268 2166
rect 3398 2170 3404 2171
rect 3398 2166 3399 2170
rect 3403 2166 3404 2170
rect 3398 2165 3404 2166
rect 3510 2170 3516 2171
rect 3510 2166 3511 2170
rect 3515 2166 3516 2170
rect 3510 2165 3516 2166
rect 110 2160 116 2161
rect 110 2156 111 2160
rect 115 2156 116 2160
rect 110 2155 116 2156
rect 1830 2160 1836 2161
rect 1830 2156 1831 2160
rect 1835 2156 1836 2160
rect 1830 2155 1836 2156
rect 1870 2152 1876 2153
rect 1870 2148 1871 2152
rect 1875 2148 1876 2152
rect 1870 2147 1876 2148
rect 3590 2152 3596 2153
rect 3590 2148 3591 2152
rect 3595 2148 3596 2152
rect 3590 2147 3596 2148
rect 110 2143 116 2144
rect 110 2139 111 2143
rect 115 2139 116 2143
rect 1830 2143 1836 2144
rect 110 2138 116 2139
rect 310 2140 316 2141
rect 310 2136 311 2140
rect 315 2136 316 2140
rect 310 2135 316 2136
rect 406 2140 412 2141
rect 406 2136 407 2140
rect 411 2136 412 2140
rect 406 2135 412 2136
rect 510 2140 516 2141
rect 510 2136 511 2140
rect 515 2136 516 2140
rect 510 2135 516 2136
rect 614 2140 620 2141
rect 614 2136 615 2140
rect 619 2136 620 2140
rect 614 2135 620 2136
rect 718 2140 724 2141
rect 718 2136 719 2140
rect 723 2136 724 2140
rect 718 2135 724 2136
rect 822 2140 828 2141
rect 822 2136 823 2140
rect 827 2136 828 2140
rect 822 2135 828 2136
rect 926 2140 932 2141
rect 926 2136 927 2140
rect 931 2136 932 2140
rect 926 2135 932 2136
rect 1030 2140 1036 2141
rect 1030 2136 1031 2140
rect 1035 2136 1036 2140
rect 1030 2135 1036 2136
rect 1142 2140 1148 2141
rect 1142 2136 1143 2140
rect 1147 2136 1148 2140
rect 1142 2135 1148 2136
rect 1254 2140 1260 2141
rect 1254 2136 1255 2140
rect 1259 2136 1260 2140
rect 1830 2139 1831 2143
rect 1835 2139 1836 2143
rect 1830 2138 1836 2139
rect 1254 2135 1260 2136
rect 1870 2135 1876 2136
rect 1870 2131 1871 2135
rect 1875 2131 1876 2135
rect 3590 2135 3596 2136
rect 1870 2130 1876 2131
rect 1958 2132 1964 2133
rect 1958 2128 1959 2132
rect 1963 2128 1964 2132
rect 1958 2127 1964 2128
rect 2070 2132 2076 2133
rect 2070 2128 2071 2132
rect 2075 2128 2076 2132
rect 2070 2127 2076 2128
rect 2206 2132 2212 2133
rect 2206 2128 2207 2132
rect 2211 2128 2212 2132
rect 2206 2127 2212 2128
rect 2358 2132 2364 2133
rect 2358 2128 2359 2132
rect 2363 2128 2364 2132
rect 2358 2127 2364 2128
rect 2518 2132 2524 2133
rect 2518 2128 2519 2132
rect 2523 2128 2524 2132
rect 2518 2127 2524 2128
rect 2678 2132 2684 2133
rect 2678 2128 2679 2132
rect 2683 2128 2684 2132
rect 2678 2127 2684 2128
rect 2838 2132 2844 2133
rect 2838 2128 2839 2132
rect 2843 2128 2844 2132
rect 2838 2127 2844 2128
rect 2982 2132 2988 2133
rect 2982 2128 2983 2132
rect 2987 2128 2988 2132
rect 2982 2127 2988 2128
rect 3118 2132 3124 2133
rect 3118 2128 3119 2132
rect 3123 2128 3124 2132
rect 3118 2127 3124 2128
rect 3254 2132 3260 2133
rect 3254 2128 3255 2132
rect 3259 2128 3260 2132
rect 3254 2127 3260 2128
rect 3390 2132 3396 2133
rect 3390 2128 3391 2132
rect 3395 2128 3396 2132
rect 3390 2127 3396 2128
rect 3502 2132 3508 2133
rect 3502 2128 3503 2132
rect 3507 2128 3508 2132
rect 3590 2131 3591 2135
rect 3595 2131 3596 2135
rect 3590 2130 3596 2131
rect 3502 2127 3508 2128
rect 278 2096 284 2097
rect 110 2093 116 2094
rect 110 2089 111 2093
rect 115 2089 116 2093
rect 278 2092 279 2096
rect 283 2092 284 2096
rect 278 2091 284 2092
rect 398 2096 404 2097
rect 398 2092 399 2096
rect 403 2092 404 2096
rect 398 2091 404 2092
rect 510 2096 516 2097
rect 510 2092 511 2096
rect 515 2092 516 2096
rect 510 2091 516 2092
rect 622 2096 628 2097
rect 622 2092 623 2096
rect 627 2092 628 2096
rect 622 2091 628 2092
rect 734 2096 740 2097
rect 734 2092 735 2096
rect 739 2092 740 2096
rect 734 2091 740 2092
rect 846 2096 852 2097
rect 846 2092 847 2096
rect 851 2092 852 2096
rect 846 2091 852 2092
rect 950 2096 956 2097
rect 950 2092 951 2096
rect 955 2092 956 2096
rect 950 2091 956 2092
rect 1046 2096 1052 2097
rect 1046 2092 1047 2096
rect 1051 2092 1052 2096
rect 1046 2091 1052 2092
rect 1142 2096 1148 2097
rect 1142 2092 1143 2096
rect 1147 2092 1148 2096
rect 1142 2091 1148 2092
rect 1238 2096 1244 2097
rect 1238 2092 1239 2096
rect 1243 2092 1244 2096
rect 1238 2091 1244 2092
rect 1342 2096 1348 2097
rect 1342 2092 1343 2096
rect 1347 2092 1348 2096
rect 1342 2091 1348 2092
rect 1830 2093 1836 2094
rect 110 2088 116 2089
rect 1830 2089 1831 2093
rect 1835 2089 1836 2093
rect 1830 2088 1836 2089
rect 2286 2088 2292 2089
rect 1870 2085 1876 2086
rect 1870 2081 1871 2085
rect 1875 2081 1876 2085
rect 2286 2084 2287 2088
rect 2291 2084 2292 2088
rect 2286 2083 2292 2084
rect 2390 2088 2396 2089
rect 2390 2084 2391 2088
rect 2395 2084 2396 2088
rect 2390 2083 2396 2084
rect 2502 2088 2508 2089
rect 2502 2084 2503 2088
rect 2507 2084 2508 2088
rect 2502 2083 2508 2084
rect 2622 2088 2628 2089
rect 2622 2084 2623 2088
rect 2627 2084 2628 2088
rect 2622 2083 2628 2084
rect 2742 2088 2748 2089
rect 2742 2084 2743 2088
rect 2747 2084 2748 2088
rect 2742 2083 2748 2084
rect 2854 2088 2860 2089
rect 2854 2084 2855 2088
rect 2859 2084 2860 2088
rect 2854 2083 2860 2084
rect 2966 2088 2972 2089
rect 2966 2084 2967 2088
rect 2971 2084 2972 2088
rect 2966 2083 2972 2084
rect 3078 2088 3084 2089
rect 3078 2084 3079 2088
rect 3083 2084 3084 2088
rect 3078 2083 3084 2084
rect 3190 2088 3196 2089
rect 3190 2084 3191 2088
rect 3195 2084 3196 2088
rect 3190 2083 3196 2084
rect 3302 2088 3308 2089
rect 3302 2084 3303 2088
rect 3307 2084 3308 2088
rect 3302 2083 3308 2084
rect 3414 2088 3420 2089
rect 3414 2084 3415 2088
rect 3419 2084 3420 2088
rect 3414 2083 3420 2084
rect 3502 2088 3508 2089
rect 3502 2084 3503 2088
rect 3507 2084 3508 2088
rect 3502 2083 3508 2084
rect 3590 2085 3596 2086
rect 1870 2080 1876 2081
rect 3590 2081 3591 2085
rect 3595 2081 3596 2085
rect 3590 2080 3596 2081
rect 110 2076 116 2077
rect 110 2072 111 2076
rect 115 2072 116 2076
rect 110 2071 116 2072
rect 1830 2076 1836 2077
rect 1830 2072 1831 2076
rect 1835 2072 1836 2076
rect 1830 2071 1836 2072
rect 1870 2068 1876 2069
rect 1870 2064 1871 2068
rect 1875 2064 1876 2068
rect 1870 2063 1876 2064
rect 3590 2068 3596 2069
rect 3590 2064 3591 2068
rect 3595 2064 3596 2068
rect 3590 2063 3596 2064
rect 286 2058 292 2059
rect 286 2054 287 2058
rect 291 2054 292 2058
rect 286 2053 292 2054
rect 406 2058 412 2059
rect 406 2054 407 2058
rect 411 2054 412 2058
rect 406 2053 412 2054
rect 518 2058 524 2059
rect 518 2054 519 2058
rect 523 2054 524 2058
rect 518 2053 524 2054
rect 630 2058 636 2059
rect 630 2054 631 2058
rect 635 2054 636 2058
rect 630 2053 636 2054
rect 742 2058 748 2059
rect 742 2054 743 2058
rect 747 2054 748 2058
rect 742 2053 748 2054
rect 854 2058 860 2059
rect 854 2054 855 2058
rect 859 2054 860 2058
rect 854 2053 860 2054
rect 958 2058 964 2059
rect 958 2054 959 2058
rect 963 2054 964 2058
rect 958 2053 964 2054
rect 1054 2058 1060 2059
rect 1054 2054 1055 2058
rect 1059 2054 1060 2058
rect 1054 2053 1060 2054
rect 1150 2058 1156 2059
rect 1150 2054 1151 2058
rect 1155 2054 1156 2058
rect 1150 2053 1156 2054
rect 1246 2058 1252 2059
rect 1246 2054 1247 2058
rect 1251 2054 1252 2058
rect 1246 2053 1252 2054
rect 1350 2058 1356 2059
rect 1350 2054 1351 2058
rect 1355 2054 1356 2058
rect 1350 2053 1356 2054
rect 2294 2050 2300 2051
rect 2294 2046 2295 2050
rect 2299 2046 2300 2050
rect 2294 2045 2300 2046
rect 2398 2050 2404 2051
rect 2398 2046 2399 2050
rect 2403 2046 2404 2050
rect 2398 2045 2404 2046
rect 2510 2050 2516 2051
rect 2510 2046 2511 2050
rect 2515 2046 2516 2050
rect 2510 2045 2516 2046
rect 2630 2050 2636 2051
rect 2630 2046 2631 2050
rect 2635 2046 2636 2050
rect 2630 2045 2636 2046
rect 2750 2050 2756 2051
rect 2750 2046 2751 2050
rect 2755 2046 2756 2050
rect 2750 2045 2756 2046
rect 2862 2050 2868 2051
rect 2862 2046 2863 2050
rect 2867 2046 2868 2050
rect 2862 2045 2868 2046
rect 2974 2050 2980 2051
rect 2974 2046 2975 2050
rect 2979 2046 2980 2050
rect 2974 2045 2980 2046
rect 3086 2050 3092 2051
rect 3086 2046 3087 2050
rect 3091 2046 3092 2050
rect 3086 2045 3092 2046
rect 3198 2050 3204 2051
rect 3198 2046 3199 2050
rect 3203 2046 3204 2050
rect 3198 2045 3204 2046
rect 3310 2050 3316 2051
rect 3310 2046 3311 2050
rect 3315 2046 3316 2050
rect 3310 2045 3316 2046
rect 3422 2050 3428 2051
rect 3422 2046 3423 2050
rect 3427 2046 3428 2050
rect 3422 2045 3428 2046
rect 3510 2050 3516 2051
rect 3510 2046 3511 2050
rect 3515 2046 3516 2050
rect 3510 2045 3516 2046
rect 182 2018 188 2019
rect 182 2014 183 2018
rect 187 2014 188 2018
rect 182 2013 188 2014
rect 326 2018 332 2019
rect 326 2014 327 2018
rect 331 2014 332 2018
rect 326 2013 332 2014
rect 470 2018 476 2019
rect 470 2014 471 2018
rect 475 2014 476 2018
rect 470 2013 476 2014
rect 622 2018 628 2019
rect 622 2014 623 2018
rect 627 2014 628 2018
rect 622 2013 628 2014
rect 766 2018 772 2019
rect 766 2014 767 2018
rect 771 2014 772 2018
rect 766 2013 772 2014
rect 910 2018 916 2019
rect 910 2014 911 2018
rect 915 2014 916 2018
rect 910 2013 916 2014
rect 1046 2018 1052 2019
rect 1046 2014 1047 2018
rect 1051 2014 1052 2018
rect 1046 2013 1052 2014
rect 1182 2018 1188 2019
rect 1182 2014 1183 2018
rect 1187 2014 1188 2018
rect 1182 2013 1188 2014
rect 1318 2018 1324 2019
rect 1318 2014 1319 2018
rect 1323 2014 1324 2018
rect 1318 2013 1324 2014
rect 1462 2018 1468 2019
rect 1462 2014 1463 2018
rect 1467 2014 1468 2018
rect 1462 2013 1468 2014
rect 2182 2014 2188 2015
rect 2182 2010 2183 2014
rect 2187 2010 2188 2014
rect 2182 2009 2188 2010
rect 2270 2014 2276 2015
rect 2270 2010 2271 2014
rect 2275 2010 2276 2014
rect 2270 2009 2276 2010
rect 2366 2014 2372 2015
rect 2366 2010 2367 2014
rect 2371 2010 2372 2014
rect 2366 2009 2372 2010
rect 2462 2014 2468 2015
rect 2462 2010 2463 2014
rect 2467 2010 2468 2014
rect 2462 2009 2468 2010
rect 2566 2014 2572 2015
rect 2566 2010 2567 2014
rect 2571 2010 2572 2014
rect 2566 2009 2572 2010
rect 2670 2014 2676 2015
rect 2670 2010 2671 2014
rect 2675 2010 2676 2014
rect 2670 2009 2676 2010
rect 2774 2014 2780 2015
rect 2774 2010 2775 2014
rect 2779 2010 2780 2014
rect 2774 2009 2780 2010
rect 2878 2014 2884 2015
rect 2878 2010 2879 2014
rect 2883 2010 2884 2014
rect 2878 2009 2884 2010
rect 2982 2014 2988 2015
rect 2982 2010 2983 2014
rect 2987 2010 2988 2014
rect 2982 2009 2988 2010
rect 3086 2014 3092 2015
rect 3086 2010 3087 2014
rect 3091 2010 3092 2014
rect 3086 2009 3092 2010
rect 3190 2014 3196 2015
rect 3190 2010 3191 2014
rect 3195 2010 3196 2014
rect 3190 2009 3196 2010
rect 110 2000 116 2001
rect 110 1996 111 2000
rect 115 1996 116 2000
rect 110 1995 116 1996
rect 1830 2000 1836 2001
rect 1830 1996 1831 2000
rect 1835 1996 1836 2000
rect 1830 1995 1836 1996
rect 1870 1996 1876 1997
rect 1870 1992 1871 1996
rect 1875 1992 1876 1996
rect 1870 1991 1876 1992
rect 3590 1996 3596 1997
rect 3590 1992 3591 1996
rect 3595 1992 3596 1996
rect 3590 1991 3596 1992
rect 110 1983 116 1984
rect 110 1979 111 1983
rect 115 1979 116 1983
rect 1830 1983 1836 1984
rect 110 1978 116 1979
rect 174 1980 180 1981
rect 174 1976 175 1980
rect 179 1976 180 1980
rect 174 1975 180 1976
rect 318 1980 324 1981
rect 318 1976 319 1980
rect 323 1976 324 1980
rect 318 1975 324 1976
rect 462 1980 468 1981
rect 462 1976 463 1980
rect 467 1976 468 1980
rect 462 1975 468 1976
rect 614 1980 620 1981
rect 614 1976 615 1980
rect 619 1976 620 1980
rect 614 1975 620 1976
rect 758 1980 764 1981
rect 758 1976 759 1980
rect 763 1976 764 1980
rect 758 1975 764 1976
rect 902 1980 908 1981
rect 902 1976 903 1980
rect 907 1976 908 1980
rect 902 1975 908 1976
rect 1038 1980 1044 1981
rect 1038 1976 1039 1980
rect 1043 1976 1044 1980
rect 1038 1975 1044 1976
rect 1174 1980 1180 1981
rect 1174 1976 1175 1980
rect 1179 1976 1180 1980
rect 1174 1975 1180 1976
rect 1310 1980 1316 1981
rect 1310 1976 1311 1980
rect 1315 1976 1316 1980
rect 1310 1975 1316 1976
rect 1454 1980 1460 1981
rect 1454 1976 1455 1980
rect 1459 1976 1460 1980
rect 1830 1979 1831 1983
rect 1835 1979 1836 1983
rect 1830 1978 1836 1979
rect 1870 1979 1876 1980
rect 1454 1975 1460 1976
rect 1870 1975 1871 1979
rect 1875 1975 1876 1979
rect 3590 1979 3596 1980
rect 1870 1974 1876 1975
rect 2174 1976 2180 1977
rect 2174 1972 2175 1976
rect 2179 1972 2180 1976
rect 2174 1971 2180 1972
rect 2262 1976 2268 1977
rect 2262 1972 2263 1976
rect 2267 1972 2268 1976
rect 2262 1971 2268 1972
rect 2358 1976 2364 1977
rect 2358 1972 2359 1976
rect 2363 1972 2364 1976
rect 2358 1971 2364 1972
rect 2454 1976 2460 1977
rect 2454 1972 2455 1976
rect 2459 1972 2460 1976
rect 2454 1971 2460 1972
rect 2558 1976 2564 1977
rect 2558 1972 2559 1976
rect 2563 1972 2564 1976
rect 2558 1971 2564 1972
rect 2662 1976 2668 1977
rect 2662 1972 2663 1976
rect 2667 1972 2668 1976
rect 2662 1971 2668 1972
rect 2766 1976 2772 1977
rect 2766 1972 2767 1976
rect 2771 1972 2772 1976
rect 2766 1971 2772 1972
rect 2870 1976 2876 1977
rect 2870 1972 2871 1976
rect 2875 1972 2876 1976
rect 2870 1971 2876 1972
rect 2974 1976 2980 1977
rect 2974 1972 2975 1976
rect 2979 1972 2980 1976
rect 2974 1971 2980 1972
rect 3078 1976 3084 1977
rect 3078 1972 3079 1976
rect 3083 1972 3084 1976
rect 3078 1971 3084 1972
rect 3182 1976 3188 1977
rect 3182 1972 3183 1976
rect 3187 1972 3188 1976
rect 3590 1975 3591 1979
rect 3595 1975 3596 1979
rect 3590 1974 3596 1975
rect 3182 1971 3188 1972
rect 134 1936 140 1937
rect 110 1933 116 1934
rect 110 1929 111 1933
rect 115 1929 116 1933
rect 134 1932 135 1936
rect 139 1932 140 1936
rect 134 1931 140 1932
rect 294 1936 300 1937
rect 294 1932 295 1936
rect 299 1932 300 1936
rect 294 1931 300 1932
rect 462 1936 468 1937
rect 462 1932 463 1936
rect 467 1932 468 1936
rect 462 1931 468 1932
rect 630 1936 636 1937
rect 630 1932 631 1936
rect 635 1932 636 1936
rect 630 1931 636 1932
rect 798 1936 804 1937
rect 798 1932 799 1936
rect 803 1932 804 1936
rect 798 1931 804 1932
rect 950 1936 956 1937
rect 950 1932 951 1936
rect 955 1932 956 1936
rect 950 1931 956 1932
rect 1094 1936 1100 1937
rect 1094 1932 1095 1936
rect 1099 1932 1100 1936
rect 1094 1931 1100 1932
rect 1230 1936 1236 1937
rect 1230 1932 1231 1936
rect 1235 1932 1236 1936
rect 1230 1931 1236 1932
rect 1358 1936 1364 1937
rect 1358 1932 1359 1936
rect 1363 1932 1364 1936
rect 1358 1931 1364 1932
rect 1486 1936 1492 1937
rect 1486 1932 1487 1936
rect 1491 1932 1492 1936
rect 1486 1931 1492 1932
rect 1622 1936 1628 1937
rect 1622 1932 1623 1936
rect 1627 1932 1628 1936
rect 1622 1931 1628 1932
rect 1830 1933 1836 1934
rect 110 1928 116 1929
rect 1830 1929 1831 1933
rect 1835 1929 1836 1933
rect 1830 1928 1836 1929
rect 1942 1928 1948 1929
rect 1870 1925 1876 1926
rect 1870 1921 1871 1925
rect 1875 1921 1876 1925
rect 1942 1924 1943 1928
rect 1947 1924 1948 1928
rect 1942 1923 1948 1924
rect 2054 1928 2060 1929
rect 2054 1924 2055 1928
rect 2059 1924 2060 1928
rect 2054 1923 2060 1924
rect 2166 1928 2172 1929
rect 2166 1924 2167 1928
rect 2171 1924 2172 1928
rect 2166 1923 2172 1924
rect 2286 1928 2292 1929
rect 2286 1924 2287 1928
rect 2291 1924 2292 1928
rect 2286 1923 2292 1924
rect 2406 1928 2412 1929
rect 2406 1924 2407 1928
rect 2411 1924 2412 1928
rect 2406 1923 2412 1924
rect 2526 1928 2532 1929
rect 2526 1924 2527 1928
rect 2531 1924 2532 1928
rect 2526 1923 2532 1924
rect 2646 1928 2652 1929
rect 2646 1924 2647 1928
rect 2651 1924 2652 1928
rect 2646 1923 2652 1924
rect 2774 1928 2780 1929
rect 2774 1924 2775 1928
rect 2779 1924 2780 1928
rect 2774 1923 2780 1924
rect 2910 1928 2916 1929
rect 2910 1924 2911 1928
rect 2915 1924 2916 1928
rect 2910 1923 2916 1924
rect 3054 1928 3060 1929
rect 3054 1924 3055 1928
rect 3059 1924 3060 1928
rect 3054 1923 3060 1924
rect 3206 1928 3212 1929
rect 3206 1924 3207 1928
rect 3211 1924 3212 1928
rect 3206 1923 3212 1924
rect 3366 1928 3372 1929
rect 3366 1924 3367 1928
rect 3371 1924 3372 1928
rect 3366 1923 3372 1924
rect 3502 1928 3508 1929
rect 3502 1924 3503 1928
rect 3507 1924 3508 1928
rect 3502 1923 3508 1924
rect 3590 1925 3596 1926
rect 1870 1920 1876 1921
rect 3590 1921 3591 1925
rect 3595 1921 3596 1925
rect 3590 1920 3596 1921
rect 110 1916 116 1917
rect 110 1912 111 1916
rect 115 1912 116 1916
rect 110 1911 116 1912
rect 1830 1916 1836 1917
rect 1830 1912 1831 1916
rect 1835 1912 1836 1916
rect 1830 1911 1836 1912
rect 1870 1908 1876 1909
rect 1870 1904 1871 1908
rect 1875 1904 1876 1908
rect 1870 1903 1876 1904
rect 3590 1908 3596 1909
rect 3590 1904 3591 1908
rect 3595 1904 3596 1908
rect 3590 1903 3596 1904
rect 142 1898 148 1899
rect 142 1894 143 1898
rect 147 1894 148 1898
rect 142 1893 148 1894
rect 302 1898 308 1899
rect 302 1894 303 1898
rect 307 1894 308 1898
rect 302 1893 308 1894
rect 470 1898 476 1899
rect 470 1894 471 1898
rect 475 1894 476 1898
rect 470 1893 476 1894
rect 638 1898 644 1899
rect 638 1894 639 1898
rect 643 1894 644 1898
rect 638 1893 644 1894
rect 806 1898 812 1899
rect 806 1894 807 1898
rect 811 1894 812 1898
rect 806 1893 812 1894
rect 958 1898 964 1899
rect 958 1894 959 1898
rect 963 1894 964 1898
rect 958 1893 964 1894
rect 1102 1898 1108 1899
rect 1102 1894 1103 1898
rect 1107 1894 1108 1898
rect 1102 1893 1108 1894
rect 1238 1898 1244 1899
rect 1238 1894 1239 1898
rect 1243 1894 1244 1898
rect 1238 1893 1244 1894
rect 1366 1898 1372 1899
rect 1366 1894 1367 1898
rect 1371 1894 1372 1898
rect 1366 1893 1372 1894
rect 1494 1898 1500 1899
rect 1494 1894 1495 1898
rect 1499 1894 1500 1898
rect 1494 1893 1500 1894
rect 1630 1898 1636 1899
rect 1630 1894 1631 1898
rect 1635 1894 1636 1898
rect 1630 1893 1636 1894
rect 1950 1890 1956 1891
rect 1950 1886 1951 1890
rect 1955 1886 1956 1890
rect 1950 1885 1956 1886
rect 2062 1890 2068 1891
rect 2062 1886 2063 1890
rect 2067 1886 2068 1890
rect 2062 1885 2068 1886
rect 2174 1890 2180 1891
rect 2174 1886 2175 1890
rect 2179 1886 2180 1890
rect 2174 1885 2180 1886
rect 2294 1890 2300 1891
rect 2294 1886 2295 1890
rect 2299 1886 2300 1890
rect 2294 1885 2300 1886
rect 2414 1890 2420 1891
rect 2414 1886 2415 1890
rect 2419 1886 2420 1890
rect 2414 1885 2420 1886
rect 2534 1890 2540 1891
rect 2534 1886 2535 1890
rect 2539 1886 2540 1890
rect 2534 1885 2540 1886
rect 2654 1890 2660 1891
rect 2654 1886 2655 1890
rect 2659 1886 2660 1890
rect 2654 1885 2660 1886
rect 2782 1890 2788 1891
rect 2782 1886 2783 1890
rect 2787 1886 2788 1890
rect 2782 1885 2788 1886
rect 2918 1890 2924 1891
rect 2918 1886 2919 1890
rect 2923 1886 2924 1890
rect 2918 1885 2924 1886
rect 3062 1890 3068 1891
rect 3062 1886 3063 1890
rect 3067 1886 3068 1890
rect 3062 1885 3068 1886
rect 3214 1890 3220 1891
rect 3214 1886 3215 1890
rect 3219 1886 3220 1890
rect 3214 1885 3220 1886
rect 3374 1890 3380 1891
rect 3374 1886 3375 1890
rect 3379 1886 3380 1890
rect 3374 1885 3380 1886
rect 3510 1890 3516 1891
rect 3510 1886 3511 1890
rect 3515 1886 3516 1890
rect 3510 1885 3516 1886
rect 142 1858 148 1859
rect 142 1854 143 1858
rect 147 1854 148 1858
rect 142 1853 148 1854
rect 318 1858 324 1859
rect 318 1854 319 1858
rect 323 1854 324 1858
rect 318 1853 324 1854
rect 518 1858 524 1859
rect 518 1854 519 1858
rect 523 1854 524 1858
rect 518 1853 524 1854
rect 710 1858 716 1859
rect 710 1854 711 1858
rect 715 1854 716 1858
rect 710 1853 716 1854
rect 886 1858 892 1859
rect 886 1854 887 1858
rect 891 1854 892 1858
rect 886 1853 892 1854
rect 1054 1858 1060 1859
rect 1054 1854 1055 1858
rect 1059 1854 1060 1858
rect 1054 1853 1060 1854
rect 1206 1858 1212 1859
rect 1206 1854 1207 1858
rect 1211 1854 1212 1858
rect 1206 1853 1212 1854
rect 1342 1858 1348 1859
rect 1342 1854 1343 1858
rect 1347 1854 1348 1858
rect 1342 1853 1348 1854
rect 1470 1858 1476 1859
rect 1470 1854 1471 1858
rect 1475 1854 1476 1858
rect 1470 1853 1476 1854
rect 1598 1858 1604 1859
rect 1598 1854 1599 1858
rect 1603 1854 1604 1858
rect 1598 1853 1604 1854
rect 1726 1858 1732 1859
rect 1726 1854 1727 1858
rect 1731 1854 1732 1858
rect 1726 1853 1732 1854
rect 1902 1854 1908 1855
rect 1902 1850 1903 1854
rect 1907 1850 1908 1854
rect 1902 1849 1908 1850
rect 1982 1854 1988 1855
rect 1982 1850 1983 1854
rect 1987 1850 1988 1854
rect 1982 1849 1988 1850
rect 2094 1854 2100 1855
rect 2094 1850 2095 1854
rect 2099 1850 2100 1854
rect 2094 1849 2100 1850
rect 2206 1854 2212 1855
rect 2206 1850 2207 1854
rect 2211 1850 2212 1854
rect 2206 1849 2212 1850
rect 2326 1854 2332 1855
rect 2326 1850 2327 1854
rect 2331 1850 2332 1854
rect 2326 1849 2332 1850
rect 2462 1854 2468 1855
rect 2462 1850 2463 1854
rect 2467 1850 2468 1854
rect 2462 1849 2468 1850
rect 2630 1854 2636 1855
rect 2630 1850 2631 1854
rect 2635 1850 2636 1854
rect 2630 1849 2636 1850
rect 2830 1854 2836 1855
rect 2830 1850 2831 1854
rect 2835 1850 2836 1854
rect 2830 1849 2836 1850
rect 3054 1854 3060 1855
rect 3054 1850 3055 1854
rect 3059 1850 3060 1854
rect 3054 1849 3060 1850
rect 3294 1854 3300 1855
rect 3294 1850 3295 1854
rect 3299 1850 3300 1854
rect 3294 1849 3300 1850
rect 3510 1854 3516 1855
rect 3510 1850 3511 1854
rect 3515 1850 3516 1854
rect 3510 1849 3516 1850
rect 110 1840 116 1841
rect 110 1836 111 1840
rect 115 1836 116 1840
rect 110 1835 116 1836
rect 1830 1840 1836 1841
rect 1830 1836 1831 1840
rect 1835 1836 1836 1840
rect 1830 1835 1836 1836
rect 1870 1836 1876 1837
rect 1870 1832 1871 1836
rect 1875 1832 1876 1836
rect 1870 1831 1876 1832
rect 3590 1836 3596 1837
rect 3590 1832 3591 1836
rect 3595 1832 3596 1836
rect 3590 1831 3596 1832
rect 110 1823 116 1824
rect 110 1819 111 1823
rect 115 1819 116 1823
rect 1830 1823 1836 1824
rect 110 1818 116 1819
rect 134 1820 140 1821
rect 134 1816 135 1820
rect 139 1816 140 1820
rect 134 1815 140 1816
rect 310 1820 316 1821
rect 310 1816 311 1820
rect 315 1816 316 1820
rect 310 1815 316 1816
rect 510 1820 516 1821
rect 510 1816 511 1820
rect 515 1816 516 1820
rect 510 1815 516 1816
rect 702 1820 708 1821
rect 702 1816 703 1820
rect 707 1816 708 1820
rect 702 1815 708 1816
rect 878 1820 884 1821
rect 878 1816 879 1820
rect 883 1816 884 1820
rect 878 1815 884 1816
rect 1046 1820 1052 1821
rect 1046 1816 1047 1820
rect 1051 1816 1052 1820
rect 1046 1815 1052 1816
rect 1198 1820 1204 1821
rect 1198 1816 1199 1820
rect 1203 1816 1204 1820
rect 1198 1815 1204 1816
rect 1334 1820 1340 1821
rect 1334 1816 1335 1820
rect 1339 1816 1340 1820
rect 1334 1815 1340 1816
rect 1462 1820 1468 1821
rect 1462 1816 1463 1820
rect 1467 1816 1468 1820
rect 1462 1815 1468 1816
rect 1590 1820 1596 1821
rect 1590 1816 1591 1820
rect 1595 1816 1596 1820
rect 1590 1815 1596 1816
rect 1718 1820 1724 1821
rect 1718 1816 1719 1820
rect 1723 1816 1724 1820
rect 1830 1819 1831 1823
rect 1835 1819 1836 1823
rect 1830 1818 1836 1819
rect 1870 1819 1876 1820
rect 1718 1815 1724 1816
rect 1870 1815 1871 1819
rect 1875 1815 1876 1819
rect 3590 1819 3596 1820
rect 1870 1814 1876 1815
rect 1894 1816 1900 1817
rect 1894 1812 1895 1816
rect 1899 1812 1900 1816
rect 1894 1811 1900 1812
rect 1974 1816 1980 1817
rect 1974 1812 1975 1816
rect 1979 1812 1980 1816
rect 1974 1811 1980 1812
rect 2086 1816 2092 1817
rect 2086 1812 2087 1816
rect 2091 1812 2092 1816
rect 2086 1811 2092 1812
rect 2198 1816 2204 1817
rect 2198 1812 2199 1816
rect 2203 1812 2204 1816
rect 2198 1811 2204 1812
rect 2318 1816 2324 1817
rect 2318 1812 2319 1816
rect 2323 1812 2324 1816
rect 2318 1811 2324 1812
rect 2454 1816 2460 1817
rect 2454 1812 2455 1816
rect 2459 1812 2460 1816
rect 2454 1811 2460 1812
rect 2622 1816 2628 1817
rect 2622 1812 2623 1816
rect 2627 1812 2628 1816
rect 2622 1811 2628 1812
rect 2822 1816 2828 1817
rect 2822 1812 2823 1816
rect 2827 1812 2828 1816
rect 2822 1811 2828 1812
rect 3046 1816 3052 1817
rect 3046 1812 3047 1816
rect 3051 1812 3052 1816
rect 3046 1811 3052 1812
rect 3286 1816 3292 1817
rect 3286 1812 3287 1816
rect 3291 1812 3292 1816
rect 3286 1811 3292 1812
rect 3502 1816 3508 1817
rect 3502 1812 3503 1816
rect 3507 1812 3508 1816
rect 3590 1815 3591 1819
rect 3595 1815 3596 1819
rect 3590 1814 3596 1815
rect 3502 1811 3508 1812
rect 134 1776 140 1777
rect 110 1773 116 1774
rect 110 1769 111 1773
rect 115 1769 116 1773
rect 134 1772 135 1776
rect 139 1772 140 1776
rect 134 1771 140 1772
rect 310 1776 316 1777
rect 310 1772 311 1776
rect 315 1772 316 1776
rect 310 1771 316 1772
rect 502 1776 508 1777
rect 502 1772 503 1776
rect 507 1772 508 1776
rect 502 1771 508 1772
rect 686 1776 692 1777
rect 686 1772 687 1776
rect 691 1772 692 1776
rect 686 1771 692 1772
rect 846 1776 852 1777
rect 846 1772 847 1776
rect 851 1772 852 1776
rect 846 1771 852 1772
rect 990 1776 996 1777
rect 990 1772 991 1776
rect 995 1772 996 1776
rect 990 1771 996 1772
rect 1126 1776 1132 1777
rect 1126 1772 1127 1776
rect 1131 1772 1132 1776
rect 1126 1771 1132 1772
rect 1246 1776 1252 1777
rect 1246 1772 1247 1776
rect 1251 1772 1252 1776
rect 1246 1771 1252 1772
rect 1358 1776 1364 1777
rect 1358 1772 1359 1776
rect 1363 1772 1364 1776
rect 1358 1771 1364 1772
rect 1462 1776 1468 1777
rect 1462 1772 1463 1776
rect 1467 1772 1468 1776
rect 1462 1771 1468 1772
rect 1558 1776 1564 1777
rect 1558 1772 1559 1776
rect 1563 1772 1564 1776
rect 1558 1771 1564 1772
rect 1662 1776 1668 1777
rect 1662 1772 1663 1776
rect 1667 1772 1668 1776
rect 1662 1771 1668 1772
rect 1742 1776 1748 1777
rect 1742 1772 1743 1776
rect 1747 1772 1748 1776
rect 1742 1771 1748 1772
rect 1830 1773 1836 1774
rect 110 1768 116 1769
rect 1830 1769 1831 1773
rect 1835 1769 1836 1773
rect 1830 1768 1836 1769
rect 110 1756 116 1757
rect 110 1752 111 1756
rect 115 1752 116 1756
rect 110 1751 116 1752
rect 1830 1756 1836 1757
rect 1830 1752 1831 1756
rect 1835 1752 1836 1756
rect 1894 1756 1900 1757
rect 1830 1751 1836 1752
rect 1870 1753 1876 1754
rect 1870 1749 1871 1753
rect 1875 1749 1876 1753
rect 1894 1752 1895 1756
rect 1899 1752 1900 1756
rect 1894 1751 1900 1752
rect 2022 1756 2028 1757
rect 2022 1752 2023 1756
rect 2027 1752 2028 1756
rect 2022 1751 2028 1752
rect 2182 1756 2188 1757
rect 2182 1752 2183 1756
rect 2187 1752 2188 1756
rect 2182 1751 2188 1752
rect 2350 1756 2356 1757
rect 2350 1752 2351 1756
rect 2355 1752 2356 1756
rect 2350 1751 2356 1752
rect 2550 1756 2556 1757
rect 2550 1752 2551 1756
rect 2555 1752 2556 1756
rect 2550 1751 2556 1752
rect 2774 1756 2780 1757
rect 2774 1752 2775 1756
rect 2779 1752 2780 1756
rect 2774 1751 2780 1752
rect 3014 1756 3020 1757
rect 3014 1752 3015 1756
rect 3019 1752 3020 1756
rect 3014 1751 3020 1752
rect 3270 1756 3276 1757
rect 3270 1752 3271 1756
rect 3275 1752 3276 1756
rect 3270 1751 3276 1752
rect 3502 1756 3508 1757
rect 3502 1752 3503 1756
rect 3507 1752 3508 1756
rect 3502 1751 3508 1752
rect 3590 1753 3596 1754
rect 1870 1748 1876 1749
rect 3590 1749 3591 1753
rect 3595 1749 3596 1753
rect 3590 1748 3596 1749
rect 142 1738 148 1739
rect 142 1734 143 1738
rect 147 1734 148 1738
rect 142 1733 148 1734
rect 318 1738 324 1739
rect 318 1734 319 1738
rect 323 1734 324 1738
rect 318 1733 324 1734
rect 510 1738 516 1739
rect 510 1734 511 1738
rect 515 1734 516 1738
rect 510 1733 516 1734
rect 694 1738 700 1739
rect 694 1734 695 1738
rect 699 1734 700 1738
rect 694 1733 700 1734
rect 854 1738 860 1739
rect 854 1734 855 1738
rect 859 1734 860 1738
rect 854 1733 860 1734
rect 998 1738 1004 1739
rect 998 1734 999 1738
rect 1003 1734 1004 1738
rect 998 1733 1004 1734
rect 1134 1738 1140 1739
rect 1134 1734 1135 1738
rect 1139 1734 1140 1738
rect 1134 1733 1140 1734
rect 1254 1738 1260 1739
rect 1254 1734 1255 1738
rect 1259 1734 1260 1738
rect 1254 1733 1260 1734
rect 1366 1738 1372 1739
rect 1366 1734 1367 1738
rect 1371 1734 1372 1738
rect 1366 1733 1372 1734
rect 1470 1738 1476 1739
rect 1470 1734 1471 1738
rect 1475 1734 1476 1738
rect 1470 1733 1476 1734
rect 1566 1738 1572 1739
rect 1566 1734 1567 1738
rect 1571 1734 1572 1738
rect 1566 1733 1572 1734
rect 1670 1738 1676 1739
rect 1670 1734 1671 1738
rect 1675 1734 1676 1738
rect 1670 1733 1676 1734
rect 1750 1738 1756 1739
rect 1750 1734 1751 1738
rect 1755 1734 1756 1738
rect 1750 1733 1756 1734
rect 1870 1736 1876 1737
rect 1870 1732 1871 1736
rect 1875 1732 1876 1736
rect 1870 1731 1876 1732
rect 3590 1736 3596 1737
rect 3590 1732 3591 1736
rect 3595 1732 3596 1736
rect 3590 1731 3596 1732
rect 1902 1718 1908 1719
rect 1902 1714 1903 1718
rect 1907 1714 1908 1718
rect 1902 1713 1908 1714
rect 2030 1718 2036 1719
rect 2030 1714 2031 1718
rect 2035 1714 2036 1718
rect 2030 1713 2036 1714
rect 2190 1718 2196 1719
rect 2190 1714 2191 1718
rect 2195 1714 2196 1718
rect 2190 1713 2196 1714
rect 2358 1718 2364 1719
rect 2358 1714 2359 1718
rect 2363 1714 2364 1718
rect 2358 1713 2364 1714
rect 2558 1718 2564 1719
rect 2558 1714 2559 1718
rect 2563 1714 2564 1718
rect 2558 1713 2564 1714
rect 2782 1718 2788 1719
rect 2782 1714 2783 1718
rect 2787 1714 2788 1718
rect 2782 1713 2788 1714
rect 3022 1718 3028 1719
rect 3022 1714 3023 1718
rect 3027 1714 3028 1718
rect 3022 1713 3028 1714
rect 3278 1718 3284 1719
rect 3278 1714 3279 1718
rect 3283 1714 3284 1718
rect 3278 1713 3284 1714
rect 3510 1718 3516 1719
rect 3510 1714 3511 1718
rect 3515 1714 3516 1718
rect 3510 1713 3516 1714
rect 142 1698 148 1699
rect 142 1694 143 1698
rect 147 1694 148 1698
rect 142 1693 148 1694
rect 238 1698 244 1699
rect 238 1694 239 1698
rect 243 1694 244 1698
rect 238 1693 244 1694
rect 366 1698 372 1699
rect 366 1694 367 1698
rect 371 1694 372 1698
rect 366 1693 372 1694
rect 486 1698 492 1699
rect 486 1694 487 1698
rect 491 1694 492 1698
rect 486 1693 492 1694
rect 606 1698 612 1699
rect 606 1694 607 1698
rect 611 1694 612 1698
rect 606 1693 612 1694
rect 718 1698 724 1699
rect 718 1694 719 1698
rect 723 1694 724 1698
rect 718 1693 724 1694
rect 822 1698 828 1699
rect 822 1694 823 1698
rect 827 1694 828 1698
rect 822 1693 828 1694
rect 926 1698 932 1699
rect 926 1694 927 1698
rect 931 1694 932 1698
rect 926 1693 932 1694
rect 1022 1698 1028 1699
rect 1022 1694 1023 1698
rect 1027 1694 1028 1698
rect 1022 1693 1028 1694
rect 1118 1698 1124 1699
rect 1118 1694 1119 1698
rect 1123 1694 1124 1698
rect 1118 1693 1124 1694
rect 1214 1698 1220 1699
rect 1214 1694 1215 1698
rect 1219 1694 1220 1698
rect 1214 1693 1220 1694
rect 1318 1698 1324 1699
rect 1318 1694 1319 1698
rect 1323 1694 1324 1698
rect 1318 1693 1324 1694
rect 1902 1686 1908 1687
rect 1902 1682 1903 1686
rect 1907 1682 1908 1686
rect 1902 1681 1908 1682
rect 1990 1686 1996 1687
rect 1990 1682 1991 1686
rect 1995 1682 1996 1686
rect 1990 1681 1996 1682
rect 2110 1686 2116 1687
rect 2110 1682 2111 1686
rect 2115 1682 2116 1686
rect 2110 1681 2116 1682
rect 2230 1686 2236 1687
rect 2230 1682 2231 1686
rect 2235 1682 2236 1686
rect 2230 1681 2236 1682
rect 2350 1686 2356 1687
rect 2350 1682 2351 1686
rect 2355 1682 2356 1686
rect 2350 1681 2356 1682
rect 2478 1686 2484 1687
rect 2478 1682 2479 1686
rect 2483 1682 2484 1686
rect 2478 1681 2484 1682
rect 2606 1686 2612 1687
rect 2606 1682 2607 1686
rect 2611 1682 2612 1686
rect 2606 1681 2612 1682
rect 2742 1686 2748 1687
rect 2742 1682 2743 1686
rect 2747 1682 2748 1686
rect 2742 1681 2748 1682
rect 2886 1686 2892 1687
rect 2886 1682 2887 1686
rect 2891 1682 2892 1686
rect 2886 1681 2892 1682
rect 3038 1686 3044 1687
rect 3038 1682 3039 1686
rect 3043 1682 3044 1686
rect 3038 1681 3044 1682
rect 3198 1686 3204 1687
rect 3198 1682 3199 1686
rect 3203 1682 3204 1686
rect 3198 1681 3204 1682
rect 3366 1686 3372 1687
rect 3366 1682 3367 1686
rect 3371 1682 3372 1686
rect 3366 1681 3372 1682
rect 3510 1686 3516 1687
rect 3510 1682 3511 1686
rect 3515 1682 3516 1686
rect 3510 1681 3516 1682
rect 110 1680 116 1681
rect 110 1676 111 1680
rect 115 1676 116 1680
rect 110 1675 116 1676
rect 1830 1680 1836 1681
rect 1830 1676 1831 1680
rect 1835 1676 1836 1680
rect 1830 1675 1836 1676
rect 1870 1668 1876 1669
rect 1870 1664 1871 1668
rect 1875 1664 1876 1668
rect 110 1663 116 1664
rect 110 1659 111 1663
rect 115 1659 116 1663
rect 1830 1663 1836 1664
rect 1870 1663 1876 1664
rect 3590 1668 3596 1669
rect 3590 1664 3591 1668
rect 3595 1664 3596 1668
rect 3590 1663 3596 1664
rect 110 1658 116 1659
rect 134 1660 140 1661
rect 134 1656 135 1660
rect 139 1656 140 1660
rect 134 1655 140 1656
rect 230 1660 236 1661
rect 230 1656 231 1660
rect 235 1656 236 1660
rect 230 1655 236 1656
rect 358 1660 364 1661
rect 358 1656 359 1660
rect 363 1656 364 1660
rect 358 1655 364 1656
rect 478 1660 484 1661
rect 478 1656 479 1660
rect 483 1656 484 1660
rect 478 1655 484 1656
rect 598 1660 604 1661
rect 598 1656 599 1660
rect 603 1656 604 1660
rect 598 1655 604 1656
rect 710 1660 716 1661
rect 710 1656 711 1660
rect 715 1656 716 1660
rect 710 1655 716 1656
rect 814 1660 820 1661
rect 814 1656 815 1660
rect 819 1656 820 1660
rect 814 1655 820 1656
rect 918 1660 924 1661
rect 918 1656 919 1660
rect 923 1656 924 1660
rect 918 1655 924 1656
rect 1014 1660 1020 1661
rect 1014 1656 1015 1660
rect 1019 1656 1020 1660
rect 1014 1655 1020 1656
rect 1110 1660 1116 1661
rect 1110 1656 1111 1660
rect 1115 1656 1116 1660
rect 1110 1655 1116 1656
rect 1206 1660 1212 1661
rect 1206 1656 1207 1660
rect 1211 1656 1212 1660
rect 1206 1655 1212 1656
rect 1310 1660 1316 1661
rect 1310 1656 1311 1660
rect 1315 1656 1316 1660
rect 1830 1659 1831 1663
rect 1835 1659 1836 1663
rect 1830 1658 1836 1659
rect 1310 1655 1316 1656
rect 1870 1651 1876 1652
rect 1870 1647 1871 1651
rect 1875 1647 1876 1651
rect 3590 1651 3596 1652
rect 1870 1646 1876 1647
rect 1894 1648 1900 1649
rect 1894 1644 1895 1648
rect 1899 1644 1900 1648
rect 1894 1643 1900 1644
rect 1982 1648 1988 1649
rect 1982 1644 1983 1648
rect 1987 1644 1988 1648
rect 1982 1643 1988 1644
rect 2102 1648 2108 1649
rect 2102 1644 2103 1648
rect 2107 1644 2108 1648
rect 2102 1643 2108 1644
rect 2222 1648 2228 1649
rect 2222 1644 2223 1648
rect 2227 1644 2228 1648
rect 2222 1643 2228 1644
rect 2342 1648 2348 1649
rect 2342 1644 2343 1648
rect 2347 1644 2348 1648
rect 2342 1643 2348 1644
rect 2470 1648 2476 1649
rect 2470 1644 2471 1648
rect 2475 1644 2476 1648
rect 2470 1643 2476 1644
rect 2598 1648 2604 1649
rect 2598 1644 2599 1648
rect 2603 1644 2604 1648
rect 2598 1643 2604 1644
rect 2734 1648 2740 1649
rect 2734 1644 2735 1648
rect 2739 1644 2740 1648
rect 2734 1643 2740 1644
rect 2878 1648 2884 1649
rect 2878 1644 2879 1648
rect 2883 1644 2884 1648
rect 2878 1643 2884 1644
rect 3030 1648 3036 1649
rect 3030 1644 3031 1648
rect 3035 1644 3036 1648
rect 3030 1643 3036 1644
rect 3190 1648 3196 1649
rect 3190 1644 3191 1648
rect 3195 1644 3196 1648
rect 3190 1643 3196 1644
rect 3358 1648 3364 1649
rect 3358 1644 3359 1648
rect 3363 1644 3364 1648
rect 3358 1643 3364 1644
rect 3502 1648 3508 1649
rect 3502 1644 3503 1648
rect 3507 1644 3508 1648
rect 3590 1647 3591 1651
rect 3595 1647 3596 1651
rect 3590 1646 3596 1647
rect 3502 1643 3508 1644
rect 174 1608 180 1609
rect 110 1605 116 1606
rect 110 1601 111 1605
rect 115 1601 116 1605
rect 174 1604 175 1608
rect 179 1604 180 1608
rect 174 1603 180 1604
rect 310 1608 316 1609
rect 310 1604 311 1608
rect 315 1604 316 1608
rect 310 1603 316 1604
rect 438 1608 444 1609
rect 438 1604 439 1608
rect 443 1604 444 1608
rect 438 1603 444 1604
rect 566 1608 572 1609
rect 566 1604 567 1608
rect 571 1604 572 1608
rect 566 1603 572 1604
rect 686 1608 692 1609
rect 686 1604 687 1608
rect 691 1604 692 1608
rect 686 1603 692 1604
rect 798 1608 804 1609
rect 798 1604 799 1608
rect 803 1604 804 1608
rect 798 1603 804 1604
rect 902 1608 908 1609
rect 902 1604 903 1608
rect 907 1604 908 1608
rect 902 1603 908 1604
rect 998 1608 1004 1609
rect 998 1604 999 1608
rect 1003 1604 1004 1608
rect 998 1603 1004 1604
rect 1094 1608 1100 1609
rect 1094 1604 1095 1608
rect 1099 1604 1100 1608
rect 1094 1603 1100 1604
rect 1198 1608 1204 1609
rect 1198 1604 1199 1608
rect 1203 1604 1204 1608
rect 1198 1603 1204 1604
rect 1302 1608 1308 1609
rect 1302 1604 1303 1608
rect 1307 1604 1308 1608
rect 1302 1603 1308 1604
rect 1830 1605 1836 1606
rect 110 1600 116 1601
rect 1830 1601 1831 1605
rect 1835 1601 1836 1605
rect 1926 1604 1932 1605
rect 1830 1600 1836 1601
rect 1870 1601 1876 1602
rect 1870 1597 1871 1601
rect 1875 1597 1876 1601
rect 1926 1600 1927 1604
rect 1931 1600 1932 1604
rect 1926 1599 1932 1600
rect 2022 1604 2028 1605
rect 2022 1600 2023 1604
rect 2027 1600 2028 1604
rect 2022 1599 2028 1600
rect 2134 1604 2140 1605
rect 2134 1600 2135 1604
rect 2139 1600 2140 1604
rect 2134 1599 2140 1600
rect 2262 1604 2268 1605
rect 2262 1600 2263 1604
rect 2267 1600 2268 1604
rect 2262 1599 2268 1600
rect 2390 1604 2396 1605
rect 2390 1600 2391 1604
rect 2395 1600 2396 1604
rect 2390 1599 2396 1600
rect 2526 1604 2532 1605
rect 2526 1600 2527 1604
rect 2531 1600 2532 1604
rect 2526 1599 2532 1600
rect 2670 1604 2676 1605
rect 2670 1600 2671 1604
rect 2675 1600 2676 1604
rect 2670 1599 2676 1600
rect 2822 1604 2828 1605
rect 2822 1600 2823 1604
rect 2827 1600 2828 1604
rect 2822 1599 2828 1600
rect 2982 1604 2988 1605
rect 2982 1600 2983 1604
rect 2987 1600 2988 1604
rect 2982 1599 2988 1600
rect 3158 1604 3164 1605
rect 3158 1600 3159 1604
rect 3163 1600 3164 1604
rect 3158 1599 3164 1600
rect 3342 1604 3348 1605
rect 3342 1600 3343 1604
rect 3347 1600 3348 1604
rect 3342 1599 3348 1600
rect 3502 1604 3508 1605
rect 3502 1600 3503 1604
rect 3507 1600 3508 1604
rect 3502 1599 3508 1600
rect 3590 1601 3596 1602
rect 1870 1596 1876 1597
rect 3590 1597 3591 1601
rect 3595 1597 3596 1601
rect 3590 1596 3596 1597
rect 110 1588 116 1589
rect 110 1584 111 1588
rect 115 1584 116 1588
rect 110 1583 116 1584
rect 1830 1588 1836 1589
rect 1830 1584 1831 1588
rect 1835 1584 1836 1588
rect 1830 1583 1836 1584
rect 1870 1584 1876 1585
rect 1870 1580 1871 1584
rect 1875 1580 1876 1584
rect 1870 1579 1876 1580
rect 3590 1584 3596 1585
rect 3590 1580 3591 1584
rect 3595 1580 3596 1584
rect 3590 1579 3596 1580
rect 182 1570 188 1571
rect 182 1566 183 1570
rect 187 1566 188 1570
rect 182 1565 188 1566
rect 318 1570 324 1571
rect 318 1566 319 1570
rect 323 1566 324 1570
rect 318 1565 324 1566
rect 446 1570 452 1571
rect 446 1566 447 1570
rect 451 1566 452 1570
rect 446 1565 452 1566
rect 574 1570 580 1571
rect 574 1566 575 1570
rect 579 1566 580 1570
rect 574 1565 580 1566
rect 694 1570 700 1571
rect 694 1566 695 1570
rect 699 1566 700 1570
rect 694 1565 700 1566
rect 806 1570 812 1571
rect 806 1566 807 1570
rect 811 1566 812 1570
rect 806 1565 812 1566
rect 910 1570 916 1571
rect 910 1566 911 1570
rect 915 1566 916 1570
rect 910 1565 916 1566
rect 1006 1570 1012 1571
rect 1006 1566 1007 1570
rect 1011 1566 1012 1570
rect 1006 1565 1012 1566
rect 1102 1570 1108 1571
rect 1102 1566 1103 1570
rect 1107 1566 1108 1570
rect 1102 1565 1108 1566
rect 1206 1570 1212 1571
rect 1206 1566 1207 1570
rect 1211 1566 1212 1570
rect 1206 1565 1212 1566
rect 1310 1570 1316 1571
rect 1310 1566 1311 1570
rect 1315 1566 1316 1570
rect 1310 1565 1316 1566
rect 1934 1566 1940 1567
rect 1934 1562 1935 1566
rect 1939 1562 1940 1566
rect 1934 1561 1940 1562
rect 2030 1566 2036 1567
rect 2030 1562 2031 1566
rect 2035 1562 2036 1566
rect 2030 1561 2036 1562
rect 2142 1566 2148 1567
rect 2142 1562 2143 1566
rect 2147 1562 2148 1566
rect 2142 1561 2148 1562
rect 2270 1566 2276 1567
rect 2270 1562 2271 1566
rect 2275 1562 2276 1566
rect 2270 1561 2276 1562
rect 2398 1566 2404 1567
rect 2398 1562 2399 1566
rect 2403 1562 2404 1566
rect 2398 1561 2404 1562
rect 2534 1566 2540 1567
rect 2534 1562 2535 1566
rect 2539 1562 2540 1566
rect 2534 1561 2540 1562
rect 2678 1566 2684 1567
rect 2678 1562 2679 1566
rect 2683 1562 2684 1566
rect 2678 1561 2684 1562
rect 2830 1566 2836 1567
rect 2830 1562 2831 1566
rect 2835 1562 2836 1566
rect 2830 1561 2836 1562
rect 2990 1566 2996 1567
rect 2990 1562 2991 1566
rect 2995 1562 2996 1566
rect 2990 1561 2996 1562
rect 3166 1566 3172 1567
rect 3166 1562 3167 1566
rect 3171 1562 3172 1566
rect 3166 1561 3172 1562
rect 3350 1566 3356 1567
rect 3350 1562 3351 1566
rect 3355 1562 3356 1566
rect 3350 1561 3356 1562
rect 3510 1566 3516 1567
rect 3510 1562 3511 1566
rect 3515 1562 3516 1566
rect 3510 1561 3516 1562
rect 238 1530 244 1531
rect 238 1526 239 1530
rect 243 1526 244 1530
rect 238 1525 244 1526
rect 342 1530 348 1531
rect 342 1526 343 1530
rect 347 1526 348 1530
rect 342 1525 348 1526
rect 462 1530 468 1531
rect 462 1526 463 1530
rect 467 1526 468 1530
rect 462 1525 468 1526
rect 590 1530 596 1531
rect 590 1526 591 1530
rect 595 1526 596 1530
rect 590 1525 596 1526
rect 718 1530 724 1531
rect 718 1526 719 1530
rect 723 1526 724 1530
rect 718 1525 724 1526
rect 854 1530 860 1531
rect 854 1526 855 1530
rect 859 1526 860 1530
rect 854 1525 860 1526
rect 982 1530 988 1531
rect 982 1526 983 1530
rect 987 1526 988 1530
rect 982 1525 988 1526
rect 1110 1530 1116 1531
rect 1110 1526 1111 1530
rect 1115 1526 1116 1530
rect 1110 1525 1116 1526
rect 1230 1530 1236 1531
rect 1230 1526 1231 1530
rect 1235 1526 1236 1530
rect 1230 1525 1236 1526
rect 1342 1530 1348 1531
rect 1342 1526 1343 1530
rect 1347 1526 1348 1530
rect 1342 1525 1348 1526
rect 1454 1530 1460 1531
rect 1454 1526 1455 1530
rect 1459 1526 1460 1530
rect 1454 1525 1460 1526
rect 1574 1530 1580 1531
rect 1574 1526 1575 1530
rect 1579 1526 1580 1530
rect 1574 1525 1580 1526
rect 2134 1526 2140 1527
rect 2134 1522 2135 1526
rect 2139 1522 2140 1526
rect 2134 1521 2140 1522
rect 2254 1526 2260 1527
rect 2254 1522 2255 1526
rect 2259 1522 2260 1526
rect 2254 1521 2260 1522
rect 2382 1526 2388 1527
rect 2382 1522 2383 1526
rect 2387 1522 2388 1526
rect 2382 1521 2388 1522
rect 2510 1526 2516 1527
rect 2510 1522 2511 1526
rect 2515 1522 2516 1526
rect 2510 1521 2516 1522
rect 2638 1526 2644 1527
rect 2638 1522 2639 1526
rect 2643 1522 2644 1526
rect 2638 1521 2644 1522
rect 2766 1526 2772 1527
rect 2766 1522 2767 1526
rect 2771 1522 2772 1526
rect 2766 1521 2772 1522
rect 2886 1526 2892 1527
rect 2886 1522 2887 1526
rect 2891 1522 2892 1526
rect 2886 1521 2892 1522
rect 3006 1526 3012 1527
rect 3006 1522 3007 1526
rect 3011 1522 3012 1526
rect 3006 1521 3012 1522
rect 3118 1526 3124 1527
rect 3118 1522 3119 1526
rect 3123 1522 3124 1526
rect 3118 1521 3124 1522
rect 3230 1526 3236 1527
rect 3230 1522 3231 1526
rect 3235 1522 3236 1526
rect 3230 1521 3236 1522
rect 3350 1526 3356 1527
rect 3350 1522 3351 1526
rect 3355 1522 3356 1526
rect 3350 1521 3356 1522
rect 110 1512 116 1513
rect 110 1508 111 1512
rect 115 1508 116 1512
rect 110 1507 116 1508
rect 1830 1512 1836 1513
rect 1830 1508 1831 1512
rect 1835 1508 1836 1512
rect 1830 1507 1836 1508
rect 1870 1508 1876 1509
rect 1870 1504 1871 1508
rect 1875 1504 1876 1508
rect 1870 1503 1876 1504
rect 3590 1508 3596 1509
rect 3590 1504 3591 1508
rect 3595 1504 3596 1508
rect 3590 1503 3596 1504
rect 110 1495 116 1496
rect 110 1491 111 1495
rect 115 1491 116 1495
rect 1830 1495 1836 1496
rect 110 1490 116 1491
rect 230 1492 236 1493
rect 230 1488 231 1492
rect 235 1488 236 1492
rect 230 1487 236 1488
rect 334 1492 340 1493
rect 334 1488 335 1492
rect 339 1488 340 1492
rect 334 1487 340 1488
rect 454 1492 460 1493
rect 454 1488 455 1492
rect 459 1488 460 1492
rect 454 1487 460 1488
rect 582 1492 588 1493
rect 582 1488 583 1492
rect 587 1488 588 1492
rect 582 1487 588 1488
rect 710 1492 716 1493
rect 710 1488 711 1492
rect 715 1488 716 1492
rect 710 1487 716 1488
rect 846 1492 852 1493
rect 846 1488 847 1492
rect 851 1488 852 1492
rect 846 1487 852 1488
rect 974 1492 980 1493
rect 974 1488 975 1492
rect 979 1488 980 1492
rect 974 1487 980 1488
rect 1102 1492 1108 1493
rect 1102 1488 1103 1492
rect 1107 1488 1108 1492
rect 1102 1487 1108 1488
rect 1222 1492 1228 1493
rect 1222 1488 1223 1492
rect 1227 1488 1228 1492
rect 1222 1487 1228 1488
rect 1334 1492 1340 1493
rect 1334 1488 1335 1492
rect 1339 1488 1340 1492
rect 1334 1487 1340 1488
rect 1446 1492 1452 1493
rect 1446 1488 1447 1492
rect 1451 1488 1452 1492
rect 1446 1487 1452 1488
rect 1566 1492 1572 1493
rect 1566 1488 1567 1492
rect 1571 1488 1572 1492
rect 1830 1491 1831 1495
rect 1835 1491 1836 1495
rect 1830 1490 1836 1491
rect 1870 1491 1876 1492
rect 1566 1487 1572 1488
rect 1870 1487 1871 1491
rect 1875 1487 1876 1491
rect 3590 1491 3596 1492
rect 1870 1486 1876 1487
rect 2126 1488 2132 1489
rect 2126 1484 2127 1488
rect 2131 1484 2132 1488
rect 2126 1483 2132 1484
rect 2246 1488 2252 1489
rect 2246 1484 2247 1488
rect 2251 1484 2252 1488
rect 2246 1483 2252 1484
rect 2374 1488 2380 1489
rect 2374 1484 2375 1488
rect 2379 1484 2380 1488
rect 2374 1483 2380 1484
rect 2502 1488 2508 1489
rect 2502 1484 2503 1488
rect 2507 1484 2508 1488
rect 2502 1483 2508 1484
rect 2630 1488 2636 1489
rect 2630 1484 2631 1488
rect 2635 1484 2636 1488
rect 2630 1483 2636 1484
rect 2758 1488 2764 1489
rect 2758 1484 2759 1488
rect 2763 1484 2764 1488
rect 2758 1483 2764 1484
rect 2878 1488 2884 1489
rect 2878 1484 2879 1488
rect 2883 1484 2884 1488
rect 2878 1483 2884 1484
rect 2998 1488 3004 1489
rect 2998 1484 2999 1488
rect 3003 1484 3004 1488
rect 2998 1483 3004 1484
rect 3110 1488 3116 1489
rect 3110 1484 3111 1488
rect 3115 1484 3116 1488
rect 3110 1483 3116 1484
rect 3222 1488 3228 1489
rect 3222 1484 3223 1488
rect 3227 1484 3228 1488
rect 3222 1483 3228 1484
rect 3342 1488 3348 1489
rect 3342 1484 3343 1488
rect 3347 1484 3348 1488
rect 3590 1487 3591 1491
rect 3595 1487 3596 1491
rect 3590 1486 3596 1487
rect 3342 1483 3348 1484
rect 278 1436 284 1437
rect 110 1433 116 1434
rect 110 1429 111 1433
rect 115 1429 116 1433
rect 278 1432 279 1436
rect 283 1432 284 1436
rect 278 1431 284 1432
rect 382 1436 388 1437
rect 382 1432 383 1436
rect 387 1432 388 1436
rect 382 1431 388 1432
rect 510 1436 516 1437
rect 510 1432 511 1436
rect 515 1432 516 1436
rect 510 1431 516 1432
rect 654 1436 660 1437
rect 654 1432 655 1436
rect 659 1432 660 1436
rect 654 1431 660 1432
rect 806 1436 812 1437
rect 806 1432 807 1436
rect 811 1432 812 1436
rect 806 1431 812 1432
rect 958 1436 964 1437
rect 958 1432 959 1436
rect 963 1432 964 1436
rect 958 1431 964 1432
rect 1110 1436 1116 1437
rect 1110 1432 1111 1436
rect 1115 1432 1116 1436
rect 1110 1431 1116 1432
rect 1246 1436 1252 1437
rect 1246 1432 1247 1436
rect 1251 1432 1252 1436
rect 1246 1431 1252 1432
rect 1382 1436 1388 1437
rect 1382 1432 1383 1436
rect 1387 1432 1388 1436
rect 1382 1431 1388 1432
rect 1510 1436 1516 1437
rect 1510 1432 1511 1436
rect 1515 1432 1516 1436
rect 1510 1431 1516 1432
rect 1638 1436 1644 1437
rect 1638 1432 1639 1436
rect 1643 1432 1644 1436
rect 1638 1431 1644 1432
rect 1742 1436 1748 1437
rect 1742 1432 1743 1436
rect 1747 1432 1748 1436
rect 2246 1436 2252 1437
rect 1742 1431 1748 1432
rect 1830 1433 1836 1434
rect 110 1428 116 1429
rect 1830 1429 1831 1433
rect 1835 1429 1836 1433
rect 1830 1428 1836 1429
rect 1870 1433 1876 1434
rect 1870 1429 1871 1433
rect 1875 1429 1876 1433
rect 2246 1432 2247 1436
rect 2251 1432 2252 1436
rect 2246 1431 2252 1432
rect 2342 1436 2348 1437
rect 2342 1432 2343 1436
rect 2347 1432 2348 1436
rect 2342 1431 2348 1432
rect 2454 1436 2460 1437
rect 2454 1432 2455 1436
rect 2459 1432 2460 1436
rect 2454 1431 2460 1432
rect 2574 1436 2580 1437
rect 2574 1432 2575 1436
rect 2579 1432 2580 1436
rect 2574 1431 2580 1432
rect 2702 1436 2708 1437
rect 2702 1432 2703 1436
rect 2707 1432 2708 1436
rect 2702 1431 2708 1432
rect 2830 1436 2836 1437
rect 2830 1432 2831 1436
rect 2835 1432 2836 1436
rect 2830 1431 2836 1432
rect 2950 1436 2956 1437
rect 2950 1432 2951 1436
rect 2955 1432 2956 1436
rect 2950 1431 2956 1432
rect 3070 1436 3076 1437
rect 3070 1432 3071 1436
rect 3075 1432 3076 1436
rect 3070 1431 3076 1432
rect 3182 1436 3188 1437
rect 3182 1432 3183 1436
rect 3187 1432 3188 1436
rect 3182 1431 3188 1432
rect 3294 1436 3300 1437
rect 3294 1432 3295 1436
rect 3299 1432 3300 1436
rect 3294 1431 3300 1432
rect 3406 1436 3412 1437
rect 3406 1432 3407 1436
rect 3411 1432 3412 1436
rect 3406 1431 3412 1432
rect 3502 1436 3508 1437
rect 3502 1432 3503 1436
rect 3507 1432 3508 1436
rect 3502 1431 3508 1432
rect 3590 1433 3596 1434
rect 1870 1428 1876 1429
rect 3590 1429 3591 1433
rect 3595 1429 3596 1433
rect 3590 1428 3596 1429
rect 110 1416 116 1417
rect 110 1412 111 1416
rect 115 1412 116 1416
rect 110 1411 116 1412
rect 1830 1416 1836 1417
rect 1830 1412 1831 1416
rect 1835 1412 1836 1416
rect 1830 1411 1836 1412
rect 1870 1416 1876 1417
rect 1870 1412 1871 1416
rect 1875 1412 1876 1416
rect 1870 1411 1876 1412
rect 3590 1416 3596 1417
rect 3590 1412 3591 1416
rect 3595 1412 3596 1416
rect 3590 1411 3596 1412
rect 286 1398 292 1399
rect 286 1394 287 1398
rect 291 1394 292 1398
rect 286 1393 292 1394
rect 390 1398 396 1399
rect 390 1394 391 1398
rect 395 1394 396 1398
rect 390 1393 396 1394
rect 518 1398 524 1399
rect 518 1394 519 1398
rect 523 1394 524 1398
rect 518 1393 524 1394
rect 662 1398 668 1399
rect 662 1394 663 1398
rect 667 1394 668 1398
rect 662 1393 668 1394
rect 814 1398 820 1399
rect 814 1394 815 1398
rect 819 1394 820 1398
rect 814 1393 820 1394
rect 966 1398 972 1399
rect 966 1394 967 1398
rect 971 1394 972 1398
rect 966 1393 972 1394
rect 1118 1398 1124 1399
rect 1118 1394 1119 1398
rect 1123 1394 1124 1398
rect 1118 1393 1124 1394
rect 1254 1398 1260 1399
rect 1254 1394 1255 1398
rect 1259 1394 1260 1398
rect 1254 1393 1260 1394
rect 1390 1398 1396 1399
rect 1390 1394 1391 1398
rect 1395 1394 1396 1398
rect 1390 1393 1396 1394
rect 1518 1398 1524 1399
rect 1518 1394 1519 1398
rect 1523 1394 1524 1398
rect 1518 1393 1524 1394
rect 1646 1398 1652 1399
rect 1646 1394 1647 1398
rect 1651 1394 1652 1398
rect 1646 1393 1652 1394
rect 1750 1398 1756 1399
rect 1750 1394 1751 1398
rect 1755 1394 1756 1398
rect 1750 1393 1756 1394
rect 2254 1398 2260 1399
rect 2254 1394 2255 1398
rect 2259 1394 2260 1398
rect 2254 1393 2260 1394
rect 2350 1398 2356 1399
rect 2350 1394 2351 1398
rect 2355 1394 2356 1398
rect 2350 1393 2356 1394
rect 2462 1398 2468 1399
rect 2462 1394 2463 1398
rect 2467 1394 2468 1398
rect 2462 1393 2468 1394
rect 2582 1398 2588 1399
rect 2582 1394 2583 1398
rect 2587 1394 2588 1398
rect 2582 1393 2588 1394
rect 2710 1398 2716 1399
rect 2710 1394 2711 1398
rect 2715 1394 2716 1398
rect 2710 1393 2716 1394
rect 2838 1398 2844 1399
rect 2838 1394 2839 1398
rect 2843 1394 2844 1398
rect 2838 1393 2844 1394
rect 2958 1398 2964 1399
rect 2958 1394 2959 1398
rect 2963 1394 2964 1398
rect 2958 1393 2964 1394
rect 3078 1398 3084 1399
rect 3078 1394 3079 1398
rect 3083 1394 3084 1398
rect 3078 1393 3084 1394
rect 3190 1398 3196 1399
rect 3190 1394 3191 1398
rect 3195 1394 3196 1398
rect 3190 1393 3196 1394
rect 3302 1398 3308 1399
rect 3302 1394 3303 1398
rect 3307 1394 3308 1398
rect 3302 1393 3308 1394
rect 3414 1398 3420 1399
rect 3414 1394 3415 1398
rect 3419 1394 3420 1398
rect 3414 1393 3420 1394
rect 3510 1398 3516 1399
rect 3510 1394 3511 1398
rect 3515 1394 3516 1398
rect 3510 1393 3516 1394
rect 2398 1358 2404 1359
rect 2398 1354 2399 1358
rect 2403 1354 2404 1358
rect 2398 1353 2404 1354
rect 2502 1358 2508 1359
rect 2502 1354 2503 1358
rect 2507 1354 2508 1358
rect 2502 1353 2508 1354
rect 2614 1358 2620 1359
rect 2614 1354 2615 1358
rect 2619 1354 2620 1358
rect 2614 1353 2620 1354
rect 2734 1358 2740 1359
rect 2734 1354 2735 1358
rect 2739 1354 2740 1358
rect 2734 1353 2740 1354
rect 2846 1358 2852 1359
rect 2846 1354 2847 1358
rect 2851 1354 2852 1358
rect 2846 1353 2852 1354
rect 2958 1358 2964 1359
rect 2958 1354 2959 1358
rect 2963 1354 2964 1358
rect 2958 1353 2964 1354
rect 3070 1358 3076 1359
rect 3070 1354 3071 1358
rect 3075 1354 3076 1358
rect 3070 1353 3076 1354
rect 3182 1358 3188 1359
rect 3182 1354 3183 1358
rect 3187 1354 3188 1358
rect 3182 1353 3188 1354
rect 3294 1358 3300 1359
rect 3294 1354 3295 1358
rect 3299 1354 3300 1358
rect 3294 1353 3300 1354
rect 3414 1358 3420 1359
rect 3414 1354 3415 1358
rect 3419 1354 3420 1358
rect 3414 1353 3420 1354
rect 222 1350 228 1351
rect 222 1346 223 1350
rect 227 1346 228 1350
rect 222 1345 228 1346
rect 334 1350 340 1351
rect 334 1346 335 1350
rect 339 1346 340 1350
rect 334 1345 340 1346
rect 470 1350 476 1351
rect 470 1346 471 1350
rect 475 1346 476 1350
rect 470 1345 476 1346
rect 622 1350 628 1351
rect 622 1346 623 1350
rect 627 1346 628 1350
rect 622 1345 628 1346
rect 782 1350 788 1351
rect 782 1346 783 1350
rect 787 1346 788 1350
rect 782 1345 788 1346
rect 942 1350 948 1351
rect 942 1346 943 1350
rect 947 1346 948 1350
rect 942 1345 948 1346
rect 1094 1350 1100 1351
rect 1094 1346 1095 1350
rect 1099 1346 1100 1350
rect 1094 1345 1100 1346
rect 1238 1350 1244 1351
rect 1238 1346 1239 1350
rect 1243 1346 1244 1350
rect 1238 1345 1244 1346
rect 1374 1350 1380 1351
rect 1374 1346 1375 1350
rect 1379 1346 1380 1350
rect 1374 1345 1380 1346
rect 1510 1350 1516 1351
rect 1510 1346 1511 1350
rect 1515 1346 1516 1350
rect 1510 1345 1516 1346
rect 1638 1350 1644 1351
rect 1638 1346 1639 1350
rect 1643 1346 1644 1350
rect 1638 1345 1644 1346
rect 1750 1350 1756 1351
rect 1750 1346 1751 1350
rect 1755 1346 1756 1350
rect 1750 1345 1756 1346
rect 1870 1340 1876 1341
rect 1870 1336 1871 1340
rect 1875 1336 1876 1340
rect 1870 1335 1876 1336
rect 3590 1340 3596 1341
rect 3590 1336 3591 1340
rect 3595 1336 3596 1340
rect 3590 1335 3596 1336
rect 110 1332 116 1333
rect 110 1328 111 1332
rect 115 1328 116 1332
rect 110 1327 116 1328
rect 1830 1332 1836 1333
rect 1830 1328 1831 1332
rect 1835 1328 1836 1332
rect 1830 1327 1836 1328
rect 1870 1323 1876 1324
rect 1870 1319 1871 1323
rect 1875 1319 1876 1323
rect 3590 1323 3596 1324
rect 1870 1318 1876 1319
rect 2390 1320 2396 1321
rect 2390 1316 2391 1320
rect 2395 1316 2396 1320
rect 110 1315 116 1316
rect 110 1311 111 1315
rect 115 1311 116 1315
rect 1830 1315 1836 1316
rect 2390 1315 2396 1316
rect 2494 1320 2500 1321
rect 2494 1316 2495 1320
rect 2499 1316 2500 1320
rect 2494 1315 2500 1316
rect 2606 1320 2612 1321
rect 2606 1316 2607 1320
rect 2611 1316 2612 1320
rect 2606 1315 2612 1316
rect 2726 1320 2732 1321
rect 2726 1316 2727 1320
rect 2731 1316 2732 1320
rect 2726 1315 2732 1316
rect 2838 1320 2844 1321
rect 2838 1316 2839 1320
rect 2843 1316 2844 1320
rect 2838 1315 2844 1316
rect 2950 1320 2956 1321
rect 2950 1316 2951 1320
rect 2955 1316 2956 1320
rect 2950 1315 2956 1316
rect 3062 1320 3068 1321
rect 3062 1316 3063 1320
rect 3067 1316 3068 1320
rect 3062 1315 3068 1316
rect 3174 1320 3180 1321
rect 3174 1316 3175 1320
rect 3179 1316 3180 1320
rect 3174 1315 3180 1316
rect 3286 1320 3292 1321
rect 3286 1316 3287 1320
rect 3291 1316 3292 1320
rect 3286 1315 3292 1316
rect 3406 1320 3412 1321
rect 3406 1316 3407 1320
rect 3411 1316 3412 1320
rect 3590 1319 3591 1323
rect 3595 1319 3596 1323
rect 3590 1318 3596 1319
rect 3406 1315 3412 1316
rect 110 1310 116 1311
rect 214 1312 220 1313
rect 214 1308 215 1312
rect 219 1308 220 1312
rect 214 1307 220 1308
rect 326 1312 332 1313
rect 326 1308 327 1312
rect 331 1308 332 1312
rect 326 1307 332 1308
rect 462 1312 468 1313
rect 462 1308 463 1312
rect 467 1308 468 1312
rect 462 1307 468 1308
rect 614 1312 620 1313
rect 614 1308 615 1312
rect 619 1308 620 1312
rect 614 1307 620 1308
rect 774 1312 780 1313
rect 774 1308 775 1312
rect 779 1308 780 1312
rect 774 1307 780 1308
rect 934 1312 940 1313
rect 934 1308 935 1312
rect 939 1308 940 1312
rect 934 1307 940 1308
rect 1086 1312 1092 1313
rect 1086 1308 1087 1312
rect 1091 1308 1092 1312
rect 1086 1307 1092 1308
rect 1230 1312 1236 1313
rect 1230 1308 1231 1312
rect 1235 1308 1236 1312
rect 1230 1307 1236 1308
rect 1366 1312 1372 1313
rect 1366 1308 1367 1312
rect 1371 1308 1372 1312
rect 1366 1307 1372 1308
rect 1502 1312 1508 1313
rect 1502 1308 1503 1312
rect 1507 1308 1508 1312
rect 1502 1307 1508 1308
rect 1630 1312 1636 1313
rect 1630 1308 1631 1312
rect 1635 1308 1636 1312
rect 1630 1307 1636 1308
rect 1742 1312 1748 1313
rect 1742 1308 1743 1312
rect 1747 1308 1748 1312
rect 1830 1311 1831 1315
rect 1835 1311 1836 1315
rect 1830 1310 1836 1311
rect 1742 1307 1748 1308
rect 134 1268 140 1269
rect 110 1265 116 1266
rect 110 1261 111 1265
rect 115 1261 116 1265
rect 134 1264 135 1268
rect 139 1264 140 1268
rect 134 1263 140 1264
rect 214 1268 220 1269
rect 214 1264 215 1268
rect 219 1264 220 1268
rect 214 1263 220 1264
rect 334 1268 340 1269
rect 334 1264 335 1268
rect 339 1264 340 1268
rect 334 1263 340 1264
rect 462 1268 468 1269
rect 462 1264 463 1268
rect 467 1264 468 1268
rect 462 1263 468 1264
rect 606 1268 612 1269
rect 606 1264 607 1268
rect 611 1264 612 1268
rect 606 1263 612 1264
rect 750 1268 756 1269
rect 750 1264 751 1268
rect 755 1264 756 1268
rect 750 1263 756 1264
rect 902 1268 908 1269
rect 902 1264 903 1268
rect 907 1264 908 1268
rect 902 1263 908 1264
rect 1046 1268 1052 1269
rect 1046 1264 1047 1268
rect 1051 1264 1052 1268
rect 1046 1263 1052 1264
rect 1182 1268 1188 1269
rect 1182 1264 1183 1268
rect 1187 1264 1188 1268
rect 1182 1263 1188 1264
rect 1302 1268 1308 1269
rect 1302 1264 1303 1268
rect 1307 1264 1308 1268
rect 1302 1263 1308 1264
rect 1422 1268 1428 1269
rect 1422 1264 1423 1268
rect 1427 1264 1428 1268
rect 1422 1263 1428 1264
rect 1534 1268 1540 1269
rect 1534 1264 1535 1268
rect 1539 1264 1540 1268
rect 1534 1263 1540 1264
rect 1646 1268 1652 1269
rect 1646 1264 1647 1268
rect 1651 1264 1652 1268
rect 1646 1263 1652 1264
rect 1742 1268 1748 1269
rect 1742 1264 1743 1268
rect 1747 1264 1748 1268
rect 1742 1263 1748 1264
rect 1830 1265 1836 1266
rect 110 1260 116 1261
rect 1830 1261 1831 1265
rect 1835 1261 1836 1265
rect 1830 1260 1836 1261
rect 1894 1260 1900 1261
rect 1870 1257 1876 1258
rect 1870 1253 1871 1257
rect 1875 1253 1876 1257
rect 1894 1256 1895 1260
rect 1899 1256 1900 1260
rect 1894 1255 1900 1256
rect 2070 1260 2076 1261
rect 2070 1256 2071 1260
rect 2075 1256 2076 1260
rect 2070 1255 2076 1256
rect 2254 1260 2260 1261
rect 2254 1256 2255 1260
rect 2259 1256 2260 1260
rect 2254 1255 2260 1256
rect 2422 1260 2428 1261
rect 2422 1256 2423 1260
rect 2427 1256 2428 1260
rect 2422 1255 2428 1256
rect 2582 1260 2588 1261
rect 2582 1256 2583 1260
rect 2587 1256 2588 1260
rect 2582 1255 2588 1256
rect 2734 1260 2740 1261
rect 2734 1256 2735 1260
rect 2739 1256 2740 1260
rect 2734 1255 2740 1256
rect 2878 1260 2884 1261
rect 2878 1256 2879 1260
rect 2883 1256 2884 1260
rect 2878 1255 2884 1256
rect 3014 1260 3020 1261
rect 3014 1256 3015 1260
rect 3019 1256 3020 1260
rect 3014 1255 3020 1256
rect 3142 1260 3148 1261
rect 3142 1256 3143 1260
rect 3147 1256 3148 1260
rect 3142 1255 3148 1256
rect 3270 1260 3276 1261
rect 3270 1256 3271 1260
rect 3275 1256 3276 1260
rect 3270 1255 3276 1256
rect 3398 1260 3404 1261
rect 3398 1256 3399 1260
rect 3403 1256 3404 1260
rect 3398 1255 3404 1256
rect 3502 1260 3508 1261
rect 3502 1256 3503 1260
rect 3507 1256 3508 1260
rect 3502 1255 3508 1256
rect 3590 1257 3596 1258
rect 1870 1252 1876 1253
rect 3590 1253 3591 1257
rect 3595 1253 3596 1257
rect 3590 1252 3596 1253
rect 110 1248 116 1249
rect 110 1244 111 1248
rect 115 1244 116 1248
rect 110 1243 116 1244
rect 1830 1248 1836 1249
rect 1830 1244 1831 1248
rect 1835 1244 1836 1248
rect 1830 1243 1836 1244
rect 1870 1240 1876 1241
rect 1870 1236 1871 1240
rect 1875 1236 1876 1240
rect 1870 1235 1876 1236
rect 3590 1240 3596 1241
rect 3590 1236 3591 1240
rect 3595 1236 3596 1240
rect 3590 1235 3596 1236
rect 142 1230 148 1231
rect 142 1226 143 1230
rect 147 1226 148 1230
rect 142 1225 148 1226
rect 222 1230 228 1231
rect 222 1226 223 1230
rect 227 1226 228 1230
rect 222 1225 228 1226
rect 342 1230 348 1231
rect 342 1226 343 1230
rect 347 1226 348 1230
rect 342 1225 348 1226
rect 470 1230 476 1231
rect 470 1226 471 1230
rect 475 1226 476 1230
rect 470 1225 476 1226
rect 614 1230 620 1231
rect 614 1226 615 1230
rect 619 1226 620 1230
rect 614 1225 620 1226
rect 758 1230 764 1231
rect 758 1226 759 1230
rect 763 1226 764 1230
rect 758 1225 764 1226
rect 910 1230 916 1231
rect 910 1226 911 1230
rect 915 1226 916 1230
rect 910 1225 916 1226
rect 1054 1230 1060 1231
rect 1054 1226 1055 1230
rect 1059 1226 1060 1230
rect 1054 1225 1060 1226
rect 1190 1230 1196 1231
rect 1190 1226 1191 1230
rect 1195 1226 1196 1230
rect 1190 1225 1196 1226
rect 1310 1230 1316 1231
rect 1310 1226 1311 1230
rect 1315 1226 1316 1230
rect 1310 1225 1316 1226
rect 1430 1230 1436 1231
rect 1430 1226 1431 1230
rect 1435 1226 1436 1230
rect 1430 1225 1436 1226
rect 1542 1230 1548 1231
rect 1542 1226 1543 1230
rect 1547 1226 1548 1230
rect 1542 1225 1548 1226
rect 1654 1230 1660 1231
rect 1654 1226 1655 1230
rect 1659 1226 1660 1230
rect 1654 1225 1660 1226
rect 1750 1230 1756 1231
rect 1750 1226 1751 1230
rect 1755 1226 1756 1230
rect 1750 1225 1756 1226
rect 1902 1222 1908 1223
rect 1902 1218 1903 1222
rect 1907 1218 1908 1222
rect 1902 1217 1908 1218
rect 2078 1222 2084 1223
rect 2078 1218 2079 1222
rect 2083 1218 2084 1222
rect 2078 1217 2084 1218
rect 2262 1222 2268 1223
rect 2262 1218 2263 1222
rect 2267 1218 2268 1222
rect 2262 1217 2268 1218
rect 2430 1222 2436 1223
rect 2430 1218 2431 1222
rect 2435 1218 2436 1222
rect 2430 1217 2436 1218
rect 2590 1222 2596 1223
rect 2590 1218 2591 1222
rect 2595 1218 2596 1222
rect 2590 1217 2596 1218
rect 2742 1222 2748 1223
rect 2742 1218 2743 1222
rect 2747 1218 2748 1222
rect 2742 1217 2748 1218
rect 2886 1222 2892 1223
rect 2886 1218 2887 1222
rect 2891 1218 2892 1222
rect 2886 1217 2892 1218
rect 3022 1222 3028 1223
rect 3022 1218 3023 1222
rect 3027 1218 3028 1222
rect 3022 1217 3028 1218
rect 3150 1222 3156 1223
rect 3150 1218 3151 1222
rect 3155 1218 3156 1222
rect 3150 1217 3156 1218
rect 3278 1222 3284 1223
rect 3278 1218 3279 1222
rect 3283 1218 3284 1222
rect 3278 1217 3284 1218
rect 3406 1222 3412 1223
rect 3406 1218 3407 1222
rect 3411 1218 3412 1222
rect 3406 1217 3412 1218
rect 3510 1222 3516 1223
rect 3510 1218 3511 1222
rect 3515 1218 3516 1222
rect 3510 1217 3516 1218
rect 142 1186 148 1187
rect 142 1182 143 1186
rect 147 1182 148 1186
rect 142 1181 148 1182
rect 254 1186 260 1187
rect 254 1182 255 1186
rect 259 1182 260 1186
rect 254 1181 260 1182
rect 382 1186 388 1187
rect 382 1182 383 1186
rect 387 1182 388 1186
rect 382 1181 388 1182
rect 502 1186 508 1187
rect 502 1182 503 1186
rect 507 1182 508 1186
rect 502 1181 508 1182
rect 614 1186 620 1187
rect 614 1182 615 1186
rect 619 1182 620 1186
rect 614 1181 620 1182
rect 718 1186 724 1187
rect 718 1182 719 1186
rect 723 1182 724 1186
rect 718 1181 724 1182
rect 814 1186 820 1187
rect 814 1182 815 1186
rect 819 1182 820 1186
rect 814 1181 820 1182
rect 910 1186 916 1187
rect 910 1182 911 1186
rect 915 1182 916 1186
rect 910 1181 916 1182
rect 998 1186 1004 1187
rect 998 1182 999 1186
rect 1003 1182 1004 1186
rect 998 1181 1004 1182
rect 1094 1186 1100 1187
rect 1094 1182 1095 1186
rect 1099 1182 1100 1186
rect 1094 1181 1100 1182
rect 1190 1186 1196 1187
rect 1190 1182 1191 1186
rect 1195 1182 1196 1186
rect 1190 1181 1196 1182
rect 1286 1186 1292 1187
rect 1286 1182 1287 1186
rect 1291 1182 1292 1186
rect 1286 1181 1292 1182
rect 1902 1182 1908 1183
rect 1902 1178 1903 1182
rect 1907 1178 1908 1182
rect 1902 1177 1908 1178
rect 1990 1182 1996 1183
rect 1990 1178 1991 1182
rect 1995 1178 1996 1182
rect 1990 1177 1996 1178
rect 2102 1182 2108 1183
rect 2102 1178 2103 1182
rect 2107 1178 2108 1182
rect 2102 1177 2108 1178
rect 2214 1182 2220 1183
rect 2214 1178 2215 1182
rect 2219 1178 2220 1182
rect 2214 1177 2220 1178
rect 2326 1182 2332 1183
rect 2326 1178 2327 1182
rect 2331 1178 2332 1182
rect 2326 1177 2332 1178
rect 2446 1182 2452 1183
rect 2446 1178 2447 1182
rect 2451 1178 2452 1182
rect 2446 1177 2452 1178
rect 2574 1182 2580 1183
rect 2574 1178 2575 1182
rect 2579 1178 2580 1182
rect 2574 1177 2580 1178
rect 2718 1182 2724 1183
rect 2718 1178 2719 1182
rect 2723 1178 2724 1182
rect 2718 1177 2724 1178
rect 2870 1182 2876 1183
rect 2870 1178 2871 1182
rect 2875 1178 2876 1182
rect 2870 1177 2876 1178
rect 3030 1182 3036 1183
rect 3030 1178 3031 1182
rect 3035 1178 3036 1182
rect 3030 1177 3036 1178
rect 3190 1182 3196 1183
rect 3190 1178 3191 1182
rect 3195 1178 3196 1182
rect 3190 1177 3196 1178
rect 3358 1182 3364 1183
rect 3358 1178 3359 1182
rect 3363 1178 3364 1182
rect 3358 1177 3364 1178
rect 3510 1182 3516 1183
rect 3510 1178 3511 1182
rect 3515 1178 3516 1182
rect 3510 1177 3516 1178
rect 110 1168 116 1169
rect 110 1164 111 1168
rect 115 1164 116 1168
rect 110 1163 116 1164
rect 1830 1168 1836 1169
rect 1830 1164 1831 1168
rect 1835 1164 1836 1168
rect 1830 1163 1836 1164
rect 1870 1164 1876 1165
rect 1870 1160 1871 1164
rect 1875 1160 1876 1164
rect 1870 1159 1876 1160
rect 3590 1164 3596 1165
rect 3590 1160 3591 1164
rect 3595 1160 3596 1164
rect 3590 1159 3596 1160
rect 110 1151 116 1152
rect 110 1147 111 1151
rect 115 1147 116 1151
rect 1830 1151 1836 1152
rect 110 1146 116 1147
rect 134 1148 140 1149
rect 134 1144 135 1148
rect 139 1144 140 1148
rect 134 1143 140 1144
rect 246 1148 252 1149
rect 246 1144 247 1148
rect 251 1144 252 1148
rect 246 1143 252 1144
rect 374 1148 380 1149
rect 374 1144 375 1148
rect 379 1144 380 1148
rect 374 1143 380 1144
rect 494 1148 500 1149
rect 494 1144 495 1148
rect 499 1144 500 1148
rect 494 1143 500 1144
rect 606 1148 612 1149
rect 606 1144 607 1148
rect 611 1144 612 1148
rect 606 1143 612 1144
rect 710 1148 716 1149
rect 710 1144 711 1148
rect 715 1144 716 1148
rect 710 1143 716 1144
rect 806 1148 812 1149
rect 806 1144 807 1148
rect 811 1144 812 1148
rect 806 1143 812 1144
rect 902 1148 908 1149
rect 902 1144 903 1148
rect 907 1144 908 1148
rect 902 1143 908 1144
rect 990 1148 996 1149
rect 990 1144 991 1148
rect 995 1144 996 1148
rect 990 1143 996 1144
rect 1086 1148 1092 1149
rect 1086 1144 1087 1148
rect 1091 1144 1092 1148
rect 1086 1143 1092 1144
rect 1182 1148 1188 1149
rect 1182 1144 1183 1148
rect 1187 1144 1188 1148
rect 1182 1143 1188 1144
rect 1278 1148 1284 1149
rect 1278 1144 1279 1148
rect 1283 1144 1284 1148
rect 1830 1147 1831 1151
rect 1835 1147 1836 1151
rect 1830 1146 1836 1147
rect 1870 1147 1876 1148
rect 1278 1143 1284 1144
rect 1870 1143 1871 1147
rect 1875 1143 1876 1147
rect 3590 1147 3596 1148
rect 1870 1142 1876 1143
rect 1894 1144 1900 1145
rect 1894 1140 1895 1144
rect 1899 1140 1900 1144
rect 1894 1139 1900 1140
rect 1982 1144 1988 1145
rect 1982 1140 1983 1144
rect 1987 1140 1988 1144
rect 1982 1139 1988 1140
rect 2094 1144 2100 1145
rect 2094 1140 2095 1144
rect 2099 1140 2100 1144
rect 2094 1139 2100 1140
rect 2206 1144 2212 1145
rect 2206 1140 2207 1144
rect 2211 1140 2212 1144
rect 2206 1139 2212 1140
rect 2318 1144 2324 1145
rect 2318 1140 2319 1144
rect 2323 1140 2324 1144
rect 2318 1139 2324 1140
rect 2438 1144 2444 1145
rect 2438 1140 2439 1144
rect 2443 1140 2444 1144
rect 2438 1139 2444 1140
rect 2566 1144 2572 1145
rect 2566 1140 2567 1144
rect 2571 1140 2572 1144
rect 2566 1139 2572 1140
rect 2710 1144 2716 1145
rect 2710 1140 2711 1144
rect 2715 1140 2716 1144
rect 2710 1139 2716 1140
rect 2862 1144 2868 1145
rect 2862 1140 2863 1144
rect 2867 1140 2868 1144
rect 2862 1139 2868 1140
rect 3022 1144 3028 1145
rect 3022 1140 3023 1144
rect 3027 1140 3028 1144
rect 3022 1139 3028 1140
rect 3182 1144 3188 1145
rect 3182 1140 3183 1144
rect 3187 1140 3188 1144
rect 3182 1139 3188 1140
rect 3350 1144 3356 1145
rect 3350 1140 3351 1144
rect 3355 1140 3356 1144
rect 3350 1139 3356 1140
rect 3502 1144 3508 1145
rect 3502 1140 3503 1144
rect 3507 1140 3508 1144
rect 3590 1143 3591 1147
rect 3595 1143 3596 1147
rect 3590 1142 3596 1143
rect 3502 1139 3508 1140
rect 134 1092 140 1093
rect 110 1089 116 1090
rect 110 1085 111 1089
rect 115 1085 116 1089
rect 134 1088 135 1092
rect 139 1088 140 1092
rect 134 1087 140 1088
rect 254 1092 260 1093
rect 254 1088 255 1092
rect 259 1088 260 1092
rect 254 1087 260 1088
rect 398 1092 404 1093
rect 398 1088 399 1092
rect 403 1088 404 1092
rect 398 1087 404 1088
rect 534 1092 540 1093
rect 534 1088 535 1092
rect 539 1088 540 1092
rect 534 1087 540 1088
rect 662 1092 668 1093
rect 662 1088 663 1092
rect 667 1088 668 1092
rect 662 1087 668 1088
rect 782 1092 788 1093
rect 782 1088 783 1092
rect 787 1088 788 1092
rect 782 1087 788 1088
rect 894 1092 900 1093
rect 894 1088 895 1092
rect 899 1088 900 1092
rect 894 1087 900 1088
rect 998 1092 1004 1093
rect 998 1088 999 1092
rect 1003 1088 1004 1092
rect 998 1087 1004 1088
rect 1094 1092 1100 1093
rect 1094 1088 1095 1092
rect 1099 1088 1100 1092
rect 1094 1087 1100 1088
rect 1190 1092 1196 1093
rect 1190 1088 1191 1092
rect 1195 1088 1196 1092
rect 1190 1087 1196 1088
rect 1294 1092 1300 1093
rect 1294 1088 1295 1092
rect 1299 1088 1300 1092
rect 1294 1087 1300 1088
rect 1398 1092 1404 1093
rect 1398 1088 1399 1092
rect 1403 1088 1404 1092
rect 1966 1092 1972 1093
rect 1398 1087 1404 1088
rect 1830 1089 1836 1090
rect 110 1084 116 1085
rect 1830 1085 1831 1089
rect 1835 1085 1836 1089
rect 1830 1084 1836 1085
rect 1870 1089 1876 1090
rect 1870 1085 1871 1089
rect 1875 1085 1876 1089
rect 1966 1088 1967 1092
rect 1971 1088 1972 1092
rect 1966 1087 1972 1088
rect 2046 1092 2052 1093
rect 2046 1088 2047 1092
rect 2051 1088 2052 1092
rect 2046 1087 2052 1088
rect 2134 1092 2140 1093
rect 2134 1088 2135 1092
rect 2139 1088 2140 1092
rect 2134 1087 2140 1088
rect 2230 1092 2236 1093
rect 2230 1088 2231 1092
rect 2235 1088 2236 1092
rect 2230 1087 2236 1088
rect 2334 1092 2340 1093
rect 2334 1088 2335 1092
rect 2339 1088 2340 1092
rect 2334 1087 2340 1088
rect 2438 1092 2444 1093
rect 2438 1088 2439 1092
rect 2443 1088 2444 1092
rect 2438 1087 2444 1088
rect 2550 1092 2556 1093
rect 2550 1088 2551 1092
rect 2555 1088 2556 1092
rect 2550 1087 2556 1088
rect 2678 1092 2684 1093
rect 2678 1088 2679 1092
rect 2683 1088 2684 1092
rect 2678 1087 2684 1088
rect 2822 1092 2828 1093
rect 2822 1088 2823 1092
rect 2827 1088 2828 1092
rect 2822 1087 2828 1088
rect 2982 1092 2988 1093
rect 2982 1088 2983 1092
rect 2987 1088 2988 1092
rect 2982 1087 2988 1088
rect 3158 1092 3164 1093
rect 3158 1088 3159 1092
rect 3163 1088 3164 1092
rect 3158 1087 3164 1088
rect 3342 1092 3348 1093
rect 3342 1088 3343 1092
rect 3347 1088 3348 1092
rect 3342 1087 3348 1088
rect 3502 1092 3508 1093
rect 3502 1088 3503 1092
rect 3507 1088 3508 1092
rect 3502 1087 3508 1088
rect 3590 1089 3596 1090
rect 1870 1084 1876 1085
rect 3590 1085 3591 1089
rect 3595 1085 3596 1089
rect 3590 1084 3596 1085
rect 110 1072 116 1073
rect 110 1068 111 1072
rect 115 1068 116 1072
rect 110 1067 116 1068
rect 1830 1072 1836 1073
rect 1830 1068 1831 1072
rect 1835 1068 1836 1072
rect 1830 1067 1836 1068
rect 1870 1072 1876 1073
rect 1870 1068 1871 1072
rect 1875 1068 1876 1072
rect 1870 1067 1876 1068
rect 3590 1072 3596 1073
rect 3590 1068 3591 1072
rect 3595 1068 3596 1072
rect 3590 1067 3596 1068
rect 142 1054 148 1055
rect 142 1050 143 1054
rect 147 1050 148 1054
rect 142 1049 148 1050
rect 262 1054 268 1055
rect 262 1050 263 1054
rect 267 1050 268 1054
rect 262 1049 268 1050
rect 406 1054 412 1055
rect 406 1050 407 1054
rect 411 1050 412 1054
rect 406 1049 412 1050
rect 542 1054 548 1055
rect 542 1050 543 1054
rect 547 1050 548 1054
rect 542 1049 548 1050
rect 670 1054 676 1055
rect 670 1050 671 1054
rect 675 1050 676 1054
rect 670 1049 676 1050
rect 790 1054 796 1055
rect 790 1050 791 1054
rect 795 1050 796 1054
rect 790 1049 796 1050
rect 902 1054 908 1055
rect 902 1050 903 1054
rect 907 1050 908 1054
rect 902 1049 908 1050
rect 1006 1054 1012 1055
rect 1006 1050 1007 1054
rect 1011 1050 1012 1054
rect 1006 1049 1012 1050
rect 1102 1054 1108 1055
rect 1102 1050 1103 1054
rect 1107 1050 1108 1054
rect 1102 1049 1108 1050
rect 1198 1054 1204 1055
rect 1198 1050 1199 1054
rect 1203 1050 1204 1054
rect 1198 1049 1204 1050
rect 1302 1054 1308 1055
rect 1302 1050 1303 1054
rect 1307 1050 1308 1054
rect 1302 1049 1308 1050
rect 1406 1054 1412 1055
rect 1406 1050 1407 1054
rect 1411 1050 1412 1054
rect 1406 1049 1412 1050
rect 1974 1054 1980 1055
rect 1974 1050 1975 1054
rect 1979 1050 1980 1054
rect 1974 1049 1980 1050
rect 2054 1054 2060 1055
rect 2054 1050 2055 1054
rect 2059 1050 2060 1054
rect 2054 1049 2060 1050
rect 2142 1054 2148 1055
rect 2142 1050 2143 1054
rect 2147 1050 2148 1054
rect 2142 1049 2148 1050
rect 2238 1054 2244 1055
rect 2238 1050 2239 1054
rect 2243 1050 2244 1054
rect 2238 1049 2244 1050
rect 2342 1054 2348 1055
rect 2342 1050 2343 1054
rect 2347 1050 2348 1054
rect 2342 1049 2348 1050
rect 2446 1054 2452 1055
rect 2446 1050 2447 1054
rect 2451 1050 2452 1054
rect 2446 1049 2452 1050
rect 2558 1054 2564 1055
rect 2558 1050 2559 1054
rect 2563 1050 2564 1054
rect 2558 1049 2564 1050
rect 2686 1054 2692 1055
rect 2686 1050 2687 1054
rect 2691 1050 2692 1054
rect 2686 1049 2692 1050
rect 2830 1054 2836 1055
rect 2830 1050 2831 1054
rect 2835 1050 2836 1054
rect 2830 1049 2836 1050
rect 2990 1054 2996 1055
rect 2990 1050 2991 1054
rect 2995 1050 2996 1054
rect 2990 1049 2996 1050
rect 3166 1054 3172 1055
rect 3166 1050 3167 1054
rect 3171 1050 3172 1054
rect 3166 1049 3172 1050
rect 3350 1054 3356 1055
rect 3350 1050 3351 1054
rect 3355 1050 3356 1054
rect 3350 1049 3356 1050
rect 3510 1054 3516 1055
rect 3510 1050 3511 1054
rect 3515 1050 3516 1054
rect 3510 1049 3516 1050
rect 142 1014 148 1015
rect 142 1010 143 1014
rect 147 1010 148 1014
rect 142 1009 148 1010
rect 270 1014 276 1015
rect 270 1010 271 1014
rect 275 1010 276 1014
rect 270 1009 276 1010
rect 422 1014 428 1015
rect 422 1010 423 1014
rect 427 1010 428 1014
rect 422 1009 428 1010
rect 582 1014 588 1015
rect 582 1010 583 1014
rect 587 1010 588 1014
rect 582 1009 588 1010
rect 734 1014 740 1015
rect 734 1010 735 1014
rect 739 1010 740 1014
rect 734 1009 740 1010
rect 886 1014 892 1015
rect 886 1010 887 1014
rect 891 1010 892 1014
rect 886 1009 892 1010
rect 1030 1014 1036 1015
rect 1030 1010 1031 1014
rect 1035 1010 1036 1014
rect 1030 1009 1036 1010
rect 1158 1014 1164 1015
rect 1158 1010 1159 1014
rect 1163 1010 1164 1014
rect 1158 1009 1164 1010
rect 1278 1014 1284 1015
rect 1278 1010 1279 1014
rect 1283 1010 1284 1014
rect 1278 1009 1284 1010
rect 1398 1014 1404 1015
rect 1398 1010 1399 1014
rect 1403 1010 1404 1014
rect 1398 1009 1404 1010
rect 1518 1014 1524 1015
rect 1518 1010 1519 1014
rect 1523 1010 1524 1014
rect 1518 1009 1524 1010
rect 1638 1014 1644 1015
rect 1638 1010 1639 1014
rect 1643 1010 1644 1014
rect 1638 1009 1644 1010
rect 2030 1014 2036 1015
rect 2030 1010 2031 1014
rect 2035 1010 2036 1014
rect 2030 1009 2036 1010
rect 2126 1014 2132 1015
rect 2126 1010 2127 1014
rect 2131 1010 2132 1014
rect 2126 1009 2132 1010
rect 2230 1014 2236 1015
rect 2230 1010 2231 1014
rect 2235 1010 2236 1014
rect 2230 1009 2236 1010
rect 2350 1014 2356 1015
rect 2350 1010 2351 1014
rect 2355 1010 2356 1014
rect 2350 1009 2356 1010
rect 2470 1014 2476 1015
rect 2470 1010 2471 1014
rect 2475 1010 2476 1014
rect 2470 1009 2476 1010
rect 2598 1014 2604 1015
rect 2598 1010 2599 1014
rect 2603 1010 2604 1014
rect 2598 1009 2604 1010
rect 2726 1014 2732 1015
rect 2726 1010 2727 1014
rect 2731 1010 2732 1014
rect 2726 1009 2732 1010
rect 2854 1014 2860 1015
rect 2854 1010 2855 1014
rect 2859 1010 2860 1014
rect 2854 1009 2860 1010
rect 2982 1014 2988 1015
rect 2982 1010 2983 1014
rect 2987 1010 2988 1014
rect 2982 1009 2988 1010
rect 3110 1014 3116 1015
rect 3110 1010 3111 1014
rect 3115 1010 3116 1014
rect 3110 1009 3116 1010
rect 3246 1014 3252 1015
rect 3246 1010 3247 1014
rect 3251 1010 3252 1014
rect 3246 1009 3252 1010
rect 3390 1014 3396 1015
rect 3390 1010 3391 1014
rect 3395 1010 3396 1014
rect 3390 1009 3396 1010
rect 3510 1014 3516 1015
rect 3510 1010 3511 1014
rect 3515 1010 3516 1014
rect 3510 1009 3516 1010
rect 110 996 116 997
rect 110 992 111 996
rect 115 992 116 996
rect 110 991 116 992
rect 1830 996 1836 997
rect 1830 992 1831 996
rect 1835 992 1836 996
rect 1830 991 1836 992
rect 1870 996 1876 997
rect 1870 992 1871 996
rect 1875 992 1876 996
rect 1870 991 1876 992
rect 3590 996 3596 997
rect 3590 992 3591 996
rect 3595 992 3596 996
rect 3590 991 3596 992
rect 110 979 116 980
rect 110 975 111 979
rect 115 975 116 979
rect 1830 979 1836 980
rect 110 974 116 975
rect 134 976 140 977
rect 134 972 135 976
rect 139 972 140 976
rect 134 971 140 972
rect 262 976 268 977
rect 262 972 263 976
rect 267 972 268 976
rect 262 971 268 972
rect 414 976 420 977
rect 414 972 415 976
rect 419 972 420 976
rect 414 971 420 972
rect 574 976 580 977
rect 574 972 575 976
rect 579 972 580 976
rect 574 971 580 972
rect 726 976 732 977
rect 726 972 727 976
rect 731 972 732 976
rect 726 971 732 972
rect 878 976 884 977
rect 878 972 879 976
rect 883 972 884 976
rect 878 971 884 972
rect 1022 976 1028 977
rect 1022 972 1023 976
rect 1027 972 1028 976
rect 1022 971 1028 972
rect 1150 976 1156 977
rect 1150 972 1151 976
rect 1155 972 1156 976
rect 1150 971 1156 972
rect 1270 976 1276 977
rect 1270 972 1271 976
rect 1275 972 1276 976
rect 1270 971 1276 972
rect 1390 976 1396 977
rect 1390 972 1391 976
rect 1395 972 1396 976
rect 1390 971 1396 972
rect 1510 976 1516 977
rect 1510 972 1511 976
rect 1515 972 1516 976
rect 1510 971 1516 972
rect 1630 976 1636 977
rect 1630 972 1631 976
rect 1635 972 1636 976
rect 1830 975 1831 979
rect 1835 975 1836 979
rect 1830 974 1836 975
rect 1870 979 1876 980
rect 1870 975 1871 979
rect 1875 975 1876 979
rect 3590 979 3596 980
rect 1870 974 1876 975
rect 2022 976 2028 977
rect 1630 971 1636 972
rect 2022 972 2023 976
rect 2027 972 2028 976
rect 2022 971 2028 972
rect 2118 976 2124 977
rect 2118 972 2119 976
rect 2123 972 2124 976
rect 2118 971 2124 972
rect 2222 976 2228 977
rect 2222 972 2223 976
rect 2227 972 2228 976
rect 2222 971 2228 972
rect 2342 976 2348 977
rect 2342 972 2343 976
rect 2347 972 2348 976
rect 2342 971 2348 972
rect 2462 976 2468 977
rect 2462 972 2463 976
rect 2467 972 2468 976
rect 2462 971 2468 972
rect 2590 976 2596 977
rect 2590 972 2591 976
rect 2595 972 2596 976
rect 2590 971 2596 972
rect 2718 976 2724 977
rect 2718 972 2719 976
rect 2723 972 2724 976
rect 2718 971 2724 972
rect 2846 976 2852 977
rect 2846 972 2847 976
rect 2851 972 2852 976
rect 2846 971 2852 972
rect 2974 976 2980 977
rect 2974 972 2975 976
rect 2979 972 2980 976
rect 2974 971 2980 972
rect 3102 976 3108 977
rect 3102 972 3103 976
rect 3107 972 3108 976
rect 3102 971 3108 972
rect 3238 976 3244 977
rect 3238 972 3239 976
rect 3243 972 3244 976
rect 3238 971 3244 972
rect 3382 976 3388 977
rect 3382 972 3383 976
rect 3387 972 3388 976
rect 3382 971 3388 972
rect 3502 976 3508 977
rect 3502 972 3503 976
rect 3507 972 3508 976
rect 3590 975 3591 979
rect 3595 975 3596 979
rect 3590 974 3596 975
rect 3502 971 3508 972
rect 134 924 140 925
rect 110 921 116 922
rect 110 917 111 921
rect 115 917 116 921
rect 134 920 135 924
rect 139 920 140 924
rect 134 919 140 920
rect 214 924 220 925
rect 214 920 215 924
rect 219 920 220 924
rect 214 919 220 920
rect 334 924 340 925
rect 334 920 335 924
rect 339 920 340 924
rect 334 919 340 920
rect 462 924 468 925
rect 462 920 463 924
rect 467 920 468 924
rect 462 919 468 920
rect 598 924 604 925
rect 598 920 599 924
rect 603 920 604 924
rect 598 919 604 920
rect 734 924 740 925
rect 734 920 735 924
rect 739 920 740 924
rect 734 919 740 920
rect 862 924 868 925
rect 862 920 863 924
rect 867 920 868 924
rect 862 919 868 920
rect 990 924 996 925
rect 990 920 991 924
rect 995 920 996 924
rect 990 919 996 920
rect 1110 924 1116 925
rect 1110 920 1111 924
rect 1115 920 1116 924
rect 1110 919 1116 920
rect 1222 924 1228 925
rect 1222 920 1223 924
rect 1227 920 1228 924
rect 1222 919 1228 920
rect 1334 924 1340 925
rect 1334 920 1335 924
rect 1339 920 1340 924
rect 1334 919 1340 920
rect 1454 924 1460 925
rect 1454 920 1455 924
rect 1459 920 1460 924
rect 1894 924 1900 925
rect 1454 919 1460 920
rect 1830 921 1836 922
rect 110 916 116 917
rect 1830 917 1831 921
rect 1835 917 1836 921
rect 1830 916 1836 917
rect 1870 921 1876 922
rect 1870 917 1871 921
rect 1875 917 1876 921
rect 1894 920 1895 924
rect 1899 920 1900 924
rect 1894 919 1900 920
rect 1982 924 1988 925
rect 1982 920 1983 924
rect 1987 920 1988 924
rect 1982 919 1988 920
rect 2110 924 2116 925
rect 2110 920 2111 924
rect 2115 920 2116 924
rect 2110 919 2116 920
rect 2262 924 2268 925
rect 2262 920 2263 924
rect 2267 920 2268 924
rect 2262 919 2268 920
rect 2422 924 2428 925
rect 2422 920 2423 924
rect 2427 920 2428 924
rect 2422 919 2428 920
rect 2582 924 2588 925
rect 2582 920 2583 924
rect 2587 920 2588 924
rect 2582 919 2588 920
rect 2734 924 2740 925
rect 2734 920 2735 924
rect 2739 920 2740 924
rect 2734 919 2740 920
rect 2878 924 2884 925
rect 2878 920 2879 924
rect 2883 920 2884 924
rect 2878 919 2884 920
rect 3014 924 3020 925
rect 3014 920 3015 924
rect 3019 920 3020 924
rect 3014 919 3020 920
rect 3142 924 3148 925
rect 3142 920 3143 924
rect 3147 920 3148 924
rect 3142 919 3148 920
rect 3270 924 3276 925
rect 3270 920 3271 924
rect 3275 920 3276 924
rect 3270 919 3276 920
rect 3398 924 3404 925
rect 3398 920 3399 924
rect 3403 920 3404 924
rect 3398 919 3404 920
rect 3502 924 3508 925
rect 3502 920 3503 924
rect 3507 920 3508 924
rect 3502 919 3508 920
rect 3590 921 3596 922
rect 1870 916 1876 917
rect 3590 917 3591 921
rect 3595 917 3596 921
rect 3590 916 3596 917
rect 110 904 116 905
rect 110 900 111 904
rect 115 900 116 904
rect 110 899 116 900
rect 1830 904 1836 905
rect 1830 900 1831 904
rect 1835 900 1836 904
rect 1830 899 1836 900
rect 1870 904 1876 905
rect 1870 900 1871 904
rect 1875 900 1876 904
rect 1870 899 1876 900
rect 3590 904 3596 905
rect 3590 900 3591 904
rect 3595 900 3596 904
rect 3590 899 3596 900
rect 142 886 148 887
rect 142 882 143 886
rect 147 882 148 886
rect 142 881 148 882
rect 222 886 228 887
rect 222 882 223 886
rect 227 882 228 886
rect 222 881 228 882
rect 342 886 348 887
rect 342 882 343 886
rect 347 882 348 886
rect 342 881 348 882
rect 470 886 476 887
rect 470 882 471 886
rect 475 882 476 886
rect 470 881 476 882
rect 606 886 612 887
rect 606 882 607 886
rect 611 882 612 886
rect 606 881 612 882
rect 742 886 748 887
rect 742 882 743 886
rect 747 882 748 886
rect 742 881 748 882
rect 870 886 876 887
rect 870 882 871 886
rect 875 882 876 886
rect 870 881 876 882
rect 998 886 1004 887
rect 998 882 999 886
rect 1003 882 1004 886
rect 998 881 1004 882
rect 1118 886 1124 887
rect 1118 882 1119 886
rect 1123 882 1124 886
rect 1118 881 1124 882
rect 1230 886 1236 887
rect 1230 882 1231 886
rect 1235 882 1236 886
rect 1230 881 1236 882
rect 1342 886 1348 887
rect 1342 882 1343 886
rect 1347 882 1348 886
rect 1342 881 1348 882
rect 1462 886 1468 887
rect 1462 882 1463 886
rect 1467 882 1468 886
rect 1462 881 1468 882
rect 1902 886 1908 887
rect 1902 882 1903 886
rect 1907 882 1908 886
rect 1902 881 1908 882
rect 1990 886 1996 887
rect 1990 882 1991 886
rect 1995 882 1996 886
rect 1990 881 1996 882
rect 2118 886 2124 887
rect 2118 882 2119 886
rect 2123 882 2124 886
rect 2118 881 2124 882
rect 2270 886 2276 887
rect 2270 882 2271 886
rect 2275 882 2276 886
rect 2270 881 2276 882
rect 2430 886 2436 887
rect 2430 882 2431 886
rect 2435 882 2436 886
rect 2430 881 2436 882
rect 2590 886 2596 887
rect 2590 882 2591 886
rect 2595 882 2596 886
rect 2590 881 2596 882
rect 2742 886 2748 887
rect 2742 882 2743 886
rect 2747 882 2748 886
rect 2742 881 2748 882
rect 2886 886 2892 887
rect 2886 882 2887 886
rect 2891 882 2892 886
rect 2886 881 2892 882
rect 3022 886 3028 887
rect 3022 882 3023 886
rect 3027 882 3028 886
rect 3022 881 3028 882
rect 3150 886 3156 887
rect 3150 882 3151 886
rect 3155 882 3156 886
rect 3150 881 3156 882
rect 3278 886 3284 887
rect 3278 882 3279 886
rect 3283 882 3284 886
rect 3278 881 3284 882
rect 3406 886 3412 887
rect 3406 882 3407 886
rect 3411 882 3412 886
rect 3406 881 3412 882
rect 3510 886 3516 887
rect 3510 882 3511 886
rect 3515 882 3516 886
rect 3510 881 3516 882
rect 1902 846 1908 847
rect 142 842 148 843
rect 142 838 143 842
rect 147 838 148 842
rect 142 837 148 838
rect 222 842 228 843
rect 222 838 223 842
rect 227 838 228 842
rect 222 837 228 838
rect 302 842 308 843
rect 302 838 303 842
rect 307 838 308 842
rect 302 837 308 838
rect 390 842 396 843
rect 390 838 391 842
rect 395 838 396 842
rect 390 837 396 838
rect 494 842 500 843
rect 494 838 495 842
rect 499 838 500 842
rect 494 837 500 838
rect 598 842 604 843
rect 598 838 599 842
rect 603 838 604 842
rect 598 837 604 838
rect 710 842 716 843
rect 710 838 711 842
rect 715 838 716 842
rect 710 837 716 838
rect 838 842 844 843
rect 838 838 839 842
rect 843 838 844 842
rect 838 837 844 838
rect 990 842 996 843
rect 990 838 991 842
rect 995 838 996 842
rect 990 837 996 838
rect 1166 842 1172 843
rect 1166 838 1167 842
rect 1171 838 1172 842
rect 1166 837 1172 838
rect 1358 842 1364 843
rect 1358 838 1359 842
rect 1363 838 1364 842
rect 1358 837 1364 838
rect 1566 842 1572 843
rect 1566 838 1567 842
rect 1571 838 1572 842
rect 1566 837 1572 838
rect 1750 842 1756 843
rect 1750 838 1751 842
rect 1755 838 1756 842
rect 1902 842 1903 846
rect 1907 842 1908 846
rect 1902 841 1908 842
rect 2038 846 2044 847
rect 2038 842 2039 846
rect 2043 842 2044 846
rect 2038 841 2044 842
rect 2214 846 2220 847
rect 2214 842 2215 846
rect 2219 842 2220 846
rect 2214 841 2220 842
rect 2390 846 2396 847
rect 2390 842 2391 846
rect 2395 842 2396 846
rect 2390 841 2396 842
rect 2566 846 2572 847
rect 2566 842 2567 846
rect 2571 842 2572 846
rect 2566 841 2572 842
rect 2734 846 2740 847
rect 2734 842 2735 846
rect 2739 842 2740 846
rect 2734 841 2740 842
rect 2886 846 2892 847
rect 2886 842 2887 846
rect 2891 842 2892 846
rect 2886 841 2892 842
rect 3030 846 3036 847
rect 3030 842 3031 846
rect 3035 842 3036 846
rect 3030 841 3036 842
rect 3158 846 3164 847
rect 3158 842 3159 846
rect 3163 842 3164 846
rect 3158 841 3164 842
rect 3286 846 3292 847
rect 3286 842 3287 846
rect 3291 842 3292 846
rect 3286 841 3292 842
rect 3406 846 3412 847
rect 3406 842 3407 846
rect 3411 842 3412 846
rect 3406 841 3412 842
rect 3510 846 3516 847
rect 3510 842 3511 846
rect 3515 842 3516 846
rect 3510 841 3516 842
rect 1750 837 1756 838
rect 1870 828 1876 829
rect 110 824 116 825
rect 110 820 111 824
rect 115 820 116 824
rect 110 819 116 820
rect 1830 824 1836 825
rect 1830 820 1831 824
rect 1835 820 1836 824
rect 1870 824 1871 828
rect 1875 824 1876 828
rect 1870 823 1876 824
rect 3590 828 3596 829
rect 3590 824 3591 828
rect 3595 824 3596 828
rect 3590 823 3596 824
rect 1830 819 1836 820
rect 1870 811 1876 812
rect 110 807 116 808
rect 110 803 111 807
rect 115 803 116 807
rect 1830 807 1836 808
rect 110 802 116 803
rect 134 804 140 805
rect 134 800 135 804
rect 139 800 140 804
rect 134 799 140 800
rect 214 804 220 805
rect 214 800 215 804
rect 219 800 220 804
rect 214 799 220 800
rect 294 804 300 805
rect 294 800 295 804
rect 299 800 300 804
rect 294 799 300 800
rect 382 804 388 805
rect 382 800 383 804
rect 387 800 388 804
rect 382 799 388 800
rect 486 804 492 805
rect 486 800 487 804
rect 491 800 492 804
rect 486 799 492 800
rect 590 804 596 805
rect 590 800 591 804
rect 595 800 596 804
rect 590 799 596 800
rect 702 804 708 805
rect 702 800 703 804
rect 707 800 708 804
rect 702 799 708 800
rect 830 804 836 805
rect 830 800 831 804
rect 835 800 836 804
rect 830 799 836 800
rect 982 804 988 805
rect 982 800 983 804
rect 987 800 988 804
rect 982 799 988 800
rect 1158 804 1164 805
rect 1158 800 1159 804
rect 1163 800 1164 804
rect 1158 799 1164 800
rect 1350 804 1356 805
rect 1350 800 1351 804
rect 1355 800 1356 804
rect 1350 799 1356 800
rect 1558 804 1564 805
rect 1558 800 1559 804
rect 1563 800 1564 804
rect 1558 799 1564 800
rect 1742 804 1748 805
rect 1742 800 1743 804
rect 1747 800 1748 804
rect 1830 803 1831 807
rect 1835 803 1836 807
rect 1870 807 1871 811
rect 1875 807 1876 811
rect 3590 811 3596 812
rect 1870 806 1876 807
rect 1894 808 1900 809
rect 1894 804 1895 808
rect 1899 804 1900 808
rect 1894 803 1900 804
rect 2030 808 2036 809
rect 2030 804 2031 808
rect 2035 804 2036 808
rect 2030 803 2036 804
rect 2206 808 2212 809
rect 2206 804 2207 808
rect 2211 804 2212 808
rect 2206 803 2212 804
rect 2382 808 2388 809
rect 2382 804 2383 808
rect 2387 804 2388 808
rect 2382 803 2388 804
rect 2558 808 2564 809
rect 2558 804 2559 808
rect 2563 804 2564 808
rect 2558 803 2564 804
rect 2726 808 2732 809
rect 2726 804 2727 808
rect 2731 804 2732 808
rect 2726 803 2732 804
rect 2878 808 2884 809
rect 2878 804 2879 808
rect 2883 804 2884 808
rect 2878 803 2884 804
rect 3022 808 3028 809
rect 3022 804 3023 808
rect 3027 804 3028 808
rect 3022 803 3028 804
rect 3150 808 3156 809
rect 3150 804 3151 808
rect 3155 804 3156 808
rect 3150 803 3156 804
rect 3278 808 3284 809
rect 3278 804 3279 808
rect 3283 804 3284 808
rect 3278 803 3284 804
rect 3398 808 3404 809
rect 3398 804 3399 808
rect 3403 804 3404 808
rect 3398 803 3404 804
rect 3502 808 3508 809
rect 3502 804 3503 808
rect 3507 804 3508 808
rect 3590 807 3591 811
rect 3595 807 3596 811
rect 3590 806 3596 807
rect 3502 803 3508 804
rect 1830 802 1836 803
rect 1742 799 1748 800
rect 198 756 204 757
rect 110 753 116 754
rect 110 749 111 753
rect 115 749 116 753
rect 198 752 199 756
rect 203 752 204 756
rect 198 751 204 752
rect 286 756 292 757
rect 286 752 287 756
rect 291 752 292 756
rect 286 751 292 752
rect 390 756 396 757
rect 390 752 391 756
rect 395 752 396 756
rect 390 751 396 752
rect 502 756 508 757
rect 502 752 503 756
rect 507 752 508 756
rect 502 751 508 752
rect 614 756 620 757
rect 614 752 615 756
rect 619 752 620 756
rect 614 751 620 752
rect 734 756 740 757
rect 734 752 735 756
rect 739 752 740 756
rect 734 751 740 752
rect 854 756 860 757
rect 854 752 855 756
rect 859 752 860 756
rect 854 751 860 752
rect 982 756 988 757
rect 982 752 983 756
rect 987 752 988 756
rect 982 751 988 752
rect 1110 756 1116 757
rect 1110 752 1111 756
rect 1115 752 1116 756
rect 1110 751 1116 752
rect 1238 756 1244 757
rect 1238 752 1239 756
rect 1243 752 1244 756
rect 1238 751 1244 752
rect 1366 756 1372 757
rect 1366 752 1367 756
rect 1371 752 1372 756
rect 1366 751 1372 752
rect 1494 756 1500 757
rect 1494 752 1495 756
rect 1499 752 1500 756
rect 1494 751 1500 752
rect 1630 756 1636 757
rect 1630 752 1631 756
rect 1635 752 1636 756
rect 1630 751 1636 752
rect 1742 756 1748 757
rect 1742 752 1743 756
rect 1747 752 1748 756
rect 1742 751 1748 752
rect 1830 753 1836 754
rect 110 748 116 749
rect 1830 749 1831 753
rect 1835 749 1836 753
rect 1830 748 1836 749
rect 2022 748 2028 749
rect 1870 745 1876 746
rect 1870 741 1871 745
rect 1875 741 1876 745
rect 2022 744 2023 748
rect 2027 744 2028 748
rect 2022 743 2028 744
rect 2190 748 2196 749
rect 2190 744 2191 748
rect 2195 744 2196 748
rect 2190 743 2196 744
rect 2358 748 2364 749
rect 2358 744 2359 748
rect 2363 744 2364 748
rect 2358 743 2364 744
rect 2518 748 2524 749
rect 2518 744 2519 748
rect 2523 744 2524 748
rect 2518 743 2524 744
rect 2678 748 2684 749
rect 2678 744 2679 748
rect 2683 744 2684 748
rect 2678 743 2684 744
rect 2830 748 2836 749
rect 2830 744 2831 748
rect 2835 744 2836 748
rect 2830 743 2836 744
rect 2974 748 2980 749
rect 2974 744 2975 748
rect 2979 744 2980 748
rect 2974 743 2980 744
rect 3110 748 3116 749
rect 3110 744 3111 748
rect 3115 744 3116 748
rect 3110 743 3116 744
rect 3246 748 3252 749
rect 3246 744 3247 748
rect 3251 744 3252 748
rect 3246 743 3252 744
rect 3382 748 3388 749
rect 3382 744 3383 748
rect 3387 744 3388 748
rect 3382 743 3388 744
rect 3502 748 3508 749
rect 3502 744 3503 748
rect 3507 744 3508 748
rect 3502 743 3508 744
rect 3590 745 3596 746
rect 1870 740 1876 741
rect 3590 741 3591 745
rect 3595 741 3596 745
rect 3590 740 3596 741
rect 110 736 116 737
rect 110 732 111 736
rect 115 732 116 736
rect 110 731 116 732
rect 1830 736 1836 737
rect 1830 732 1831 736
rect 1835 732 1836 736
rect 1830 731 1836 732
rect 1870 728 1876 729
rect 1870 724 1871 728
rect 1875 724 1876 728
rect 1870 723 1876 724
rect 3590 728 3596 729
rect 3590 724 3591 728
rect 3595 724 3596 728
rect 3590 723 3596 724
rect 206 718 212 719
rect 206 714 207 718
rect 211 714 212 718
rect 206 713 212 714
rect 294 718 300 719
rect 294 714 295 718
rect 299 714 300 718
rect 294 713 300 714
rect 398 718 404 719
rect 398 714 399 718
rect 403 714 404 718
rect 398 713 404 714
rect 510 718 516 719
rect 510 714 511 718
rect 515 714 516 718
rect 510 713 516 714
rect 622 718 628 719
rect 622 714 623 718
rect 627 714 628 718
rect 622 713 628 714
rect 742 718 748 719
rect 742 714 743 718
rect 747 714 748 718
rect 742 713 748 714
rect 862 718 868 719
rect 862 714 863 718
rect 867 714 868 718
rect 862 713 868 714
rect 990 718 996 719
rect 990 714 991 718
rect 995 714 996 718
rect 990 713 996 714
rect 1118 718 1124 719
rect 1118 714 1119 718
rect 1123 714 1124 718
rect 1118 713 1124 714
rect 1246 718 1252 719
rect 1246 714 1247 718
rect 1251 714 1252 718
rect 1246 713 1252 714
rect 1374 718 1380 719
rect 1374 714 1375 718
rect 1379 714 1380 718
rect 1374 713 1380 714
rect 1502 718 1508 719
rect 1502 714 1503 718
rect 1507 714 1508 718
rect 1502 713 1508 714
rect 1638 718 1644 719
rect 1638 714 1639 718
rect 1643 714 1644 718
rect 1638 713 1644 714
rect 1750 718 1756 719
rect 1750 714 1751 718
rect 1755 714 1756 718
rect 1750 713 1756 714
rect 2030 710 2036 711
rect 2030 706 2031 710
rect 2035 706 2036 710
rect 2030 705 2036 706
rect 2198 710 2204 711
rect 2198 706 2199 710
rect 2203 706 2204 710
rect 2198 705 2204 706
rect 2366 710 2372 711
rect 2366 706 2367 710
rect 2371 706 2372 710
rect 2366 705 2372 706
rect 2526 710 2532 711
rect 2526 706 2527 710
rect 2531 706 2532 710
rect 2526 705 2532 706
rect 2686 710 2692 711
rect 2686 706 2687 710
rect 2691 706 2692 710
rect 2686 705 2692 706
rect 2838 710 2844 711
rect 2838 706 2839 710
rect 2843 706 2844 710
rect 2838 705 2844 706
rect 2982 710 2988 711
rect 2982 706 2983 710
rect 2987 706 2988 710
rect 2982 705 2988 706
rect 3118 710 3124 711
rect 3118 706 3119 710
rect 3123 706 3124 710
rect 3118 705 3124 706
rect 3254 710 3260 711
rect 3254 706 3255 710
rect 3259 706 3260 710
rect 3254 705 3260 706
rect 3390 710 3396 711
rect 3390 706 3391 710
rect 3395 706 3396 710
rect 3390 705 3396 706
rect 3510 710 3516 711
rect 3510 706 3511 710
rect 3515 706 3516 710
rect 3510 705 3516 706
rect 2094 674 2100 675
rect 382 670 388 671
rect 382 666 383 670
rect 387 666 388 670
rect 382 665 388 666
rect 478 670 484 671
rect 478 666 479 670
rect 483 666 484 670
rect 478 665 484 666
rect 590 670 596 671
rect 590 666 591 670
rect 595 666 596 670
rect 590 665 596 666
rect 718 670 724 671
rect 718 666 719 670
rect 723 666 724 670
rect 718 665 724 666
rect 854 670 860 671
rect 854 666 855 670
rect 859 666 860 670
rect 854 665 860 666
rect 990 670 996 671
rect 990 666 991 670
rect 995 666 996 670
rect 990 665 996 666
rect 1126 670 1132 671
rect 1126 666 1127 670
rect 1131 666 1132 670
rect 1126 665 1132 666
rect 1254 670 1260 671
rect 1254 666 1255 670
rect 1259 666 1260 670
rect 1254 665 1260 666
rect 1382 670 1388 671
rect 1382 666 1383 670
rect 1387 666 1388 670
rect 1382 665 1388 666
rect 1502 670 1508 671
rect 1502 666 1503 670
rect 1507 666 1508 670
rect 1502 665 1508 666
rect 1630 670 1636 671
rect 1630 666 1631 670
rect 1635 666 1636 670
rect 1630 665 1636 666
rect 1750 670 1756 671
rect 1750 666 1751 670
rect 1755 666 1756 670
rect 2094 670 2095 674
rect 2099 670 2100 674
rect 2094 669 2100 670
rect 2174 674 2180 675
rect 2174 670 2175 674
rect 2179 670 2180 674
rect 2174 669 2180 670
rect 2262 674 2268 675
rect 2262 670 2263 674
rect 2267 670 2268 674
rect 2262 669 2268 670
rect 2358 674 2364 675
rect 2358 670 2359 674
rect 2363 670 2364 674
rect 2358 669 2364 670
rect 2462 674 2468 675
rect 2462 670 2463 674
rect 2467 670 2468 674
rect 2462 669 2468 670
rect 2566 674 2572 675
rect 2566 670 2567 674
rect 2571 670 2572 674
rect 2566 669 2572 670
rect 2678 674 2684 675
rect 2678 670 2679 674
rect 2683 670 2684 674
rect 2678 669 2684 670
rect 2798 674 2804 675
rect 2798 670 2799 674
rect 2803 670 2804 674
rect 2798 669 2804 670
rect 2926 674 2932 675
rect 2926 670 2927 674
rect 2931 670 2932 674
rect 2926 669 2932 670
rect 3070 674 3076 675
rect 3070 670 3071 674
rect 3075 670 3076 674
rect 3070 669 3076 670
rect 3222 674 3228 675
rect 3222 670 3223 674
rect 3227 670 3228 674
rect 3222 669 3228 670
rect 3374 674 3380 675
rect 3374 670 3375 674
rect 3379 670 3380 674
rect 3374 669 3380 670
rect 3510 674 3516 675
rect 3510 670 3511 674
rect 3515 670 3516 674
rect 3510 669 3516 670
rect 1750 665 1756 666
rect 1870 656 1876 657
rect 110 652 116 653
rect 110 648 111 652
rect 115 648 116 652
rect 110 647 116 648
rect 1830 652 1836 653
rect 1830 648 1831 652
rect 1835 648 1836 652
rect 1870 652 1871 656
rect 1875 652 1876 656
rect 1870 651 1876 652
rect 3590 656 3596 657
rect 3590 652 3591 656
rect 3595 652 3596 656
rect 3590 651 3596 652
rect 1830 647 1836 648
rect 1870 639 1876 640
rect 110 635 116 636
rect 110 631 111 635
rect 115 631 116 635
rect 1830 635 1836 636
rect 110 630 116 631
rect 374 632 380 633
rect 374 628 375 632
rect 379 628 380 632
rect 374 627 380 628
rect 470 632 476 633
rect 470 628 471 632
rect 475 628 476 632
rect 470 627 476 628
rect 582 632 588 633
rect 582 628 583 632
rect 587 628 588 632
rect 582 627 588 628
rect 710 632 716 633
rect 710 628 711 632
rect 715 628 716 632
rect 710 627 716 628
rect 846 632 852 633
rect 846 628 847 632
rect 851 628 852 632
rect 846 627 852 628
rect 982 632 988 633
rect 982 628 983 632
rect 987 628 988 632
rect 982 627 988 628
rect 1118 632 1124 633
rect 1118 628 1119 632
rect 1123 628 1124 632
rect 1118 627 1124 628
rect 1246 632 1252 633
rect 1246 628 1247 632
rect 1251 628 1252 632
rect 1246 627 1252 628
rect 1374 632 1380 633
rect 1374 628 1375 632
rect 1379 628 1380 632
rect 1374 627 1380 628
rect 1494 632 1500 633
rect 1494 628 1495 632
rect 1499 628 1500 632
rect 1494 627 1500 628
rect 1622 632 1628 633
rect 1622 628 1623 632
rect 1627 628 1628 632
rect 1622 627 1628 628
rect 1742 632 1748 633
rect 1742 628 1743 632
rect 1747 628 1748 632
rect 1830 631 1831 635
rect 1835 631 1836 635
rect 1870 635 1871 639
rect 1875 635 1876 639
rect 3590 639 3596 640
rect 1870 634 1876 635
rect 2086 636 2092 637
rect 2086 632 2087 636
rect 2091 632 2092 636
rect 2086 631 2092 632
rect 2166 636 2172 637
rect 2166 632 2167 636
rect 2171 632 2172 636
rect 2166 631 2172 632
rect 2254 636 2260 637
rect 2254 632 2255 636
rect 2259 632 2260 636
rect 2254 631 2260 632
rect 2350 636 2356 637
rect 2350 632 2351 636
rect 2355 632 2356 636
rect 2350 631 2356 632
rect 2454 636 2460 637
rect 2454 632 2455 636
rect 2459 632 2460 636
rect 2454 631 2460 632
rect 2558 636 2564 637
rect 2558 632 2559 636
rect 2563 632 2564 636
rect 2558 631 2564 632
rect 2670 636 2676 637
rect 2670 632 2671 636
rect 2675 632 2676 636
rect 2670 631 2676 632
rect 2790 636 2796 637
rect 2790 632 2791 636
rect 2795 632 2796 636
rect 2790 631 2796 632
rect 2918 636 2924 637
rect 2918 632 2919 636
rect 2923 632 2924 636
rect 2918 631 2924 632
rect 3062 636 3068 637
rect 3062 632 3063 636
rect 3067 632 3068 636
rect 3062 631 3068 632
rect 3214 636 3220 637
rect 3214 632 3215 636
rect 3219 632 3220 636
rect 3214 631 3220 632
rect 3366 636 3372 637
rect 3366 632 3367 636
rect 3371 632 3372 636
rect 3366 631 3372 632
rect 3502 636 3508 637
rect 3502 632 3503 636
rect 3507 632 3508 636
rect 3590 635 3591 639
rect 3595 635 3596 639
rect 3590 634 3596 635
rect 3502 631 3508 632
rect 1830 630 1836 631
rect 1742 627 1748 628
rect 598 580 604 581
rect 110 577 116 578
rect 110 573 111 577
rect 115 573 116 577
rect 598 576 599 580
rect 603 576 604 580
rect 598 575 604 576
rect 686 580 692 581
rect 686 576 687 580
rect 691 576 692 580
rect 686 575 692 576
rect 782 580 788 581
rect 782 576 783 580
rect 787 576 788 580
rect 782 575 788 576
rect 886 580 892 581
rect 886 576 887 580
rect 891 576 892 580
rect 886 575 892 576
rect 990 580 996 581
rect 990 576 991 580
rect 995 576 996 580
rect 990 575 996 576
rect 1094 580 1100 581
rect 1094 576 1095 580
rect 1099 576 1100 580
rect 1094 575 1100 576
rect 1198 580 1204 581
rect 1198 576 1199 580
rect 1203 576 1204 580
rect 1198 575 1204 576
rect 1302 580 1308 581
rect 1302 576 1303 580
rect 1307 576 1308 580
rect 1302 575 1308 576
rect 1398 580 1404 581
rect 1398 576 1399 580
rect 1403 576 1404 580
rect 1398 575 1404 576
rect 1502 580 1508 581
rect 1502 576 1503 580
rect 1507 576 1508 580
rect 1502 575 1508 576
rect 1606 580 1612 581
rect 1606 576 1607 580
rect 1611 576 1612 580
rect 1606 575 1612 576
rect 1710 580 1716 581
rect 1710 576 1711 580
rect 1715 576 1716 580
rect 2166 580 2172 581
rect 1710 575 1716 576
rect 1830 577 1836 578
rect 110 572 116 573
rect 1830 573 1831 577
rect 1835 573 1836 577
rect 1830 572 1836 573
rect 1870 577 1876 578
rect 1870 573 1871 577
rect 1875 573 1876 577
rect 2166 576 2167 580
rect 2171 576 2172 580
rect 2166 575 2172 576
rect 2246 580 2252 581
rect 2246 576 2247 580
rect 2251 576 2252 580
rect 2246 575 2252 576
rect 2326 580 2332 581
rect 2326 576 2327 580
rect 2331 576 2332 580
rect 2326 575 2332 576
rect 2406 580 2412 581
rect 2406 576 2407 580
rect 2411 576 2412 580
rect 2406 575 2412 576
rect 2486 580 2492 581
rect 2486 576 2487 580
rect 2491 576 2492 580
rect 2486 575 2492 576
rect 2566 580 2572 581
rect 2566 576 2567 580
rect 2571 576 2572 580
rect 2566 575 2572 576
rect 2646 580 2652 581
rect 2646 576 2647 580
rect 2651 576 2652 580
rect 2646 575 2652 576
rect 2742 580 2748 581
rect 2742 576 2743 580
rect 2747 576 2748 580
rect 2742 575 2748 576
rect 2862 580 2868 581
rect 2862 576 2863 580
rect 2867 576 2868 580
rect 2862 575 2868 576
rect 2998 580 3004 581
rect 2998 576 2999 580
rect 3003 576 3004 580
rect 2998 575 3004 576
rect 3158 580 3164 581
rect 3158 576 3159 580
rect 3163 576 3164 580
rect 3158 575 3164 576
rect 3326 580 3332 581
rect 3326 576 3327 580
rect 3331 576 3332 580
rect 3326 575 3332 576
rect 3494 580 3500 581
rect 3494 576 3495 580
rect 3499 576 3500 580
rect 3494 575 3500 576
rect 3590 577 3596 578
rect 1870 572 1876 573
rect 3590 573 3591 577
rect 3595 573 3596 577
rect 3590 572 3596 573
rect 110 560 116 561
rect 110 556 111 560
rect 115 556 116 560
rect 110 555 116 556
rect 1830 560 1836 561
rect 1830 556 1831 560
rect 1835 556 1836 560
rect 1830 555 1836 556
rect 1870 560 1876 561
rect 1870 556 1871 560
rect 1875 556 1876 560
rect 1870 555 1876 556
rect 3590 560 3596 561
rect 3590 556 3591 560
rect 3595 556 3596 560
rect 3590 555 3596 556
rect 606 542 612 543
rect 606 538 607 542
rect 611 538 612 542
rect 606 537 612 538
rect 694 542 700 543
rect 694 538 695 542
rect 699 538 700 542
rect 694 537 700 538
rect 790 542 796 543
rect 790 538 791 542
rect 795 538 796 542
rect 790 537 796 538
rect 894 542 900 543
rect 894 538 895 542
rect 899 538 900 542
rect 894 537 900 538
rect 998 542 1004 543
rect 998 538 999 542
rect 1003 538 1004 542
rect 998 537 1004 538
rect 1102 542 1108 543
rect 1102 538 1103 542
rect 1107 538 1108 542
rect 1102 537 1108 538
rect 1206 542 1212 543
rect 1206 538 1207 542
rect 1211 538 1212 542
rect 1206 537 1212 538
rect 1310 542 1316 543
rect 1310 538 1311 542
rect 1315 538 1316 542
rect 1310 537 1316 538
rect 1406 542 1412 543
rect 1406 538 1407 542
rect 1411 538 1412 542
rect 1406 537 1412 538
rect 1510 542 1516 543
rect 1510 538 1511 542
rect 1515 538 1516 542
rect 1510 537 1516 538
rect 1614 542 1620 543
rect 1614 538 1615 542
rect 1619 538 1620 542
rect 1614 537 1620 538
rect 1718 542 1724 543
rect 1718 538 1719 542
rect 1723 538 1724 542
rect 1718 537 1724 538
rect 2174 542 2180 543
rect 2174 538 2175 542
rect 2179 538 2180 542
rect 2174 537 2180 538
rect 2254 542 2260 543
rect 2254 538 2255 542
rect 2259 538 2260 542
rect 2254 537 2260 538
rect 2334 542 2340 543
rect 2334 538 2335 542
rect 2339 538 2340 542
rect 2334 537 2340 538
rect 2414 542 2420 543
rect 2414 538 2415 542
rect 2419 538 2420 542
rect 2414 537 2420 538
rect 2494 542 2500 543
rect 2494 538 2495 542
rect 2499 538 2500 542
rect 2494 537 2500 538
rect 2574 542 2580 543
rect 2574 538 2575 542
rect 2579 538 2580 542
rect 2574 537 2580 538
rect 2654 542 2660 543
rect 2654 538 2655 542
rect 2659 538 2660 542
rect 2654 537 2660 538
rect 2750 542 2756 543
rect 2750 538 2751 542
rect 2755 538 2756 542
rect 2750 537 2756 538
rect 2870 542 2876 543
rect 2870 538 2871 542
rect 2875 538 2876 542
rect 2870 537 2876 538
rect 3006 542 3012 543
rect 3006 538 3007 542
rect 3011 538 3012 542
rect 3006 537 3012 538
rect 3166 542 3172 543
rect 3166 538 3167 542
rect 3171 538 3172 542
rect 3166 537 3172 538
rect 3334 542 3340 543
rect 3334 538 3335 542
rect 3339 538 3340 542
rect 3334 537 3340 538
rect 3502 542 3508 543
rect 3502 538 3503 542
rect 3507 538 3508 542
rect 3502 537 3508 538
rect 366 502 372 503
rect 366 498 367 502
rect 371 498 372 502
rect 366 497 372 498
rect 462 502 468 503
rect 462 498 463 502
rect 467 498 468 502
rect 462 497 468 498
rect 574 502 580 503
rect 574 498 575 502
rect 579 498 580 502
rect 574 497 580 498
rect 702 502 708 503
rect 702 498 703 502
rect 707 498 708 502
rect 702 497 708 498
rect 838 502 844 503
rect 838 498 839 502
rect 843 498 844 502
rect 838 497 844 498
rect 974 502 980 503
rect 974 498 975 502
rect 979 498 980 502
rect 974 497 980 498
rect 1110 502 1116 503
rect 1110 498 1111 502
rect 1115 498 1116 502
rect 1110 497 1116 498
rect 1238 502 1244 503
rect 1238 498 1239 502
rect 1243 498 1244 502
rect 1238 497 1244 498
rect 1358 502 1364 503
rect 1358 498 1359 502
rect 1363 498 1364 502
rect 1358 497 1364 498
rect 1470 502 1476 503
rect 1470 498 1471 502
rect 1475 498 1476 502
rect 1470 497 1476 498
rect 1582 502 1588 503
rect 1582 498 1583 502
rect 1587 498 1588 502
rect 1582 497 1588 498
rect 1702 502 1708 503
rect 1702 498 1703 502
rect 1707 498 1708 502
rect 1702 497 1708 498
rect 2158 502 2164 503
rect 2158 498 2159 502
rect 2163 498 2164 502
rect 2158 497 2164 498
rect 2238 502 2244 503
rect 2238 498 2239 502
rect 2243 498 2244 502
rect 2238 497 2244 498
rect 2318 502 2324 503
rect 2318 498 2319 502
rect 2323 498 2324 502
rect 2318 497 2324 498
rect 2398 502 2404 503
rect 2398 498 2399 502
rect 2403 498 2404 502
rect 2398 497 2404 498
rect 2478 502 2484 503
rect 2478 498 2479 502
rect 2483 498 2484 502
rect 2478 497 2484 498
rect 2558 502 2564 503
rect 2558 498 2559 502
rect 2563 498 2564 502
rect 2558 497 2564 498
rect 2638 502 2644 503
rect 2638 498 2639 502
rect 2643 498 2644 502
rect 2638 497 2644 498
rect 2734 502 2740 503
rect 2734 498 2735 502
rect 2739 498 2740 502
rect 2734 497 2740 498
rect 2854 502 2860 503
rect 2854 498 2855 502
rect 2859 498 2860 502
rect 2854 497 2860 498
rect 2990 502 2996 503
rect 2990 498 2991 502
rect 2995 498 2996 502
rect 2990 497 2996 498
rect 3142 502 3148 503
rect 3142 498 3143 502
rect 3147 498 3148 502
rect 3142 497 3148 498
rect 3310 502 3316 503
rect 3310 498 3311 502
rect 3315 498 3316 502
rect 3310 497 3316 498
rect 3478 502 3484 503
rect 3478 498 3479 502
rect 3483 498 3484 502
rect 3478 497 3484 498
rect 110 484 116 485
rect 110 480 111 484
rect 115 480 116 484
rect 110 479 116 480
rect 1830 484 1836 485
rect 1830 480 1831 484
rect 1835 480 1836 484
rect 1830 479 1836 480
rect 1870 484 1876 485
rect 1870 480 1871 484
rect 1875 480 1876 484
rect 1870 479 1876 480
rect 3590 484 3596 485
rect 3590 480 3591 484
rect 3595 480 3596 484
rect 3590 479 3596 480
rect 110 467 116 468
rect 110 463 111 467
rect 115 463 116 467
rect 1830 467 1836 468
rect 110 462 116 463
rect 358 464 364 465
rect 358 460 359 464
rect 363 460 364 464
rect 358 459 364 460
rect 454 464 460 465
rect 454 460 455 464
rect 459 460 460 464
rect 454 459 460 460
rect 566 464 572 465
rect 566 460 567 464
rect 571 460 572 464
rect 566 459 572 460
rect 694 464 700 465
rect 694 460 695 464
rect 699 460 700 464
rect 694 459 700 460
rect 830 464 836 465
rect 830 460 831 464
rect 835 460 836 464
rect 830 459 836 460
rect 966 464 972 465
rect 966 460 967 464
rect 971 460 972 464
rect 966 459 972 460
rect 1102 464 1108 465
rect 1102 460 1103 464
rect 1107 460 1108 464
rect 1102 459 1108 460
rect 1230 464 1236 465
rect 1230 460 1231 464
rect 1235 460 1236 464
rect 1230 459 1236 460
rect 1350 464 1356 465
rect 1350 460 1351 464
rect 1355 460 1356 464
rect 1350 459 1356 460
rect 1462 464 1468 465
rect 1462 460 1463 464
rect 1467 460 1468 464
rect 1462 459 1468 460
rect 1574 464 1580 465
rect 1574 460 1575 464
rect 1579 460 1580 464
rect 1574 459 1580 460
rect 1694 464 1700 465
rect 1694 460 1695 464
rect 1699 460 1700 464
rect 1830 463 1831 467
rect 1835 463 1836 467
rect 1830 462 1836 463
rect 1870 467 1876 468
rect 1870 463 1871 467
rect 1875 463 1876 467
rect 3590 467 3596 468
rect 1870 462 1876 463
rect 2150 464 2156 465
rect 1694 459 1700 460
rect 2150 460 2151 464
rect 2155 460 2156 464
rect 2150 459 2156 460
rect 2230 464 2236 465
rect 2230 460 2231 464
rect 2235 460 2236 464
rect 2230 459 2236 460
rect 2310 464 2316 465
rect 2310 460 2311 464
rect 2315 460 2316 464
rect 2310 459 2316 460
rect 2390 464 2396 465
rect 2390 460 2391 464
rect 2395 460 2396 464
rect 2390 459 2396 460
rect 2470 464 2476 465
rect 2470 460 2471 464
rect 2475 460 2476 464
rect 2470 459 2476 460
rect 2550 464 2556 465
rect 2550 460 2551 464
rect 2555 460 2556 464
rect 2550 459 2556 460
rect 2630 464 2636 465
rect 2630 460 2631 464
rect 2635 460 2636 464
rect 2630 459 2636 460
rect 2726 464 2732 465
rect 2726 460 2727 464
rect 2731 460 2732 464
rect 2726 459 2732 460
rect 2846 464 2852 465
rect 2846 460 2847 464
rect 2851 460 2852 464
rect 2846 459 2852 460
rect 2982 464 2988 465
rect 2982 460 2983 464
rect 2987 460 2988 464
rect 2982 459 2988 460
rect 3134 464 3140 465
rect 3134 460 3135 464
rect 3139 460 3140 464
rect 3134 459 3140 460
rect 3302 464 3308 465
rect 3302 460 3303 464
rect 3307 460 3308 464
rect 3302 459 3308 460
rect 3470 464 3476 465
rect 3470 460 3471 464
rect 3475 460 3476 464
rect 3590 463 3591 467
rect 3595 463 3596 467
rect 3590 462 3596 463
rect 3470 459 3476 460
rect 134 408 140 409
rect 110 405 116 406
rect 110 401 111 405
rect 115 401 116 405
rect 134 404 135 408
rect 139 404 140 408
rect 134 403 140 404
rect 222 408 228 409
rect 222 404 223 408
rect 227 404 228 408
rect 222 403 228 404
rect 358 408 364 409
rect 358 404 359 408
rect 363 404 364 408
rect 358 403 364 404
rect 510 408 516 409
rect 510 404 511 408
rect 515 404 516 408
rect 510 403 516 404
rect 678 408 684 409
rect 678 404 679 408
rect 683 404 684 408
rect 678 403 684 404
rect 838 408 844 409
rect 838 404 839 408
rect 843 404 844 408
rect 838 403 844 404
rect 998 408 1004 409
rect 998 404 999 408
rect 1003 404 1004 408
rect 998 403 1004 404
rect 1142 408 1148 409
rect 1142 404 1143 408
rect 1147 404 1148 408
rect 1142 403 1148 404
rect 1278 408 1284 409
rect 1278 404 1279 408
rect 1283 404 1284 408
rect 1278 403 1284 404
rect 1414 408 1420 409
rect 1414 404 1415 408
rect 1419 404 1420 408
rect 1414 403 1420 404
rect 1550 408 1556 409
rect 1550 404 1551 408
rect 1555 404 1556 408
rect 1550 403 1556 404
rect 1686 408 1692 409
rect 1686 404 1687 408
rect 1691 404 1692 408
rect 2158 408 2164 409
rect 1686 403 1692 404
rect 1830 405 1836 406
rect 110 400 116 401
rect 1830 401 1831 405
rect 1835 401 1836 405
rect 1830 400 1836 401
rect 1870 405 1876 406
rect 1870 401 1871 405
rect 1875 401 1876 405
rect 2158 404 2159 408
rect 2163 404 2164 408
rect 2158 403 2164 404
rect 2238 408 2244 409
rect 2238 404 2239 408
rect 2243 404 2244 408
rect 2238 403 2244 404
rect 2318 408 2324 409
rect 2318 404 2319 408
rect 2323 404 2324 408
rect 2318 403 2324 404
rect 2398 408 2404 409
rect 2398 404 2399 408
rect 2403 404 2404 408
rect 2398 403 2404 404
rect 2478 408 2484 409
rect 2478 404 2479 408
rect 2483 404 2484 408
rect 2478 403 2484 404
rect 2558 408 2564 409
rect 2558 404 2559 408
rect 2563 404 2564 408
rect 2558 403 2564 404
rect 2638 408 2644 409
rect 2638 404 2639 408
rect 2643 404 2644 408
rect 2638 403 2644 404
rect 2734 408 2740 409
rect 2734 404 2735 408
rect 2739 404 2740 408
rect 2734 403 2740 404
rect 2838 408 2844 409
rect 2838 404 2839 408
rect 2843 404 2844 408
rect 2838 403 2844 404
rect 2958 408 2964 409
rect 2958 404 2959 408
rect 2963 404 2964 408
rect 2958 403 2964 404
rect 3086 408 3092 409
rect 3086 404 3087 408
rect 3091 404 3092 408
rect 3086 403 3092 404
rect 3230 408 3236 409
rect 3230 404 3231 408
rect 3235 404 3236 408
rect 3230 403 3236 404
rect 3374 408 3380 409
rect 3374 404 3375 408
rect 3379 404 3380 408
rect 3374 403 3380 404
rect 3502 408 3508 409
rect 3502 404 3503 408
rect 3507 404 3508 408
rect 3502 403 3508 404
rect 3590 405 3596 406
rect 1870 400 1876 401
rect 3590 401 3591 405
rect 3595 401 3596 405
rect 3590 400 3596 401
rect 110 388 116 389
rect 110 384 111 388
rect 115 384 116 388
rect 110 383 116 384
rect 1830 388 1836 389
rect 1830 384 1831 388
rect 1835 384 1836 388
rect 1830 383 1836 384
rect 1870 388 1876 389
rect 1870 384 1871 388
rect 1875 384 1876 388
rect 1870 383 1876 384
rect 3590 388 3596 389
rect 3590 384 3591 388
rect 3595 384 3596 388
rect 3590 383 3596 384
rect 142 370 148 371
rect 142 366 143 370
rect 147 366 148 370
rect 142 365 148 366
rect 230 370 236 371
rect 230 366 231 370
rect 235 366 236 370
rect 230 365 236 366
rect 366 370 372 371
rect 366 366 367 370
rect 371 366 372 370
rect 366 365 372 366
rect 518 370 524 371
rect 518 366 519 370
rect 523 366 524 370
rect 518 365 524 366
rect 686 370 692 371
rect 686 366 687 370
rect 691 366 692 370
rect 686 365 692 366
rect 846 370 852 371
rect 846 366 847 370
rect 851 366 852 370
rect 846 365 852 366
rect 1006 370 1012 371
rect 1006 366 1007 370
rect 1011 366 1012 370
rect 1006 365 1012 366
rect 1150 370 1156 371
rect 1150 366 1151 370
rect 1155 366 1156 370
rect 1150 365 1156 366
rect 1286 370 1292 371
rect 1286 366 1287 370
rect 1291 366 1292 370
rect 1286 365 1292 366
rect 1422 370 1428 371
rect 1422 366 1423 370
rect 1427 366 1428 370
rect 1422 365 1428 366
rect 1558 370 1564 371
rect 1558 366 1559 370
rect 1563 366 1564 370
rect 1558 365 1564 366
rect 1694 370 1700 371
rect 1694 366 1695 370
rect 1699 366 1700 370
rect 1694 365 1700 366
rect 2166 370 2172 371
rect 2166 366 2167 370
rect 2171 366 2172 370
rect 2166 365 2172 366
rect 2246 370 2252 371
rect 2246 366 2247 370
rect 2251 366 2252 370
rect 2246 365 2252 366
rect 2326 370 2332 371
rect 2326 366 2327 370
rect 2331 366 2332 370
rect 2326 365 2332 366
rect 2406 370 2412 371
rect 2406 366 2407 370
rect 2411 366 2412 370
rect 2406 365 2412 366
rect 2486 370 2492 371
rect 2486 366 2487 370
rect 2491 366 2492 370
rect 2486 365 2492 366
rect 2566 370 2572 371
rect 2566 366 2567 370
rect 2571 366 2572 370
rect 2566 365 2572 366
rect 2646 370 2652 371
rect 2646 366 2647 370
rect 2651 366 2652 370
rect 2646 365 2652 366
rect 2742 370 2748 371
rect 2742 366 2743 370
rect 2747 366 2748 370
rect 2742 365 2748 366
rect 2846 370 2852 371
rect 2846 366 2847 370
rect 2851 366 2852 370
rect 2846 365 2852 366
rect 2966 370 2972 371
rect 2966 366 2967 370
rect 2971 366 2972 370
rect 2966 365 2972 366
rect 3094 370 3100 371
rect 3094 366 3095 370
rect 3099 366 3100 370
rect 3094 365 3100 366
rect 3238 370 3244 371
rect 3238 366 3239 370
rect 3243 366 3244 370
rect 3238 365 3244 366
rect 3382 370 3388 371
rect 3382 366 3383 370
rect 3387 366 3388 370
rect 3382 365 3388 366
rect 3510 370 3516 371
rect 3510 366 3511 370
rect 3515 366 3516 370
rect 3510 365 3516 366
rect 142 330 148 331
rect 142 326 143 330
rect 147 326 148 330
rect 142 325 148 326
rect 278 330 284 331
rect 278 326 279 330
rect 283 326 284 330
rect 278 325 284 326
rect 454 330 460 331
rect 454 326 455 330
rect 459 326 460 330
rect 454 325 460 326
rect 638 330 644 331
rect 638 326 639 330
rect 643 326 644 330
rect 638 325 644 326
rect 822 330 828 331
rect 822 326 823 330
rect 827 326 828 330
rect 822 325 828 326
rect 998 330 1004 331
rect 998 326 999 330
rect 1003 326 1004 330
rect 998 325 1004 326
rect 1166 330 1172 331
rect 1166 326 1167 330
rect 1171 326 1172 330
rect 1166 325 1172 326
rect 1326 330 1332 331
rect 1326 326 1327 330
rect 1331 326 1332 330
rect 1326 325 1332 326
rect 1478 330 1484 331
rect 1478 326 1479 330
rect 1483 326 1484 330
rect 1478 325 1484 326
rect 1622 330 1628 331
rect 1622 326 1623 330
rect 1627 326 1628 330
rect 1622 325 1628 326
rect 1750 330 1756 331
rect 1750 326 1751 330
rect 1755 326 1756 330
rect 1750 325 1756 326
rect 2030 326 2036 327
rect 2030 322 2031 326
rect 2035 322 2036 326
rect 2030 321 2036 322
rect 2118 326 2124 327
rect 2118 322 2119 326
rect 2123 322 2124 326
rect 2118 321 2124 322
rect 2222 326 2228 327
rect 2222 322 2223 326
rect 2227 322 2228 326
rect 2222 321 2228 322
rect 2334 326 2340 327
rect 2334 322 2335 326
rect 2339 322 2340 326
rect 2334 321 2340 322
rect 2446 326 2452 327
rect 2446 322 2447 326
rect 2451 322 2452 326
rect 2446 321 2452 322
rect 2566 326 2572 327
rect 2566 322 2567 326
rect 2571 322 2572 326
rect 2566 321 2572 322
rect 2694 326 2700 327
rect 2694 322 2695 326
rect 2699 322 2700 326
rect 2694 321 2700 322
rect 2838 326 2844 327
rect 2838 322 2839 326
rect 2843 322 2844 326
rect 2838 321 2844 322
rect 2998 326 3004 327
rect 2998 322 2999 326
rect 3003 322 3004 326
rect 2998 321 3004 322
rect 3166 326 3172 327
rect 3166 322 3167 326
rect 3171 322 3172 326
rect 3166 321 3172 322
rect 3342 326 3348 327
rect 3342 322 3343 326
rect 3347 322 3348 326
rect 3342 321 3348 322
rect 3510 326 3516 327
rect 3510 322 3511 326
rect 3515 322 3516 326
rect 3510 321 3516 322
rect 110 312 116 313
rect 110 308 111 312
rect 115 308 116 312
rect 110 307 116 308
rect 1830 312 1836 313
rect 1830 308 1831 312
rect 1835 308 1836 312
rect 1830 307 1836 308
rect 1870 308 1876 309
rect 1870 304 1871 308
rect 1875 304 1876 308
rect 1870 303 1876 304
rect 3590 308 3596 309
rect 3590 304 3591 308
rect 3595 304 3596 308
rect 3590 303 3596 304
rect 110 295 116 296
rect 110 291 111 295
rect 115 291 116 295
rect 1830 295 1836 296
rect 110 290 116 291
rect 134 292 140 293
rect 134 288 135 292
rect 139 288 140 292
rect 134 287 140 288
rect 270 292 276 293
rect 270 288 271 292
rect 275 288 276 292
rect 270 287 276 288
rect 446 292 452 293
rect 446 288 447 292
rect 451 288 452 292
rect 446 287 452 288
rect 630 292 636 293
rect 630 288 631 292
rect 635 288 636 292
rect 630 287 636 288
rect 814 292 820 293
rect 814 288 815 292
rect 819 288 820 292
rect 814 287 820 288
rect 990 292 996 293
rect 990 288 991 292
rect 995 288 996 292
rect 990 287 996 288
rect 1158 292 1164 293
rect 1158 288 1159 292
rect 1163 288 1164 292
rect 1158 287 1164 288
rect 1318 292 1324 293
rect 1318 288 1319 292
rect 1323 288 1324 292
rect 1318 287 1324 288
rect 1470 292 1476 293
rect 1470 288 1471 292
rect 1475 288 1476 292
rect 1470 287 1476 288
rect 1614 292 1620 293
rect 1614 288 1615 292
rect 1619 288 1620 292
rect 1614 287 1620 288
rect 1742 292 1748 293
rect 1742 288 1743 292
rect 1747 288 1748 292
rect 1830 291 1831 295
rect 1835 291 1836 295
rect 1830 290 1836 291
rect 1870 291 1876 292
rect 1742 287 1748 288
rect 1870 287 1871 291
rect 1875 287 1876 291
rect 3590 291 3596 292
rect 1870 286 1876 287
rect 2022 288 2028 289
rect 2022 284 2023 288
rect 2027 284 2028 288
rect 2022 283 2028 284
rect 2110 288 2116 289
rect 2110 284 2111 288
rect 2115 284 2116 288
rect 2110 283 2116 284
rect 2214 288 2220 289
rect 2214 284 2215 288
rect 2219 284 2220 288
rect 2214 283 2220 284
rect 2326 288 2332 289
rect 2326 284 2327 288
rect 2331 284 2332 288
rect 2326 283 2332 284
rect 2438 288 2444 289
rect 2438 284 2439 288
rect 2443 284 2444 288
rect 2438 283 2444 284
rect 2558 288 2564 289
rect 2558 284 2559 288
rect 2563 284 2564 288
rect 2558 283 2564 284
rect 2686 288 2692 289
rect 2686 284 2687 288
rect 2691 284 2692 288
rect 2686 283 2692 284
rect 2830 288 2836 289
rect 2830 284 2831 288
rect 2835 284 2836 288
rect 2830 283 2836 284
rect 2990 288 2996 289
rect 2990 284 2991 288
rect 2995 284 2996 288
rect 2990 283 2996 284
rect 3158 288 3164 289
rect 3158 284 3159 288
rect 3163 284 3164 288
rect 3158 283 3164 284
rect 3334 288 3340 289
rect 3334 284 3335 288
rect 3339 284 3340 288
rect 3334 283 3340 284
rect 3502 288 3508 289
rect 3502 284 3503 288
rect 3507 284 3508 288
rect 3590 287 3591 291
rect 3595 287 3596 291
rect 3590 286 3596 287
rect 3502 283 3508 284
rect 302 244 308 245
rect 110 241 116 242
rect 110 237 111 241
rect 115 237 116 241
rect 302 240 303 244
rect 307 240 308 244
rect 302 239 308 240
rect 390 244 396 245
rect 390 240 391 244
rect 395 240 396 244
rect 390 239 396 240
rect 494 244 500 245
rect 494 240 495 244
rect 499 240 500 244
rect 494 239 500 240
rect 598 244 604 245
rect 598 240 599 244
rect 603 240 604 244
rect 598 239 604 240
rect 710 244 716 245
rect 710 240 711 244
rect 715 240 716 244
rect 710 239 716 240
rect 822 244 828 245
rect 822 240 823 244
rect 827 240 828 244
rect 822 239 828 240
rect 942 244 948 245
rect 942 240 943 244
rect 947 240 948 244
rect 942 239 948 240
rect 1062 244 1068 245
rect 1062 240 1063 244
rect 1067 240 1068 244
rect 1062 239 1068 240
rect 1174 244 1180 245
rect 1174 240 1175 244
rect 1179 240 1180 244
rect 1174 239 1180 240
rect 1286 244 1292 245
rect 1286 240 1287 244
rect 1291 240 1292 244
rect 1286 239 1292 240
rect 1406 244 1412 245
rect 1406 240 1407 244
rect 1411 240 1412 244
rect 1406 239 1412 240
rect 1526 244 1532 245
rect 1526 240 1527 244
rect 1531 240 1532 244
rect 1526 239 1532 240
rect 1646 244 1652 245
rect 1646 240 1647 244
rect 1651 240 1652 244
rect 1646 239 1652 240
rect 1742 244 1748 245
rect 1742 240 1743 244
rect 1747 240 1748 244
rect 1742 239 1748 240
rect 1830 241 1836 242
rect 110 236 116 237
rect 1830 237 1831 241
rect 1835 237 1836 241
rect 2070 240 2076 241
rect 1830 236 1836 237
rect 1870 237 1876 238
rect 1870 233 1871 237
rect 1875 233 1876 237
rect 2070 236 2071 240
rect 2075 236 2076 240
rect 2070 235 2076 236
rect 2318 240 2324 241
rect 2318 236 2319 240
rect 2323 236 2324 240
rect 2318 235 2324 236
rect 2542 240 2548 241
rect 2542 236 2543 240
rect 2547 236 2548 240
rect 2542 235 2548 236
rect 2742 240 2748 241
rect 2742 236 2743 240
rect 2747 236 2748 240
rect 2742 235 2748 236
rect 2926 240 2932 241
rect 2926 236 2927 240
rect 2931 236 2932 240
rect 2926 235 2932 236
rect 3086 240 3092 241
rect 3086 236 3087 240
rect 3091 236 3092 240
rect 3086 235 3092 236
rect 3238 240 3244 241
rect 3238 236 3239 240
rect 3243 236 3244 240
rect 3238 235 3244 236
rect 3382 240 3388 241
rect 3382 236 3383 240
rect 3387 236 3388 240
rect 3382 235 3388 236
rect 3502 240 3508 241
rect 3502 236 3503 240
rect 3507 236 3508 240
rect 3502 235 3508 236
rect 3590 237 3596 238
rect 1870 232 1876 233
rect 3590 233 3591 237
rect 3595 233 3596 237
rect 3590 232 3596 233
rect 110 224 116 225
rect 110 220 111 224
rect 115 220 116 224
rect 110 219 116 220
rect 1830 224 1836 225
rect 1830 220 1831 224
rect 1835 220 1836 224
rect 1830 219 1836 220
rect 1870 220 1876 221
rect 1870 216 1871 220
rect 1875 216 1876 220
rect 1870 215 1876 216
rect 3590 220 3596 221
rect 3590 216 3591 220
rect 3595 216 3596 220
rect 3590 215 3596 216
rect 310 206 316 207
rect 310 202 311 206
rect 315 202 316 206
rect 310 201 316 202
rect 398 206 404 207
rect 398 202 399 206
rect 403 202 404 206
rect 398 201 404 202
rect 502 206 508 207
rect 502 202 503 206
rect 507 202 508 206
rect 502 201 508 202
rect 606 206 612 207
rect 606 202 607 206
rect 611 202 612 206
rect 606 201 612 202
rect 718 206 724 207
rect 718 202 719 206
rect 723 202 724 206
rect 718 201 724 202
rect 830 206 836 207
rect 830 202 831 206
rect 835 202 836 206
rect 830 201 836 202
rect 950 206 956 207
rect 950 202 951 206
rect 955 202 956 206
rect 950 201 956 202
rect 1070 206 1076 207
rect 1070 202 1071 206
rect 1075 202 1076 206
rect 1070 201 1076 202
rect 1182 206 1188 207
rect 1182 202 1183 206
rect 1187 202 1188 206
rect 1182 201 1188 202
rect 1294 206 1300 207
rect 1294 202 1295 206
rect 1299 202 1300 206
rect 1294 201 1300 202
rect 1414 206 1420 207
rect 1414 202 1415 206
rect 1419 202 1420 206
rect 1414 201 1420 202
rect 1534 206 1540 207
rect 1534 202 1535 206
rect 1539 202 1540 206
rect 1534 201 1540 202
rect 1654 206 1660 207
rect 1654 202 1655 206
rect 1659 202 1660 206
rect 1654 201 1660 202
rect 1750 206 1756 207
rect 1750 202 1751 206
rect 1755 202 1756 206
rect 1750 201 1756 202
rect 2078 202 2084 203
rect 2078 198 2079 202
rect 2083 198 2084 202
rect 2078 197 2084 198
rect 2326 202 2332 203
rect 2326 198 2327 202
rect 2331 198 2332 202
rect 2326 197 2332 198
rect 2550 202 2556 203
rect 2550 198 2551 202
rect 2555 198 2556 202
rect 2550 197 2556 198
rect 2750 202 2756 203
rect 2750 198 2751 202
rect 2755 198 2756 202
rect 2750 197 2756 198
rect 2934 202 2940 203
rect 2934 198 2935 202
rect 2939 198 2940 202
rect 2934 197 2940 198
rect 3094 202 3100 203
rect 3094 198 3095 202
rect 3099 198 3100 202
rect 3094 197 3100 198
rect 3246 202 3252 203
rect 3246 198 3247 202
rect 3251 198 3252 202
rect 3246 197 3252 198
rect 3390 202 3396 203
rect 3390 198 3391 202
rect 3395 198 3396 202
rect 3390 197 3396 198
rect 3510 202 3516 203
rect 3510 198 3511 202
rect 3515 198 3516 202
rect 3510 197 3516 198
rect 262 150 268 151
rect 262 146 263 150
rect 267 146 268 150
rect 262 145 268 146
rect 342 150 348 151
rect 342 146 343 150
rect 347 146 348 150
rect 342 145 348 146
rect 422 150 428 151
rect 422 146 423 150
rect 427 146 428 150
rect 422 145 428 146
rect 502 150 508 151
rect 502 146 503 150
rect 507 146 508 150
rect 502 145 508 146
rect 582 150 588 151
rect 582 146 583 150
rect 587 146 588 150
rect 582 145 588 146
rect 662 150 668 151
rect 662 146 663 150
rect 667 146 668 150
rect 662 145 668 146
rect 742 150 748 151
rect 742 146 743 150
rect 747 146 748 150
rect 742 145 748 146
rect 822 150 828 151
rect 822 146 823 150
rect 827 146 828 150
rect 822 145 828 146
rect 902 150 908 151
rect 902 146 903 150
rect 907 146 908 150
rect 902 145 908 146
rect 982 150 988 151
rect 982 146 983 150
rect 987 146 988 150
rect 982 145 988 146
rect 1062 150 1068 151
rect 1062 146 1063 150
rect 1067 146 1068 150
rect 1062 145 1068 146
rect 1142 150 1148 151
rect 1142 146 1143 150
rect 1147 146 1148 150
rect 1142 145 1148 146
rect 1222 150 1228 151
rect 1222 146 1223 150
rect 1227 146 1228 150
rect 1222 145 1228 146
rect 1302 150 1308 151
rect 1302 146 1303 150
rect 1307 146 1308 150
rect 1302 145 1308 146
rect 1382 150 1388 151
rect 1382 146 1383 150
rect 1387 146 1388 150
rect 1382 145 1388 146
rect 1462 150 1468 151
rect 1462 146 1463 150
rect 1467 146 1468 150
rect 1462 145 1468 146
rect 1542 150 1548 151
rect 1542 146 1543 150
rect 1547 146 1548 150
rect 1542 145 1548 146
rect 1902 146 1908 147
rect 1902 142 1903 146
rect 1907 142 1908 146
rect 1902 141 1908 142
rect 1982 146 1988 147
rect 1982 142 1983 146
rect 1987 142 1988 146
rect 1982 141 1988 142
rect 2062 146 2068 147
rect 2062 142 2063 146
rect 2067 142 2068 146
rect 2062 141 2068 142
rect 2142 146 2148 147
rect 2142 142 2143 146
rect 2147 142 2148 146
rect 2142 141 2148 142
rect 2222 146 2228 147
rect 2222 142 2223 146
rect 2227 142 2228 146
rect 2222 141 2228 142
rect 2302 146 2308 147
rect 2302 142 2303 146
rect 2307 142 2308 146
rect 2302 141 2308 142
rect 2398 146 2404 147
rect 2398 142 2399 146
rect 2403 142 2404 146
rect 2398 141 2404 142
rect 2502 146 2508 147
rect 2502 142 2503 146
rect 2507 142 2508 146
rect 2502 141 2508 142
rect 2606 146 2612 147
rect 2606 142 2607 146
rect 2611 142 2612 146
rect 2606 141 2612 142
rect 2710 146 2716 147
rect 2710 142 2711 146
rect 2715 142 2716 146
rect 2710 141 2716 142
rect 2814 146 2820 147
rect 2814 142 2815 146
rect 2819 142 2820 146
rect 2814 141 2820 142
rect 2910 146 2916 147
rect 2910 142 2911 146
rect 2915 142 2916 146
rect 2910 141 2916 142
rect 2998 146 3004 147
rect 2998 142 2999 146
rect 3003 142 3004 146
rect 2998 141 3004 142
rect 3086 146 3092 147
rect 3086 142 3087 146
rect 3091 142 3092 146
rect 3086 141 3092 142
rect 3174 146 3180 147
rect 3174 142 3175 146
rect 3179 142 3180 146
rect 3174 141 3180 142
rect 3262 146 3268 147
rect 3262 142 3263 146
rect 3267 142 3268 146
rect 3262 141 3268 142
rect 3350 146 3356 147
rect 3350 142 3351 146
rect 3355 142 3356 146
rect 3350 141 3356 142
rect 3430 146 3436 147
rect 3430 142 3431 146
rect 3435 142 3436 146
rect 3430 141 3436 142
rect 3510 146 3516 147
rect 3510 142 3511 146
rect 3515 142 3516 146
rect 3510 141 3516 142
rect 110 132 116 133
rect 110 128 111 132
rect 115 128 116 132
rect 110 127 116 128
rect 1830 132 1836 133
rect 1830 128 1831 132
rect 1835 128 1836 132
rect 1830 127 1836 128
rect 1870 128 1876 129
rect 1870 124 1871 128
rect 1875 124 1876 128
rect 1870 123 1876 124
rect 3590 128 3596 129
rect 3590 124 3591 128
rect 3595 124 3596 128
rect 3590 123 3596 124
rect 110 115 116 116
rect 110 111 111 115
rect 115 111 116 115
rect 1830 115 1836 116
rect 110 110 116 111
rect 254 112 260 113
rect 254 108 255 112
rect 259 108 260 112
rect 254 107 260 108
rect 334 112 340 113
rect 334 108 335 112
rect 339 108 340 112
rect 334 107 340 108
rect 414 112 420 113
rect 414 108 415 112
rect 419 108 420 112
rect 414 107 420 108
rect 494 112 500 113
rect 494 108 495 112
rect 499 108 500 112
rect 494 107 500 108
rect 574 112 580 113
rect 574 108 575 112
rect 579 108 580 112
rect 574 107 580 108
rect 654 112 660 113
rect 654 108 655 112
rect 659 108 660 112
rect 654 107 660 108
rect 734 112 740 113
rect 734 108 735 112
rect 739 108 740 112
rect 734 107 740 108
rect 814 112 820 113
rect 814 108 815 112
rect 819 108 820 112
rect 814 107 820 108
rect 894 112 900 113
rect 894 108 895 112
rect 899 108 900 112
rect 894 107 900 108
rect 974 112 980 113
rect 974 108 975 112
rect 979 108 980 112
rect 974 107 980 108
rect 1054 112 1060 113
rect 1054 108 1055 112
rect 1059 108 1060 112
rect 1054 107 1060 108
rect 1134 112 1140 113
rect 1134 108 1135 112
rect 1139 108 1140 112
rect 1134 107 1140 108
rect 1214 112 1220 113
rect 1214 108 1215 112
rect 1219 108 1220 112
rect 1214 107 1220 108
rect 1294 112 1300 113
rect 1294 108 1295 112
rect 1299 108 1300 112
rect 1294 107 1300 108
rect 1374 112 1380 113
rect 1374 108 1375 112
rect 1379 108 1380 112
rect 1374 107 1380 108
rect 1454 112 1460 113
rect 1454 108 1455 112
rect 1459 108 1460 112
rect 1454 107 1460 108
rect 1534 112 1540 113
rect 1534 108 1535 112
rect 1539 108 1540 112
rect 1830 111 1831 115
rect 1835 111 1836 115
rect 1830 110 1836 111
rect 1870 111 1876 112
rect 1534 107 1540 108
rect 1870 107 1871 111
rect 1875 107 1876 111
rect 3590 111 3596 112
rect 1870 106 1876 107
rect 1894 108 1900 109
rect 1894 104 1895 108
rect 1899 104 1900 108
rect 1894 103 1900 104
rect 1974 108 1980 109
rect 1974 104 1975 108
rect 1979 104 1980 108
rect 1974 103 1980 104
rect 2054 108 2060 109
rect 2054 104 2055 108
rect 2059 104 2060 108
rect 2054 103 2060 104
rect 2134 108 2140 109
rect 2134 104 2135 108
rect 2139 104 2140 108
rect 2134 103 2140 104
rect 2214 108 2220 109
rect 2214 104 2215 108
rect 2219 104 2220 108
rect 2214 103 2220 104
rect 2294 108 2300 109
rect 2294 104 2295 108
rect 2299 104 2300 108
rect 2294 103 2300 104
rect 2390 108 2396 109
rect 2390 104 2391 108
rect 2395 104 2396 108
rect 2390 103 2396 104
rect 2494 108 2500 109
rect 2494 104 2495 108
rect 2499 104 2500 108
rect 2494 103 2500 104
rect 2598 108 2604 109
rect 2598 104 2599 108
rect 2603 104 2604 108
rect 2598 103 2604 104
rect 2702 108 2708 109
rect 2702 104 2703 108
rect 2707 104 2708 108
rect 2702 103 2708 104
rect 2806 108 2812 109
rect 2806 104 2807 108
rect 2811 104 2812 108
rect 2806 103 2812 104
rect 2902 108 2908 109
rect 2902 104 2903 108
rect 2907 104 2908 108
rect 2902 103 2908 104
rect 2990 108 2996 109
rect 2990 104 2991 108
rect 2995 104 2996 108
rect 2990 103 2996 104
rect 3078 108 3084 109
rect 3078 104 3079 108
rect 3083 104 3084 108
rect 3078 103 3084 104
rect 3166 108 3172 109
rect 3166 104 3167 108
rect 3171 104 3172 108
rect 3166 103 3172 104
rect 3254 108 3260 109
rect 3254 104 3255 108
rect 3259 104 3260 108
rect 3254 103 3260 104
rect 3342 108 3348 109
rect 3342 104 3343 108
rect 3347 104 3348 108
rect 3342 103 3348 104
rect 3422 108 3428 109
rect 3422 104 3423 108
rect 3427 104 3428 108
rect 3422 103 3428 104
rect 3502 108 3508 109
rect 3502 104 3503 108
rect 3507 104 3508 108
rect 3590 107 3591 111
rect 3595 107 3596 111
rect 3590 106 3596 107
rect 3502 103 3508 104
<< m3c >>
rect 143 3638 147 3642
rect 223 3638 227 3642
rect 351 3638 355 3642
rect 495 3638 499 3642
rect 647 3638 651 3642
rect 807 3638 811 3642
rect 975 3638 979 3642
rect 1151 3638 1155 3642
rect 1335 3638 1339 3642
rect 111 3620 115 3624
rect 1831 3620 1835 3624
rect 1927 3610 1931 3614
rect 2007 3610 2011 3614
rect 2103 3610 2107 3614
rect 2207 3610 2211 3614
rect 2319 3610 2323 3614
rect 2431 3610 2435 3614
rect 2551 3610 2555 3614
rect 2663 3610 2667 3614
rect 2775 3610 2779 3614
rect 2879 3610 2883 3614
rect 2983 3610 2987 3614
rect 3095 3610 3099 3614
rect 3207 3610 3211 3614
rect 111 3603 115 3607
rect 135 3600 139 3604
rect 215 3600 219 3604
rect 343 3600 347 3604
rect 487 3600 491 3604
rect 639 3600 643 3604
rect 799 3600 803 3604
rect 967 3600 971 3604
rect 1143 3600 1147 3604
rect 1327 3600 1331 3604
rect 1831 3603 1835 3607
rect 1871 3592 1875 3596
rect 3591 3592 3595 3596
rect 1871 3575 1875 3579
rect 1919 3572 1923 3576
rect 1999 3572 2003 3576
rect 2095 3572 2099 3576
rect 2199 3572 2203 3576
rect 2311 3572 2315 3576
rect 2423 3572 2427 3576
rect 2543 3572 2547 3576
rect 2655 3572 2659 3576
rect 2767 3572 2771 3576
rect 2871 3572 2875 3576
rect 2975 3572 2979 3576
rect 3087 3572 3091 3576
rect 3199 3572 3203 3576
rect 3591 3575 3595 3579
rect 111 3553 115 3557
rect 239 3556 243 3560
rect 359 3556 363 3560
rect 479 3556 483 3560
rect 607 3556 611 3560
rect 735 3556 739 3560
rect 863 3556 867 3560
rect 983 3556 987 3560
rect 1095 3556 1099 3560
rect 1207 3556 1211 3560
rect 1319 3556 1323 3560
rect 1439 3556 1443 3560
rect 1831 3553 1835 3557
rect 111 3536 115 3540
rect 1831 3536 1835 3540
rect 1871 3525 1875 3529
rect 1943 3528 1947 3532
rect 2127 3528 2131 3532
rect 2303 3528 2307 3532
rect 2479 3528 2483 3532
rect 2647 3528 2651 3532
rect 2815 3528 2819 3532
rect 2975 3528 2979 3532
rect 3135 3528 3139 3532
rect 3303 3528 3307 3532
rect 3591 3525 3595 3529
rect 247 3518 251 3522
rect 367 3518 371 3522
rect 487 3518 491 3522
rect 615 3518 619 3522
rect 743 3518 747 3522
rect 871 3518 875 3522
rect 991 3518 995 3522
rect 1103 3518 1107 3522
rect 1215 3518 1219 3522
rect 1327 3518 1331 3522
rect 1447 3518 1451 3522
rect 1871 3508 1875 3512
rect 3591 3508 3595 3512
rect 167 3486 171 3490
rect 287 3486 291 3490
rect 415 3486 419 3490
rect 551 3486 555 3490
rect 687 3486 691 3490
rect 823 3486 827 3490
rect 951 3486 955 3490
rect 1071 3486 1075 3490
rect 1183 3486 1187 3490
rect 1303 3486 1307 3490
rect 1423 3486 1427 3490
rect 1951 3490 1955 3494
rect 2135 3490 2139 3494
rect 2311 3490 2315 3494
rect 2487 3490 2491 3494
rect 2655 3490 2659 3494
rect 2823 3490 2827 3494
rect 2983 3490 2987 3494
rect 3143 3490 3147 3494
rect 3311 3490 3315 3494
rect 111 3468 115 3472
rect 1831 3468 1835 3472
rect 1959 3458 1963 3462
rect 2079 3458 2083 3462
rect 2199 3458 2203 3462
rect 2335 3458 2339 3462
rect 2479 3458 2483 3462
rect 2631 3458 2635 3462
rect 2791 3458 2795 3462
rect 2959 3458 2963 3462
rect 3127 3458 3131 3462
rect 3303 3458 3307 3462
rect 111 3451 115 3455
rect 159 3448 163 3452
rect 279 3448 283 3452
rect 407 3448 411 3452
rect 543 3448 547 3452
rect 679 3448 683 3452
rect 815 3448 819 3452
rect 943 3448 947 3452
rect 1063 3448 1067 3452
rect 1175 3448 1179 3452
rect 1295 3448 1299 3452
rect 1415 3448 1419 3452
rect 1831 3451 1835 3455
rect 1871 3440 1875 3444
rect 3591 3440 3595 3444
rect 1871 3423 1875 3427
rect 1951 3420 1955 3424
rect 2071 3420 2075 3424
rect 2191 3420 2195 3424
rect 2327 3420 2331 3424
rect 2471 3420 2475 3424
rect 2623 3420 2627 3424
rect 2783 3420 2787 3424
rect 2951 3420 2955 3424
rect 3119 3420 3123 3424
rect 3295 3420 3299 3424
rect 3591 3423 3595 3427
rect 111 3393 115 3397
rect 135 3396 139 3400
rect 247 3396 251 3400
rect 375 3396 379 3400
rect 503 3396 507 3400
rect 639 3396 643 3400
rect 775 3396 779 3400
rect 903 3396 907 3400
rect 1031 3396 1035 3400
rect 1159 3396 1163 3400
rect 1287 3396 1291 3400
rect 1415 3396 1419 3400
rect 1831 3393 1835 3397
rect 111 3376 115 3380
rect 1831 3376 1835 3380
rect 1871 3365 1875 3369
rect 1975 3368 1979 3372
rect 2135 3368 2139 3372
rect 2287 3368 2291 3372
rect 2431 3368 2435 3372
rect 2559 3368 2563 3372
rect 2679 3368 2683 3372
rect 2791 3368 2795 3372
rect 2895 3368 2899 3372
rect 2991 3368 2995 3372
rect 3079 3368 3083 3372
rect 3167 3368 3171 3372
rect 3255 3368 3259 3372
rect 3343 3368 3347 3372
rect 3423 3368 3427 3372
rect 3503 3368 3507 3372
rect 3591 3365 3595 3369
rect 143 3358 147 3362
rect 255 3358 259 3362
rect 383 3358 387 3362
rect 511 3358 515 3362
rect 647 3358 651 3362
rect 783 3358 787 3362
rect 911 3358 915 3362
rect 1039 3358 1043 3362
rect 1167 3358 1171 3362
rect 1295 3358 1299 3362
rect 1423 3358 1427 3362
rect 1871 3348 1875 3352
rect 3591 3348 3595 3352
rect 1983 3330 1987 3334
rect 2143 3330 2147 3334
rect 2295 3330 2299 3334
rect 2439 3330 2443 3334
rect 2567 3330 2571 3334
rect 2687 3330 2691 3334
rect 2799 3330 2803 3334
rect 2903 3330 2907 3334
rect 2999 3330 3003 3334
rect 3087 3330 3091 3334
rect 3175 3330 3179 3334
rect 3263 3330 3267 3334
rect 3351 3330 3355 3334
rect 3431 3330 3435 3334
rect 3511 3330 3515 3334
rect 271 3322 275 3326
rect 391 3322 395 3326
rect 519 3322 523 3326
rect 655 3322 659 3326
rect 791 3322 795 3326
rect 919 3322 923 3326
rect 1055 3322 1059 3326
rect 1191 3322 1195 3326
rect 1327 3322 1331 3326
rect 1463 3322 1467 3326
rect 111 3304 115 3308
rect 1831 3304 1835 3308
rect 1935 3294 1939 3298
rect 2071 3294 2075 3298
rect 2207 3294 2211 3298
rect 2367 3294 2371 3298
rect 2551 3294 2555 3298
rect 2767 3294 2771 3298
rect 3007 3294 3011 3298
rect 3255 3294 3259 3298
rect 3511 3294 3515 3298
rect 111 3287 115 3291
rect 263 3284 267 3288
rect 383 3284 387 3288
rect 511 3284 515 3288
rect 647 3284 651 3288
rect 783 3284 787 3288
rect 911 3284 915 3288
rect 1047 3284 1051 3288
rect 1183 3284 1187 3288
rect 1319 3284 1323 3288
rect 1455 3284 1459 3288
rect 1831 3287 1835 3291
rect 1871 3276 1875 3280
rect 3591 3276 3595 3280
rect 1871 3259 1875 3263
rect 1927 3256 1931 3260
rect 2063 3256 2067 3260
rect 2199 3256 2203 3260
rect 2359 3256 2363 3260
rect 2543 3256 2547 3260
rect 2759 3256 2763 3260
rect 2999 3256 3003 3260
rect 3247 3256 3251 3260
rect 3503 3256 3507 3260
rect 3591 3259 3595 3263
rect 111 3233 115 3237
rect 383 3236 387 3240
rect 471 3236 475 3240
rect 575 3236 579 3240
rect 687 3236 691 3240
rect 807 3236 811 3240
rect 935 3236 939 3240
rect 1063 3236 1067 3240
rect 1191 3236 1195 3240
rect 1319 3236 1323 3240
rect 1447 3236 1451 3240
rect 1575 3236 1579 3240
rect 1831 3233 1835 3237
rect 111 3216 115 3220
rect 1831 3216 1835 3220
rect 1871 3205 1875 3209
rect 1895 3208 1899 3212
rect 2007 3208 2011 3212
rect 2143 3208 2147 3212
rect 2279 3208 2283 3212
rect 2415 3208 2419 3212
rect 2567 3208 2571 3212
rect 2727 3208 2731 3212
rect 2911 3208 2915 3212
rect 3103 3208 3107 3212
rect 3311 3208 3315 3212
rect 3503 3208 3507 3212
rect 3591 3205 3595 3209
rect 391 3198 395 3202
rect 479 3198 483 3202
rect 583 3198 587 3202
rect 695 3198 699 3202
rect 815 3198 819 3202
rect 943 3198 947 3202
rect 1071 3198 1075 3202
rect 1199 3198 1203 3202
rect 1327 3198 1331 3202
rect 1455 3198 1459 3202
rect 1583 3198 1587 3202
rect 1871 3188 1875 3192
rect 3591 3188 3595 3192
rect 1903 3170 1907 3174
rect 2015 3170 2019 3174
rect 2151 3170 2155 3174
rect 2287 3170 2291 3174
rect 2423 3170 2427 3174
rect 2575 3170 2579 3174
rect 2735 3170 2739 3174
rect 2919 3170 2923 3174
rect 3111 3170 3115 3174
rect 3319 3170 3323 3174
rect 3511 3170 3515 3174
rect 383 3158 387 3162
rect 463 3158 467 3162
rect 543 3158 547 3162
rect 623 3158 627 3162
rect 711 3158 715 3162
rect 815 3158 819 3162
rect 927 3158 931 3162
rect 1039 3158 1043 3162
rect 1159 3158 1163 3162
rect 1271 3158 1275 3162
rect 1383 3158 1387 3162
rect 1495 3158 1499 3162
rect 1615 3158 1619 3162
rect 1735 3158 1739 3162
rect 111 3140 115 3144
rect 1831 3140 1835 3144
rect 1903 3138 1907 3142
rect 2079 3138 2083 3142
rect 2271 3138 2275 3142
rect 2455 3138 2459 3142
rect 2623 3138 2627 3142
rect 2783 3138 2787 3142
rect 2935 3138 2939 3142
rect 3079 3138 3083 3142
rect 3231 3138 3235 3142
rect 111 3123 115 3127
rect 375 3120 379 3124
rect 455 3120 459 3124
rect 535 3120 539 3124
rect 615 3120 619 3124
rect 703 3120 707 3124
rect 807 3120 811 3124
rect 919 3120 923 3124
rect 1031 3120 1035 3124
rect 1151 3120 1155 3124
rect 1263 3120 1267 3124
rect 1375 3120 1379 3124
rect 1487 3120 1491 3124
rect 1607 3120 1611 3124
rect 1727 3120 1731 3124
rect 1831 3123 1835 3127
rect 1871 3120 1875 3124
rect 3591 3120 3595 3124
rect 1871 3103 1875 3107
rect 1895 3100 1899 3104
rect 2071 3100 2075 3104
rect 2263 3100 2267 3104
rect 2447 3100 2451 3104
rect 2615 3100 2619 3104
rect 2775 3100 2779 3104
rect 2927 3100 2931 3104
rect 3071 3100 3075 3104
rect 3223 3100 3227 3104
rect 3591 3103 3595 3107
rect 111 3073 115 3077
rect 943 3076 947 3080
rect 1023 3076 1027 3080
rect 1103 3076 1107 3080
rect 1183 3076 1187 3080
rect 1263 3076 1267 3080
rect 1343 3076 1347 3080
rect 1423 3076 1427 3080
rect 1503 3076 1507 3080
rect 1583 3076 1587 3080
rect 1663 3076 1667 3080
rect 1743 3076 1747 3080
rect 1831 3073 1835 3077
rect 111 3056 115 3060
rect 1831 3056 1835 3060
rect 1871 3045 1875 3049
rect 1991 3048 1995 3052
rect 2247 3048 2251 3052
rect 2487 3048 2491 3052
rect 2703 3048 2707 3052
rect 2895 3048 2899 3052
rect 3063 3048 3067 3052
rect 3223 3048 3227 3052
rect 3375 3048 3379 3052
rect 3503 3048 3507 3052
rect 3591 3045 3595 3049
rect 951 3038 955 3042
rect 1031 3038 1035 3042
rect 1111 3038 1115 3042
rect 1191 3038 1195 3042
rect 1271 3038 1275 3042
rect 1351 3038 1355 3042
rect 1431 3038 1435 3042
rect 1511 3038 1515 3042
rect 1591 3038 1595 3042
rect 1671 3038 1675 3042
rect 1751 3038 1755 3042
rect 1871 3028 1875 3032
rect 3591 3028 3595 3032
rect 1999 3010 2003 3014
rect 2255 3010 2259 3014
rect 2495 3010 2499 3014
rect 2711 3010 2715 3014
rect 2903 3010 2907 3014
rect 3071 3010 3075 3014
rect 3231 3010 3235 3014
rect 3383 3010 3387 3014
rect 3511 3010 3515 3014
rect 207 2990 211 2994
rect 327 2990 331 2994
rect 471 2990 475 2994
rect 631 2990 635 2994
rect 807 2990 811 2994
rect 983 2990 987 2994
rect 1151 2990 1155 2994
rect 1311 2990 1315 2994
rect 1463 2990 1467 2994
rect 1615 2990 1619 2994
rect 1751 2990 1755 2994
rect 111 2972 115 2976
rect 1831 2972 1835 2976
rect 1903 2974 1907 2978
rect 2143 2974 2147 2978
rect 2391 2974 2395 2978
rect 2607 2974 2611 2978
rect 2799 2974 2803 2978
rect 2967 2974 2971 2978
rect 3119 2974 3123 2978
rect 3263 2974 3267 2978
rect 3399 2974 3403 2978
rect 3511 2974 3515 2978
rect 111 2955 115 2959
rect 199 2952 203 2956
rect 319 2952 323 2956
rect 463 2952 467 2956
rect 623 2952 627 2956
rect 799 2952 803 2956
rect 975 2952 979 2956
rect 1143 2952 1147 2956
rect 1303 2952 1307 2956
rect 1455 2952 1459 2956
rect 1607 2952 1611 2956
rect 1743 2952 1747 2956
rect 1831 2955 1835 2959
rect 1871 2956 1875 2960
rect 3591 2956 3595 2960
rect 1871 2939 1875 2943
rect 1895 2936 1899 2940
rect 2135 2936 2139 2940
rect 2383 2936 2387 2940
rect 2599 2936 2603 2940
rect 2791 2936 2795 2940
rect 2959 2936 2963 2940
rect 3111 2936 3115 2940
rect 3255 2936 3259 2940
rect 3391 2936 3395 2940
rect 3503 2936 3507 2940
rect 3591 2939 3595 2943
rect 111 2905 115 2909
rect 247 2908 251 2912
rect 351 2908 355 2912
rect 471 2908 475 2912
rect 607 2908 611 2912
rect 751 2908 755 2912
rect 895 2908 899 2912
rect 1031 2908 1035 2912
rect 1159 2908 1163 2912
rect 1279 2908 1283 2912
rect 1399 2908 1403 2912
rect 1519 2908 1523 2912
rect 1639 2908 1643 2912
rect 1831 2905 1835 2909
rect 111 2888 115 2892
rect 1831 2888 1835 2892
rect 1871 2877 1875 2881
rect 2351 2880 2355 2884
rect 2447 2880 2451 2884
rect 2551 2880 2555 2884
rect 2655 2880 2659 2884
rect 2759 2880 2763 2884
rect 2871 2880 2875 2884
rect 2983 2880 2987 2884
rect 3095 2880 3099 2884
rect 3207 2880 3211 2884
rect 3591 2877 3595 2881
rect 255 2870 259 2874
rect 359 2870 363 2874
rect 479 2870 483 2874
rect 615 2870 619 2874
rect 759 2870 763 2874
rect 903 2870 907 2874
rect 1039 2870 1043 2874
rect 1167 2870 1171 2874
rect 1287 2870 1291 2874
rect 1407 2870 1411 2874
rect 1527 2870 1531 2874
rect 1647 2870 1651 2874
rect 1871 2860 1875 2864
rect 3591 2860 3595 2864
rect 151 2838 155 2842
rect 279 2838 283 2842
rect 407 2838 411 2842
rect 543 2838 547 2842
rect 671 2838 675 2842
rect 799 2838 803 2842
rect 919 2838 923 2842
rect 1039 2838 1043 2842
rect 1151 2838 1155 2842
rect 1271 2838 1275 2842
rect 1391 2838 1395 2842
rect 2359 2842 2363 2846
rect 2455 2842 2459 2846
rect 2559 2842 2563 2846
rect 2663 2842 2667 2846
rect 2767 2842 2771 2846
rect 2879 2842 2883 2846
rect 2991 2842 2995 2846
rect 3103 2842 3107 2846
rect 3215 2842 3219 2846
rect 111 2820 115 2824
rect 1831 2820 1835 2824
rect 2239 2810 2243 2814
rect 2319 2810 2323 2814
rect 2399 2810 2403 2814
rect 2479 2810 2483 2814
rect 2567 2810 2571 2814
rect 2671 2810 2675 2814
rect 2807 2810 2811 2814
rect 2967 2810 2971 2814
rect 3143 2810 3147 2814
rect 3335 2810 3339 2814
rect 3511 2810 3515 2814
rect 111 2803 115 2807
rect 143 2800 147 2804
rect 271 2800 275 2804
rect 399 2800 403 2804
rect 535 2800 539 2804
rect 663 2800 667 2804
rect 791 2800 795 2804
rect 911 2800 915 2804
rect 1031 2800 1035 2804
rect 1143 2800 1147 2804
rect 1263 2800 1267 2804
rect 1383 2800 1387 2804
rect 1831 2803 1835 2807
rect 1871 2792 1875 2796
rect 3591 2792 3595 2796
rect 1871 2775 1875 2779
rect 2231 2772 2235 2776
rect 2311 2772 2315 2776
rect 2391 2772 2395 2776
rect 2471 2772 2475 2776
rect 2559 2772 2563 2776
rect 2663 2772 2667 2776
rect 2799 2772 2803 2776
rect 2959 2772 2963 2776
rect 3135 2772 3139 2776
rect 3327 2772 3331 2776
rect 3503 2772 3507 2776
rect 3591 2775 3595 2779
rect 111 2745 115 2749
rect 143 2748 147 2752
rect 295 2748 299 2752
rect 439 2748 443 2752
rect 567 2748 571 2752
rect 687 2748 691 2752
rect 799 2748 803 2752
rect 903 2748 907 2752
rect 1007 2748 1011 2752
rect 1103 2748 1107 2752
rect 1199 2748 1203 2752
rect 1303 2748 1307 2752
rect 1831 2745 1835 2749
rect 111 2728 115 2732
rect 1831 2728 1835 2732
rect 151 2710 155 2714
rect 303 2710 307 2714
rect 447 2710 451 2714
rect 575 2710 579 2714
rect 695 2710 699 2714
rect 807 2710 811 2714
rect 911 2710 915 2714
rect 1015 2710 1019 2714
rect 1111 2710 1115 2714
rect 1207 2710 1211 2714
rect 1311 2710 1315 2714
rect 1871 2713 1875 2717
rect 2047 2716 2051 2720
rect 2135 2716 2139 2720
rect 2231 2716 2235 2720
rect 2327 2716 2331 2720
rect 2423 2716 2427 2720
rect 2519 2716 2523 2720
rect 2615 2716 2619 2720
rect 2727 2716 2731 2720
rect 2855 2716 2859 2720
rect 3007 2716 3011 2720
rect 3175 2716 3179 2720
rect 3351 2716 3355 2720
rect 3503 2716 3507 2720
rect 3591 2713 3595 2717
rect 1871 2696 1875 2700
rect 3591 2696 3595 2700
rect 143 2674 147 2678
rect 263 2674 267 2678
rect 407 2674 411 2678
rect 543 2674 547 2678
rect 671 2674 675 2678
rect 791 2674 795 2678
rect 903 2674 907 2678
rect 1015 2674 1019 2678
rect 1119 2674 1123 2678
rect 1215 2674 1219 2678
rect 1319 2674 1323 2678
rect 1423 2674 1427 2678
rect 2055 2678 2059 2682
rect 2143 2678 2147 2682
rect 2239 2678 2243 2682
rect 2335 2678 2339 2682
rect 2431 2678 2435 2682
rect 2527 2678 2531 2682
rect 2623 2678 2627 2682
rect 2735 2678 2739 2682
rect 2863 2678 2867 2682
rect 3015 2678 3019 2682
rect 3183 2678 3187 2682
rect 3359 2678 3363 2682
rect 3511 2678 3515 2682
rect 111 2656 115 2660
rect 1831 2656 1835 2660
rect 2071 2646 2075 2650
rect 2295 2646 2299 2650
rect 2567 2646 2571 2650
rect 2871 2646 2875 2650
rect 3199 2646 3203 2650
rect 3511 2646 3515 2650
rect 111 2639 115 2643
rect 135 2636 139 2640
rect 255 2636 259 2640
rect 399 2636 403 2640
rect 535 2636 539 2640
rect 663 2636 667 2640
rect 783 2636 787 2640
rect 895 2636 899 2640
rect 1007 2636 1011 2640
rect 1111 2636 1115 2640
rect 1207 2636 1211 2640
rect 1311 2636 1315 2640
rect 1415 2636 1419 2640
rect 1831 2639 1835 2643
rect 1871 2628 1875 2632
rect 3591 2628 3595 2632
rect 1871 2611 1875 2615
rect 2063 2608 2067 2612
rect 2287 2608 2291 2612
rect 2559 2608 2563 2612
rect 2863 2608 2867 2612
rect 3191 2608 3195 2612
rect 3503 2608 3507 2612
rect 3591 2611 3595 2615
rect 111 2581 115 2585
rect 143 2584 147 2588
rect 311 2584 315 2588
rect 479 2584 483 2588
rect 639 2584 643 2588
rect 791 2584 795 2588
rect 927 2584 931 2588
rect 1055 2584 1059 2588
rect 1175 2584 1179 2588
rect 1295 2584 1299 2588
rect 1407 2584 1411 2588
rect 1527 2584 1531 2588
rect 1831 2581 1835 2585
rect 111 2564 115 2568
rect 1831 2564 1835 2568
rect 1871 2557 1875 2561
rect 2167 2560 2171 2564
rect 2263 2560 2267 2564
rect 2367 2560 2371 2564
rect 2479 2560 2483 2564
rect 2591 2560 2595 2564
rect 2695 2560 2699 2564
rect 2799 2560 2803 2564
rect 2903 2560 2907 2564
rect 3015 2560 3019 2564
rect 3135 2560 3139 2564
rect 3263 2560 3267 2564
rect 3391 2560 3395 2564
rect 3503 2560 3507 2564
rect 3591 2557 3595 2561
rect 151 2546 155 2550
rect 319 2546 323 2550
rect 487 2546 491 2550
rect 647 2546 651 2550
rect 799 2546 803 2550
rect 935 2546 939 2550
rect 1063 2546 1067 2550
rect 1183 2546 1187 2550
rect 1303 2546 1307 2550
rect 1415 2546 1419 2550
rect 1535 2546 1539 2550
rect 1871 2540 1875 2544
rect 3591 2540 3595 2544
rect 2175 2522 2179 2526
rect 2271 2522 2275 2526
rect 2375 2522 2379 2526
rect 2487 2522 2491 2526
rect 2599 2522 2603 2526
rect 2703 2522 2707 2526
rect 2807 2522 2811 2526
rect 2911 2522 2915 2526
rect 3023 2522 3027 2526
rect 3143 2522 3147 2526
rect 3271 2522 3275 2526
rect 3399 2522 3403 2526
rect 3511 2522 3515 2526
rect 143 2506 147 2510
rect 295 2506 299 2510
rect 447 2506 451 2510
rect 591 2506 595 2510
rect 735 2506 739 2510
rect 879 2506 883 2510
rect 1015 2506 1019 2510
rect 1143 2506 1147 2510
rect 1271 2506 1275 2510
rect 1399 2506 1403 2510
rect 1535 2506 1539 2510
rect 111 2488 115 2492
rect 1831 2488 1835 2492
rect 2135 2490 2139 2494
rect 2223 2490 2227 2494
rect 2319 2490 2323 2494
rect 2423 2490 2427 2494
rect 2535 2490 2539 2494
rect 2655 2490 2659 2494
rect 2783 2490 2787 2494
rect 2919 2490 2923 2494
rect 3063 2490 3067 2494
rect 3215 2490 3219 2494
rect 3375 2490 3379 2494
rect 3511 2490 3515 2494
rect 111 2471 115 2475
rect 135 2468 139 2472
rect 287 2468 291 2472
rect 439 2468 443 2472
rect 583 2468 587 2472
rect 727 2468 731 2472
rect 871 2468 875 2472
rect 1007 2468 1011 2472
rect 1135 2468 1139 2472
rect 1263 2468 1267 2472
rect 1391 2468 1395 2472
rect 1527 2468 1531 2472
rect 1831 2471 1835 2475
rect 1871 2472 1875 2476
rect 3591 2472 3595 2476
rect 1871 2455 1875 2459
rect 2127 2452 2131 2456
rect 2215 2452 2219 2456
rect 2311 2452 2315 2456
rect 2415 2452 2419 2456
rect 2527 2452 2531 2456
rect 2647 2452 2651 2456
rect 2775 2452 2779 2456
rect 2911 2452 2915 2456
rect 3055 2452 3059 2456
rect 3207 2452 3211 2456
rect 3367 2452 3371 2456
rect 3503 2452 3507 2456
rect 3591 2455 3595 2459
rect 111 2417 115 2421
rect 199 2420 203 2424
rect 351 2420 355 2424
rect 495 2420 499 2424
rect 639 2420 643 2424
rect 783 2420 787 2424
rect 919 2420 923 2424
rect 1047 2420 1051 2424
rect 1175 2420 1179 2424
rect 1311 2420 1315 2424
rect 1447 2420 1451 2424
rect 1831 2417 1835 2421
rect 111 2400 115 2404
rect 1831 2400 1835 2404
rect 1871 2397 1875 2401
rect 1975 2400 1979 2404
rect 2087 2400 2091 2404
rect 2207 2400 2211 2404
rect 2335 2400 2339 2404
rect 2479 2400 2483 2404
rect 2631 2400 2635 2404
rect 2791 2400 2795 2404
rect 2967 2400 2971 2404
rect 3151 2400 3155 2404
rect 3335 2400 3339 2404
rect 3503 2400 3507 2404
rect 3591 2397 3595 2401
rect 207 2382 211 2386
rect 359 2382 363 2386
rect 503 2382 507 2386
rect 647 2382 651 2386
rect 791 2382 795 2386
rect 927 2382 931 2386
rect 1055 2382 1059 2386
rect 1183 2382 1187 2386
rect 1319 2382 1323 2386
rect 1455 2382 1459 2386
rect 1871 2380 1875 2384
rect 3591 2380 3595 2384
rect 1983 2362 1987 2366
rect 2095 2362 2099 2366
rect 2215 2362 2219 2366
rect 2343 2362 2347 2366
rect 2487 2362 2491 2366
rect 2639 2362 2643 2366
rect 2799 2362 2803 2366
rect 2975 2362 2979 2366
rect 3159 2362 3163 2366
rect 3343 2362 3347 2366
rect 3511 2362 3515 2366
rect 223 2342 227 2346
rect 327 2342 331 2346
rect 439 2342 443 2346
rect 559 2342 563 2346
rect 679 2342 683 2346
rect 799 2342 803 2346
rect 911 2342 915 2346
rect 1023 2342 1027 2346
rect 1135 2342 1139 2346
rect 1247 2342 1251 2346
rect 1367 2342 1371 2346
rect 111 2324 115 2328
rect 1831 2324 1835 2328
rect 1903 2326 1907 2330
rect 2015 2326 2019 2330
rect 2167 2326 2171 2330
rect 2319 2326 2323 2330
rect 2471 2326 2475 2330
rect 2623 2326 2627 2330
rect 2775 2326 2779 2330
rect 2927 2326 2931 2330
rect 3087 2326 3091 2330
rect 3247 2326 3251 2330
rect 3415 2326 3419 2330
rect 111 2307 115 2311
rect 215 2304 219 2308
rect 319 2304 323 2308
rect 431 2304 435 2308
rect 551 2304 555 2308
rect 671 2304 675 2308
rect 791 2304 795 2308
rect 903 2304 907 2308
rect 1015 2304 1019 2308
rect 1127 2304 1131 2308
rect 1239 2304 1243 2308
rect 1359 2304 1363 2308
rect 1831 2307 1835 2311
rect 1871 2308 1875 2312
rect 3591 2308 3595 2312
rect 1871 2291 1875 2295
rect 1895 2288 1899 2292
rect 2007 2288 2011 2292
rect 2159 2288 2163 2292
rect 2311 2288 2315 2292
rect 2463 2288 2467 2292
rect 2615 2288 2619 2292
rect 2767 2288 2771 2292
rect 2919 2288 2923 2292
rect 3079 2288 3083 2292
rect 3239 2288 3243 2292
rect 3407 2288 3411 2292
rect 3591 2291 3595 2295
rect 111 2245 115 2249
rect 311 2248 315 2252
rect 407 2248 411 2252
rect 503 2248 507 2252
rect 607 2248 611 2252
rect 711 2248 715 2252
rect 815 2248 819 2252
rect 911 2248 915 2252
rect 1007 2248 1011 2252
rect 1103 2248 1107 2252
rect 1199 2248 1203 2252
rect 1303 2248 1307 2252
rect 1831 2245 1835 2249
rect 1871 2241 1875 2245
rect 1895 2244 1899 2248
rect 2031 2244 2035 2248
rect 2207 2244 2211 2248
rect 2391 2244 2395 2248
rect 2575 2244 2579 2248
rect 2767 2244 2771 2248
rect 2951 2244 2955 2248
rect 3143 2244 3147 2248
rect 3335 2244 3339 2248
rect 3503 2244 3507 2248
rect 3591 2241 3595 2245
rect 111 2228 115 2232
rect 1831 2228 1835 2232
rect 1871 2224 1875 2228
rect 3591 2224 3595 2228
rect 319 2210 323 2214
rect 415 2210 419 2214
rect 511 2210 515 2214
rect 615 2210 619 2214
rect 719 2210 723 2214
rect 823 2210 827 2214
rect 919 2210 923 2214
rect 1015 2210 1019 2214
rect 1111 2210 1115 2214
rect 1207 2210 1211 2214
rect 1311 2210 1315 2214
rect 1903 2206 1907 2210
rect 2039 2206 2043 2210
rect 2215 2206 2219 2210
rect 2399 2206 2403 2210
rect 2583 2206 2587 2210
rect 2775 2206 2779 2210
rect 2959 2206 2963 2210
rect 3151 2206 3155 2210
rect 3343 2206 3347 2210
rect 3511 2206 3515 2210
rect 319 2174 323 2178
rect 415 2174 419 2178
rect 519 2174 523 2178
rect 623 2174 627 2178
rect 727 2174 731 2178
rect 831 2174 835 2178
rect 935 2174 939 2178
rect 1039 2174 1043 2178
rect 1151 2174 1155 2178
rect 1263 2174 1267 2178
rect 1967 2166 1971 2170
rect 2079 2166 2083 2170
rect 2215 2166 2219 2170
rect 2367 2166 2371 2170
rect 2527 2166 2531 2170
rect 2687 2166 2691 2170
rect 2847 2166 2851 2170
rect 2991 2166 2995 2170
rect 3127 2166 3131 2170
rect 3263 2166 3267 2170
rect 3399 2166 3403 2170
rect 3511 2166 3515 2170
rect 111 2156 115 2160
rect 1831 2156 1835 2160
rect 1871 2148 1875 2152
rect 3591 2148 3595 2152
rect 111 2139 115 2143
rect 311 2136 315 2140
rect 407 2136 411 2140
rect 511 2136 515 2140
rect 615 2136 619 2140
rect 719 2136 723 2140
rect 823 2136 827 2140
rect 927 2136 931 2140
rect 1031 2136 1035 2140
rect 1143 2136 1147 2140
rect 1255 2136 1259 2140
rect 1831 2139 1835 2143
rect 1871 2131 1875 2135
rect 1959 2128 1963 2132
rect 2071 2128 2075 2132
rect 2207 2128 2211 2132
rect 2359 2128 2363 2132
rect 2519 2128 2523 2132
rect 2679 2128 2683 2132
rect 2839 2128 2843 2132
rect 2983 2128 2987 2132
rect 3119 2128 3123 2132
rect 3255 2128 3259 2132
rect 3391 2128 3395 2132
rect 3503 2128 3507 2132
rect 3591 2131 3595 2135
rect 111 2089 115 2093
rect 279 2092 283 2096
rect 399 2092 403 2096
rect 511 2092 515 2096
rect 623 2092 627 2096
rect 735 2092 739 2096
rect 847 2092 851 2096
rect 951 2092 955 2096
rect 1047 2092 1051 2096
rect 1143 2092 1147 2096
rect 1239 2092 1243 2096
rect 1343 2092 1347 2096
rect 1831 2089 1835 2093
rect 1871 2081 1875 2085
rect 2287 2084 2291 2088
rect 2391 2084 2395 2088
rect 2503 2084 2507 2088
rect 2623 2084 2627 2088
rect 2743 2084 2747 2088
rect 2855 2084 2859 2088
rect 2967 2084 2971 2088
rect 3079 2084 3083 2088
rect 3191 2084 3195 2088
rect 3303 2084 3307 2088
rect 3415 2084 3419 2088
rect 3503 2084 3507 2088
rect 3591 2081 3595 2085
rect 111 2072 115 2076
rect 1831 2072 1835 2076
rect 1871 2064 1875 2068
rect 3591 2064 3595 2068
rect 287 2054 291 2058
rect 407 2054 411 2058
rect 519 2054 523 2058
rect 631 2054 635 2058
rect 743 2054 747 2058
rect 855 2054 859 2058
rect 959 2054 963 2058
rect 1055 2054 1059 2058
rect 1151 2054 1155 2058
rect 1247 2054 1251 2058
rect 1351 2054 1355 2058
rect 2295 2046 2299 2050
rect 2399 2046 2403 2050
rect 2511 2046 2515 2050
rect 2631 2046 2635 2050
rect 2751 2046 2755 2050
rect 2863 2046 2867 2050
rect 2975 2046 2979 2050
rect 3087 2046 3091 2050
rect 3199 2046 3203 2050
rect 3311 2046 3315 2050
rect 3423 2046 3427 2050
rect 3511 2046 3515 2050
rect 183 2014 187 2018
rect 327 2014 331 2018
rect 471 2014 475 2018
rect 623 2014 627 2018
rect 767 2014 771 2018
rect 911 2014 915 2018
rect 1047 2014 1051 2018
rect 1183 2014 1187 2018
rect 1319 2014 1323 2018
rect 1463 2014 1467 2018
rect 2183 2010 2187 2014
rect 2271 2010 2275 2014
rect 2367 2010 2371 2014
rect 2463 2010 2467 2014
rect 2567 2010 2571 2014
rect 2671 2010 2675 2014
rect 2775 2010 2779 2014
rect 2879 2010 2883 2014
rect 2983 2010 2987 2014
rect 3087 2010 3091 2014
rect 3191 2010 3195 2014
rect 111 1996 115 2000
rect 1831 1996 1835 2000
rect 1871 1992 1875 1996
rect 3591 1992 3595 1996
rect 111 1979 115 1983
rect 175 1976 179 1980
rect 319 1976 323 1980
rect 463 1976 467 1980
rect 615 1976 619 1980
rect 759 1976 763 1980
rect 903 1976 907 1980
rect 1039 1976 1043 1980
rect 1175 1976 1179 1980
rect 1311 1976 1315 1980
rect 1455 1976 1459 1980
rect 1831 1979 1835 1983
rect 1871 1975 1875 1979
rect 2175 1972 2179 1976
rect 2263 1972 2267 1976
rect 2359 1972 2363 1976
rect 2455 1972 2459 1976
rect 2559 1972 2563 1976
rect 2663 1972 2667 1976
rect 2767 1972 2771 1976
rect 2871 1972 2875 1976
rect 2975 1972 2979 1976
rect 3079 1972 3083 1976
rect 3183 1972 3187 1976
rect 3591 1975 3595 1979
rect 111 1929 115 1933
rect 135 1932 139 1936
rect 295 1932 299 1936
rect 463 1932 467 1936
rect 631 1932 635 1936
rect 799 1932 803 1936
rect 951 1932 955 1936
rect 1095 1932 1099 1936
rect 1231 1932 1235 1936
rect 1359 1932 1363 1936
rect 1487 1932 1491 1936
rect 1623 1932 1627 1936
rect 1831 1929 1835 1933
rect 1871 1921 1875 1925
rect 1943 1924 1947 1928
rect 2055 1924 2059 1928
rect 2167 1924 2171 1928
rect 2287 1924 2291 1928
rect 2407 1924 2411 1928
rect 2527 1924 2531 1928
rect 2647 1924 2651 1928
rect 2775 1924 2779 1928
rect 2911 1924 2915 1928
rect 3055 1924 3059 1928
rect 3207 1924 3211 1928
rect 3367 1924 3371 1928
rect 3503 1924 3507 1928
rect 3591 1921 3595 1925
rect 111 1912 115 1916
rect 1831 1912 1835 1916
rect 1871 1904 1875 1908
rect 3591 1904 3595 1908
rect 143 1894 147 1898
rect 303 1894 307 1898
rect 471 1894 475 1898
rect 639 1894 643 1898
rect 807 1894 811 1898
rect 959 1894 963 1898
rect 1103 1894 1107 1898
rect 1239 1894 1243 1898
rect 1367 1894 1371 1898
rect 1495 1894 1499 1898
rect 1631 1894 1635 1898
rect 1951 1886 1955 1890
rect 2063 1886 2067 1890
rect 2175 1886 2179 1890
rect 2295 1886 2299 1890
rect 2415 1886 2419 1890
rect 2535 1886 2539 1890
rect 2655 1886 2659 1890
rect 2783 1886 2787 1890
rect 2919 1886 2923 1890
rect 3063 1886 3067 1890
rect 3215 1886 3219 1890
rect 3375 1886 3379 1890
rect 3511 1886 3515 1890
rect 143 1854 147 1858
rect 319 1854 323 1858
rect 519 1854 523 1858
rect 711 1854 715 1858
rect 887 1854 891 1858
rect 1055 1854 1059 1858
rect 1207 1854 1211 1858
rect 1343 1854 1347 1858
rect 1471 1854 1475 1858
rect 1599 1854 1603 1858
rect 1727 1854 1731 1858
rect 1903 1850 1907 1854
rect 1983 1850 1987 1854
rect 2095 1850 2099 1854
rect 2207 1850 2211 1854
rect 2327 1850 2331 1854
rect 2463 1850 2467 1854
rect 2631 1850 2635 1854
rect 2831 1850 2835 1854
rect 3055 1850 3059 1854
rect 3295 1850 3299 1854
rect 3511 1850 3515 1854
rect 111 1836 115 1840
rect 1831 1836 1835 1840
rect 1871 1832 1875 1836
rect 3591 1832 3595 1836
rect 111 1819 115 1823
rect 135 1816 139 1820
rect 311 1816 315 1820
rect 511 1816 515 1820
rect 703 1816 707 1820
rect 879 1816 883 1820
rect 1047 1816 1051 1820
rect 1199 1816 1203 1820
rect 1335 1816 1339 1820
rect 1463 1816 1467 1820
rect 1591 1816 1595 1820
rect 1719 1816 1723 1820
rect 1831 1819 1835 1823
rect 1871 1815 1875 1819
rect 1895 1812 1899 1816
rect 1975 1812 1979 1816
rect 2087 1812 2091 1816
rect 2199 1812 2203 1816
rect 2319 1812 2323 1816
rect 2455 1812 2459 1816
rect 2623 1812 2627 1816
rect 2823 1812 2827 1816
rect 3047 1812 3051 1816
rect 3287 1812 3291 1816
rect 3503 1812 3507 1816
rect 3591 1815 3595 1819
rect 111 1769 115 1773
rect 135 1772 139 1776
rect 311 1772 315 1776
rect 503 1772 507 1776
rect 687 1772 691 1776
rect 847 1772 851 1776
rect 991 1772 995 1776
rect 1127 1772 1131 1776
rect 1247 1772 1251 1776
rect 1359 1772 1363 1776
rect 1463 1772 1467 1776
rect 1559 1772 1563 1776
rect 1663 1772 1667 1776
rect 1743 1772 1747 1776
rect 1831 1769 1835 1773
rect 111 1752 115 1756
rect 1831 1752 1835 1756
rect 1871 1749 1875 1753
rect 1895 1752 1899 1756
rect 2023 1752 2027 1756
rect 2183 1752 2187 1756
rect 2351 1752 2355 1756
rect 2551 1752 2555 1756
rect 2775 1752 2779 1756
rect 3015 1752 3019 1756
rect 3271 1752 3275 1756
rect 3503 1752 3507 1756
rect 3591 1749 3595 1753
rect 143 1734 147 1738
rect 319 1734 323 1738
rect 511 1734 515 1738
rect 695 1734 699 1738
rect 855 1734 859 1738
rect 999 1734 1003 1738
rect 1135 1734 1139 1738
rect 1255 1734 1259 1738
rect 1367 1734 1371 1738
rect 1471 1734 1475 1738
rect 1567 1734 1571 1738
rect 1671 1734 1675 1738
rect 1751 1734 1755 1738
rect 1871 1732 1875 1736
rect 3591 1732 3595 1736
rect 1903 1714 1907 1718
rect 2031 1714 2035 1718
rect 2191 1714 2195 1718
rect 2359 1714 2363 1718
rect 2559 1714 2563 1718
rect 2783 1714 2787 1718
rect 3023 1714 3027 1718
rect 3279 1714 3283 1718
rect 3511 1714 3515 1718
rect 143 1694 147 1698
rect 239 1694 243 1698
rect 367 1694 371 1698
rect 487 1694 491 1698
rect 607 1694 611 1698
rect 719 1694 723 1698
rect 823 1694 827 1698
rect 927 1694 931 1698
rect 1023 1694 1027 1698
rect 1119 1694 1123 1698
rect 1215 1694 1219 1698
rect 1319 1694 1323 1698
rect 1903 1682 1907 1686
rect 1991 1682 1995 1686
rect 2111 1682 2115 1686
rect 2231 1682 2235 1686
rect 2351 1682 2355 1686
rect 2479 1682 2483 1686
rect 2607 1682 2611 1686
rect 2743 1682 2747 1686
rect 2887 1682 2891 1686
rect 3039 1682 3043 1686
rect 3199 1682 3203 1686
rect 3367 1682 3371 1686
rect 3511 1682 3515 1686
rect 111 1676 115 1680
rect 1831 1676 1835 1680
rect 1871 1664 1875 1668
rect 111 1659 115 1663
rect 3591 1664 3595 1668
rect 135 1656 139 1660
rect 231 1656 235 1660
rect 359 1656 363 1660
rect 479 1656 483 1660
rect 599 1656 603 1660
rect 711 1656 715 1660
rect 815 1656 819 1660
rect 919 1656 923 1660
rect 1015 1656 1019 1660
rect 1111 1656 1115 1660
rect 1207 1656 1211 1660
rect 1311 1656 1315 1660
rect 1831 1659 1835 1663
rect 1871 1647 1875 1651
rect 1895 1644 1899 1648
rect 1983 1644 1987 1648
rect 2103 1644 2107 1648
rect 2223 1644 2227 1648
rect 2343 1644 2347 1648
rect 2471 1644 2475 1648
rect 2599 1644 2603 1648
rect 2735 1644 2739 1648
rect 2879 1644 2883 1648
rect 3031 1644 3035 1648
rect 3191 1644 3195 1648
rect 3359 1644 3363 1648
rect 3503 1644 3507 1648
rect 3591 1647 3595 1651
rect 111 1601 115 1605
rect 175 1604 179 1608
rect 311 1604 315 1608
rect 439 1604 443 1608
rect 567 1604 571 1608
rect 687 1604 691 1608
rect 799 1604 803 1608
rect 903 1604 907 1608
rect 999 1604 1003 1608
rect 1095 1604 1099 1608
rect 1199 1604 1203 1608
rect 1303 1604 1307 1608
rect 1831 1601 1835 1605
rect 1871 1597 1875 1601
rect 1927 1600 1931 1604
rect 2023 1600 2027 1604
rect 2135 1600 2139 1604
rect 2263 1600 2267 1604
rect 2391 1600 2395 1604
rect 2527 1600 2531 1604
rect 2671 1600 2675 1604
rect 2823 1600 2827 1604
rect 2983 1600 2987 1604
rect 3159 1600 3163 1604
rect 3343 1600 3347 1604
rect 3503 1600 3507 1604
rect 3591 1597 3595 1601
rect 111 1584 115 1588
rect 1831 1584 1835 1588
rect 1871 1580 1875 1584
rect 3591 1580 3595 1584
rect 183 1566 187 1570
rect 319 1566 323 1570
rect 447 1566 451 1570
rect 575 1566 579 1570
rect 695 1566 699 1570
rect 807 1566 811 1570
rect 911 1566 915 1570
rect 1007 1566 1011 1570
rect 1103 1566 1107 1570
rect 1207 1566 1211 1570
rect 1311 1566 1315 1570
rect 1935 1562 1939 1566
rect 2031 1562 2035 1566
rect 2143 1562 2147 1566
rect 2271 1562 2275 1566
rect 2399 1562 2403 1566
rect 2535 1562 2539 1566
rect 2679 1562 2683 1566
rect 2831 1562 2835 1566
rect 2991 1562 2995 1566
rect 3167 1562 3171 1566
rect 3351 1562 3355 1566
rect 3511 1562 3515 1566
rect 239 1526 243 1530
rect 343 1526 347 1530
rect 463 1526 467 1530
rect 591 1526 595 1530
rect 719 1526 723 1530
rect 855 1526 859 1530
rect 983 1526 987 1530
rect 1111 1526 1115 1530
rect 1231 1526 1235 1530
rect 1343 1526 1347 1530
rect 1455 1526 1459 1530
rect 1575 1526 1579 1530
rect 2135 1522 2139 1526
rect 2255 1522 2259 1526
rect 2383 1522 2387 1526
rect 2511 1522 2515 1526
rect 2639 1522 2643 1526
rect 2767 1522 2771 1526
rect 2887 1522 2891 1526
rect 3007 1522 3011 1526
rect 3119 1522 3123 1526
rect 3231 1522 3235 1526
rect 3351 1522 3355 1526
rect 111 1508 115 1512
rect 1831 1508 1835 1512
rect 1871 1504 1875 1508
rect 3591 1504 3595 1508
rect 111 1491 115 1495
rect 231 1488 235 1492
rect 335 1488 339 1492
rect 455 1488 459 1492
rect 583 1488 587 1492
rect 711 1488 715 1492
rect 847 1488 851 1492
rect 975 1488 979 1492
rect 1103 1488 1107 1492
rect 1223 1488 1227 1492
rect 1335 1488 1339 1492
rect 1447 1488 1451 1492
rect 1567 1488 1571 1492
rect 1831 1491 1835 1495
rect 1871 1487 1875 1491
rect 2127 1484 2131 1488
rect 2247 1484 2251 1488
rect 2375 1484 2379 1488
rect 2503 1484 2507 1488
rect 2631 1484 2635 1488
rect 2759 1484 2763 1488
rect 2879 1484 2883 1488
rect 2999 1484 3003 1488
rect 3111 1484 3115 1488
rect 3223 1484 3227 1488
rect 3343 1484 3347 1488
rect 3591 1487 3595 1491
rect 111 1429 115 1433
rect 279 1432 283 1436
rect 383 1432 387 1436
rect 511 1432 515 1436
rect 655 1432 659 1436
rect 807 1432 811 1436
rect 959 1432 963 1436
rect 1111 1432 1115 1436
rect 1247 1432 1251 1436
rect 1383 1432 1387 1436
rect 1511 1432 1515 1436
rect 1639 1432 1643 1436
rect 1743 1432 1747 1436
rect 1831 1429 1835 1433
rect 1871 1429 1875 1433
rect 2247 1432 2251 1436
rect 2343 1432 2347 1436
rect 2455 1432 2459 1436
rect 2575 1432 2579 1436
rect 2703 1432 2707 1436
rect 2831 1432 2835 1436
rect 2951 1432 2955 1436
rect 3071 1432 3075 1436
rect 3183 1432 3187 1436
rect 3295 1432 3299 1436
rect 3407 1432 3411 1436
rect 3503 1432 3507 1436
rect 3591 1429 3595 1433
rect 111 1412 115 1416
rect 1831 1412 1835 1416
rect 1871 1412 1875 1416
rect 3591 1412 3595 1416
rect 287 1394 291 1398
rect 391 1394 395 1398
rect 519 1394 523 1398
rect 663 1394 667 1398
rect 815 1394 819 1398
rect 967 1394 971 1398
rect 1119 1394 1123 1398
rect 1255 1394 1259 1398
rect 1391 1394 1395 1398
rect 1519 1394 1523 1398
rect 1647 1394 1651 1398
rect 1751 1394 1755 1398
rect 2255 1394 2259 1398
rect 2351 1394 2355 1398
rect 2463 1394 2467 1398
rect 2583 1394 2587 1398
rect 2711 1394 2715 1398
rect 2839 1394 2843 1398
rect 2959 1394 2963 1398
rect 3079 1394 3083 1398
rect 3191 1394 3195 1398
rect 3303 1394 3307 1398
rect 3415 1394 3419 1398
rect 3511 1394 3515 1398
rect 2399 1354 2403 1358
rect 2503 1354 2507 1358
rect 2615 1354 2619 1358
rect 2735 1354 2739 1358
rect 2847 1354 2851 1358
rect 2959 1354 2963 1358
rect 3071 1354 3075 1358
rect 3183 1354 3187 1358
rect 3295 1354 3299 1358
rect 3415 1354 3419 1358
rect 223 1346 227 1350
rect 335 1346 339 1350
rect 471 1346 475 1350
rect 623 1346 627 1350
rect 783 1346 787 1350
rect 943 1346 947 1350
rect 1095 1346 1099 1350
rect 1239 1346 1243 1350
rect 1375 1346 1379 1350
rect 1511 1346 1515 1350
rect 1639 1346 1643 1350
rect 1751 1346 1755 1350
rect 1871 1336 1875 1340
rect 3591 1336 3595 1340
rect 111 1328 115 1332
rect 1831 1328 1835 1332
rect 1871 1319 1875 1323
rect 2391 1316 2395 1320
rect 111 1311 115 1315
rect 2495 1316 2499 1320
rect 2607 1316 2611 1320
rect 2727 1316 2731 1320
rect 2839 1316 2843 1320
rect 2951 1316 2955 1320
rect 3063 1316 3067 1320
rect 3175 1316 3179 1320
rect 3287 1316 3291 1320
rect 3407 1316 3411 1320
rect 3591 1319 3595 1323
rect 215 1308 219 1312
rect 327 1308 331 1312
rect 463 1308 467 1312
rect 615 1308 619 1312
rect 775 1308 779 1312
rect 935 1308 939 1312
rect 1087 1308 1091 1312
rect 1231 1308 1235 1312
rect 1367 1308 1371 1312
rect 1503 1308 1507 1312
rect 1631 1308 1635 1312
rect 1743 1308 1747 1312
rect 1831 1311 1835 1315
rect 111 1261 115 1265
rect 135 1264 139 1268
rect 215 1264 219 1268
rect 335 1264 339 1268
rect 463 1264 467 1268
rect 607 1264 611 1268
rect 751 1264 755 1268
rect 903 1264 907 1268
rect 1047 1264 1051 1268
rect 1183 1264 1187 1268
rect 1303 1264 1307 1268
rect 1423 1264 1427 1268
rect 1535 1264 1539 1268
rect 1647 1264 1651 1268
rect 1743 1264 1747 1268
rect 1831 1261 1835 1265
rect 1871 1253 1875 1257
rect 1895 1256 1899 1260
rect 2071 1256 2075 1260
rect 2255 1256 2259 1260
rect 2423 1256 2427 1260
rect 2583 1256 2587 1260
rect 2735 1256 2739 1260
rect 2879 1256 2883 1260
rect 3015 1256 3019 1260
rect 3143 1256 3147 1260
rect 3271 1256 3275 1260
rect 3399 1256 3403 1260
rect 3503 1256 3507 1260
rect 3591 1253 3595 1257
rect 111 1244 115 1248
rect 1831 1244 1835 1248
rect 1871 1236 1875 1240
rect 3591 1236 3595 1240
rect 143 1226 147 1230
rect 223 1226 227 1230
rect 343 1226 347 1230
rect 471 1226 475 1230
rect 615 1226 619 1230
rect 759 1226 763 1230
rect 911 1226 915 1230
rect 1055 1226 1059 1230
rect 1191 1226 1195 1230
rect 1311 1226 1315 1230
rect 1431 1226 1435 1230
rect 1543 1226 1547 1230
rect 1655 1226 1659 1230
rect 1751 1226 1755 1230
rect 1903 1218 1907 1222
rect 2079 1218 2083 1222
rect 2263 1218 2267 1222
rect 2431 1218 2435 1222
rect 2591 1218 2595 1222
rect 2743 1218 2747 1222
rect 2887 1218 2891 1222
rect 3023 1218 3027 1222
rect 3151 1218 3155 1222
rect 3279 1218 3283 1222
rect 3407 1218 3411 1222
rect 3511 1218 3515 1222
rect 143 1182 147 1186
rect 255 1182 259 1186
rect 383 1182 387 1186
rect 503 1182 507 1186
rect 615 1182 619 1186
rect 719 1182 723 1186
rect 815 1182 819 1186
rect 911 1182 915 1186
rect 999 1182 1003 1186
rect 1095 1182 1099 1186
rect 1191 1182 1195 1186
rect 1287 1182 1291 1186
rect 1903 1178 1907 1182
rect 1991 1178 1995 1182
rect 2103 1178 2107 1182
rect 2215 1178 2219 1182
rect 2327 1178 2331 1182
rect 2447 1178 2451 1182
rect 2575 1178 2579 1182
rect 2719 1178 2723 1182
rect 2871 1178 2875 1182
rect 3031 1178 3035 1182
rect 3191 1178 3195 1182
rect 3359 1178 3363 1182
rect 3511 1178 3515 1182
rect 111 1164 115 1168
rect 1831 1164 1835 1168
rect 1871 1160 1875 1164
rect 3591 1160 3595 1164
rect 111 1147 115 1151
rect 135 1144 139 1148
rect 247 1144 251 1148
rect 375 1144 379 1148
rect 495 1144 499 1148
rect 607 1144 611 1148
rect 711 1144 715 1148
rect 807 1144 811 1148
rect 903 1144 907 1148
rect 991 1144 995 1148
rect 1087 1144 1091 1148
rect 1183 1144 1187 1148
rect 1279 1144 1283 1148
rect 1831 1147 1835 1151
rect 1871 1143 1875 1147
rect 1895 1140 1899 1144
rect 1983 1140 1987 1144
rect 2095 1140 2099 1144
rect 2207 1140 2211 1144
rect 2319 1140 2323 1144
rect 2439 1140 2443 1144
rect 2567 1140 2571 1144
rect 2711 1140 2715 1144
rect 2863 1140 2867 1144
rect 3023 1140 3027 1144
rect 3183 1140 3187 1144
rect 3351 1140 3355 1144
rect 3503 1140 3507 1144
rect 3591 1143 3595 1147
rect 111 1085 115 1089
rect 135 1088 139 1092
rect 255 1088 259 1092
rect 399 1088 403 1092
rect 535 1088 539 1092
rect 663 1088 667 1092
rect 783 1088 787 1092
rect 895 1088 899 1092
rect 999 1088 1003 1092
rect 1095 1088 1099 1092
rect 1191 1088 1195 1092
rect 1295 1088 1299 1092
rect 1399 1088 1403 1092
rect 1831 1085 1835 1089
rect 1871 1085 1875 1089
rect 1967 1088 1971 1092
rect 2047 1088 2051 1092
rect 2135 1088 2139 1092
rect 2231 1088 2235 1092
rect 2335 1088 2339 1092
rect 2439 1088 2443 1092
rect 2551 1088 2555 1092
rect 2679 1088 2683 1092
rect 2823 1088 2827 1092
rect 2983 1088 2987 1092
rect 3159 1088 3163 1092
rect 3343 1088 3347 1092
rect 3503 1088 3507 1092
rect 3591 1085 3595 1089
rect 111 1068 115 1072
rect 1831 1068 1835 1072
rect 1871 1068 1875 1072
rect 3591 1068 3595 1072
rect 143 1050 147 1054
rect 263 1050 267 1054
rect 407 1050 411 1054
rect 543 1050 547 1054
rect 671 1050 675 1054
rect 791 1050 795 1054
rect 903 1050 907 1054
rect 1007 1050 1011 1054
rect 1103 1050 1107 1054
rect 1199 1050 1203 1054
rect 1303 1050 1307 1054
rect 1407 1050 1411 1054
rect 1975 1050 1979 1054
rect 2055 1050 2059 1054
rect 2143 1050 2147 1054
rect 2239 1050 2243 1054
rect 2343 1050 2347 1054
rect 2447 1050 2451 1054
rect 2559 1050 2563 1054
rect 2687 1050 2691 1054
rect 2831 1050 2835 1054
rect 2991 1050 2995 1054
rect 3167 1050 3171 1054
rect 3351 1050 3355 1054
rect 3511 1050 3515 1054
rect 143 1010 147 1014
rect 271 1010 275 1014
rect 423 1010 427 1014
rect 583 1010 587 1014
rect 735 1010 739 1014
rect 887 1010 891 1014
rect 1031 1010 1035 1014
rect 1159 1010 1163 1014
rect 1279 1010 1283 1014
rect 1399 1010 1403 1014
rect 1519 1010 1523 1014
rect 1639 1010 1643 1014
rect 2031 1010 2035 1014
rect 2127 1010 2131 1014
rect 2231 1010 2235 1014
rect 2351 1010 2355 1014
rect 2471 1010 2475 1014
rect 2599 1010 2603 1014
rect 2727 1010 2731 1014
rect 2855 1010 2859 1014
rect 2983 1010 2987 1014
rect 3111 1010 3115 1014
rect 3247 1010 3251 1014
rect 3391 1010 3395 1014
rect 3511 1010 3515 1014
rect 111 992 115 996
rect 1831 992 1835 996
rect 1871 992 1875 996
rect 3591 992 3595 996
rect 111 975 115 979
rect 135 972 139 976
rect 263 972 267 976
rect 415 972 419 976
rect 575 972 579 976
rect 727 972 731 976
rect 879 972 883 976
rect 1023 972 1027 976
rect 1151 972 1155 976
rect 1271 972 1275 976
rect 1391 972 1395 976
rect 1511 972 1515 976
rect 1631 972 1635 976
rect 1831 975 1835 979
rect 1871 975 1875 979
rect 2023 972 2027 976
rect 2119 972 2123 976
rect 2223 972 2227 976
rect 2343 972 2347 976
rect 2463 972 2467 976
rect 2591 972 2595 976
rect 2719 972 2723 976
rect 2847 972 2851 976
rect 2975 972 2979 976
rect 3103 972 3107 976
rect 3239 972 3243 976
rect 3383 972 3387 976
rect 3503 972 3507 976
rect 3591 975 3595 979
rect 111 917 115 921
rect 135 920 139 924
rect 215 920 219 924
rect 335 920 339 924
rect 463 920 467 924
rect 599 920 603 924
rect 735 920 739 924
rect 863 920 867 924
rect 991 920 995 924
rect 1111 920 1115 924
rect 1223 920 1227 924
rect 1335 920 1339 924
rect 1455 920 1459 924
rect 1831 917 1835 921
rect 1871 917 1875 921
rect 1895 920 1899 924
rect 1983 920 1987 924
rect 2111 920 2115 924
rect 2263 920 2267 924
rect 2423 920 2427 924
rect 2583 920 2587 924
rect 2735 920 2739 924
rect 2879 920 2883 924
rect 3015 920 3019 924
rect 3143 920 3147 924
rect 3271 920 3275 924
rect 3399 920 3403 924
rect 3503 920 3507 924
rect 3591 917 3595 921
rect 111 900 115 904
rect 1831 900 1835 904
rect 1871 900 1875 904
rect 3591 900 3595 904
rect 143 882 147 886
rect 223 882 227 886
rect 343 882 347 886
rect 471 882 475 886
rect 607 882 611 886
rect 743 882 747 886
rect 871 882 875 886
rect 999 882 1003 886
rect 1119 882 1123 886
rect 1231 882 1235 886
rect 1343 882 1347 886
rect 1463 882 1467 886
rect 1903 882 1907 886
rect 1991 882 1995 886
rect 2119 882 2123 886
rect 2271 882 2275 886
rect 2431 882 2435 886
rect 2591 882 2595 886
rect 2743 882 2747 886
rect 2887 882 2891 886
rect 3023 882 3027 886
rect 3151 882 3155 886
rect 3279 882 3283 886
rect 3407 882 3411 886
rect 3511 882 3515 886
rect 143 838 147 842
rect 223 838 227 842
rect 303 838 307 842
rect 391 838 395 842
rect 495 838 499 842
rect 599 838 603 842
rect 711 838 715 842
rect 839 838 843 842
rect 991 838 995 842
rect 1167 838 1171 842
rect 1359 838 1363 842
rect 1567 838 1571 842
rect 1751 838 1755 842
rect 1903 842 1907 846
rect 2039 842 2043 846
rect 2215 842 2219 846
rect 2391 842 2395 846
rect 2567 842 2571 846
rect 2735 842 2739 846
rect 2887 842 2891 846
rect 3031 842 3035 846
rect 3159 842 3163 846
rect 3287 842 3291 846
rect 3407 842 3411 846
rect 3511 842 3515 846
rect 111 820 115 824
rect 1831 820 1835 824
rect 1871 824 1875 828
rect 3591 824 3595 828
rect 111 803 115 807
rect 135 800 139 804
rect 215 800 219 804
rect 295 800 299 804
rect 383 800 387 804
rect 487 800 491 804
rect 591 800 595 804
rect 703 800 707 804
rect 831 800 835 804
rect 983 800 987 804
rect 1159 800 1163 804
rect 1351 800 1355 804
rect 1559 800 1563 804
rect 1743 800 1747 804
rect 1831 803 1835 807
rect 1871 807 1875 811
rect 1895 804 1899 808
rect 2031 804 2035 808
rect 2207 804 2211 808
rect 2383 804 2387 808
rect 2559 804 2563 808
rect 2727 804 2731 808
rect 2879 804 2883 808
rect 3023 804 3027 808
rect 3151 804 3155 808
rect 3279 804 3283 808
rect 3399 804 3403 808
rect 3503 804 3507 808
rect 3591 807 3595 811
rect 111 749 115 753
rect 199 752 203 756
rect 287 752 291 756
rect 391 752 395 756
rect 503 752 507 756
rect 615 752 619 756
rect 735 752 739 756
rect 855 752 859 756
rect 983 752 987 756
rect 1111 752 1115 756
rect 1239 752 1243 756
rect 1367 752 1371 756
rect 1495 752 1499 756
rect 1631 752 1635 756
rect 1743 752 1747 756
rect 1831 749 1835 753
rect 1871 741 1875 745
rect 2023 744 2027 748
rect 2191 744 2195 748
rect 2359 744 2363 748
rect 2519 744 2523 748
rect 2679 744 2683 748
rect 2831 744 2835 748
rect 2975 744 2979 748
rect 3111 744 3115 748
rect 3247 744 3251 748
rect 3383 744 3387 748
rect 3503 744 3507 748
rect 3591 741 3595 745
rect 111 732 115 736
rect 1831 732 1835 736
rect 1871 724 1875 728
rect 3591 724 3595 728
rect 207 714 211 718
rect 295 714 299 718
rect 399 714 403 718
rect 511 714 515 718
rect 623 714 627 718
rect 743 714 747 718
rect 863 714 867 718
rect 991 714 995 718
rect 1119 714 1123 718
rect 1247 714 1251 718
rect 1375 714 1379 718
rect 1503 714 1507 718
rect 1639 714 1643 718
rect 1751 714 1755 718
rect 2031 706 2035 710
rect 2199 706 2203 710
rect 2367 706 2371 710
rect 2527 706 2531 710
rect 2687 706 2691 710
rect 2839 706 2843 710
rect 2983 706 2987 710
rect 3119 706 3123 710
rect 3255 706 3259 710
rect 3391 706 3395 710
rect 3511 706 3515 710
rect 383 666 387 670
rect 479 666 483 670
rect 591 666 595 670
rect 719 666 723 670
rect 855 666 859 670
rect 991 666 995 670
rect 1127 666 1131 670
rect 1255 666 1259 670
rect 1383 666 1387 670
rect 1503 666 1507 670
rect 1631 666 1635 670
rect 1751 666 1755 670
rect 2095 670 2099 674
rect 2175 670 2179 674
rect 2263 670 2267 674
rect 2359 670 2363 674
rect 2463 670 2467 674
rect 2567 670 2571 674
rect 2679 670 2683 674
rect 2799 670 2803 674
rect 2927 670 2931 674
rect 3071 670 3075 674
rect 3223 670 3227 674
rect 3375 670 3379 674
rect 3511 670 3515 674
rect 111 648 115 652
rect 1831 648 1835 652
rect 1871 652 1875 656
rect 3591 652 3595 656
rect 111 631 115 635
rect 375 628 379 632
rect 471 628 475 632
rect 583 628 587 632
rect 711 628 715 632
rect 847 628 851 632
rect 983 628 987 632
rect 1119 628 1123 632
rect 1247 628 1251 632
rect 1375 628 1379 632
rect 1495 628 1499 632
rect 1623 628 1627 632
rect 1743 628 1747 632
rect 1831 631 1835 635
rect 1871 635 1875 639
rect 2087 632 2091 636
rect 2167 632 2171 636
rect 2255 632 2259 636
rect 2351 632 2355 636
rect 2455 632 2459 636
rect 2559 632 2563 636
rect 2671 632 2675 636
rect 2791 632 2795 636
rect 2919 632 2923 636
rect 3063 632 3067 636
rect 3215 632 3219 636
rect 3367 632 3371 636
rect 3503 632 3507 636
rect 3591 635 3595 639
rect 111 573 115 577
rect 599 576 603 580
rect 687 576 691 580
rect 783 576 787 580
rect 887 576 891 580
rect 991 576 995 580
rect 1095 576 1099 580
rect 1199 576 1203 580
rect 1303 576 1307 580
rect 1399 576 1403 580
rect 1503 576 1507 580
rect 1607 576 1611 580
rect 1711 576 1715 580
rect 1831 573 1835 577
rect 1871 573 1875 577
rect 2167 576 2171 580
rect 2247 576 2251 580
rect 2327 576 2331 580
rect 2407 576 2411 580
rect 2487 576 2491 580
rect 2567 576 2571 580
rect 2647 576 2651 580
rect 2743 576 2747 580
rect 2863 576 2867 580
rect 2999 576 3003 580
rect 3159 576 3163 580
rect 3327 576 3331 580
rect 3495 576 3499 580
rect 3591 573 3595 577
rect 111 556 115 560
rect 1831 556 1835 560
rect 1871 556 1875 560
rect 3591 556 3595 560
rect 607 538 611 542
rect 695 538 699 542
rect 791 538 795 542
rect 895 538 899 542
rect 999 538 1003 542
rect 1103 538 1107 542
rect 1207 538 1211 542
rect 1311 538 1315 542
rect 1407 538 1411 542
rect 1511 538 1515 542
rect 1615 538 1619 542
rect 1719 538 1723 542
rect 2175 538 2179 542
rect 2255 538 2259 542
rect 2335 538 2339 542
rect 2415 538 2419 542
rect 2495 538 2499 542
rect 2575 538 2579 542
rect 2655 538 2659 542
rect 2751 538 2755 542
rect 2871 538 2875 542
rect 3007 538 3011 542
rect 3167 538 3171 542
rect 3335 538 3339 542
rect 3503 538 3507 542
rect 367 498 371 502
rect 463 498 467 502
rect 575 498 579 502
rect 703 498 707 502
rect 839 498 843 502
rect 975 498 979 502
rect 1111 498 1115 502
rect 1239 498 1243 502
rect 1359 498 1363 502
rect 1471 498 1475 502
rect 1583 498 1587 502
rect 1703 498 1707 502
rect 2159 498 2163 502
rect 2239 498 2243 502
rect 2319 498 2323 502
rect 2399 498 2403 502
rect 2479 498 2483 502
rect 2559 498 2563 502
rect 2639 498 2643 502
rect 2735 498 2739 502
rect 2855 498 2859 502
rect 2991 498 2995 502
rect 3143 498 3147 502
rect 3311 498 3315 502
rect 3479 498 3483 502
rect 111 480 115 484
rect 1831 480 1835 484
rect 1871 480 1875 484
rect 3591 480 3595 484
rect 111 463 115 467
rect 359 460 363 464
rect 455 460 459 464
rect 567 460 571 464
rect 695 460 699 464
rect 831 460 835 464
rect 967 460 971 464
rect 1103 460 1107 464
rect 1231 460 1235 464
rect 1351 460 1355 464
rect 1463 460 1467 464
rect 1575 460 1579 464
rect 1695 460 1699 464
rect 1831 463 1835 467
rect 1871 463 1875 467
rect 2151 460 2155 464
rect 2231 460 2235 464
rect 2311 460 2315 464
rect 2391 460 2395 464
rect 2471 460 2475 464
rect 2551 460 2555 464
rect 2631 460 2635 464
rect 2727 460 2731 464
rect 2847 460 2851 464
rect 2983 460 2987 464
rect 3135 460 3139 464
rect 3303 460 3307 464
rect 3471 460 3475 464
rect 3591 463 3595 467
rect 111 401 115 405
rect 135 404 139 408
rect 223 404 227 408
rect 359 404 363 408
rect 511 404 515 408
rect 679 404 683 408
rect 839 404 843 408
rect 999 404 1003 408
rect 1143 404 1147 408
rect 1279 404 1283 408
rect 1415 404 1419 408
rect 1551 404 1555 408
rect 1687 404 1691 408
rect 1831 401 1835 405
rect 1871 401 1875 405
rect 2159 404 2163 408
rect 2239 404 2243 408
rect 2319 404 2323 408
rect 2399 404 2403 408
rect 2479 404 2483 408
rect 2559 404 2563 408
rect 2639 404 2643 408
rect 2735 404 2739 408
rect 2839 404 2843 408
rect 2959 404 2963 408
rect 3087 404 3091 408
rect 3231 404 3235 408
rect 3375 404 3379 408
rect 3503 404 3507 408
rect 3591 401 3595 405
rect 111 384 115 388
rect 1831 384 1835 388
rect 1871 384 1875 388
rect 3591 384 3595 388
rect 143 366 147 370
rect 231 366 235 370
rect 367 366 371 370
rect 519 366 523 370
rect 687 366 691 370
rect 847 366 851 370
rect 1007 366 1011 370
rect 1151 366 1155 370
rect 1287 366 1291 370
rect 1423 366 1427 370
rect 1559 366 1563 370
rect 1695 366 1699 370
rect 2167 366 2171 370
rect 2247 366 2251 370
rect 2327 366 2331 370
rect 2407 366 2411 370
rect 2487 366 2491 370
rect 2567 366 2571 370
rect 2647 366 2651 370
rect 2743 366 2747 370
rect 2847 366 2851 370
rect 2967 366 2971 370
rect 3095 366 3099 370
rect 3239 366 3243 370
rect 3383 366 3387 370
rect 3511 366 3515 370
rect 143 326 147 330
rect 279 326 283 330
rect 455 326 459 330
rect 639 326 643 330
rect 823 326 827 330
rect 999 326 1003 330
rect 1167 326 1171 330
rect 1327 326 1331 330
rect 1479 326 1483 330
rect 1623 326 1627 330
rect 1751 326 1755 330
rect 2031 322 2035 326
rect 2119 322 2123 326
rect 2223 322 2227 326
rect 2335 322 2339 326
rect 2447 322 2451 326
rect 2567 322 2571 326
rect 2695 322 2699 326
rect 2839 322 2843 326
rect 2999 322 3003 326
rect 3167 322 3171 326
rect 3343 322 3347 326
rect 3511 322 3515 326
rect 111 308 115 312
rect 1831 308 1835 312
rect 1871 304 1875 308
rect 3591 304 3595 308
rect 111 291 115 295
rect 135 288 139 292
rect 271 288 275 292
rect 447 288 451 292
rect 631 288 635 292
rect 815 288 819 292
rect 991 288 995 292
rect 1159 288 1163 292
rect 1319 288 1323 292
rect 1471 288 1475 292
rect 1615 288 1619 292
rect 1743 288 1747 292
rect 1831 291 1835 295
rect 1871 287 1875 291
rect 2023 284 2027 288
rect 2111 284 2115 288
rect 2215 284 2219 288
rect 2327 284 2331 288
rect 2439 284 2443 288
rect 2559 284 2563 288
rect 2687 284 2691 288
rect 2831 284 2835 288
rect 2991 284 2995 288
rect 3159 284 3163 288
rect 3335 284 3339 288
rect 3503 284 3507 288
rect 3591 287 3595 291
rect 111 237 115 241
rect 303 240 307 244
rect 391 240 395 244
rect 495 240 499 244
rect 599 240 603 244
rect 711 240 715 244
rect 823 240 827 244
rect 943 240 947 244
rect 1063 240 1067 244
rect 1175 240 1179 244
rect 1287 240 1291 244
rect 1407 240 1411 244
rect 1527 240 1531 244
rect 1647 240 1651 244
rect 1743 240 1747 244
rect 1831 237 1835 241
rect 1871 233 1875 237
rect 2071 236 2075 240
rect 2319 236 2323 240
rect 2543 236 2547 240
rect 2743 236 2747 240
rect 2927 236 2931 240
rect 3087 236 3091 240
rect 3239 236 3243 240
rect 3383 236 3387 240
rect 3503 236 3507 240
rect 3591 233 3595 237
rect 111 220 115 224
rect 1831 220 1835 224
rect 1871 216 1875 220
rect 3591 216 3595 220
rect 311 202 315 206
rect 399 202 403 206
rect 503 202 507 206
rect 607 202 611 206
rect 719 202 723 206
rect 831 202 835 206
rect 951 202 955 206
rect 1071 202 1075 206
rect 1183 202 1187 206
rect 1295 202 1299 206
rect 1415 202 1419 206
rect 1535 202 1539 206
rect 1655 202 1659 206
rect 1751 202 1755 206
rect 2079 198 2083 202
rect 2327 198 2331 202
rect 2551 198 2555 202
rect 2751 198 2755 202
rect 2935 198 2939 202
rect 3095 198 3099 202
rect 3247 198 3251 202
rect 3391 198 3395 202
rect 3511 198 3515 202
rect 263 146 267 150
rect 343 146 347 150
rect 423 146 427 150
rect 503 146 507 150
rect 583 146 587 150
rect 663 146 667 150
rect 743 146 747 150
rect 823 146 827 150
rect 903 146 907 150
rect 983 146 987 150
rect 1063 146 1067 150
rect 1143 146 1147 150
rect 1223 146 1227 150
rect 1303 146 1307 150
rect 1383 146 1387 150
rect 1463 146 1467 150
rect 1543 146 1547 150
rect 1903 142 1907 146
rect 1983 142 1987 146
rect 2063 142 2067 146
rect 2143 142 2147 146
rect 2223 142 2227 146
rect 2303 142 2307 146
rect 2399 142 2403 146
rect 2503 142 2507 146
rect 2607 142 2611 146
rect 2711 142 2715 146
rect 2815 142 2819 146
rect 2911 142 2915 146
rect 2999 142 3003 146
rect 3087 142 3091 146
rect 3175 142 3179 146
rect 3263 142 3267 146
rect 3351 142 3355 146
rect 3431 142 3435 146
rect 3511 142 3515 146
rect 111 128 115 132
rect 1831 128 1835 132
rect 1871 124 1875 128
rect 3591 124 3595 128
rect 111 111 115 115
rect 255 108 259 112
rect 335 108 339 112
rect 415 108 419 112
rect 495 108 499 112
rect 575 108 579 112
rect 655 108 659 112
rect 735 108 739 112
rect 815 108 819 112
rect 895 108 899 112
rect 975 108 979 112
rect 1055 108 1059 112
rect 1135 108 1139 112
rect 1215 108 1219 112
rect 1295 108 1299 112
rect 1375 108 1379 112
rect 1455 108 1459 112
rect 1535 108 1539 112
rect 1831 111 1835 115
rect 1871 107 1875 111
rect 1895 104 1899 108
rect 1975 104 1979 108
rect 2055 104 2059 108
rect 2135 104 2139 108
rect 2215 104 2219 108
rect 2295 104 2299 108
rect 2391 104 2395 108
rect 2495 104 2499 108
rect 2599 104 2603 108
rect 2703 104 2707 108
rect 2807 104 2811 108
rect 2903 104 2907 108
rect 2991 104 2995 108
rect 3079 104 3083 108
rect 3167 104 3171 108
rect 3255 104 3259 108
rect 3343 104 3347 108
rect 3423 104 3427 108
rect 3503 104 3507 108
rect 3591 107 3595 111
<< m3 >>
rect 111 3658 115 3659
rect 111 3653 115 3654
rect 143 3658 147 3659
rect 143 3653 147 3654
rect 223 3658 227 3659
rect 223 3653 227 3654
rect 351 3658 355 3659
rect 351 3653 355 3654
rect 495 3658 499 3659
rect 495 3653 499 3654
rect 647 3658 651 3659
rect 647 3653 651 3654
rect 807 3658 811 3659
rect 807 3653 811 3654
rect 975 3658 979 3659
rect 975 3653 979 3654
rect 1151 3658 1155 3659
rect 1151 3653 1155 3654
rect 1335 3658 1339 3659
rect 1335 3653 1339 3654
rect 1831 3658 1835 3659
rect 1831 3653 1835 3654
rect 112 3625 114 3653
rect 144 3643 146 3653
rect 224 3643 226 3653
rect 352 3643 354 3653
rect 496 3643 498 3653
rect 648 3643 650 3653
rect 808 3643 810 3653
rect 976 3643 978 3653
rect 1152 3643 1154 3653
rect 1336 3643 1338 3653
rect 142 3642 148 3643
rect 142 3638 143 3642
rect 147 3638 148 3642
rect 142 3637 148 3638
rect 222 3642 228 3643
rect 222 3638 223 3642
rect 227 3638 228 3642
rect 222 3637 228 3638
rect 350 3642 356 3643
rect 350 3638 351 3642
rect 355 3638 356 3642
rect 350 3637 356 3638
rect 494 3642 500 3643
rect 494 3638 495 3642
rect 499 3638 500 3642
rect 494 3637 500 3638
rect 646 3642 652 3643
rect 646 3638 647 3642
rect 651 3638 652 3642
rect 646 3637 652 3638
rect 806 3642 812 3643
rect 806 3638 807 3642
rect 811 3638 812 3642
rect 806 3637 812 3638
rect 974 3642 980 3643
rect 974 3638 975 3642
rect 979 3638 980 3642
rect 974 3637 980 3638
rect 1150 3642 1156 3643
rect 1150 3638 1151 3642
rect 1155 3638 1156 3642
rect 1150 3637 1156 3638
rect 1334 3642 1340 3643
rect 1334 3638 1335 3642
rect 1339 3638 1340 3642
rect 1334 3637 1340 3638
rect 1832 3625 1834 3653
rect 1871 3630 1875 3631
rect 1871 3625 1875 3626
rect 1927 3630 1931 3631
rect 1927 3625 1931 3626
rect 2007 3630 2011 3631
rect 2007 3625 2011 3626
rect 2103 3630 2107 3631
rect 2103 3625 2107 3626
rect 2207 3630 2211 3631
rect 2207 3625 2211 3626
rect 2319 3630 2323 3631
rect 2319 3625 2323 3626
rect 2431 3630 2435 3631
rect 2431 3625 2435 3626
rect 2551 3630 2555 3631
rect 2551 3625 2555 3626
rect 2663 3630 2667 3631
rect 2663 3625 2667 3626
rect 2775 3630 2779 3631
rect 2775 3625 2779 3626
rect 2879 3630 2883 3631
rect 2879 3625 2883 3626
rect 2983 3630 2987 3631
rect 2983 3625 2987 3626
rect 3095 3630 3099 3631
rect 3095 3625 3099 3626
rect 3207 3630 3211 3631
rect 3207 3625 3211 3626
rect 3591 3630 3595 3631
rect 3591 3625 3595 3626
rect 110 3624 116 3625
rect 110 3620 111 3624
rect 115 3620 116 3624
rect 110 3619 116 3620
rect 1830 3624 1836 3625
rect 1830 3620 1831 3624
rect 1835 3620 1836 3624
rect 1830 3619 1836 3620
rect 110 3607 116 3608
rect 110 3603 111 3607
rect 115 3603 116 3607
rect 1830 3607 1836 3608
rect 110 3602 116 3603
rect 134 3604 140 3605
rect 112 3583 114 3602
rect 134 3600 135 3604
rect 139 3600 140 3604
rect 134 3599 140 3600
rect 214 3604 220 3605
rect 214 3600 215 3604
rect 219 3600 220 3604
rect 214 3599 220 3600
rect 342 3604 348 3605
rect 342 3600 343 3604
rect 347 3600 348 3604
rect 342 3599 348 3600
rect 486 3604 492 3605
rect 486 3600 487 3604
rect 491 3600 492 3604
rect 486 3599 492 3600
rect 638 3604 644 3605
rect 638 3600 639 3604
rect 643 3600 644 3604
rect 638 3599 644 3600
rect 798 3604 804 3605
rect 798 3600 799 3604
rect 803 3600 804 3604
rect 798 3599 804 3600
rect 966 3604 972 3605
rect 966 3600 967 3604
rect 971 3600 972 3604
rect 966 3599 972 3600
rect 1142 3604 1148 3605
rect 1142 3600 1143 3604
rect 1147 3600 1148 3604
rect 1142 3599 1148 3600
rect 1326 3604 1332 3605
rect 1326 3600 1327 3604
rect 1331 3600 1332 3604
rect 1830 3603 1831 3607
rect 1835 3603 1836 3607
rect 1830 3602 1836 3603
rect 1326 3599 1332 3600
rect 136 3583 138 3599
rect 216 3583 218 3599
rect 344 3583 346 3599
rect 488 3583 490 3599
rect 640 3583 642 3599
rect 800 3583 802 3599
rect 968 3583 970 3599
rect 1144 3583 1146 3599
rect 1328 3583 1330 3599
rect 1832 3583 1834 3602
rect 1872 3597 1874 3625
rect 1928 3615 1930 3625
rect 2008 3615 2010 3625
rect 2104 3615 2106 3625
rect 2208 3615 2210 3625
rect 2320 3615 2322 3625
rect 2432 3615 2434 3625
rect 2552 3615 2554 3625
rect 2664 3615 2666 3625
rect 2776 3615 2778 3625
rect 2880 3615 2882 3625
rect 2984 3615 2986 3625
rect 3096 3615 3098 3625
rect 3208 3615 3210 3625
rect 1926 3614 1932 3615
rect 1926 3610 1927 3614
rect 1931 3610 1932 3614
rect 1926 3609 1932 3610
rect 2006 3614 2012 3615
rect 2006 3610 2007 3614
rect 2011 3610 2012 3614
rect 2006 3609 2012 3610
rect 2102 3614 2108 3615
rect 2102 3610 2103 3614
rect 2107 3610 2108 3614
rect 2102 3609 2108 3610
rect 2206 3614 2212 3615
rect 2206 3610 2207 3614
rect 2211 3610 2212 3614
rect 2206 3609 2212 3610
rect 2318 3614 2324 3615
rect 2318 3610 2319 3614
rect 2323 3610 2324 3614
rect 2318 3609 2324 3610
rect 2430 3614 2436 3615
rect 2430 3610 2431 3614
rect 2435 3610 2436 3614
rect 2430 3609 2436 3610
rect 2550 3614 2556 3615
rect 2550 3610 2551 3614
rect 2555 3610 2556 3614
rect 2550 3609 2556 3610
rect 2662 3614 2668 3615
rect 2662 3610 2663 3614
rect 2667 3610 2668 3614
rect 2662 3609 2668 3610
rect 2774 3614 2780 3615
rect 2774 3610 2775 3614
rect 2779 3610 2780 3614
rect 2774 3609 2780 3610
rect 2878 3614 2884 3615
rect 2878 3610 2879 3614
rect 2883 3610 2884 3614
rect 2878 3609 2884 3610
rect 2982 3614 2988 3615
rect 2982 3610 2983 3614
rect 2987 3610 2988 3614
rect 2982 3609 2988 3610
rect 3094 3614 3100 3615
rect 3094 3610 3095 3614
rect 3099 3610 3100 3614
rect 3094 3609 3100 3610
rect 3206 3614 3212 3615
rect 3206 3610 3207 3614
rect 3211 3610 3212 3614
rect 3206 3609 3212 3610
rect 3592 3597 3594 3625
rect 1870 3596 1876 3597
rect 1870 3592 1871 3596
rect 1875 3592 1876 3596
rect 1870 3591 1876 3592
rect 3590 3596 3596 3597
rect 3590 3592 3591 3596
rect 3595 3592 3596 3596
rect 3590 3591 3596 3592
rect 111 3582 115 3583
rect 111 3577 115 3578
rect 135 3582 139 3583
rect 135 3577 139 3578
rect 215 3582 219 3583
rect 215 3577 219 3578
rect 239 3582 243 3583
rect 239 3577 243 3578
rect 343 3582 347 3583
rect 343 3577 347 3578
rect 359 3582 363 3583
rect 359 3577 363 3578
rect 479 3582 483 3583
rect 479 3577 483 3578
rect 487 3582 491 3583
rect 487 3577 491 3578
rect 607 3582 611 3583
rect 607 3577 611 3578
rect 639 3582 643 3583
rect 639 3577 643 3578
rect 735 3582 739 3583
rect 735 3577 739 3578
rect 799 3582 803 3583
rect 799 3577 803 3578
rect 863 3582 867 3583
rect 863 3577 867 3578
rect 967 3582 971 3583
rect 967 3577 971 3578
rect 983 3582 987 3583
rect 983 3577 987 3578
rect 1095 3582 1099 3583
rect 1095 3577 1099 3578
rect 1143 3582 1147 3583
rect 1143 3577 1147 3578
rect 1207 3582 1211 3583
rect 1207 3577 1211 3578
rect 1319 3582 1323 3583
rect 1319 3577 1323 3578
rect 1327 3582 1331 3583
rect 1327 3577 1331 3578
rect 1439 3582 1443 3583
rect 1439 3577 1443 3578
rect 1831 3582 1835 3583
rect 1831 3577 1835 3578
rect 1870 3579 1876 3580
rect 112 3558 114 3577
rect 240 3561 242 3577
rect 360 3561 362 3577
rect 480 3561 482 3577
rect 608 3561 610 3577
rect 736 3561 738 3577
rect 864 3561 866 3577
rect 984 3561 986 3577
rect 1096 3561 1098 3577
rect 1208 3561 1210 3577
rect 1320 3561 1322 3577
rect 1440 3561 1442 3577
rect 238 3560 244 3561
rect 110 3557 116 3558
rect 110 3553 111 3557
rect 115 3553 116 3557
rect 238 3556 239 3560
rect 243 3556 244 3560
rect 238 3555 244 3556
rect 358 3560 364 3561
rect 358 3556 359 3560
rect 363 3556 364 3560
rect 358 3555 364 3556
rect 478 3560 484 3561
rect 478 3556 479 3560
rect 483 3556 484 3560
rect 478 3555 484 3556
rect 606 3560 612 3561
rect 606 3556 607 3560
rect 611 3556 612 3560
rect 606 3555 612 3556
rect 734 3560 740 3561
rect 734 3556 735 3560
rect 739 3556 740 3560
rect 734 3555 740 3556
rect 862 3560 868 3561
rect 862 3556 863 3560
rect 867 3556 868 3560
rect 862 3555 868 3556
rect 982 3560 988 3561
rect 982 3556 983 3560
rect 987 3556 988 3560
rect 982 3555 988 3556
rect 1094 3560 1100 3561
rect 1094 3556 1095 3560
rect 1099 3556 1100 3560
rect 1094 3555 1100 3556
rect 1206 3560 1212 3561
rect 1206 3556 1207 3560
rect 1211 3556 1212 3560
rect 1206 3555 1212 3556
rect 1318 3560 1324 3561
rect 1318 3556 1319 3560
rect 1323 3556 1324 3560
rect 1318 3555 1324 3556
rect 1438 3560 1444 3561
rect 1438 3556 1439 3560
rect 1443 3556 1444 3560
rect 1832 3558 1834 3577
rect 1870 3575 1871 3579
rect 1875 3575 1876 3579
rect 3590 3579 3596 3580
rect 1870 3574 1876 3575
rect 1918 3576 1924 3577
rect 1438 3555 1444 3556
rect 1830 3557 1836 3558
rect 110 3552 116 3553
rect 1830 3553 1831 3557
rect 1835 3553 1836 3557
rect 1872 3555 1874 3574
rect 1918 3572 1919 3576
rect 1923 3572 1924 3576
rect 1918 3571 1924 3572
rect 1998 3576 2004 3577
rect 1998 3572 1999 3576
rect 2003 3572 2004 3576
rect 1998 3571 2004 3572
rect 2094 3576 2100 3577
rect 2094 3572 2095 3576
rect 2099 3572 2100 3576
rect 2094 3571 2100 3572
rect 2198 3576 2204 3577
rect 2198 3572 2199 3576
rect 2203 3572 2204 3576
rect 2198 3571 2204 3572
rect 2310 3576 2316 3577
rect 2310 3572 2311 3576
rect 2315 3572 2316 3576
rect 2310 3571 2316 3572
rect 2422 3576 2428 3577
rect 2422 3572 2423 3576
rect 2427 3572 2428 3576
rect 2422 3571 2428 3572
rect 2542 3576 2548 3577
rect 2542 3572 2543 3576
rect 2547 3572 2548 3576
rect 2542 3571 2548 3572
rect 2654 3576 2660 3577
rect 2654 3572 2655 3576
rect 2659 3572 2660 3576
rect 2654 3571 2660 3572
rect 2766 3576 2772 3577
rect 2766 3572 2767 3576
rect 2771 3572 2772 3576
rect 2766 3571 2772 3572
rect 2870 3576 2876 3577
rect 2870 3572 2871 3576
rect 2875 3572 2876 3576
rect 2870 3571 2876 3572
rect 2974 3576 2980 3577
rect 2974 3572 2975 3576
rect 2979 3572 2980 3576
rect 2974 3571 2980 3572
rect 3086 3576 3092 3577
rect 3086 3572 3087 3576
rect 3091 3572 3092 3576
rect 3086 3571 3092 3572
rect 3198 3576 3204 3577
rect 3198 3572 3199 3576
rect 3203 3572 3204 3576
rect 3590 3575 3591 3579
rect 3595 3575 3596 3579
rect 3590 3574 3596 3575
rect 3198 3571 3204 3572
rect 1920 3555 1922 3571
rect 2000 3555 2002 3571
rect 2096 3555 2098 3571
rect 2200 3555 2202 3571
rect 2312 3555 2314 3571
rect 2424 3555 2426 3571
rect 2544 3555 2546 3571
rect 2656 3555 2658 3571
rect 2768 3555 2770 3571
rect 2872 3555 2874 3571
rect 2976 3555 2978 3571
rect 3088 3555 3090 3571
rect 3200 3555 3202 3571
rect 3592 3555 3594 3574
rect 1830 3552 1836 3553
rect 1871 3554 1875 3555
rect 1871 3549 1875 3550
rect 1919 3554 1923 3555
rect 1919 3549 1923 3550
rect 1943 3554 1947 3555
rect 1943 3549 1947 3550
rect 1999 3554 2003 3555
rect 1999 3549 2003 3550
rect 2095 3554 2099 3555
rect 2095 3549 2099 3550
rect 2127 3554 2131 3555
rect 2127 3549 2131 3550
rect 2199 3554 2203 3555
rect 2199 3549 2203 3550
rect 2303 3554 2307 3555
rect 2303 3549 2307 3550
rect 2311 3554 2315 3555
rect 2311 3549 2315 3550
rect 2423 3554 2427 3555
rect 2423 3549 2427 3550
rect 2479 3554 2483 3555
rect 2479 3549 2483 3550
rect 2543 3554 2547 3555
rect 2543 3549 2547 3550
rect 2647 3554 2651 3555
rect 2647 3549 2651 3550
rect 2655 3554 2659 3555
rect 2655 3549 2659 3550
rect 2767 3554 2771 3555
rect 2767 3549 2771 3550
rect 2815 3554 2819 3555
rect 2815 3549 2819 3550
rect 2871 3554 2875 3555
rect 2871 3549 2875 3550
rect 2975 3554 2979 3555
rect 2975 3549 2979 3550
rect 3087 3554 3091 3555
rect 3087 3549 3091 3550
rect 3135 3554 3139 3555
rect 3135 3549 3139 3550
rect 3199 3554 3203 3555
rect 3199 3549 3203 3550
rect 3303 3554 3307 3555
rect 3303 3549 3307 3550
rect 3591 3554 3595 3555
rect 3591 3549 3595 3550
rect 110 3540 116 3541
rect 110 3536 111 3540
rect 115 3536 116 3540
rect 110 3535 116 3536
rect 1830 3540 1836 3541
rect 1830 3536 1831 3540
rect 1835 3536 1836 3540
rect 1830 3535 1836 3536
rect 112 3507 114 3535
rect 246 3522 252 3523
rect 246 3518 247 3522
rect 251 3518 252 3522
rect 246 3517 252 3518
rect 366 3522 372 3523
rect 366 3518 367 3522
rect 371 3518 372 3522
rect 366 3517 372 3518
rect 486 3522 492 3523
rect 486 3518 487 3522
rect 491 3518 492 3522
rect 486 3517 492 3518
rect 614 3522 620 3523
rect 614 3518 615 3522
rect 619 3518 620 3522
rect 614 3517 620 3518
rect 742 3522 748 3523
rect 742 3518 743 3522
rect 747 3518 748 3522
rect 742 3517 748 3518
rect 870 3522 876 3523
rect 870 3518 871 3522
rect 875 3518 876 3522
rect 870 3517 876 3518
rect 990 3522 996 3523
rect 990 3518 991 3522
rect 995 3518 996 3522
rect 990 3517 996 3518
rect 1102 3522 1108 3523
rect 1102 3518 1103 3522
rect 1107 3518 1108 3522
rect 1102 3517 1108 3518
rect 1214 3522 1220 3523
rect 1214 3518 1215 3522
rect 1219 3518 1220 3522
rect 1214 3517 1220 3518
rect 1326 3522 1332 3523
rect 1326 3518 1327 3522
rect 1331 3518 1332 3522
rect 1326 3517 1332 3518
rect 1446 3522 1452 3523
rect 1446 3518 1447 3522
rect 1451 3518 1452 3522
rect 1446 3517 1452 3518
rect 248 3507 250 3517
rect 368 3507 370 3517
rect 488 3507 490 3517
rect 616 3507 618 3517
rect 744 3507 746 3517
rect 872 3507 874 3517
rect 992 3507 994 3517
rect 1104 3507 1106 3517
rect 1216 3507 1218 3517
rect 1328 3507 1330 3517
rect 1448 3507 1450 3517
rect 1832 3507 1834 3535
rect 1872 3530 1874 3549
rect 1944 3533 1946 3549
rect 2128 3533 2130 3549
rect 2304 3533 2306 3549
rect 2480 3533 2482 3549
rect 2648 3533 2650 3549
rect 2816 3533 2818 3549
rect 2976 3533 2978 3549
rect 3136 3533 3138 3549
rect 3304 3533 3306 3549
rect 1942 3532 1948 3533
rect 1870 3529 1876 3530
rect 1870 3525 1871 3529
rect 1875 3525 1876 3529
rect 1942 3528 1943 3532
rect 1947 3528 1948 3532
rect 1942 3527 1948 3528
rect 2126 3532 2132 3533
rect 2126 3528 2127 3532
rect 2131 3528 2132 3532
rect 2126 3527 2132 3528
rect 2302 3532 2308 3533
rect 2302 3528 2303 3532
rect 2307 3528 2308 3532
rect 2302 3527 2308 3528
rect 2478 3532 2484 3533
rect 2478 3528 2479 3532
rect 2483 3528 2484 3532
rect 2478 3527 2484 3528
rect 2646 3532 2652 3533
rect 2646 3528 2647 3532
rect 2651 3528 2652 3532
rect 2646 3527 2652 3528
rect 2814 3532 2820 3533
rect 2814 3528 2815 3532
rect 2819 3528 2820 3532
rect 2814 3527 2820 3528
rect 2974 3532 2980 3533
rect 2974 3528 2975 3532
rect 2979 3528 2980 3532
rect 2974 3527 2980 3528
rect 3134 3532 3140 3533
rect 3134 3528 3135 3532
rect 3139 3528 3140 3532
rect 3134 3527 3140 3528
rect 3302 3532 3308 3533
rect 3302 3528 3303 3532
rect 3307 3528 3308 3532
rect 3592 3530 3594 3549
rect 3302 3527 3308 3528
rect 3590 3529 3596 3530
rect 1870 3524 1876 3525
rect 3590 3525 3591 3529
rect 3595 3525 3596 3529
rect 3590 3524 3596 3525
rect 1870 3512 1876 3513
rect 1870 3508 1871 3512
rect 1875 3508 1876 3512
rect 1870 3507 1876 3508
rect 3590 3512 3596 3513
rect 3590 3508 3591 3512
rect 3595 3508 3596 3512
rect 3590 3507 3596 3508
rect 111 3506 115 3507
rect 111 3501 115 3502
rect 167 3506 171 3507
rect 167 3501 171 3502
rect 247 3506 251 3507
rect 247 3501 251 3502
rect 287 3506 291 3507
rect 287 3501 291 3502
rect 367 3506 371 3507
rect 367 3501 371 3502
rect 415 3506 419 3507
rect 415 3501 419 3502
rect 487 3506 491 3507
rect 487 3501 491 3502
rect 551 3506 555 3507
rect 551 3501 555 3502
rect 615 3506 619 3507
rect 615 3501 619 3502
rect 687 3506 691 3507
rect 687 3501 691 3502
rect 743 3506 747 3507
rect 743 3501 747 3502
rect 823 3506 827 3507
rect 823 3501 827 3502
rect 871 3506 875 3507
rect 871 3501 875 3502
rect 951 3506 955 3507
rect 951 3501 955 3502
rect 991 3506 995 3507
rect 991 3501 995 3502
rect 1071 3506 1075 3507
rect 1071 3501 1075 3502
rect 1103 3506 1107 3507
rect 1103 3501 1107 3502
rect 1183 3506 1187 3507
rect 1183 3501 1187 3502
rect 1215 3506 1219 3507
rect 1215 3501 1219 3502
rect 1303 3506 1307 3507
rect 1303 3501 1307 3502
rect 1327 3506 1331 3507
rect 1327 3501 1331 3502
rect 1423 3506 1427 3507
rect 1423 3501 1427 3502
rect 1447 3506 1451 3507
rect 1447 3501 1451 3502
rect 1831 3506 1835 3507
rect 1831 3501 1835 3502
rect 112 3473 114 3501
rect 168 3491 170 3501
rect 288 3491 290 3501
rect 416 3491 418 3501
rect 552 3491 554 3501
rect 688 3491 690 3501
rect 824 3491 826 3501
rect 952 3491 954 3501
rect 1072 3491 1074 3501
rect 1184 3491 1186 3501
rect 1304 3491 1306 3501
rect 1424 3491 1426 3501
rect 166 3490 172 3491
rect 166 3486 167 3490
rect 171 3486 172 3490
rect 166 3485 172 3486
rect 286 3490 292 3491
rect 286 3486 287 3490
rect 291 3486 292 3490
rect 286 3485 292 3486
rect 414 3490 420 3491
rect 414 3486 415 3490
rect 419 3486 420 3490
rect 414 3485 420 3486
rect 550 3490 556 3491
rect 550 3486 551 3490
rect 555 3486 556 3490
rect 550 3485 556 3486
rect 686 3490 692 3491
rect 686 3486 687 3490
rect 691 3486 692 3490
rect 686 3485 692 3486
rect 822 3490 828 3491
rect 822 3486 823 3490
rect 827 3486 828 3490
rect 822 3485 828 3486
rect 950 3490 956 3491
rect 950 3486 951 3490
rect 955 3486 956 3490
rect 950 3485 956 3486
rect 1070 3490 1076 3491
rect 1070 3486 1071 3490
rect 1075 3486 1076 3490
rect 1070 3485 1076 3486
rect 1182 3490 1188 3491
rect 1182 3486 1183 3490
rect 1187 3486 1188 3490
rect 1182 3485 1188 3486
rect 1302 3490 1308 3491
rect 1302 3486 1303 3490
rect 1307 3486 1308 3490
rect 1302 3485 1308 3486
rect 1422 3490 1428 3491
rect 1422 3486 1423 3490
rect 1427 3486 1428 3490
rect 1422 3485 1428 3486
rect 1832 3473 1834 3501
rect 1872 3479 1874 3507
rect 1950 3494 1956 3495
rect 1950 3490 1951 3494
rect 1955 3490 1956 3494
rect 1950 3489 1956 3490
rect 2134 3494 2140 3495
rect 2134 3490 2135 3494
rect 2139 3490 2140 3494
rect 2134 3489 2140 3490
rect 2310 3494 2316 3495
rect 2310 3490 2311 3494
rect 2315 3490 2316 3494
rect 2310 3489 2316 3490
rect 2486 3494 2492 3495
rect 2486 3490 2487 3494
rect 2491 3490 2492 3494
rect 2486 3489 2492 3490
rect 2654 3494 2660 3495
rect 2654 3490 2655 3494
rect 2659 3490 2660 3494
rect 2654 3489 2660 3490
rect 2822 3494 2828 3495
rect 2822 3490 2823 3494
rect 2827 3490 2828 3494
rect 2822 3489 2828 3490
rect 2982 3494 2988 3495
rect 2982 3490 2983 3494
rect 2987 3490 2988 3494
rect 2982 3489 2988 3490
rect 3142 3494 3148 3495
rect 3142 3490 3143 3494
rect 3147 3490 3148 3494
rect 3142 3489 3148 3490
rect 3310 3494 3316 3495
rect 3310 3490 3311 3494
rect 3315 3490 3316 3494
rect 3310 3489 3316 3490
rect 1952 3479 1954 3489
rect 2136 3479 2138 3489
rect 2312 3479 2314 3489
rect 2488 3479 2490 3489
rect 2656 3479 2658 3489
rect 2824 3479 2826 3489
rect 2984 3479 2986 3489
rect 3144 3479 3146 3489
rect 3312 3479 3314 3489
rect 3592 3479 3594 3507
rect 1871 3478 1875 3479
rect 1871 3473 1875 3474
rect 1951 3478 1955 3479
rect 1951 3473 1955 3474
rect 1959 3478 1963 3479
rect 1959 3473 1963 3474
rect 2079 3478 2083 3479
rect 2079 3473 2083 3474
rect 2135 3478 2139 3479
rect 2135 3473 2139 3474
rect 2199 3478 2203 3479
rect 2199 3473 2203 3474
rect 2311 3478 2315 3479
rect 2311 3473 2315 3474
rect 2335 3478 2339 3479
rect 2335 3473 2339 3474
rect 2479 3478 2483 3479
rect 2479 3473 2483 3474
rect 2487 3478 2491 3479
rect 2487 3473 2491 3474
rect 2631 3478 2635 3479
rect 2631 3473 2635 3474
rect 2655 3478 2659 3479
rect 2655 3473 2659 3474
rect 2791 3478 2795 3479
rect 2791 3473 2795 3474
rect 2823 3478 2827 3479
rect 2823 3473 2827 3474
rect 2959 3478 2963 3479
rect 2959 3473 2963 3474
rect 2983 3478 2987 3479
rect 2983 3473 2987 3474
rect 3127 3478 3131 3479
rect 3127 3473 3131 3474
rect 3143 3478 3147 3479
rect 3143 3473 3147 3474
rect 3303 3478 3307 3479
rect 3303 3473 3307 3474
rect 3311 3478 3315 3479
rect 3311 3473 3315 3474
rect 3591 3478 3595 3479
rect 3591 3473 3595 3474
rect 110 3472 116 3473
rect 110 3468 111 3472
rect 115 3468 116 3472
rect 110 3467 116 3468
rect 1830 3472 1836 3473
rect 1830 3468 1831 3472
rect 1835 3468 1836 3472
rect 1830 3467 1836 3468
rect 110 3455 116 3456
rect 110 3451 111 3455
rect 115 3451 116 3455
rect 1830 3455 1836 3456
rect 110 3450 116 3451
rect 158 3452 164 3453
rect 112 3423 114 3450
rect 158 3448 159 3452
rect 163 3448 164 3452
rect 158 3447 164 3448
rect 278 3452 284 3453
rect 278 3448 279 3452
rect 283 3448 284 3452
rect 278 3447 284 3448
rect 406 3452 412 3453
rect 406 3448 407 3452
rect 411 3448 412 3452
rect 406 3447 412 3448
rect 542 3452 548 3453
rect 542 3448 543 3452
rect 547 3448 548 3452
rect 542 3447 548 3448
rect 678 3452 684 3453
rect 678 3448 679 3452
rect 683 3448 684 3452
rect 678 3447 684 3448
rect 814 3452 820 3453
rect 814 3448 815 3452
rect 819 3448 820 3452
rect 814 3447 820 3448
rect 942 3452 948 3453
rect 942 3448 943 3452
rect 947 3448 948 3452
rect 942 3447 948 3448
rect 1062 3452 1068 3453
rect 1062 3448 1063 3452
rect 1067 3448 1068 3452
rect 1062 3447 1068 3448
rect 1174 3452 1180 3453
rect 1174 3448 1175 3452
rect 1179 3448 1180 3452
rect 1174 3447 1180 3448
rect 1294 3452 1300 3453
rect 1294 3448 1295 3452
rect 1299 3448 1300 3452
rect 1294 3447 1300 3448
rect 1414 3452 1420 3453
rect 1414 3448 1415 3452
rect 1419 3448 1420 3452
rect 1830 3451 1831 3455
rect 1835 3451 1836 3455
rect 1830 3450 1836 3451
rect 1414 3447 1420 3448
rect 160 3423 162 3447
rect 280 3423 282 3447
rect 408 3423 410 3447
rect 544 3423 546 3447
rect 680 3423 682 3447
rect 816 3423 818 3447
rect 944 3423 946 3447
rect 1064 3423 1066 3447
rect 1176 3423 1178 3447
rect 1296 3423 1298 3447
rect 1416 3423 1418 3447
rect 1832 3423 1834 3450
rect 1872 3445 1874 3473
rect 1960 3463 1962 3473
rect 2080 3463 2082 3473
rect 2200 3463 2202 3473
rect 2336 3463 2338 3473
rect 2480 3463 2482 3473
rect 2632 3463 2634 3473
rect 2792 3463 2794 3473
rect 2960 3463 2962 3473
rect 3128 3463 3130 3473
rect 3304 3463 3306 3473
rect 1958 3462 1964 3463
rect 1958 3458 1959 3462
rect 1963 3458 1964 3462
rect 1958 3457 1964 3458
rect 2078 3462 2084 3463
rect 2078 3458 2079 3462
rect 2083 3458 2084 3462
rect 2078 3457 2084 3458
rect 2198 3462 2204 3463
rect 2198 3458 2199 3462
rect 2203 3458 2204 3462
rect 2198 3457 2204 3458
rect 2334 3462 2340 3463
rect 2334 3458 2335 3462
rect 2339 3458 2340 3462
rect 2334 3457 2340 3458
rect 2478 3462 2484 3463
rect 2478 3458 2479 3462
rect 2483 3458 2484 3462
rect 2478 3457 2484 3458
rect 2630 3462 2636 3463
rect 2630 3458 2631 3462
rect 2635 3458 2636 3462
rect 2630 3457 2636 3458
rect 2790 3462 2796 3463
rect 2790 3458 2791 3462
rect 2795 3458 2796 3462
rect 2790 3457 2796 3458
rect 2958 3462 2964 3463
rect 2958 3458 2959 3462
rect 2963 3458 2964 3462
rect 2958 3457 2964 3458
rect 3126 3462 3132 3463
rect 3126 3458 3127 3462
rect 3131 3458 3132 3462
rect 3126 3457 3132 3458
rect 3302 3462 3308 3463
rect 3302 3458 3303 3462
rect 3307 3458 3308 3462
rect 3302 3457 3308 3458
rect 3592 3445 3594 3473
rect 1870 3444 1876 3445
rect 1870 3440 1871 3444
rect 1875 3440 1876 3444
rect 1870 3439 1876 3440
rect 3590 3444 3596 3445
rect 3590 3440 3591 3444
rect 3595 3440 3596 3444
rect 3590 3439 3596 3440
rect 1870 3427 1876 3428
rect 1870 3423 1871 3427
rect 1875 3423 1876 3427
rect 3590 3427 3596 3428
rect 111 3422 115 3423
rect 111 3417 115 3418
rect 135 3422 139 3423
rect 135 3417 139 3418
rect 159 3422 163 3423
rect 159 3417 163 3418
rect 247 3422 251 3423
rect 247 3417 251 3418
rect 279 3422 283 3423
rect 279 3417 283 3418
rect 375 3422 379 3423
rect 375 3417 379 3418
rect 407 3422 411 3423
rect 407 3417 411 3418
rect 503 3422 507 3423
rect 503 3417 507 3418
rect 543 3422 547 3423
rect 543 3417 547 3418
rect 639 3422 643 3423
rect 639 3417 643 3418
rect 679 3422 683 3423
rect 679 3417 683 3418
rect 775 3422 779 3423
rect 775 3417 779 3418
rect 815 3422 819 3423
rect 815 3417 819 3418
rect 903 3422 907 3423
rect 903 3417 907 3418
rect 943 3422 947 3423
rect 943 3417 947 3418
rect 1031 3422 1035 3423
rect 1031 3417 1035 3418
rect 1063 3422 1067 3423
rect 1063 3417 1067 3418
rect 1159 3422 1163 3423
rect 1159 3417 1163 3418
rect 1175 3422 1179 3423
rect 1175 3417 1179 3418
rect 1287 3422 1291 3423
rect 1287 3417 1291 3418
rect 1295 3422 1299 3423
rect 1295 3417 1299 3418
rect 1415 3422 1419 3423
rect 1415 3417 1419 3418
rect 1831 3422 1835 3423
rect 1870 3422 1876 3423
rect 1950 3424 1956 3425
rect 1831 3417 1835 3418
rect 112 3398 114 3417
rect 136 3401 138 3417
rect 248 3401 250 3417
rect 376 3401 378 3417
rect 504 3401 506 3417
rect 640 3401 642 3417
rect 776 3401 778 3417
rect 904 3401 906 3417
rect 1032 3401 1034 3417
rect 1160 3401 1162 3417
rect 1288 3401 1290 3417
rect 1416 3401 1418 3417
rect 134 3400 140 3401
rect 110 3397 116 3398
rect 110 3393 111 3397
rect 115 3393 116 3397
rect 134 3396 135 3400
rect 139 3396 140 3400
rect 134 3395 140 3396
rect 246 3400 252 3401
rect 246 3396 247 3400
rect 251 3396 252 3400
rect 246 3395 252 3396
rect 374 3400 380 3401
rect 374 3396 375 3400
rect 379 3396 380 3400
rect 374 3395 380 3396
rect 502 3400 508 3401
rect 502 3396 503 3400
rect 507 3396 508 3400
rect 502 3395 508 3396
rect 638 3400 644 3401
rect 638 3396 639 3400
rect 643 3396 644 3400
rect 638 3395 644 3396
rect 774 3400 780 3401
rect 774 3396 775 3400
rect 779 3396 780 3400
rect 774 3395 780 3396
rect 902 3400 908 3401
rect 902 3396 903 3400
rect 907 3396 908 3400
rect 902 3395 908 3396
rect 1030 3400 1036 3401
rect 1030 3396 1031 3400
rect 1035 3396 1036 3400
rect 1030 3395 1036 3396
rect 1158 3400 1164 3401
rect 1158 3396 1159 3400
rect 1163 3396 1164 3400
rect 1158 3395 1164 3396
rect 1286 3400 1292 3401
rect 1286 3396 1287 3400
rect 1291 3396 1292 3400
rect 1286 3395 1292 3396
rect 1414 3400 1420 3401
rect 1414 3396 1415 3400
rect 1419 3396 1420 3400
rect 1832 3398 1834 3417
rect 1414 3395 1420 3396
rect 1830 3397 1836 3398
rect 110 3392 116 3393
rect 1830 3393 1831 3397
rect 1835 3393 1836 3397
rect 1872 3395 1874 3422
rect 1950 3420 1951 3424
rect 1955 3420 1956 3424
rect 1950 3419 1956 3420
rect 2070 3424 2076 3425
rect 2070 3420 2071 3424
rect 2075 3420 2076 3424
rect 2070 3419 2076 3420
rect 2190 3424 2196 3425
rect 2190 3420 2191 3424
rect 2195 3420 2196 3424
rect 2190 3419 2196 3420
rect 2326 3424 2332 3425
rect 2326 3420 2327 3424
rect 2331 3420 2332 3424
rect 2326 3419 2332 3420
rect 2470 3424 2476 3425
rect 2470 3420 2471 3424
rect 2475 3420 2476 3424
rect 2470 3419 2476 3420
rect 2622 3424 2628 3425
rect 2622 3420 2623 3424
rect 2627 3420 2628 3424
rect 2622 3419 2628 3420
rect 2782 3424 2788 3425
rect 2782 3420 2783 3424
rect 2787 3420 2788 3424
rect 2782 3419 2788 3420
rect 2950 3424 2956 3425
rect 2950 3420 2951 3424
rect 2955 3420 2956 3424
rect 2950 3419 2956 3420
rect 3118 3424 3124 3425
rect 3118 3420 3119 3424
rect 3123 3420 3124 3424
rect 3118 3419 3124 3420
rect 3294 3424 3300 3425
rect 3294 3420 3295 3424
rect 3299 3420 3300 3424
rect 3590 3423 3591 3427
rect 3595 3423 3596 3427
rect 3590 3422 3596 3423
rect 3294 3419 3300 3420
rect 1952 3395 1954 3419
rect 2072 3395 2074 3419
rect 2192 3395 2194 3419
rect 2328 3395 2330 3419
rect 2472 3395 2474 3419
rect 2624 3395 2626 3419
rect 2784 3395 2786 3419
rect 2952 3395 2954 3419
rect 3120 3395 3122 3419
rect 3296 3395 3298 3419
rect 3592 3395 3594 3422
rect 1830 3392 1836 3393
rect 1871 3394 1875 3395
rect 1871 3389 1875 3390
rect 1951 3394 1955 3395
rect 1951 3389 1955 3390
rect 1975 3394 1979 3395
rect 1975 3389 1979 3390
rect 2071 3394 2075 3395
rect 2071 3389 2075 3390
rect 2135 3394 2139 3395
rect 2135 3389 2139 3390
rect 2191 3394 2195 3395
rect 2191 3389 2195 3390
rect 2287 3394 2291 3395
rect 2287 3389 2291 3390
rect 2327 3394 2331 3395
rect 2327 3389 2331 3390
rect 2431 3394 2435 3395
rect 2431 3389 2435 3390
rect 2471 3394 2475 3395
rect 2471 3389 2475 3390
rect 2559 3394 2563 3395
rect 2559 3389 2563 3390
rect 2623 3394 2627 3395
rect 2623 3389 2627 3390
rect 2679 3394 2683 3395
rect 2679 3389 2683 3390
rect 2783 3394 2787 3395
rect 2783 3389 2787 3390
rect 2791 3394 2795 3395
rect 2791 3389 2795 3390
rect 2895 3394 2899 3395
rect 2895 3389 2899 3390
rect 2951 3394 2955 3395
rect 2951 3389 2955 3390
rect 2991 3394 2995 3395
rect 2991 3389 2995 3390
rect 3079 3394 3083 3395
rect 3079 3389 3083 3390
rect 3119 3394 3123 3395
rect 3119 3389 3123 3390
rect 3167 3394 3171 3395
rect 3167 3389 3171 3390
rect 3255 3394 3259 3395
rect 3255 3389 3259 3390
rect 3295 3394 3299 3395
rect 3295 3389 3299 3390
rect 3343 3394 3347 3395
rect 3343 3389 3347 3390
rect 3423 3394 3427 3395
rect 3423 3389 3427 3390
rect 3503 3394 3507 3395
rect 3503 3389 3507 3390
rect 3591 3394 3595 3395
rect 3591 3389 3595 3390
rect 110 3380 116 3381
rect 110 3376 111 3380
rect 115 3376 116 3380
rect 110 3375 116 3376
rect 1830 3380 1836 3381
rect 1830 3376 1831 3380
rect 1835 3376 1836 3380
rect 1830 3375 1836 3376
rect 112 3343 114 3375
rect 142 3362 148 3363
rect 142 3358 143 3362
rect 147 3358 148 3362
rect 142 3357 148 3358
rect 254 3362 260 3363
rect 254 3358 255 3362
rect 259 3358 260 3362
rect 254 3357 260 3358
rect 382 3362 388 3363
rect 382 3358 383 3362
rect 387 3358 388 3362
rect 382 3357 388 3358
rect 510 3362 516 3363
rect 510 3358 511 3362
rect 515 3358 516 3362
rect 510 3357 516 3358
rect 646 3362 652 3363
rect 646 3358 647 3362
rect 651 3358 652 3362
rect 646 3357 652 3358
rect 782 3362 788 3363
rect 782 3358 783 3362
rect 787 3358 788 3362
rect 782 3357 788 3358
rect 910 3362 916 3363
rect 910 3358 911 3362
rect 915 3358 916 3362
rect 910 3357 916 3358
rect 1038 3362 1044 3363
rect 1038 3358 1039 3362
rect 1043 3358 1044 3362
rect 1038 3357 1044 3358
rect 1166 3362 1172 3363
rect 1166 3358 1167 3362
rect 1171 3358 1172 3362
rect 1166 3357 1172 3358
rect 1294 3362 1300 3363
rect 1294 3358 1295 3362
rect 1299 3358 1300 3362
rect 1294 3357 1300 3358
rect 1422 3362 1428 3363
rect 1422 3358 1423 3362
rect 1427 3358 1428 3362
rect 1422 3357 1428 3358
rect 144 3343 146 3357
rect 256 3343 258 3357
rect 384 3343 386 3357
rect 512 3343 514 3357
rect 648 3343 650 3357
rect 784 3343 786 3357
rect 912 3343 914 3357
rect 1040 3343 1042 3357
rect 1168 3343 1170 3357
rect 1296 3343 1298 3357
rect 1424 3343 1426 3357
rect 1832 3343 1834 3375
rect 1872 3370 1874 3389
rect 1976 3373 1978 3389
rect 2136 3373 2138 3389
rect 2288 3373 2290 3389
rect 2432 3373 2434 3389
rect 2560 3373 2562 3389
rect 2680 3373 2682 3389
rect 2792 3373 2794 3389
rect 2896 3373 2898 3389
rect 2992 3373 2994 3389
rect 3080 3373 3082 3389
rect 3168 3373 3170 3389
rect 3256 3373 3258 3389
rect 3344 3373 3346 3389
rect 3424 3373 3426 3389
rect 3504 3373 3506 3389
rect 1974 3372 1980 3373
rect 1870 3369 1876 3370
rect 1870 3365 1871 3369
rect 1875 3365 1876 3369
rect 1974 3368 1975 3372
rect 1979 3368 1980 3372
rect 1974 3367 1980 3368
rect 2134 3372 2140 3373
rect 2134 3368 2135 3372
rect 2139 3368 2140 3372
rect 2134 3367 2140 3368
rect 2286 3372 2292 3373
rect 2286 3368 2287 3372
rect 2291 3368 2292 3372
rect 2286 3367 2292 3368
rect 2430 3372 2436 3373
rect 2430 3368 2431 3372
rect 2435 3368 2436 3372
rect 2430 3367 2436 3368
rect 2558 3372 2564 3373
rect 2558 3368 2559 3372
rect 2563 3368 2564 3372
rect 2558 3367 2564 3368
rect 2678 3372 2684 3373
rect 2678 3368 2679 3372
rect 2683 3368 2684 3372
rect 2678 3367 2684 3368
rect 2790 3372 2796 3373
rect 2790 3368 2791 3372
rect 2795 3368 2796 3372
rect 2790 3367 2796 3368
rect 2894 3372 2900 3373
rect 2894 3368 2895 3372
rect 2899 3368 2900 3372
rect 2894 3367 2900 3368
rect 2990 3372 2996 3373
rect 2990 3368 2991 3372
rect 2995 3368 2996 3372
rect 2990 3367 2996 3368
rect 3078 3372 3084 3373
rect 3078 3368 3079 3372
rect 3083 3368 3084 3372
rect 3078 3367 3084 3368
rect 3166 3372 3172 3373
rect 3166 3368 3167 3372
rect 3171 3368 3172 3372
rect 3166 3367 3172 3368
rect 3254 3372 3260 3373
rect 3254 3368 3255 3372
rect 3259 3368 3260 3372
rect 3254 3367 3260 3368
rect 3342 3372 3348 3373
rect 3342 3368 3343 3372
rect 3347 3368 3348 3372
rect 3342 3367 3348 3368
rect 3422 3372 3428 3373
rect 3422 3368 3423 3372
rect 3427 3368 3428 3372
rect 3422 3367 3428 3368
rect 3502 3372 3508 3373
rect 3502 3368 3503 3372
rect 3507 3368 3508 3372
rect 3592 3370 3594 3389
rect 3502 3367 3508 3368
rect 3590 3369 3596 3370
rect 1870 3364 1876 3365
rect 3590 3365 3591 3369
rect 3595 3365 3596 3369
rect 3590 3364 3596 3365
rect 1870 3352 1876 3353
rect 1870 3348 1871 3352
rect 1875 3348 1876 3352
rect 1870 3347 1876 3348
rect 3590 3352 3596 3353
rect 3590 3348 3591 3352
rect 3595 3348 3596 3352
rect 3590 3347 3596 3348
rect 111 3342 115 3343
rect 111 3337 115 3338
rect 143 3342 147 3343
rect 143 3337 147 3338
rect 255 3342 259 3343
rect 255 3337 259 3338
rect 271 3342 275 3343
rect 271 3337 275 3338
rect 383 3342 387 3343
rect 383 3337 387 3338
rect 391 3342 395 3343
rect 391 3337 395 3338
rect 511 3342 515 3343
rect 511 3337 515 3338
rect 519 3342 523 3343
rect 519 3337 523 3338
rect 647 3342 651 3343
rect 647 3337 651 3338
rect 655 3342 659 3343
rect 655 3337 659 3338
rect 783 3342 787 3343
rect 783 3337 787 3338
rect 791 3342 795 3343
rect 791 3337 795 3338
rect 911 3342 915 3343
rect 911 3337 915 3338
rect 919 3342 923 3343
rect 919 3337 923 3338
rect 1039 3342 1043 3343
rect 1039 3337 1043 3338
rect 1055 3342 1059 3343
rect 1055 3337 1059 3338
rect 1167 3342 1171 3343
rect 1167 3337 1171 3338
rect 1191 3342 1195 3343
rect 1191 3337 1195 3338
rect 1295 3342 1299 3343
rect 1295 3337 1299 3338
rect 1327 3342 1331 3343
rect 1327 3337 1331 3338
rect 1423 3342 1427 3343
rect 1423 3337 1427 3338
rect 1463 3342 1467 3343
rect 1463 3337 1467 3338
rect 1831 3342 1835 3343
rect 1831 3337 1835 3338
rect 112 3309 114 3337
rect 272 3327 274 3337
rect 392 3327 394 3337
rect 520 3327 522 3337
rect 656 3327 658 3337
rect 792 3327 794 3337
rect 920 3327 922 3337
rect 1056 3327 1058 3337
rect 1192 3327 1194 3337
rect 1328 3327 1330 3337
rect 1464 3327 1466 3337
rect 270 3326 276 3327
rect 270 3322 271 3326
rect 275 3322 276 3326
rect 270 3321 276 3322
rect 390 3326 396 3327
rect 390 3322 391 3326
rect 395 3322 396 3326
rect 390 3321 396 3322
rect 518 3326 524 3327
rect 518 3322 519 3326
rect 523 3322 524 3326
rect 518 3321 524 3322
rect 654 3326 660 3327
rect 654 3322 655 3326
rect 659 3322 660 3326
rect 654 3321 660 3322
rect 790 3326 796 3327
rect 790 3322 791 3326
rect 795 3322 796 3326
rect 790 3321 796 3322
rect 918 3326 924 3327
rect 918 3322 919 3326
rect 923 3322 924 3326
rect 918 3321 924 3322
rect 1054 3326 1060 3327
rect 1054 3322 1055 3326
rect 1059 3322 1060 3326
rect 1054 3321 1060 3322
rect 1190 3326 1196 3327
rect 1190 3322 1191 3326
rect 1195 3322 1196 3326
rect 1190 3321 1196 3322
rect 1326 3326 1332 3327
rect 1326 3322 1327 3326
rect 1331 3322 1332 3326
rect 1326 3321 1332 3322
rect 1462 3326 1468 3327
rect 1462 3322 1463 3326
rect 1467 3322 1468 3326
rect 1462 3321 1468 3322
rect 1832 3309 1834 3337
rect 1872 3315 1874 3347
rect 1982 3334 1988 3335
rect 1982 3330 1983 3334
rect 1987 3330 1988 3334
rect 1982 3329 1988 3330
rect 2142 3334 2148 3335
rect 2142 3330 2143 3334
rect 2147 3330 2148 3334
rect 2142 3329 2148 3330
rect 2294 3334 2300 3335
rect 2294 3330 2295 3334
rect 2299 3330 2300 3334
rect 2294 3329 2300 3330
rect 2438 3334 2444 3335
rect 2438 3330 2439 3334
rect 2443 3330 2444 3334
rect 2438 3329 2444 3330
rect 2566 3334 2572 3335
rect 2566 3330 2567 3334
rect 2571 3330 2572 3334
rect 2566 3329 2572 3330
rect 2686 3334 2692 3335
rect 2686 3330 2687 3334
rect 2691 3330 2692 3334
rect 2686 3329 2692 3330
rect 2798 3334 2804 3335
rect 2798 3330 2799 3334
rect 2803 3330 2804 3334
rect 2798 3329 2804 3330
rect 2902 3334 2908 3335
rect 2902 3330 2903 3334
rect 2907 3330 2908 3334
rect 2902 3329 2908 3330
rect 2998 3334 3004 3335
rect 2998 3330 2999 3334
rect 3003 3330 3004 3334
rect 2998 3329 3004 3330
rect 3086 3334 3092 3335
rect 3086 3330 3087 3334
rect 3091 3330 3092 3334
rect 3086 3329 3092 3330
rect 3174 3334 3180 3335
rect 3174 3330 3175 3334
rect 3179 3330 3180 3334
rect 3174 3329 3180 3330
rect 3262 3334 3268 3335
rect 3262 3330 3263 3334
rect 3267 3330 3268 3334
rect 3262 3329 3268 3330
rect 3350 3334 3356 3335
rect 3350 3330 3351 3334
rect 3355 3330 3356 3334
rect 3350 3329 3356 3330
rect 3430 3334 3436 3335
rect 3430 3330 3431 3334
rect 3435 3330 3436 3334
rect 3430 3329 3436 3330
rect 3510 3334 3516 3335
rect 3510 3330 3511 3334
rect 3515 3330 3516 3334
rect 3510 3329 3516 3330
rect 1984 3315 1986 3329
rect 2144 3315 2146 3329
rect 2296 3315 2298 3329
rect 2440 3315 2442 3329
rect 2568 3315 2570 3329
rect 2688 3315 2690 3329
rect 2800 3315 2802 3329
rect 2904 3315 2906 3329
rect 3000 3315 3002 3329
rect 3088 3315 3090 3329
rect 3176 3315 3178 3329
rect 3264 3315 3266 3329
rect 3352 3315 3354 3329
rect 3432 3315 3434 3329
rect 3512 3315 3514 3329
rect 3592 3315 3594 3347
rect 1871 3314 1875 3315
rect 1871 3309 1875 3310
rect 1935 3314 1939 3315
rect 1935 3309 1939 3310
rect 1983 3314 1987 3315
rect 1983 3309 1987 3310
rect 2071 3314 2075 3315
rect 2071 3309 2075 3310
rect 2143 3314 2147 3315
rect 2143 3309 2147 3310
rect 2207 3314 2211 3315
rect 2207 3309 2211 3310
rect 2295 3314 2299 3315
rect 2295 3309 2299 3310
rect 2367 3314 2371 3315
rect 2367 3309 2371 3310
rect 2439 3314 2443 3315
rect 2439 3309 2443 3310
rect 2551 3314 2555 3315
rect 2551 3309 2555 3310
rect 2567 3314 2571 3315
rect 2567 3309 2571 3310
rect 2687 3314 2691 3315
rect 2687 3309 2691 3310
rect 2767 3314 2771 3315
rect 2767 3309 2771 3310
rect 2799 3314 2803 3315
rect 2799 3309 2803 3310
rect 2903 3314 2907 3315
rect 2903 3309 2907 3310
rect 2999 3314 3003 3315
rect 2999 3309 3003 3310
rect 3007 3314 3011 3315
rect 3007 3309 3011 3310
rect 3087 3314 3091 3315
rect 3087 3309 3091 3310
rect 3175 3314 3179 3315
rect 3175 3309 3179 3310
rect 3255 3314 3259 3315
rect 3255 3309 3259 3310
rect 3263 3314 3267 3315
rect 3263 3309 3267 3310
rect 3351 3314 3355 3315
rect 3351 3309 3355 3310
rect 3431 3314 3435 3315
rect 3431 3309 3435 3310
rect 3511 3314 3515 3315
rect 3511 3309 3515 3310
rect 3591 3314 3595 3315
rect 3591 3309 3595 3310
rect 110 3308 116 3309
rect 110 3304 111 3308
rect 115 3304 116 3308
rect 110 3303 116 3304
rect 1830 3308 1836 3309
rect 1830 3304 1831 3308
rect 1835 3304 1836 3308
rect 1830 3303 1836 3304
rect 110 3291 116 3292
rect 110 3287 111 3291
rect 115 3287 116 3291
rect 1830 3291 1836 3292
rect 110 3286 116 3287
rect 262 3288 268 3289
rect 112 3263 114 3286
rect 262 3284 263 3288
rect 267 3284 268 3288
rect 262 3283 268 3284
rect 382 3288 388 3289
rect 382 3284 383 3288
rect 387 3284 388 3288
rect 382 3283 388 3284
rect 510 3288 516 3289
rect 510 3284 511 3288
rect 515 3284 516 3288
rect 510 3283 516 3284
rect 646 3288 652 3289
rect 646 3284 647 3288
rect 651 3284 652 3288
rect 646 3283 652 3284
rect 782 3288 788 3289
rect 782 3284 783 3288
rect 787 3284 788 3288
rect 782 3283 788 3284
rect 910 3288 916 3289
rect 910 3284 911 3288
rect 915 3284 916 3288
rect 910 3283 916 3284
rect 1046 3288 1052 3289
rect 1046 3284 1047 3288
rect 1051 3284 1052 3288
rect 1046 3283 1052 3284
rect 1182 3288 1188 3289
rect 1182 3284 1183 3288
rect 1187 3284 1188 3288
rect 1182 3283 1188 3284
rect 1318 3288 1324 3289
rect 1318 3284 1319 3288
rect 1323 3284 1324 3288
rect 1318 3283 1324 3284
rect 1454 3288 1460 3289
rect 1454 3284 1455 3288
rect 1459 3284 1460 3288
rect 1830 3287 1831 3291
rect 1835 3287 1836 3291
rect 1830 3286 1836 3287
rect 1454 3283 1460 3284
rect 264 3263 266 3283
rect 384 3263 386 3283
rect 512 3263 514 3283
rect 648 3263 650 3283
rect 784 3263 786 3283
rect 912 3263 914 3283
rect 1048 3263 1050 3283
rect 1184 3263 1186 3283
rect 1320 3263 1322 3283
rect 1456 3263 1458 3283
rect 1832 3263 1834 3286
rect 1872 3281 1874 3309
rect 1936 3299 1938 3309
rect 2072 3299 2074 3309
rect 2208 3299 2210 3309
rect 2368 3299 2370 3309
rect 2552 3299 2554 3309
rect 2768 3299 2770 3309
rect 3008 3299 3010 3309
rect 3256 3299 3258 3309
rect 3512 3299 3514 3309
rect 1934 3298 1940 3299
rect 1934 3294 1935 3298
rect 1939 3294 1940 3298
rect 1934 3293 1940 3294
rect 2070 3298 2076 3299
rect 2070 3294 2071 3298
rect 2075 3294 2076 3298
rect 2070 3293 2076 3294
rect 2206 3298 2212 3299
rect 2206 3294 2207 3298
rect 2211 3294 2212 3298
rect 2206 3293 2212 3294
rect 2366 3298 2372 3299
rect 2366 3294 2367 3298
rect 2371 3294 2372 3298
rect 2366 3293 2372 3294
rect 2550 3298 2556 3299
rect 2550 3294 2551 3298
rect 2555 3294 2556 3298
rect 2550 3293 2556 3294
rect 2766 3298 2772 3299
rect 2766 3294 2767 3298
rect 2771 3294 2772 3298
rect 2766 3293 2772 3294
rect 3006 3298 3012 3299
rect 3006 3294 3007 3298
rect 3011 3294 3012 3298
rect 3006 3293 3012 3294
rect 3254 3298 3260 3299
rect 3254 3294 3255 3298
rect 3259 3294 3260 3298
rect 3254 3293 3260 3294
rect 3510 3298 3516 3299
rect 3510 3294 3511 3298
rect 3515 3294 3516 3298
rect 3510 3293 3516 3294
rect 3592 3281 3594 3309
rect 1870 3280 1876 3281
rect 1870 3276 1871 3280
rect 1875 3276 1876 3280
rect 1870 3275 1876 3276
rect 3590 3280 3596 3281
rect 3590 3276 3591 3280
rect 3595 3276 3596 3280
rect 3590 3275 3596 3276
rect 1870 3263 1876 3264
rect 111 3262 115 3263
rect 111 3257 115 3258
rect 263 3262 267 3263
rect 263 3257 267 3258
rect 383 3262 387 3263
rect 383 3257 387 3258
rect 471 3262 475 3263
rect 471 3257 475 3258
rect 511 3262 515 3263
rect 511 3257 515 3258
rect 575 3262 579 3263
rect 575 3257 579 3258
rect 647 3262 651 3263
rect 647 3257 651 3258
rect 687 3262 691 3263
rect 687 3257 691 3258
rect 783 3262 787 3263
rect 783 3257 787 3258
rect 807 3262 811 3263
rect 807 3257 811 3258
rect 911 3262 915 3263
rect 911 3257 915 3258
rect 935 3262 939 3263
rect 935 3257 939 3258
rect 1047 3262 1051 3263
rect 1047 3257 1051 3258
rect 1063 3262 1067 3263
rect 1063 3257 1067 3258
rect 1183 3262 1187 3263
rect 1183 3257 1187 3258
rect 1191 3262 1195 3263
rect 1191 3257 1195 3258
rect 1319 3262 1323 3263
rect 1319 3257 1323 3258
rect 1447 3262 1451 3263
rect 1447 3257 1451 3258
rect 1455 3262 1459 3263
rect 1455 3257 1459 3258
rect 1575 3262 1579 3263
rect 1575 3257 1579 3258
rect 1831 3262 1835 3263
rect 1870 3259 1871 3263
rect 1875 3259 1876 3263
rect 3590 3263 3596 3264
rect 1870 3258 1876 3259
rect 1926 3260 1932 3261
rect 1831 3257 1835 3258
rect 112 3238 114 3257
rect 384 3241 386 3257
rect 472 3241 474 3257
rect 576 3241 578 3257
rect 688 3241 690 3257
rect 808 3241 810 3257
rect 936 3241 938 3257
rect 1064 3241 1066 3257
rect 1192 3241 1194 3257
rect 1320 3241 1322 3257
rect 1448 3241 1450 3257
rect 1576 3241 1578 3257
rect 382 3240 388 3241
rect 110 3237 116 3238
rect 110 3233 111 3237
rect 115 3233 116 3237
rect 382 3236 383 3240
rect 387 3236 388 3240
rect 382 3235 388 3236
rect 470 3240 476 3241
rect 470 3236 471 3240
rect 475 3236 476 3240
rect 470 3235 476 3236
rect 574 3240 580 3241
rect 574 3236 575 3240
rect 579 3236 580 3240
rect 574 3235 580 3236
rect 686 3240 692 3241
rect 686 3236 687 3240
rect 691 3236 692 3240
rect 686 3235 692 3236
rect 806 3240 812 3241
rect 806 3236 807 3240
rect 811 3236 812 3240
rect 806 3235 812 3236
rect 934 3240 940 3241
rect 934 3236 935 3240
rect 939 3236 940 3240
rect 934 3235 940 3236
rect 1062 3240 1068 3241
rect 1062 3236 1063 3240
rect 1067 3236 1068 3240
rect 1062 3235 1068 3236
rect 1190 3240 1196 3241
rect 1190 3236 1191 3240
rect 1195 3236 1196 3240
rect 1190 3235 1196 3236
rect 1318 3240 1324 3241
rect 1318 3236 1319 3240
rect 1323 3236 1324 3240
rect 1318 3235 1324 3236
rect 1446 3240 1452 3241
rect 1446 3236 1447 3240
rect 1451 3236 1452 3240
rect 1446 3235 1452 3236
rect 1574 3240 1580 3241
rect 1574 3236 1575 3240
rect 1579 3236 1580 3240
rect 1832 3238 1834 3257
rect 1574 3235 1580 3236
rect 1830 3237 1836 3238
rect 110 3232 116 3233
rect 1830 3233 1831 3237
rect 1835 3233 1836 3237
rect 1872 3235 1874 3258
rect 1926 3256 1927 3260
rect 1931 3256 1932 3260
rect 1926 3255 1932 3256
rect 2062 3260 2068 3261
rect 2062 3256 2063 3260
rect 2067 3256 2068 3260
rect 2062 3255 2068 3256
rect 2198 3260 2204 3261
rect 2198 3256 2199 3260
rect 2203 3256 2204 3260
rect 2198 3255 2204 3256
rect 2358 3260 2364 3261
rect 2358 3256 2359 3260
rect 2363 3256 2364 3260
rect 2358 3255 2364 3256
rect 2542 3260 2548 3261
rect 2542 3256 2543 3260
rect 2547 3256 2548 3260
rect 2542 3255 2548 3256
rect 2758 3260 2764 3261
rect 2758 3256 2759 3260
rect 2763 3256 2764 3260
rect 2758 3255 2764 3256
rect 2998 3260 3004 3261
rect 2998 3256 2999 3260
rect 3003 3256 3004 3260
rect 2998 3255 3004 3256
rect 3246 3260 3252 3261
rect 3246 3256 3247 3260
rect 3251 3256 3252 3260
rect 3246 3255 3252 3256
rect 3502 3260 3508 3261
rect 3502 3256 3503 3260
rect 3507 3256 3508 3260
rect 3590 3259 3591 3263
rect 3595 3259 3596 3263
rect 3590 3258 3596 3259
rect 3502 3255 3508 3256
rect 1928 3235 1930 3255
rect 2064 3235 2066 3255
rect 2200 3235 2202 3255
rect 2360 3235 2362 3255
rect 2544 3235 2546 3255
rect 2760 3235 2762 3255
rect 3000 3235 3002 3255
rect 3248 3235 3250 3255
rect 3504 3235 3506 3255
rect 3592 3235 3594 3258
rect 1830 3232 1836 3233
rect 1871 3234 1875 3235
rect 1871 3229 1875 3230
rect 1895 3234 1899 3235
rect 1895 3229 1899 3230
rect 1927 3234 1931 3235
rect 1927 3229 1931 3230
rect 2007 3234 2011 3235
rect 2007 3229 2011 3230
rect 2063 3234 2067 3235
rect 2063 3229 2067 3230
rect 2143 3234 2147 3235
rect 2143 3229 2147 3230
rect 2199 3234 2203 3235
rect 2199 3229 2203 3230
rect 2279 3234 2283 3235
rect 2279 3229 2283 3230
rect 2359 3234 2363 3235
rect 2359 3229 2363 3230
rect 2415 3234 2419 3235
rect 2415 3229 2419 3230
rect 2543 3234 2547 3235
rect 2543 3229 2547 3230
rect 2567 3234 2571 3235
rect 2567 3229 2571 3230
rect 2727 3234 2731 3235
rect 2727 3229 2731 3230
rect 2759 3234 2763 3235
rect 2759 3229 2763 3230
rect 2911 3234 2915 3235
rect 2911 3229 2915 3230
rect 2999 3234 3003 3235
rect 2999 3229 3003 3230
rect 3103 3234 3107 3235
rect 3103 3229 3107 3230
rect 3247 3234 3251 3235
rect 3247 3229 3251 3230
rect 3311 3234 3315 3235
rect 3311 3229 3315 3230
rect 3503 3234 3507 3235
rect 3503 3229 3507 3230
rect 3591 3234 3595 3235
rect 3591 3229 3595 3230
rect 110 3220 116 3221
rect 110 3216 111 3220
rect 115 3216 116 3220
rect 110 3215 116 3216
rect 1830 3220 1836 3221
rect 1830 3216 1831 3220
rect 1835 3216 1836 3220
rect 1830 3215 1836 3216
rect 112 3179 114 3215
rect 390 3202 396 3203
rect 390 3198 391 3202
rect 395 3198 396 3202
rect 390 3197 396 3198
rect 478 3202 484 3203
rect 478 3198 479 3202
rect 483 3198 484 3202
rect 478 3197 484 3198
rect 582 3202 588 3203
rect 582 3198 583 3202
rect 587 3198 588 3202
rect 582 3197 588 3198
rect 694 3202 700 3203
rect 694 3198 695 3202
rect 699 3198 700 3202
rect 694 3197 700 3198
rect 814 3202 820 3203
rect 814 3198 815 3202
rect 819 3198 820 3202
rect 814 3197 820 3198
rect 942 3202 948 3203
rect 942 3198 943 3202
rect 947 3198 948 3202
rect 942 3197 948 3198
rect 1070 3202 1076 3203
rect 1070 3198 1071 3202
rect 1075 3198 1076 3202
rect 1070 3197 1076 3198
rect 1198 3202 1204 3203
rect 1198 3198 1199 3202
rect 1203 3198 1204 3202
rect 1198 3197 1204 3198
rect 1326 3202 1332 3203
rect 1326 3198 1327 3202
rect 1331 3198 1332 3202
rect 1326 3197 1332 3198
rect 1454 3202 1460 3203
rect 1454 3198 1455 3202
rect 1459 3198 1460 3202
rect 1454 3197 1460 3198
rect 1582 3202 1588 3203
rect 1582 3198 1583 3202
rect 1587 3198 1588 3202
rect 1582 3197 1588 3198
rect 392 3179 394 3197
rect 480 3179 482 3197
rect 584 3179 586 3197
rect 696 3179 698 3197
rect 816 3179 818 3197
rect 944 3179 946 3197
rect 1072 3179 1074 3197
rect 1200 3179 1202 3197
rect 1328 3179 1330 3197
rect 1456 3179 1458 3197
rect 1584 3179 1586 3197
rect 1832 3179 1834 3215
rect 1872 3210 1874 3229
rect 1896 3213 1898 3229
rect 2008 3213 2010 3229
rect 2144 3213 2146 3229
rect 2280 3213 2282 3229
rect 2416 3213 2418 3229
rect 2568 3213 2570 3229
rect 2728 3213 2730 3229
rect 2912 3213 2914 3229
rect 3104 3213 3106 3229
rect 3312 3213 3314 3229
rect 3504 3213 3506 3229
rect 1894 3212 1900 3213
rect 1870 3209 1876 3210
rect 1870 3205 1871 3209
rect 1875 3205 1876 3209
rect 1894 3208 1895 3212
rect 1899 3208 1900 3212
rect 1894 3207 1900 3208
rect 2006 3212 2012 3213
rect 2006 3208 2007 3212
rect 2011 3208 2012 3212
rect 2006 3207 2012 3208
rect 2142 3212 2148 3213
rect 2142 3208 2143 3212
rect 2147 3208 2148 3212
rect 2142 3207 2148 3208
rect 2278 3212 2284 3213
rect 2278 3208 2279 3212
rect 2283 3208 2284 3212
rect 2278 3207 2284 3208
rect 2414 3212 2420 3213
rect 2414 3208 2415 3212
rect 2419 3208 2420 3212
rect 2414 3207 2420 3208
rect 2566 3212 2572 3213
rect 2566 3208 2567 3212
rect 2571 3208 2572 3212
rect 2566 3207 2572 3208
rect 2726 3212 2732 3213
rect 2726 3208 2727 3212
rect 2731 3208 2732 3212
rect 2726 3207 2732 3208
rect 2910 3212 2916 3213
rect 2910 3208 2911 3212
rect 2915 3208 2916 3212
rect 2910 3207 2916 3208
rect 3102 3212 3108 3213
rect 3102 3208 3103 3212
rect 3107 3208 3108 3212
rect 3102 3207 3108 3208
rect 3310 3212 3316 3213
rect 3310 3208 3311 3212
rect 3315 3208 3316 3212
rect 3310 3207 3316 3208
rect 3502 3212 3508 3213
rect 3502 3208 3503 3212
rect 3507 3208 3508 3212
rect 3592 3210 3594 3229
rect 3502 3207 3508 3208
rect 3590 3209 3596 3210
rect 1870 3204 1876 3205
rect 3590 3205 3591 3209
rect 3595 3205 3596 3209
rect 3590 3204 3596 3205
rect 1870 3192 1876 3193
rect 1870 3188 1871 3192
rect 1875 3188 1876 3192
rect 1870 3187 1876 3188
rect 3590 3192 3596 3193
rect 3590 3188 3591 3192
rect 3595 3188 3596 3192
rect 3590 3187 3596 3188
rect 111 3178 115 3179
rect 111 3173 115 3174
rect 383 3178 387 3179
rect 383 3173 387 3174
rect 391 3178 395 3179
rect 391 3173 395 3174
rect 463 3178 467 3179
rect 463 3173 467 3174
rect 479 3178 483 3179
rect 479 3173 483 3174
rect 543 3178 547 3179
rect 543 3173 547 3174
rect 583 3178 587 3179
rect 583 3173 587 3174
rect 623 3178 627 3179
rect 623 3173 627 3174
rect 695 3178 699 3179
rect 695 3173 699 3174
rect 711 3178 715 3179
rect 711 3173 715 3174
rect 815 3178 819 3179
rect 815 3173 819 3174
rect 927 3178 931 3179
rect 927 3173 931 3174
rect 943 3178 947 3179
rect 943 3173 947 3174
rect 1039 3178 1043 3179
rect 1039 3173 1043 3174
rect 1071 3178 1075 3179
rect 1071 3173 1075 3174
rect 1159 3178 1163 3179
rect 1159 3173 1163 3174
rect 1199 3178 1203 3179
rect 1199 3173 1203 3174
rect 1271 3178 1275 3179
rect 1271 3173 1275 3174
rect 1327 3178 1331 3179
rect 1327 3173 1331 3174
rect 1383 3178 1387 3179
rect 1383 3173 1387 3174
rect 1455 3178 1459 3179
rect 1455 3173 1459 3174
rect 1495 3178 1499 3179
rect 1495 3173 1499 3174
rect 1583 3178 1587 3179
rect 1583 3173 1587 3174
rect 1615 3178 1619 3179
rect 1615 3173 1619 3174
rect 1735 3178 1739 3179
rect 1735 3173 1739 3174
rect 1831 3178 1835 3179
rect 1831 3173 1835 3174
rect 112 3145 114 3173
rect 384 3163 386 3173
rect 464 3163 466 3173
rect 544 3163 546 3173
rect 624 3163 626 3173
rect 712 3163 714 3173
rect 816 3163 818 3173
rect 928 3163 930 3173
rect 1040 3163 1042 3173
rect 1160 3163 1162 3173
rect 1272 3163 1274 3173
rect 1384 3163 1386 3173
rect 1496 3163 1498 3173
rect 1616 3163 1618 3173
rect 1736 3163 1738 3173
rect 382 3162 388 3163
rect 382 3158 383 3162
rect 387 3158 388 3162
rect 382 3157 388 3158
rect 462 3162 468 3163
rect 462 3158 463 3162
rect 467 3158 468 3162
rect 462 3157 468 3158
rect 542 3162 548 3163
rect 542 3158 543 3162
rect 547 3158 548 3162
rect 542 3157 548 3158
rect 622 3162 628 3163
rect 622 3158 623 3162
rect 627 3158 628 3162
rect 622 3157 628 3158
rect 710 3162 716 3163
rect 710 3158 711 3162
rect 715 3158 716 3162
rect 710 3157 716 3158
rect 814 3162 820 3163
rect 814 3158 815 3162
rect 819 3158 820 3162
rect 814 3157 820 3158
rect 926 3162 932 3163
rect 926 3158 927 3162
rect 931 3158 932 3162
rect 926 3157 932 3158
rect 1038 3162 1044 3163
rect 1038 3158 1039 3162
rect 1043 3158 1044 3162
rect 1038 3157 1044 3158
rect 1158 3162 1164 3163
rect 1158 3158 1159 3162
rect 1163 3158 1164 3162
rect 1158 3157 1164 3158
rect 1270 3162 1276 3163
rect 1270 3158 1271 3162
rect 1275 3158 1276 3162
rect 1270 3157 1276 3158
rect 1382 3162 1388 3163
rect 1382 3158 1383 3162
rect 1387 3158 1388 3162
rect 1382 3157 1388 3158
rect 1494 3162 1500 3163
rect 1494 3158 1495 3162
rect 1499 3158 1500 3162
rect 1494 3157 1500 3158
rect 1614 3162 1620 3163
rect 1614 3158 1615 3162
rect 1619 3158 1620 3162
rect 1614 3157 1620 3158
rect 1734 3162 1740 3163
rect 1734 3158 1735 3162
rect 1739 3158 1740 3162
rect 1734 3157 1740 3158
rect 1832 3145 1834 3173
rect 1872 3159 1874 3187
rect 1902 3174 1908 3175
rect 1902 3170 1903 3174
rect 1907 3170 1908 3174
rect 1902 3169 1908 3170
rect 2014 3174 2020 3175
rect 2014 3170 2015 3174
rect 2019 3170 2020 3174
rect 2014 3169 2020 3170
rect 2150 3174 2156 3175
rect 2150 3170 2151 3174
rect 2155 3170 2156 3174
rect 2150 3169 2156 3170
rect 2286 3174 2292 3175
rect 2286 3170 2287 3174
rect 2291 3170 2292 3174
rect 2286 3169 2292 3170
rect 2422 3174 2428 3175
rect 2422 3170 2423 3174
rect 2427 3170 2428 3174
rect 2422 3169 2428 3170
rect 2574 3174 2580 3175
rect 2574 3170 2575 3174
rect 2579 3170 2580 3174
rect 2574 3169 2580 3170
rect 2734 3174 2740 3175
rect 2734 3170 2735 3174
rect 2739 3170 2740 3174
rect 2734 3169 2740 3170
rect 2918 3174 2924 3175
rect 2918 3170 2919 3174
rect 2923 3170 2924 3174
rect 2918 3169 2924 3170
rect 3110 3174 3116 3175
rect 3110 3170 3111 3174
rect 3115 3170 3116 3174
rect 3110 3169 3116 3170
rect 3318 3174 3324 3175
rect 3318 3170 3319 3174
rect 3323 3170 3324 3174
rect 3318 3169 3324 3170
rect 3510 3174 3516 3175
rect 3510 3170 3511 3174
rect 3515 3170 3516 3174
rect 3510 3169 3516 3170
rect 1904 3159 1906 3169
rect 2016 3159 2018 3169
rect 2152 3159 2154 3169
rect 2288 3159 2290 3169
rect 2424 3159 2426 3169
rect 2576 3159 2578 3169
rect 2736 3159 2738 3169
rect 2920 3159 2922 3169
rect 3112 3159 3114 3169
rect 3320 3159 3322 3169
rect 3512 3159 3514 3169
rect 3592 3159 3594 3187
rect 1871 3158 1875 3159
rect 1871 3153 1875 3154
rect 1903 3158 1907 3159
rect 1903 3153 1907 3154
rect 2015 3158 2019 3159
rect 2015 3153 2019 3154
rect 2079 3158 2083 3159
rect 2079 3153 2083 3154
rect 2151 3158 2155 3159
rect 2151 3153 2155 3154
rect 2271 3158 2275 3159
rect 2271 3153 2275 3154
rect 2287 3158 2291 3159
rect 2287 3153 2291 3154
rect 2423 3158 2427 3159
rect 2423 3153 2427 3154
rect 2455 3158 2459 3159
rect 2455 3153 2459 3154
rect 2575 3158 2579 3159
rect 2575 3153 2579 3154
rect 2623 3158 2627 3159
rect 2623 3153 2627 3154
rect 2735 3158 2739 3159
rect 2735 3153 2739 3154
rect 2783 3158 2787 3159
rect 2783 3153 2787 3154
rect 2919 3158 2923 3159
rect 2919 3153 2923 3154
rect 2935 3158 2939 3159
rect 2935 3153 2939 3154
rect 3079 3158 3083 3159
rect 3079 3153 3083 3154
rect 3111 3158 3115 3159
rect 3111 3153 3115 3154
rect 3231 3158 3235 3159
rect 3231 3153 3235 3154
rect 3319 3158 3323 3159
rect 3319 3153 3323 3154
rect 3511 3158 3515 3159
rect 3511 3153 3515 3154
rect 3591 3158 3595 3159
rect 3591 3153 3595 3154
rect 110 3144 116 3145
rect 110 3140 111 3144
rect 115 3140 116 3144
rect 110 3139 116 3140
rect 1830 3144 1836 3145
rect 1830 3140 1831 3144
rect 1835 3140 1836 3144
rect 1830 3139 1836 3140
rect 110 3127 116 3128
rect 110 3123 111 3127
rect 115 3123 116 3127
rect 1830 3127 1836 3128
rect 110 3122 116 3123
rect 374 3124 380 3125
rect 112 3103 114 3122
rect 374 3120 375 3124
rect 379 3120 380 3124
rect 374 3119 380 3120
rect 454 3124 460 3125
rect 454 3120 455 3124
rect 459 3120 460 3124
rect 454 3119 460 3120
rect 534 3124 540 3125
rect 534 3120 535 3124
rect 539 3120 540 3124
rect 534 3119 540 3120
rect 614 3124 620 3125
rect 614 3120 615 3124
rect 619 3120 620 3124
rect 614 3119 620 3120
rect 702 3124 708 3125
rect 702 3120 703 3124
rect 707 3120 708 3124
rect 702 3119 708 3120
rect 806 3124 812 3125
rect 806 3120 807 3124
rect 811 3120 812 3124
rect 806 3119 812 3120
rect 918 3124 924 3125
rect 918 3120 919 3124
rect 923 3120 924 3124
rect 918 3119 924 3120
rect 1030 3124 1036 3125
rect 1030 3120 1031 3124
rect 1035 3120 1036 3124
rect 1030 3119 1036 3120
rect 1150 3124 1156 3125
rect 1150 3120 1151 3124
rect 1155 3120 1156 3124
rect 1150 3119 1156 3120
rect 1262 3124 1268 3125
rect 1262 3120 1263 3124
rect 1267 3120 1268 3124
rect 1262 3119 1268 3120
rect 1374 3124 1380 3125
rect 1374 3120 1375 3124
rect 1379 3120 1380 3124
rect 1374 3119 1380 3120
rect 1486 3124 1492 3125
rect 1486 3120 1487 3124
rect 1491 3120 1492 3124
rect 1486 3119 1492 3120
rect 1606 3124 1612 3125
rect 1606 3120 1607 3124
rect 1611 3120 1612 3124
rect 1606 3119 1612 3120
rect 1726 3124 1732 3125
rect 1726 3120 1727 3124
rect 1731 3120 1732 3124
rect 1830 3123 1831 3127
rect 1835 3123 1836 3127
rect 1872 3125 1874 3153
rect 1904 3143 1906 3153
rect 2080 3143 2082 3153
rect 2272 3143 2274 3153
rect 2456 3143 2458 3153
rect 2624 3143 2626 3153
rect 2784 3143 2786 3153
rect 2936 3143 2938 3153
rect 3080 3143 3082 3153
rect 3232 3143 3234 3153
rect 1902 3142 1908 3143
rect 1902 3138 1903 3142
rect 1907 3138 1908 3142
rect 1902 3137 1908 3138
rect 2078 3142 2084 3143
rect 2078 3138 2079 3142
rect 2083 3138 2084 3142
rect 2078 3137 2084 3138
rect 2270 3142 2276 3143
rect 2270 3138 2271 3142
rect 2275 3138 2276 3142
rect 2270 3137 2276 3138
rect 2454 3142 2460 3143
rect 2454 3138 2455 3142
rect 2459 3138 2460 3142
rect 2454 3137 2460 3138
rect 2622 3142 2628 3143
rect 2622 3138 2623 3142
rect 2627 3138 2628 3142
rect 2622 3137 2628 3138
rect 2782 3142 2788 3143
rect 2782 3138 2783 3142
rect 2787 3138 2788 3142
rect 2782 3137 2788 3138
rect 2934 3142 2940 3143
rect 2934 3138 2935 3142
rect 2939 3138 2940 3142
rect 2934 3137 2940 3138
rect 3078 3142 3084 3143
rect 3078 3138 3079 3142
rect 3083 3138 3084 3142
rect 3078 3137 3084 3138
rect 3230 3142 3236 3143
rect 3230 3138 3231 3142
rect 3235 3138 3236 3142
rect 3230 3137 3236 3138
rect 3592 3125 3594 3153
rect 1830 3122 1836 3123
rect 1870 3124 1876 3125
rect 1726 3119 1732 3120
rect 376 3103 378 3119
rect 456 3103 458 3119
rect 536 3103 538 3119
rect 616 3103 618 3119
rect 704 3103 706 3119
rect 808 3103 810 3119
rect 920 3103 922 3119
rect 1032 3103 1034 3119
rect 1152 3103 1154 3119
rect 1264 3103 1266 3119
rect 1376 3103 1378 3119
rect 1488 3103 1490 3119
rect 1608 3103 1610 3119
rect 1728 3103 1730 3119
rect 1832 3103 1834 3122
rect 1870 3120 1871 3124
rect 1875 3120 1876 3124
rect 1870 3119 1876 3120
rect 3590 3124 3596 3125
rect 3590 3120 3591 3124
rect 3595 3120 3596 3124
rect 3590 3119 3596 3120
rect 1870 3107 1876 3108
rect 1870 3103 1871 3107
rect 1875 3103 1876 3107
rect 3590 3107 3596 3108
rect 111 3102 115 3103
rect 111 3097 115 3098
rect 375 3102 379 3103
rect 375 3097 379 3098
rect 455 3102 459 3103
rect 455 3097 459 3098
rect 535 3102 539 3103
rect 535 3097 539 3098
rect 615 3102 619 3103
rect 615 3097 619 3098
rect 703 3102 707 3103
rect 703 3097 707 3098
rect 807 3102 811 3103
rect 807 3097 811 3098
rect 919 3102 923 3103
rect 919 3097 923 3098
rect 943 3102 947 3103
rect 943 3097 947 3098
rect 1023 3102 1027 3103
rect 1023 3097 1027 3098
rect 1031 3102 1035 3103
rect 1031 3097 1035 3098
rect 1103 3102 1107 3103
rect 1103 3097 1107 3098
rect 1151 3102 1155 3103
rect 1151 3097 1155 3098
rect 1183 3102 1187 3103
rect 1183 3097 1187 3098
rect 1263 3102 1267 3103
rect 1263 3097 1267 3098
rect 1343 3102 1347 3103
rect 1343 3097 1347 3098
rect 1375 3102 1379 3103
rect 1375 3097 1379 3098
rect 1423 3102 1427 3103
rect 1423 3097 1427 3098
rect 1487 3102 1491 3103
rect 1487 3097 1491 3098
rect 1503 3102 1507 3103
rect 1503 3097 1507 3098
rect 1583 3102 1587 3103
rect 1583 3097 1587 3098
rect 1607 3102 1611 3103
rect 1607 3097 1611 3098
rect 1663 3102 1667 3103
rect 1663 3097 1667 3098
rect 1727 3102 1731 3103
rect 1727 3097 1731 3098
rect 1743 3102 1747 3103
rect 1743 3097 1747 3098
rect 1831 3102 1835 3103
rect 1870 3102 1876 3103
rect 1894 3104 1900 3105
rect 1831 3097 1835 3098
rect 112 3078 114 3097
rect 944 3081 946 3097
rect 1024 3081 1026 3097
rect 1104 3081 1106 3097
rect 1184 3081 1186 3097
rect 1264 3081 1266 3097
rect 1344 3081 1346 3097
rect 1424 3081 1426 3097
rect 1504 3081 1506 3097
rect 1584 3081 1586 3097
rect 1664 3081 1666 3097
rect 1744 3081 1746 3097
rect 942 3080 948 3081
rect 110 3077 116 3078
rect 110 3073 111 3077
rect 115 3073 116 3077
rect 942 3076 943 3080
rect 947 3076 948 3080
rect 942 3075 948 3076
rect 1022 3080 1028 3081
rect 1022 3076 1023 3080
rect 1027 3076 1028 3080
rect 1022 3075 1028 3076
rect 1102 3080 1108 3081
rect 1102 3076 1103 3080
rect 1107 3076 1108 3080
rect 1102 3075 1108 3076
rect 1182 3080 1188 3081
rect 1182 3076 1183 3080
rect 1187 3076 1188 3080
rect 1182 3075 1188 3076
rect 1262 3080 1268 3081
rect 1262 3076 1263 3080
rect 1267 3076 1268 3080
rect 1262 3075 1268 3076
rect 1342 3080 1348 3081
rect 1342 3076 1343 3080
rect 1347 3076 1348 3080
rect 1342 3075 1348 3076
rect 1422 3080 1428 3081
rect 1422 3076 1423 3080
rect 1427 3076 1428 3080
rect 1422 3075 1428 3076
rect 1502 3080 1508 3081
rect 1502 3076 1503 3080
rect 1507 3076 1508 3080
rect 1502 3075 1508 3076
rect 1582 3080 1588 3081
rect 1582 3076 1583 3080
rect 1587 3076 1588 3080
rect 1582 3075 1588 3076
rect 1662 3080 1668 3081
rect 1662 3076 1663 3080
rect 1667 3076 1668 3080
rect 1662 3075 1668 3076
rect 1742 3080 1748 3081
rect 1742 3076 1743 3080
rect 1747 3076 1748 3080
rect 1832 3078 1834 3097
rect 1742 3075 1748 3076
rect 1830 3077 1836 3078
rect 110 3072 116 3073
rect 1830 3073 1831 3077
rect 1835 3073 1836 3077
rect 1872 3075 1874 3102
rect 1894 3100 1895 3104
rect 1899 3100 1900 3104
rect 1894 3099 1900 3100
rect 2070 3104 2076 3105
rect 2070 3100 2071 3104
rect 2075 3100 2076 3104
rect 2070 3099 2076 3100
rect 2262 3104 2268 3105
rect 2262 3100 2263 3104
rect 2267 3100 2268 3104
rect 2262 3099 2268 3100
rect 2446 3104 2452 3105
rect 2446 3100 2447 3104
rect 2451 3100 2452 3104
rect 2446 3099 2452 3100
rect 2614 3104 2620 3105
rect 2614 3100 2615 3104
rect 2619 3100 2620 3104
rect 2614 3099 2620 3100
rect 2774 3104 2780 3105
rect 2774 3100 2775 3104
rect 2779 3100 2780 3104
rect 2774 3099 2780 3100
rect 2926 3104 2932 3105
rect 2926 3100 2927 3104
rect 2931 3100 2932 3104
rect 2926 3099 2932 3100
rect 3070 3104 3076 3105
rect 3070 3100 3071 3104
rect 3075 3100 3076 3104
rect 3070 3099 3076 3100
rect 3222 3104 3228 3105
rect 3222 3100 3223 3104
rect 3227 3100 3228 3104
rect 3590 3103 3591 3107
rect 3595 3103 3596 3107
rect 3590 3102 3596 3103
rect 3222 3099 3228 3100
rect 1896 3075 1898 3099
rect 2072 3075 2074 3099
rect 2264 3075 2266 3099
rect 2448 3075 2450 3099
rect 2616 3075 2618 3099
rect 2776 3075 2778 3099
rect 2928 3075 2930 3099
rect 3072 3075 3074 3099
rect 3224 3075 3226 3099
rect 3592 3075 3594 3102
rect 1830 3072 1836 3073
rect 1871 3074 1875 3075
rect 1871 3069 1875 3070
rect 1895 3074 1899 3075
rect 1895 3069 1899 3070
rect 1991 3074 1995 3075
rect 1991 3069 1995 3070
rect 2071 3074 2075 3075
rect 2071 3069 2075 3070
rect 2247 3074 2251 3075
rect 2247 3069 2251 3070
rect 2263 3074 2267 3075
rect 2263 3069 2267 3070
rect 2447 3074 2451 3075
rect 2447 3069 2451 3070
rect 2487 3074 2491 3075
rect 2487 3069 2491 3070
rect 2615 3074 2619 3075
rect 2615 3069 2619 3070
rect 2703 3074 2707 3075
rect 2703 3069 2707 3070
rect 2775 3074 2779 3075
rect 2775 3069 2779 3070
rect 2895 3074 2899 3075
rect 2895 3069 2899 3070
rect 2927 3074 2931 3075
rect 2927 3069 2931 3070
rect 3063 3074 3067 3075
rect 3063 3069 3067 3070
rect 3071 3074 3075 3075
rect 3071 3069 3075 3070
rect 3223 3074 3227 3075
rect 3223 3069 3227 3070
rect 3375 3074 3379 3075
rect 3375 3069 3379 3070
rect 3503 3074 3507 3075
rect 3503 3069 3507 3070
rect 3591 3074 3595 3075
rect 3591 3069 3595 3070
rect 110 3060 116 3061
rect 110 3056 111 3060
rect 115 3056 116 3060
rect 110 3055 116 3056
rect 1830 3060 1836 3061
rect 1830 3056 1831 3060
rect 1835 3056 1836 3060
rect 1830 3055 1836 3056
rect 112 3011 114 3055
rect 950 3042 956 3043
rect 950 3038 951 3042
rect 955 3038 956 3042
rect 950 3037 956 3038
rect 1030 3042 1036 3043
rect 1030 3038 1031 3042
rect 1035 3038 1036 3042
rect 1030 3037 1036 3038
rect 1110 3042 1116 3043
rect 1110 3038 1111 3042
rect 1115 3038 1116 3042
rect 1110 3037 1116 3038
rect 1190 3042 1196 3043
rect 1190 3038 1191 3042
rect 1195 3038 1196 3042
rect 1190 3037 1196 3038
rect 1270 3042 1276 3043
rect 1270 3038 1271 3042
rect 1275 3038 1276 3042
rect 1270 3037 1276 3038
rect 1350 3042 1356 3043
rect 1350 3038 1351 3042
rect 1355 3038 1356 3042
rect 1350 3037 1356 3038
rect 1430 3042 1436 3043
rect 1430 3038 1431 3042
rect 1435 3038 1436 3042
rect 1430 3037 1436 3038
rect 1510 3042 1516 3043
rect 1510 3038 1511 3042
rect 1515 3038 1516 3042
rect 1510 3037 1516 3038
rect 1590 3042 1596 3043
rect 1590 3038 1591 3042
rect 1595 3038 1596 3042
rect 1590 3037 1596 3038
rect 1670 3042 1676 3043
rect 1670 3038 1671 3042
rect 1675 3038 1676 3042
rect 1670 3037 1676 3038
rect 1750 3042 1756 3043
rect 1750 3038 1751 3042
rect 1755 3038 1756 3042
rect 1750 3037 1756 3038
rect 952 3011 954 3037
rect 1032 3011 1034 3037
rect 1112 3011 1114 3037
rect 1192 3011 1194 3037
rect 1272 3011 1274 3037
rect 1352 3011 1354 3037
rect 1432 3011 1434 3037
rect 1512 3011 1514 3037
rect 1592 3011 1594 3037
rect 1672 3011 1674 3037
rect 1752 3011 1754 3037
rect 1832 3011 1834 3055
rect 1872 3050 1874 3069
rect 1992 3053 1994 3069
rect 2248 3053 2250 3069
rect 2488 3053 2490 3069
rect 2704 3053 2706 3069
rect 2896 3053 2898 3069
rect 3064 3053 3066 3069
rect 3224 3053 3226 3069
rect 3376 3053 3378 3069
rect 3504 3053 3506 3069
rect 1990 3052 1996 3053
rect 1870 3049 1876 3050
rect 1870 3045 1871 3049
rect 1875 3045 1876 3049
rect 1990 3048 1991 3052
rect 1995 3048 1996 3052
rect 1990 3047 1996 3048
rect 2246 3052 2252 3053
rect 2246 3048 2247 3052
rect 2251 3048 2252 3052
rect 2246 3047 2252 3048
rect 2486 3052 2492 3053
rect 2486 3048 2487 3052
rect 2491 3048 2492 3052
rect 2486 3047 2492 3048
rect 2702 3052 2708 3053
rect 2702 3048 2703 3052
rect 2707 3048 2708 3052
rect 2702 3047 2708 3048
rect 2894 3052 2900 3053
rect 2894 3048 2895 3052
rect 2899 3048 2900 3052
rect 2894 3047 2900 3048
rect 3062 3052 3068 3053
rect 3062 3048 3063 3052
rect 3067 3048 3068 3052
rect 3062 3047 3068 3048
rect 3222 3052 3228 3053
rect 3222 3048 3223 3052
rect 3227 3048 3228 3052
rect 3222 3047 3228 3048
rect 3374 3052 3380 3053
rect 3374 3048 3375 3052
rect 3379 3048 3380 3052
rect 3374 3047 3380 3048
rect 3502 3052 3508 3053
rect 3502 3048 3503 3052
rect 3507 3048 3508 3052
rect 3592 3050 3594 3069
rect 3502 3047 3508 3048
rect 3590 3049 3596 3050
rect 1870 3044 1876 3045
rect 3590 3045 3591 3049
rect 3595 3045 3596 3049
rect 3590 3044 3596 3045
rect 1870 3032 1876 3033
rect 1870 3028 1871 3032
rect 1875 3028 1876 3032
rect 1870 3027 1876 3028
rect 3590 3032 3596 3033
rect 3590 3028 3591 3032
rect 3595 3028 3596 3032
rect 3590 3027 3596 3028
rect 111 3010 115 3011
rect 111 3005 115 3006
rect 207 3010 211 3011
rect 207 3005 211 3006
rect 327 3010 331 3011
rect 327 3005 331 3006
rect 471 3010 475 3011
rect 471 3005 475 3006
rect 631 3010 635 3011
rect 631 3005 635 3006
rect 807 3010 811 3011
rect 807 3005 811 3006
rect 951 3010 955 3011
rect 951 3005 955 3006
rect 983 3010 987 3011
rect 983 3005 987 3006
rect 1031 3010 1035 3011
rect 1031 3005 1035 3006
rect 1111 3010 1115 3011
rect 1111 3005 1115 3006
rect 1151 3010 1155 3011
rect 1151 3005 1155 3006
rect 1191 3010 1195 3011
rect 1191 3005 1195 3006
rect 1271 3010 1275 3011
rect 1271 3005 1275 3006
rect 1311 3010 1315 3011
rect 1311 3005 1315 3006
rect 1351 3010 1355 3011
rect 1351 3005 1355 3006
rect 1431 3010 1435 3011
rect 1431 3005 1435 3006
rect 1463 3010 1467 3011
rect 1463 3005 1467 3006
rect 1511 3010 1515 3011
rect 1511 3005 1515 3006
rect 1591 3010 1595 3011
rect 1591 3005 1595 3006
rect 1615 3010 1619 3011
rect 1615 3005 1619 3006
rect 1671 3010 1675 3011
rect 1671 3005 1675 3006
rect 1751 3010 1755 3011
rect 1751 3005 1755 3006
rect 1831 3010 1835 3011
rect 1831 3005 1835 3006
rect 112 2977 114 3005
rect 208 2995 210 3005
rect 328 2995 330 3005
rect 472 2995 474 3005
rect 632 2995 634 3005
rect 808 2995 810 3005
rect 984 2995 986 3005
rect 1152 2995 1154 3005
rect 1312 2995 1314 3005
rect 1464 2995 1466 3005
rect 1616 2995 1618 3005
rect 1752 2995 1754 3005
rect 206 2994 212 2995
rect 206 2990 207 2994
rect 211 2990 212 2994
rect 206 2989 212 2990
rect 326 2994 332 2995
rect 326 2990 327 2994
rect 331 2990 332 2994
rect 326 2989 332 2990
rect 470 2994 476 2995
rect 470 2990 471 2994
rect 475 2990 476 2994
rect 470 2989 476 2990
rect 630 2994 636 2995
rect 630 2990 631 2994
rect 635 2990 636 2994
rect 630 2989 636 2990
rect 806 2994 812 2995
rect 806 2990 807 2994
rect 811 2990 812 2994
rect 806 2989 812 2990
rect 982 2994 988 2995
rect 982 2990 983 2994
rect 987 2990 988 2994
rect 982 2989 988 2990
rect 1150 2994 1156 2995
rect 1150 2990 1151 2994
rect 1155 2990 1156 2994
rect 1150 2989 1156 2990
rect 1310 2994 1316 2995
rect 1310 2990 1311 2994
rect 1315 2990 1316 2994
rect 1310 2989 1316 2990
rect 1462 2994 1468 2995
rect 1462 2990 1463 2994
rect 1467 2990 1468 2994
rect 1462 2989 1468 2990
rect 1614 2994 1620 2995
rect 1614 2990 1615 2994
rect 1619 2990 1620 2994
rect 1614 2989 1620 2990
rect 1750 2994 1756 2995
rect 1750 2990 1751 2994
rect 1755 2990 1756 2994
rect 1750 2989 1756 2990
rect 1832 2977 1834 3005
rect 1872 2995 1874 3027
rect 1998 3014 2004 3015
rect 1998 3010 1999 3014
rect 2003 3010 2004 3014
rect 1998 3009 2004 3010
rect 2254 3014 2260 3015
rect 2254 3010 2255 3014
rect 2259 3010 2260 3014
rect 2254 3009 2260 3010
rect 2494 3014 2500 3015
rect 2494 3010 2495 3014
rect 2499 3010 2500 3014
rect 2494 3009 2500 3010
rect 2710 3014 2716 3015
rect 2710 3010 2711 3014
rect 2715 3010 2716 3014
rect 2710 3009 2716 3010
rect 2902 3014 2908 3015
rect 2902 3010 2903 3014
rect 2907 3010 2908 3014
rect 2902 3009 2908 3010
rect 3070 3014 3076 3015
rect 3070 3010 3071 3014
rect 3075 3010 3076 3014
rect 3070 3009 3076 3010
rect 3230 3014 3236 3015
rect 3230 3010 3231 3014
rect 3235 3010 3236 3014
rect 3230 3009 3236 3010
rect 3382 3014 3388 3015
rect 3382 3010 3383 3014
rect 3387 3010 3388 3014
rect 3382 3009 3388 3010
rect 3510 3014 3516 3015
rect 3510 3010 3511 3014
rect 3515 3010 3516 3014
rect 3510 3009 3516 3010
rect 2000 2995 2002 3009
rect 2256 2995 2258 3009
rect 2496 2995 2498 3009
rect 2712 2995 2714 3009
rect 2904 2995 2906 3009
rect 3072 2995 3074 3009
rect 3232 2995 3234 3009
rect 3384 2995 3386 3009
rect 3512 2995 3514 3009
rect 3592 2995 3594 3027
rect 1871 2994 1875 2995
rect 1871 2989 1875 2990
rect 1903 2994 1907 2995
rect 1903 2989 1907 2990
rect 1999 2994 2003 2995
rect 1999 2989 2003 2990
rect 2143 2994 2147 2995
rect 2143 2989 2147 2990
rect 2255 2994 2259 2995
rect 2255 2989 2259 2990
rect 2391 2994 2395 2995
rect 2391 2989 2395 2990
rect 2495 2994 2499 2995
rect 2495 2989 2499 2990
rect 2607 2994 2611 2995
rect 2607 2989 2611 2990
rect 2711 2994 2715 2995
rect 2711 2989 2715 2990
rect 2799 2994 2803 2995
rect 2799 2989 2803 2990
rect 2903 2994 2907 2995
rect 2903 2989 2907 2990
rect 2967 2994 2971 2995
rect 2967 2989 2971 2990
rect 3071 2994 3075 2995
rect 3071 2989 3075 2990
rect 3119 2994 3123 2995
rect 3119 2989 3123 2990
rect 3231 2994 3235 2995
rect 3231 2989 3235 2990
rect 3263 2994 3267 2995
rect 3263 2989 3267 2990
rect 3383 2994 3387 2995
rect 3383 2989 3387 2990
rect 3399 2994 3403 2995
rect 3399 2989 3403 2990
rect 3511 2994 3515 2995
rect 3511 2989 3515 2990
rect 3591 2994 3595 2995
rect 3591 2989 3595 2990
rect 110 2976 116 2977
rect 110 2972 111 2976
rect 115 2972 116 2976
rect 110 2971 116 2972
rect 1830 2976 1836 2977
rect 1830 2972 1831 2976
rect 1835 2972 1836 2976
rect 1830 2971 1836 2972
rect 1872 2961 1874 2989
rect 1904 2979 1906 2989
rect 2144 2979 2146 2989
rect 2392 2979 2394 2989
rect 2608 2979 2610 2989
rect 2800 2979 2802 2989
rect 2968 2979 2970 2989
rect 3120 2979 3122 2989
rect 3264 2979 3266 2989
rect 3400 2979 3402 2989
rect 3512 2979 3514 2989
rect 1902 2978 1908 2979
rect 1902 2974 1903 2978
rect 1907 2974 1908 2978
rect 1902 2973 1908 2974
rect 2142 2978 2148 2979
rect 2142 2974 2143 2978
rect 2147 2974 2148 2978
rect 2142 2973 2148 2974
rect 2390 2978 2396 2979
rect 2390 2974 2391 2978
rect 2395 2974 2396 2978
rect 2390 2973 2396 2974
rect 2606 2978 2612 2979
rect 2606 2974 2607 2978
rect 2611 2974 2612 2978
rect 2606 2973 2612 2974
rect 2798 2978 2804 2979
rect 2798 2974 2799 2978
rect 2803 2974 2804 2978
rect 2798 2973 2804 2974
rect 2966 2978 2972 2979
rect 2966 2974 2967 2978
rect 2971 2974 2972 2978
rect 2966 2973 2972 2974
rect 3118 2978 3124 2979
rect 3118 2974 3119 2978
rect 3123 2974 3124 2978
rect 3118 2973 3124 2974
rect 3262 2978 3268 2979
rect 3262 2974 3263 2978
rect 3267 2974 3268 2978
rect 3262 2973 3268 2974
rect 3398 2978 3404 2979
rect 3398 2974 3399 2978
rect 3403 2974 3404 2978
rect 3398 2973 3404 2974
rect 3510 2978 3516 2979
rect 3510 2974 3511 2978
rect 3515 2974 3516 2978
rect 3510 2973 3516 2974
rect 3592 2961 3594 2989
rect 1870 2960 1876 2961
rect 110 2959 116 2960
rect 110 2955 111 2959
rect 115 2955 116 2959
rect 1830 2959 1836 2960
rect 110 2954 116 2955
rect 198 2956 204 2957
rect 112 2935 114 2954
rect 198 2952 199 2956
rect 203 2952 204 2956
rect 198 2951 204 2952
rect 318 2956 324 2957
rect 318 2952 319 2956
rect 323 2952 324 2956
rect 318 2951 324 2952
rect 462 2956 468 2957
rect 462 2952 463 2956
rect 467 2952 468 2956
rect 462 2951 468 2952
rect 622 2956 628 2957
rect 622 2952 623 2956
rect 627 2952 628 2956
rect 622 2951 628 2952
rect 798 2956 804 2957
rect 798 2952 799 2956
rect 803 2952 804 2956
rect 798 2951 804 2952
rect 974 2956 980 2957
rect 974 2952 975 2956
rect 979 2952 980 2956
rect 974 2951 980 2952
rect 1142 2956 1148 2957
rect 1142 2952 1143 2956
rect 1147 2952 1148 2956
rect 1142 2951 1148 2952
rect 1302 2956 1308 2957
rect 1302 2952 1303 2956
rect 1307 2952 1308 2956
rect 1302 2951 1308 2952
rect 1454 2956 1460 2957
rect 1454 2952 1455 2956
rect 1459 2952 1460 2956
rect 1454 2951 1460 2952
rect 1606 2956 1612 2957
rect 1606 2952 1607 2956
rect 1611 2952 1612 2956
rect 1606 2951 1612 2952
rect 1742 2956 1748 2957
rect 1742 2952 1743 2956
rect 1747 2952 1748 2956
rect 1830 2955 1831 2959
rect 1835 2955 1836 2959
rect 1870 2956 1871 2960
rect 1875 2956 1876 2960
rect 1870 2955 1876 2956
rect 3590 2960 3596 2961
rect 3590 2956 3591 2960
rect 3595 2956 3596 2960
rect 3590 2955 3596 2956
rect 1830 2954 1836 2955
rect 1742 2951 1748 2952
rect 200 2935 202 2951
rect 320 2935 322 2951
rect 464 2935 466 2951
rect 624 2935 626 2951
rect 800 2935 802 2951
rect 976 2935 978 2951
rect 1144 2935 1146 2951
rect 1304 2935 1306 2951
rect 1456 2935 1458 2951
rect 1608 2935 1610 2951
rect 1744 2935 1746 2951
rect 1832 2935 1834 2954
rect 1870 2943 1876 2944
rect 1870 2939 1871 2943
rect 1875 2939 1876 2943
rect 3590 2943 3596 2944
rect 1870 2938 1876 2939
rect 1894 2940 1900 2941
rect 111 2934 115 2935
rect 111 2929 115 2930
rect 199 2934 203 2935
rect 199 2929 203 2930
rect 247 2934 251 2935
rect 247 2929 251 2930
rect 319 2934 323 2935
rect 319 2929 323 2930
rect 351 2934 355 2935
rect 351 2929 355 2930
rect 463 2934 467 2935
rect 463 2929 467 2930
rect 471 2934 475 2935
rect 471 2929 475 2930
rect 607 2934 611 2935
rect 607 2929 611 2930
rect 623 2934 627 2935
rect 623 2929 627 2930
rect 751 2934 755 2935
rect 751 2929 755 2930
rect 799 2934 803 2935
rect 799 2929 803 2930
rect 895 2934 899 2935
rect 895 2929 899 2930
rect 975 2934 979 2935
rect 975 2929 979 2930
rect 1031 2934 1035 2935
rect 1031 2929 1035 2930
rect 1143 2934 1147 2935
rect 1143 2929 1147 2930
rect 1159 2934 1163 2935
rect 1159 2929 1163 2930
rect 1279 2934 1283 2935
rect 1279 2929 1283 2930
rect 1303 2934 1307 2935
rect 1303 2929 1307 2930
rect 1399 2934 1403 2935
rect 1399 2929 1403 2930
rect 1455 2934 1459 2935
rect 1455 2929 1459 2930
rect 1519 2934 1523 2935
rect 1519 2929 1523 2930
rect 1607 2934 1611 2935
rect 1607 2929 1611 2930
rect 1639 2934 1643 2935
rect 1639 2929 1643 2930
rect 1743 2934 1747 2935
rect 1743 2929 1747 2930
rect 1831 2934 1835 2935
rect 1831 2929 1835 2930
rect 112 2910 114 2929
rect 248 2913 250 2929
rect 352 2913 354 2929
rect 472 2913 474 2929
rect 608 2913 610 2929
rect 752 2913 754 2929
rect 896 2913 898 2929
rect 1032 2913 1034 2929
rect 1160 2913 1162 2929
rect 1280 2913 1282 2929
rect 1400 2913 1402 2929
rect 1520 2913 1522 2929
rect 1640 2913 1642 2929
rect 246 2912 252 2913
rect 110 2909 116 2910
rect 110 2905 111 2909
rect 115 2905 116 2909
rect 246 2908 247 2912
rect 251 2908 252 2912
rect 246 2907 252 2908
rect 350 2912 356 2913
rect 350 2908 351 2912
rect 355 2908 356 2912
rect 350 2907 356 2908
rect 470 2912 476 2913
rect 470 2908 471 2912
rect 475 2908 476 2912
rect 470 2907 476 2908
rect 606 2912 612 2913
rect 606 2908 607 2912
rect 611 2908 612 2912
rect 606 2907 612 2908
rect 750 2912 756 2913
rect 750 2908 751 2912
rect 755 2908 756 2912
rect 750 2907 756 2908
rect 894 2912 900 2913
rect 894 2908 895 2912
rect 899 2908 900 2912
rect 894 2907 900 2908
rect 1030 2912 1036 2913
rect 1030 2908 1031 2912
rect 1035 2908 1036 2912
rect 1030 2907 1036 2908
rect 1158 2912 1164 2913
rect 1158 2908 1159 2912
rect 1163 2908 1164 2912
rect 1158 2907 1164 2908
rect 1278 2912 1284 2913
rect 1278 2908 1279 2912
rect 1283 2908 1284 2912
rect 1278 2907 1284 2908
rect 1398 2912 1404 2913
rect 1398 2908 1399 2912
rect 1403 2908 1404 2912
rect 1398 2907 1404 2908
rect 1518 2912 1524 2913
rect 1518 2908 1519 2912
rect 1523 2908 1524 2912
rect 1518 2907 1524 2908
rect 1638 2912 1644 2913
rect 1638 2908 1639 2912
rect 1643 2908 1644 2912
rect 1832 2910 1834 2929
rect 1638 2907 1644 2908
rect 1830 2909 1836 2910
rect 110 2904 116 2905
rect 1830 2905 1831 2909
rect 1835 2905 1836 2909
rect 1872 2907 1874 2938
rect 1894 2936 1895 2940
rect 1899 2936 1900 2940
rect 1894 2935 1900 2936
rect 2134 2940 2140 2941
rect 2134 2936 2135 2940
rect 2139 2936 2140 2940
rect 2134 2935 2140 2936
rect 2382 2940 2388 2941
rect 2382 2936 2383 2940
rect 2387 2936 2388 2940
rect 2382 2935 2388 2936
rect 2598 2940 2604 2941
rect 2598 2936 2599 2940
rect 2603 2936 2604 2940
rect 2598 2935 2604 2936
rect 2790 2940 2796 2941
rect 2790 2936 2791 2940
rect 2795 2936 2796 2940
rect 2790 2935 2796 2936
rect 2958 2940 2964 2941
rect 2958 2936 2959 2940
rect 2963 2936 2964 2940
rect 2958 2935 2964 2936
rect 3110 2940 3116 2941
rect 3110 2936 3111 2940
rect 3115 2936 3116 2940
rect 3110 2935 3116 2936
rect 3254 2940 3260 2941
rect 3254 2936 3255 2940
rect 3259 2936 3260 2940
rect 3254 2935 3260 2936
rect 3390 2940 3396 2941
rect 3390 2936 3391 2940
rect 3395 2936 3396 2940
rect 3390 2935 3396 2936
rect 3502 2940 3508 2941
rect 3502 2936 3503 2940
rect 3507 2936 3508 2940
rect 3590 2939 3591 2943
rect 3595 2939 3596 2943
rect 3590 2938 3596 2939
rect 3502 2935 3508 2936
rect 1896 2907 1898 2935
rect 2136 2907 2138 2935
rect 2384 2907 2386 2935
rect 2600 2907 2602 2935
rect 2792 2907 2794 2935
rect 2960 2907 2962 2935
rect 3112 2907 3114 2935
rect 3256 2907 3258 2935
rect 3392 2907 3394 2935
rect 3504 2907 3506 2935
rect 3592 2907 3594 2938
rect 1830 2904 1836 2905
rect 1871 2906 1875 2907
rect 1871 2901 1875 2902
rect 1895 2906 1899 2907
rect 1895 2901 1899 2902
rect 2135 2906 2139 2907
rect 2135 2901 2139 2902
rect 2351 2906 2355 2907
rect 2351 2901 2355 2902
rect 2383 2906 2387 2907
rect 2383 2901 2387 2902
rect 2447 2906 2451 2907
rect 2447 2901 2451 2902
rect 2551 2906 2555 2907
rect 2551 2901 2555 2902
rect 2599 2906 2603 2907
rect 2599 2901 2603 2902
rect 2655 2906 2659 2907
rect 2655 2901 2659 2902
rect 2759 2906 2763 2907
rect 2759 2901 2763 2902
rect 2791 2906 2795 2907
rect 2791 2901 2795 2902
rect 2871 2906 2875 2907
rect 2871 2901 2875 2902
rect 2959 2906 2963 2907
rect 2959 2901 2963 2902
rect 2983 2906 2987 2907
rect 2983 2901 2987 2902
rect 3095 2906 3099 2907
rect 3095 2901 3099 2902
rect 3111 2906 3115 2907
rect 3111 2901 3115 2902
rect 3207 2906 3211 2907
rect 3207 2901 3211 2902
rect 3255 2906 3259 2907
rect 3255 2901 3259 2902
rect 3391 2906 3395 2907
rect 3391 2901 3395 2902
rect 3503 2906 3507 2907
rect 3503 2901 3507 2902
rect 3591 2906 3595 2907
rect 3591 2901 3595 2902
rect 110 2892 116 2893
rect 110 2888 111 2892
rect 115 2888 116 2892
rect 110 2887 116 2888
rect 1830 2892 1836 2893
rect 1830 2888 1831 2892
rect 1835 2888 1836 2892
rect 1830 2887 1836 2888
rect 112 2859 114 2887
rect 254 2874 260 2875
rect 254 2870 255 2874
rect 259 2870 260 2874
rect 254 2869 260 2870
rect 358 2874 364 2875
rect 358 2870 359 2874
rect 363 2870 364 2874
rect 358 2869 364 2870
rect 478 2874 484 2875
rect 478 2870 479 2874
rect 483 2870 484 2874
rect 478 2869 484 2870
rect 614 2874 620 2875
rect 614 2870 615 2874
rect 619 2870 620 2874
rect 614 2869 620 2870
rect 758 2874 764 2875
rect 758 2870 759 2874
rect 763 2870 764 2874
rect 758 2869 764 2870
rect 902 2874 908 2875
rect 902 2870 903 2874
rect 907 2870 908 2874
rect 902 2869 908 2870
rect 1038 2874 1044 2875
rect 1038 2870 1039 2874
rect 1043 2870 1044 2874
rect 1038 2869 1044 2870
rect 1166 2874 1172 2875
rect 1166 2870 1167 2874
rect 1171 2870 1172 2874
rect 1166 2869 1172 2870
rect 1286 2874 1292 2875
rect 1286 2870 1287 2874
rect 1291 2870 1292 2874
rect 1286 2869 1292 2870
rect 1406 2874 1412 2875
rect 1406 2870 1407 2874
rect 1411 2870 1412 2874
rect 1406 2869 1412 2870
rect 1526 2874 1532 2875
rect 1526 2870 1527 2874
rect 1531 2870 1532 2874
rect 1526 2869 1532 2870
rect 1646 2874 1652 2875
rect 1646 2870 1647 2874
rect 1651 2870 1652 2874
rect 1646 2869 1652 2870
rect 256 2859 258 2869
rect 360 2859 362 2869
rect 480 2859 482 2869
rect 616 2859 618 2869
rect 760 2859 762 2869
rect 904 2859 906 2869
rect 1040 2859 1042 2869
rect 1168 2859 1170 2869
rect 1288 2859 1290 2869
rect 1408 2859 1410 2869
rect 1528 2859 1530 2869
rect 1648 2859 1650 2869
rect 1832 2859 1834 2887
rect 1872 2882 1874 2901
rect 2352 2885 2354 2901
rect 2448 2885 2450 2901
rect 2552 2885 2554 2901
rect 2656 2885 2658 2901
rect 2760 2885 2762 2901
rect 2872 2885 2874 2901
rect 2984 2885 2986 2901
rect 3096 2885 3098 2901
rect 3208 2885 3210 2901
rect 2350 2884 2356 2885
rect 1870 2881 1876 2882
rect 1870 2877 1871 2881
rect 1875 2877 1876 2881
rect 2350 2880 2351 2884
rect 2355 2880 2356 2884
rect 2350 2879 2356 2880
rect 2446 2884 2452 2885
rect 2446 2880 2447 2884
rect 2451 2880 2452 2884
rect 2446 2879 2452 2880
rect 2550 2884 2556 2885
rect 2550 2880 2551 2884
rect 2555 2880 2556 2884
rect 2550 2879 2556 2880
rect 2654 2884 2660 2885
rect 2654 2880 2655 2884
rect 2659 2880 2660 2884
rect 2654 2879 2660 2880
rect 2758 2884 2764 2885
rect 2758 2880 2759 2884
rect 2763 2880 2764 2884
rect 2758 2879 2764 2880
rect 2870 2884 2876 2885
rect 2870 2880 2871 2884
rect 2875 2880 2876 2884
rect 2870 2879 2876 2880
rect 2982 2884 2988 2885
rect 2982 2880 2983 2884
rect 2987 2880 2988 2884
rect 2982 2879 2988 2880
rect 3094 2884 3100 2885
rect 3094 2880 3095 2884
rect 3099 2880 3100 2884
rect 3094 2879 3100 2880
rect 3206 2884 3212 2885
rect 3206 2880 3207 2884
rect 3211 2880 3212 2884
rect 3592 2882 3594 2901
rect 3206 2879 3212 2880
rect 3590 2881 3596 2882
rect 1870 2876 1876 2877
rect 3590 2877 3591 2881
rect 3595 2877 3596 2881
rect 3590 2876 3596 2877
rect 1870 2864 1876 2865
rect 1870 2860 1871 2864
rect 1875 2860 1876 2864
rect 1870 2859 1876 2860
rect 3590 2864 3596 2865
rect 3590 2860 3591 2864
rect 3595 2860 3596 2864
rect 3590 2859 3596 2860
rect 111 2858 115 2859
rect 111 2853 115 2854
rect 151 2858 155 2859
rect 151 2853 155 2854
rect 255 2858 259 2859
rect 255 2853 259 2854
rect 279 2858 283 2859
rect 279 2853 283 2854
rect 359 2858 363 2859
rect 359 2853 363 2854
rect 407 2858 411 2859
rect 407 2853 411 2854
rect 479 2858 483 2859
rect 479 2853 483 2854
rect 543 2858 547 2859
rect 543 2853 547 2854
rect 615 2858 619 2859
rect 615 2853 619 2854
rect 671 2858 675 2859
rect 671 2853 675 2854
rect 759 2858 763 2859
rect 759 2853 763 2854
rect 799 2858 803 2859
rect 799 2853 803 2854
rect 903 2858 907 2859
rect 903 2853 907 2854
rect 919 2858 923 2859
rect 919 2853 923 2854
rect 1039 2858 1043 2859
rect 1039 2853 1043 2854
rect 1151 2858 1155 2859
rect 1151 2853 1155 2854
rect 1167 2858 1171 2859
rect 1167 2853 1171 2854
rect 1271 2858 1275 2859
rect 1271 2853 1275 2854
rect 1287 2858 1291 2859
rect 1287 2853 1291 2854
rect 1391 2858 1395 2859
rect 1391 2853 1395 2854
rect 1407 2858 1411 2859
rect 1407 2853 1411 2854
rect 1527 2858 1531 2859
rect 1527 2853 1531 2854
rect 1647 2858 1651 2859
rect 1647 2853 1651 2854
rect 1831 2858 1835 2859
rect 1831 2853 1835 2854
rect 112 2825 114 2853
rect 152 2843 154 2853
rect 280 2843 282 2853
rect 408 2843 410 2853
rect 544 2843 546 2853
rect 672 2843 674 2853
rect 800 2843 802 2853
rect 920 2843 922 2853
rect 1040 2843 1042 2853
rect 1152 2843 1154 2853
rect 1272 2843 1274 2853
rect 1392 2843 1394 2853
rect 150 2842 156 2843
rect 150 2838 151 2842
rect 155 2838 156 2842
rect 150 2837 156 2838
rect 278 2842 284 2843
rect 278 2838 279 2842
rect 283 2838 284 2842
rect 278 2837 284 2838
rect 406 2842 412 2843
rect 406 2838 407 2842
rect 411 2838 412 2842
rect 406 2837 412 2838
rect 542 2842 548 2843
rect 542 2838 543 2842
rect 547 2838 548 2842
rect 542 2837 548 2838
rect 670 2842 676 2843
rect 670 2838 671 2842
rect 675 2838 676 2842
rect 670 2837 676 2838
rect 798 2842 804 2843
rect 798 2838 799 2842
rect 803 2838 804 2842
rect 798 2837 804 2838
rect 918 2842 924 2843
rect 918 2838 919 2842
rect 923 2838 924 2842
rect 918 2837 924 2838
rect 1038 2842 1044 2843
rect 1038 2838 1039 2842
rect 1043 2838 1044 2842
rect 1038 2837 1044 2838
rect 1150 2842 1156 2843
rect 1150 2838 1151 2842
rect 1155 2838 1156 2842
rect 1150 2837 1156 2838
rect 1270 2842 1276 2843
rect 1270 2838 1271 2842
rect 1275 2838 1276 2842
rect 1270 2837 1276 2838
rect 1390 2842 1396 2843
rect 1390 2838 1391 2842
rect 1395 2838 1396 2842
rect 1390 2837 1396 2838
rect 1832 2825 1834 2853
rect 1872 2831 1874 2859
rect 2358 2846 2364 2847
rect 2358 2842 2359 2846
rect 2363 2842 2364 2846
rect 2358 2841 2364 2842
rect 2454 2846 2460 2847
rect 2454 2842 2455 2846
rect 2459 2842 2460 2846
rect 2454 2841 2460 2842
rect 2558 2846 2564 2847
rect 2558 2842 2559 2846
rect 2563 2842 2564 2846
rect 2558 2841 2564 2842
rect 2662 2846 2668 2847
rect 2662 2842 2663 2846
rect 2667 2842 2668 2846
rect 2662 2841 2668 2842
rect 2766 2846 2772 2847
rect 2766 2842 2767 2846
rect 2771 2842 2772 2846
rect 2766 2841 2772 2842
rect 2878 2846 2884 2847
rect 2878 2842 2879 2846
rect 2883 2842 2884 2846
rect 2878 2841 2884 2842
rect 2990 2846 2996 2847
rect 2990 2842 2991 2846
rect 2995 2842 2996 2846
rect 2990 2841 2996 2842
rect 3102 2846 3108 2847
rect 3102 2842 3103 2846
rect 3107 2842 3108 2846
rect 3102 2841 3108 2842
rect 3214 2846 3220 2847
rect 3214 2842 3215 2846
rect 3219 2842 3220 2846
rect 3214 2841 3220 2842
rect 2360 2831 2362 2841
rect 2456 2831 2458 2841
rect 2560 2831 2562 2841
rect 2664 2831 2666 2841
rect 2768 2831 2770 2841
rect 2880 2831 2882 2841
rect 2992 2831 2994 2841
rect 3104 2831 3106 2841
rect 3216 2831 3218 2841
rect 3592 2831 3594 2859
rect 1871 2830 1875 2831
rect 1871 2825 1875 2826
rect 2239 2830 2243 2831
rect 2239 2825 2243 2826
rect 2319 2830 2323 2831
rect 2319 2825 2323 2826
rect 2359 2830 2363 2831
rect 2359 2825 2363 2826
rect 2399 2830 2403 2831
rect 2399 2825 2403 2826
rect 2455 2830 2459 2831
rect 2455 2825 2459 2826
rect 2479 2830 2483 2831
rect 2479 2825 2483 2826
rect 2559 2830 2563 2831
rect 2559 2825 2563 2826
rect 2567 2830 2571 2831
rect 2567 2825 2571 2826
rect 2663 2830 2667 2831
rect 2663 2825 2667 2826
rect 2671 2830 2675 2831
rect 2671 2825 2675 2826
rect 2767 2830 2771 2831
rect 2767 2825 2771 2826
rect 2807 2830 2811 2831
rect 2807 2825 2811 2826
rect 2879 2830 2883 2831
rect 2879 2825 2883 2826
rect 2967 2830 2971 2831
rect 2967 2825 2971 2826
rect 2991 2830 2995 2831
rect 2991 2825 2995 2826
rect 3103 2830 3107 2831
rect 3103 2825 3107 2826
rect 3143 2830 3147 2831
rect 3143 2825 3147 2826
rect 3215 2830 3219 2831
rect 3215 2825 3219 2826
rect 3335 2830 3339 2831
rect 3335 2825 3339 2826
rect 3511 2830 3515 2831
rect 3511 2825 3515 2826
rect 3591 2830 3595 2831
rect 3591 2825 3595 2826
rect 110 2824 116 2825
rect 110 2820 111 2824
rect 115 2820 116 2824
rect 110 2819 116 2820
rect 1830 2824 1836 2825
rect 1830 2820 1831 2824
rect 1835 2820 1836 2824
rect 1830 2819 1836 2820
rect 110 2807 116 2808
rect 110 2803 111 2807
rect 115 2803 116 2807
rect 1830 2807 1836 2808
rect 110 2802 116 2803
rect 142 2804 148 2805
rect 112 2775 114 2802
rect 142 2800 143 2804
rect 147 2800 148 2804
rect 142 2799 148 2800
rect 270 2804 276 2805
rect 270 2800 271 2804
rect 275 2800 276 2804
rect 270 2799 276 2800
rect 398 2804 404 2805
rect 398 2800 399 2804
rect 403 2800 404 2804
rect 398 2799 404 2800
rect 534 2804 540 2805
rect 534 2800 535 2804
rect 539 2800 540 2804
rect 534 2799 540 2800
rect 662 2804 668 2805
rect 662 2800 663 2804
rect 667 2800 668 2804
rect 662 2799 668 2800
rect 790 2804 796 2805
rect 790 2800 791 2804
rect 795 2800 796 2804
rect 790 2799 796 2800
rect 910 2804 916 2805
rect 910 2800 911 2804
rect 915 2800 916 2804
rect 910 2799 916 2800
rect 1030 2804 1036 2805
rect 1030 2800 1031 2804
rect 1035 2800 1036 2804
rect 1030 2799 1036 2800
rect 1142 2804 1148 2805
rect 1142 2800 1143 2804
rect 1147 2800 1148 2804
rect 1142 2799 1148 2800
rect 1262 2804 1268 2805
rect 1262 2800 1263 2804
rect 1267 2800 1268 2804
rect 1262 2799 1268 2800
rect 1382 2804 1388 2805
rect 1382 2800 1383 2804
rect 1387 2800 1388 2804
rect 1830 2803 1831 2807
rect 1835 2803 1836 2807
rect 1830 2802 1836 2803
rect 1382 2799 1388 2800
rect 144 2775 146 2799
rect 272 2775 274 2799
rect 400 2775 402 2799
rect 536 2775 538 2799
rect 664 2775 666 2799
rect 792 2775 794 2799
rect 912 2775 914 2799
rect 1032 2775 1034 2799
rect 1144 2775 1146 2799
rect 1264 2775 1266 2799
rect 1384 2775 1386 2799
rect 1832 2775 1834 2802
rect 1872 2797 1874 2825
rect 2240 2815 2242 2825
rect 2320 2815 2322 2825
rect 2400 2815 2402 2825
rect 2480 2815 2482 2825
rect 2568 2815 2570 2825
rect 2672 2815 2674 2825
rect 2808 2815 2810 2825
rect 2968 2815 2970 2825
rect 3144 2815 3146 2825
rect 3336 2815 3338 2825
rect 3512 2815 3514 2825
rect 2238 2814 2244 2815
rect 2238 2810 2239 2814
rect 2243 2810 2244 2814
rect 2238 2809 2244 2810
rect 2318 2814 2324 2815
rect 2318 2810 2319 2814
rect 2323 2810 2324 2814
rect 2318 2809 2324 2810
rect 2398 2814 2404 2815
rect 2398 2810 2399 2814
rect 2403 2810 2404 2814
rect 2398 2809 2404 2810
rect 2478 2814 2484 2815
rect 2478 2810 2479 2814
rect 2483 2810 2484 2814
rect 2478 2809 2484 2810
rect 2566 2814 2572 2815
rect 2566 2810 2567 2814
rect 2571 2810 2572 2814
rect 2566 2809 2572 2810
rect 2670 2814 2676 2815
rect 2670 2810 2671 2814
rect 2675 2810 2676 2814
rect 2670 2809 2676 2810
rect 2806 2814 2812 2815
rect 2806 2810 2807 2814
rect 2811 2810 2812 2814
rect 2806 2809 2812 2810
rect 2966 2814 2972 2815
rect 2966 2810 2967 2814
rect 2971 2810 2972 2814
rect 2966 2809 2972 2810
rect 3142 2814 3148 2815
rect 3142 2810 3143 2814
rect 3147 2810 3148 2814
rect 3142 2809 3148 2810
rect 3334 2814 3340 2815
rect 3334 2810 3335 2814
rect 3339 2810 3340 2814
rect 3334 2809 3340 2810
rect 3510 2814 3516 2815
rect 3510 2810 3511 2814
rect 3515 2810 3516 2814
rect 3510 2809 3516 2810
rect 3592 2797 3594 2825
rect 1870 2796 1876 2797
rect 1870 2792 1871 2796
rect 1875 2792 1876 2796
rect 1870 2791 1876 2792
rect 3590 2796 3596 2797
rect 3590 2792 3591 2796
rect 3595 2792 3596 2796
rect 3590 2791 3596 2792
rect 1870 2779 1876 2780
rect 1870 2775 1871 2779
rect 1875 2775 1876 2779
rect 3590 2779 3596 2780
rect 111 2774 115 2775
rect 111 2769 115 2770
rect 143 2774 147 2775
rect 143 2769 147 2770
rect 271 2774 275 2775
rect 271 2769 275 2770
rect 295 2774 299 2775
rect 295 2769 299 2770
rect 399 2774 403 2775
rect 399 2769 403 2770
rect 439 2774 443 2775
rect 439 2769 443 2770
rect 535 2774 539 2775
rect 535 2769 539 2770
rect 567 2774 571 2775
rect 567 2769 571 2770
rect 663 2774 667 2775
rect 663 2769 667 2770
rect 687 2774 691 2775
rect 687 2769 691 2770
rect 791 2774 795 2775
rect 791 2769 795 2770
rect 799 2774 803 2775
rect 799 2769 803 2770
rect 903 2774 907 2775
rect 903 2769 907 2770
rect 911 2774 915 2775
rect 911 2769 915 2770
rect 1007 2774 1011 2775
rect 1007 2769 1011 2770
rect 1031 2774 1035 2775
rect 1031 2769 1035 2770
rect 1103 2774 1107 2775
rect 1103 2769 1107 2770
rect 1143 2774 1147 2775
rect 1143 2769 1147 2770
rect 1199 2774 1203 2775
rect 1199 2769 1203 2770
rect 1263 2774 1267 2775
rect 1263 2769 1267 2770
rect 1303 2774 1307 2775
rect 1303 2769 1307 2770
rect 1383 2774 1387 2775
rect 1383 2769 1387 2770
rect 1831 2774 1835 2775
rect 1870 2774 1876 2775
rect 2230 2776 2236 2777
rect 1831 2769 1835 2770
rect 112 2750 114 2769
rect 144 2753 146 2769
rect 296 2753 298 2769
rect 440 2753 442 2769
rect 568 2753 570 2769
rect 688 2753 690 2769
rect 800 2753 802 2769
rect 904 2753 906 2769
rect 1008 2753 1010 2769
rect 1104 2753 1106 2769
rect 1200 2753 1202 2769
rect 1304 2753 1306 2769
rect 142 2752 148 2753
rect 110 2749 116 2750
rect 110 2745 111 2749
rect 115 2745 116 2749
rect 142 2748 143 2752
rect 147 2748 148 2752
rect 142 2747 148 2748
rect 294 2752 300 2753
rect 294 2748 295 2752
rect 299 2748 300 2752
rect 294 2747 300 2748
rect 438 2752 444 2753
rect 438 2748 439 2752
rect 443 2748 444 2752
rect 438 2747 444 2748
rect 566 2752 572 2753
rect 566 2748 567 2752
rect 571 2748 572 2752
rect 566 2747 572 2748
rect 686 2752 692 2753
rect 686 2748 687 2752
rect 691 2748 692 2752
rect 686 2747 692 2748
rect 798 2752 804 2753
rect 798 2748 799 2752
rect 803 2748 804 2752
rect 798 2747 804 2748
rect 902 2752 908 2753
rect 902 2748 903 2752
rect 907 2748 908 2752
rect 902 2747 908 2748
rect 1006 2752 1012 2753
rect 1006 2748 1007 2752
rect 1011 2748 1012 2752
rect 1006 2747 1012 2748
rect 1102 2752 1108 2753
rect 1102 2748 1103 2752
rect 1107 2748 1108 2752
rect 1102 2747 1108 2748
rect 1198 2752 1204 2753
rect 1198 2748 1199 2752
rect 1203 2748 1204 2752
rect 1198 2747 1204 2748
rect 1302 2752 1308 2753
rect 1302 2748 1303 2752
rect 1307 2748 1308 2752
rect 1832 2750 1834 2769
rect 1302 2747 1308 2748
rect 1830 2749 1836 2750
rect 110 2744 116 2745
rect 1830 2745 1831 2749
rect 1835 2745 1836 2749
rect 1830 2744 1836 2745
rect 1872 2743 1874 2774
rect 2230 2772 2231 2776
rect 2235 2772 2236 2776
rect 2230 2771 2236 2772
rect 2310 2776 2316 2777
rect 2310 2772 2311 2776
rect 2315 2772 2316 2776
rect 2310 2771 2316 2772
rect 2390 2776 2396 2777
rect 2390 2772 2391 2776
rect 2395 2772 2396 2776
rect 2390 2771 2396 2772
rect 2470 2776 2476 2777
rect 2470 2772 2471 2776
rect 2475 2772 2476 2776
rect 2470 2771 2476 2772
rect 2558 2776 2564 2777
rect 2558 2772 2559 2776
rect 2563 2772 2564 2776
rect 2558 2771 2564 2772
rect 2662 2776 2668 2777
rect 2662 2772 2663 2776
rect 2667 2772 2668 2776
rect 2662 2771 2668 2772
rect 2798 2776 2804 2777
rect 2798 2772 2799 2776
rect 2803 2772 2804 2776
rect 2798 2771 2804 2772
rect 2958 2776 2964 2777
rect 2958 2772 2959 2776
rect 2963 2772 2964 2776
rect 2958 2771 2964 2772
rect 3134 2776 3140 2777
rect 3134 2772 3135 2776
rect 3139 2772 3140 2776
rect 3134 2771 3140 2772
rect 3326 2776 3332 2777
rect 3326 2772 3327 2776
rect 3331 2772 3332 2776
rect 3326 2771 3332 2772
rect 3502 2776 3508 2777
rect 3502 2772 3503 2776
rect 3507 2772 3508 2776
rect 3590 2775 3591 2779
rect 3595 2775 3596 2779
rect 3590 2774 3596 2775
rect 3502 2771 3508 2772
rect 2232 2743 2234 2771
rect 2312 2743 2314 2771
rect 2392 2743 2394 2771
rect 2472 2743 2474 2771
rect 2560 2743 2562 2771
rect 2664 2743 2666 2771
rect 2800 2743 2802 2771
rect 2960 2743 2962 2771
rect 3136 2743 3138 2771
rect 3328 2743 3330 2771
rect 3504 2743 3506 2771
rect 3592 2743 3594 2774
rect 1871 2742 1875 2743
rect 1871 2737 1875 2738
rect 2047 2742 2051 2743
rect 2047 2737 2051 2738
rect 2135 2742 2139 2743
rect 2135 2737 2139 2738
rect 2231 2742 2235 2743
rect 2231 2737 2235 2738
rect 2311 2742 2315 2743
rect 2311 2737 2315 2738
rect 2327 2742 2331 2743
rect 2327 2737 2331 2738
rect 2391 2742 2395 2743
rect 2391 2737 2395 2738
rect 2423 2742 2427 2743
rect 2423 2737 2427 2738
rect 2471 2742 2475 2743
rect 2471 2737 2475 2738
rect 2519 2742 2523 2743
rect 2519 2737 2523 2738
rect 2559 2742 2563 2743
rect 2559 2737 2563 2738
rect 2615 2742 2619 2743
rect 2615 2737 2619 2738
rect 2663 2742 2667 2743
rect 2663 2737 2667 2738
rect 2727 2742 2731 2743
rect 2727 2737 2731 2738
rect 2799 2742 2803 2743
rect 2799 2737 2803 2738
rect 2855 2742 2859 2743
rect 2855 2737 2859 2738
rect 2959 2742 2963 2743
rect 2959 2737 2963 2738
rect 3007 2742 3011 2743
rect 3007 2737 3011 2738
rect 3135 2742 3139 2743
rect 3135 2737 3139 2738
rect 3175 2742 3179 2743
rect 3175 2737 3179 2738
rect 3327 2742 3331 2743
rect 3327 2737 3331 2738
rect 3351 2742 3355 2743
rect 3351 2737 3355 2738
rect 3503 2742 3507 2743
rect 3503 2737 3507 2738
rect 3591 2742 3595 2743
rect 3591 2737 3595 2738
rect 110 2732 116 2733
rect 110 2728 111 2732
rect 115 2728 116 2732
rect 110 2727 116 2728
rect 1830 2732 1836 2733
rect 1830 2728 1831 2732
rect 1835 2728 1836 2732
rect 1830 2727 1836 2728
rect 112 2695 114 2727
rect 150 2714 156 2715
rect 150 2710 151 2714
rect 155 2710 156 2714
rect 150 2709 156 2710
rect 302 2714 308 2715
rect 302 2710 303 2714
rect 307 2710 308 2714
rect 302 2709 308 2710
rect 446 2714 452 2715
rect 446 2710 447 2714
rect 451 2710 452 2714
rect 446 2709 452 2710
rect 574 2714 580 2715
rect 574 2710 575 2714
rect 579 2710 580 2714
rect 574 2709 580 2710
rect 694 2714 700 2715
rect 694 2710 695 2714
rect 699 2710 700 2714
rect 694 2709 700 2710
rect 806 2714 812 2715
rect 806 2710 807 2714
rect 811 2710 812 2714
rect 806 2709 812 2710
rect 910 2714 916 2715
rect 910 2710 911 2714
rect 915 2710 916 2714
rect 910 2709 916 2710
rect 1014 2714 1020 2715
rect 1014 2710 1015 2714
rect 1019 2710 1020 2714
rect 1014 2709 1020 2710
rect 1110 2714 1116 2715
rect 1110 2710 1111 2714
rect 1115 2710 1116 2714
rect 1110 2709 1116 2710
rect 1206 2714 1212 2715
rect 1206 2710 1207 2714
rect 1211 2710 1212 2714
rect 1206 2709 1212 2710
rect 1310 2714 1316 2715
rect 1310 2710 1311 2714
rect 1315 2710 1316 2714
rect 1310 2709 1316 2710
rect 152 2695 154 2709
rect 304 2695 306 2709
rect 448 2695 450 2709
rect 576 2695 578 2709
rect 696 2695 698 2709
rect 808 2695 810 2709
rect 912 2695 914 2709
rect 1016 2695 1018 2709
rect 1112 2695 1114 2709
rect 1208 2695 1210 2709
rect 1312 2695 1314 2709
rect 1832 2695 1834 2727
rect 1872 2718 1874 2737
rect 2048 2721 2050 2737
rect 2136 2721 2138 2737
rect 2232 2721 2234 2737
rect 2328 2721 2330 2737
rect 2424 2721 2426 2737
rect 2520 2721 2522 2737
rect 2616 2721 2618 2737
rect 2728 2721 2730 2737
rect 2856 2721 2858 2737
rect 3008 2721 3010 2737
rect 3176 2721 3178 2737
rect 3352 2721 3354 2737
rect 3504 2721 3506 2737
rect 2046 2720 2052 2721
rect 1870 2717 1876 2718
rect 1870 2713 1871 2717
rect 1875 2713 1876 2717
rect 2046 2716 2047 2720
rect 2051 2716 2052 2720
rect 2046 2715 2052 2716
rect 2134 2720 2140 2721
rect 2134 2716 2135 2720
rect 2139 2716 2140 2720
rect 2134 2715 2140 2716
rect 2230 2720 2236 2721
rect 2230 2716 2231 2720
rect 2235 2716 2236 2720
rect 2230 2715 2236 2716
rect 2326 2720 2332 2721
rect 2326 2716 2327 2720
rect 2331 2716 2332 2720
rect 2326 2715 2332 2716
rect 2422 2720 2428 2721
rect 2422 2716 2423 2720
rect 2427 2716 2428 2720
rect 2422 2715 2428 2716
rect 2518 2720 2524 2721
rect 2518 2716 2519 2720
rect 2523 2716 2524 2720
rect 2518 2715 2524 2716
rect 2614 2720 2620 2721
rect 2614 2716 2615 2720
rect 2619 2716 2620 2720
rect 2614 2715 2620 2716
rect 2726 2720 2732 2721
rect 2726 2716 2727 2720
rect 2731 2716 2732 2720
rect 2726 2715 2732 2716
rect 2854 2720 2860 2721
rect 2854 2716 2855 2720
rect 2859 2716 2860 2720
rect 2854 2715 2860 2716
rect 3006 2720 3012 2721
rect 3006 2716 3007 2720
rect 3011 2716 3012 2720
rect 3006 2715 3012 2716
rect 3174 2720 3180 2721
rect 3174 2716 3175 2720
rect 3179 2716 3180 2720
rect 3174 2715 3180 2716
rect 3350 2720 3356 2721
rect 3350 2716 3351 2720
rect 3355 2716 3356 2720
rect 3350 2715 3356 2716
rect 3502 2720 3508 2721
rect 3502 2716 3503 2720
rect 3507 2716 3508 2720
rect 3592 2718 3594 2737
rect 3502 2715 3508 2716
rect 3590 2717 3596 2718
rect 1870 2712 1876 2713
rect 3590 2713 3591 2717
rect 3595 2713 3596 2717
rect 3590 2712 3596 2713
rect 1870 2700 1876 2701
rect 1870 2696 1871 2700
rect 1875 2696 1876 2700
rect 1870 2695 1876 2696
rect 3590 2700 3596 2701
rect 3590 2696 3591 2700
rect 3595 2696 3596 2700
rect 3590 2695 3596 2696
rect 111 2694 115 2695
rect 111 2689 115 2690
rect 143 2694 147 2695
rect 143 2689 147 2690
rect 151 2694 155 2695
rect 151 2689 155 2690
rect 263 2694 267 2695
rect 263 2689 267 2690
rect 303 2694 307 2695
rect 303 2689 307 2690
rect 407 2694 411 2695
rect 407 2689 411 2690
rect 447 2694 451 2695
rect 447 2689 451 2690
rect 543 2694 547 2695
rect 543 2689 547 2690
rect 575 2694 579 2695
rect 575 2689 579 2690
rect 671 2694 675 2695
rect 671 2689 675 2690
rect 695 2694 699 2695
rect 695 2689 699 2690
rect 791 2694 795 2695
rect 791 2689 795 2690
rect 807 2694 811 2695
rect 807 2689 811 2690
rect 903 2694 907 2695
rect 903 2689 907 2690
rect 911 2694 915 2695
rect 911 2689 915 2690
rect 1015 2694 1019 2695
rect 1015 2689 1019 2690
rect 1111 2694 1115 2695
rect 1111 2689 1115 2690
rect 1119 2694 1123 2695
rect 1119 2689 1123 2690
rect 1207 2694 1211 2695
rect 1207 2689 1211 2690
rect 1215 2694 1219 2695
rect 1215 2689 1219 2690
rect 1311 2694 1315 2695
rect 1311 2689 1315 2690
rect 1319 2694 1323 2695
rect 1319 2689 1323 2690
rect 1423 2694 1427 2695
rect 1423 2689 1427 2690
rect 1831 2694 1835 2695
rect 1831 2689 1835 2690
rect 112 2661 114 2689
rect 144 2679 146 2689
rect 264 2679 266 2689
rect 408 2679 410 2689
rect 544 2679 546 2689
rect 672 2679 674 2689
rect 792 2679 794 2689
rect 904 2679 906 2689
rect 1016 2679 1018 2689
rect 1120 2679 1122 2689
rect 1216 2679 1218 2689
rect 1320 2679 1322 2689
rect 1424 2679 1426 2689
rect 142 2678 148 2679
rect 142 2674 143 2678
rect 147 2674 148 2678
rect 142 2673 148 2674
rect 262 2678 268 2679
rect 262 2674 263 2678
rect 267 2674 268 2678
rect 262 2673 268 2674
rect 406 2678 412 2679
rect 406 2674 407 2678
rect 411 2674 412 2678
rect 406 2673 412 2674
rect 542 2678 548 2679
rect 542 2674 543 2678
rect 547 2674 548 2678
rect 542 2673 548 2674
rect 670 2678 676 2679
rect 670 2674 671 2678
rect 675 2674 676 2678
rect 670 2673 676 2674
rect 790 2678 796 2679
rect 790 2674 791 2678
rect 795 2674 796 2678
rect 790 2673 796 2674
rect 902 2678 908 2679
rect 902 2674 903 2678
rect 907 2674 908 2678
rect 902 2673 908 2674
rect 1014 2678 1020 2679
rect 1014 2674 1015 2678
rect 1019 2674 1020 2678
rect 1014 2673 1020 2674
rect 1118 2678 1124 2679
rect 1118 2674 1119 2678
rect 1123 2674 1124 2678
rect 1118 2673 1124 2674
rect 1214 2678 1220 2679
rect 1214 2674 1215 2678
rect 1219 2674 1220 2678
rect 1214 2673 1220 2674
rect 1318 2678 1324 2679
rect 1318 2674 1319 2678
rect 1323 2674 1324 2678
rect 1318 2673 1324 2674
rect 1422 2678 1428 2679
rect 1422 2674 1423 2678
rect 1427 2674 1428 2678
rect 1422 2673 1428 2674
rect 1832 2661 1834 2689
rect 1872 2667 1874 2695
rect 2054 2682 2060 2683
rect 2054 2678 2055 2682
rect 2059 2678 2060 2682
rect 2054 2677 2060 2678
rect 2142 2682 2148 2683
rect 2142 2678 2143 2682
rect 2147 2678 2148 2682
rect 2142 2677 2148 2678
rect 2238 2682 2244 2683
rect 2238 2678 2239 2682
rect 2243 2678 2244 2682
rect 2238 2677 2244 2678
rect 2334 2682 2340 2683
rect 2334 2678 2335 2682
rect 2339 2678 2340 2682
rect 2334 2677 2340 2678
rect 2430 2682 2436 2683
rect 2430 2678 2431 2682
rect 2435 2678 2436 2682
rect 2430 2677 2436 2678
rect 2526 2682 2532 2683
rect 2526 2678 2527 2682
rect 2531 2678 2532 2682
rect 2526 2677 2532 2678
rect 2622 2682 2628 2683
rect 2622 2678 2623 2682
rect 2627 2678 2628 2682
rect 2622 2677 2628 2678
rect 2734 2682 2740 2683
rect 2734 2678 2735 2682
rect 2739 2678 2740 2682
rect 2734 2677 2740 2678
rect 2862 2682 2868 2683
rect 2862 2678 2863 2682
rect 2867 2678 2868 2682
rect 2862 2677 2868 2678
rect 3014 2682 3020 2683
rect 3014 2678 3015 2682
rect 3019 2678 3020 2682
rect 3014 2677 3020 2678
rect 3182 2682 3188 2683
rect 3182 2678 3183 2682
rect 3187 2678 3188 2682
rect 3182 2677 3188 2678
rect 3358 2682 3364 2683
rect 3358 2678 3359 2682
rect 3363 2678 3364 2682
rect 3358 2677 3364 2678
rect 3510 2682 3516 2683
rect 3510 2678 3511 2682
rect 3515 2678 3516 2682
rect 3510 2677 3516 2678
rect 2056 2667 2058 2677
rect 2144 2667 2146 2677
rect 2240 2667 2242 2677
rect 2336 2667 2338 2677
rect 2432 2667 2434 2677
rect 2528 2667 2530 2677
rect 2624 2667 2626 2677
rect 2736 2667 2738 2677
rect 2864 2667 2866 2677
rect 3016 2667 3018 2677
rect 3184 2667 3186 2677
rect 3360 2667 3362 2677
rect 3512 2667 3514 2677
rect 3592 2667 3594 2695
rect 1871 2666 1875 2667
rect 1871 2661 1875 2662
rect 2055 2666 2059 2667
rect 2055 2661 2059 2662
rect 2071 2666 2075 2667
rect 2071 2661 2075 2662
rect 2143 2666 2147 2667
rect 2143 2661 2147 2662
rect 2239 2666 2243 2667
rect 2239 2661 2243 2662
rect 2295 2666 2299 2667
rect 2295 2661 2299 2662
rect 2335 2666 2339 2667
rect 2335 2661 2339 2662
rect 2431 2666 2435 2667
rect 2431 2661 2435 2662
rect 2527 2666 2531 2667
rect 2527 2661 2531 2662
rect 2567 2666 2571 2667
rect 2567 2661 2571 2662
rect 2623 2666 2627 2667
rect 2623 2661 2627 2662
rect 2735 2666 2739 2667
rect 2735 2661 2739 2662
rect 2863 2666 2867 2667
rect 2863 2661 2867 2662
rect 2871 2666 2875 2667
rect 2871 2661 2875 2662
rect 3015 2666 3019 2667
rect 3015 2661 3019 2662
rect 3183 2666 3187 2667
rect 3183 2661 3187 2662
rect 3199 2666 3203 2667
rect 3199 2661 3203 2662
rect 3359 2666 3363 2667
rect 3359 2661 3363 2662
rect 3511 2666 3515 2667
rect 3511 2661 3515 2662
rect 3591 2666 3595 2667
rect 3591 2661 3595 2662
rect 110 2660 116 2661
rect 110 2656 111 2660
rect 115 2656 116 2660
rect 110 2655 116 2656
rect 1830 2660 1836 2661
rect 1830 2656 1831 2660
rect 1835 2656 1836 2660
rect 1830 2655 1836 2656
rect 110 2643 116 2644
rect 110 2639 111 2643
rect 115 2639 116 2643
rect 1830 2643 1836 2644
rect 110 2638 116 2639
rect 134 2640 140 2641
rect 112 2611 114 2638
rect 134 2636 135 2640
rect 139 2636 140 2640
rect 134 2635 140 2636
rect 254 2640 260 2641
rect 254 2636 255 2640
rect 259 2636 260 2640
rect 254 2635 260 2636
rect 398 2640 404 2641
rect 398 2636 399 2640
rect 403 2636 404 2640
rect 398 2635 404 2636
rect 534 2640 540 2641
rect 534 2636 535 2640
rect 539 2636 540 2640
rect 534 2635 540 2636
rect 662 2640 668 2641
rect 662 2636 663 2640
rect 667 2636 668 2640
rect 662 2635 668 2636
rect 782 2640 788 2641
rect 782 2636 783 2640
rect 787 2636 788 2640
rect 782 2635 788 2636
rect 894 2640 900 2641
rect 894 2636 895 2640
rect 899 2636 900 2640
rect 894 2635 900 2636
rect 1006 2640 1012 2641
rect 1006 2636 1007 2640
rect 1011 2636 1012 2640
rect 1006 2635 1012 2636
rect 1110 2640 1116 2641
rect 1110 2636 1111 2640
rect 1115 2636 1116 2640
rect 1110 2635 1116 2636
rect 1206 2640 1212 2641
rect 1206 2636 1207 2640
rect 1211 2636 1212 2640
rect 1206 2635 1212 2636
rect 1310 2640 1316 2641
rect 1310 2636 1311 2640
rect 1315 2636 1316 2640
rect 1310 2635 1316 2636
rect 1414 2640 1420 2641
rect 1414 2636 1415 2640
rect 1419 2636 1420 2640
rect 1830 2639 1831 2643
rect 1835 2639 1836 2643
rect 1830 2638 1836 2639
rect 1414 2635 1420 2636
rect 136 2611 138 2635
rect 256 2611 258 2635
rect 400 2611 402 2635
rect 536 2611 538 2635
rect 664 2611 666 2635
rect 784 2611 786 2635
rect 896 2611 898 2635
rect 1008 2611 1010 2635
rect 1112 2611 1114 2635
rect 1208 2611 1210 2635
rect 1312 2611 1314 2635
rect 1416 2611 1418 2635
rect 1832 2611 1834 2638
rect 1872 2633 1874 2661
rect 2072 2651 2074 2661
rect 2296 2651 2298 2661
rect 2568 2651 2570 2661
rect 2872 2651 2874 2661
rect 3200 2651 3202 2661
rect 3512 2651 3514 2661
rect 2070 2650 2076 2651
rect 2070 2646 2071 2650
rect 2075 2646 2076 2650
rect 2070 2645 2076 2646
rect 2294 2650 2300 2651
rect 2294 2646 2295 2650
rect 2299 2646 2300 2650
rect 2294 2645 2300 2646
rect 2566 2650 2572 2651
rect 2566 2646 2567 2650
rect 2571 2646 2572 2650
rect 2566 2645 2572 2646
rect 2870 2650 2876 2651
rect 2870 2646 2871 2650
rect 2875 2646 2876 2650
rect 2870 2645 2876 2646
rect 3198 2650 3204 2651
rect 3198 2646 3199 2650
rect 3203 2646 3204 2650
rect 3198 2645 3204 2646
rect 3510 2650 3516 2651
rect 3510 2646 3511 2650
rect 3515 2646 3516 2650
rect 3510 2645 3516 2646
rect 3592 2633 3594 2661
rect 1870 2632 1876 2633
rect 1870 2628 1871 2632
rect 1875 2628 1876 2632
rect 1870 2627 1876 2628
rect 3590 2632 3596 2633
rect 3590 2628 3591 2632
rect 3595 2628 3596 2632
rect 3590 2627 3596 2628
rect 1870 2615 1876 2616
rect 1870 2611 1871 2615
rect 1875 2611 1876 2615
rect 3590 2615 3596 2616
rect 111 2610 115 2611
rect 111 2605 115 2606
rect 135 2610 139 2611
rect 135 2605 139 2606
rect 143 2610 147 2611
rect 143 2605 147 2606
rect 255 2610 259 2611
rect 255 2605 259 2606
rect 311 2610 315 2611
rect 311 2605 315 2606
rect 399 2610 403 2611
rect 399 2605 403 2606
rect 479 2610 483 2611
rect 479 2605 483 2606
rect 535 2610 539 2611
rect 535 2605 539 2606
rect 639 2610 643 2611
rect 639 2605 643 2606
rect 663 2610 667 2611
rect 663 2605 667 2606
rect 783 2610 787 2611
rect 783 2605 787 2606
rect 791 2610 795 2611
rect 791 2605 795 2606
rect 895 2610 899 2611
rect 895 2605 899 2606
rect 927 2610 931 2611
rect 927 2605 931 2606
rect 1007 2610 1011 2611
rect 1007 2605 1011 2606
rect 1055 2610 1059 2611
rect 1055 2605 1059 2606
rect 1111 2610 1115 2611
rect 1111 2605 1115 2606
rect 1175 2610 1179 2611
rect 1175 2605 1179 2606
rect 1207 2610 1211 2611
rect 1207 2605 1211 2606
rect 1295 2610 1299 2611
rect 1295 2605 1299 2606
rect 1311 2610 1315 2611
rect 1311 2605 1315 2606
rect 1407 2610 1411 2611
rect 1407 2605 1411 2606
rect 1415 2610 1419 2611
rect 1415 2605 1419 2606
rect 1527 2610 1531 2611
rect 1527 2605 1531 2606
rect 1831 2610 1835 2611
rect 1870 2610 1876 2611
rect 2062 2612 2068 2613
rect 1831 2605 1835 2606
rect 112 2586 114 2605
rect 144 2589 146 2605
rect 312 2589 314 2605
rect 480 2589 482 2605
rect 640 2589 642 2605
rect 792 2589 794 2605
rect 928 2589 930 2605
rect 1056 2589 1058 2605
rect 1176 2589 1178 2605
rect 1296 2589 1298 2605
rect 1408 2589 1410 2605
rect 1528 2589 1530 2605
rect 142 2588 148 2589
rect 110 2585 116 2586
rect 110 2581 111 2585
rect 115 2581 116 2585
rect 142 2584 143 2588
rect 147 2584 148 2588
rect 142 2583 148 2584
rect 310 2588 316 2589
rect 310 2584 311 2588
rect 315 2584 316 2588
rect 310 2583 316 2584
rect 478 2588 484 2589
rect 478 2584 479 2588
rect 483 2584 484 2588
rect 478 2583 484 2584
rect 638 2588 644 2589
rect 638 2584 639 2588
rect 643 2584 644 2588
rect 638 2583 644 2584
rect 790 2588 796 2589
rect 790 2584 791 2588
rect 795 2584 796 2588
rect 790 2583 796 2584
rect 926 2588 932 2589
rect 926 2584 927 2588
rect 931 2584 932 2588
rect 926 2583 932 2584
rect 1054 2588 1060 2589
rect 1054 2584 1055 2588
rect 1059 2584 1060 2588
rect 1054 2583 1060 2584
rect 1174 2588 1180 2589
rect 1174 2584 1175 2588
rect 1179 2584 1180 2588
rect 1174 2583 1180 2584
rect 1294 2588 1300 2589
rect 1294 2584 1295 2588
rect 1299 2584 1300 2588
rect 1294 2583 1300 2584
rect 1406 2588 1412 2589
rect 1406 2584 1407 2588
rect 1411 2584 1412 2588
rect 1406 2583 1412 2584
rect 1526 2588 1532 2589
rect 1526 2584 1527 2588
rect 1531 2584 1532 2588
rect 1832 2586 1834 2605
rect 1872 2587 1874 2610
rect 2062 2608 2063 2612
rect 2067 2608 2068 2612
rect 2062 2607 2068 2608
rect 2286 2612 2292 2613
rect 2286 2608 2287 2612
rect 2291 2608 2292 2612
rect 2286 2607 2292 2608
rect 2558 2612 2564 2613
rect 2558 2608 2559 2612
rect 2563 2608 2564 2612
rect 2558 2607 2564 2608
rect 2862 2612 2868 2613
rect 2862 2608 2863 2612
rect 2867 2608 2868 2612
rect 2862 2607 2868 2608
rect 3190 2612 3196 2613
rect 3190 2608 3191 2612
rect 3195 2608 3196 2612
rect 3190 2607 3196 2608
rect 3502 2612 3508 2613
rect 3502 2608 3503 2612
rect 3507 2608 3508 2612
rect 3590 2611 3591 2615
rect 3595 2611 3596 2615
rect 3590 2610 3596 2611
rect 3502 2607 3508 2608
rect 2064 2587 2066 2607
rect 2288 2587 2290 2607
rect 2560 2587 2562 2607
rect 2864 2587 2866 2607
rect 3192 2587 3194 2607
rect 3504 2587 3506 2607
rect 3592 2587 3594 2610
rect 1871 2586 1875 2587
rect 1526 2583 1532 2584
rect 1830 2585 1836 2586
rect 110 2580 116 2581
rect 1830 2581 1831 2585
rect 1835 2581 1836 2585
rect 1871 2581 1875 2582
rect 2063 2586 2067 2587
rect 2063 2581 2067 2582
rect 2167 2586 2171 2587
rect 2167 2581 2171 2582
rect 2263 2586 2267 2587
rect 2263 2581 2267 2582
rect 2287 2586 2291 2587
rect 2287 2581 2291 2582
rect 2367 2586 2371 2587
rect 2367 2581 2371 2582
rect 2479 2586 2483 2587
rect 2479 2581 2483 2582
rect 2559 2586 2563 2587
rect 2559 2581 2563 2582
rect 2591 2586 2595 2587
rect 2591 2581 2595 2582
rect 2695 2586 2699 2587
rect 2695 2581 2699 2582
rect 2799 2586 2803 2587
rect 2799 2581 2803 2582
rect 2863 2586 2867 2587
rect 2863 2581 2867 2582
rect 2903 2586 2907 2587
rect 2903 2581 2907 2582
rect 3015 2586 3019 2587
rect 3015 2581 3019 2582
rect 3135 2586 3139 2587
rect 3135 2581 3139 2582
rect 3191 2586 3195 2587
rect 3191 2581 3195 2582
rect 3263 2586 3267 2587
rect 3263 2581 3267 2582
rect 3391 2586 3395 2587
rect 3391 2581 3395 2582
rect 3503 2586 3507 2587
rect 3503 2581 3507 2582
rect 3591 2586 3595 2587
rect 3591 2581 3595 2582
rect 1830 2580 1836 2581
rect 110 2568 116 2569
rect 110 2564 111 2568
rect 115 2564 116 2568
rect 110 2563 116 2564
rect 1830 2568 1836 2569
rect 1830 2564 1831 2568
rect 1835 2564 1836 2568
rect 1830 2563 1836 2564
rect 112 2527 114 2563
rect 150 2550 156 2551
rect 150 2546 151 2550
rect 155 2546 156 2550
rect 150 2545 156 2546
rect 318 2550 324 2551
rect 318 2546 319 2550
rect 323 2546 324 2550
rect 318 2545 324 2546
rect 486 2550 492 2551
rect 486 2546 487 2550
rect 491 2546 492 2550
rect 486 2545 492 2546
rect 646 2550 652 2551
rect 646 2546 647 2550
rect 651 2546 652 2550
rect 646 2545 652 2546
rect 798 2550 804 2551
rect 798 2546 799 2550
rect 803 2546 804 2550
rect 798 2545 804 2546
rect 934 2550 940 2551
rect 934 2546 935 2550
rect 939 2546 940 2550
rect 934 2545 940 2546
rect 1062 2550 1068 2551
rect 1062 2546 1063 2550
rect 1067 2546 1068 2550
rect 1062 2545 1068 2546
rect 1182 2550 1188 2551
rect 1182 2546 1183 2550
rect 1187 2546 1188 2550
rect 1182 2545 1188 2546
rect 1302 2550 1308 2551
rect 1302 2546 1303 2550
rect 1307 2546 1308 2550
rect 1302 2545 1308 2546
rect 1414 2550 1420 2551
rect 1414 2546 1415 2550
rect 1419 2546 1420 2550
rect 1414 2545 1420 2546
rect 1534 2550 1540 2551
rect 1534 2546 1535 2550
rect 1539 2546 1540 2550
rect 1534 2545 1540 2546
rect 152 2527 154 2545
rect 320 2527 322 2545
rect 488 2527 490 2545
rect 648 2527 650 2545
rect 800 2527 802 2545
rect 936 2527 938 2545
rect 1064 2527 1066 2545
rect 1184 2527 1186 2545
rect 1304 2527 1306 2545
rect 1416 2527 1418 2545
rect 1536 2527 1538 2545
rect 1832 2527 1834 2563
rect 1872 2562 1874 2581
rect 2168 2565 2170 2581
rect 2264 2565 2266 2581
rect 2368 2565 2370 2581
rect 2480 2565 2482 2581
rect 2592 2565 2594 2581
rect 2696 2565 2698 2581
rect 2800 2565 2802 2581
rect 2904 2565 2906 2581
rect 3016 2565 3018 2581
rect 3136 2565 3138 2581
rect 3264 2565 3266 2581
rect 3392 2565 3394 2581
rect 3504 2565 3506 2581
rect 2166 2564 2172 2565
rect 1870 2561 1876 2562
rect 1870 2557 1871 2561
rect 1875 2557 1876 2561
rect 2166 2560 2167 2564
rect 2171 2560 2172 2564
rect 2166 2559 2172 2560
rect 2262 2564 2268 2565
rect 2262 2560 2263 2564
rect 2267 2560 2268 2564
rect 2262 2559 2268 2560
rect 2366 2564 2372 2565
rect 2366 2560 2367 2564
rect 2371 2560 2372 2564
rect 2366 2559 2372 2560
rect 2478 2564 2484 2565
rect 2478 2560 2479 2564
rect 2483 2560 2484 2564
rect 2478 2559 2484 2560
rect 2590 2564 2596 2565
rect 2590 2560 2591 2564
rect 2595 2560 2596 2564
rect 2590 2559 2596 2560
rect 2694 2564 2700 2565
rect 2694 2560 2695 2564
rect 2699 2560 2700 2564
rect 2694 2559 2700 2560
rect 2798 2564 2804 2565
rect 2798 2560 2799 2564
rect 2803 2560 2804 2564
rect 2798 2559 2804 2560
rect 2902 2564 2908 2565
rect 2902 2560 2903 2564
rect 2907 2560 2908 2564
rect 2902 2559 2908 2560
rect 3014 2564 3020 2565
rect 3014 2560 3015 2564
rect 3019 2560 3020 2564
rect 3014 2559 3020 2560
rect 3134 2564 3140 2565
rect 3134 2560 3135 2564
rect 3139 2560 3140 2564
rect 3134 2559 3140 2560
rect 3262 2564 3268 2565
rect 3262 2560 3263 2564
rect 3267 2560 3268 2564
rect 3262 2559 3268 2560
rect 3390 2564 3396 2565
rect 3390 2560 3391 2564
rect 3395 2560 3396 2564
rect 3390 2559 3396 2560
rect 3502 2564 3508 2565
rect 3502 2560 3503 2564
rect 3507 2560 3508 2564
rect 3592 2562 3594 2581
rect 3502 2559 3508 2560
rect 3590 2561 3596 2562
rect 1870 2556 1876 2557
rect 3590 2557 3591 2561
rect 3595 2557 3596 2561
rect 3590 2556 3596 2557
rect 1870 2544 1876 2545
rect 1870 2540 1871 2544
rect 1875 2540 1876 2544
rect 1870 2539 1876 2540
rect 3590 2544 3596 2545
rect 3590 2540 3591 2544
rect 3595 2540 3596 2544
rect 3590 2539 3596 2540
rect 111 2526 115 2527
rect 111 2521 115 2522
rect 143 2526 147 2527
rect 143 2521 147 2522
rect 151 2526 155 2527
rect 151 2521 155 2522
rect 295 2526 299 2527
rect 295 2521 299 2522
rect 319 2526 323 2527
rect 319 2521 323 2522
rect 447 2526 451 2527
rect 447 2521 451 2522
rect 487 2526 491 2527
rect 487 2521 491 2522
rect 591 2526 595 2527
rect 591 2521 595 2522
rect 647 2526 651 2527
rect 647 2521 651 2522
rect 735 2526 739 2527
rect 735 2521 739 2522
rect 799 2526 803 2527
rect 799 2521 803 2522
rect 879 2526 883 2527
rect 879 2521 883 2522
rect 935 2526 939 2527
rect 935 2521 939 2522
rect 1015 2526 1019 2527
rect 1015 2521 1019 2522
rect 1063 2526 1067 2527
rect 1063 2521 1067 2522
rect 1143 2526 1147 2527
rect 1143 2521 1147 2522
rect 1183 2526 1187 2527
rect 1183 2521 1187 2522
rect 1271 2526 1275 2527
rect 1271 2521 1275 2522
rect 1303 2526 1307 2527
rect 1303 2521 1307 2522
rect 1399 2526 1403 2527
rect 1399 2521 1403 2522
rect 1415 2526 1419 2527
rect 1415 2521 1419 2522
rect 1535 2526 1539 2527
rect 1535 2521 1539 2522
rect 1831 2526 1835 2527
rect 1831 2521 1835 2522
rect 112 2493 114 2521
rect 144 2511 146 2521
rect 296 2511 298 2521
rect 448 2511 450 2521
rect 592 2511 594 2521
rect 736 2511 738 2521
rect 880 2511 882 2521
rect 1016 2511 1018 2521
rect 1144 2511 1146 2521
rect 1272 2511 1274 2521
rect 1400 2511 1402 2521
rect 1536 2511 1538 2521
rect 142 2510 148 2511
rect 142 2506 143 2510
rect 147 2506 148 2510
rect 142 2505 148 2506
rect 294 2510 300 2511
rect 294 2506 295 2510
rect 299 2506 300 2510
rect 294 2505 300 2506
rect 446 2510 452 2511
rect 446 2506 447 2510
rect 451 2506 452 2510
rect 446 2505 452 2506
rect 590 2510 596 2511
rect 590 2506 591 2510
rect 595 2506 596 2510
rect 590 2505 596 2506
rect 734 2510 740 2511
rect 734 2506 735 2510
rect 739 2506 740 2510
rect 734 2505 740 2506
rect 878 2510 884 2511
rect 878 2506 879 2510
rect 883 2506 884 2510
rect 878 2505 884 2506
rect 1014 2510 1020 2511
rect 1014 2506 1015 2510
rect 1019 2506 1020 2510
rect 1014 2505 1020 2506
rect 1142 2510 1148 2511
rect 1142 2506 1143 2510
rect 1147 2506 1148 2510
rect 1142 2505 1148 2506
rect 1270 2510 1276 2511
rect 1270 2506 1271 2510
rect 1275 2506 1276 2510
rect 1270 2505 1276 2506
rect 1398 2510 1404 2511
rect 1398 2506 1399 2510
rect 1403 2506 1404 2510
rect 1398 2505 1404 2506
rect 1534 2510 1540 2511
rect 1534 2506 1535 2510
rect 1539 2506 1540 2510
rect 1534 2505 1540 2506
rect 1832 2493 1834 2521
rect 1872 2511 1874 2539
rect 2174 2526 2180 2527
rect 2174 2522 2175 2526
rect 2179 2522 2180 2526
rect 2174 2521 2180 2522
rect 2270 2526 2276 2527
rect 2270 2522 2271 2526
rect 2275 2522 2276 2526
rect 2270 2521 2276 2522
rect 2374 2526 2380 2527
rect 2374 2522 2375 2526
rect 2379 2522 2380 2526
rect 2374 2521 2380 2522
rect 2486 2526 2492 2527
rect 2486 2522 2487 2526
rect 2491 2522 2492 2526
rect 2486 2521 2492 2522
rect 2598 2526 2604 2527
rect 2598 2522 2599 2526
rect 2603 2522 2604 2526
rect 2598 2521 2604 2522
rect 2702 2526 2708 2527
rect 2702 2522 2703 2526
rect 2707 2522 2708 2526
rect 2702 2521 2708 2522
rect 2806 2526 2812 2527
rect 2806 2522 2807 2526
rect 2811 2522 2812 2526
rect 2806 2521 2812 2522
rect 2910 2526 2916 2527
rect 2910 2522 2911 2526
rect 2915 2522 2916 2526
rect 2910 2521 2916 2522
rect 3022 2526 3028 2527
rect 3022 2522 3023 2526
rect 3027 2522 3028 2526
rect 3022 2521 3028 2522
rect 3142 2526 3148 2527
rect 3142 2522 3143 2526
rect 3147 2522 3148 2526
rect 3142 2521 3148 2522
rect 3270 2526 3276 2527
rect 3270 2522 3271 2526
rect 3275 2522 3276 2526
rect 3270 2521 3276 2522
rect 3398 2526 3404 2527
rect 3398 2522 3399 2526
rect 3403 2522 3404 2526
rect 3398 2521 3404 2522
rect 3510 2526 3516 2527
rect 3510 2522 3511 2526
rect 3515 2522 3516 2526
rect 3510 2521 3516 2522
rect 2176 2511 2178 2521
rect 2272 2511 2274 2521
rect 2376 2511 2378 2521
rect 2488 2511 2490 2521
rect 2600 2511 2602 2521
rect 2704 2511 2706 2521
rect 2808 2511 2810 2521
rect 2912 2511 2914 2521
rect 3024 2511 3026 2521
rect 3144 2511 3146 2521
rect 3272 2511 3274 2521
rect 3400 2511 3402 2521
rect 3512 2511 3514 2521
rect 3592 2511 3594 2539
rect 1871 2510 1875 2511
rect 1871 2505 1875 2506
rect 2135 2510 2139 2511
rect 2135 2505 2139 2506
rect 2175 2510 2179 2511
rect 2175 2505 2179 2506
rect 2223 2510 2227 2511
rect 2223 2505 2227 2506
rect 2271 2510 2275 2511
rect 2271 2505 2275 2506
rect 2319 2510 2323 2511
rect 2319 2505 2323 2506
rect 2375 2510 2379 2511
rect 2375 2505 2379 2506
rect 2423 2510 2427 2511
rect 2423 2505 2427 2506
rect 2487 2510 2491 2511
rect 2487 2505 2491 2506
rect 2535 2510 2539 2511
rect 2535 2505 2539 2506
rect 2599 2510 2603 2511
rect 2599 2505 2603 2506
rect 2655 2510 2659 2511
rect 2655 2505 2659 2506
rect 2703 2510 2707 2511
rect 2703 2505 2707 2506
rect 2783 2510 2787 2511
rect 2783 2505 2787 2506
rect 2807 2510 2811 2511
rect 2807 2505 2811 2506
rect 2911 2510 2915 2511
rect 2911 2505 2915 2506
rect 2919 2510 2923 2511
rect 2919 2505 2923 2506
rect 3023 2510 3027 2511
rect 3023 2505 3027 2506
rect 3063 2510 3067 2511
rect 3063 2505 3067 2506
rect 3143 2510 3147 2511
rect 3143 2505 3147 2506
rect 3215 2510 3219 2511
rect 3215 2505 3219 2506
rect 3271 2510 3275 2511
rect 3271 2505 3275 2506
rect 3375 2510 3379 2511
rect 3375 2505 3379 2506
rect 3399 2510 3403 2511
rect 3399 2505 3403 2506
rect 3511 2510 3515 2511
rect 3511 2505 3515 2506
rect 3591 2510 3595 2511
rect 3591 2505 3595 2506
rect 110 2492 116 2493
rect 110 2488 111 2492
rect 115 2488 116 2492
rect 110 2487 116 2488
rect 1830 2492 1836 2493
rect 1830 2488 1831 2492
rect 1835 2488 1836 2492
rect 1830 2487 1836 2488
rect 1872 2477 1874 2505
rect 2136 2495 2138 2505
rect 2224 2495 2226 2505
rect 2320 2495 2322 2505
rect 2424 2495 2426 2505
rect 2536 2495 2538 2505
rect 2656 2495 2658 2505
rect 2784 2495 2786 2505
rect 2920 2495 2922 2505
rect 3064 2495 3066 2505
rect 3216 2495 3218 2505
rect 3376 2495 3378 2505
rect 3512 2495 3514 2505
rect 2134 2494 2140 2495
rect 2134 2490 2135 2494
rect 2139 2490 2140 2494
rect 2134 2489 2140 2490
rect 2222 2494 2228 2495
rect 2222 2490 2223 2494
rect 2227 2490 2228 2494
rect 2222 2489 2228 2490
rect 2318 2494 2324 2495
rect 2318 2490 2319 2494
rect 2323 2490 2324 2494
rect 2318 2489 2324 2490
rect 2422 2494 2428 2495
rect 2422 2490 2423 2494
rect 2427 2490 2428 2494
rect 2422 2489 2428 2490
rect 2534 2494 2540 2495
rect 2534 2490 2535 2494
rect 2539 2490 2540 2494
rect 2534 2489 2540 2490
rect 2654 2494 2660 2495
rect 2654 2490 2655 2494
rect 2659 2490 2660 2494
rect 2654 2489 2660 2490
rect 2782 2494 2788 2495
rect 2782 2490 2783 2494
rect 2787 2490 2788 2494
rect 2782 2489 2788 2490
rect 2918 2494 2924 2495
rect 2918 2490 2919 2494
rect 2923 2490 2924 2494
rect 2918 2489 2924 2490
rect 3062 2494 3068 2495
rect 3062 2490 3063 2494
rect 3067 2490 3068 2494
rect 3062 2489 3068 2490
rect 3214 2494 3220 2495
rect 3214 2490 3215 2494
rect 3219 2490 3220 2494
rect 3214 2489 3220 2490
rect 3374 2494 3380 2495
rect 3374 2490 3375 2494
rect 3379 2490 3380 2494
rect 3374 2489 3380 2490
rect 3510 2494 3516 2495
rect 3510 2490 3511 2494
rect 3515 2490 3516 2494
rect 3510 2489 3516 2490
rect 3592 2477 3594 2505
rect 1870 2476 1876 2477
rect 110 2475 116 2476
rect 110 2471 111 2475
rect 115 2471 116 2475
rect 1830 2475 1836 2476
rect 110 2470 116 2471
rect 134 2472 140 2473
rect 112 2447 114 2470
rect 134 2468 135 2472
rect 139 2468 140 2472
rect 134 2467 140 2468
rect 286 2472 292 2473
rect 286 2468 287 2472
rect 291 2468 292 2472
rect 286 2467 292 2468
rect 438 2472 444 2473
rect 438 2468 439 2472
rect 443 2468 444 2472
rect 438 2467 444 2468
rect 582 2472 588 2473
rect 582 2468 583 2472
rect 587 2468 588 2472
rect 582 2467 588 2468
rect 726 2472 732 2473
rect 726 2468 727 2472
rect 731 2468 732 2472
rect 726 2467 732 2468
rect 870 2472 876 2473
rect 870 2468 871 2472
rect 875 2468 876 2472
rect 870 2467 876 2468
rect 1006 2472 1012 2473
rect 1006 2468 1007 2472
rect 1011 2468 1012 2472
rect 1006 2467 1012 2468
rect 1134 2472 1140 2473
rect 1134 2468 1135 2472
rect 1139 2468 1140 2472
rect 1134 2467 1140 2468
rect 1262 2472 1268 2473
rect 1262 2468 1263 2472
rect 1267 2468 1268 2472
rect 1262 2467 1268 2468
rect 1390 2472 1396 2473
rect 1390 2468 1391 2472
rect 1395 2468 1396 2472
rect 1390 2467 1396 2468
rect 1526 2472 1532 2473
rect 1526 2468 1527 2472
rect 1531 2468 1532 2472
rect 1830 2471 1831 2475
rect 1835 2471 1836 2475
rect 1870 2472 1871 2476
rect 1875 2472 1876 2476
rect 1870 2471 1876 2472
rect 3590 2476 3596 2477
rect 3590 2472 3591 2476
rect 3595 2472 3596 2476
rect 3590 2471 3596 2472
rect 1830 2470 1836 2471
rect 1526 2467 1532 2468
rect 136 2447 138 2467
rect 288 2447 290 2467
rect 440 2447 442 2467
rect 584 2447 586 2467
rect 728 2447 730 2467
rect 872 2447 874 2467
rect 1008 2447 1010 2467
rect 1136 2447 1138 2467
rect 1264 2447 1266 2467
rect 1392 2447 1394 2467
rect 1528 2447 1530 2467
rect 1832 2447 1834 2470
rect 1870 2459 1876 2460
rect 1870 2455 1871 2459
rect 1875 2455 1876 2459
rect 3590 2459 3596 2460
rect 1870 2454 1876 2455
rect 2126 2456 2132 2457
rect 111 2446 115 2447
rect 111 2441 115 2442
rect 135 2446 139 2447
rect 135 2441 139 2442
rect 199 2446 203 2447
rect 199 2441 203 2442
rect 287 2446 291 2447
rect 287 2441 291 2442
rect 351 2446 355 2447
rect 351 2441 355 2442
rect 439 2446 443 2447
rect 439 2441 443 2442
rect 495 2446 499 2447
rect 495 2441 499 2442
rect 583 2446 587 2447
rect 583 2441 587 2442
rect 639 2446 643 2447
rect 639 2441 643 2442
rect 727 2446 731 2447
rect 727 2441 731 2442
rect 783 2446 787 2447
rect 783 2441 787 2442
rect 871 2446 875 2447
rect 871 2441 875 2442
rect 919 2446 923 2447
rect 919 2441 923 2442
rect 1007 2446 1011 2447
rect 1007 2441 1011 2442
rect 1047 2446 1051 2447
rect 1047 2441 1051 2442
rect 1135 2446 1139 2447
rect 1135 2441 1139 2442
rect 1175 2446 1179 2447
rect 1175 2441 1179 2442
rect 1263 2446 1267 2447
rect 1263 2441 1267 2442
rect 1311 2446 1315 2447
rect 1311 2441 1315 2442
rect 1391 2446 1395 2447
rect 1391 2441 1395 2442
rect 1447 2446 1451 2447
rect 1447 2441 1451 2442
rect 1527 2446 1531 2447
rect 1527 2441 1531 2442
rect 1831 2446 1835 2447
rect 1831 2441 1835 2442
rect 112 2422 114 2441
rect 200 2425 202 2441
rect 352 2425 354 2441
rect 496 2425 498 2441
rect 640 2425 642 2441
rect 784 2425 786 2441
rect 920 2425 922 2441
rect 1048 2425 1050 2441
rect 1176 2425 1178 2441
rect 1312 2425 1314 2441
rect 1448 2425 1450 2441
rect 198 2424 204 2425
rect 110 2421 116 2422
rect 110 2417 111 2421
rect 115 2417 116 2421
rect 198 2420 199 2424
rect 203 2420 204 2424
rect 198 2419 204 2420
rect 350 2424 356 2425
rect 350 2420 351 2424
rect 355 2420 356 2424
rect 350 2419 356 2420
rect 494 2424 500 2425
rect 494 2420 495 2424
rect 499 2420 500 2424
rect 494 2419 500 2420
rect 638 2424 644 2425
rect 638 2420 639 2424
rect 643 2420 644 2424
rect 638 2419 644 2420
rect 782 2424 788 2425
rect 782 2420 783 2424
rect 787 2420 788 2424
rect 782 2419 788 2420
rect 918 2424 924 2425
rect 918 2420 919 2424
rect 923 2420 924 2424
rect 918 2419 924 2420
rect 1046 2424 1052 2425
rect 1046 2420 1047 2424
rect 1051 2420 1052 2424
rect 1046 2419 1052 2420
rect 1174 2424 1180 2425
rect 1174 2420 1175 2424
rect 1179 2420 1180 2424
rect 1174 2419 1180 2420
rect 1310 2424 1316 2425
rect 1310 2420 1311 2424
rect 1315 2420 1316 2424
rect 1310 2419 1316 2420
rect 1446 2424 1452 2425
rect 1446 2420 1447 2424
rect 1451 2420 1452 2424
rect 1832 2422 1834 2441
rect 1872 2427 1874 2454
rect 2126 2452 2127 2456
rect 2131 2452 2132 2456
rect 2126 2451 2132 2452
rect 2214 2456 2220 2457
rect 2214 2452 2215 2456
rect 2219 2452 2220 2456
rect 2214 2451 2220 2452
rect 2310 2456 2316 2457
rect 2310 2452 2311 2456
rect 2315 2452 2316 2456
rect 2310 2451 2316 2452
rect 2414 2456 2420 2457
rect 2414 2452 2415 2456
rect 2419 2452 2420 2456
rect 2414 2451 2420 2452
rect 2526 2456 2532 2457
rect 2526 2452 2527 2456
rect 2531 2452 2532 2456
rect 2526 2451 2532 2452
rect 2646 2456 2652 2457
rect 2646 2452 2647 2456
rect 2651 2452 2652 2456
rect 2646 2451 2652 2452
rect 2774 2456 2780 2457
rect 2774 2452 2775 2456
rect 2779 2452 2780 2456
rect 2774 2451 2780 2452
rect 2910 2456 2916 2457
rect 2910 2452 2911 2456
rect 2915 2452 2916 2456
rect 2910 2451 2916 2452
rect 3054 2456 3060 2457
rect 3054 2452 3055 2456
rect 3059 2452 3060 2456
rect 3054 2451 3060 2452
rect 3206 2456 3212 2457
rect 3206 2452 3207 2456
rect 3211 2452 3212 2456
rect 3206 2451 3212 2452
rect 3366 2456 3372 2457
rect 3366 2452 3367 2456
rect 3371 2452 3372 2456
rect 3366 2451 3372 2452
rect 3502 2456 3508 2457
rect 3502 2452 3503 2456
rect 3507 2452 3508 2456
rect 3590 2455 3591 2459
rect 3595 2455 3596 2459
rect 3590 2454 3596 2455
rect 3502 2451 3508 2452
rect 2128 2427 2130 2451
rect 2216 2427 2218 2451
rect 2312 2427 2314 2451
rect 2416 2427 2418 2451
rect 2528 2427 2530 2451
rect 2648 2427 2650 2451
rect 2776 2427 2778 2451
rect 2912 2427 2914 2451
rect 3056 2427 3058 2451
rect 3208 2427 3210 2451
rect 3368 2427 3370 2451
rect 3504 2427 3506 2451
rect 3592 2427 3594 2454
rect 1871 2426 1875 2427
rect 1446 2419 1452 2420
rect 1830 2421 1836 2422
rect 1871 2421 1875 2422
rect 1975 2426 1979 2427
rect 1975 2421 1979 2422
rect 2087 2426 2091 2427
rect 2087 2421 2091 2422
rect 2127 2426 2131 2427
rect 2127 2421 2131 2422
rect 2207 2426 2211 2427
rect 2207 2421 2211 2422
rect 2215 2426 2219 2427
rect 2215 2421 2219 2422
rect 2311 2426 2315 2427
rect 2311 2421 2315 2422
rect 2335 2426 2339 2427
rect 2335 2421 2339 2422
rect 2415 2426 2419 2427
rect 2415 2421 2419 2422
rect 2479 2426 2483 2427
rect 2479 2421 2483 2422
rect 2527 2426 2531 2427
rect 2527 2421 2531 2422
rect 2631 2426 2635 2427
rect 2631 2421 2635 2422
rect 2647 2426 2651 2427
rect 2647 2421 2651 2422
rect 2775 2426 2779 2427
rect 2775 2421 2779 2422
rect 2791 2426 2795 2427
rect 2791 2421 2795 2422
rect 2911 2426 2915 2427
rect 2911 2421 2915 2422
rect 2967 2426 2971 2427
rect 2967 2421 2971 2422
rect 3055 2426 3059 2427
rect 3055 2421 3059 2422
rect 3151 2426 3155 2427
rect 3151 2421 3155 2422
rect 3207 2426 3211 2427
rect 3207 2421 3211 2422
rect 3335 2426 3339 2427
rect 3335 2421 3339 2422
rect 3367 2426 3371 2427
rect 3367 2421 3371 2422
rect 3503 2426 3507 2427
rect 3503 2421 3507 2422
rect 3591 2426 3595 2427
rect 3591 2421 3595 2422
rect 110 2416 116 2417
rect 1830 2417 1831 2421
rect 1835 2417 1836 2421
rect 1830 2416 1836 2417
rect 110 2404 116 2405
rect 110 2400 111 2404
rect 115 2400 116 2404
rect 110 2399 116 2400
rect 1830 2404 1836 2405
rect 1830 2400 1831 2404
rect 1835 2400 1836 2404
rect 1872 2402 1874 2421
rect 1976 2405 1978 2421
rect 2088 2405 2090 2421
rect 2208 2405 2210 2421
rect 2336 2405 2338 2421
rect 2480 2405 2482 2421
rect 2632 2405 2634 2421
rect 2792 2405 2794 2421
rect 2968 2405 2970 2421
rect 3152 2405 3154 2421
rect 3336 2405 3338 2421
rect 3504 2405 3506 2421
rect 1974 2404 1980 2405
rect 1830 2399 1836 2400
rect 1870 2401 1876 2402
rect 112 2363 114 2399
rect 206 2386 212 2387
rect 206 2382 207 2386
rect 211 2382 212 2386
rect 206 2381 212 2382
rect 358 2386 364 2387
rect 358 2382 359 2386
rect 363 2382 364 2386
rect 358 2381 364 2382
rect 502 2386 508 2387
rect 502 2382 503 2386
rect 507 2382 508 2386
rect 502 2381 508 2382
rect 646 2386 652 2387
rect 646 2382 647 2386
rect 651 2382 652 2386
rect 646 2381 652 2382
rect 790 2386 796 2387
rect 790 2382 791 2386
rect 795 2382 796 2386
rect 790 2381 796 2382
rect 926 2386 932 2387
rect 926 2382 927 2386
rect 931 2382 932 2386
rect 926 2381 932 2382
rect 1054 2386 1060 2387
rect 1054 2382 1055 2386
rect 1059 2382 1060 2386
rect 1054 2381 1060 2382
rect 1182 2386 1188 2387
rect 1182 2382 1183 2386
rect 1187 2382 1188 2386
rect 1182 2381 1188 2382
rect 1318 2386 1324 2387
rect 1318 2382 1319 2386
rect 1323 2382 1324 2386
rect 1318 2381 1324 2382
rect 1454 2386 1460 2387
rect 1454 2382 1455 2386
rect 1459 2382 1460 2386
rect 1454 2381 1460 2382
rect 208 2363 210 2381
rect 360 2363 362 2381
rect 504 2363 506 2381
rect 648 2363 650 2381
rect 792 2363 794 2381
rect 928 2363 930 2381
rect 1056 2363 1058 2381
rect 1184 2363 1186 2381
rect 1320 2363 1322 2381
rect 1456 2363 1458 2381
rect 1832 2363 1834 2399
rect 1870 2397 1871 2401
rect 1875 2397 1876 2401
rect 1974 2400 1975 2404
rect 1979 2400 1980 2404
rect 1974 2399 1980 2400
rect 2086 2404 2092 2405
rect 2086 2400 2087 2404
rect 2091 2400 2092 2404
rect 2086 2399 2092 2400
rect 2206 2404 2212 2405
rect 2206 2400 2207 2404
rect 2211 2400 2212 2404
rect 2206 2399 2212 2400
rect 2334 2404 2340 2405
rect 2334 2400 2335 2404
rect 2339 2400 2340 2404
rect 2334 2399 2340 2400
rect 2478 2404 2484 2405
rect 2478 2400 2479 2404
rect 2483 2400 2484 2404
rect 2478 2399 2484 2400
rect 2630 2404 2636 2405
rect 2630 2400 2631 2404
rect 2635 2400 2636 2404
rect 2630 2399 2636 2400
rect 2790 2404 2796 2405
rect 2790 2400 2791 2404
rect 2795 2400 2796 2404
rect 2790 2399 2796 2400
rect 2966 2404 2972 2405
rect 2966 2400 2967 2404
rect 2971 2400 2972 2404
rect 2966 2399 2972 2400
rect 3150 2404 3156 2405
rect 3150 2400 3151 2404
rect 3155 2400 3156 2404
rect 3150 2399 3156 2400
rect 3334 2404 3340 2405
rect 3334 2400 3335 2404
rect 3339 2400 3340 2404
rect 3334 2399 3340 2400
rect 3502 2404 3508 2405
rect 3502 2400 3503 2404
rect 3507 2400 3508 2404
rect 3592 2402 3594 2421
rect 3502 2399 3508 2400
rect 3590 2401 3596 2402
rect 1870 2396 1876 2397
rect 3590 2397 3591 2401
rect 3595 2397 3596 2401
rect 3590 2396 3596 2397
rect 1870 2384 1876 2385
rect 1870 2380 1871 2384
rect 1875 2380 1876 2384
rect 1870 2379 1876 2380
rect 3590 2384 3596 2385
rect 3590 2380 3591 2384
rect 3595 2380 3596 2384
rect 3590 2379 3596 2380
rect 111 2362 115 2363
rect 111 2357 115 2358
rect 207 2362 211 2363
rect 207 2357 211 2358
rect 223 2362 227 2363
rect 223 2357 227 2358
rect 327 2362 331 2363
rect 327 2357 331 2358
rect 359 2362 363 2363
rect 359 2357 363 2358
rect 439 2362 443 2363
rect 439 2357 443 2358
rect 503 2362 507 2363
rect 503 2357 507 2358
rect 559 2362 563 2363
rect 559 2357 563 2358
rect 647 2362 651 2363
rect 647 2357 651 2358
rect 679 2362 683 2363
rect 679 2357 683 2358
rect 791 2362 795 2363
rect 791 2357 795 2358
rect 799 2362 803 2363
rect 799 2357 803 2358
rect 911 2362 915 2363
rect 911 2357 915 2358
rect 927 2362 931 2363
rect 927 2357 931 2358
rect 1023 2362 1027 2363
rect 1023 2357 1027 2358
rect 1055 2362 1059 2363
rect 1055 2357 1059 2358
rect 1135 2362 1139 2363
rect 1135 2357 1139 2358
rect 1183 2362 1187 2363
rect 1183 2357 1187 2358
rect 1247 2362 1251 2363
rect 1247 2357 1251 2358
rect 1319 2362 1323 2363
rect 1319 2357 1323 2358
rect 1367 2362 1371 2363
rect 1367 2357 1371 2358
rect 1455 2362 1459 2363
rect 1455 2357 1459 2358
rect 1831 2362 1835 2363
rect 1831 2357 1835 2358
rect 112 2329 114 2357
rect 224 2347 226 2357
rect 328 2347 330 2357
rect 440 2347 442 2357
rect 560 2347 562 2357
rect 680 2347 682 2357
rect 800 2347 802 2357
rect 912 2347 914 2357
rect 1024 2347 1026 2357
rect 1136 2347 1138 2357
rect 1248 2347 1250 2357
rect 1368 2347 1370 2357
rect 222 2346 228 2347
rect 222 2342 223 2346
rect 227 2342 228 2346
rect 222 2341 228 2342
rect 326 2346 332 2347
rect 326 2342 327 2346
rect 331 2342 332 2346
rect 326 2341 332 2342
rect 438 2346 444 2347
rect 438 2342 439 2346
rect 443 2342 444 2346
rect 438 2341 444 2342
rect 558 2346 564 2347
rect 558 2342 559 2346
rect 563 2342 564 2346
rect 558 2341 564 2342
rect 678 2346 684 2347
rect 678 2342 679 2346
rect 683 2342 684 2346
rect 678 2341 684 2342
rect 798 2346 804 2347
rect 798 2342 799 2346
rect 803 2342 804 2346
rect 798 2341 804 2342
rect 910 2346 916 2347
rect 910 2342 911 2346
rect 915 2342 916 2346
rect 910 2341 916 2342
rect 1022 2346 1028 2347
rect 1022 2342 1023 2346
rect 1027 2342 1028 2346
rect 1022 2341 1028 2342
rect 1134 2346 1140 2347
rect 1134 2342 1135 2346
rect 1139 2342 1140 2346
rect 1134 2341 1140 2342
rect 1246 2346 1252 2347
rect 1246 2342 1247 2346
rect 1251 2342 1252 2346
rect 1246 2341 1252 2342
rect 1366 2346 1372 2347
rect 1366 2342 1367 2346
rect 1371 2342 1372 2346
rect 1366 2341 1372 2342
rect 1832 2329 1834 2357
rect 1872 2347 1874 2379
rect 1982 2366 1988 2367
rect 1982 2362 1983 2366
rect 1987 2362 1988 2366
rect 1982 2361 1988 2362
rect 2094 2366 2100 2367
rect 2094 2362 2095 2366
rect 2099 2362 2100 2366
rect 2094 2361 2100 2362
rect 2214 2366 2220 2367
rect 2214 2362 2215 2366
rect 2219 2362 2220 2366
rect 2214 2361 2220 2362
rect 2342 2366 2348 2367
rect 2342 2362 2343 2366
rect 2347 2362 2348 2366
rect 2342 2361 2348 2362
rect 2486 2366 2492 2367
rect 2486 2362 2487 2366
rect 2491 2362 2492 2366
rect 2486 2361 2492 2362
rect 2638 2366 2644 2367
rect 2638 2362 2639 2366
rect 2643 2362 2644 2366
rect 2638 2361 2644 2362
rect 2798 2366 2804 2367
rect 2798 2362 2799 2366
rect 2803 2362 2804 2366
rect 2798 2361 2804 2362
rect 2974 2366 2980 2367
rect 2974 2362 2975 2366
rect 2979 2362 2980 2366
rect 2974 2361 2980 2362
rect 3158 2366 3164 2367
rect 3158 2362 3159 2366
rect 3163 2362 3164 2366
rect 3158 2361 3164 2362
rect 3342 2366 3348 2367
rect 3342 2362 3343 2366
rect 3347 2362 3348 2366
rect 3342 2361 3348 2362
rect 3510 2366 3516 2367
rect 3510 2362 3511 2366
rect 3515 2362 3516 2366
rect 3510 2361 3516 2362
rect 1984 2347 1986 2361
rect 2096 2347 2098 2361
rect 2216 2347 2218 2361
rect 2344 2347 2346 2361
rect 2488 2347 2490 2361
rect 2640 2347 2642 2361
rect 2800 2347 2802 2361
rect 2976 2347 2978 2361
rect 3160 2347 3162 2361
rect 3344 2347 3346 2361
rect 3512 2347 3514 2361
rect 3592 2347 3594 2379
rect 1871 2346 1875 2347
rect 1871 2341 1875 2342
rect 1903 2346 1907 2347
rect 1903 2341 1907 2342
rect 1983 2346 1987 2347
rect 1983 2341 1987 2342
rect 2015 2346 2019 2347
rect 2015 2341 2019 2342
rect 2095 2346 2099 2347
rect 2095 2341 2099 2342
rect 2167 2346 2171 2347
rect 2167 2341 2171 2342
rect 2215 2346 2219 2347
rect 2215 2341 2219 2342
rect 2319 2346 2323 2347
rect 2319 2341 2323 2342
rect 2343 2346 2347 2347
rect 2343 2341 2347 2342
rect 2471 2346 2475 2347
rect 2471 2341 2475 2342
rect 2487 2346 2491 2347
rect 2487 2341 2491 2342
rect 2623 2346 2627 2347
rect 2623 2341 2627 2342
rect 2639 2346 2643 2347
rect 2639 2341 2643 2342
rect 2775 2346 2779 2347
rect 2775 2341 2779 2342
rect 2799 2346 2803 2347
rect 2799 2341 2803 2342
rect 2927 2346 2931 2347
rect 2927 2341 2931 2342
rect 2975 2346 2979 2347
rect 2975 2341 2979 2342
rect 3087 2346 3091 2347
rect 3087 2341 3091 2342
rect 3159 2346 3163 2347
rect 3159 2341 3163 2342
rect 3247 2346 3251 2347
rect 3247 2341 3251 2342
rect 3343 2346 3347 2347
rect 3343 2341 3347 2342
rect 3415 2346 3419 2347
rect 3415 2341 3419 2342
rect 3511 2346 3515 2347
rect 3511 2341 3515 2342
rect 3591 2346 3595 2347
rect 3591 2341 3595 2342
rect 110 2328 116 2329
rect 110 2324 111 2328
rect 115 2324 116 2328
rect 110 2323 116 2324
rect 1830 2328 1836 2329
rect 1830 2324 1831 2328
rect 1835 2324 1836 2328
rect 1830 2323 1836 2324
rect 1872 2313 1874 2341
rect 1904 2331 1906 2341
rect 2016 2331 2018 2341
rect 2168 2331 2170 2341
rect 2320 2331 2322 2341
rect 2472 2331 2474 2341
rect 2624 2331 2626 2341
rect 2776 2331 2778 2341
rect 2928 2331 2930 2341
rect 3088 2331 3090 2341
rect 3248 2331 3250 2341
rect 3416 2331 3418 2341
rect 1902 2330 1908 2331
rect 1902 2326 1903 2330
rect 1907 2326 1908 2330
rect 1902 2325 1908 2326
rect 2014 2330 2020 2331
rect 2014 2326 2015 2330
rect 2019 2326 2020 2330
rect 2014 2325 2020 2326
rect 2166 2330 2172 2331
rect 2166 2326 2167 2330
rect 2171 2326 2172 2330
rect 2166 2325 2172 2326
rect 2318 2330 2324 2331
rect 2318 2326 2319 2330
rect 2323 2326 2324 2330
rect 2318 2325 2324 2326
rect 2470 2330 2476 2331
rect 2470 2326 2471 2330
rect 2475 2326 2476 2330
rect 2470 2325 2476 2326
rect 2622 2330 2628 2331
rect 2622 2326 2623 2330
rect 2627 2326 2628 2330
rect 2622 2325 2628 2326
rect 2774 2330 2780 2331
rect 2774 2326 2775 2330
rect 2779 2326 2780 2330
rect 2774 2325 2780 2326
rect 2926 2330 2932 2331
rect 2926 2326 2927 2330
rect 2931 2326 2932 2330
rect 2926 2325 2932 2326
rect 3086 2330 3092 2331
rect 3086 2326 3087 2330
rect 3091 2326 3092 2330
rect 3086 2325 3092 2326
rect 3246 2330 3252 2331
rect 3246 2326 3247 2330
rect 3251 2326 3252 2330
rect 3246 2325 3252 2326
rect 3414 2330 3420 2331
rect 3414 2326 3415 2330
rect 3419 2326 3420 2330
rect 3414 2325 3420 2326
rect 3592 2313 3594 2341
rect 1870 2312 1876 2313
rect 110 2311 116 2312
rect 110 2307 111 2311
rect 115 2307 116 2311
rect 1830 2311 1836 2312
rect 110 2306 116 2307
rect 214 2308 220 2309
rect 112 2275 114 2306
rect 214 2304 215 2308
rect 219 2304 220 2308
rect 214 2303 220 2304
rect 318 2308 324 2309
rect 318 2304 319 2308
rect 323 2304 324 2308
rect 318 2303 324 2304
rect 430 2308 436 2309
rect 430 2304 431 2308
rect 435 2304 436 2308
rect 430 2303 436 2304
rect 550 2308 556 2309
rect 550 2304 551 2308
rect 555 2304 556 2308
rect 550 2303 556 2304
rect 670 2308 676 2309
rect 670 2304 671 2308
rect 675 2304 676 2308
rect 670 2303 676 2304
rect 790 2308 796 2309
rect 790 2304 791 2308
rect 795 2304 796 2308
rect 790 2303 796 2304
rect 902 2308 908 2309
rect 902 2304 903 2308
rect 907 2304 908 2308
rect 902 2303 908 2304
rect 1014 2308 1020 2309
rect 1014 2304 1015 2308
rect 1019 2304 1020 2308
rect 1014 2303 1020 2304
rect 1126 2308 1132 2309
rect 1126 2304 1127 2308
rect 1131 2304 1132 2308
rect 1126 2303 1132 2304
rect 1238 2308 1244 2309
rect 1238 2304 1239 2308
rect 1243 2304 1244 2308
rect 1238 2303 1244 2304
rect 1358 2308 1364 2309
rect 1358 2304 1359 2308
rect 1363 2304 1364 2308
rect 1830 2307 1831 2311
rect 1835 2307 1836 2311
rect 1870 2308 1871 2312
rect 1875 2308 1876 2312
rect 1870 2307 1876 2308
rect 3590 2312 3596 2313
rect 3590 2308 3591 2312
rect 3595 2308 3596 2312
rect 3590 2307 3596 2308
rect 1830 2306 1836 2307
rect 1358 2303 1364 2304
rect 216 2275 218 2303
rect 320 2275 322 2303
rect 432 2275 434 2303
rect 552 2275 554 2303
rect 672 2275 674 2303
rect 792 2275 794 2303
rect 904 2275 906 2303
rect 1016 2275 1018 2303
rect 1128 2275 1130 2303
rect 1240 2275 1242 2303
rect 1360 2275 1362 2303
rect 1832 2275 1834 2306
rect 1870 2295 1876 2296
rect 1870 2291 1871 2295
rect 1875 2291 1876 2295
rect 3590 2295 3596 2296
rect 1870 2290 1876 2291
rect 1894 2292 1900 2293
rect 111 2274 115 2275
rect 111 2269 115 2270
rect 215 2274 219 2275
rect 215 2269 219 2270
rect 311 2274 315 2275
rect 311 2269 315 2270
rect 319 2274 323 2275
rect 319 2269 323 2270
rect 407 2274 411 2275
rect 407 2269 411 2270
rect 431 2274 435 2275
rect 431 2269 435 2270
rect 503 2274 507 2275
rect 503 2269 507 2270
rect 551 2274 555 2275
rect 551 2269 555 2270
rect 607 2274 611 2275
rect 607 2269 611 2270
rect 671 2274 675 2275
rect 671 2269 675 2270
rect 711 2274 715 2275
rect 711 2269 715 2270
rect 791 2274 795 2275
rect 791 2269 795 2270
rect 815 2274 819 2275
rect 815 2269 819 2270
rect 903 2274 907 2275
rect 903 2269 907 2270
rect 911 2274 915 2275
rect 911 2269 915 2270
rect 1007 2274 1011 2275
rect 1007 2269 1011 2270
rect 1015 2274 1019 2275
rect 1015 2269 1019 2270
rect 1103 2274 1107 2275
rect 1103 2269 1107 2270
rect 1127 2274 1131 2275
rect 1127 2269 1131 2270
rect 1199 2274 1203 2275
rect 1199 2269 1203 2270
rect 1239 2274 1243 2275
rect 1239 2269 1243 2270
rect 1303 2274 1307 2275
rect 1303 2269 1307 2270
rect 1359 2274 1363 2275
rect 1359 2269 1363 2270
rect 1831 2274 1835 2275
rect 1872 2271 1874 2290
rect 1894 2288 1895 2292
rect 1899 2288 1900 2292
rect 1894 2287 1900 2288
rect 2006 2292 2012 2293
rect 2006 2288 2007 2292
rect 2011 2288 2012 2292
rect 2006 2287 2012 2288
rect 2158 2292 2164 2293
rect 2158 2288 2159 2292
rect 2163 2288 2164 2292
rect 2158 2287 2164 2288
rect 2310 2292 2316 2293
rect 2310 2288 2311 2292
rect 2315 2288 2316 2292
rect 2310 2287 2316 2288
rect 2462 2292 2468 2293
rect 2462 2288 2463 2292
rect 2467 2288 2468 2292
rect 2462 2287 2468 2288
rect 2614 2292 2620 2293
rect 2614 2288 2615 2292
rect 2619 2288 2620 2292
rect 2614 2287 2620 2288
rect 2766 2292 2772 2293
rect 2766 2288 2767 2292
rect 2771 2288 2772 2292
rect 2766 2287 2772 2288
rect 2918 2292 2924 2293
rect 2918 2288 2919 2292
rect 2923 2288 2924 2292
rect 2918 2287 2924 2288
rect 3078 2292 3084 2293
rect 3078 2288 3079 2292
rect 3083 2288 3084 2292
rect 3078 2287 3084 2288
rect 3238 2292 3244 2293
rect 3238 2288 3239 2292
rect 3243 2288 3244 2292
rect 3238 2287 3244 2288
rect 3406 2292 3412 2293
rect 3406 2288 3407 2292
rect 3411 2288 3412 2292
rect 3590 2291 3591 2295
rect 3595 2291 3596 2295
rect 3590 2290 3596 2291
rect 3406 2287 3412 2288
rect 1896 2271 1898 2287
rect 2008 2271 2010 2287
rect 2160 2271 2162 2287
rect 2312 2271 2314 2287
rect 2464 2271 2466 2287
rect 2616 2271 2618 2287
rect 2768 2271 2770 2287
rect 2920 2271 2922 2287
rect 3080 2271 3082 2287
rect 3240 2271 3242 2287
rect 3408 2271 3410 2287
rect 3592 2271 3594 2290
rect 1831 2269 1835 2270
rect 1871 2270 1875 2271
rect 112 2250 114 2269
rect 312 2253 314 2269
rect 408 2253 410 2269
rect 504 2253 506 2269
rect 608 2253 610 2269
rect 712 2253 714 2269
rect 816 2253 818 2269
rect 912 2253 914 2269
rect 1008 2253 1010 2269
rect 1104 2253 1106 2269
rect 1200 2253 1202 2269
rect 1304 2253 1306 2269
rect 310 2252 316 2253
rect 110 2249 116 2250
rect 110 2245 111 2249
rect 115 2245 116 2249
rect 310 2248 311 2252
rect 315 2248 316 2252
rect 310 2247 316 2248
rect 406 2252 412 2253
rect 406 2248 407 2252
rect 411 2248 412 2252
rect 406 2247 412 2248
rect 502 2252 508 2253
rect 502 2248 503 2252
rect 507 2248 508 2252
rect 502 2247 508 2248
rect 606 2252 612 2253
rect 606 2248 607 2252
rect 611 2248 612 2252
rect 606 2247 612 2248
rect 710 2252 716 2253
rect 710 2248 711 2252
rect 715 2248 716 2252
rect 710 2247 716 2248
rect 814 2252 820 2253
rect 814 2248 815 2252
rect 819 2248 820 2252
rect 814 2247 820 2248
rect 910 2252 916 2253
rect 910 2248 911 2252
rect 915 2248 916 2252
rect 910 2247 916 2248
rect 1006 2252 1012 2253
rect 1006 2248 1007 2252
rect 1011 2248 1012 2252
rect 1006 2247 1012 2248
rect 1102 2252 1108 2253
rect 1102 2248 1103 2252
rect 1107 2248 1108 2252
rect 1102 2247 1108 2248
rect 1198 2252 1204 2253
rect 1198 2248 1199 2252
rect 1203 2248 1204 2252
rect 1198 2247 1204 2248
rect 1302 2252 1308 2253
rect 1302 2248 1303 2252
rect 1307 2248 1308 2252
rect 1832 2250 1834 2269
rect 1871 2265 1875 2266
rect 1895 2270 1899 2271
rect 1895 2265 1899 2266
rect 2007 2270 2011 2271
rect 2007 2265 2011 2266
rect 2031 2270 2035 2271
rect 2031 2265 2035 2266
rect 2159 2270 2163 2271
rect 2159 2265 2163 2266
rect 2207 2270 2211 2271
rect 2207 2265 2211 2266
rect 2311 2270 2315 2271
rect 2311 2265 2315 2266
rect 2391 2270 2395 2271
rect 2391 2265 2395 2266
rect 2463 2270 2467 2271
rect 2463 2265 2467 2266
rect 2575 2270 2579 2271
rect 2575 2265 2579 2266
rect 2615 2270 2619 2271
rect 2615 2265 2619 2266
rect 2767 2270 2771 2271
rect 2767 2265 2771 2266
rect 2919 2270 2923 2271
rect 2919 2265 2923 2266
rect 2951 2270 2955 2271
rect 2951 2265 2955 2266
rect 3079 2270 3083 2271
rect 3079 2265 3083 2266
rect 3143 2270 3147 2271
rect 3143 2265 3147 2266
rect 3239 2270 3243 2271
rect 3239 2265 3243 2266
rect 3335 2270 3339 2271
rect 3335 2265 3339 2266
rect 3407 2270 3411 2271
rect 3407 2265 3411 2266
rect 3503 2270 3507 2271
rect 3503 2265 3507 2266
rect 3591 2270 3595 2271
rect 3591 2265 3595 2266
rect 1302 2247 1308 2248
rect 1830 2249 1836 2250
rect 110 2244 116 2245
rect 1830 2245 1831 2249
rect 1835 2245 1836 2249
rect 1872 2246 1874 2265
rect 1896 2249 1898 2265
rect 2032 2249 2034 2265
rect 2208 2249 2210 2265
rect 2392 2249 2394 2265
rect 2576 2249 2578 2265
rect 2768 2249 2770 2265
rect 2952 2249 2954 2265
rect 3144 2249 3146 2265
rect 3336 2249 3338 2265
rect 3504 2249 3506 2265
rect 1894 2248 1900 2249
rect 1830 2244 1836 2245
rect 1870 2245 1876 2246
rect 1870 2241 1871 2245
rect 1875 2241 1876 2245
rect 1894 2244 1895 2248
rect 1899 2244 1900 2248
rect 1894 2243 1900 2244
rect 2030 2248 2036 2249
rect 2030 2244 2031 2248
rect 2035 2244 2036 2248
rect 2030 2243 2036 2244
rect 2206 2248 2212 2249
rect 2206 2244 2207 2248
rect 2211 2244 2212 2248
rect 2206 2243 2212 2244
rect 2390 2248 2396 2249
rect 2390 2244 2391 2248
rect 2395 2244 2396 2248
rect 2390 2243 2396 2244
rect 2574 2248 2580 2249
rect 2574 2244 2575 2248
rect 2579 2244 2580 2248
rect 2574 2243 2580 2244
rect 2766 2248 2772 2249
rect 2766 2244 2767 2248
rect 2771 2244 2772 2248
rect 2766 2243 2772 2244
rect 2950 2248 2956 2249
rect 2950 2244 2951 2248
rect 2955 2244 2956 2248
rect 2950 2243 2956 2244
rect 3142 2248 3148 2249
rect 3142 2244 3143 2248
rect 3147 2244 3148 2248
rect 3142 2243 3148 2244
rect 3334 2248 3340 2249
rect 3334 2244 3335 2248
rect 3339 2244 3340 2248
rect 3334 2243 3340 2244
rect 3502 2248 3508 2249
rect 3502 2244 3503 2248
rect 3507 2244 3508 2248
rect 3592 2246 3594 2265
rect 3502 2243 3508 2244
rect 3590 2245 3596 2246
rect 1870 2240 1876 2241
rect 3590 2241 3591 2245
rect 3595 2241 3596 2245
rect 3590 2240 3596 2241
rect 110 2232 116 2233
rect 110 2228 111 2232
rect 115 2228 116 2232
rect 110 2227 116 2228
rect 1830 2232 1836 2233
rect 1830 2228 1831 2232
rect 1835 2228 1836 2232
rect 1830 2227 1836 2228
rect 1870 2228 1876 2229
rect 112 2195 114 2227
rect 318 2214 324 2215
rect 318 2210 319 2214
rect 323 2210 324 2214
rect 318 2209 324 2210
rect 414 2214 420 2215
rect 414 2210 415 2214
rect 419 2210 420 2214
rect 414 2209 420 2210
rect 510 2214 516 2215
rect 510 2210 511 2214
rect 515 2210 516 2214
rect 510 2209 516 2210
rect 614 2214 620 2215
rect 614 2210 615 2214
rect 619 2210 620 2214
rect 614 2209 620 2210
rect 718 2214 724 2215
rect 718 2210 719 2214
rect 723 2210 724 2214
rect 718 2209 724 2210
rect 822 2214 828 2215
rect 822 2210 823 2214
rect 827 2210 828 2214
rect 822 2209 828 2210
rect 918 2214 924 2215
rect 918 2210 919 2214
rect 923 2210 924 2214
rect 918 2209 924 2210
rect 1014 2214 1020 2215
rect 1014 2210 1015 2214
rect 1019 2210 1020 2214
rect 1014 2209 1020 2210
rect 1110 2214 1116 2215
rect 1110 2210 1111 2214
rect 1115 2210 1116 2214
rect 1110 2209 1116 2210
rect 1206 2214 1212 2215
rect 1206 2210 1207 2214
rect 1211 2210 1212 2214
rect 1206 2209 1212 2210
rect 1310 2214 1316 2215
rect 1310 2210 1311 2214
rect 1315 2210 1316 2214
rect 1310 2209 1316 2210
rect 320 2195 322 2209
rect 416 2195 418 2209
rect 512 2195 514 2209
rect 616 2195 618 2209
rect 720 2195 722 2209
rect 824 2195 826 2209
rect 920 2195 922 2209
rect 1016 2195 1018 2209
rect 1112 2195 1114 2209
rect 1208 2195 1210 2209
rect 1312 2195 1314 2209
rect 1832 2195 1834 2227
rect 1870 2224 1871 2228
rect 1875 2224 1876 2228
rect 1870 2223 1876 2224
rect 3590 2228 3596 2229
rect 3590 2224 3591 2228
rect 3595 2224 3596 2228
rect 3590 2223 3596 2224
rect 111 2194 115 2195
rect 111 2189 115 2190
rect 319 2194 323 2195
rect 319 2189 323 2190
rect 415 2194 419 2195
rect 415 2189 419 2190
rect 511 2194 515 2195
rect 511 2189 515 2190
rect 519 2194 523 2195
rect 519 2189 523 2190
rect 615 2194 619 2195
rect 615 2189 619 2190
rect 623 2194 627 2195
rect 623 2189 627 2190
rect 719 2194 723 2195
rect 719 2189 723 2190
rect 727 2194 731 2195
rect 727 2189 731 2190
rect 823 2194 827 2195
rect 823 2189 827 2190
rect 831 2194 835 2195
rect 831 2189 835 2190
rect 919 2194 923 2195
rect 919 2189 923 2190
rect 935 2194 939 2195
rect 935 2189 939 2190
rect 1015 2194 1019 2195
rect 1015 2189 1019 2190
rect 1039 2194 1043 2195
rect 1039 2189 1043 2190
rect 1111 2194 1115 2195
rect 1111 2189 1115 2190
rect 1151 2194 1155 2195
rect 1151 2189 1155 2190
rect 1207 2194 1211 2195
rect 1207 2189 1211 2190
rect 1263 2194 1267 2195
rect 1263 2189 1267 2190
rect 1311 2194 1315 2195
rect 1311 2189 1315 2190
rect 1831 2194 1835 2195
rect 1831 2189 1835 2190
rect 112 2161 114 2189
rect 320 2179 322 2189
rect 416 2179 418 2189
rect 520 2179 522 2189
rect 624 2179 626 2189
rect 728 2179 730 2189
rect 832 2179 834 2189
rect 936 2179 938 2189
rect 1040 2179 1042 2189
rect 1152 2179 1154 2189
rect 1264 2179 1266 2189
rect 318 2178 324 2179
rect 318 2174 319 2178
rect 323 2174 324 2178
rect 318 2173 324 2174
rect 414 2178 420 2179
rect 414 2174 415 2178
rect 419 2174 420 2178
rect 414 2173 420 2174
rect 518 2178 524 2179
rect 518 2174 519 2178
rect 523 2174 524 2178
rect 518 2173 524 2174
rect 622 2178 628 2179
rect 622 2174 623 2178
rect 627 2174 628 2178
rect 622 2173 628 2174
rect 726 2178 732 2179
rect 726 2174 727 2178
rect 731 2174 732 2178
rect 726 2173 732 2174
rect 830 2178 836 2179
rect 830 2174 831 2178
rect 835 2174 836 2178
rect 830 2173 836 2174
rect 934 2178 940 2179
rect 934 2174 935 2178
rect 939 2174 940 2178
rect 934 2173 940 2174
rect 1038 2178 1044 2179
rect 1038 2174 1039 2178
rect 1043 2174 1044 2178
rect 1038 2173 1044 2174
rect 1150 2178 1156 2179
rect 1150 2174 1151 2178
rect 1155 2174 1156 2178
rect 1150 2173 1156 2174
rect 1262 2178 1268 2179
rect 1262 2174 1263 2178
rect 1267 2174 1268 2178
rect 1262 2173 1268 2174
rect 1832 2161 1834 2189
rect 1872 2187 1874 2223
rect 1902 2210 1908 2211
rect 1902 2206 1903 2210
rect 1907 2206 1908 2210
rect 1902 2205 1908 2206
rect 2038 2210 2044 2211
rect 2038 2206 2039 2210
rect 2043 2206 2044 2210
rect 2038 2205 2044 2206
rect 2214 2210 2220 2211
rect 2214 2206 2215 2210
rect 2219 2206 2220 2210
rect 2214 2205 2220 2206
rect 2398 2210 2404 2211
rect 2398 2206 2399 2210
rect 2403 2206 2404 2210
rect 2398 2205 2404 2206
rect 2582 2210 2588 2211
rect 2582 2206 2583 2210
rect 2587 2206 2588 2210
rect 2582 2205 2588 2206
rect 2774 2210 2780 2211
rect 2774 2206 2775 2210
rect 2779 2206 2780 2210
rect 2774 2205 2780 2206
rect 2958 2210 2964 2211
rect 2958 2206 2959 2210
rect 2963 2206 2964 2210
rect 2958 2205 2964 2206
rect 3150 2210 3156 2211
rect 3150 2206 3151 2210
rect 3155 2206 3156 2210
rect 3150 2205 3156 2206
rect 3342 2210 3348 2211
rect 3342 2206 3343 2210
rect 3347 2206 3348 2210
rect 3342 2205 3348 2206
rect 3510 2210 3516 2211
rect 3510 2206 3511 2210
rect 3515 2206 3516 2210
rect 3510 2205 3516 2206
rect 1904 2187 1906 2205
rect 2040 2187 2042 2205
rect 2216 2187 2218 2205
rect 2400 2187 2402 2205
rect 2584 2187 2586 2205
rect 2776 2187 2778 2205
rect 2960 2187 2962 2205
rect 3152 2187 3154 2205
rect 3344 2187 3346 2205
rect 3512 2187 3514 2205
rect 3592 2187 3594 2223
rect 1871 2186 1875 2187
rect 1871 2181 1875 2182
rect 1903 2186 1907 2187
rect 1903 2181 1907 2182
rect 1967 2186 1971 2187
rect 1967 2181 1971 2182
rect 2039 2186 2043 2187
rect 2039 2181 2043 2182
rect 2079 2186 2083 2187
rect 2079 2181 2083 2182
rect 2215 2186 2219 2187
rect 2215 2181 2219 2182
rect 2367 2186 2371 2187
rect 2367 2181 2371 2182
rect 2399 2186 2403 2187
rect 2399 2181 2403 2182
rect 2527 2186 2531 2187
rect 2527 2181 2531 2182
rect 2583 2186 2587 2187
rect 2583 2181 2587 2182
rect 2687 2186 2691 2187
rect 2687 2181 2691 2182
rect 2775 2186 2779 2187
rect 2775 2181 2779 2182
rect 2847 2186 2851 2187
rect 2847 2181 2851 2182
rect 2959 2186 2963 2187
rect 2959 2181 2963 2182
rect 2991 2186 2995 2187
rect 2991 2181 2995 2182
rect 3127 2186 3131 2187
rect 3127 2181 3131 2182
rect 3151 2186 3155 2187
rect 3151 2181 3155 2182
rect 3263 2186 3267 2187
rect 3263 2181 3267 2182
rect 3343 2186 3347 2187
rect 3343 2181 3347 2182
rect 3399 2186 3403 2187
rect 3399 2181 3403 2182
rect 3511 2186 3515 2187
rect 3511 2181 3515 2182
rect 3591 2186 3595 2187
rect 3591 2181 3595 2182
rect 110 2160 116 2161
rect 110 2156 111 2160
rect 115 2156 116 2160
rect 110 2155 116 2156
rect 1830 2160 1836 2161
rect 1830 2156 1831 2160
rect 1835 2156 1836 2160
rect 1830 2155 1836 2156
rect 1872 2153 1874 2181
rect 1968 2171 1970 2181
rect 2080 2171 2082 2181
rect 2216 2171 2218 2181
rect 2368 2171 2370 2181
rect 2528 2171 2530 2181
rect 2688 2171 2690 2181
rect 2848 2171 2850 2181
rect 2992 2171 2994 2181
rect 3128 2171 3130 2181
rect 3264 2171 3266 2181
rect 3400 2171 3402 2181
rect 3512 2171 3514 2181
rect 1966 2170 1972 2171
rect 1966 2166 1967 2170
rect 1971 2166 1972 2170
rect 1966 2165 1972 2166
rect 2078 2170 2084 2171
rect 2078 2166 2079 2170
rect 2083 2166 2084 2170
rect 2078 2165 2084 2166
rect 2214 2170 2220 2171
rect 2214 2166 2215 2170
rect 2219 2166 2220 2170
rect 2214 2165 2220 2166
rect 2366 2170 2372 2171
rect 2366 2166 2367 2170
rect 2371 2166 2372 2170
rect 2366 2165 2372 2166
rect 2526 2170 2532 2171
rect 2526 2166 2527 2170
rect 2531 2166 2532 2170
rect 2526 2165 2532 2166
rect 2686 2170 2692 2171
rect 2686 2166 2687 2170
rect 2691 2166 2692 2170
rect 2686 2165 2692 2166
rect 2846 2170 2852 2171
rect 2846 2166 2847 2170
rect 2851 2166 2852 2170
rect 2846 2165 2852 2166
rect 2990 2170 2996 2171
rect 2990 2166 2991 2170
rect 2995 2166 2996 2170
rect 2990 2165 2996 2166
rect 3126 2170 3132 2171
rect 3126 2166 3127 2170
rect 3131 2166 3132 2170
rect 3126 2165 3132 2166
rect 3262 2170 3268 2171
rect 3262 2166 3263 2170
rect 3267 2166 3268 2170
rect 3262 2165 3268 2166
rect 3398 2170 3404 2171
rect 3398 2166 3399 2170
rect 3403 2166 3404 2170
rect 3398 2165 3404 2166
rect 3510 2170 3516 2171
rect 3510 2166 3511 2170
rect 3515 2166 3516 2170
rect 3510 2165 3516 2166
rect 3592 2153 3594 2181
rect 1870 2152 1876 2153
rect 1870 2148 1871 2152
rect 1875 2148 1876 2152
rect 1870 2147 1876 2148
rect 3590 2152 3596 2153
rect 3590 2148 3591 2152
rect 3595 2148 3596 2152
rect 3590 2147 3596 2148
rect 110 2143 116 2144
rect 110 2139 111 2143
rect 115 2139 116 2143
rect 1830 2143 1836 2144
rect 110 2138 116 2139
rect 310 2140 316 2141
rect 112 2119 114 2138
rect 310 2136 311 2140
rect 315 2136 316 2140
rect 310 2135 316 2136
rect 406 2140 412 2141
rect 406 2136 407 2140
rect 411 2136 412 2140
rect 406 2135 412 2136
rect 510 2140 516 2141
rect 510 2136 511 2140
rect 515 2136 516 2140
rect 510 2135 516 2136
rect 614 2140 620 2141
rect 614 2136 615 2140
rect 619 2136 620 2140
rect 614 2135 620 2136
rect 718 2140 724 2141
rect 718 2136 719 2140
rect 723 2136 724 2140
rect 718 2135 724 2136
rect 822 2140 828 2141
rect 822 2136 823 2140
rect 827 2136 828 2140
rect 822 2135 828 2136
rect 926 2140 932 2141
rect 926 2136 927 2140
rect 931 2136 932 2140
rect 926 2135 932 2136
rect 1030 2140 1036 2141
rect 1030 2136 1031 2140
rect 1035 2136 1036 2140
rect 1030 2135 1036 2136
rect 1142 2140 1148 2141
rect 1142 2136 1143 2140
rect 1147 2136 1148 2140
rect 1142 2135 1148 2136
rect 1254 2140 1260 2141
rect 1254 2136 1255 2140
rect 1259 2136 1260 2140
rect 1830 2139 1831 2143
rect 1835 2139 1836 2143
rect 1830 2138 1836 2139
rect 1254 2135 1260 2136
rect 312 2119 314 2135
rect 408 2119 410 2135
rect 512 2119 514 2135
rect 616 2119 618 2135
rect 720 2119 722 2135
rect 824 2119 826 2135
rect 928 2119 930 2135
rect 1032 2119 1034 2135
rect 1144 2119 1146 2135
rect 1256 2119 1258 2135
rect 1832 2119 1834 2138
rect 1870 2135 1876 2136
rect 1870 2131 1871 2135
rect 1875 2131 1876 2135
rect 3590 2135 3596 2136
rect 1870 2130 1876 2131
rect 1958 2132 1964 2133
rect 111 2118 115 2119
rect 111 2113 115 2114
rect 279 2118 283 2119
rect 279 2113 283 2114
rect 311 2118 315 2119
rect 311 2113 315 2114
rect 399 2118 403 2119
rect 399 2113 403 2114
rect 407 2118 411 2119
rect 407 2113 411 2114
rect 511 2118 515 2119
rect 511 2113 515 2114
rect 615 2118 619 2119
rect 615 2113 619 2114
rect 623 2118 627 2119
rect 623 2113 627 2114
rect 719 2118 723 2119
rect 719 2113 723 2114
rect 735 2118 739 2119
rect 735 2113 739 2114
rect 823 2118 827 2119
rect 823 2113 827 2114
rect 847 2118 851 2119
rect 847 2113 851 2114
rect 927 2118 931 2119
rect 927 2113 931 2114
rect 951 2118 955 2119
rect 951 2113 955 2114
rect 1031 2118 1035 2119
rect 1031 2113 1035 2114
rect 1047 2118 1051 2119
rect 1047 2113 1051 2114
rect 1143 2118 1147 2119
rect 1143 2113 1147 2114
rect 1239 2118 1243 2119
rect 1239 2113 1243 2114
rect 1255 2118 1259 2119
rect 1255 2113 1259 2114
rect 1343 2118 1347 2119
rect 1343 2113 1347 2114
rect 1831 2118 1835 2119
rect 1831 2113 1835 2114
rect 112 2094 114 2113
rect 280 2097 282 2113
rect 400 2097 402 2113
rect 512 2097 514 2113
rect 624 2097 626 2113
rect 736 2097 738 2113
rect 848 2097 850 2113
rect 952 2097 954 2113
rect 1048 2097 1050 2113
rect 1144 2097 1146 2113
rect 1240 2097 1242 2113
rect 1344 2097 1346 2113
rect 278 2096 284 2097
rect 110 2093 116 2094
rect 110 2089 111 2093
rect 115 2089 116 2093
rect 278 2092 279 2096
rect 283 2092 284 2096
rect 278 2091 284 2092
rect 398 2096 404 2097
rect 398 2092 399 2096
rect 403 2092 404 2096
rect 398 2091 404 2092
rect 510 2096 516 2097
rect 510 2092 511 2096
rect 515 2092 516 2096
rect 510 2091 516 2092
rect 622 2096 628 2097
rect 622 2092 623 2096
rect 627 2092 628 2096
rect 622 2091 628 2092
rect 734 2096 740 2097
rect 734 2092 735 2096
rect 739 2092 740 2096
rect 734 2091 740 2092
rect 846 2096 852 2097
rect 846 2092 847 2096
rect 851 2092 852 2096
rect 846 2091 852 2092
rect 950 2096 956 2097
rect 950 2092 951 2096
rect 955 2092 956 2096
rect 950 2091 956 2092
rect 1046 2096 1052 2097
rect 1046 2092 1047 2096
rect 1051 2092 1052 2096
rect 1046 2091 1052 2092
rect 1142 2096 1148 2097
rect 1142 2092 1143 2096
rect 1147 2092 1148 2096
rect 1142 2091 1148 2092
rect 1238 2096 1244 2097
rect 1238 2092 1239 2096
rect 1243 2092 1244 2096
rect 1238 2091 1244 2092
rect 1342 2096 1348 2097
rect 1342 2092 1343 2096
rect 1347 2092 1348 2096
rect 1832 2094 1834 2113
rect 1872 2111 1874 2130
rect 1958 2128 1959 2132
rect 1963 2128 1964 2132
rect 1958 2127 1964 2128
rect 2070 2132 2076 2133
rect 2070 2128 2071 2132
rect 2075 2128 2076 2132
rect 2070 2127 2076 2128
rect 2206 2132 2212 2133
rect 2206 2128 2207 2132
rect 2211 2128 2212 2132
rect 2206 2127 2212 2128
rect 2358 2132 2364 2133
rect 2358 2128 2359 2132
rect 2363 2128 2364 2132
rect 2358 2127 2364 2128
rect 2518 2132 2524 2133
rect 2518 2128 2519 2132
rect 2523 2128 2524 2132
rect 2518 2127 2524 2128
rect 2678 2132 2684 2133
rect 2678 2128 2679 2132
rect 2683 2128 2684 2132
rect 2678 2127 2684 2128
rect 2838 2132 2844 2133
rect 2838 2128 2839 2132
rect 2843 2128 2844 2132
rect 2838 2127 2844 2128
rect 2982 2132 2988 2133
rect 2982 2128 2983 2132
rect 2987 2128 2988 2132
rect 2982 2127 2988 2128
rect 3118 2132 3124 2133
rect 3118 2128 3119 2132
rect 3123 2128 3124 2132
rect 3118 2127 3124 2128
rect 3254 2132 3260 2133
rect 3254 2128 3255 2132
rect 3259 2128 3260 2132
rect 3254 2127 3260 2128
rect 3390 2132 3396 2133
rect 3390 2128 3391 2132
rect 3395 2128 3396 2132
rect 3390 2127 3396 2128
rect 3502 2132 3508 2133
rect 3502 2128 3503 2132
rect 3507 2128 3508 2132
rect 3590 2131 3591 2135
rect 3595 2131 3596 2135
rect 3590 2130 3596 2131
rect 3502 2127 3508 2128
rect 1960 2111 1962 2127
rect 2072 2111 2074 2127
rect 2208 2111 2210 2127
rect 2360 2111 2362 2127
rect 2520 2111 2522 2127
rect 2680 2111 2682 2127
rect 2840 2111 2842 2127
rect 2984 2111 2986 2127
rect 3120 2111 3122 2127
rect 3256 2111 3258 2127
rect 3392 2111 3394 2127
rect 3504 2111 3506 2127
rect 3592 2111 3594 2130
rect 1871 2110 1875 2111
rect 1871 2105 1875 2106
rect 1959 2110 1963 2111
rect 1959 2105 1963 2106
rect 2071 2110 2075 2111
rect 2071 2105 2075 2106
rect 2207 2110 2211 2111
rect 2207 2105 2211 2106
rect 2287 2110 2291 2111
rect 2287 2105 2291 2106
rect 2359 2110 2363 2111
rect 2359 2105 2363 2106
rect 2391 2110 2395 2111
rect 2391 2105 2395 2106
rect 2503 2110 2507 2111
rect 2503 2105 2507 2106
rect 2519 2110 2523 2111
rect 2519 2105 2523 2106
rect 2623 2110 2627 2111
rect 2623 2105 2627 2106
rect 2679 2110 2683 2111
rect 2679 2105 2683 2106
rect 2743 2110 2747 2111
rect 2743 2105 2747 2106
rect 2839 2110 2843 2111
rect 2839 2105 2843 2106
rect 2855 2110 2859 2111
rect 2855 2105 2859 2106
rect 2967 2110 2971 2111
rect 2967 2105 2971 2106
rect 2983 2110 2987 2111
rect 2983 2105 2987 2106
rect 3079 2110 3083 2111
rect 3079 2105 3083 2106
rect 3119 2110 3123 2111
rect 3119 2105 3123 2106
rect 3191 2110 3195 2111
rect 3191 2105 3195 2106
rect 3255 2110 3259 2111
rect 3255 2105 3259 2106
rect 3303 2110 3307 2111
rect 3303 2105 3307 2106
rect 3391 2110 3395 2111
rect 3391 2105 3395 2106
rect 3415 2110 3419 2111
rect 3415 2105 3419 2106
rect 3503 2110 3507 2111
rect 3503 2105 3507 2106
rect 3591 2110 3595 2111
rect 3591 2105 3595 2106
rect 1342 2091 1348 2092
rect 1830 2093 1836 2094
rect 110 2088 116 2089
rect 1830 2089 1831 2093
rect 1835 2089 1836 2093
rect 1830 2088 1836 2089
rect 1872 2086 1874 2105
rect 2288 2089 2290 2105
rect 2392 2089 2394 2105
rect 2504 2089 2506 2105
rect 2624 2089 2626 2105
rect 2744 2089 2746 2105
rect 2856 2089 2858 2105
rect 2968 2089 2970 2105
rect 3080 2089 3082 2105
rect 3192 2089 3194 2105
rect 3304 2089 3306 2105
rect 3416 2089 3418 2105
rect 3504 2089 3506 2105
rect 2286 2088 2292 2089
rect 1870 2085 1876 2086
rect 1870 2081 1871 2085
rect 1875 2081 1876 2085
rect 2286 2084 2287 2088
rect 2291 2084 2292 2088
rect 2286 2083 2292 2084
rect 2390 2088 2396 2089
rect 2390 2084 2391 2088
rect 2395 2084 2396 2088
rect 2390 2083 2396 2084
rect 2502 2088 2508 2089
rect 2502 2084 2503 2088
rect 2507 2084 2508 2088
rect 2502 2083 2508 2084
rect 2622 2088 2628 2089
rect 2622 2084 2623 2088
rect 2627 2084 2628 2088
rect 2622 2083 2628 2084
rect 2742 2088 2748 2089
rect 2742 2084 2743 2088
rect 2747 2084 2748 2088
rect 2742 2083 2748 2084
rect 2854 2088 2860 2089
rect 2854 2084 2855 2088
rect 2859 2084 2860 2088
rect 2854 2083 2860 2084
rect 2966 2088 2972 2089
rect 2966 2084 2967 2088
rect 2971 2084 2972 2088
rect 2966 2083 2972 2084
rect 3078 2088 3084 2089
rect 3078 2084 3079 2088
rect 3083 2084 3084 2088
rect 3078 2083 3084 2084
rect 3190 2088 3196 2089
rect 3190 2084 3191 2088
rect 3195 2084 3196 2088
rect 3190 2083 3196 2084
rect 3302 2088 3308 2089
rect 3302 2084 3303 2088
rect 3307 2084 3308 2088
rect 3302 2083 3308 2084
rect 3414 2088 3420 2089
rect 3414 2084 3415 2088
rect 3419 2084 3420 2088
rect 3414 2083 3420 2084
rect 3502 2088 3508 2089
rect 3502 2084 3503 2088
rect 3507 2084 3508 2088
rect 3592 2086 3594 2105
rect 3502 2083 3508 2084
rect 3590 2085 3596 2086
rect 1870 2080 1876 2081
rect 3590 2081 3591 2085
rect 3595 2081 3596 2085
rect 3590 2080 3596 2081
rect 110 2076 116 2077
rect 110 2072 111 2076
rect 115 2072 116 2076
rect 110 2071 116 2072
rect 1830 2076 1836 2077
rect 1830 2072 1831 2076
rect 1835 2072 1836 2076
rect 1830 2071 1836 2072
rect 112 2035 114 2071
rect 286 2058 292 2059
rect 286 2054 287 2058
rect 291 2054 292 2058
rect 286 2053 292 2054
rect 406 2058 412 2059
rect 406 2054 407 2058
rect 411 2054 412 2058
rect 406 2053 412 2054
rect 518 2058 524 2059
rect 518 2054 519 2058
rect 523 2054 524 2058
rect 518 2053 524 2054
rect 630 2058 636 2059
rect 630 2054 631 2058
rect 635 2054 636 2058
rect 630 2053 636 2054
rect 742 2058 748 2059
rect 742 2054 743 2058
rect 747 2054 748 2058
rect 742 2053 748 2054
rect 854 2058 860 2059
rect 854 2054 855 2058
rect 859 2054 860 2058
rect 854 2053 860 2054
rect 958 2058 964 2059
rect 958 2054 959 2058
rect 963 2054 964 2058
rect 958 2053 964 2054
rect 1054 2058 1060 2059
rect 1054 2054 1055 2058
rect 1059 2054 1060 2058
rect 1054 2053 1060 2054
rect 1150 2058 1156 2059
rect 1150 2054 1151 2058
rect 1155 2054 1156 2058
rect 1150 2053 1156 2054
rect 1246 2058 1252 2059
rect 1246 2054 1247 2058
rect 1251 2054 1252 2058
rect 1246 2053 1252 2054
rect 1350 2058 1356 2059
rect 1350 2054 1351 2058
rect 1355 2054 1356 2058
rect 1350 2053 1356 2054
rect 288 2035 290 2053
rect 408 2035 410 2053
rect 520 2035 522 2053
rect 632 2035 634 2053
rect 744 2035 746 2053
rect 856 2035 858 2053
rect 960 2035 962 2053
rect 1056 2035 1058 2053
rect 1152 2035 1154 2053
rect 1248 2035 1250 2053
rect 1352 2035 1354 2053
rect 1832 2035 1834 2071
rect 1870 2068 1876 2069
rect 1870 2064 1871 2068
rect 1875 2064 1876 2068
rect 1870 2063 1876 2064
rect 3590 2068 3596 2069
rect 3590 2064 3591 2068
rect 3595 2064 3596 2068
rect 3590 2063 3596 2064
rect 111 2034 115 2035
rect 111 2029 115 2030
rect 183 2034 187 2035
rect 183 2029 187 2030
rect 287 2034 291 2035
rect 287 2029 291 2030
rect 327 2034 331 2035
rect 327 2029 331 2030
rect 407 2034 411 2035
rect 407 2029 411 2030
rect 471 2034 475 2035
rect 471 2029 475 2030
rect 519 2034 523 2035
rect 519 2029 523 2030
rect 623 2034 627 2035
rect 623 2029 627 2030
rect 631 2034 635 2035
rect 631 2029 635 2030
rect 743 2034 747 2035
rect 743 2029 747 2030
rect 767 2034 771 2035
rect 767 2029 771 2030
rect 855 2034 859 2035
rect 855 2029 859 2030
rect 911 2034 915 2035
rect 911 2029 915 2030
rect 959 2034 963 2035
rect 959 2029 963 2030
rect 1047 2034 1051 2035
rect 1047 2029 1051 2030
rect 1055 2034 1059 2035
rect 1055 2029 1059 2030
rect 1151 2034 1155 2035
rect 1151 2029 1155 2030
rect 1183 2034 1187 2035
rect 1183 2029 1187 2030
rect 1247 2034 1251 2035
rect 1247 2029 1251 2030
rect 1319 2034 1323 2035
rect 1319 2029 1323 2030
rect 1351 2034 1355 2035
rect 1351 2029 1355 2030
rect 1463 2034 1467 2035
rect 1463 2029 1467 2030
rect 1831 2034 1835 2035
rect 1872 2031 1874 2063
rect 2294 2050 2300 2051
rect 2294 2046 2295 2050
rect 2299 2046 2300 2050
rect 2294 2045 2300 2046
rect 2398 2050 2404 2051
rect 2398 2046 2399 2050
rect 2403 2046 2404 2050
rect 2398 2045 2404 2046
rect 2510 2050 2516 2051
rect 2510 2046 2511 2050
rect 2515 2046 2516 2050
rect 2510 2045 2516 2046
rect 2630 2050 2636 2051
rect 2630 2046 2631 2050
rect 2635 2046 2636 2050
rect 2630 2045 2636 2046
rect 2750 2050 2756 2051
rect 2750 2046 2751 2050
rect 2755 2046 2756 2050
rect 2750 2045 2756 2046
rect 2862 2050 2868 2051
rect 2862 2046 2863 2050
rect 2867 2046 2868 2050
rect 2862 2045 2868 2046
rect 2974 2050 2980 2051
rect 2974 2046 2975 2050
rect 2979 2046 2980 2050
rect 2974 2045 2980 2046
rect 3086 2050 3092 2051
rect 3086 2046 3087 2050
rect 3091 2046 3092 2050
rect 3086 2045 3092 2046
rect 3198 2050 3204 2051
rect 3198 2046 3199 2050
rect 3203 2046 3204 2050
rect 3198 2045 3204 2046
rect 3310 2050 3316 2051
rect 3310 2046 3311 2050
rect 3315 2046 3316 2050
rect 3310 2045 3316 2046
rect 3422 2050 3428 2051
rect 3422 2046 3423 2050
rect 3427 2046 3428 2050
rect 3422 2045 3428 2046
rect 3510 2050 3516 2051
rect 3510 2046 3511 2050
rect 3515 2046 3516 2050
rect 3510 2045 3516 2046
rect 2296 2031 2298 2045
rect 2400 2031 2402 2045
rect 2512 2031 2514 2045
rect 2632 2031 2634 2045
rect 2752 2031 2754 2045
rect 2864 2031 2866 2045
rect 2976 2031 2978 2045
rect 3088 2031 3090 2045
rect 3200 2031 3202 2045
rect 3312 2031 3314 2045
rect 3424 2031 3426 2045
rect 3512 2031 3514 2045
rect 3592 2031 3594 2063
rect 1831 2029 1835 2030
rect 1871 2030 1875 2031
rect 112 2001 114 2029
rect 184 2019 186 2029
rect 328 2019 330 2029
rect 472 2019 474 2029
rect 624 2019 626 2029
rect 768 2019 770 2029
rect 912 2019 914 2029
rect 1048 2019 1050 2029
rect 1184 2019 1186 2029
rect 1320 2019 1322 2029
rect 1464 2019 1466 2029
rect 182 2018 188 2019
rect 182 2014 183 2018
rect 187 2014 188 2018
rect 182 2013 188 2014
rect 326 2018 332 2019
rect 326 2014 327 2018
rect 331 2014 332 2018
rect 326 2013 332 2014
rect 470 2018 476 2019
rect 470 2014 471 2018
rect 475 2014 476 2018
rect 470 2013 476 2014
rect 622 2018 628 2019
rect 622 2014 623 2018
rect 627 2014 628 2018
rect 622 2013 628 2014
rect 766 2018 772 2019
rect 766 2014 767 2018
rect 771 2014 772 2018
rect 766 2013 772 2014
rect 910 2018 916 2019
rect 910 2014 911 2018
rect 915 2014 916 2018
rect 910 2013 916 2014
rect 1046 2018 1052 2019
rect 1046 2014 1047 2018
rect 1051 2014 1052 2018
rect 1046 2013 1052 2014
rect 1182 2018 1188 2019
rect 1182 2014 1183 2018
rect 1187 2014 1188 2018
rect 1182 2013 1188 2014
rect 1318 2018 1324 2019
rect 1318 2014 1319 2018
rect 1323 2014 1324 2018
rect 1318 2013 1324 2014
rect 1462 2018 1468 2019
rect 1462 2014 1463 2018
rect 1467 2014 1468 2018
rect 1462 2013 1468 2014
rect 1832 2001 1834 2029
rect 1871 2025 1875 2026
rect 2183 2030 2187 2031
rect 2183 2025 2187 2026
rect 2271 2030 2275 2031
rect 2271 2025 2275 2026
rect 2295 2030 2299 2031
rect 2295 2025 2299 2026
rect 2367 2030 2371 2031
rect 2367 2025 2371 2026
rect 2399 2030 2403 2031
rect 2399 2025 2403 2026
rect 2463 2030 2467 2031
rect 2463 2025 2467 2026
rect 2511 2030 2515 2031
rect 2511 2025 2515 2026
rect 2567 2030 2571 2031
rect 2567 2025 2571 2026
rect 2631 2030 2635 2031
rect 2631 2025 2635 2026
rect 2671 2030 2675 2031
rect 2671 2025 2675 2026
rect 2751 2030 2755 2031
rect 2751 2025 2755 2026
rect 2775 2030 2779 2031
rect 2775 2025 2779 2026
rect 2863 2030 2867 2031
rect 2863 2025 2867 2026
rect 2879 2030 2883 2031
rect 2879 2025 2883 2026
rect 2975 2030 2979 2031
rect 2975 2025 2979 2026
rect 2983 2030 2987 2031
rect 2983 2025 2987 2026
rect 3087 2030 3091 2031
rect 3087 2025 3091 2026
rect 3191 2030 3195 2031
rect 3191 2025 3195 2026
rect 3199 2030 3203 2031
rect 3199 2025 3203 2026
rect 3311 2030 3315 2031
rect 3311 2025 3315 2026
rect 3423 2030 3427 2031
rect 3423 2025 3427 2026
rect 3511 2030 3515 2031
rect 3511 2025 3515 2026
rect 3591 2030 3595 2031
rect 3591 2025 3595 2026
rect 110 2000 116 2001
rect 110 1996 111 2000
rect 115 1996 116 2000
rect 110 1995 116 1996
rect 1830 2000 1836 2001
rect 1830 1996 1831 2000
rect 1835 1996 1836 2000
rect 1872 1997 1874 2025
rect 2184 2015 2186 2025
rect 2272 2015 2274 2025
rect 2368 2015 2370 2025
rect 2464 2015 2466 2025
rect 2568 2015 2570 2025
rect 2672 2015 2674 2025
rect 2776 2015 2778 2025
rect 2880 2015 2882 2025
rect 2984 2015 2986 2025
rect 3088 2015 3090 2025
rect 3192 2015 3194 2025
rect 2182 2014 2188 2015
rect 2182 2010 2183 2014
rect 2187 2010 2188 2014
rect 2182 2009 2188 2010
rect 2270 2014 2276 2015
rect 2270 2010 2271 2014
rect 2275 2010 2276 2014
rect 2270 2009 2276 2010
rect 2366 2014 2372 2015
rect 2366 2010 2367 2014
rect 2371 2010 2372 2014
rect 2366 2009 2372 2010
rect 2462 2014 2468 2015
rect 2462 2010 2463 2014
rect 2467 2010 2468 2014
rect 2462 2009 2468 2010
rect 2566 2014 2572 2015
rect 2566 2010 2567 2014
rect 2571 2010 2572 2014
rect 2566 2009 2572 2010
rect 2670 2014 2676 2015
rect 2670 2010 2671 2014
rect 2675 2010 2676 2014
rect 2670 2009 2676 2010
rect 2774 2014 2780 2015
rect 2774 2010 2775 2014
rect 2779 2010 2780 2014
rect 2774 2009 2780 2010
rect 2878 2014 2884 2015
rect 2878 2010 2879 2014
rect 2883 2010 2884 2014
rect 2878 2009 2884 2010
rect 2982 2014 2988 2015
rect 2982 2010 2983 2014
rect 2987 2010 2988 2014
rect 2982 2009 2988 2010
rect 3086 2014 3092 2015
rect 3086 2010 3087 2014
rect 3091 2010 3092 2014
rect 3086 2009 3092 2010
rect 3190 2014 3196 2015
rect 3190 2010 3191 2014
rect 3195 2010 3196 2014
rect 3190 2009 3196 2010
rect 3592 1997 3594 2025
rect 1830 1995 1836 1996
rect 1870 1996 1876 1997
rect 1870 1992 1871 1996
rect 1875 1992 1876 1996
rect 1870 1991 1876 1992
rect 3590 1996 3596 1997
rect 3590 1992 3591 1996
rect 3595 1992 3596 1996
rect 3590 1991 3596 1992
rect 110 1983 116 1984
rect 110 1979 111 1983
rect 115 1979 116 1983
rect 1830 1983 1836 1984
rect 110 1978 116 1979
rect 174 1980 180 1981
rect 112 1959 114 1978
rect 174 1976 175 1980
rect 179 1976 180 1980
rect 174 1975 180 1976
rect 318 1980 324 1981
rect 318 1976 319 1980
rect 323 1976 324 1980
rect 318 1975 324 1976
rect 462 1980 468 1981
rect 462 1976 463 1980
rect 467 1976 468 1980
rect 462 1975 468 1976
rect 614 1980 620 1981
rect 614 1976 615 1980
rect 619 1976 620 1980
rect 614 1975 620 1976
rect 758 1980 764 1981
rect 758 1976 759 1980
rect 763 1976 764 1980
rect 758 1975 764 1976
rect 902 1980 908 1981
rect 902 1976 903 1980
rect 907 1976 908 1980
rect 902 1975 908 1976
rect 1038 1980 1044 1981
rect 1038 1976 1039 1980
rect 1043 1976 1044 1980
rect 1038 1975 1044 1976
rect 1174 1980 1180 1981
rect 1174 1976 1175 1980
rect 1179 1976 1180 1980
rect 1174 1975 1180 1976
rect 1310 1980 1316 1981
rect 1310 1976 1311 1980
rect 1315 1976 1316 1980
rect 1310 1975 1316 1976
rect 1454 1980 1460 1981
rect 1454 1976 1455 1980
rect 1459 1976 1460 1980
rect 1830 1979 1831 1983
rect 1835 1979 1836 1983
rect 1830 1978 1836 1979
rect 1870 1979 1876 1980
rect 1454 1975 1460 1976
rect 176 1959 178 1975
rect 320 1959 322 1975
rect 464 1959 466 1975
rect 616 1959 618 1975
rect 760 1959 762 1975
rect 904 1959 906 1975
rect 1040 1959 1042 1975
rect 1176 1959 1178 1975
rect 1312 1959 1314 1975
rect 1456 1959 1458 1975
rect 1832 1959 1834 1978
rect 1870 1975 1871 1979
rect 1875 1975 1876 1979
rect 3590 1979 3596 1980
rect 1870 1974 1876 1975
rect 2174 1976 2180 1977
rect 111 1958 115 1959
rect 111 1953 115 1954
rect 135 1958 139 1959
rect 135 1953 139 1954
rect 175 1958 179 1959
rect 175 1953 179 1954
rect 295 1958 299 1959
rect 295 1953 299 1954
rect 319 1958 323 1959
rect 319 1953 323 1954
rect 463 1958 467 1959
rect 463 1953 467 1954
rect 615 1958 619 1959
rect 615 1953 619 1954
rect 631 1958 635 1959
rect 631 1953 635 1954
rect 759 1958 763 1959
rect 759 1953 763 1954
rect 799 1958 803 1959
rect 799 1953 803 1954
rect 903 1958 907 1959
rect 903 1953 907 1954
rect 951 1958 955 1959
rect 951 1953 955 1954
rect 1039 1958 1043 1959
rect 1039 1953 1043 1954
rect 1095 1958 1099 1959
rect 1095 1953 1099 1954
rect 1175 1958 1179 1959
rect 1175 1953 1179 1954
rect 1231 1958 1235 1959
rect 1231 1953 1235 1954
rect 1311 1958 1315 1959
rect 1311 1953 1315 1954
rect 1359 1958 1363 1959
rect 1359 1953 1363 1954
rect 1455 1958 1459 1959
rect 1455 1953 1459 1954
rect 1487 1958 1491 1959
rect 1487 1953 1491 1954
rect 1623 1958 1627 1959
rect 1623 1953 1627 1954
rect 1831 1958 1835 1959
rect 1831 1953 1835 1954
rect 112 1934 114 1953
rect 136 1937 138 1953
rect 296 1937 298 1953
rect 464 1937 466 1953
rect 632 1937 634 1953
rect 800 1937 802 1953
rect 952 1937 954 1953
rect 1096 1937 1098 1953
rect 1232 1937 1234 1953
rect 1360 1937 1362 1953
rect 1488 1937 1490 1953
rect 1624 1937 1626 1953
rect 134 1936 140 1937
rect 110 1933 116 1934
rect 110 1929 111 1933
rect 115 1929 116 1933
rect 134 1932 135 1936
rect 139 1932 140 1936
rect 134 1931 140 1932
rect 294 1936 300 1937
rect 294 1932 295 1936
rect 299 1932 300 1936
rect 294 1931 300 1932
rect 462 1936 468 1937
rect 462 1932 463 1936
rect 467 1932 468 1936
rect 462 1931 468 1932
rect 630 1936 636 1937
rect 630 1932 631 1936
rect 635 1932 636 1936
rect 630 1931 636 1932
rect 798 1936 804 1937
rect 798 1932 799 1936
rect 803 1932 804 1936
rect 798 1931 804 1932
rect 950 1936 956 1937
rect 950 1932 951 1936
rect 955 1932 956 1936
rect 950 1931 956 1932
rect 1094 1936 1100 1937
rect 1094 1932 1095 1936
rect 1099 1932 1100 1936
rect 1094 1931 1100 1932
rect 1230 1936 1236 1937
rect 1230 1932 1231 1936
rect 1235 1932 1236 1936
rect 1230 1931 1236 1932
rect 1358 1936 1364 1937
rect 1358 1932 1359 1936
rect 1363 1932 1364 1936
rect 1358 1931 1364 1932
rect 1486 1936 1492 1937
rect 1486 1932 1487 1936
rect 1491 1932 1492 1936
rect 1486 1931 1492 1932
rect 1622 1936 1628 1937
rect 1622 1932 1623 1936
rect 1627 1932 1628 1936
rect 1832 1934 1834 1953
rect 1872 1951 1874 1974
rect 2174 1972 2175 1976
rect 2179 1972 2180 1976
rect 2174 1971 2180 1972
rect 2262 1976 2268 1977
rect 2262 1972 2263 1976
rect 2267 1972 2268 1976
rect 2262 1971 2268 1972
rect 2358 1976 2364 1977
rect 2358 1972 2359 1976
rect 2363 1972 2364 1976
rect 2358 1971 2364 1972
rect 2454 1976 2460 1977
rect 2454 1972 2455 1976
rect 2459 1972 2460 1976
rect 2454 1971 2460 1972
rect 2558 1976 2564 1977
rect 2558 1972 2559 1976
rect 2563 1972 2564 1976
rect 2558 1971 2564 1972
rect 2662 1976 2668 1977
rect 2662 1972 2663 1976
rect 2667 1972 2668 1976
rect 2662 1971 2668 1972
rect 2766 1976 2772 1977
rect 2766 1972 2767 1976
rect 2771 1972 2772 1976
rect 2766 1971 2772 1972
rect 2870 1976 2876 1977
rect 2870 1972 2871 1976
rect 2875 1972 2876 1976
rect 2870 1971 2876 1972
rect 2974 1976 2980 1977
rect 2974 1972 2975 1976
rect 2979 1972 2980 1976
rect 2974 1971 2980 1972
rect 3078 1976 3084 1977
rect 3078 1972 3079 1976
rect 3083 1972 3084 1976
rect 3078 1971 3084 1972
rect 3182 1976 3188 1977
rect 3182 1972 3183 1976
rect 3187 1972 3188 1976
rect 3590 1975 3591 1979
rect 3595 1975 3596 1979
rect 3590 1974 3596 1975
rect 3182 1971 3188 1972
rect 2176 1951 2178 1971
rect 2264 1951 2266 1971
rect 2360 1951 2362 1971
rect 2456 1951 2458 1971
rect 2560 1951 2562 1971
rect 2664 1951 2666 1971
rect 2768 1951 2770 1971
rect 2872 1951 2874 1971
rect 2976 1951 2978 1971
rect 3080 1951 3082 1971
rect 3184 1951 3186 1971
rect 3592 1951 3594 1974
rect 1871 1950 1875 1951
rect 1871 1945 1875 1946
rect 1943 1950 1947 1951
rect 1943 1945 1947 1946
rect 2055 1950 2059 1951
rect 2055 1945 2059 1946
rect 2167 1950 2171 1951
rect 2167 1945 2171 1946
rect 2175 1950 2179 1951
rect 2175 1945 2179 1946
rect 2263 1950 2267 1951
rect 2263 1945 2267 1946
rect 2287 1950 2291 1951
rect 2287 1945 2291 1946
rect 2359 1950 2363 1951
rect 2359 1945 2363 1946
rect 2407 1950 2411 1951
rect 2407 1945 2411 1946
rect 2455 1950 2459 1951
rect 2455 1945 2459 1946
rect 2527 1950 2531 1951
rect 2527 1945 2531 1946
rect 2559 1950 2563 1951
rect 2559 1945 2563 1946
rect 2647 1950 2651 1951
rect 2647 1945 2651 1946
rect 2663 1950 2667 1951
rect 2663 1945 2667 1946
rect 2767 1950 2771 1951
rect 2767 1945 2771 1946
rect 2775 1950 2779 1951
rect 2775 1945 2779 1946
rect 2871 1950 2875 1951
rect 2871 1945 2875 1946
rect 2911 1950 2915 1951
rect 2911 1945 2915 1946
rect 2975 1950 2979 1951
rect 2975 1945 2979 1946
rect 3055 1950 3059 1951
rect 3055 1945 3059 1946
rect 3079 1950 3083 1951
rect 3079 1945 3083 1946
rect 3183 1950 3187 1951
rect 3183 1945 3187 1946
rect 3207 1950 3211 1951
rect 3207 1945 3211 1946
rect 3367 1950 3371 1951
rect 3367 1945 3371 1946
rect 3503 1950 3507 1951
rect 3503 1945 3507 1946
rect 3591 1950 3595 1951
rect 3591 1945 3595 1946
rect 1622 1931 1628 1932
rect 1830 1933 1836 1934
rect 110 1928 116 1929
rect 1830 1929 1831 1933
rect 1835 1929 1836 1933
rect 1830 1928 1836 1929
rect 1872 1926 1874 1945
rect 1944 1929 1946 1945
rect 2056 1929 2058 1945
rect 2168 1929 2170 1945
rect 2288 1929 2290 1945
rect 2408 1929 2410 1945
rect 2528 1929 2530 1945
rect 2648 1929 2650 1945
rect 2776 1929 2778 1945
rect 2912 1929 2914 1945
rect 3056 1929 3058 1945
rect 3208 1929 3210 1945
rect 3368 1929 3370 1945
rect 3504 1929 3506 1945
rect 1942 1928 1948 1929
rect 1870 1925 1876 1926
rect 1870 1921 1871 1925
rect 1875 1921 1876 1925
rect 1942 1924 1943 1928
rect 1947 1924 1948 1928
rect 1942 1923 1948 1924
rect 2054 1928 2060 1929
rect 2054 1924 2055 1928
rect 2059 1924 2060 1928
rect 2054 1923 2060 1924
rect 2166 1928 2172 1929
rect 2166 1924 2167 1928
rect 2171 1924 2172 1928
rect 2166 1923 2172 1924
rect 2286 1928 2292 1929
rect 2286 1924 2287 1928
rect 2291 1924 2292 1928
rect 2286 1923 2292 1924
rect 2406 1928 2412 1929
rect 2406 1924 2407 1928
rect 2411 1924 2412 1928
rect 2406 1923 2412 1924
rect 2526 1928 2532 1929
rect 2526 1924 2527 1928
rect 2531 1924 2532 1928
rect 2526 1923 2532 1924
rect 2646 1928 2652 1929
rect 2646 1924 2647 1928
rect 2651 1924 2652 1928
rect 2646 1923 2652 1924
rect 2774 1928 2780 1929
rect 2774 1924 2775 1928
rect 2779 1924 2780 1928
rect 2774 1923 2780 1924
rect 2910 1928 2916 1929
rect 2910 1924 2911 1928
rect 2915 1924 2916 1928
rect 2910 1923 2916 1924
rect 3054 1928 3060 1929
rect 3054 1924 3055 1928
rect 3059 1924 3060 1928
rect 3054 1923 3060 1924
rect 3206 1928 3212 1929
rect 3206 1924 3207 1928
rect 3211 1924 3212 1928
rect 3206 1923 3212 1924
rect 3366 1928 3372 1929
rect 3366 1924 3367 1928
rect 3371 1924 3372 1928
rect 3366 1923 3372 1924
rect 3502 1928 3508 1929
rect 3502 1924 3503 1928
rect 3507 1924 3508 1928
rect 3592 1926 3594 1945
rect 3502 1923 3508 1924
rect 3590 1925 3596 1926
rect 1870 1920 1876 1921
rect 3590 1921 3591 1925
rect 3595 1921 3596 1925
rect 3590 1920 3596 1921
rect 110 1916 116 1917
rect 110 1912 111 1916
rect 115 1912 116 1916
rect 110 1911 116 1912
rect 1830 1916 1836 1917
rect 1830 1912 1831 1916
rect 1835 1912 1836 1916
rect 1830 1911 1836 1912
rect 112 1875 114 1911
rect 142 1898 148 1899
rect 142 1894 143 1898
rect 147 1894 148 1898
rect 142 1893 148 1894
rect 302 1898 308 1899
rect 302 1894 303 1898
rect 307 1894 308 1898
rect 302 1893 308 1894
rect 470 1898 476 1899
rect 470 1894 471 1898
rect 475 1894 476 1898
rect 470 1893 476 1894
rect 638 1898 644 1899
rect 638 1894 639 1898
rect 643 1894 644 1898
rect 638 1893 644 1894
rect 806 1898 812 1899
rect 806 1894 807 1898
rect 811 1894 812 1898
rect 806 1893 812 1894
rect 958 1898 964 1899
rect 958 1894 959 1898
rect 963 1894 964 1898
rect 958 1893 964 1894
rect 1102 1898 1108 1899
rect 1102 1894 1103 1898
rect 1107 1894 1108 1898
rect 1102 1893 1108 1894
rect 1238 1898 1244 1899
rect 1238 1894 1239 1898
rect 1243 1894 1244 1898
rect 1238 1893 1244 1894
rect 1366 1898 1372 1899
rect 1366 1894 1367 1898
rect 1371 1894 1372 1898
rect 1366 1893 1372 1894
rect 1494 1898 1500 1899
rect 1494 1894 1495 1898
rect 1499 1894 1500 1898
rect 1494 1893 1500 1894
rect 1630 1898 1636 1899
rect 1630 1894 1631 1898
rect 1635 1894 1636 1898
rect 1630 1893 1636 1894
rect 144 1875 146 1893
rect 304 1875 306 1893
rect 472 1875 474 1893
rect 640 1875 642 1893
rect 808 1875 810 1893
rect 960 1875 962 1893
rect 1104 1875 1106 1893
rect 1240 1875 1242 1893
rect 1368 1875 1370 1893
rect 1496 1875 1498 1893
rect 1632 1875 1634 1893
rect 1832 1875 1834 1911
rect 1870 1908 1876 1909
rect 1870 1904 1871 1908
rect 1875 1904 1876 1908
rect 1870 1903 1876 1904
rect 3590 1908 3596 1909
rect 3590 1904 3591 1908
rect 3595 1904 3596 1908
rect 3590 1903 3596 1904
rect 111 1874 115 1875
rect 111 1869 115 1870
rect 143 1874 147 1875
rect 143 1869 147 1870
rect 303 1874 307 1875
rect 303 1869 307 1870
rect 319 1874 323 1875
rect 319 1869 323 1870
rect 471 1874 475 1875
rect 471 1869 475 1870
rect 519 1874 523 1875
rect 519 1869 523 1870
rect 639 1874 643 1875
rect 639 1869 643 1870
rect 711 1874 715 1875
rect 711 1869 715 1870
rect 807 1874 811 1875
rect 807 1869 811 1870
rect 887 1874 891 1875
rect 887 1869 891 1870
rect 959 1874 963 1875
rect 959 1869 963 1870
rect 1055 1874 1059 1875
rect 1055 1869 1059 1870
rect 1103 1874 1107 1875
rect 1103 1869 1107 1870
rect 1207 1874 1211 1875
rect 1207 1869 1211 1870
rect 1239 1874 1243 1875
rect 1239 1869 1243 1870
rect 1343 1874 1347 1875
rect 1343 1869 1347 1870
rect 1367 1874 1371 1875
rect 1367 1869 1371 1870
rect 1471 1874 1475 1875
rect 1471 1869 1475 1870
rect 1495 1874 1499 1875
rect 1495 1869 1499 1870
rect 1599 1874 1603 1875
rect 1599 1869 1603 1870
rect 1631 1874 1635 1875
rect 1631 1869 1635 1870
rect 1727 1874 1731 1875
rect 1727 1869 1731 1870
rect 1831 1874 1835 1875
rect 1872 1871 1874 1903
rect 1950 1890 1956 1891
rect 1950 1886 1951 1890
rect 1955 1886 1956 1890
rect 1950 1885 1956 1886
rect 2062 1890 2068 1891
rect 2062 1886 2063 1890
rect 2067 1886 2068 1890
rect 2062 1885 2068 1886
rect 2174 1890 2180 1891
rect 2174 1886 2175 1890
rect 2179 1886 2180 1890
rect 2174 1885 2180 1886
rect 2294 1890 2300 1891
rect 2294 1886 2295 1890
rect 2299 1886 2300 1890
rect 2294 1885 2300 1886
rect 2414 1890 2420 1891
rect 2414 1886 2415 1890
rect 2419 1886 2420 1890
rect 2414 1885 2420 1886
rect 2534 1890 2540 1891
rect 2534 1886 2535 1890
rect 2539 1886 2540 1890
rect 2534 1885 2540 1886
rect 2654 1890 2660 1891
rect 2654 1886 2655 1890
rect 2659 1886 2660 1890
rect 2654 1885 2660 1886
rect 2782 1890 2788 1891
rect 2782 1886 2783 1890
rect 2787 1886 2788 1890
rect 2782 1885 2788 1886
rect 2918 1890 2924 1891
rect 2918 1886 2919 1890
rect 2923 1886 2924 1890
rect 2918 1885 2924 1886
rect 3062 1890 3068 1891
rect 3062 1886 3063 1890
rect 3067 1886 3068 1890
rect 3062 1885 3068 1886
rect 3214 1890 3220 1891
rect 3214 1886 3215 1890
rect 3219 1886 3220 1890
rect 3214 1885 3220 1886
rect 3374 1890 3380 1891
rect 3374 1886 3375 1890
rect 3379 1886 3380 1890
rect 3374 1885 3380 1886
rect 3510 1890 3516 1891
rect 3510 1886 3511 1890
rect 3515 1886 3516 1890
rect 3510 1885 3516 1886
rect 1952 1871 1954 1885
rect 2064 1871 2066 1885
rect 2176 1871 2178 1885
rect 2296 1871 2298 1885
rect 2416 1871 2418 1885
rect 2536 1871 2538 1885
rect 2656 1871 2658 1885
rect 2784 1871 2786 1885
rect 2920 1871 2922 1885
rect 3064 1871 3066 1885
rect 3216 1871 3218 1885
rect 3376 1871 3378 1885
rect 3512 1871 3514 1885
rect 3592 1871 3594 1903
rect 1831 1869 1835 1870
rect 1871 1870 1875 1871
rect 112 1841 114 1869
rect 144 1859 146 1869
rect 320 1859 322 1869
rect 520 1859 522 1869
rect 712 1859 714 1869
rect 888 1859 890 1869
rect 1056 1859 1058 1869
rect 1208 1859 1210 1869
rect 1344 1859 1346 1869
rect 1472 1859 1474 1869
rect 1600 1859 1602 1869
rect 1728 1859 1730 1869
rect 142 1858 148 1859
rect 142 1854 143 1858
rect 147 1854 148 1858
rect 142 1853 148 1854
rect 318 1858 324 1859
rect 318 1854 319 1858
rect 323 1854 324 1858
rect 318 1853 324 1854
rect 518 1858 524 1859
rect 518 1854 519 1858
rect 523 1854 524 1858
rect 518 1853 524 1854
rect 710 1858 716 1859
rect 710 1854 711 1858
rect 715 1854 716 1858
rect 710 1853 716 1854
rect 886 1858 892 1859
rect 886 1854 887 1858
rect 891 1854 892 1858
rect 886 1853 892 1854
rect 1054 1858 1060 1859
rect 1054 1854 1055 1858
rect 1059 1854 1060 1858
rect 1054 1853 1060 1854
rect 1206 1858 1212 1859
rect 1206 1854 1207 1858
rect 1211 1854 1212 1858
rect 1206 1853 1212 1854
rect 1342 1858 1348 1859
rect 1342 1854 1343 1858
rect 1347 1854 1348 1858
rect 1342 1853 1348 1854
rect 1470 1858 1476 1859
rect 1470 1854 1471 1858
rect 1475 1854 1476 1858
rect 1470 1853 1476 1854
rect 1598 1858 1604 1859
rect 1598 1854 1599 1858
rect 1603 1854 1604 1858
rect 1598 1853 1604 1854
rect 1726 1858 1732 1859
rect 1726 1854 1727 1858
rect 1731 1854 1732 1858
rect 1726 1853 1732 1854
rect 1832 1841 1834 1869
rect 1871 1865 1875 1866
rect 1903 1870 1907 1871
rect 1903 1865 1907 1866
rect 1951 1870 1955 1871
rect 1951 1865 1955 1866
rect 1983 1870 1987 1871
rect 1983 1865 1987 1866
rect 2063 1870 2067 1871
rect 2063 1865 2067 1866
rect 2095 1870 2099 1871
rect 2095 1865 2099 1866
rect 2175 1870 2179 1871
rect 2175 1865 2179 1866
rect 2207 1870 2211 1871
rect 2207 1865 2211 1866
rect 2295 1870 2299 1871
rect 2295 1865 2299 1866
rect 2327 1870 2331 1871
rect 2327 1865 2331 1866
rect 2415 1870 2419 1871
rect 2415 1865 2419 1866
rect 2463 1870 2467 1871
rect 2463 1865 2467 1866
rect 2535 1870 2539 1871
rect 2535 1865 2539 1866
rect 2631 1870 2635 1871
rect 2631 1865 2635 1866
rect 2655 1870 2659 1871
rect 2655 1865 2659 1866
rect 2783 1870 2787 1871
rect 2783 1865 2787 1866
rect 2831 1870 2835 1871
rect 2831 1865 2835 1866
rect 2919 1870 2923 1871
rect 2919 1865 2923 1866
rect 3055 1870 3059 1871
rect 3055 1865 3059 1866
rect 3063 1870 3067 1871
rect 3063 1865 3067 1866
rect 3215 1870 3219 1871
rect 3215 1865 3219 1866
rect 3295 1870 3299 1871
rect 3295 1865 3299 1866
rect 3375 1870 3379 1871
rect 3375 1865 3379 1866
rect 3511 1870 3515 1871
rect 3511 1865 3515 1866
rect 3591 1870 3595 1871
rect 3591 1865 3595 1866
rect 110 1840 116 1841
rect 110 1836 111 1840
rect 115 1836 116 1840
rect 110 1835 116 1836
rect 1830 1840 1836 1841
rect 1830 1836 1831 1840
rect 1835 1836 1836 1840
rect 1872 1837 1874 1865
rect 1904 1855 1906 1865
rect 1984 1855 1986 1865
rect 2096 1855 2098 1865
rect 2208 1855 2210 1865
rect 2328 1855 2330 1865
rect 2464 1855 2466 1865
rect 2632 1855 2634 1865
rect 2832 1855 2834 1865
rect 3056 1855 3058 1865
rect 3296 1855 3298 1865
rect 3512 1855 3514 1865
rect 1902 1854 1908 1855
rect 1902 1850 1903 1854
rect 1907 1850 1908 1854
rect 1902 1849 1908 1850
rect 1982 1854 1988 1855
rect 1982 1850 1983 1854
rect 1987 1850 1988 1854
rect 1982 1849 1988 1850
rect 2094 1854 2100 1855
rect 2094 1850 2095 1854
rect 2099 1850 2100 1854
rect 2094 1849 2100 1850
rect 2206 1854 2212 1855
rect 2206 1850 2207 1854
rect 2211 1850 2212 1854
rect 2206 1849 2212 1850
rect 2326 1854 2332 1855
rect 2326 1850 2327 1854
rect 2331 1850 2332 1854
rect 2326 1849 2332 1850
rect 2462 1854 2468 1855
rect 2462 1850 2463 1854
rect 2467 1850 2468 1854
rect 2462 1849 2468 1850
rect 2630 1854 2636 1855
rect 2630 1850 2631 1854
rect 2635 1850 2636 1854
rect 2630 1849 2636 1850
rect 2830 1854 2836 1855
rect 2830 1850 2831 1854
rect 2835 1850 2836 1854
rect 2830 1849 2836 1850
rect 3054 1854 3060 1855
rect 3054 1850 3055 1854
rect 3059 1850 3060 1854
rect 3054 1849 3060 1850
rect 3294 1854 3300 1855
rect 3294 1850 3295 1854
rect 3299 1850 3300 1854
rect 3294 1849 3300 1850
rect 3510 1854 3516 1855
rect 3510 1850 3511 1854
rect 3515 1850 3516 1854
rect 3510 1849 3516 1850
rect 3592 1837 3594 1865
rect 1830 1835 1836 1836
rect 1870 1836 1876 1837
rect 1870 1832 1871 1836
rect 1875 1832 1876 1836
rect 1870 1831 1876 1832
rect 3590 1836 3596 1837
rect 3590 1832 3591 1836
rect 3595 1832 3596 1836
rect 3590 1831 3596 1832
rect 110 1823 116 1824
rect 110 1819 111 1823
rect 115 1819 116 1823
rect 1830 1823 1836 1824
rect 110 1818 116 1819
rect 134 1820 140 1821
rect 112 1799 114 1818
rect 134 1816 135 1820
rect 139 1816 140 1820
rect 134 1815 140 1816
rect 310 1820 316 1821
rect 310 1816 311 1820
rect 315 1816 316 1820
rect 310 1815 316 1816
rect 510 1820 516 1821
rect 510 1816 511 1820
rect 515 1816 516 1820
rect 510 1815 516 1816
rect 702 1820 708 1821
rect 702 1816 703 1820
rect 707 1816 708 1820
rect 702 1815 708 1816
rect 878 1820 884 1821
rect 878 1816 879 1820
rect 883 1816 884 1820
rect 878 1815 884 1816
rect 1046 1820 1052 1821
rect 1046 1816 1047 1820
rect 1051 1816 1052 1820
rect 1046 1815 1052 1816
rect 1198 1820 1204 1821
rect 1198 1816 1199 1820
rect 1203 1816 1204 1820
rect 1198 1815 1204 1816
rect 1334 1820 1340 1821
rect 1334 1816 1335 1820
rect 1339 1816 1340 1820
rect 1334 1815 1340 1816
rect 1462 1820 1468 1821
rect 1462 1816 1463 1820
rect 1467 1816 1468 1820
rect 1462 1815 1468 1816
rect 1590 1820 1596 1821
rect 1590 1816 1591 1820
rect 1595 1816 1596 1820
rect 1590 1815 1596 1816
rect 1718 1820 1724 1821
rect 1718 1816 1719 1820
rect 1723 1816 1724 1820
rect 1830 1819 1831 1823
rect 1835 1819 1836 1823
rect 1830 1818 1836 1819
rect 1870 1819 1876 1820
rect 1718 1815 1724 1816
rect 136 1799 138 1815
rect 312 1799 314 1815
rect 512 1799 514 1815
rect 704 1799 706 1815
rect 880 1799 882 1815
rect 1048 1799 1050 1815
rect 1200 1799 1202 1815
rect 1336 1799 1338 1815
rect 1464 1799 1466 1815
rect 1592 1799 1594 1815
rect 1720 1799 1722 1815
rect 1832 1799 1834 1818
rect 1870 1815 1871 1819
rect 1875 1815 1876 1819
rect 3590 1819 3596 1820
rect 1870 1814 1876 1815
rect 1894 1816 1900 1817
rect 111 1798 115 1799
rect 111 1793 115 1794
rect 135 1798 139 1799
rect 135 1793 139 1794
rect 311 1798 315 1799
rect 311 1793 315 1794
rect 503 1798 507 1799
rect 503 1793 507 1794
rect 511 1798 515 1799
rect 511 1793 515 1794
rect 687 1798 691 1799
rect 687 1793 691 1794
rect 703 1798 707 1799
rect 703 1793 707 1794
rect 847 1798 851 1799
rect 847 1793 851 1794
rect 879 1798 883 1799
rect 879 1793 883 1794
rect 991 1798 995 1799
rect 991 1793 995 1794
rect 1047 1798 1051 1799
rect 1047 1793 1051 1794
rect 1127 1798 1131 1799
rect 1127 1793 1131 1794
rect 1199 1798 1203 1799
rect 1199 1793 1203 1794
rect 1247 1798 1251 1799
rect 1247 1793 1251 1794
rect 1335 1798 1339 1799
rect 1335 1793 1339 1794
rect 1359 1798 1363 1799
rect 1359 1793 1363 1794
rect 1463 1798 1467 1799
rect 1463 1793 1467 1794
rect 1559 1798 1563 1799
rect 1559 1793 1563 1794
rect 1591 1798 1595 1799
rect 1591 1793 1595 1794
rect 1663 1798 1667 1799
rect 1663 1793 1667 1794
rect 1719 1798 1723 1799
rect 1719 1793 1723 1794
rect 1743 1798 1747 1799
rect 1743 1793 1747 1794
rect 1831 1798 1835 1799
rect 1831 1793 1835 1794
rect 112 1774 114 1793
rect 136 1777 138 1793
rect 312 1777 314 1793
rect 504 1777 506 1793
rect 688 1777 690 1793
rect 848 1777 850 1793
rect 992 1777 994 1793
rect 1128 1777 1130 1793
rect 1248 1777 1250 1793
rect 1360 1777 1362 1793
rect 1464 1777 1466 1793
rect 1560 1777 1562 1793
rect 1664 1777 1666 1793
rect 1744 1777 1746 1793
rect 134 1776 140 1777
rect 110 1773 116 1774
rect 110 1769 111 1773
rect 115 1769 116 1773
rect 134 1772 135 1776
rect 139 1772 140 1776
rect 134 1771 140 1772
rect 310 1776 316 1777
rect 310 1772 311 1776
rect 315 1772 316 1776
rect 310 1771 316 1772
rect 502 1776 508 1777
rect 502 1772 503 1776
rect 507 1772 508 1776
rect 502 1771 508 1772
rect 686 1776 692 1777
rect 686 1772 687 1776
rect 691 1772 692 1776
rect 686 1771 692 1772
rect 846 1776 852 1777
rect 846 1772 847 1776
rect 851 1772 852 1776
rect 846 1771 852 1772
rect 990 1776 996 1777
rect 990 1772 991 1776
rect 995 1772 996 1776
rect 990 1771 996 1772
rect 1126 1776 1132 1777
rect 1126 1772 1127 1776
rect 1131 1772 1132 1776
rect 1126 1771 1132 1772
rect 1246 1776 1252 1777
rect 1246 1772 1247 1776
rect 1251 1772 1252 1776
rect 1246 1771 1252 1772
rect 1358 1776 1364 1777
rect 1358 1772 1359 1776
rect 1363 1772 1364 1776
rect 1358 1771 1364 1772
rect 1462 1776 1468 1777
rect 1462 1772 1463 1776
rect 1467 1772 1468 1776
rect 1462 1771 1468 1772
rect 1558 1776 1564 1777
rect 1558 1772 1559 1776
rect 1563 1772 1564 1776
rect 1558 1771 1564 1772
rect 1662 1776 1668 1777
rect 1662 1772 1663 1776
rect 1667 1772 1668 1776
rect 1662 1771 1668 1772
rect 1742 1776 1748 1777
rect 1742 1772 1743 1776
rect 1747 1772 1748 1776
rect 1832 1774 1834 1793
rect 1872 1779 1874 1814
rect 1894 1812 1895 1816
rect 1899 1812 1900 1816
rect 1894 1811 1900 1812
rect 1974 1816 1980 1817
rect 1974 1812 1975 1816
rect 1979 1812 1980 1816
rect 1974 1811 1980 1812
rect 2086 1816 2092 1817
rect 2086 1812 2087 1816
rect 2091 1812 2092 1816
rect 2086 1811 2092 1812
rect 2198 1816 2204 1817
rect 2198 1812 2199 1816
rect 2203 1812 2204 1816
rect 2198 1811 2204 1812
rect 2318 1816 2324 1817
rect 2318 1812 2319 1816
rect 2323 1812 2324 1816
rect 2318 1811 2324 1812
rect 2454 1816 2460 1817
rect 2454 1812 2455 1816
rect 2459 1812 2460 1816
rect 2454 1811 2460 1812
rect 2622 1816 2628 1817
rect 2622 1812 2623 1816
rect 2627 1812 2628 1816
rect 2622 1811 2628 1812
rect 2822 1816 2828 1817
rect 2822 1812 2823 1816
rect 2827 1812 2828 1816
rect 2822 1811 2828 1812
rect 3046 1816 3052 1817
rect 3046 1812 3047 1816
rect 3051 1812 3052 1816
rect 3046 1811 3052 1812
rect 3286 1816 3292 1817
rect 3286 1812 3287 1816
rect 3291 1812 3292 1816
rect 3286 1811 3292 1812
rect 3502 1816 3508 1817
rect 3502 1812 3503 1816
rect 3507 1812 3508 1816
rect 3590 1815 3591 1819
rect 3595 1815 3596 1819
rect 3590 1814 3596 1815
rect 3502 1811 3508 1812
rect 1896 1779 1898 1811
rect 1976 1779 1978 1811
rect 2088 1779 2090 1811
rect 2200 1779 2202 1811
rect 2320 1779 2322 1811
rect 2456 1779 2458 1811
rect 2624 1779 2626 1811
rect 2824 1779 2826 1811
rect 3048 1779 3050 1811
rect 3288 1779 3290 1811
rect 3504 1779 3506 1811
rect 3592 1779 3594 1814
rect 1871 1778 1875 1779
rect 1742 1771 1748 1772
rect 1830 1773 1836 1774
rect 1871 1773 1875 1774
rect 1895 1778 1899 1779
rect 1895 1773 1899 1774
rect 1975 1778 1979 1779
rect 1975 1773 1979 1774
rect 2023 1778 2027 1779
rect 2023 1773 2027 1774
rect 2087 1778 2091 1779
rect 2087 1773 2091 1774
rect 2183 1778 2187 1779
rect 2183 1773 2187 1774
rect 2199 1778 2203 1779
rect 2199 1773 2203 1774
rect 2319 1778 2323 1779
rect 2319 1773 2323 1774
rect 2351 1778 2355 1779
rect 2351 1773 2355 1774
rect 2455 1778 2459 1779
rect 2455 1773 2459 1774
rect 2551 1778 2555 1779
rect 2551 1773 2555 1774
rect 2623 1778 2627 1779
rect 2623 1773 2627 1774
rect 2775 1778 2779 1779
rect 2775 1773 2779 1774
rect 2823 1778 2827 1779
rect 2823 1773 2827 1774
rect 3015 1778 3019 1779
rect 3015 1773 3019 1774
rect 3047 1778 3051 1779
rect 3047 1773 3051 1774
rect 3271 1778 3275 1779
rect 3271 1773 3275 1774
rect 3287 1778 3291 1779
rect 3287 1773 3291 1774
rect 3503 1778 3507 1779
rect 3503 1773 3507 1774
rect 3591 1778 3595 1779
rect 3591 1773 3595 1774
rect 110 1768 116 1769
rect 1830 1769 1831 1773
rect 1835 1769 1836 1773
rect 1830 1768 1836 1769
rect 110 1756 116 1757
rect 110 1752 111 1756
rect 115 1752 116 1756
rect 110 1751 116 1752
rect 1830 1756 1836 1757
rect 1830 1752 1831 1756
rect 1835 1752 1836 1756
rect 1872 1754 1874 1773
rect 1896 1757 1898 1773
rect 2024 1757 2026 1773
rect 2184 1757 2186 1773
rect 2352 1757 2354 1773
rect 2552 1757 2554 1773
rect 2776 1757 2778 1773
rect 3016 1757 3018 1773
rect 3272 1757 3274 1773
rect 3504 1757 3506 1773
rect 1894 1756 1900 1757
rect 1830 1751 1836 1752
rect 1870 1753 1876 1754
rect 112 1715 114 1751
rect 142 1738 148 1739
rect 142 1734 143 1738
rect 147 1734 148 1738
rect 142 1733 148 1734
rect 318 1738 324 1739
rect 318 1734 319 1738
rect 323 1734 324 1738
rect 318 1733 324 1734
rect 510 1738 516 1739
rect 510 1734 511 1738
rect 515 1734 516 1738
rect 510 1733 516 1734
rect 694 1738 700 1739
rect 694 1734 695 1738
rect 699 1734 700 1738
rect 694 1733 700 1734
rect 854 1738 860 1739
rect 854 1734 855 1738
rect 859 1734 860 1738
rect 854 1733 860 1734
rect 998 1738 1004 1739
rect 998 1734 999 1738
rect 1003 1734 1004 1738
rect 998 1733 1004 1734
rect 1134 1738 1140 1739
rect 1134 1734 1135 1738
rect 1139 1734 1140 1738
rect 1134 1733 1140 1734
rect 1254 1738 1260 1739
rect 1254 1734 1255 1738
rect 1259 1734 1260 1738
rect 1254 1733 1260 1734
rect 1366 1738 1372 1739
rect 1366 1734 1367 1738
rect 1371 1734 1372 1738
rect 1366 1733 1372 1734
rect 1470 1738 1476 1739
rect 1470 1734 1471 1738
rect 1475 1734 1476 1738
rect 1470 1733 1476 1734
rect 1566 1738 1572 1739
rect 1566 1734 1567 1738
rect 1571 1734 1572 1738
rect 1566 1733 1572 1734
rect 1670 1738 1676 1739
rect 1670 1734 1671 1738
rect 1675 1734 1676 1738
rect 1670 1733 1676 1734
rect 1750 1738 1756 1739
rect 1750 1734 1751 1738
rect 1755 1734 1756 1738
rect 1750 1733 1756 1734
rect 144 1715 146 1733
rect 320 1715 322 1733
rect 512 1715 514 1733
rect 696 1715 698 1733
rect 856 1715 858 1733
rect 1000 1715 1002 1733
rect 1136 1715 1138 1733
rect 1256 1715 1258 1733
rect 1368 1715 1370 1733
rect 1472 1715 1474 1733
rect 1568 1715 1570 1733
rect 1672 1715 1674 1733
rect 1752 1715 1754 1733
rect 1832 1715 1834 1751
rect 1870 1749 1871 1753
rect 1875 1749 1876 1753
rect 1894 1752 1895 1756
rect 1899 1752 1900 1756
rect 1894 1751 1900 1752
rect 2022 1756 2028 1757
rect 2022 1752 2023 1756
rect 2027 1752 2028 1756
rect 2022 1751 2028 1752
rect 2182 1756 2188 1757
rect 2182 1752 2183 1756
rect 2187 1752 2188 1756
rect 2182 1751 2188 1752
rect 2350 1756 2356 1757
rect 2350 1752 2351 1756
rect 2355 1752 2356 1756
rect 2350 1751 2356 1752
rect 2550 1756 2556 1757
rect 2550 1752 2551 1756
rect 2555 1752 2556 1756
rect 2550 1751 2556 1752
rect 2774 1756 2780 1757
rect 2774 1752 2775 1756
rect 2779 1752 2780 1756
rect 2774 1751 2780 1752
rect 3014 1756 3020 1757
rect 3014 1752 3015 1756
rect 3019 1752 3020 1756
rect 3014 1751 3020 1752
rect 3270 1756 3276 1757
rect 3270 1752 3271 1756
rect 3275 1752 3276 1756
rect 3270 1751 3276 1752
rect 3502 1756 3508 1757
rect 3502 1752 3503 1756
rect 3507 1752 3508 1756
rect 3592 1754 3594 1773
rect 3502 1751 3508 1752
rect 3590 1753 3596 1754
rect 1870 1748 1876 1749
rect 3590 1749 3591 1753
rect 3595 1749 3596 1753
rect 3590 1748 3596 1749
rect 1870 1736 1876 1737
rect 1870 1732 1871 1736
rect 1875 1732 1876 1736
rect 1870 1731 1876 1732
rect 3590 1736 3596 1737
rect 3590 1732 3591 1736
rect 3595 1732 3596 1736
rect 3590 1731 3596 1732
rect 111 1714 115 1715
rect 111 1709 115 1710
rect 143 1714 147 1715
rect 143 1709 147 1710
rect 239 1714 243 1715
rect 239 1709 243 1710
rect 319 1714 323 1715
rect 319 1709 323 1710
rect 367 1714 371 1715
rect 367 1709 371 1710
rect 487 1714 491 1715
rect 487 1709 491 1710
rect 511 1714 515 1715
rect 511 1709 515 1710
rect 607 1714 611 1715
rect 607 1709 611 1710
rect 695 1714 699 1715
rect 695 1709 699 1710
rect 719 1714 723 1715
rect 719 1709 723 1710
rect 823 1714 827 1715
rect 823 1709 827 1710
rect 855 1714 859 1715
rect 855 1709 859 1710
rect 927 1714 931 1715
rect 927 1709 931 1710
rect 999 1714 1003 1715
rect 999 1709 1003 1710
rect 1023 1714 1027 1715
rect 1023 1709 1027 1710
rect 1119 1714 1123 1715
rect 1119 1709 1123 1710
rect 1135 1714 1139 1715
rect 1135 1709 1139 1710
rect 1215 1714 1219 1715
rect 1215 1709 1219 1710
rect 1255 1714 1259 1715
rect 1255 1709 1259 1710
rect 1319 1714 1323 1715
rect 1319 1709 1323 1710
rect 1367 1714 1371 1715
rect 1367 1709 1371 1710
rect 1471 1714 1475 1715
rect 1471 1709 1475 1710
rect 1567 1714 1571 1715
rect 1567 1709 1571 1710
rect 1671 1714 1675 1715
rect 1671 1709 1675 1710
rect 1751 1714 1755 1715
rect 1751 1709 1755 1710
rect 1831 1714 1835 1715
rect 1831 1709 1835 1710
rect 112 1681 114 1709
rect 144 1699 146 1709
rect 240 1699 242 1709
rect 368 1699 370 1709
rect 488 1699 490 1709
rect 608 1699 610 1709
rect 720 1699 722 1709
rect 824 1699 826 1709
rect 928 1699 930 1709
rect 1024 1699 1026 1709
rect 1120 1699 1122 1709
rect 1216 1699 1218 1709
rect 1320 1699 1322 1709
rect 142 1698 148 1699
rect 142 1694 143 1698
rect 147 1694 148 1698
rect 142 1693 148 1694
rect 238 1698 244 1699
rect 238 1694 239 1698
rect 243 1694 244 1698
rect 238 1693 244 1694
rect 366 1698 372 1699
rect 366 1694 367 1698
rect 371 1694 372 1698
rect 366 1693 372 1694
rect 486 1698 492 1699
rect 486 1694 487 1698
rect 491 1694 492 1698
rect 486 1693 492 1694
rect 606 1698 612 1699
rect 606 1694 607 1698
rect 611 1694 612 1698
rect 606 1693 612 1694
rect 718 1698 724 1699
rect 718 1694 719 1698
rect 723 1694 724 1698
rect 718 1693 724 1694
rect 822 1698 828 1699
rect 822 1694 823 1698
rect 827 1694 828 1698
rect 822 1693 828 1694
rect 926 1698 932 1699
rect 926 1694 927 1698
rect 931 1694 932 1698
rect 926 1693 932 1694
rect 1022 1698 1028 1699
rect 1022 1694 1023 1698
rect 1027 1694 1028 1698
rect 1022 1693 1028 1694
rect 1118 1698 1124 1699
rect 1118 1694 1119 1698
rect 1123 1694 1124 1698
rect 1118 1693 1124 1694
rect 1214 1698 1220 1699
rect 1214 1694 1215 1698
rect 1219 1694 1220 1698
rect 1214 1693 1220 1694
rect 1318 1698 1324 1699
rect 1318 1694 1319 1698
rect 1323 1694 1324 1698
rect 1318 1693 1324 1694
rect 1832 1681 1834 1709
rect 1872 1703 1874 1731
rect 1902 1718 1908 1719
rect 1902 1714 1903 1718
rect 1907 1714 1908 1718
rect 1902 1713 1908 1714
rect 2030 1718 2036 1719
rect 2030 1714 2031 1718
rect 2035 1714 2036 1718
rect 2030 1713 2036 1714
rect 2190 1718 2196 1719
rect 2190 1714 2191 1718
rect 2195 1714 2196 1718
rect 2190 1713 2196 1714
rect 2358 1718 2364 1719
rect 2358 1714 2359 1718
rect 2363 1714 2364 1718
rect 2358 1713 2364 1714
rect 2558 1718 2564 1719
rect 2558 1714 2559 1718
rect 2563 1714 2564 1718
rect 2558 1713 2564 1714
rect 2782 1718 2788 1719
rect 2782 1714 2783 1718
rect 2787 1714 2788 1718
rect 2782 1713 2788 1714
rect 3022 1718 3028 1719
rect 3022 1714 3023 1718
rect 3027 1714 3028 1718
rect 3022 1713 3028 1714
rect 3278 1718 3284 1719
rect 3278 1714 3279 1718
rect 3283 1714 3284 1718
rect 3278 1713 3284 1714
rect 3510 1718 3516 1719
rect 3510 1714 3511 1718
rect 3515 1714 3516 1718
rect 3510 1713 3516 1714
rect 1904 1703 1906 1713
rect 2032 1703 2034 1713
rect 2192 1703 2194 1713
rect 2360 1703 2362 1713
rect 2560 1703 2562 1713
rect 2784 1703 2786 1713
rect 3024 1703 3026 1713
rect 3280 1703 3282 1713
rect 3512 1703 3514 1713
rect 3592 1703 3594 1731
rect 1871 1702 1875 1703
rect 1871 1697 1875 1698
rect 1903 1702 1907 1703
rect 1903 1697 1907 1698
rect 1991 1702 1995 1703
rect 1991 1697 1995 1698
rect 2031 1702 2035 1703
rect 2031 1697 2035 1698
rect 2111 1702 2115 1703
rect 2111 1697 2115 1698
rect 2191 1702 2195 1703
rect 2191 1697 2195 1698
rect 2231 1702 2235 1703
rect 2231 1697 2235 1698
rect 2351 1702 2355 1703
rect 2351 1697 2355 1698
rect 2359 1702 2363 1703
rect 2359 1697 2363 1698
rect 2479 1702 2483 1703
rect 2479 1697 2483 1698
rect 2559 1702 2563 1703
rect 2559 1697 2563 1698
rect 2607 1702 2611 1703
rect 2607 1697 2611 1698
rect 2743 1702 2747 1703
rect 2743 1697 2747 1698
rect 2783 1702 2787 1703
rect 2783 1697 2787 1698
rect 2887 1702 2891 1703
rect 2887 1697 2891 1698
rect 3023 1702 3027 1703
rect 3023 1697 3027 1698
rect 3039 1702 3043 1703
rect 3039 1697 3043 1698
rect 3199 1702 3203 1703
rect 3199 1697 3203 1698
rect 3279 1702 3283 1703
rect 3279 1697 3283 1698
rect 3367 1702 3371 1703
rect 3367 1697 3371 1698
rect 3511 1702 3515 1703
rect 3511 1697 3515 1698
rect 3591 1702 3595 1703
rect 3591 1697 3595 1698
rect 110 1680 116 1681
rect 110 1676 111 1680
rect 115 1676 116 1680
rect 110 1675 116 1676
rect 1830 1680 1836 1681
rect 1830 1676 1831 1680
rect 1835 1676 1836 1680
rect 1830 1675 1836 1676
rect 1872 1669 1874 1697
rect 1904 1687 1906 1697
rect 1992 1687 1994 1697
rect 2112 1687 2114 1697
rect 2232 1687 2234 1697
rect 2352 1687 2354 1697
rect 2480 1687 2482 1697
rect 2608 1687 2610 1697
rect 2744 1687 2746 1697
rect 2888 1687 2890 1697
rect 3040 1687 3042 1697
rect 3200 1687 3202 1697
rect 3368 1687 3370 1697
rect 3512 1687 3514 1697
rect 1902 1686 1908 1687
rect 1902 1682 1903 1686
rect 1907 1682 1908 1686
rect 1902 1681 1908 1682
rect 1990 1686 1996 1687
rect 1990 1682 1991 1686
rect 1995 1682 1996 1686
rect 1990 1681 1996 1682
rect 2110 1686 2116 1687
rect 2110 1682 2111 1686
rect 2115 1682 2116 1686
rect 2110 1681 2116 1682
rect 2230 1686 2236 1687
rect 2230 1682 2231 1686
rect 2235 1682 2236 1686
rect 2230 1681 2236 1682
rect 2350 1686 2356 1687
rect 2350 1682 2351 1686
rect 2355 1682 2356 1686
rect 2350 1681 2356 1682
rect 2478 1686 2484 1687
rect 2478 1682 2479 1686
rect 2483 1682 2484 1686
rect 2478 1681 2484 1682
rect 2606 1686 2612 1687
rect 2606 1682 2607 1686
rect 2611 1682 2612 1686
rect 2606 1681 2612 1682
rect 2742 1686 2748 1687
rect 2742 1682 2743 1686
rect 2747 1682 2748 1686
rect 2742 1681 2748 1682
rect 2886 1686 2892 1687
rect 2886 1682 2887 1686
rect 2891 1682 2892 1686
rect 2886 1681 2892 1682
rect 3038 1686 3044 1687
rect 3038 1682 3039 1686
rect 3043 1682 3044 1686
rect 3038 1681 3044 1682
rect 3198 1686 3204 1687
rect 3198 1682 3199 1686
rect 3203 1682 3204 1686
rect 3198 1681 3204 1682
rect 3366 1686 3372 1687
rect 3366 1682 3367 1686
rect 3371 1682 3372 1686
rect 3366 1681 3372 1682
rect 3510 1686 3516 1687
rect 3510 1682 3511 1686
rect 3515 1682 3516 1686
rect 3510 1681 3516 1682
rect 3592 1669 3594 1697
rect 1870 1668 1876 1669
rect 1870 1664 1871 1668
rect 1875 1664 1876 1668
rect 110 1663 116 1664
rect 110 1659 111 1663
rect 115 1659 116 1663
rect 1830 1663 1836 1664
rect 1870 1663 1876 1664
rect 3590 1668 3596 1669
rect 3590 1664 3591 1668
rect 3595 1664 3596 1668
rect 3590 1663 3596 1664
rect 110 1658 116 1659
rect 134 1660 140 1661
rect 112 1631 114 1658
rect 134 1656 135 1660
rect 139 1656 140 1660
rect 134 1655 140 1656
rect 230 1660 236 1661
rect 230 1656 231 1660
rect 235 1656 236 1660
rect 230 1655 236 1656
rect 358 1660 364 1661
rect 358 1656 359 1660
rect 363 1656 364 1660
rect 358 1655 364 1656
rect 478 1660 484 1661
rect 478 1656 479 1660
rect 483 1656 484 1660
rect 478 1655 484 1656
rect 598 1660 604 1661
rect 598 1656 599 1660
rect 603 1656 604 1660
rect 598 1655 604 1656
rect 710 1660 716 1661
rect 710 1656 711 1660
rect 715 1656 716 1660
rect 710 1655 716 1656
rect 814 1660 820 1661
rect 814 1656 815 1660
rect 819 1656 820 1660
rect 814 1655 820 1656
rect 918 1660 924 1661
rect 918 1656 919 1660
rect 923 1656 924 1660
rect 918 1655 924 1656
rect 1014 1660 1020 1661
rect 1014 1656 1015 1660
rect 1019 1656 1020 1660
rect 1014 1655 1020 1656
rect 1110 1660 1116 1661
rect 1110 1656 1111 1660
rect 1115 1656 1116 1660
rect 1110 1655 1116 1656
rect 1206 1660 1212 1661
rect 1206 1656 1207 1660
rect 1211 1656 1212 1660
rect 1206 1655 1212 1656
rect 1310 1660 1316 1661
rect 1310 1656 1311 1660
rect 1315 1656 1316 1660
rect 1830 1659 1831 1663
rect 1835 1659 1836 1663
rect 1830 1658 1836 1659
rect 1310 1655 1316 1656
rect 136 1631 138 1655
rect 232 1631 234 1655
rect 360 1631 362 1655
rect 480 1631 482 1655
rect 600 1631 602 1655
rect 712 1631 714 1655
rect 816 1631 818 1655
rect 920 1631 922 1655
rect 1016 1631 1018 1655
rect 1112 1631 1114 1655
rect 1208 1631 1210 1655
rect 1312 1631 1314 1655
rect 1832 1631 1834 1658
rect 1870 1651 1876 1652
rect 1870 1647 1871 1651
rect 1875 1647 1876 1651
rect 3590 1651 3596 1652
rect 1870 1646 1876 1647
rect 1894 1648 1900 1649
rect 111 1630 115 1631
rect 111 1625 115 1626
rect 135 1630 139 1631
rect 135 1625 139 1626
rect 175 1630 179 1631
rect 175 1625 179 1626
rect 231 1630 235 1631
rect 231 1625 235 1626
rect 311 1630 315 1631
rect 311 1625 315 1626
rect 359 1630 363 1631
rect 359 1625 363 1626
rect 439 1630 443 1631
rect 439 1625 443 1626
rect 479 1630 483 1631
rect 479 1625 483 1626
rect 567 1630 571 1631
rect 567 1625 571 1626
rect 599 1630 603 1631
rect 599 1625 603 1626
rect 687 1630 691 1631
rect 687 1625 691 1626
rect 711 1630 715 1631
rect 711 1625 715 1626
rect 799 1630 803 1631
rect 799 1625 803 1626
rect 815 1630 819 1631
rect 815 1625 819 1626
rect 903 1630 907 1631
rect 903 1625 907 1626
rect 919 1630 923 1631
rect 919 1625 923 1626
rect 999 1630 1003 1631
rect 999 1625 1003 1626
rect 1015 1630 1019 1631
rect 1015 1625 1019 1626
rect 1095 1630 1099 1631
rect 1095 1625 1099 1626
rect 1111 1630 1115 1631
rect 1111 1625 1115 1626
rect 1199 1630 1203 1631
rect 1199 1625 1203 1626
rect 1207 1630 1211 1631
rect 1207 1625 1211 1626
rect 1303 1630 1307 1631
rect 1303 1625 1307 1626
rect 1311 1630 1315 1631
rect 1311 1625 1315 1626
rect 1831 1630 1835 1631
rect 1872 1627 1874 1646
rect 1894 1644 1895 1648
rect 1899 1644 1900 1648
rect 1894 1643 1900 1644
rect 1982 1648 1988 1649
rect 1982 1644 1983 1648
rect 1987 1644 1988 1648
rect 1982 1643 1988 1644
rect 2102 1648 2108 1649
rect 2102 1644 2103 1648
rect 2107 1644 2108 1648
rect 2102 1643 2108 1644
rect 2222 1648 2228 1649
rect 2222 1644 2223 1648
rect 2227 1644 2228 1648
rect 2222 1643 2228 1644
rect 2342 1648 2348 1649
rect 2342 1644 2343 1648
rect 2347 1644 2348 1648
rect 2342 1643 2348 1644
rect 2470 1648 2476 1649
rect 2470 1644 2471 1648
rect 2475 1644 2476 1648
rect 2470 1643 2476 1644
rect 2598 1648 2604 1649
rect 2598 1644 2599 1648
rect 2603 1644 2604 1648
rect 2598 1643 2604 1644
rect 2734 1648 2740 1649
rect 2734 1644 2735 1648
rect 2739 1644 2740 1648
rect 2734 1643 2740 1644
rect 2878 1648 2884 1649
rect 2878 1644 2879 1648
rect 2883 1644 2884 1648
rect 2878 1643 2884 1644
rect 3030 1648 3036 1649
rect 3030 1644 3031 1648
rect 3035 1644 3036 1648
rect 3030 1643 3036 1644
rect 3190 1648 3196 1649
rect 3190 1644 3191 1648
rect 3195 1644 3196 1648
rect 3190 1643 3196 1644
rect 3358 1648 3364 1649
rect 3358 1644 3359 1648
rect 3363 1644 3364 1648
rect 3358 1643 3364 1644
rect 3502 1648 3508 1649
rect 3502 1644 3503 1648
rect 3507 1644 3508 1648
rect 3590 1647 3591 1651
rect 3595 1647 3596 1651
rect 3590 1646 3596 1647
rect 3502 1643 3508 1644
rect 1896 1627 1898 1643
rect 1984 1627 1986 1643
rect 2104 1627 2106 1643
rect 2224 1627 2226 1643
rect 2344 1627 2346 1643
rect 2472 1627 2474 1643
rect 2600 1627 2602 1643
rect 2736 1627 2738 1643
rect 2880 1627 2882 1643
rect 3032 1627 3034 1643
rect 3192 1627 3194 1643
rect 3360 1627 3362 1643
rect 3504 1627 3506 1643
rect 3592 1627 3594 1646
rect 1831 1625 1835 1626
rect 1871 1626 1875 1627
rect 112 1606 114 1625
rect 176 1609 178 1625
rect 312 1609 314 1625
rect 440 1609 442 1625
rect 568 1609 570 1625
rect 688 1609 690 1625
rect 800 1609 802 1625
rect 904 1609 906 1625
rect 1000 1609 1002 1625
rect 1096 1609 1098 1625
rect 1200 1609 1202 1625
rect 1304 1609 1306 1625
rect 174 1608 180 1609
rect 110 1605 116 1606
rect 110 1601 111 1605
rect 115 1601 116 1605
rect 174 1604 175 1608
rect 179 1604 180 1608
rect 174 1603 180 1604
rect 310 1608 316 1609
rect 310 1604 311 1608
rect 315 1604 316 1608
rect 310 1603 316 1604
rect 438 1608 444 1609
rect 438 1604 439 1608
rect 443 1604 444 1608
rect 438 1603 444 1604
rect 566 1608 572 1609
rect 566 1604 567 1608
rect 571 1604 572 1608
rect 566 1603 572 1604
rect 686 1608 692 1609
rect 686 1604 687 1608
rect 691 1604 692 1608
rect 686 1603 692 1604
rect 798 1608 804 1609
rect 798 1604 799 1608
rect 803 1604 804 1608
rect 798 1603 804 1604
rect 902 1608 908 1609
rect 902 1604 903 1608
rect 907 1604 908 1608
rect 902 1603 908 1604
rect 998 1608 1004 1609
rect 998 1604 999 1608
rect 1003 1604 1004 1608
rect 998 1603 1004 1604
rect 1094 1608 1100 1609
rect 1094 1604 1095 1608
rect 1099 1604 1100 1608
rect 1094 1603 1100 1604
rect 1198 1608 1204 1609
rect 1198 1604 1199 1608
rect 1203 1604 1204 1608
rect 1198 1603 1204 1604
rect 1302 1608 1308 1609
rect 1302 1604 1303 1608
rect 1307 1604 1308 1608
rect 1832 1606 1834 1625
rect 1871 1621 1875 1622
rect 1895 1626 1899 1627
rect 1895 1621 1899 1622
rect 1927 1626 1931 1627
rect 1927 1621 1931 1622
rect 1983 1626 1987 1627
rect 1983 1621 1987 1622
rect 2023 1626 2027 1627
rect 2023 1621 2027 1622
rect 2103 1626 2107 1627
rect 2103 1621 2107 1622
rect 2135 1626 2139 1627
rect 2135 1621 2139 1622
rect 2223 1626 2227 1627
rect 2223 1621 2227 1622
rect 2263 1626 2267 1627
rect 2263 1621 2267 1622
rect 2343 1626 2347 1627
rect 2343 1621 2347 1622
rect 2391 1626 2395 1627
rect 2391 1621 2395 1622
rect 2471 1626 2475 1627
rect 2471 1621 2475 1622
rect 2527 1626 2531 1627
rect 2527 1621 2531 1622
rect 2599 1626 2603 1627
rect 2599 1621 2603 1622
rect 2671 1626 2675 1627
rect 2671 1621 2675 1622
rect 2735 1626 2739 1627
rect 2735 1621 2739 1622
rect 2823 1626 2827 1627
rect 2823 1621 2827 1622
rect 2879 1626 2883 1627
rect 2879 1621 2883 1622
rect 2983 1626 2987 1627
rect 2983 1621 2987 1622
rect 3031 1626 3035 1627
rect 3031 1621 3035 1622
rect 3159 1626 3163 1627
rect 3159 1621 3163 1622
rect 3191 1626 3195 1627
rect 3191 1621 3195 1622
rect 3343 1626 3347 1627
rect 3343 1621 3347 1622
rect 3359 1626 3363 1627
rect 3359 1621 3363 1622
rect 3503 1626 3507 1627
rect 3503 1621 3507 1622
rect 3591 1626 3595 1627
rect 3591 1621 3595 1622
rect 1302 1603 1308 1604
rect 1830 1605 1836 1606
rect 110 1600 116 1601
rect 1830 1601 1831 1605
rect 1835 1601 1836 1605
rect 1872 1602 1874 1621
rect 1928 1605 1930 1621
rect 2024 1605 2026 1621
rect 2136 1605 2138 1621
rect 2264 1605 2266 1621
rect 2392 1605 2394 1621
rect 2528 1605 2530 1621
rect 2672 1605 2674 1621
rect 2824 1605 2826 1621
rect 2984 1605 2986 1621
rect 3160 1605 3162 1621
rect 3344 1605 3346 1621
rect 3504 1605 3506 1621
rect 1926 1604 1932 1605
rect 1830 1600 1836 1601
rect 1870 1601 1876 1602
rect 1870 1597 1871 1601
rect 1875 1597 1876 1601
rect 1926 1600 1927 1604
rect 1931 1600 1932 1604
rect 1926 1599 1932 1600
rect 2022 1604 2028 1605
rect 2022 1600 2023 1604
rect 2027 1600 2028 1604
rect 2022 1599 2028 1600
rect 2134 1604 2140 1605
rect 2134 1600 2135 1604
rect 2139 1600 2140 1604
rect 2134 1599 2140 1600
rect 2262 1604 2268 1605
rect 2262 1600 2263 1604
rect 2267 1600 2268 1604
rect 2262 1599 2268 1600
rect 2390 1604 2396 1605
rect 2390 1600 2391 1604
rect 2395 1600 2396 1604
rect 2390 1599 2396 1600
rect 2526 1604 2532 1605
rect 2526 1600 2527 1604
rect 2531 1600 2532 1604
rect 2526 1599 2532 1600
rect 2670 1604 2676 1605
rect 2670 1600 2671 1604
rect 2675 1600 2676 1604
rect 2670 1599 2676 1600
rect 2822 1604 2828 1605
rect 2822 1600 2823 1604
rect 2827 1600 2828 1604
rect 2822 1599 2828 1600
rect 2982 1604 2988 1605
rect 2982 1600 2983 1604
rect 2987 1600 2988 1604
rect 2982 1599 2988 1600
rect 3158 1604 3164 1605
rect 3158 1600 3159 1604
rect 3163 1600 3164 1604
rect 3158 1599 3164 1600
rect 3342 1604 3348 1605
rect 3342 1600 3343 1604
rect 3347 1600 3348 1604
rect 3342 1599 3348 1600
rect 3502 1604 3508 1605
rect 3502 1600 3503 1604
rect 3507 1600 3508 1604
rect 3592 1602 3594 1621
rect 3502 1599 3508 1600
rect 3590 1601 3596 1602
rect 1870 1596 1876 1597
rect 3590 1597 3591 1601
rect 3595 1597 3596 1601
rect 3590 1596 3596 1597
rect 110 1588 116 1589
rect 110 1584 111 1588
rect 115 1584 116 1588
rect 110 1583 116 1584
rect 1830 1588 1836 1589
rect 1830 1584 1831 1588
rect 1835 1584 1836 1588
rect 1830 1583 1836 1584
rect 1870 1584 1876 1585
rect 112 1547 114 1583
rect 182 1570 188 1571
rect 182 1566 183 1570
rect 187 1566 188 1570
rect 182 1565 188 1566
rect 318 1570 324 1571
rect 318 1566 319 1570
rect 323 1566 324 1570
rect 318 1565 324 1566
rect 446 1570 452 1571
rect 446 1566 447 1570
rect 451 1566 452 1570
rect 446 1565 452 1566
rect 574 1570 580 1571
rect 574 1566 575 1570
rect 579 1566 580 1570
rect 574 1565 580 1566
rect 694 1570 700 1571
rect 694 1566 695 1570
rect 699 1566 700 1570
rect 694 1565 700 1566
rect 806 1570 812 1571
rect 806 1566 807 1570
rect 811 1566 812 1570
rect 806 1565 812 1566
rect 910 1570 916 1571
rect 910 1566 911 1570
rect 915 1566 916 1570
rect 910 1565 916 1566
rect 1006 1570 1012 1571
rect 1006 1566 1007 1570
rect 1011 1566 1012 1570
rect 1006 1565 1012 1566
rect 1102 1570 1108 1571
rect 1102 1566 1103 1570
rect 1107 1566 1108 1570
rect 1102 1565 1108 1566
rect 1206 1570 1212 1571
rect 1206 1566 1207 1570
rect 1211 1566 1212 1570
rect 1206 1565 1212 1566
rect 1310 1570 1316 1571
rect 1310 1566 1311 1570
rect 1315 1566 1316 1570
rect 1310 1565 1316 1566
rect 184 1547 186 1565
rect 320 1547 322 1565
rect 448 1547 450 1565
rect 576 1547 578 1565
rect 696 1547 698 1565
rect 808 1547 810 1565
rect 912 1547 914 1565
rect 1008 1547 1010 1565
rect 1104 1547 1106 1565
rect 1208 1547 1210 1565
rect 1312 1547 1314 1565
rect 1832 1547 1834 1583
rect 1870 1580 1871 1584
rect 1875 1580 1876 1584
rect 1870 1579 1876 1580
rect 3590 1584 3596 1585
rect 3590 1580 3591 1584
rect 3595 1580 3596 1584
rect 3590 1579 3596 1580
rect 111 1546 115 1547
rect 111 1541 115 1542
rect 183 1546 187 1547
rect 183 1541 187 1542
rect 239 1546 243 1547
rect 239 1541 243 1542
rect 319 1546 323 1547
rect 319 1541 323 1542
rect 343 1546 347 1547
rect 343 1541 347 1542
rect 447 1546 451 1547
rect 447 1541 451 1542
rect 463 1546 467 1547
rect 463 1541 467 1542
rect 575 1546 579 1547
rect 575 1541 579 1542
rect 591 1546 595 1547
rect 591 1541 595 1542
rect 695 1546 699 1547
rect 695 1541 699 1542
rect 719 1546 723 1547
rect 719 1541 723 1542
rect 807 1546 811 1547
rect 807 1541 811 1542
rect 855 1546 859 1547
rect 855 1541 859 1542
rect 911 1546 915 1547
rect 911 1541 915 1542
rect 983 1546 987 1547
rect 983 1541 987 1542
rect 1007 1546 1011 1547
rect 1007 1541 1011 1542
rect 1103 1546 1107 1547
rect 1103 1541 1107 1542
rect 1111 1546 1115 1547
rect 1111 1541 1115 1542
rect 1207 1546 1211 1547
rect 1207 1541 1211 1542
rect 1231 1546 1235 1547
rect 1231 1541 1235 1542
rect 1311 1546 1315 1547
rect 1311 1541 1315 1542
rect 1343 1546 1347 1547
rect 1343 1541 1347 1542
rect 1455 1546 1459 1547
rect 1455 1541 1459 1542
rect 1575 1546 1579 1547
rect 1575 1541 1579 1542
rect 1831 1546 1835 1547
rect 1872 1543 1874 1579
rect 1934 1566 1940 1567
rect 1934 1562 1935 1566
rect 1939 1562 1940 1566
rect 1934 1561 1940 1562
rect 2030 1566 2036 1567
rect 2030 1562 2031 1566
rect 2035 1562 2036 1566
rect 2030 1561 2036 1562
rect 2142 1566 2148 1567
rect 2142 1562 2143 1566
rect 2147 1562 2148 1566
rect 2142 1561 2148 1562
rect 2270 1566 2276 1567
rect 2270 1562 2271 1566
rect 2275 1562 2276 1566
rect 2270 1561 2276 1562
rect 2398 1566 2404 1567
rect 2398 1562 2399 1566
rect 2403 1562 2404 1566
rect 2398 1561 2404 1562
rect 2534 1566 2540 1567
rect 2534 1562 2535 1566
rect 2539 1562 2540 1566
rect 2534 1561 2540 1562
rect 2678 1566 2684 1567
rect 2678 1562 2679 1566
rect 2683 1562 2684 1566
rect 2678 1561 2684 1562
rect 2830 1566 2836 1567
rect 2830 1562 2831 1566
rect 2835 1562 2836 1566
rect 2830 1561 2836 1562
rect 2990 1566 2996 1567
rect 2990 1562 2991 1566
rect 2995 1562 2996 1566
rect 2990 1561 2996 1562
rect 3166 1566 3172 1567
rect 3166 1562 3167 1566
rect 3171 1562 3172 1566
rect 3166 1561 3172 1562
rect 3350 1566 3356 1567
rect 3350 1562 3351 1566
rect 3355 1562 3356 1566
rect 3350 1561 3356 1562
rect 3510 1566 3516 1567
rect 3510 1562 3511 1566
rect 3515 1562 3516 1566
rect 3510 1561 3516 1562
rect 1936 1543 1938 1561
rect 2032 1543 2034 1561
rect 2144 1543 2146 1561
rect 2272 1543 2274 1561
rect 2400 1543 2402 1561
rect 2536 1543 2538 1561
rect 2680 1543 2682 1561
rect 2832 1543 2834 1561
rect 2992 1543 2994 1561
rect 3168 1543 3170 1561
rect 3352 1543 3354 1561
rect 3512 1543 3514 1561
rect 3592 1543 3594 1579
rect 1831 1541 1835 1542
rect 1871 1542 1875 1543
rect 112 1513 114 1541
rect 240 1531 242 1541
rect 344 1531 346 1541
rect 464 1531 466 1541
rect 592 1531 594 1541
rect 720 1531 722 1541
rect 856 1531 858 1541
rect 984 1531 986 1541
rect 1112 1531 1114 1541
rect 1232 1531 1234 1541
rect 1344 1531 1346 1541
rect 1456 1531 1458 1541
rect 1576 1531 1578 1541
rect 238 1530 244 1531
rect 238 1526 239 1530
rect 243 1526 244 1530
rect 238 1525 244 1526
rect 342 1530 348 1531
rect 342 1526 343 1530
rect 347 1526 348 1530
rect 342 1525 348 1526
rect 462 1530 468 1531
rect 462 1526 463 1530
rect 467 1526 468 1530
rect 462 1525 468 1526
rect 590 1530 596 1531
rect 590 1526 591 1530
rect 595 1526 596 1530
rect 590 1525 596 1526
rect 718 1530 724 1531
rect 718 1526 719 1530
rect 723 1526 724 1530
rect 718 1525 724 1526
rect 854 1530 860 1531
rect 854 1526 855 1530
rect 859 1526 860 1530
rect 854 1525 860 1526
rect 982 1530 988 1531
rect 982 1526 983 1530
rect 987 1526 988 1530
rect 982 1525 988 1526
rect 1110 1530 1116 1531
rect 1110 1526 1111 1530
rect 1115 1526 1116 1530
rect 1110 1525 1116 1526
rect 1230 1530 1236 1531
rect 1230 1526 1231 1530
rect 1235 1526 1236 1530
rect 1230 1525 1236 1526
rect 1342 1530 1348 1531
rect 1342 1526 1343 1530
rect 1347 1526 1348 1530
rect 1342 1525 1348 1526
rect 1454 1530 1460 1531
rect 1454 1526 1455 1530
rect 1459 1526 1460 1530
rect 1454 1525 1460 1526
rect 1574 1530 1580 1531
rect 1574 1526 1575 1530
rect 1579 1526 1580 1530
rect 1574 1525 1580 1526
rect 1832 1513 1834 1541
rect 1871 1537 1875 1538
rect 1935 1542 1939 1543
rect 1935 1537 1939 1538
rect 2031 1542 2035 1543
rect 2031 1537 2035 1538
rect 2135 1542 2139 1543
rect 2135 1537 2139 1538
rect 2143 1542 2147 1543
rect 2143 1537 2147 1538
rect 2255 1542 2259 1543
rect 2255 1537 2259 1538
rect 2271 1542 2275 1543
rect 2271 1537 2275 1538
rect 2383 1542 2387 1543
rect 2383 1537 2387 1538
rect 2399 1542 2403 1543
rect 2399 1537 2403 1538
rect 2511 1542 2515 1543
rect 2511 1537 2515 1538
rect 2535 1542 2539 1543
rect 2535 1537 2539 1538
rect 2639 1542 2643 1543
rect 2639 1537 2643 1538
rect 2679 1542 2683 1543
rect 2679 1537 2683 1538
rect 2767 1542 2771 1543
rect 2767 1537 2771 1538
rect 2831 1542 2835 1543
rect 2831 1537 2835 1538
rect 2887 1542 2891 1543
rect 2887 1537 2891 1538
rect 2991 1542 2995 1543
rect 2991 1537 2995 1538
rect 3007 1542 3011 1543
rect 3007 1537 3011 1538
rect 3119 1542 3123 1543
rect 3119 1537 3123 1538
rect 3167 1542 3171 1543
rect 3167 1537 3171 1538
rect 3231 1542 3235 1543
rect 3231 1537 3235 1538
rect 3351 1542 3355 1543
rect 3351 1537 3355 1538
rect 3511 1542 3515 1543
rect 3511 1537 3515 1538
rect 3591 1542 3595 1543
rect 3591 1537 3595 1538
rect 110 1512 116 1513
rect 110 1508 111 1512
rect 115 1508 116 1512
rect 110 1507 116 1508
rect 1830 1512 1836 1513
rect 1830 1508 1831 1512
rect 1835 1508 1836 1512
rect 1872 1509 1874 1537
rect 2136 1527 2138 1537
rect 2256 1527 2258 1537
rect 2384 1527 2386 1537
rect 2512 1527 2514 1537
rect 2640 1527 2642 1537
rect 2768 1527 2770 1537
rect 2888 1527 2890 1537
rect 3008 1527 3010 1537
rect 3120 1527 3122 1537
rect 3232 1527 3234 1537
rect 3352 1527 3354 1537
rect 2134 1526 2140 1527
rect 2134 1522 2135 1526
rect 2139 1522 2140 1526
rect 2134 1521 2140 1522
rect 2254 1526 2260 1527
rect 2254 1522 2255 1526
rect 2259 1522 2260 1526
rect 2254 1521 2260 1522
rect 2382 1526 2388 1527
rect 2382 1522 2383 1526
rect 2387 1522 2388 1526
rect 2382 1521 2388 1522
rect 2510 1526 2516 1527
rect 2510 1522 2511 1526
rect 2515 1522 2516 1526
rect 2510 1521 2516 1522
rect 2638 1526 2644 1527
rect 2638 1522 2639 1526
rect 2643 1522 2644 1526
rect 2638 1521 2644 1522
rect 2766 1526 2772 1527
rect 2766 1522 2767 1526
rect 2771 1522 2772 1526
rect 2766 1521 2772 1522
rect 2886 1526 2892 1527
rect 2886 1522 2887 1526
rect 2891 1522 2892 1526
rect 2886 1521 2892 1522
rect 3006 1526 3012 1527
rect 3006 1522 3007 1526
rect 3011 1522 3012 1526
rect 3006 1521 3012 1522
rect 3118 1526 3124 1527
rect 3118 1522 3119 1526
rect 3123 1522 3124 1526
rect 3118 1521 3124 1522
rect 3230 1526 3236 1527
rect 3230 1522 3231 1526
rect 3235 1522 3236 1526
rect 3230 1521 3236 1522
rect 3350 1526 3356 1527
rect 3350 1522 3351 1526
rect 3355 1522 3356 1526
rect 3350 1521 3356 1522
rect 3592 1509 3594 1537
rect 1830 1507 1836 1508
rect 1870 1508 1876 1509
rect 1870 1504 1871 1508
rect 1875 1504 1876 1508
rect 1870 1503 1876 1504
rect 3590 1508 3596 1509
rect 3590 1504 3591 1508
rect 3595 1504 3596 1508
rect 3590 1503 3596 1504
rect 110 1495 116 1496
rect 110 1491 111 1495
rect 115 1491 116 1495
rect 1830 1495 1836 1496
rect 110 1490 116 1491
rect 230 1492 236 1493
rect 112 1459 114 1490
rect 230 1488 231 1492
rect 235 1488 236 1492
rect 230 1487 236 1488
rect 334 1492 340 1493
rect 334 1488 335 1492
rect 339 1488 340 1492
rect 334 1487 340 1488
rect 454 1492 460 1493
rect 454 1488 455 1492
rect 459 1488 460 1492
rect 454 1487 460 1488
rect 582 1492 588 1493
rect 582 1488 583 1492
rect 587 1488 588 1492
rect 582 1487 588 1488
rect 710 1492 716 1493
rect 710 1488 711 1492
rect 715 1488 716 1492
rect 710 1487 716 1488
rect 846 1492 852 1493
rect 846 1488 847 1492
rect 851 1488 852 1492
rect 846 1487 852 1488
rect 974 1492 980 1493
rect 974 1488 975 1492
rect 979 1488 980 1492
rect 974 1487 980 1488
rect 1102 1492 1108 1493
rect 1102 1488 1103 1492
rect 1107 1488 1108 1492
rect 1102 1487 1108 1488
rect 1222 1492 1228 1493
rect 1222 1488 1223 1492
rect 1227 1488 1228 1492
rect 1222 1487 1228 1488
rect 1334 1492 1340 1493
rect 1334 1488 1335 1492
rect 1339 1488 1340 1492
rect 1334 1487 1340 1488
rect 1446 1492 1452 1493
rect 1446 1488 1447 1492
rect 1451 1488 1452 1492
rect 1446 1487 1452 1488
rect 1566 1492 1572 1493
rect 1566 1488 1567 1492
rect 1571 1488 1572 1492
rect 1830 1491 1831 1495
rect 1835 1491 1836 1495
rect 1830 1490 1836 1491
rect 1870 1491 1876 1492
rect 1566 1487 1572 1488
rect 232 1459 234 1487
rect 336 1459 338 1487
rect 456 1459 458 1487
rect 584 1459 586 1487
rect 712 1459 714 1487
rect 848 1459 850 1487
rect 976 1459 978 1487
rect 1104 1459 1106 1487
rect 1224 1459 1226 1487
rect 1336 1459 1338 1487
rect 1448 1459 1450 1487
rect 1568 1459 1570 1487
rect 1832 1459 1834 1490
rect 1870 1487 1871 1491
rect 1875 1487 1876 1491
rect 3590 1491 3596 1492
rect 1870 1486 1876 1487
rect 2126 1488 2132 1489
rect 1872 1459 1874 1486
rect 2126 1484 2127 1488
rect 2131 1484 2132 1488
rect 2126 1483 2132 1484
rect 2246 1488 2252 1489
rect 2246 1484 2247 1488
rect 2251 1484 2252 1488
rect 2246 1483 2252 1484
rect 2374 1488 2380 1489
rect 2374 1484 2375 1488
rect 2379 1484 2380 1488
rect 2374 1483 2380 1484
rect 2502 1488 2508 1489
rect 2502 1484 2503 1488
rect 2507 1484 2508 1488
rect 2502 1483 2508 1484
rect 2630 1488 2636 1489
rect 2630 1484 2631 1488
rect 2635 1484 2636 1488
rect 2630 1483 2636 1484
rect 2758 1488 2764 1489
rect 2758 1484 2759 1488
rect 2763 1484 2764 1488
rect 2758 1483 2764 1484
rect 2878 1488 2884 1489
rect 2878 1484 2879 1488
rect 2883 1484 2884 1488
rect 2878 1483 2884 1484
rect 2998 1488 3004 1489
rect 2998 1484 2999 1488
rect 3003 1484 3004 1488
rect 2998 1483 3004 1484
rect 3110 1488 3116 1489
rect 3110 1484 3111 1488
rect 3115 1484 3116 1488
rect 3110 1483 3116 1484
rect 3222 1488 3228 1489
rect 3222 1484 3223 1488
rect 3227 1484 3228 1488
rect 3222 1483 3228 1484
rect 3342 1488 3348 1489
rect 3342 1484 3343 1488
rect 3347 1484 3348 1488
rect 3590 1487 3591 1491
rect 3595 1487 3596 1491
rect 3590 1486 3596 1487
rect 3342 1483 3348 1484
rect 2128 1459 2130 1483
rect 2248 1459 2250 1483
rect 2376 1459 2378 1483
rect 2504 1459 2506 1483
rect 2632 1459 2634 1483
rect 2760 1459 2762 1483
rect 2880 1459 2882 1483
rect 3000 1459 3002 1483
rect 3112 1459 3114 1483
rect 3224 1459 3226 1483
rect 3344 1459 3346 1483
rect 3592 1459 3594 1486
rect 111 1458 115 1459
rect 111 1453 115 1454
rect 231 1458 235 1459
rect 231 1453 235 1454
rect 279 1458 283 1459
rect 279 1453 283 1454
rect 335 1458 339 1459
rect 335 1453 339 1454
rect 383 1458 387 1459
rect 383 1453 387 1454
rect 455 1458 459 1459
rect 455 1453 459 1454
rect 511 1458 515 1459
rect 511 1453 515 1454
rect 583 1458 587 1459
rect 583 1453 587 1454
rect 655 1458 659 1459
rect 655 1453 659 1454
rect 711 1458 715 1459
rect 711 1453 715 1454
rect 807 1458 811 1459
rect 807 1453 811 1454
rect 847 1458 851 1459
rect 847 1453 851 1454
rect 959 1458 963 1459
rect 959 1453 963 1454
rect 975 1458 979 1459
rect 975 1453 979 1454
rect 1103 1458 1107 1459
rect 1103 1453 1107 1454
rect 1111 1458 1115 1459
rect 1111 1453 1115 1454
rect 1223 1458 1227 1459
rect 1223 1453 1227 1454
rect 1247 1458 1251 1459
rect 1247 1453 1251 1454
rect 1335 1458 1339 1459
rect 1335 1453 1339 1454
rect 1383 1458 1387 1459
rect 1383 1453 1387 1454
rect 1447 1458 1451 1459
rect 1447 1453 1451 1454
rect 1511 1458 1515 1459
rect 1511 1453 1515 1454
rect 1567 1458 1571 1459
rect 1567 1453 1571 1454
rect 1639 1458 1643 1459
rect 1639 1453 1643 1454
rect 1743 1458 1747 1459
rect 1743 1453 1747 1454
rect 1831 1458 1835 1459
rect 1831 1453 1835 1454
rect 1871 1458 1875 1459
rect 1871 1453 1875 1454
rect 2127 1458 2131 1459
rect 2127 1453 2131 1454
rect 2247 1458 2251 1459
rect 2247 1453 2251 1454
rect 2343 1458 2347 1459
rect 2343 1453 2347 1454
rect 2375 1458 2379 1459
rect 2375 1453 2379 1454
rect 2455 1458 2459 1459
rect 2455 1453 2459 1454
rect 2503 1458 2507 1459
rect 2503 1453 2507 1454
rect 2575 1458 2579 1459
rect 2575 1453 2579 1454
rect 2631 1458 2635 1459
rect 2631 1453 2635 1454
rect 2703 1458 2707 1459
rect 2703 1453 2707 1454
rect 2759 1458 2763 1459
rect 2759 1453 2763 1454
rect 2831 1458 2835 1459
rect 2831 1453 2835 1454
rect 2879 1458 2883 1459
rect 2879 1453 2883 1454
rect 2951 1458 2955 1459
rect 2951 1453 2955 1454
rect 2999 1458 3003 1459
rect 2999 1453 3003 1454
rect 3071 1458 3075 1459
rect 3071 1453 3075 1454
rect 3111 1458 3115 1459
rect 3111 1453 3115 1454
rect 3183 1458 3187 1459
rect 3183 1453 3187 1454
rect 3223 1458 3227 1459
rect 3223 1453 3227 1454
rect 3295 1458 3299 1459
rect 3295 1453 3299 1454
rect 3343 1458 3347 1459
rect 3343 1453 3347 1454
rect 3407 1458 3411 1459
rect 3407 1453 3411 1454
rect 3503 1458 3507 1459
rect 3503 1453 3507 1454
rect 3591 1458 3595 1459
rect 3591 1453 3595 1454
rect 112 1434 114 1453
rect 280 1437 282 1453
rect 384 1437 386 1453
rect 512 1437 514 1453
rect 656 1437 658 1453
rect 808 1437 810 1453
rect 960 1437 962 1453
rect 1112 1437 1114 1453
rect 1248 1437 1250 1453
rect 1384 1437 1386 1453
rect 1512 1437 1514 1453
rect 1640 1437 1642 1453
rect 1744 1437 1746 1453
rect 278 1436 284 1437
rect 110 1433 116 1434
rect 110 1429 111 1433
rect 115 1429 116 1433
rect 278 1432 279 1436
rect 283 1432 284 1436
rect 278 1431 284 1432
rect 382 1436 388 1437
rect 382 1432 383 1436
rect 387 1432 388 1436
rect 382 1431 388 1432
rect 510 1436 516 1437
rect 510 1432 511 1436
rect 515 1432 516 1436
rect 510 1431 516 1432
rect 654 1436 660 1437
rect 654 1432 655 1436
rect 659 1432 660 1436
rect 654 1431 660 1432
rect 806 1436 812 1437
rect 806 1432 807 1436
rect 811 1432 812 1436
rect 806 1431 812 1432
rect 958 1436 964 1437
rect 958 1432 959 1436
rect 963 1432 964 1436
rect 958 1431 964 1432
rect 1110 1436 1116 1437
rect 1110 1432 1111 1436
rect 1115 1432 1116 1436
rect 1110 1431 1116 1432
rect 1246 1436 1252 1437
rect 1246 1432 1247 1436
rect 1251 1432 1252 1436
rect 1246 1431 1252 1432
rect 1382 1436 1388 1437
rect 1382 1432 1383 1436
rect 1387 1432 1388 1436
rect 1382 1431 1388 1432
rect 1510 1436 1516 1437
rect 1510 1432 1511 1436
rect 1515 1432 1516 1436
rect 1510 1431 1516 1432
rect 1638 1436 1644 1437
rect 1638 1432 1639 1436
rect 1643 1432 1644 1436
rect 1638 1431 1644 1432
rect 1742 1436 1748 1437
rect 1742 1432 1743 1436
rect 1747 1432 1748 1436
rect 1832 1434 1834 1453
rect 1872 1434 1874 1453
rect 2248 1437 2250 1453
rect 2344 1437 2346 1453
rect 2456 1437 2458 1453
rect 2576 1437 2578 1453
rect 2704 1437 2706 1453
rect 2832 1437 2834 1453
rect 2952 1437 2954 1453
rect 3072 1437 3074 1453
rect 3184 1437 3186 1453
rect 3296 1437 3298 1453
rect 3408 1437 3410 1453
rect 3504 1437 3506 1453
rect 2246 1436 2252 1437
rect 1742 1431 1748 1432
rect 1830 1433 1836 1434
rect 110 1428 116 1429
rect 1830 1429 1831 1433
rect 1835 1429 1836 1433
rect 1830 1428 1836 1429
rect 1870 1433 1876 1434
rect 1870 1429 1871 1433
rect 1875 1429 1876 1433
rect 2246 1432 2247 1436
rect 2251 1432 2252 1436
rect 2246 1431 2252 1432
rect 2342 1436 2348 1437
rect 2342 1432 2343 1436
rect 2347 1432 2348 1436
rect 2342 1431 2348 1432
rect 2454 1436 2460 1437
rect 2454 1432 2455 1436
rect 2459 1432 2460 1436
rect 2454 1431 2460 1432
rect 2574 1436 2580 1437
rect 2574 1432 2575 1436
rect 2579 1432 2580 1436
rect 2574 1431 2580 1432
rect 2702 1436 2708 1437
rect 2702 1432 2703 1436
rect 2707 1432 2708 1436
rect 2702 1431 2708 1432
rect 2830 1436 2836 1437
rect 2830 1432 2831 1436
rect 2835 1432 2836 1436
rect 2830 1431 2836 1432
rect 2950 1436 2956 1437
rect 2950 1432 2951 1436
rect 2955 1432 2956 1436
rect 2950 1431 2956 1432
rect 3070 1436 3076 1437
rect 3070 1432 3071 1436
rect 3075 1432 3076 1436
rect 3070 1431 3076 1432
rect 3182 1436 3188 1437
rect 3182 1432 3183 1436
rect 3187 1432 3188 1436
rect 3182 1431 3188 1432
rect 3294 1436 3300 1437
rect 3294 1432 3295 1436
rect 3299 1432 3300 1436
rect 3294 1431 3300 1432
rect 3406 1436 3412 1437
rect 3406 1432 3407 1436
rect 3411 1432 3412 1436
rect 3406 1431 3412 1432
rect 3502 1436 3508 1437
rect 3502 1432 3503 1436
rect 3507 1432 3508 1436
rect 3592 1434 3594 1453
rect 3502 1431 3508 1432
rect 3590 1433 3596 1434
rect 1870 1428 1876 1429
rect 3590 1429 3591 1433
rect 3595 1429 3596 1433
rect 3590 1428 3596 1429
rect 110 1416 116 1417
rect 110 1412 111 1416
rect 115 1412 116 1416
rect 110 1411 116 1412
rect 1830 1416 1836 1417
rect 1830 1412 1831 1416
rect 1835 1412 1836 1416
rect 1830 1411 1836 1412
rect 1870 1416 1876 1417
rect 1870 1412 1871 1416
rect 1875 1412 1876 1416
rect 1870 1411 1876 1412
rect 3590 1416 3596 1417
rect 3590 1412 3591 1416
rect 3595 1412 3596 1416
rect 3590 1411 3596 1412
rect 112 1367 114 1411
rect 286 1398 292 1399
rect 286 1394 287 1398
rect 291 1394 292 1398
rect 286 1393 292 1394
rect 390 1398 396 1399
rect 390 1394 391 1398
rect 395 1394 396 1398
rect 390 1393 396 1394
rect 518 1398 524 1399
rect 518 1394 519 1398
rect 523 1394 524 1398
rect 518 1393 524 1394
rect 662 1398 668 1399
rect 662 1394 663 1398
rect 667 1394 668 1398
rect 662 1393 668 1394
rect 814 1398 820 1399
rect 814 1394 815 1398
rect 819 1394 820 1398
rect 814 1393 820 1394
rect 966 1398 972 1399
rect 966 1394 967 1398
rect 971 1394 972 1398
rect 966 1393 972 1394
rect 1118 1398 1124 1399
rect 1118 1394 1119 1398
rect 1123 1394 1124 1398
rect 1118 1393 1124 1394
rect 1254 1398 1260 1399
rect 1254 1394 1255 1398
rect 1259 1394 1260 1398
rect 1254 1393 1260 1394
rect 1390 1398 1396 1399
rect 1390 1394 1391 1398
rect 1395 1394 1396 1398
rect 1390 1393 1396 1394
rect 1518 1398 1524 1399
rect 1518 1394 1519 1398
rect 1523 1394 1524 1398
rect 1518 1393 1524 1394
rect 1646 1398 1652 1399
rect 1646 1394 1647 1398
rect 1651 1394 1652 1398
rect 1646 1393 1652 1394
rect 1750 1398 1756 1399
rect 1750 1394 1751 1398
rect 1755 1394 1756 1398
rect 1750 1393 1756 1394
rect 288 1367 290 1393
rect 392 1367 394 1393
rect 520 1367 522 1393
rect 664 1367 666 1393
rect 816 1367 818 1393
rect 968 1367 970 1393
rect 1120 1367 1122 1393
rect 1256 1367 1258 1393
rect 1392 1367 1394 1393
rect 1520 1367 1522 1393
rect 1648 1367 1650 1393
rect 1752 1367 1754 1393
rect 1832 1367 1834 1411
rect 1872 1375 1874 1411
rect 2254 1398 2260 1399
rect 2254 1394 2255 1398
rect 2259 1394 2260 1398
rect 2254 1393 2260 1394
rect 2350 1398 2356 1399
rect 2350 1394 2351 1398
rect 2355 1394 2356 1398
rect 2350 1393 2356 1394
rect 2462 1398 2468 1399
rect 2462 1394 2463 1398
rect 2467 1394 2468 1398
rect 2462 1393 2468 1394
rect 2582 1398 2588 1399
rect 2582 1394 2583 1398
rect 2587 1394 2588 1398
rect 2582 1393 2588 1394
rect 2710 1398 2716 1399
rect 2710 1394 2711 1398
rect 2715 1394 2716 1398
rect 2710 1393 2716 1394
rect 2838 1398 2844 1399
rect 2838 1394 2839 1398
rect 2843 1394 2844 1398
rect 2838 1393 2844 1394
rect 2958 1398 2964 1399
rect 2958 1394 2959 1398
rect 2963 1394 2964 1398
rect 2958 1393 2964 1394
rect 3078 1398 3084 1399
rect 3078 1394 3079 1398
rect 3083 1394 3084 1398
rect 3078 1393 3084 1394
rect 3190 1398 3196 1399
rect 3190 1394 3191 1398
rect 3195 1394 3196 1398
rect 3190 1393 3196 1394
rect 3302 1398 3308 1399
rect 3302 1394 3303 1398
rect 3307 1394 3308 1398
rect 3302 1393 3308 1394
rect 3414 1398 3420 1399
rect 3414 1394 3415 1398
rect 3419 1394 3420 1398
rect 3414 1393 3420 1394
rect 3510 1398 3516 1399
rect 3510 1394 3511 1398
rect 3515 1394 3516 1398
rect 3510 1393 3516 1394
rect 2256 1375 2258 1393
rect 2352 1375 2354 1393
rect 2464 1375 2466 1393
rect 2584 1375 2586 1393
rect 2712 1375 2714 1393
rect 2840 1375 2842 1393
rect 2960 1375 2962 1393
rect 3080 1375 3082 1393
rect 3192 1375 3194 1393
rect 3304 1375 3306 1393
rect 3416 1375 3418 1393
rect 3512 1375 3514 1393
rect 3592 1375 3594 1411
rect 1871 1374 1875 1375
rect 1871 1369 1875 1370
rect 2255 1374 2259 1375
rect 2255 1369 2259 1370
rect 2351 1374 2355 1375
rect 2351 1369 2355 1370
rect 2399 1374 2403 1375
rect 2399 1369 2403 1370
rect 2463 1374 2467 1375
rect 2463 1369 2467 1370
rect 2503 1374 2507 1375
rect 2503 1369 2507 1370
rect 2583 1374 2587 1375
rect 2583 1369 2587 1370
rect 2615 1374 2619 1375
rect 2615 1369 2619 1370
rect 2711 1374 2715 1375
rect 2711 1369 2715 1370
rect 2735 1374 2739 1375
rect 2735 1369 2739 1370
rect 2839 1374 2843 1375
rect 2839 1369 2843 1370
rect 2847 1374 2851 1375
rect 2847 1369 2851 1370
rect 2959 1374 2963 1375
rect 2959 1369 2963 1370
rect 3071 1374 3075 1375
rect 3071 1369 3075 1370
rect 3079 1374 3083 1375
rect 3079 1369 3083 1370
rect 3183 1374 3187 1375
rect 3183 1369 3187 1370
rect 3191 1374 3195 1375
rect 3191 1369 3195 1370
rect 3295 1374 3299 1375
rect 3295 1369 3299 1370
rect 3303 1374 3307 1375
rect 3303 1369 3307 1370
rect 3415 1374 3419 1375
rect 3415 1369 3419 1370
rect 3511 1374 3515 1375
rect 3511 1369 3515 1370
rect 3591 1374 3595 1375
rect 3591 1369 3595 1370
rect 111 1366 115 1367
rect 111 1361 115 1362
rect 223 1366 227 1367
rect 223 1361 227 1362
rect 287 1366 291 1367
rect 287 1361 291 1362
rect 335 1366 339 1367
rect 335 1361 339 1362
rect 391 1366 395 1367
rect 391 1361 395 1362
rect 471 1366 475 1367
rect 471 1361 475 1362
rect 519 1366 523 1367
rect 519 1361 523 1362
rect 623 1366 627 1367
rect 623 1361 627 1362
rect 663 1366 667 1367
rect 663 1361 667 1362
rect 783 1366 787 1367
rect 783 1361 787 1362
rect 815 1366 819 1367
rect 815 1361 819 1362
rect 943 1366 947 1367
rect 943 1361 947 1362
rect 967 1366 971 1367
rect 967 1361 971 1362
rect 1095 1366 1099 1367
rect 1095 1361 1099 1362
rect 1119 1366 1123 1367
rect 1119 1361 1123 1362
rect 1239 1366 1243 1367
rect 1239 1361 1243 1362
rect 1255 1366 1259 1367
rect 1255 1361 1259 1362
rect 1375 1366 1379 1367
rect 1375 1361 1379 1362
rect 1391 1366 1395 1367
rect 1391 1361 1395 1362
rect 1511 1366 1515 1367
rect 1511 1361 1515 1362
rect 1519 1366 1523 1367
rect 1519 1361 1523 1362
rect 1639 1366 1643 1367
rect 1639 1361 1643 1362
rect 1647 1366 1651 1367
rect 1647 1361 1651 1362
rect 1751 1366 1755 1367
rect 1751 1361 1755 1362
rect 1831 1366 1835 1367
rect 1831 1361 1835 1362
rect 112 1333 114 1361
rect 224 1351 226 1361
rect 336 1351 338 1361
rect 472 1351 474 1361
rect 624 1351 626 1361
rect 784 1351 786 1361
rect 944 1351 946 1361
rect 1096 1351 1098 1361
rect 1240 1351 1242 1361
rect 1376 1351 1378 1361
rect 1512 1351 1514 1361
rect 1640 1351 1642 1361
rect 1752 1351 1754 1361
rect 222 1350 228 1351
rect 222 1346 223 1350
rect 227 1346 228 1350
rect 222 1345 228 1346
rect 334 1350 340 1351
rect 334 1346 335 1350
rect 339 1346 340 1350
rect 334 1345 340 1346
rect 470 1350 476 1351
rect 470 1346 471 1350
rect 475 1346 476 1350
rect 470 1345 476 1346
rect 622 1350 628 1351
rect 622 1346 623 1350
rect 627 1346 628 1350
rect 622 1345 628 1346
rect 782 1350 788 1351
rect 782 1346 783 1350
rect 787 1346 788 1350
rect 782 1345 788 1346
rect 942 1350 948 1351
rect 942 1346 943 1350
rect 947 1346 948 1350
rect 942 1345 948 1346
rect 1094 1350 1100 1351
rect 1094 1346 1095 1350
rect 1099 1346 1100 1350
rect 1094 1345 1100 1346
rect 1238 1350 1244 1351
rect 1238 1346 1239 1350
rect 1243 1346 1244 1350
rect 1238 1345 1244 1346
rect 1374 1350 1380 1351
rect 1374 1346 1375 1350
rect 1379 1346 1380 1350
rect 1374 1345 1380 1346
rect 1510 1350 1516 1351
rect 1510 1346 1511 1350
rect 1515 1346 1516 1350
rect 1510 1345 1516 1346
rect 1638 1350 1644 1351
rect 1638 1346 1639 1350
rect 1643 1346 1644 1350
rect 1638 1345 1644 1346
rect 1750 1350 1756 1351
rect 1750 1346 1751 1350
rect 1755 1346 1756 1350
rect 1750 1345 1756 1346
rect 1832 1333 1834 1361
rect 1872 1341 1874 1369
rect 2400 1359 2402 1369
rect 2504 1359 2506 1369
rect 2616 1359 2618 1369
rect 2736 1359 2738 1369
rect 2848 1359 2850 1369
rect 2960 1359 2962 1369
rect 3072 1359 3074 1369
rect 3184 1359 3186 1369
rect 3296 1359 3298 1369
rect 3416 1359 3418 1369
rect 2398 1358 2404 1359
rect 2398 1354 2399 1358
rect 2403 1354 2404 1358
rect 2398 1353 2404 1354
rect 2502 1358 2508 1359
rect 2502 1354 2503 1358
rect 2507 1354 2508 1358
rect 2502 1353 2508 1354
rect 2614 1358 2620 1359
rect 2614 1354 2615 1358
rect 2619 1354 2620 1358
rect 2614 1353 2620 1354
rect 2734 1358 2740 1359
rect 2734 1354 2735 1358
rect 2739 1354 2740 1358
rect 2734 1353 2740 1354
rect 2846 1358 2852 1359
rect 2846 1354 2847 1358
rect 2851 1354 2852 1358
rect 2846 1353 2852 1354
rect 2958 1358 2964 1359
rect 2958 1354 2959 1358
rect 2963 1354 2964 1358
rect 2958 1353 2964 1354
rect 3070 1358 3076 1359
rect 3070 1354 3071 1358
rect 3075 1354 3076 1358
rect 3070 1353 3076 1354
rect 3182 1358 3188 1359
rect 3182 1354 3183 1358
rect 3187 1354 3188 1358
rect 3182 1353 3188 1354
rect 3294 1358 3300 1359
rect 3294 1354 3295 1358
rect 3299 1354 3300 1358
rect 3294 1353 3300 1354
rect 3414 1358 3420 1359
rect 3414 1354 3415 1358
rect 3419 1354 3420 1358
rect 3414 1353 3420 1354
rect 3592 1341 3594 1369
rect 1870 1340 1876 1341
rect 1870 1336 1871 1340
rect 1875 1336 1876 1340
rect 1870 1335 1876 1336
rect 3590 1340 3596 1341
rect 3590 1336 3591 1340
rect 3595 1336 3596 1340
rect 3590 1335 3596 1336
rect 110 1332 116 1333
rect 110 1328 111 1332
rect 115 1328 116 1332
rect 110 1327 116 1328
rect 1830 1332 1836 1333
rect 1830 1328 1831 1332
rect 1835 1328 1836 1332
rect 1830 1327 1836 1328
rect 1870 1323 1876 1324
rect 1870 1319 1871 1323
rect 1875 1319 1876 1323
rect 3590 1323 3596 1324
rect 1870 1318 1876 1319
rect 2390 1320 2396 1321
rect 110 1315 116 1316
rect 110 1311 111 1315
rect 115 1311 116 1315
rect 1830 1315 1836 1316
rect 110 1310 116 1311
rect 214 1312 220 1313
rect 112 1291 114 1310
rect 214 1308 215 1312
rect 219 1308 220 1312
rect 214 1307 220 1308
rect 326 1312 332 1313
rect 326 1308 327 1312
rect 331 1308 332 1312
rect 326 1307 332 1308
rect 462 1312 468 1313
rect 462 1308 463 1312
rect 467 1308 468 1312
rect 462 1307 468 1308
rect 614 1312 620 1313
rect 614 1308 615 1312
rect 619 1308 620 1312
rect 614 1307 620 1308
rect 774 1312 780 1313
rect 774 1308 775 1312
rect 779 1308 780 1312
rect 774 1307 780 1308
rect 934 1312 940 1313
rect 934 1308 935 1312
rect 939 1308 940 1312
rect 934 1307 940 1308
rect 1086 1312 1092 1313
rect 1086 1308 1087 1312
rect 1091 1308 1092 1312
rect 1086 1307 1092 1308
rect 1230 1312 1236 1313
rect 1230 1308 1231 1312
rect 1235 1308 1236 1312
rect 1230 1307 1236 1308
rect 1366 1312 1372 1313
rect 1366 1308 1367 1312
rect 1371 1308 1372 1312
rect 1366 1307 1372 1308
rect 1502 1312 1508 1313
rect 1502 1308 1503 1312
rect 1507 1308 1508 1312
rect 1502 1307 1508 1308
rect 1630 1312 1636 1313
rect 1630 1308 1631 1312
rect 1635 1308 1636 1312
rect 1630 1307 1636 1308
rect 1742 1312 1748 1313
rect 1742 1308 1743 1312
rect 1747 1308 1748 1312
rect 1830 1311 1831 1315
rect 1835 1311 1836 1315
rect 1830 1310 1836 1311
rect 1742 1307 1748 1308
rect 216 1291 218 1307
rect 328 1291 330 1307
rect 464 1291 466 1307
rect 616 1291 618 1307
rect 776 1291 778 1307
rect 936 1291 938 1307
rect 1088 1291 1090 1307
rect 1232 1291 1234 1307
rect 1368 1291 1370 1307
rect 1504 1291 1506 1307
rect 1632 1291 1634 1307
rect 1744 1291 1746 1307
rect 1832 1291 1834 1310
rect 111 1290 115 1291
rect 111 1285 115 1286
rect 135 1290 139 1291
rect 135 1285 139 1286
rect 215 1290 219 1291
rect 215 1285 219 1286
rect 327 1290 331 1291
rect 327 1285 331 1286
rect 335 1290 339 1291
rect 335 1285 339 1286
rect 463 1290 467 1291
rect 463 1285 467 1286
rect 607 1290 611 1291
rect 607 1285 611 1286
rect 615 1290 619 1291
rect 615 1285 619 1286
rect 751 1290 755 1291
rect 751 1285 755 1286
rect 775 1290 779 1291
rect 775 1285 779 1286
rect 903 1290 907 1291
rect 903 1285 907 1286
rect 935 1290 939 1291
rect 935 1285 939 1286
rect 1047 1290 1051 1291
rect 1047 1285 1051 1286
rect 1087 1290 1091 1291
rect 1087 1285 1091 1286
rect 1183 1290 1187 1291
rect 1183 1285 1187 1286
rect 1231 1290 1235 1291
rect 1231 1285 1235 1286
rect 1303 1290 1307 1291
rect 1303 1285 1307 1286
rect 1367 1290 1371 1291
rect 1367 1285 1371 1286
rect 1423 1290 1427 1291
rect 1423 1285 1427 1286
rect 1503 1290 1507 1291
rect 1503 1285 1507 1286
rect 1535 1290 1539 1291
rect 1535 1285 1539 1286
rect 1631 1290 1635 1291
rect 1631 1285 1635 1286
rect 1647 1290 1651 1291
rect 1647 1285 1651 1286
rect 1743 1290 1747 1291
rect 1743 1285 1747 1286
rect 1831 1290 1835 1291
rect 1831 1285 1835 1286
rect 112 1266 114 1285
rect 136 1269 138 1285
rect 216 1269 218 1285
rect 336 1269 338 1285
rect 464 1269 466 1285
rect 608 1269 610 1285
rect 752 1269 754 1285
rect 904 1269 906 1285
rect 1048 1269 1050 1285
rect 1184 1269 1186 1285
rect 1304 1269 1306 1285
rect 1424 1269 1426 1285
rect 1536 1269 1538 1285
rect 1648 1269 1650 1285
rect 1744 1269 1746 1285
rect 134 1268 140 1269
rect 110 1265 116 1266
rect 110 1261 111 1265
rect 115 1261 116 1265
rect 134 1264 135 1268
rect 139 1264 140 1268
rect 134 1263 140 1264
rect 214 1268 220 1269
rect 214 1264 215 1268
rect 219 1264 220 1268
rect 214 1263 220 1264
rect 334 1268 340 1269
rect 334 1264 335 1268
rect 339 1264 340 1268
rect 334 1263 340 1264
rect 462 1268 468 1269
rect 462 1264 463 1268
rect 467 1264 468 1268
rect 462 1263 468 1264
rect 606 1268 612 1269
rect 606 1264 607 1268
rect 611 1264 612 1268
rect 606 1263 612 1264
rect 750 1268 756 1269
rect 750 1264 751 1268
rect 755 1264 756 1268
rect 750 1263 756 1264
rect 902 1268 908 1269
rect 902 1264 903 1268
rect 907 1264 908 1268
rect 902 1263 908 1264
rect 1046 1268 1052 1269
rect 1046 1264 1047 1268
rect 1051 1264 1052 1268
rect 1046 1263 1052 1264
rect 1182 1268 1188 1269
rect 1182 1264 1183 1268
rect 1187 1264 1188 1268
rect 1182 1263 1188 1264
rect 1302 1268 1308 1269
rect 1302 1264 1303 1268
rect 1307 1264 1308 1268
rect 1302 1263 1308 1264
rect 1422 1268 1428 1269
rect 1422 1264 1423 1268
rect 1427 1264 1428 1268
rect 1422 1263 1428 1264
rect 1534 1268 1540 1269
rect 1534 1264 1535 1268
rect 1539 1264 1540 1268
rect 1534 1263 1540 1264
rect 1646 1268 1652 1269
rect 1646 1264 1647 1268
rect 1651 1264 1652 1268
rect 1646 1263 1652 1264
rect 1742 1268 1748 1269
rect 1742 1264 1743 1268
rect 1747 1264 1748 1268
rect 1832 1266 1834 1285
rect 1872 1283 1874 1318
rect 2390 1316 2391 1320
rect 2395 1316 2396 1320
rect 2390 1315 2396 1316
rect 2494 1320 2500 1321
rect 2494 1316 2495 1320
rect 2499 1316 2500 1320
rect 2494 1315 2500 1316
rect 2606 1320 2612 1321
rect 2606 1316 2607 1320
rect 2611 1316 2612 1320
rect 2606 1315 2612 1316
rect 2726 1320 2732 1321
rect 2726 1316 2727 1320
rect 2731 1316 2732 1320
rect 2726 1315 2732 1316
rect 2838 1320 2844 1321
rect 2838 1316 2839 1320
rect 2843 1316 2844 1320
rect 2838 1315 2844 1316
rect 2950 1320 2956 1321
rect 2950 1316 2951 1320
rect 2955 1316 2956 1320
rect 2950 1315 2956 1316
rect 3062 1320 3068 1321
rect 3062 1316 3063 1320
rect 3067 1316 3068 1320
rect 3062 1315 3068 1316
rect 3174 1320 3180 1321
rect 3174 1316 3175 1320
rect 3179 1316 3180 1320
rect 3174 1315 3180 1316
rect 3286 1320 3292 1321
rect 3286 1316 3287 1320
rect 3291 1316 3292 1320
rect 3286 1315 3292 1316
rect 3406 1320 3412 1321
rect 3406 1316 3407 1320
rect 3411 1316 3412 1320
rect 3590 1319 3591 1323
rect 3595 1319 3596 1323
rect 3590 1318 3596 1319
rect 3406 1315 3412 1316
rect 2392 1283 2394 1315
rect 2496 1283 2498 1315
rect 2608 1283 2610 1315
rect 2728 1283 2730 1315
rect 2840 1283 2842 1315
rect 2952 1283 2954 1315
rect 3064 1283 3066 1315
rect 3176 1283 3178 1315
rect 3288 1283 3290 1315
rect 3408 1283 3410 1315
rect 3592 1283 3594 1318
rect 1871 1282 1875 1283
rect 1871 1277 1875 1278
rect 1895 1282 1899 1283
rect 1895 1277 1899 1278
rect 2071 1282 2075 1283
rect 2071 1277 2075 1278
rect 2255 1282 2259 1283
rect 2255 1277 2259 1278
rect 2391 1282 2395 1283
rect 2391 1277 2395 1278
rect 2423 1282 2427 1283
rect 2423 1277 2427 1278
rect 2495 1282 2499 1283
rect 2495 1277 2499 1278
rect 2583 1282 2587 1283
rect 2583 1277 2587 1278
rect 2607 1282 2611 1283
rect 2607 1277 2611 1278
rect 2727 1282 2731 1283
rect 2727 1277 2731 1278
rect 2735 1282 2739 1283
rect 2735 1277 2739 1278
rect 2839 1282 2843 1283
rect 2839 1277 2843 1278
rect 2879 1282 2883 1283
rect 2879 1277 2883 1278
rect 2951 1282 2955 1283
rect 2951 1277 2955 1278
rect 3015 1282 3019 1283
rect 3015 1277 3019 1278
rect 3063 1282 3067 1283
rect 3063 1277 3067 1278
rect 3143 1282 3147 1283
rect 3143 1277 3147 1278
rect 3175 1282 3179 1283
rect 3175 1277 3179 1278
rect 3271 1282 3275 1283
rect 3271 1277 3275 1278
rect 3287 1282 3291 1283
rect 3287 1277 3291 1278
rect 3399 1282 3403 1283
rect 3399 1277 3403 1278
rect 3407 1282 3411 1283
rect 3407 1277 3411 1278
rect 3503 1282 3507 1283
rect 3503 1277 3507 1278
rect 3591 1282 3595 1283
rect 3591 1277 3595 1278
rect 1742 1263 1748 1264
rect 1830 1265 1836 1266
rect 110 1260 116 1261
rect 1830 1261 1831 1265
rect 1835 1261 1836 1265
rect 1830 1260 1836 1261
rect 1872 1258 1874 1277
rect 1896 1261 1898 1277
rect 2072 1261 2074 1277
rect 2256 1261 2258 1277
rect 2424 1261 2426 1277
rect 2584 1261 2586 1277
rect 2736 1261 2738 1277
rect 2880 1261 2882 1277
rect 3016 1261 3018 1277
rect 3144 1261 3146 1277
rect 3272 1261 3274 1277
rect 3400 1261 3402 1277
rect 3504 1261 3506 1277
rect 1894 1260 1900 1261
rect 1870 1257 1876 1258
rect 1870 1253 1871 1257
rect 1875 1253 1876 1257
rect 1894 1256 1895 1260
rect 1899 1256 1900 1260
rect 1894 1255 1900 1256
rect 2070 1260 2076 1261
rect 2070 1256 2071 1260
rect 2075 1256 2076 1260
rect 2070 1255 2076 1256
rect 2254 1260 2260 1261
rect 2254 1256 2255 1260
rect 2259 1256 2260 1260
rect 2254 1255 2260 1256
rect 2422 1260 2428 1261
rect 2422 1256 2423 1260
rect 2427 1256 2428 1260
rect 2422 1255 2428 1256
rect 2582 1260 2588 1261
rect 2582 1256 2583 1260
rect 2587 1256 2588 1260
rect 2582 1255 2588 1256
rect 2734 1260 2740 1261
rect 2734 1256 2735 1260
rect 2739 1256 2740 1260
rect 2734 1255 2740 1256
rect 2878 1260 2884 1261
rect 2878 1256 2879 1260
rect 2883 1256 2884 1260
rect 2878 1255 2884 1256
rect 3014 1260 3020 1261
rect 3014 1256 3015 1260
rect 3019 1256 3020 1260
rect 3014 1255 3020 1256
rect 3142 1260 3148 1261
rect 3142 1256 3143 1260
rect 3147 1256 3148 1260
rect 3142 1255 3148 1256
rect 3270 1260 3276 1261
rect 3270 1256 3271 1260
rect 3275 1256 3276 1260
rect 3270 1255 3276 1256
rect 3398 1260 3404 1261
rect 3398 1256 3399 1260
rect 3403 1256 3404 1260
rect 3398 1255 3404 1256
rect 3502 1260 3508 1261
rect 3502 1256 3503 1260
rect 3507 1256 3508 1260
rect 3592 1258 3594 1277
rect 3502 1255 3508 1256
rect 3590 1257 3596 1258
rect 1870 1252 1876 1253
rect 3590 1253 3591 1257
rect 3595 1253 3596 1257
rect 3590 1252 3596 1253
rect 110 1248 116 1249
rect 110 1244 111 1248
rect 115 1244 116 1248
rect 110 1243 116 1244
rect 1830 1248 1836 1249
rect 1830 1244 1831 1248
rect 1835 1244 1836 1248
rect 1830 1243 1836 1244
rect 112 1203 114 1243
rect 142 1230 148 1231
rect 142 1226 143 1230
rect 147 1226 148 1230
rect 142 1225 148 1226
rect 222 1230 228 1231
rect 222 1226 223 1230
rect 227 1226 228 1230
rect 222 1225 228 1226
rect 342 1230 348 1231
rect 342 1226 343 1230
rect 347 1226 348 1230
rect 342 1225 348 1226
rect 470 1230 476 1231
rect 470 1226 471 1230
rect 475 1226 476 1230
rect 470 1225 476 1226
rect 614 1230 620 1231
rect 614 1226 615 1230
rect 619 1226 620 1230
rect 614 1225 620 1226
rect 758 1230 764 1231
rect 758 1226 759 1230
rect 763 1226 764 1230
rect 758 1225 764 1226
rect 910 1230 916 1231
rect 910 1226 911 1230
rect 915 1226 916 1230
rect 910 1225 916 1226
rect 1054 1230 1060 1231
rect 1054 1226 1055 1230
rect 1059 1226 1060 1230
rect 1054 1225 1060 1226
rect 1190 1230 1196 1231
rect 1190 1226 1191 1230
rect 1195 1226 1196 1230
rect 1190 1225 1196 1226
rect 1310 1230 1316 1231
rect 1310 1226 1311 1230
rect 1315 1226 1316 1230
rect 1310 1225 1316 1226
rect 1430 1230 1436 1231
rect 1430 1226 1431 1230
rect 1435 1226 1436 1230
rect 1430 1225 1436 1226
rect 1542 1230 1548 1231
rect 1542 1226 1543 1230
rect 1547 1226 1548 1230
rect 1542 1225 1548 1226
rect 1654 1230 1660 1231
rect 1654 1226 1655 1230
rect 1659 1226 1660 1230
rect 1654 1225 1660 1226
rect 1750 1230 1756 1231
rect 1750 1226 1751 1230
rect 1755 1226 1756 1230
rect 1750 1225 1756 1226
rect 144 1203 146 1225
rect 224 1203 226 1225
rect 344 1203 346 1225
rect 472 1203 474 1225
rect 616 1203 618 1225
rect 760 1203 762 1225
rect 912 1203 914 1225
rect 1056 1203 1058 1225
rect 1192 1203 1194 1225
rect 1312 1203 1314 1225
rect 1432 1203 1434 1225
rect 1544 1203 1546 1225
rect 1656 1203 1658 1225
rect 1752 1203 1754 1225
rect 1832 1203 1834 1243
rect 1870 1240 1876 1241
rect 1870 1236 1871 1240
rect 1875 1236 1876 1240
rect 1870 1235 1876 1236
rect 3590 1240 3596 1241
rect 3590 1236 3591 1240
rect 3595 1236 3596 1240
rect 3590 1235 3596 1236
rect 111 1202 115 1203
rect 111 1197 115 1198
rect 143 1202 147 1203
rect 143 1197 147 1198
rect 223 1202 227 1203
rect 223 1197 227 1198
rect 255 1202 259 1203
rect 255 1197 259 1198
rect 343 1202 347 1203
rect 343 1197 347 1198
rect 383 1202 387 1203
rect 383 1197 387 1198
rect 471 1202 475 1203
rect 471 1197 475 1198
rect 503 1202 507 1203
rect 503 1197 507 1198
rect 615 1202 619 1203
rect 615 1197 619 1198
rect 719 1202 723 1203
rect 719 1197 723 1198
rect 759 1202 763 1203
rect 759 1197 763 1198
rect 815 1202 819 1203
rect 815 1197 819 1198
rect 911 1202 915 1203
rect 911 1197 915 1198
rect 999 1202 1003 1203
rect 999 1197 1003 1198
rect 1055 1202 1059 1203
rect 1055 1197 1059 1198
rect 1095 1202 1099 1203
rect 1095 1197 1099 1198
rect 1191 1202 1195 1203
rect 1191 1197 1195 1198
rect 1287 1202 1291 1203
rect 1287 1197 1291 1198
rect 1311 1202 1315 1203
rect 1311 1197 1315 1198
rect 1431 1202 1435 1203
rect 1431 1197 1435 1198
rect 1543 1202 1547 1203
rect 1543 1197 1547 1198
rect 1655 1202 1659 1203
rect 1655 1197 1659 1198
rect 1751 1202 1755 1203
rect 1751 1197 1755 1198
rect 1831 1202 1835 1203
rect 1872 1199 1874 1235
rect 1902 1222 1908 1223
rect 1902 1218 1903 1222
rect 1907 1218 1908 1222
rect 1902 1217 1908 1218
rect 2078 1222 2084 1223
rect 2078 1218 2079 1222
rect 2083 1218 2084 1222
rect 2078 1217 2084 1218
rect 2262 1222 2268 1223
rect 2262 1218 2263 1222
rect 2267 1218 2268 1222
rect 2262 1217 2268 1218
rect 2430 1222 2436 1223
rect 2430 1218 2431 1222
rect 2435 1218 2436 1222
rect 2430 1217 2436 1218
rect 2590 1222 2596 1223
rect 2590 1218 2591 1222
rect 2595 1218 2596 1222
rect 2590 1217 2596 1218
rect 2742 1222 2748 1223
rect 2742 1218 2743 1222
rect 2747 1218 2748 1222
rect 2742 1217 2748 1218
rect 2886 1222 2892 1223
rect 2886 1218 2887 1222
rect 2891 1218 2892 1222
rect 2886 1217 2892 1218
rect 3022 1222 3028 1223
rect 3022 1218 3023 1222
rect 3027 1218 3028 1222
rect 3022 1217 3028 1218
rect 3150 1222 3156 1223
rect 3150 1218 3151 1222
rect 3155 1218 3156 1222
rect 3150 1217 3156 1218
rect 3278 1222 3284 1223
rect 3278 1218 3279 1222
rect 3283 1218 3284 1222
rect 3278 1217 3284 1218
rect 3406 1222 3412 1223
rect 3406 1218 3407 1222
rect 3411 1218 3412 1222
rect 3406 1217 3412 1218
rect 3510 1222 3516 1223
rect 3510 1218 3511 1222
rect 3515 1218 3516 1222
rect 3510 1217 3516 1218
rect 1904 1199 1906 1217
rect 2080 1199 2082 1217
rect 2264 1199 2266 1217
rect 2432 1199 2434 1217
rect 2592 1199 2594 1217
rect 2744 1199 2746 1217
rect 2888 1199 2890 1217
rect 3024 1199 3026 1217
rect 3152 1199 3154 1217
rect 3280 1199 3282 1217
rect 3408 1199 3410 1217
rect 3512 1199 3514 1217
rect 3592 1199 3594 1235
rect 1831 1197 1835 1198
rect 1871 1198 1875 1199
rect 112 1169 114 1197
rect 144 1187 146 1197
rect 256 1187 258 1197
rect 384 1187 386 1197
rect 504 1187 506 1197
rect 616 1187 618 1197
rect 720 1187 722 1197
rect 816 1187 818 1197
rect 912 1187 914 1197
rect 1000 1187 1002 1197
rect 1096 1187 1098 1197
rect 1192 1187 1194 1197
rect 1288 1187 1290 1197
rect 142 1186 148 1187
rect 142 1182 143 1186
rect 147 1182 148 1186
rect 142 1181 148 1182
rect 254 1186 260 1187
rect 254 1182 255 1186
rect 259 1182 260 1186
rect 254 1181 260 1182
rect 382 1186 388 1187
rect 382 1182 383 1186
rect 387 1182 388 1186
rect 382 1181 388 1182
rect 502 1186 508 1187
rect 502 1182 503 1186
rect 507 1182 508 1186
rect 502 1181 508 1182
rect 614 1186 620 1187
rect 614 1182 615 1186
rect 619 1182 620 1186
rect 614 1181 620 1182
rect 718 1186 724 1187
rect 718 1182 719 1186
rect 723 1182 724 1186
rect 718 1181 724 1182
rect 814 1186 820 1187
rect 814 1182 815 1186
rect 819 1182 820 1186
rect 814 1181 820 1182
rect 910 1186 916 1187
rect 910 1182 911 1186
rect 915 1182 916 1186
rect 910 1181 916 1182
rect 998 1186 1004 1187
rect 998 1182 999 1186
rect 1003 1182 1004 1186
rect 998 1181 1004 1182
rect 1094 1186 1100 1187
rect 1094 1182 1095 1186
rect 1099 1182 1100 1186
rect 1094 1181 1100 1182
rect 1190 1186 1196 1187
rect 1190 1182 1191 1186
rect 1195 1182 1196 1186
rect 1190 1181 1196 1182
rect 1286 1186 1292 1187
rect 1286 1182 1287 1186
rect 1291 1182 1292 1186
rect 1286 1181 1292 1182
rect 1832 1169 1834 1197
rect 1871 1193 1875 1194
rect 1903 1198 1907 1199
rect 1903 1193 1907 1194
rect 1991 1198 1995 1199
rect 1991 1193 1995 1194
rect 2079 1198 2083 1199
rect 2079 1193 2083 1194
rect 2103 1198 2107 1199
rect 2103 1193 2107 1194
rect 2215 1198 2219 1199
rect 2215 1193 2219 1194
rect 2263 1198 2267 1199
rect 2263 1193 2267 1194
rect 2327 1198 2331 1199
rect 2327 1193 2331 1194
rect 2431 1198 2435 1199
rect 2431 1193 2435 1194
rect 2447 1198 2451 1199
rect 2447 1193 2451 1194
rect 2575 1198 2579 1199
rect 2575 1193 2579 1194
rect 2591 1198 2595 1199
rect 2591 1193 2595 1194
rect 2719 1198 2723 1199
rect 2719 1193 2723 1194
rect 2743 1198 2747 1199
rect 2743 1193 2747 1194
rect 2871 1198 2875 1199
rect 2871 1193 2875 1194
rect 2887 1198 2891 1199
rect 2887 1193 2891 1194
rect 3023 1198 3027 1199
rect 3023 1193 3027 1194
rect 3031 1198 3035 1199
rect 3031 1193 3035 1194
rect 3151 1198 3155 1199
rect 3151 1193 3155 1194
rect 3191 1198 3195 1199
rect 3191 1193 3195 1194
rect 3279 1198 3283 1199
rect 3279 1193 3283 1194
rect 3359 1198 3363 1199
rect 3359 1193 3363 1194
rect 3407 1198 3411 1199
rect 3407 1193 3411 1194
rect 3511 1198 3515 1199
rect 3511 1193 3515 1194
rect 3591 1198 3595 1199
rect 3591 1193 3595 1194
rect 110 1168 116 1169
rect 110 1164 111 1168
rect 115 1164 116 1168
rect 110 1163 116 1164
rect 1830 1168 1836 1169
rect 1830 1164 1831 1168
rect 1835 1164 1836 1168
rect 1872 1165 1874 1193
rect 1904 1183 1906 1193
rect 1992 1183 1994 1193
rect 2104 1183 2106 1193
rect 2216 1183 2218 1193
rect 2328 1183 2330 1193
rect 2448 1183 2450 1193
rect 2576 1183 2578 1193
rect 2720 1183 2722 1193
rect 2872 1183 2874 1193
rect 3032 1183 3034 1193
rect 3192 1183 3194 1193
rect 3360 1183 3362 1193
rect 3512 1183 3514 1193
rect 1902 1182 1908 1183
rect 1902 1178 1903 1182
rect 1907 1178 1908 1182
rect 1902 1177 1908 1178
rect 1990 1182 1996 1183
rect 1990 1178 1991 1182
rect 1995 1178 1996 1182
rect 1990 1177 1996 1178
rect 2102 1182 2108 1183
rect 2102 1178 2103 1182
rect 2107 1178 2108 1182
rect 2102 1177 2108 1178
rect 2214 1182 2220 1183
rect 2214 1178 2215 1182
rect 2219 1178 2220 1182
rect 2214 1177 2220 1178
rect 2326 1182 2332 1183
rect 2326 1178 2327 1182
rect 2331 1178 2332 1182
rect 2326 1177 2332 1178
rect 2446 1182 2452 1183
rect 2446 1178 2447 1182
rect 2451 1178 2452 1182
rect 2446 1177 2452 1178
rect 2574 1182 2580 1183
rect 2574 1178 2575 1182
rect 2579 1178 2580 1182
rect 2574 1177 2580 1178
rect 2718 1182 2724 1183
rect 2718 1178 2719 1182
rect 2723 1178 2724 1182
rect 2718 1177 2724 1178
rect 2870 1182 2876 1183
rect 2870 1178 2871 1182
rect 2875 1178 2876 1182
rect 2870 1177 2876 1178
rect 3030 1182 3036 1183
rect 3030 1178 3031 1182
rect 3035 1178 3036 1182
rect 3030 1177 3036 1178
rect 3190 1182 3196 1183
rect 3190 1178 3191 1182
rect 3195 1178 3196 1182
rect 3190 1177 3196 1178
rect 3358 1182 3364 1183
rect 3358 1178 3359 1182
rect 3363 1178 3364 1182
rect 3358 1177 3364 1178
rect 3510 1182 3516 1183
rect 3510 1178 3511 1182
rect 3515 1178 3516 1182
rect 3510 1177 3516 1178
rect 3592 1165 3594 1193
rect 1830 1163 1836 1164
rect 1870 1164 1876 1165
rect 1870 1160 1871 1164
rect 1875 1160 1876 1164
rect 1870 1159 1876 1160
rect 3590 1164 3596 1165
rect 3590 1160 3591 1164
rect 3595 1160 3596 1164
rect 3590 1159 3596 1160
rect 110 1151 116 1152
rect 110 1147 111 1151
rect 115 1147 116 1151
rect 1830 1151 1836 1152
rect 110 1146 116 1147
rect 134 1148 140 1149
rect 112 1115 114 1146
rect 134 1144 135 1148
rect 139 1144 140 1148
rect 134 1143 140 1144
rect 246 1148 252 1149
rect 246 1144 247 1148
rect 251 1144 252 1148
rect 246 1143 252 1144
rect 374 1148 380 1149
rect 374 1144 375 1148
rect 379 1144 380 1148
rect 374 1143 380 1144
rect 494 1148 500 1149
rect 494 1144 495 1148
rect 499 1144 500 1148
rect 494 1143 500 1144
rect 606 1148 612 1149
rect 606 1144 607 1148
rect 611 1144 612 1148
rect 606 1143 612 1144
rect 710 1148 716 1149
rect 710 1144 711 1148
rect 715 1144 716 1148
rect 710 1143 716 1144
rect 806 1148 812 1149
rect 806 1144 807 1148
rect 811 1144 812 1148
rect 806 1143 812 1144
rect 902 1148 908 1149
rect 902 1144 903 1148
rect 907 1144 908 1148
rect 902 1143 908 1144
rect 990 1148 996 1149
rect 990 1144 991 1148
rect 995 1144 996 1148
rect 990 1143 996 1144
rect 1086 1148 1092 1149
rect 1086 1144 1087 1148
rect 1091 1144 1092 1148
rect 1086 1143 1092 1144
rect 1182 1148 1188 1149
rect 1182 1144 1183 1148
rect 1187 1144 1188 1148
rect 1182 1143 1188 1144
rect 1278 1148 1284 1149
rect 1278 1144 1279 1148
rect 1283 1144 1284 1148
rect 1830 1147 1831 1151
rect 1835 1147 1836 1151
rect 1830 1146 1836 1147
rect 1870 1147 1876 1148
rect 1278 1143 1284 1144
rect 136 1115 138 1143
rect 248 1115 250 1143
rect 376 1115 378 1143
rect 496 1115 498 1143
rect 608 1115 610 1143
rect 712 1115 714 1143
rect 808 1115 810 1143
rect 904 1115 906 1143
rect 992 1115 994 1143
rect 1088 1115 1090 1143
rect 1184 1115 1186 1143
rect 1280 1115 1282 1143
rect 1832 1115 1834 1146
rect 1870 1143 1871 1147
rect 1875 1143 1876 1147
rect 3590 1147 3596 1148
rect 1870 1142 1876 1143
rect 1894 1144 1900 1145
rect 1872 1115 1874 1142
rect 1894 1140 1895 1144
rect 1899 1140 1900 1144
rect 1894 1139 1900 1140
rect 1982 1144 1988 1145
rect 1982 1140 1983 1144
rect 1987 1140 1988 1144
rect 1982 1139 1988 1140
rect 2094 1144 2100 1145
rect 2094 1140 2095 1144
rect 2099 1140 2100 1144
rect 2094 1139 2100 1140
rect 2206 1144 2212 1145
rect 2206 1140 2207 1144
rect 2211 1140 2212 1144
rect 2206 1139 2212 1140
rect 2318 1144 2324 1145
rect 2318 1140 2319 1144
rect 2323 1140 2324 1144
rect 2318 1139 2324 1140
rect 2438 1144 2444 1145
rect 2438 1140 2439 1144
rect 2443 1140 2444 1144
rect 2438 1139 2444 1140
rect 2566 1144 2572 1145
rect 2566 1140 2567 1144
rect 2571 1140 2572 1144
rect 2566 1139 2572 1140
rect 2710 1144 2716 1145
rect 2710 1140 2711 1144
rect 2715 1140 2716 1144
rect 2710 1139 2716 1140
rect 2862 1144 2868 1145
rect 2862 1140 2863 1144
rect 2867 1140 2868 1144
rect 2862 1139 2868 1140
rect 3022 1144 3028 1145
rect 3022 1140 3023 1144
rect 3027 1140 3028 1144
rect 3022 1139 3028 1140
rect 3182 1144 3188 1145
rect 3182 1140 3183 1144
rect 3187 1140 3188 1144
rect 3182 1139 3188 1140
rect 3350 1144 3356 1145
rect 3350 1140 3351 1144
rect 3355 1140 3356 1144
rect 3350 1139 3356 1140
rect 3502 1144 3508 1145
rect 3502 1140 3503 1144
rect 3507 1140 3508 1144
rect 3590 1143 3591 1147
rect 3595 1143 3596 1147
rect 3590 1142 3596 1143
rect 3502 1139 3508 1140
rect 1896 1115 1898 1139
rect 1984 1115 1986 1139
rect 2096 1115 2098 1139
rect 2208 1115 2210 1139
rect 2320 1115 2322 1139
rect 2440 1115 2442 1139
rect 2568 1115 2570 1139
rect 2712 1115 2714 1139
rect 2864 1115 2866 1139
rect 3024 1115 3026 1139
rect 3184 1115 3186 1139
rect 3352 1115 3354 1139
rect 3504 1115 3506 1139
rect 3592 1115 3594 1142
rect 111 1114 115 1115
rect 111 1109 115 1110
rect 135 1114 139 1115
rect 135 1109 139 1110
rect 247 1114 251 1115
rect 247 1109 251 1110
rect 255 1114 259 1115
rect 255 1109 259 1110
rect 375 1114 379 1115
rect 375 1109 379 1110
rect 399 1114 403 1115
rect 399 1109 403 1110
rect 495 1114 499 1115
rect 495 1109 499 1110
rect 535 1114 539 1115
rect 535 1109 539 1110
rect 607 1114 611 1115
rect 607 1109 611 1110
rect 663 1114 667 1115
rect 663 1109 667 1110
rect 711 1114 715 1115
rect 711 1109 715 1110
rect 783 1114 787 1115
rect 783 1109 787 1110
rect 807 1114 811 1115
rect 807 1109 811 1110
rect 895 1114 899 1115
rect 895 1109 899 1110
rect 903 1114 907 1115
rect 903 1109 907 1110
rect 991 1114 995 1115
rect 991 1109 995 1110
rect 999 1114 1003 1115
rect 999 1109 1003 1110
rect 1087 1114 1091 1115
rect 1087 1109 1091 1110
rect 1095 1114 1099 1115
rect 1095 1109 1099 1110
rect 1183 1114 1187 1115
rect 1183 1109 1187 1110
rect 1191 1114 1195 1115
rect 1191 1109 1195 1110
rect 1279 1114 1283 1115
rect 1279 1109 1283 1110
rect 1295 1114 1299 1115
rect 1295 1109 1299 1110
rect 1399 1114 1403 1115
rect 1399 1109 1403 1110
rect 1831 1114 1835 1115
rect 1831 1109 1835 1110
rect 1871 1114 1875 1115
rect 1871 1109 1875 1110
rect 1895 1114 1899 1115
rect 1895 1109 1899 1110
rect 1967 1114 1971 1115
rect 1967 1109 1971 1110
rect 1983 1114 1987 1115
rect 1983 1109 1987 1110
rect 2047 1114 2051 1115
rect 2047 1109 2051 1110
rect 2095 1114 2099 1115
rect 2095 1109 2099 1110
rect 2135 1114 2139 1115
rect 2135 1109 2139 1110
rect 2207 1114 2211 1115
rect 2207 1109 2211 1110
rect 2231 1114 2235 1115
rect 2231 1109 2235 1110
rect 2319 1114 2323 1115
rect 2319 1109 2323 1110
rect 2335 1114 2339 1115
rect 2335 1109 2339 1110
rect 2439 1114 2443 1115
rect 2439 1109 2443 1110
rect 2551 1114 2555 1115
rect 2551 1109 2555 1110
rect 2567 1114 2571 1115
rect 2567 1109 2571 1110
rect 2679 1114 2683 1115
rect 2679 1109 2683 1110
rect 2711 1114 2715 1115
rect 2711 1109 2715 1110
rect 2823 1114 2827 1115
rect 2823 1109 2827 1110
rect 2863 1114 2867 1115
rect 2863 1109 2867 1110
rect 2983 1114 2987 1115
rect 2983 1109 2987 1110
rect 3023 1114 3027 1115
rect 3023 1109 3027 1110
rect 3159 1114 3163 1115
rect 3159 1109 3163 1110
rect 3183 1114 3187 1115
rect 3183 1109 3187 1110
rect 3343 1114 3347 1115
rect 3343 1109 3347 1110
rect 3351 1114 3355 1115
rect 3351 1109 3355 1110
rect 3503 1114 3507 1115
rect 3503 1109 3507 1110
rect 3591 1114 3595 1115
rect 3591 1109 3595 1110
rect 112 1090 114 1109
rect 136 1093 138 1109
rect 256 1093 258 1109
rect 400 1093 402 1109
rect 536 1093 538 1109
rect 664 1093 666 1109
rect 784 1093 786 1109
rect 896 1093 898 1109
rect 1000 1093 1002 1109
rect 1096 1093 1098 1109
rect 1192 1093 1194 1109
rect 1296 1093 1298 1109
rect 1400 1093 1402 1109
rect 134 1092 140 1093
rect 110 1089 116 1090
rect 110 1085 111 1089
rect 115 1085 116 1089
rect 134 1088 135 1092
rect 139 1088 140 1092
rect 134 1087 140 1088
rect 254 1092 260 1093
rect 254 1088 255 1092
rect 259 1088 260 1092
rect 254 1087 260 1088
rect 398 1092 404 1093
rect 398 1088 399 1092
rect 403 1088 404 1092
rect 398 1087 404 1088
rect 534 1092 540 1093
rect 534 1088 535 1092
rect 539 1088 540 1092
rect 534 1087 540 1088
rect 662 1092 668 1093
rect 662 1088 663 1092
rect 667 1088 668 1092
rect 662 1087 668 1088
rect 782 1092 788 1093
rect 782 1088 783 1092
rect 787 1088 788 1092
rect 782 1087 788 1088
rect 894 1092 900 1093
rect 894 1088 895 1092
rect 899 1088 900 1092
rect 894 1087 900 1088
rect 998 1092 1004 1093
rect 998 1088 999 1092
rect 1003 1088 1004 1092
rect 998 1087 1004 1088
rect 1094 1092 1100 1093
rect 1094 1088 1095 1092
rect 1099 1088 1100 1092
rect 1094 1087 1100 1088
rect 1190 1092 1196 1093
rect 1190 1088 1191 1092
rect 1195 1088 1196 1092
rect 1190 1087 1196 1088
rect 1294 1092 1300 1093
rect 1294 1088 1295 1092
rect 1299 1088 1300 1092
rect 1294 1087 1300 1088
rect 1398 1092 1404 1093
rect 1398 1088 1399 1092
rect 1403 1088 1404 1092
rect 1832 1090 1834 1109
rect 1872 1090 1874 1109
rect 1968 1093 1970 1109
rect 2048 1093 2050 1109
rect 2136 1093 2138 1109
rect 2232 1093 2234 1109
rect 2336 1093 2338 1109
rect 2440 1093 2442 1109
rect 2552 1093 2554 1109
rect 2680 1093 2682 1109
rect 2824 1093 2826 1109
rect 2984 1093 2986 1109
rect 3160 1093 3162 1109
rect 3344 1093 3346 1109
rect 3504 1093 3506 1109
rect 1966 1092 1972 1093
rect 1398 1087 1404 1088
rect 1830 1089 1836 1090
rect 110 1084 116 1085
rect 1830 1085 1831 1089
rect 1835 1085 1836 1089
rect 1830 1084 1836 1085
rect 1870 1089 1876 1090
rect 1870 1085 1871 1089
rect 1875 1085 1876 1089
rect 1966 1088 1967 1092
rect 1971 1088 1972 1092
rect 1966 1087 1972 1088
rect 2046 1092 2052 1093
rect 2046 1088 2047 1092
rect 2051 1088 2052 1092
rect 2046 1087 2052 1088
rect 2134 1092 2140 1093
rect 2134 1088 2135 1092
rect 2139 1088 2140 1092
rect 2134 1087 2140 1088
rect 2230 1092 2236 1093
rect 2230 1088 2231 1092
rect 2235 1088 2236 1092
rect 2230 1087 2236 1088
rect 2334 1092 2340 1093
rect 2334 1088 2335 1092
rect 2339 1088 2340 1092
rect 2334 1087 2340 1088
rect 2438 1092 2444 1093
rect 2438 1088 2439 1092
rect 2443 1088 2444 1092
rect 2438 1087 2444 1088
rect 2550 1092 2556 1093
rect 2550 1088 2551 1092
rect 2555 1088 2556 1092
rect 2550 1087 2556 1088
rect 2678 1092 2684 1093
rect 2678 1088 2679 1092
rect 2683 1088 2684 1092
rect 2678 1087 2684 1088
rect 2822 1092 2828 1093
rect 2822 1088 2823 1092
rect 2827 1088 2828 1092
rect 2822 1087 2828 1088
rect 2982 1092 2988 1093
rect 2982 1088 2983 1092
rect 2987 1088 2988 1092
rect 2982 1087 2988 1088
rect 3158 1092 3164 1093
rect 3158 1088 3159 1092
rect 3163 1088 3164 1092
rect 3158 1087 3164 1088
rect 3342 1092 3348 1093
rect 3342 1088 3343 1092
rect 3347 1088 3348 1092
rect 3342 1087 3348 1088
rect 3502 1092 3508 1093
rect 3502 1088 3503 1092
rect 3507 1088 3508 1092
rect 3592 1090 3594 1109
rect 3502 1087 3508 1088
rect 3590 1089 3596 1090
rect 1870 1084 1876 1085
rect 3590 1085 3591 1089
rect 3595 1085 3596 1089
rect 3590 1084 3596 1085
rect 110 1072 116 1073
rect 110 1068 111 1072
rect 115 1068 116 1072
rect 110 1067 116 1068
rect 1830 1072 1836 1073
rect 1830 1068 1831 1072
rect 1835 1068 1836 1072
rect 1830 1067 1836 1068
rect 1870 1072 1876 1073
rect 1870 1068 1871 1072
rect 1875 1068 1876 1072
rect 1870 1067 1876 1068
rect 3590 1072 3596 1073
rect 3590 1068 3591 1072
rect 3595 1068 3596 1072
rect 3590 1067 3596 1068
rect 112 1031 114 1067
rect 142 1054 148 1055
rect 142 1050 143 1054
rect 147 1050 148 1054
rect 142 1049 148 1050
rect 262 1054 268 1055
rect 262 1050 263 1054
rect 267 1050 268 1054
rect 262 1049 268 1050
rect 406 1054 412 1055
rect 406 1050 407 1054
rect 411 1050 412 1054
rect 406 1049 412 1050
rect 542 1054 548 1055
rect 542 1050 543 1054
rect 547 1050 548 1054
rect 542 1049 548 1050
rect 670 1054 676 1055
rect 670 1050 671 1054
rect 675 1050 676 1054
rect 670 1049 676 1050
rect 790 1054 796 1055
rect 790 1050 791 1054
rect 795 1050 796 1054
rect 790 1049 796 1050
rect 902 1054 908 1055
rect 902 1050 903 1054
rect 907 1050 908 1054
rect 902 1049 908 1050
rect 1006 1054 1012 1055
rect 1006 1050 1007 1054
rect 1011 1050 1012 1054
rect 1006 1049 1012 1050
rect 1102 1054 1108 1055
rect 1102 1050 1103 1054
rect 1107 1050 1108 1054
rect 1102 1049 1108 1050
rect 1198 1054 1204 1055
rect 1198 1050 1199 1054
rect 1203 1050 1204 1054
rect 1198 1049 1204 1050
rect 1302 1054 1308 1055
rect 1302 1050 1303 1054
rect 1307 1050 1308 1054
rect 1302 1049 1308 1050
rect 1406 1054 1412 1055
rect 1406 1050 1407 1054
rect 1411 1050 1412 1054
rect 1406 1049 1412 1050
rect 144 1031 146 1049
rect 264 1031 266 1049
rect 408 1031 410 1049
rect 544 1031 546 1049
rect 672 1031 674 1049
rect 792 1031 794 1049
rect 904 1031 906 1049
rect 1008 1031 1010 1049
rect 1104 1031 1106 1049
rect 1200 1031 1202 1049
rect 1304 1031 1306 1049
rect 1408 1031 1410 1049
rect 1832 1031 1834 1067
rect 1872 1031 1874 1067
rect 1974 1054 1980 1055
rect 1974 1050 1975 1054
rect 1979 1050 1980 1054
rect 1974 1049 1980 1050
rect 2054 1054 2060 1055
rect 2054 1050 2055 1054
rect 2059 1050 2060 1054
rect 2054 1049 2060 1050
rect 2142 1054 2148 1055
rect 2142 1050 2143 1054
rect 2147 1050 2148 1054
rect 2142 1049 2148 1050
rect 2238 1054 2244 1055
rect 2238 1050 2239 1054
rect 2243 1050 2244 1054
rect 2238 1049 2244 1050
rect 2342 1054 2348 1055
rect 2342 1050 2343 1054
rect 2347 1050 2348 1054
rect 2342 1049 2348 1050
rect 2446 1054 2452 1055
rect 2446 1050 2447 1054
rect 2451 1050 2452 1054
rect 2446 1049 2452 1050
rect 2558 1054 2564 1055
rect 2558 1050 2559 1054
rect 2563 1050 2564 1054
rect 2558 1049 2564 1050
rect 2686 1054 2692 1055
rect 2686 1050 2687 1054
rect 2691 1050 2692 1054
rect 2686 1049 2692 1050
rect 2830 1054 2836 1055
rect 2830 1050 2831 1054
rect 2835 1050 2836 1054
rect 2830 1049 2836 1050
rect 2990 1054 2996 1055
rect 2990 1050 2991 1054
rect 2995 1050 2996 1054
rect 2990 1049 2996 1050
rect 3166 1054 3172 1055
rect 3166 1050 3167 1054
rect 3171 1050 3172 1054
rect 3166 1049 3172 1050
rect 3350 1054 3356 1055
rect 3350 1050 3351 1054
rect 3355 1050 3356 1054
rect 3350 1049 3356 1050
rect 3510 1054 3516 1055
rect 3510 1050 3511 1054
rect 3515 1050 3516 1054
rect 3510 1049 3516 1050
rect 1976 1031 1978 1049
rect 2056 1031 2058 1049
rect 2144 1031 2146 1049
rect 2240 1031 2242 1049
rect 2344 1031 2346 1049
rect 2448 1031 2450 1049
rect 2560 1031 2562 1049
rect 2688 1031 2690 1049
rect 2832 1031 2834 1049
rect 2992 1031 2994 1049
rect 3168 1031 3170 1049
rect 3352 1031 3354 1049
rect 3512 1031 3514 1049
rect 3592 1031 3594 1067
rect 111 1030 115 1031
rect 111 1025 115 1026
rect 143 1030 147 1031
rect 143 1025 147 1026
rect 263 1030 267 1031
rect 263 1025 267 1026
rect 271 1030 275 1031
rect 271 1025 275 1026
rect 407 1030 411 1031
rect 407 1025 411 1026
rect 423 1030 427 1031
rect 423 1025 427 1026
rect 543 1030 547 1031
rect 543 1025 547 1026
rect 583 1030 587 1031
rect 583 1025 587 1026
rect 671 1030 675 1031
rect 671 1025 675 1026
rect 735 1030 739 1031
rect 735 1025 739 1026
rect 791 1030 795 1031
rect 791 1025 795 1026
rect 887 1030 891 1031
rect 887 1025 891 1026
rect 903 1030 907 1031
rect 903 1025 907 1026
rect 1007 1030 1011 1031
rect 1007 1025 1011 1026
rect 1031 1030 1035 1031
rect 1031 1025 1035 1026
rect 1103 1030 1107 1031
rect 1103 1025 1107 1026
rect 1159 1030 1163 1031
rect 1159 1025 1163 1026
rect 1199 1030 1203 1031
rect 1199 1025 1203 1026
rect 1279 1030 1283 1031
rect 1279 1025 1283 1026
rect 1303 1030 1307 1031
rect 1303 1025 1307 1026
rect 1399 1030 1403 1031
rect 1399 1025 1403 1026
rect 1407 1030 1411 1031
rect 1407 1025 1411 1026
rect 1519 1030 1523 1031
rect 1519 1025 1523 1026
rect 1639 1030 1643 1031
rect 1639 1025 1643 1026
rect 1831 1030 1835 1031
rect 1831 1025 1835 1026
rect 1871 1030 1875 1031
rect 1871 1025 1875 1026
rect 1975 1030 1979 1031
rect 1975 1025 1979 1026
rect 2031 1030 2035 1031
rect 2031 1025 2035 1026
rect 2055 1030 2059 1031
rect 2055 1025 2059 1026
rect 2127 1030 2131 1031
rect 2127 1025 2131 1026
rect 2143 1030 2147 1031
rect 2143 1025 2147 1026
rect 2231 1030 2235 1031
rect 2231 1025 2235 1026
rect 2239 1030 2243 1031
rect 2239 1025 2243 1026
rect 2343 1030 2347 1031
rect 2343 1025 2347 1026
rect 2351 1030 2355 1031
rect 2351 1025 2355 1026
rect 2447 1030 2451 1031
rect 2447 1025 2451 1026
rect 2471 1030 2475 1031
rect 2471 1025 2475 1026
rect 2559 1030 2563 1031
rect 2559 1025 2563 1026
rect 2599 1030 2603 1031
rect 2599 1025 2603 1026
rect 2687 1030 2691 1031
rect 2687 1025 2691 1026
rect 2727 1030 2731 1031
rect 2727 1025 2731 1026
rect 2831 1030 2835 1031
rect 2831 1025 2835 1026
rect 2855 1030 2859 1031
rect 2855 1025 2859 1026
rect 2983 1030 2987 1031
rect 2983 1025 2987 1026
rect 2991 1030 2995 1031
rect 2991 1025 2995 1026
rect 3111 1030 3115 1031
rect 3111 1025 3115 1026
rect 3167 1030 3171 1031
rect 3167 1025 3171 1026
rect 3247 1030 3251 1031
rect 3247 1025 3251 1026
rect 3351 1030 3355 1031
rect 3351 1025 3355 1026
rect 3391 1030 3395 1031
rect 3391 1025 3395 1026
rect 3511 1030 3515 1031
rect 3511 1025 3515 1026
rect 3591 1030 3595 1031
rect 3591 1025 3595 1026
rect 112 997 114 1025
rect 144 1015 146 1025
rect 272 1015 274 1025
rect 424 1015 426 1025
rect 584 1015 586 1025
rect 736 1015 738 1025
rect 888 1015 890 1025
rect 1032 1015 1034 1025
rect 1160 1015 1162 1025
rect 1280 1015 1282 1025
rect 1400 1015 1402 1025
rect 1520 1015 1522 1025
rect 1640 1015 1642 1025
rect 142 1014 148 1015
rect 142 1010 143 1014
rect 147 1010 148 1014
rect 142 1009 148 1010
rect 270 1014 276 1015
rect 270 1010 271 1014
rect 275 1010 276 1014
rect 270 1009 276 1010
rect 422 1014 428 1015
rect 422 1010 423 1014
rect 427 1010 428 1014
rect 422 1009 428 1010
rect 582 1014 588 1015
rect 582 1010 583 1014
rect 587 1010 588 1014
rect 582 1009 588 1010
rect 734 1014 740 1015
rect 734 1010 735 1014
rect 739 1010 740 1014
rect 734 1009 740 1010
rect 886 1014 892 1015
rect 886 1010 887 1014
rect 891 1010 892 1014
rect 886 1009 892 1010
rect 1030 1014 1036 1015
rect 1030 1010 1031 1014
rect 1035 1010 1036 1014
rect 1030 1009 1036 1010
rect 1158 1014 1164 1015
rect 1158 1010 1159 1014
rect 1163 1010 1164 1014
rect 1158 1009 1164 1010
rect 1278 1014 1284 1015
rect 1278 1010 1279 1014
rect 1283 1010 1284 1014
rect 1278 1009 1284 1010
rect 1398 1014 1404 1015
rect 1398 1010 1399 1014
rect 1403 1010 1404 1014
rect 1398 1009 1404 1010
rect 1518 1014 1524 1015
rect 1518 1010 1519 1014
rect 1523 1010 1524 1014
rect 1518 1009 1524 1010
rect 1638 1014 1644 1015
rect 1638 1010 1639 1014
rect 1643 1010 1644 1014
rect 1638 1009 1644 1010
rect 1832 997 1834 1025
rect 1872 997 1874 1025
rect 2032 1015 2034 1025
rect 2128 1015 2130 1025
rect 2232 1015 2234 1025
rect 2352 1015 2354 1025
rect 2472 1015 2474 1025
rect 2600 1015 2602 1025
rect 2728 1015 2730 1025
rect 2856 1015 2858 1025
rect 2984 1015 2986 1025
rect 3112 1015 3114 1025
rect 3248 1015 3250 1025
rect 3392 1015 3394 1025
rect 3512 1015 3514 1025
rect 2030 1014 2036 1015
rect 2030 1010 2031 1014
rect 2035 1010 2036 1014
rect 2030 1009 2036 1010
rect 2126 1014 2132 1015
rect 2126 1010 2127 1014
rect 2131 1010 2132 1014
rect 2126 1009 2132 1010
rect 2230 1014 2236 1015
rect 2230 1010 2231 1014
rect 2235 1010 2236 1014
rect 2230 1009 2236 1010
rect 2350 1014 2356 1015
rect 2350 1010 2351 1014
rect 2355 1010 2356 1014
rect 2350 1009 2356 1010
rect 2470 1014 2476 1015
rect 2470 1010 2471 1014
rect 2475 1010 2476 1014
rect 2470 1009 2476 1010
rect 2598 1014 2604 1015
rect 2598 1010 2599 1014
rect 2603 1010 2604 1014
rect 2598 1009 2604 1010
rect 2726 1014 2732 1015
rect 2726 1010 2727 1014
rect 2731 1010 2732 1014
rect 2726 1009 2732 1010
rect 2854 1014 2860 1015
rect 2854 1010 2855 1014
rect 2859 1010 2860 1014
rect 2854 1009 2860 1010
rect 2982 1014 2988 1015
rect 2982 1010 2983 1014
rect 2987 1010 2988 1014
rect 2982 1009 2988 1010
rect 3110 1014 3116 1015
rect 3110 1010 3111 1014
rect 3115 1010 3116 1014
rect 3110 1009 3116 1010
rect 3246 1014 3252 1015
rect 3246 1010 3247 1014
rect 3251 1010 3252 1014
rect 3246 1009 3252 1010
rect 3390 1014 3396 1015
rect 3390 1010 3391 1014
rect 3395 1010 3396 1014
rect 3390 1009 3396 1010
rect 3510 1014 3516 1015
rect 3510 1010 3511 1014
rect 3515 1010 3516 1014
rect 3510 1009 3516 1010
rect 3592 997 3594 1025
rect 110 996 116 997
rect 110 992 111 996
rect 115 992 116 996
rect 110 991 116 992
rect 1830 996 1836 997
rect 1830 992 1831 996
rect 1835 992 1836 996
rect 1830 991 1836 992
rect 1870 996 1876 997
rect 1870 992 1871 996
rect 1875 992 1876 996
rect 1870 991 1876 992
rect 3590 996 3596 997
rect 3590 992 3591 996
rect 3595 992 3596 996
rect 3590 991 3596 992
rect 110 979 116 980
rect 110 975 111 979
rect 115 975 116 979
rect 1830 979 1836 980
rect 110 974 116 975
rect 134 976 140 977
rect 112 947 114 974
rect 134 972 135 976
rect 139 972 140 976
rect 134 971 140 972
rect 262 976 268 977
rect 262 972 263 976
rect 267 972 268 976
rect 262 971 268 972
rect 414 976 420 977
rect 414 972 415 976
rect 419 972 420 976
rect 414 971 420 972
rect 574 976 580 977
rect 574 972 575 976
rect 579 972 580 976
rect 574 971 580 972
rect 726 976 732 977
rect 726 972 727 976
rect 731 972 732 976
rect 726 971 732 972
rect 878 976 884 977
rect 878 972 879 976
rect 883 972 884 976
rect 878 971 884 972
rect 1022 976 1028 977
rect 1022 972 1023 976
rect 1027 972 1028 976
rect 1022 971 1028 972
rect 1150 976 1156 977
rect 1150 972 1151 976
rect 1155 972 1156 976
rect 1150 971 1156 972
rect 1270 976 1276 977
rect 1270 972 1271 976
rect 1275 972 1276 976
rect 1270 971 1276 972
rect 1390 976 1396 977
rect 1390 972 1391 976
rect 1395 972 1396 976
rect 1390 971 1396 972
rect 1510 976 1516 977
rect 1510 972 1511 976
rect 1515 972 1516 976
rect 1510 971 1516 972
rect 1630 976 1636 977
rect 1630 972 1631 976
rect 1635 972 1636 976
rect 1830 975 1831 979
rect 1835 975 1836 979
rect 1830 974 1836 975
rect 1870 979 1876 980
rect 1870 975 1871 979
rect 1875 975 1876 979
rect 3590 979 3596 980
rect 1870 974 1876 975
rect 2022 976 2028 977
rect 1630 971 1636 972
rect 136 947 138 971
rect 264 947 266 971
rect 416 947 418 971
rect 576 947 578 971
rect 728 947 730 971
rect 880 947 882 971
rect 1024 947 1026 971
rect 1152 947 1154 971
rect 1272 947 1274 971
rect 1392 947 1394 971
rect 1512 947 1514 971
rect 1632 947 1634 971
rect 1832 947 1834 974
rect 1872 947 1874 974
rect 2022 972 2023 976
rect 2027 972 2028 976
rect 2022 971 2028 972
rect 2118 976 2124 977
rect 2118 972 2119 976
rect 2123 972 2124 976
rect 2118 971 2124 972
rect 2222 976 2228 977
rect 2222 972 2223 976
rect 2227 972 2228 976
rect 2222 971 2228 972
rect 2342 976 2348 977
rect 2342 972 2343 976
rect 2347 972 2348 976
rect 2342 971 2348 972
rect 2462 976 2468 977
rect 2462 972 2463 976
rect 2467 972 2468 976
rect 2462 971 2468 972
rect 2590 976 2596 977
rect 2590 972 2591 976
rect 2595 972 2596 976
rect 2590 971 2596 972
rect 2718 976 2724 977
rect 2718 972 2719 976
rect 2723 972 2724 976
rect 2718 971 2724 972
rect 2846 976 2852 977
rect 2846 972 2847 976
rect 2851 972 2852 976
rect 2846 971 2852 972
rect 2974 976 2980 977
rect 2974 972 2975 976
rect 2979 972 2980 976
rect 2974 971 2980 972
rect 3102 976 3108 977
rect 3102 972 3103 976
rect 3107 972 3108 976
rect 3102 971 3108 972
rect 3238 976 3244 977
rect 3238 972 3239 976
rect 3243 972 3244 976
rect 3238 971 3244 972
rect 3382 976 3388 977
rect 3382 972 3383 976
rect 3387 972 3388 976
rect 3382 971 3388 972
rect 3502 976 3508 977
rect 3502 972 3503 976
rect 3507 972 3508 976
rect 3590 975 3591 979
rect 3595 975 3596 979
rect 3590 974 3596 975
rect 3502 971 3508 972
rect 2024 947 2026 971
rect 2120 947 2122 971
rect 2224 947 2226 971
rect 2344 947 2346 971
rect 2464 947 2466 971
rect 2592 947 2594 971
rect 2720 947 2722 971
rect 2848 947 2850 971
rect 2976 947 2978 971
rect 3104 947 3106 971
rect 3240 947 3242 971
rect 3384 947 3386 971
rect 3504 947 3506 971
rect 3592 947 3594 974
rect 111 946 115 947
rect 111 941 115 942
rect 135 946 139 947
rect 135 941 139 942
rect 215 946 219 947
rect 215 941 219 942
rect 263 946 267 947
rect 263 941 267 942
rect 335 946 339 947
rect 335 941 339 942
rect 415 946 419 947
rect 415 941 419 942
rect 463 946 467 947
rect 463 941 467 942
rect 575 946 579 947
rect 575 941 579 942
rect 599 946 603 947
rect 599 941 603 942
rect 727 946 731 947
rect 727 941 731 942
rect 735 946 739 947
rect 735 941 739 942
rect 863 946 867 947
rect 863 941 867 942
rect 879 946 883 947
rect 879 941 883 942
rect 991 946 995 947
rect 991 941 995 942
rect 1023 946 1027 947
rect 1023 941 1027 942
rect 1111 946 1115 947
rect 1111 941 1115 942
rect 1151 946 1155 947
rect 1151 941 1155 942
rect 1223 946 1227 947
rect 1223 941 1227 942
rect 1271 946 1275 947
rect 1271 941 1275 942
rect 1335 946 1339 947
rect 1335 941 1339 942
rect 1391 946 1395 947
rect 1391 941 1395 942
rect 1455 946 1459 947
rect 1455 941 1459 942
rect 1511 946 1515 947
rect 1511 941 1515 942
rect 1631 946 1635 947
rect 1631 941 1635 942
rect 1831 946 1835 947
rect 1831 941 1835 942
rect 1871 946 1875 947
rect 1871 941 1875 942
rect 1895 946 1899 947
rect 1895 941 1899 942
rect 1983 946 1987 947
rect 1983 941 1987 942
rect 2023 946 2027 947
rect 2023 941 2027 942
rect 2111 946 2115 947
rect 2111 941 2115 942
rect 2119 946 2123 947
rect 2119 941 2123 942
rect 2223 946 2227 947
rect 2223 941 2227 942
rect 2263 946 2267 947
rect 2263 941 2267 942
rect 2343 946 2347 947
rect 2343 941 2347 942
rect 2423 946 2427 947
rect 2423 941 2427 942
rect 2463 946 2467 947
rect 2463 941 2467 942
rect 2583 946 2587 947
rect 2583 941 2587 942
rect 2591 946 2595 947
rect 2591 941 2595 942
rect 2719 946 2723 947
rect 2719 941 2723 942
rect 2735 946 2739 947
rect 2735 941 2739 942
rect 2847 946 2851 947
rect 2847 941 2851 942
rect 2879 946 2883 947
rect 2879 941 2883 942
rect 2975 946 2979 947
rect 2975 941 2979 942
rect 3015 946 3019 947
rect 3015 941 3019 942
rect 3103 946 3107 947
rect 3103 941 3107 942
rect 3143 946 3147 947
rect 3143 941 3147 942
rect 3239 946 3243 947
rect 3239 941 3243 942
rect 3271 946 3275 947
rect 3271 941 3275 942
rect 3383 946 3387 947
rect 3383 941 3387 942
rect 3399 946 3403 947
rect 3399 941 3403 942
rect 3503 946 3507 947
rect 3503 941 3507 942
rect 3591 946 3595 947
rect 3591 941 3595 942
rect 112 922 114 941
rect 136 925 138 941
rect 216 925 218 941
rect 336 925 338 941
rect 464 925 466 941
rect 600 925 602 941
rect 736 925 738 941
rect 864 925 866 941
rect 992 925 994 941
rect 1112 925 1114 941
rect 1224 925 1226 941
rect 1336 925 1338 941
rect 1456 925 1458 941
rect 134 924 140 925
rect 110 921 116 922
rect 110 917 111 921
rect 115 917 116 921
rect 134 920 135 924
rect 139 920 140 924
rect 134 919 140 920
rect 214 924 220 925
rect 214 920 215 924
rect 219 920 220 924
rect 214 919 220 920
rect 334 924 340 925
rect 334 920 335 924
rect 339 920 340 924
rect 334 919 340 920
rect 462 924 468 925
rect 462 920 463 924
rect 467 920 468 924
rect 462 919 468 920
rect 598 924 604 925
rect 598 920 599 924
rect 603 920 604 924
rect 598 919 604 920
rect 734 924 740 925
rect 734 920 735 924
rect 739 920 740 924
rect 734 919 740 920
rect 862 924 868 925
rect 862 920 863 924
rect 867 920 868 924
rect 862 919 868 920
rect 990 924 996 925
rect 990 920 991 924
rect 995 920 996 924
rect 990 919 996 920
rect 1110 924 1116 925
rect 1110 920 1111 924
rect 1115 920 1116 924
rect 1110 919 1116 920
rect 1222 924 1228 925
rect 1222 920 1223 924
rect 1227 920 1228 924
rect 1222 919 1228 920
rect 1334 924 1340 925
rect 1334 920 1335 924
rect 1339 920 1340 924
rect 1334 919 1340 920
rect 1454 924 1460 925
rect 1454 920 1455 924
rect 1459 920 1460 924
rect 1832 922 1834 941
rect 1872 922 1874 941
rect 1896 925 1898 941
rect 1984 925 1986 941
rect 2112 925 2114 941
rect 2264 925 2266 941
rect 2424 925 2426 941
rect 2584 925 2586 941
rect 2736 925 2738 941
rect 2880 925 2882 941
rect 3016 925 3018 941
rect 3144 925 3146 941
rect 3272 925 3274 941
rect 3400 925 3402 941
rect 3504 925 3506 941
rect 1894 924 1900 925
rect 1454 919 1460 920
rect 1830 921 1836 922
rect 110 916 116 917
rect 1830 917 1831 921
rect 1835 917 1836 921
rect 1830 916 1836 917
rect 1870 921 1876 922
rect 1870 917 1871 921
rect 1875 917 1876 921
rect 1894 920 1895 924
rect 1899 920 1900 924
rect 1894 919 1900 920
rect 1982 924 1988 925
rect 1982 920 1983 924
rect 1987 920 1988 924
rect 1982 919 1988 920
rect 2110 924 2116 925
rect 2110 920 2111 924
rect 2115 920 2116 924
rect 2110 919 2116 920
rect 2262 924 2268 925
rect 2262 920 2263 924
rect 2267 920 2268 924
rect 2262 919 2268 920
rect 2422 924 2428 925
rect 2422 920 2423 924
rect 2427 920 2428 924
rect 2422 919 2428 920
rect 2582 924 2588 925
rect 2582 920 2583 924
rect 2587 920 2588 924
rect 2582 919 2588 920
rect 2734 924 2740 925
rect 2734 920 2735 924
rect 2739 920 2740 924
rect 2734 919 2740 920
rect 2878 924 2884 925
rect 2878 920 2879 924
rect 2883 920 2884 924
rect 2878 919 2884 920
rect 3014 924 3020 925
rect 3014 920 3015 924
rect 3019 920 3020 924
rect 3014 919 3020 920
rect 3142 924 3148 925
rect 3142 920 3143 924
rect 3147 920 3148 924
rect 3142 919 3148 920
rect 3270 924 3276 925
rect 3270 920 3271 924
rect 3275 920 3276 924
rect 3270 919 3276 920
rect 3398 924 3404 925
rect 3398 920 3399 924
rect 3403 920 3404 924
rect 3398 919 3404 920
rect 3502 924 3508 925
rect 3502 920 3503 924
rect 3507 920 3508 924
rect 3592 922 3594 941
rect 3502 919 3508 920
rect 3590 921 3596 922
rect 1870 916 1876 917
rect 3590 917 3591 921
rect 3595 917 3596 921
rect 3590 916 3596 917
rect 110 904 116 905
rect 110 900 111 904
rect 115 900 116 904
rect 110 899 116 900
rect 1830 904 1836 905
rect 1830 900 1831 904
rect 1835 900 1836 904
rect 1830 899 1836 900
rect 1870 904 1876 905
rect 1870 900 1871 904
rect 1875 900 1876 904
rect 1870 899 1876 900
rect 3590 904 3596 905
rect 3590 900 3591 904
rect 3595 900 3596 904
rect 3590 899 3596 900
rect 112 859 114 899
rect 142 886 148 887
rect 142 882 143 886
rect 147 882 148 886
rect 142 881 148 882
rect 222 886 228 887
rect 222 882 223 886
rect 227 882 228 886
rect 222 881 228 882
rect 342 886 348 887
rect 342 882 343 886
rect 347 882 348 886
rect 342 881 348 882
rect 470 886 476 887
rect 470 882 471 886
rect 475 882 476 886
rect 470 881 476 882
rect 606 886 612 887
rect 606 882 607 886
rect 611 882 612 886
rect 606 881 612 882
rect 742 886 748 887
rect 742 882 743 886
rect 747 882 748 886
rect 742 881 748 882
rect 870 886 876 887
rect 870 882 871 886
rect 875 882 876 886
rect 870 881 876 882
rect 998 886 1004 887
rect 998 882 999 886
rect 1003 882 1004 886
rect 998 881 1004 882
rect 1118 886 1124 887
rect 1118 882 1119 886
rect 1123 882 1124 886
rect 1118 881 1124 882
rect 1230 886 1236 887
rect 1230 882 1231 886
rect 1235 882 1236 886
rect 1230 881 1236 882
rect 1342 886 1348 887
rect 1342 882 1343 886
rect 1347 882 1348 886
rect 1342 881 1348 882
rect 1462 886 1468 887
rect 1462 882 1463 886
rect 1467 882 1468 886
rect 1462 881 1468 882
rect 144 859 146 881
rect 224 859 226 881
rect 344 859 346 881
rect 472 859 474 881
rect 608 859 610 881
rect 744 859 746 881
rect 872 859 874 881
rect 1000 859 1002 881
rect 1120 859 1122 881
rect 1232 859 1234 881
rect 1344 859 1346 881
rect 1464 859 1466 881
rect 1832 859 1834 899
rect 1872 863 1874 899
rect 1902 886 1908 887
rect 1902 882 1903 886
rect 1907 882 1908 886
rect 1902 881 1908 882
rect 1990 886 1996 887
rect 1990 882 1991 886
rect 1995 882 1996 886
rect 1990 881 1996 882
rect 2118 886 2124 887
rect 2118 882 2119 886
rect 2123 882 2124 886
rect 2118 881 2124 882
rect 2270 886 2276 887
rect 2270 882 2271 886
rect 2275 882 2276 886
rect 2270 881 2276 882
rect 2430 886 2436 887
rect 2430 882 2431 886
rect 2435 882 2436 886
rect 2430 881 2436 882
rect 2590 886 2596 887
rect 2590 882 2591 886
rect 2595 882 2596 886
rect 2590 881 2596 882
rect 2742 886 2748 887
rect 2742 882 2743 886
rect 2747 882 2748 886
rect 2742 881 2748 882
rect 2886 886 2892 887
rect 2886 882 2887 886
rect 2891 882 2892 886
rect 2886 881 2892 882
rect 3022 886 3028 887
rect 3022 882 3023 886
rect 3027 882 3028 886
rect 3022 881 3028 882
rect 3150 886 3156 887
rect 3150 882 3151 886
rect 3155 882 3156 886
rect 3150 881 3156 882
rect 3278 886 3284 887
rect 3278 882 3279 886
rect 3283 882 3284 886
rect 3278 881 3284 882
rect 3406 886 3412 887
rect 3406 882 3407 886
rect 3411 882 3412 886
rect 3406 881 3412 882
rect 3510 886 3516 887
rect 3510 882 3511 886
rect 3515 882 3516 886
rect 3510 881 3516 882
rect 1904 863 1906 881
rect 1992 863 1994 881
rect 2120 863 2122 881
rect 2272 863 2274 881
rect 2432 863 2434 881
rect 2592 863 2594 881
rect 2744 863 2746 881
rect 2888 863 2890 881
rect 3024 863 3026 881
rect 3152 863 3154 881
rect 3280 863 3282 881
rect 3408 863 3410 881
rect 3512 863 3514 881
rect 3592 863 3594 899
rect 1871 862 1875 863
rect 111 858 115 859
rect 111 853 115 854
rect 143 858 147 859
rect 143 853 147 854
rect 223 858 227 859
rect 223 853 227 854
rect 303 858 307 859
rect 303 853 307 854
rect 343 858 347 859
rect 343 853 347 854
rect 391 858 395 859
rect 391 853 395 854
rect 471 858 475 859
rect 471 853 475 854
rect 495 858 499 859
rect 495 853 499 854
rect 599 858 603 859
rect 599 853 603 854
rect 607 858 611 859
rect 607 853 611 854
rect 711 858 715 859
rect 711 853 715 854
rect 743 858 747 859
rect 743 853 747 854
rect 839 858 843 859
rect 839 853 843 854
rect 871 858 875 859
rect 871 853 875 854
rect 991 858 995 859
rect 991 853 995 854
rect 999 858 1003 859
rect 999 853 1003 854
rect 1119 858 1123 859
rect 1119 853 1123 854
rect 1167 858 1171 859
rect 1167 853 1171 854
rect 1231 858 1235 859
rect 1231 853 1235 854
rect 1343 858 1347 859
rect 1343 853 1347 854
rect 1359 858 1363 859
rect 1359 853 1363 854
rect 1463 858 1467 859
rect 1463 853 1467 854
rect 1567 858 1571 859
rect 1567 853 1571 854
rect 1751 858 1755 859
rect 1751 853 1755 854
rect 1831 858 1835 859
rect 1871 857 1875 858
rect 1903 862 1907 863
rect 1903 857 1907 858
rect 1991 862 1995 863
rect 1991 857 1995 858
rect 2039 862 2043 863
rect 2039 857 2043 858
rect 2119 862 2123 863
rect 2119 857 2123 858
rect 2215 862 2219 863
rect 2215 857 2219 858
rect 2271 862 2275 863
rect 2271 857 2275 858
rect 2391 862 2395 863
rect 2391 857 2395 858
rect 2431 862 2435 863
rect 2431 857 2435 858
rect 2567 862 2571 863
rect 2567 857 2571 858
rect 2591 862 2595 863
rect 2591 857 2595 858
rect 2735 862 2739 863
rect 2735 857 2739 858
rect 2743 862 2747 863
rect 2743 857 2747 858
rect 2887 862 2891 863
rect 2887 857 2891 858
rect 3023 862 3027 863
rect 3023 857 3027 858
rect 3031 862 3035 863
rect 3031 857 3035 858
rect 3151 862 3155 863
rect 3151 857 3155 858
rect 3159 862 3163 863
rect 3159 857 3163 858
rect 3279 862 3283 863
rect 3279 857 3283 858
rect 3287 862 3291 863
rect 3287 857 3291 858
rect 3407 862 3411 863
rect 3407 857 3411 858
rect 3511 862 3515 863
rect 3511 857 3515 858
rect 3591 862 3595 863
rect 3591 857 3595 858
rect 1831 853 1835 854
rect 112 825 114 853
rect 144 843 146 853
rect 224 843 226 853
rect 304 843 306 853
rect 392 843 394 853
rect 496 843 498 853
rect 600 843 602 853
rect 712 843 714 853
rect 840 843 842 853
rect 992 843 994 853
rect 1168 843 1170 853
rect 1360 843 1362 853
rect 1568 843 1570 853
rect 1752 843 1754 853
rect 142 842 148 843
rect 142 838 143 842
rect 147 838 148 842
rect 142 837 148 838
rect 222 842 228 843
rect 222 838 223 842
rect 227 838 228 842
rect 222 837 228 838
rect 302 842 308 843
rect 302 838 303 842
rect 307 838 308 842
rect 302 837 308 838
rect 390 842 396 843
rect 390 838 391 842
rect 395 838 396 842
rect 390 837 396 838
rect 494 842 500 843
rect 494 838 495 842
rect 499 838 500 842
rect 494 837 500 838
rect 598 842 604 843
rect 598 838 599 842
rect 603 838 604 842
rect 598 837 604 838
rect 710 842 716 843
rect 710 838 711 842
rect 715 838 716 842
rect 710 837 716 838
rect 838 842 844 843
rect 838 838 839 842
rect 843 838 844 842
rect 838 837 844 838
rect 990 842 996 843
rect 990 838 991 842
rect 995 838 996 842
rect 990 837 996 838
rect 1166 842 1172 843
rect 1166 838 1167 842
rect 1171 838 1172 842
rect 1166 837 1172 838
rect 1358 842 1364 843
rect 1358 838 1359 842
rect 1363 838 1364 842
rect 1358 837 1364 838
rect 1566 842 1572 843
rect 1566 838 1567 842
rect 1571 838 1572 842
rect 1566 837 1572 838
rect 1750 842 1756 843
rect 1750 838 1751 842
rect 1755 838 1756 842
rect 1750 837 1756 838
rect 1832 825 1834 853
rect 1872 829 1874 857
rect 1904 847 1906 857
rect 2040 847 2042 857
rect 2216 847 2218 857
rect 2392 847 2394 857
rect 2568 847 2570 857
rect 2736 847 2738 857
rect 2888 847 2890 857
rect 3032 847 3034 857
rect 3160 847 3162 857
rect 3288 847 3290 857
rect 3408 847 3410 857
rect 3512 847 3514 857
rect 1902 846 1908 847
rect 1902 842 1903 846
rect 1907 842 1908 846
rect 1902 841 1908 842
rect 2038 846 2044 847
rect 2038 842 2039 846
rect 2043 842 2044 846
rect 2038 841 2044 842
rect 2214 846 2220 847
rect 2214 842 2215 846
rect 2219 842 2220 846
rect 2214 841 2220 842
rect 2390 846 2396 847
rect 2390 842 2391 846
rect 2395 842 2396 846
rect 2390 841 2396 842
rect 2566 846 2572 847
rect 2566 842 2567 846
rect 2571 842 2572 846
rect 2566 841 2572 842
rect 2734 846 2740 847
rect 2734 842 2735 846
rect 2739 842 2740 846
rect 2734 841 2740 842
rect 2886 846 2892 847
rect 2886 842 2887 846
rect 2891 842 2892 846
rect 2886 841 2892 842
rect 3030 846 3036 847
rect 3030 842 3031 846
rect 3035 842 3036 846
rect 3030 841 3036 842
rect 3158 846 3164 847
rect 3158 842 3159 846
rect 3163 842 3164 846
rect 3158 841 3164 842
rect 3286 846 3292 847
rect 3286 842 3287 846
rect 3291 842 3292 846
rect 3286 841 3292 842
rect 3406 846 3412 847
rect 3406 842 3407 846
rect 3411 842 3412 846
rect 3406 841 3412 842
rect 3510 846 3516 847
rect 3510 842 3511 846
rect 3515 842 3516 846
rect 3510 841 3516 842
rect 3592 829 3594 857
rect 1870 828 1876 829
rect 110 824 116 825
rect 110 820 111 824
rect 115 820 116 824
rect 110 819 116 820
rect 1830 824 1836 825
rect 1830 820 1831 824
rect 1835 820 1836 824
rect 1870 824 1871 828
rect 1875 824 1876 828
rect 1870 823 1876 824
rect 3590 828 3596 829
rect 3590 824 3591 828
rect 3595 824 3596 828
rect 3590 823 3596 824
rect 1830 819 1836 820
rect 1870 811 1876 812
rect 110 807 116 808
rect 110 803 111 807
rect 115 803 116 807
rect 1830 807 1836 808
rect 110 802 116 803
rect 134 804 140 805
rect 112 779 114 802
rect 134 800 135 804
rect 139 800 140 804
rect 134 799 140 800
rect 214 804 220 805
rect 214 800 215 804
rect 219 800 220 804
rect 214 799 220 800
rect 294 804 300 805
rect 294 800 295 804
rect 299 800 300 804
rect 294 799 300 800
rect 382 804 388 805
rect 382 800 383 804
rect 387 800 388 804
rect 382 799 388 800
rect 486 804 492 805
rect 486 800 487 804
rect 491 800 492 804
rect 486 799 492 800
rect 590 804 596 805
rect 590 800 591 804
rect 595 800 596 804
rect 590 799 596 800
rect 702 804 708 805
rect 702 800 703 804
rect 707 800 708 804
rect 702 799 708 800
rect 830 804 836 805
rect 830 800 831 804
rect 835 800 836 804
rect 830 799 836 800
rect 982 804 988 805
rect 982 800 983 804
rect 987 800 988 804
rect 982 799 988 800
rect 1158 804 1164 805
rect 1158 800 1159 804
rect 1163 800 1164 804
rect 1158 799 1164 800
rect 1350 804 1356 805
rect 1350 800 1351 804
rect 1355 800 1356 804
rect 1350 799 1356 800
rect 1558 804 1564 805
rect 1558 800 1559 804
rect 1563 800 1564 804
rect 1558 799 1564 800
rect 1742 804 1748 805
rect 1742 800 1743 804
rect 1747 800 1748 804
rect 1830 803 1831 807
rect 1835 803 1836 807
rect 1870 807 1871 811
rect 1875 807 1876 811
rect 3590 811 3596 812
rect 1870 806 1876 807
rect 1894 808 1900 809
rect 1830 802 1836 803
rect 1742 799 1748 800
rect 136 779 138 799
rect 216 779 218 799
rect 296 779 298 799
rect 384 779 386 799
rect 488 779 490 799
rect 592 779 594 799
rect 704 779 706 799
rect 832 779 834 799
rect 984 779 986 799
rect 1160 779 1162 799
rect 1352 779 1354 799
rect 1560 779 1562 799
rect 1744 779 1746 799
rect 1832 779 1834 802
rect 111 778 115 779
rect 111 773 115 774
rect 135 778 139 779
rect 135 773 139 774
rect 199 778 203 779
rect 199 773 203 774
rect 215 778 219 779
rect 215 773 219 774
rect 287 778 291 779
rect 287 773 291 774
rect 295 778 299 779
rect 295 773 299 774
rect 383 778 387 779
rect 383 773 387 774
rect 391 778 395 779
rect 391 773 395 774
rect 487 778 491 779
rect 487 773 491 774
rect 503 778 507 779
rect 503 773 507 774
rect 591 778 595 779
rect 591 773 595 774
rect 615 778 619 779
rect 615 773 619 774
rect 703 778 707 779
rect 703 773 707 774
rect 735 778 739 779
rect 735 773 739 774
rect 831 778 835 779
rect 831 773 835 774
rect 855 778 859 779
rect 855 773 859 774
rect 983 778 987 779
rect 983 773 987 774
rect 1111 778 1115 779
rect 1111 773 1115 774
rect 1159 778 1163 779
rect 1159 773 1163 774
rect 1239 778 1243 779
rect 1239 773 1243 774
rect 1351 778 1355 779
rect 1351 773 1355 774
rect 1367 778 1371 779
rect 1367 773 1371 774
rect 1495 778 1499 779
rect 1495 773 1499 774
rect 1559 778 1563 779
rect 1559 773 1563 774
rect 1631 778 1635 779
rect 1631 773 1635 774
rect 1743 778 1747 779
rect 1743 773 1747 774
rect 1831 778 1835 779
rect 1831 773 1835 774
rect 112 754 114 773
rect 200 757 202 773
rect 288 757 290 773
rect 392 757 394 773
rect 504 757 506 773
rect 616 757 618 773
rect 736 757 738 773
rect 856 757 858 773
rect 984 757 986 773
rect 1112 757 1114 773
rect 1240 757 1242 773
rect 1368 757 1370 773
rect 1496 757 1498 773
rect 1632 757 1634 773
rect 1744 757 1746 773
rect 198 756 204 757
rect 110 753 116 754
rect 110 749 111 753
rect 115 749 116 753
rect 198 752 199 756
rect 203 752 204 756
rect 198 751 204 752
rect 286 756 292 757
rect 286 752 287 756
rect 291 752 292 756
rect 286 751 292 752
rect 390 756 396 757
rect 390 752 391 756
rect 395 752 396 756
rect 390 751 396 752
rect 502 756 508 757
rect 502 752 503 756
rect 507 752 508 756
rect 502 751 508 752
rect 614 756 620 757
rect 614 752 615 756
rect 619 752 620 756
rect 614 751 620 752
rect 734 756 740 757
rect 734 752 735 756
rect 739 752 740 756
rect 734 751 740 752
rect 854 756 860 757
rect 854 752 855 756
rect 859 752 860 756
rect 854 751 860 752
rect 982 756 988 757
rect 982 752 983 756
rect 987 752 988 756
rect 982 751 988 752
rect 1110 756 1116 757
rect 1110 752 1111 756
rect 1115 752 1116 756
rect 1110 751 1116 752
rect 1238 756 1244 757
rect 1238 752 1239 756
rect 1243 752 1244 756
rect 1238 751 1244 752
rect 1366 756 1372 757
rect 1366 752 1367 756
rect 1371 752 1372 756
rect 1366 751 1372 752
rect 1494 756 1500 757
rect 1494 752 1495 756
rect 1499 752 1500 756
rect 1494 751 1500 752
rect 1630 756 1636 757
rect 1630 752 1631 756
rect 1635 752 1636 756
rect 1630 751 1636 752
rect 1742 756 1748 757
rect 1742 752 1743 756
rect 1747 752 1748 756
rect 1832 754 1834 773
rect 1872 771 1874 806
rect 1894 804 1895 808
rect 1899 804 1900 808
rect 1894 803 1900 804
rect 2030 808 2036 809
rect 2030 804 2031 808
rect 2035 804 2036 808
rect 2030 803 2036 804
rect 2206 808 2212 809
rect 2206 804 2207 808
rect 2211 804 2212 808
rect 2206 803 2212 804
rect 2382 808 2388 809
rect 2382 804 2383 808
rect 2387 804 2388 808
rect 2382 803 2388 804
rect 2558 808 2564 809
rect 2558 804 2559 808
rect 2563 804 2564 808
rect 2558 803 2564 804
rect 2726 808 2732 809
rect 2726 804 2727 808
rect 2731 804 2732 808
rect 2726 803 2732 804
rect 2878 808 2884 809
rect 2878 804 2879 808
rect 2883 804 2884 808
rect 2878 803 2884 804
rect 3022 808 3028 809
rect 3022 804 3023 808
rect 3027 804 3028 808
rect 3022 803 3028 804
rect 3150 808 3156 809
rect 3150 804 3151 808
rect 3155 804 3156 808
rect 3150 803 3156 804
rect 3278 808 3284 809
rect 3278 804 3279 808
rect 3283 804 3284 808
rect 3278 803 3284 804
rect 3398 808 3404 809
rect 3398 804 3399 808
rect 3403 804 3404 808
rect 3398 803 3404 804
rect 3502 808 3508 809
rect 3502 804 3503 808
rect 3507 804 3508 808
rect 3590 807 3591 811
rect 3595 807 3596 811
rect 3590 806 3596 807
rect 3502 803 3508 804
rect 1896 771 1898 803
rect 2032 771 2034 803
rect 2208 771 2210 803
rect 2384 771 2386 803
rect 2560 771 2562 803
rect 2728 771 2730 803
rect 2880 771 2882 803
rect 3024 771 3026 803
rect 3152 771 3154 803
rect 3280 771 3282 803
rect 3400 771 3402 803
rect 3504 771 3506 803
rect 3592 771 3594 806
rect 1871 770 1875 771
rect 1871 765 1875 766
rect 1895 770 1899 771
rect 1895 765 1899 766
rect 2023 770 2027 771
rect 2023 765 2027 766
rect 2031 770 2035 771
rect 2031 765 2035 766
rect 2191 770 2195 771
rect 2191 765 2195 766
rect 2207 770 2211 771
rect 2207 765 2211 766
rect 2359 770 2363 771
rect 2359 765 2363 766
rect 2383 770 2387 771
rect 2383 765 2387 766
rect 2519 770 2523 771
rect 2519 765 2523 766
rect 2559 770 2563 771
rect 2559 765 2563 766
rect 2679 770 2683 771
rect 2679 765 2683 766
rect 2727 770 2731 771
rect 2727 765 2731 766
rect 2831 770 2835 771
rect 2831 765 2835 766
rect 2879 770 2883 771
rect 2879 765 2883 766
rect 2975 770 2979 771
rect 2975 765 2979 766
rect 3023 770 3027 771
rect 3023 765 3027 766
rect 3111 770 3115 771
rect 3111 765 3115 766
rect 3151 770 3155 771
rect 3151 765 3155 766
rect 3247 770 3251 771
rect 3247 765 3251 766
rect 3279 770 3283 771
rect 3279 765 3283 766
rect 3383 770 3387 771
rect 3383 765 3387 766
rect 3399 770 3403 771
rect 3399 765 3403 766
rect 3503 770 3507 771
rect 3503 765 3507 766
rect 3591 770 3595 771
rect 3591 765 3595 766
rect 1742 751 1748 752
rect 1830 753 1836 754
rect 110 748 116 749
rect 1830 749 1831 753
rect 1835 749 1836 753
rect 1830 748 1836 749
rect 1872 746 1874 765
rect 2024 749 2026 765
rect 2192 749 2194 765
rect 2360 749 2362 765
rect 2520 749 2522 765
rect 2680 749 2682 765
rect 2832 749 2834 765
rect 2976 749 2978 765
rect 3112 749 3114 765
rect 3248 749 3250 765
rect 3384 749 3386 765
rect 3504 749 3506 765
rect 2022 748 2028 749
rect 1870 745 1876 746
rect 1870 741 1871 745
rect 1875 741 1876 745
rect 2022 744 2023 748
rect 2027 744 2028 748
rect 2022 743 2028 744
rect 2190 748 2196 749
rect 2190 744 2191 748
rect 2195 744 2196 748
rect 2190 743 2196 744
rect 2358 748 2364 749
rect 2358 744 2359 748
rect 2363 744 2364 748
rect 2358 743 2364 744
rect 2518 748 2524 749
rect 2518 744 2519 748
rect 2523 744 2524 748
rect 2518 743 2524 744
rect 2678 748 2684 749
rect 2678 744 2679 748
rect 2683 744 2684 748
rect 2678 743 2684 744
rect 2830 748 2836 749
rect 2830 744 2831 748
rect 2835 744 2836 748
rect 2830 743 2836 744
rect 2974 748 2980 749
rect 2974 744 2975 748
rect 2979 744 2980 748
rect 2974 743 2980 744
rect 3110 748 3116 749
rect 3110 744 3111 748
rect 3115 744 3116 748
rect 3110 743 3116 744
rect 3246 748 3252 749
rect 3246 744 3247 748
rect 3251 744 3252 748
rect 3246 743 3252 744
rect 3382 748 3388 749
rect 3382 744 3383 748
rect 3387 744 3388 748
rect 3382 743 3388 744
rect 3502 748 3508 749
rect 3502 744 3503 748
rect 3507 744 3508 748
rect 3592 746 3594 765
rect 3502 743 3508 744
rect 3590 745 3596 746
rect 1870 740 1876 741
rect 3590 741 3591 745
rect 3595 741 3596 745
rect 3590 740 3596 741
rect 110 736 116 737
rect 110 732 111 736
rect 115 732 116 736
rect 110 731 116 732
rect 1830 736 1836 737
rect 1830 732 1831 736
rect 1835 732 1836 736
rect 1830 731 1836 732
rect 112 687 114 731
rect 206 718 212 719
rect 206 714 207 718
rect 211 714 212 718
rect 206 713 212 714
rect 294 718 300 719
rect 294 714 295 718
rect 299 714 300 718
rect 294 713 300 714
rect 398 718 404 719
rect 398 714 399 718
rect 403 714 404 718
rect 398 713 404 714
rect 510 718 516 719
rect 510 714 511 718
rect 515 714 516 718
rect 510 713 516 714
rect 622 718 628 719
rect 622 714 623 718
rect 627 714 628 718
rect 622 713 628 714
rect 742 718 748 719
rect 742 714 743 718
rect 747 714 748 718
rect 742 713 748 714
rect 862 718 868 719
rect 862 714 863 718
rect 867 714 868 718
rect 862 713 868 714
rect 990 718 996 719
rect 990 714 991 718
rect 995 714 996 718
rect 990 713 996 714
rect 1118 718 1124 719
rect 1118 714 1119 718
rect 1123 714 1124 718
rect 1118 713 1124 714
rect 1246 718 1252 719
rect 1246 714 1247 718
rect 1251 714 1252 718
rect 1246 713 1252 714
rect 1374 718 1380 719
rect 1374 714 1375 718
rect 1379 714 1380 718
rect 1374 713 1380 714
rect 1502 718 1508 719
rect 1502 714 1503 718
rect 1507 714 1508 718
rect 1502 713 1508 714
rect 1638 718 1644 719
rect 1638 714 1639 718
rect 1643 714 1644 718
rect 1638 713 1644 714
rect 1750 718 1756 719
rect 1750 714 1751 718
rect 1755 714 1756 718
rect 1750 713 1756 714
rect 208 687 210 713
rect 296 687 298 713
rect 400 687 402 713
rect 512 687 514 713
rect 624 687 626 713
rect 744 687 746 713
rect 864 687 866 713
rect 992 687 994 713
rect 1120 687 1122 713
rect 1248 687 1250 713
rect 1376 687 1378 713
rect 1504 687 1506 713
rect 1640 687 1642 713
rect 1752 687 1754 713
rect 1832 687 1834 731
rect 1870 728 1876 729
rect 1870 724 1871 728
rect 1875 724 1876 728
rect 1870 723 1876 724
rect 3590 728 3596 729
rect 3590 724 3591 728
rect 3595 724 3596 728
rect 3590 723 3596 724
rect 1872 691 1874 723
rect 2030 710 2036 711
rect 2030 706 2031 710
rect 2035 706 2036 710
rect 2030 705 2036 706
rect 2198 710 2204 711
rect 2198 706 2199 710
rect 2203 706 2204 710
rect 2198 705 2204 706
rect 2366 710 2372 711
rect 2366 706 2367 710
rect 2371 706 2372 710
rect 2366 705 2372 706
rect 2526 710 2532 711
rect 2526 706 2527 710
rect 2531 706 2532 710
rect 2526 705 2532 706
rect 2686 710 2692 711
rect 2686 706 2687 710
rect 2691 706 2692 710
rect 2686 705 2692 706
rect 2838 710 2844 711
rect 2838 706 2839 710
rect 2843 706 2844 710
rect 2838 705 2844 706
rect 2982 710 2988 711
rect 2982 706 2983 710
rect 2987 706 2988 710
rect 2982 705 2988 706
rect 3118 710 3124 711
rect 3118 706 3119 710
rect 3123 706 3124 710
rect 3118 705 3124 706
rect 3254 710 3260 711
rect 3254 706 3255 710
rect 3259 706 3260 710
rect 3254 705 3260 706
rect 3390 710 3396 711
rect 3390 706 3391 710
rect 3395 706 3396 710
rect 3390 705 3396 706
rect 3510 710 3516 711
rect 3510 706 3511 710
rect 3515 706 3516 710
rect 3510 705 3516 706
rect 2032 691 2034 705
rect 2200 691 2202 705
rect 2368 691 2370 705
rect 2528 691 2530 705
rect 2688 691 2690 705
rect 2840 691 2842 705
rect 2984 691 2986 705
rect 3120 691 3122 705
rect 3256 691 3258 705
rect 3392 691 3394 705
rect 3512 691 3514 705
rect 3592 691 3594 723
rect 1871 690 1875 691
rect 111 686 115 687
rect 111 681 115 682
rect 207 686 211 687
rect 207 681 211 682
rect 295 686 299 687
rect 295 681 299 682
rect 383 686 387 687
rect 383 681 387 682
rect 399 686 403 687
rect 399 681 403 682
rect 479 686 483 687
rect 479 681 483 682
rect 511 686 515 687
rect 511 681 515 682
rect 591 686 595 687
rect 591 681 595 682
rect 623 686 627 687
rect 623 681 627 682
rect 719 686 723 687
rect 719 681 723 682
rect 743 686 747 687
rect 743 681 747 682
rect 855 686 859 687
rect 855 681 859 682
rect 863 686 867 687
rect 863 681 867 682
rect 991 686 995 687
rect 991 681 995 682
rect 1119 686 1123 687
rect 1119 681 1123 682
rect 1127 686 1131 687
rect 1127 681 1131 682
rect 1247 686 1251 687
rect 1247 681 1251 682
rect 1255 686 1259 687
rect 1255 681 1259 682
rect 1375 686 1379 687
rect 1375 681 1379 682
rect 1383 686 1387 687
rect 1383 681 1387 682
rect 1503 686 1507 687
rect 1503 681 1507 682
rect 1631 686 1635 687
rect 1631 681 1635 682
rect 1639 686 1643 687
rect 1639 681 1643 682
rect 1751 686 1755 687
rect 1751 681 1755 682
rect 1831 686 1835 687
rect 1871 685 1875 686
rect 2031 690 2035 691
rect 2031 685 2035 686
rect 2095 690 2099 691
rect 2095 685 2099 686
rect 2175 690 2179 691
rect 2175 685 2179 686
rect 2199 690 2203 691
rect 2199 685 2203 686
rect 2263 690 2267 691
rect 2263 685 2267 686
rect 2359 690 2363 691
rect 2359 685 2363 686
rect 2367 690 2371 691
rect 2367 685 2371 686
rect 2463 690 2467 691
rect 2463 685 2467 686
rect 2527 690 2531 691
rect 2527 685 2531 686
rect 2567 690 2571 691
rect 2567 685 2571 686
rect 2679 690 2683 691
rect 2679 685 2683 686
rect 2687 690 2691 691
rect 2687 685 2691 686
rect 2799 690 2803 691
rect 2799 685 2803 686
rect 2839 690 2843 691
rect 2839 685 2843 686
rect 2927 690 2931 691
rect 2927 685 2931 686
rect 2983 690 2987 691
rect 2983 685 2987 686
rect 3071 690 3075 691
rect 3071 685 3075 686
rect 3119 690 3123 691
rect 3119 685 3123 686
rect 3223 690 3227 691
rect 3223 685 3227 686
rect 3255 690 3259 691
rect 3255 685 3259 686
rect 3375 690 3379 691
rect 3375 685 3379 686
rect 3391 690 3395 691
rect 3391 685 3395 686
rect 3511 690 3515 691
rect 3511 685 3515 686
rect 3591 690 3595 691
rect 3591 685 3595 686
rect 1831 681 1835 682
rect 112 653 114 681
rect 384 671 386 681
rect 480 671 482 681
rect 592 671 594 681
rect 720 671 722 681
rect 856 671 858 681
rect 992 671 994 681
rect 1128 671 1130 681
rect 1256 671 1258 681
rect 1384 671 1386 681
rect 1504 671 1506 681
rect 1632 671 1634 681
rect 1752 671 1754 681
rect 382 670 388 671
rect 382 666 383 670
rect 387 666 388 670
rect 382 665 388 666
rect 478 670 484 671
rect 478 666 479 670
rect 483 666 484 670
rect 478 665 484 666
rect 590 670 596 671
rect 590 666 591 670
rect 595 666 596 670
rect 590 665 596 666
rect 718 670 724 671
rect 718 666 719 670
rect 723 666 724 670
rect 718 665 724 666
rect 854 670 860 671
rect 854 666 855 670
rect 859 666 860 670
rect 854 665 860 666
rect 990 670 996 671
rect 990 666 991 670
rect 995 666 996 670
rect 990 665 996 666
rect 1126 670 1132 671
rect 1126 666 1127 670
rect 1131 666 1132 670
rect 1126 665 1132 666
rect 1254 670 1260 671
rect 1254 666 1255 670
rect 1259 666 1260 670
rect 1254 665 1260 666
rect 1382 670 1388 671
rect 1382 666 1383 670
rect 1387 666 1388 670
rect 1382 665 1388 666
rect 1502 670 1508 671
rect 1502 666 1503 670
rect 1507 666 1508 670
rect 1502 665 1508 666
rect 1630 670 1636 671
rect 1630 666 1631 670
rect 1635 666 1636 670
rect 1630 665 1636 666
rect 1750 670 1756 671
rect 1750 666 1751 670
rect 1755 666 1756 670
rect 1750 665 1756 666
rect 1832 653 1834 681
rect 1872 657 1874 685
rect 2096 675 2098 685
rect 2176 675 2178 685
rect 2264 675 2266 685
rect 2360 675 2362 685
rect 2464 675 2466 685
rect 2568 675 2570 685
rect 2680 675 2682 685
rect 2800 675 2802 685
rect 2928 675 2930 685
rect 3072 675 3074 685
rect 3224 675 3226 685
rect 3376 675 3378 685
rect 3512 675 3514 685
rect 2094 674 2100 675
rect 2094 670 2095 674
rect 2099 670 2100 674
rect 2094 669 2100 670
rect 2174 674 2180 675
rect 2174 670 2175 674
rect 2179 670 2180 674
rect 2174 669 2180 670
rect 2262 674 2268 675
rect 2262 670 2263 674
rect 2267 670 2268 674
rect 2262 669 2268 670
rect 2358 674 2364 675
rect 2358 670 2359 674
rect 2363 670 2364 674
rect 2358 669 2364 670
rect 2462 674 2468 675
rect 2462 670 2463 674
rect 2467 670 2468 674
rect 2462 669 2468 670
rect 2566 674 2572 675
rect 2566 670 2567 674
rect 2571 670 2572 674
rect 2566 669 2572 670
rect 2678 674 2684 675
rect 2678 670 2679 674
rect 2683 670 2684 674
rect 2678 669 2684 670
rect 2798 674 2804 675
rect 2798 670 2799 674
rect 2803 670 2804 674
rect 2798 669 2804 670
rect 2926 674 2932 675
rect 2926 670 2927 674
rect 2931 670 2932 674
rect 2926 669 2932 670
rect 3070 674 3076 675
rect 3070 670 3071 674
rect 3075 670 3076 674
rect 3070 669 3076 670
rect 3222 674 3228 675
rect 3222 670 3223 674
rect 3227 670 3228 674
rect 3222 669 3228 670
rect 3374 674 3380 675
rect 3374 670 3375 674
rect 3379 670 3380 674
rect 3374 669 3380 670
rect 3510 674 3516 675
rect 3510 670 3511 674
rect 3515 670 3516 674
rect 3510 669 3516 670
rect 3592 657 3594 685
rect 1870 656 1876 657
rect 110 652 116 653
rect 110 648 111 652
rect 115 648 116 652
rect 110 647 116 648
rect 1830 652 1836 653
rect 1830 648 1831 652
rect 1835 648 1836 652
rect 1870 652 1871 656
rect 1875 652 1876 656
rect 1870 651 1876 652
rect 3590 656 3596 657
rect 3590 652 3591 656
rect 3595 652 3596 656
rect 3590 651 3596 652
rect 1830 647 1836 648
rect 1870 639 1876 640
rect 110 635 116 636
rect 110 631 111 635
rect 115 631 116 635
rect 1830 635 1836 636
rect 110 630 116 631
rect 374 632 380 633
rect 112 603 114 630
rect 374 628 375 632
rect 379 628 380 632
rect 374 627 380 628
rect 470 632 476 633
rect 470 628 471 632
rect 475 628 476 632
rect 470 627 476 628
rect 582 632 588 633
rect 582 628 583 632
rect 587 628 588 632
rect 582 627 588 628
rect 710 632 716 633
rect 710 628 711 632
rect 715 628 716 632
rect 710 627 716 628
rect 846 632 852 633
rect 846 628 847 632
rect 851 628 852 632
rect 846 627 852 628
rect 982 632 988 633
rect 982 628 983 632
rect 987 628 988 632
rect 982 627 988 628
rect 1118 632 1124 633
rect 1118 628 1119 632
rect 1123 628 1124 632
rect 1118 627 1124 628
rect 1246 632 1252 633
rect 1246 628 1247 632
rect 1251 628 1252 632
rect 1246 627 1252 628
rect 1374 632 1380 633
rect 1374 628 1375 632
rect 1379 628 1380 632
rect 1374 627 1380 628
rect 1494 632 1500 633
rect 1494 628 1495 632
rect 1499 628 1500 632
rect 1494 627 1500 628
rect 1622 632 1628 633
rect 1622 628 1623 632
rect 1627 628 1628 632
rect 1622 627 1628 628
rect 1742 632 1748 633
rect 1742 628 1743 632
rect 1747 628 1748 632
rect 1830 631 1831 635
rect 1835 631 1836 635
rect 1870 635 1871 639
rect 1875 635 1876 639
rect 3590 639 3596 640
rect 1870 634 1876 635
rect 2086 636 2092 637
rect 1830 630 1836 631
rect 1742 627 1748 628
rect 376 603 378 627
rect 472 603 474 627
rect 584 603 586 627
rect 712 603 714 627
rect 848 603 850 627
rect 984 603 986 627
rect 1120 603 1122 627
rect 1248 603 1250 627
rect 1376 603 1378 627
rect 1496 603 1498 627
rect 1624 603 1626 627
rect 1744 603 1746 627
rect 1832 603 1834 630
rect 1872 603 1874 634
rect 2086 632 2087 636
rect 2091 632 2092 636
rect 2086 631 2092 632
rect 2166 636 2172 637
rect 2166 632 2167 636
rect 2171 632 2172 636
rect 2166 631 2172 632
rect 2254 636 2260 637
rect 2254 632 2255 636
rect 2259 632 2260 636
rect 2254 631 2260 632
rect 2350 636 2356 637
rect 2350 632 2351 636
rect 2355 632 2356 636
rect 2350 631 2356 632
rect 2454 636 2460 637
rect 2454 632 2455 636
rect 2459 632 2460 636
rect 2454 631 2460 632
rect 2558 636 2564 637
rect 2558 632 2559 636
rect 2563 632 2564 636
rect 2558 631 2564 632
rect 2670 636 2676 637
rect 2670 632 2671 636
rect 2675 632 2676 636
rect 2670 631 2676 632
rect 2790 636 2796 637
rect 2790 632 2791 636
rect 2795 632 2796 636
rect 2790 631 2796 632
rect 2918 636 2924 637
rect 2918 632 2919 636
rect 2923 632 2924 636
rect 2918 631 2924 632
rect 3062 636 3068 637
rect 3062 632 3063 636
rect 3067 632 3068 636
rect 3062 631 3068 632
rect 3214 636 3220 637
rect 3214 632 3215 636
rect 3219 632 3220 636
rect 3214 631 3220 632
rect 3366 636 3372 637
rect 3366 632 3367 636
rect 3371 632 3372 636
rect 3366 631 3372 632
rect 3502 636 3508 637
rect 3502 632 3503 636
rect 3507 632 3508 636
rect 3590 635 3591 639
rect 3595 635 3596 639
rect 3590 634 3596 635
rect 3502 631 3508 632
rect 2088 603 2090 631
rect 2168 603 2170 631
rect 2256 603 2258 631
rect 2352 603 2354 631
rect 2456 603 2458 631
rect 2560 603 2562 631
rect 2672 603 2674 631
rect 2792 603 2794 631
rect 2920 603 2922 631
rect 3064 603 3066 631
rect 3216 603 3218 631
rect 3368 603 3370 631
rect 3504 603 3506 631
rect 3592 603 3594 634
rect 111 602 115 603
rect 111 597 115 598
rect 375 602 379 603
rect 375 597 379 598
rect 471 602 475 603
rect 471 597 475 598
rect 583 602 587 603
rect 583 597 587 598
rect 599 602 603 603
rect 599 597 603 598
rect 687 602 691 603
rect 687 597 691 598
rect 711 602 715 603
rect 711 597 715 598
rect 783 602 787 603
rect 783 597 787 598
rect 847 602 851 603
rect 847 597 851 598
rect 887 602 891 603
rect 887 597 891 598
rect 983 602 987 603
rect 983 597 987 598
rect 991 602 995 603
rect 991 597 995 598
rect 1095 602 1099 603
rect 1095 597 1099 598
rect 1119 602 1123 603
rect 1119 597 1123 598
rect 1199 602 1203 603
rect 1199 597 1203 598
rect 1247 602 1251 603
rect 1247 597 1251 598
rect 1303 602 1307 603
rect 1303 597 1307 598
rect 1375 602 1379 603
rect 1375 597 1379 598
rect 1399 602 1403 603
rect 1399 597 1403 598
rect 1495 602 1499 603
rect 1495 597 1499 598
rect 1503 602 1507 603
rect 1503 597 1507 598
rect 1607 602 1611 603
rect 1607 597 1611 598
rect 1623 602 1627 603
rect 1623 597 1627 598
rect 1711 602 1715 603
rect 1711 597 1715 598
rect 1743 602 1747 603
rect 1743 597 1747 598
rect 1831 602 1835 603
rect 1831 597 1835 598
rect 1871 602 1875 603
rect 1871 597 1875 598
rect 2087 602 2091 603
rect 2087 597 2091 598
rect 2167 602 2171 603
rect 2167 597 2171 598
rect 2247 602 2251 603
rect 2247 597 2251 598
rect 2255 602 2259 603
rect 2255 597 2259 598
rect 2327 602 2331 603
rect 2327 597 2331 598
rect 2351 602 2355 603
rect 2351 597 2355 598
rect 2407 602 2411 603
rect 2407 597 2411 598
rect 2455 602 2459 603
rect 2455 597 2459 598
rect 2487 602 2491 603
rect 2487 597 2491 598
rect 2559 602 2563 603
rect 2559 597 2563 598
rect 2567 602 2571 603
rect 2567 597 2571 598
rect 2647 602 2651 603
rect 2647 597 2651 598
rect 2671 602 2675 603
rect 2671 597 2675 598
rect 2743 602 2747 603
rect 2743 597 2747 598
rect 2791 602 2795 603
rect 2791 597 2795 598
rect 2863 602 2867 603
rect 2863 597 2867 598
rect 2919 602 2923 603
rect 2919 597 2923 598
rect 2999 602 3003 603
rect 2999 597 3003 598
rect 3063 602 3067 603
rect 3063 597 3067 598
rect 3159 602 3163 603
rect 3159 597 3163 598
rect 3215 602 3219 603
rect 3215 597 3219 598
rect 3327 602 3331 603
rect 3327 597 3331 598
rect 3367 602 3371 603
rect 3367 597 3371 598
rect 3495 602 3499 603
rect 3495 597 3499 598
rect 3503 602 3507 603
rect 3503 597 3507 598
rect 3591 602 3595 603
rect 3591 597 3595 598
rect 112 578 114 597
rect 600 581 602 597
rect 688 581 690 597
rect 784 581 786 597
rect 888 581 890 597
rect 992 581 994 597
rect 1096 581 1098 597
rect 1200 581 1202 597
rect 1304 581 1306 597
rect 1400 581 1402 597
rect 1504 581 1506 597
rect 1608 581 1610 597
rect 1712 581 1714 597
rect 598 580 604 581
rect 110 577 116 578
rect 110 573 111 577
rect 115 573 116 577
rect 598 576 599 580
rect 603 576 604 580
rect 598 575 604 576
rect 686 580 692 581
rect 686 576 687 580
rect 691 576 692 580
rect 686 575 692 576
rect 782 580 788 581
rect 782 576 783 580
rect 787 576 788 580
rect 782 575 788 576
rect 886 580 892 581
rect 886 576 887 580
rect 891 576 892 580
rect 886 575 892 576
rect 990 580 996 581
rect 990 576 991 580
rect 995 576 996 580
rect 990 575 996 576
rect 1094 580 1100 581
rect 1094 576 1095 580
rect 1099 576 1100 580
rect 1094 575 1100 576
rect 1198 580 1204 581
rect 1198 576 1199 580
rect 1203 576 1204 580
rect 1198 575 1204 576
rect 1302 580 1308 581
rect 1302 576 1303 580
rect 1307 576 1308 580
rect 1302 575 1308 576
rect 1398 580 1404 581
rect 1398 576 1399 580
rect 1403 576 1404 580
rect 1398 575 1404 576
rect 1502 580 1508 581
rect 1502 576 1503 580
rect 1507 576 1508 580
rect 1502 575 1508 576
rect 1606 580 1612 581
rect 1606 576 1607 580
rect 1611 576 1612 580
rect 1606 575 1612 576
rect 1710 580 1716 581
rect 1710 576 1711 580
rect 1715 576 1716 580
rect 1832 578 1834 597
rect 1872 578 1874 597
rect 2168 581 2170 597
rect 2248 581 2250 597
rect 2328 581 2330 597
rect 2408 581 2410 597
rect 2488 581 2490 597
rect 2568 581 2570 597
rect 2648 581 2650 597
rect 2744 581 2746 597
rect 2864 581 2866 597
rect 3000 581 3002 597
rect 3160 581 3162 597
rect 3328 581 3330 597
rect 3496 581 3498 597
rect 2166 580 2172 581
rect 1710 575 1716 576
rect 1830 577 1836 578
rect 110 572 116 573
rect 1830 573 1831 577
rect 1835 573 1836 577
rect 1830 572 1836 573
rect 1870 577 1876 578
rect 1870 573 1871 577
rect 1875 573 1876 577
rect 2166 576 2167 580
rect 2171 576 2172 580
rect 2166 575 2172 576
rect 2246 580 2252 581
rect 2246 576 2247 580
rect 2251 576 2252 580
rect 2246 575 2252 576
rect 2326 580 2332 581
rect 2326 576 2327 580
rect 2331 576 2332 580
rect 2326 575 2332 576
rect 2406 580 2412 581
rect 2406 576 2407 580
rect 2411 576 2412 580
rect 2406 575 2412 576
rect 2486 580 2492 581
rect 2486 576 2487 580
rect 2491 576 2492 580
rect 2486 575 2492 576
rect 2566 580 2572 581
rect 2566 576 2567 580
rect 2571 576 2572 580
rect 2566 575 2572 576
rect 2646 580 2652 581
rect 2646 576 2647 580
rect 2651 576 2652 580
rect 2646 575 2652 576
rect 2742 580 2748 581
rect 2742 576 2743 580
rect 2747 576 2748 580
rect 2742 575 2748 576
rect 2862 580 2868 581
rect 2862 576 2863 580
rect 2867 576 2868 580
rect 2862 575 2868 576
rect 2998 580 3004 581
rect 2998 576 2999 580
rect 3003 576 3004 580
rect 2998 575 3004 576
rect 3158 580 3164 581
rect 3158 576 3159 580
rect 3163 576 3164 580
rect 3158 575 3164 576
rect 3326 580 3332 581
rect 3326 576 3327 580
rect 3331 576 3332 580
rect 3326 575 3332 576
rect 3494 580 3500 581
rect 3494 576 3495 580
rect 3499 576 3500 580
rect 3592 578 3594 597
rect 3494 575 3500 576
rect 3590 577 3596 578
rect 1870 572 1876 573
rect 3590 573 3591 577
rect 3595 573 3596 577
rect 3590 572 3596 573
rect 110 560 116 561
rect 110 556 111 560
rect 115 556 116 560
rect 110 555 116 556
rect 1830 560 1836 561
rect 1830 556 1831 560
rect 1835 556 1836 560
rect 1830 555 1836 556
rect 1870 560 1876 561
rect 1870 556 1871 560
rect 1875 556 1876 560
rect 1870 555 1876 556
rect 3590 560 3596 561
rect 3590 556 3591 560
rect 3595 556 3596 560
rect 3590 555 3596 556
rect 112 519 114 555
rect 606 542 612 543
rect 606 538 607 542
rect 611 538 612 542
rect 606 537 612 538
rect 694 542 700 543
rect 694 538 695 542
rect 699 538 700 542
rect 694 537 700 538
rect 790 542 796 543
rect 790 538 791 542
rect 795 538 796 542
rect 790 537 796 538
rect 894 542 900 543
rect 894 538 895 542
rect 899 538 900 542
rect 894 537 900 538
rect 998 542 1004 543
rect 998 538 999 542
rect 1003 538 1004 542
rect 998 537 1004 538
rect 1102 542 1108 543
rect 1102 538 1103 542
rect 1107 538 1108 542
rect 1102 537 1108 538
rect 1206 542 1212 543
rect 1206 538 1207 542
rect 1211 538 1212 542
rect 1206 537 1212 538
rect 1310 542 1316 543
rect 1310 538 1311 542
rect 1315 538 1316 542
rect 1310 537 1316 538
rect 1406 542 1412 543
rect 1406 538 1407 542
rect 1411 538 1412 542
rect 1406 537 1412 538
rect 1510 542 1516 543
rect 1510 538 1511 542
rect 1515 538 1516 542
rect 1510 537 1516 538
rect 1614 542 1620 543
rect 1614 538 1615 542
rect 1619 538 1620 542
rect 1614 537 1620 538
rect 1718 542 1724 543
rect 1718 538 1719 542
rect 1723 538 1724 542
rect 1718 537 1724 538
rect 608 519 610 537
rect 696 519 698 537
rect 792 519 794 537
rect 896 519 898 537
rect 1000 519 1002 537
rect 1104 519 1106 537
rect 1208 519 1210 537
rect 1312 519 1314 537
rect 1408 519 1410 537
rect 1512 519 1514 537
rect 1616 519 1618 537
rect 1720 519 1722 537
rect 1832 519 1834 555
rect 1872 519 1874 555
rect 2174 542 2180 543
rect 2174 538 2175 542
rect 2179 538 2180 542
rect 2174 537 2180 538
rect 2254 542 2260 543
rect 2254 538 2255 542
rect 2259 538 2260 542
rect 2254 537 2260 538
rect 2334 542 2340 543
rect 2334 538 2335 542
rect 2339 538 2340 542
rect 2334 537 2340 538
rect 2414 542 2420 543
rect 2414 538 2415 542
rect 2419 538 2420 542
rect 2414 537 2420 538
rect 2494 542 2500 543
rect 2494 538 2495 542
rect 2499 538 2500 542
rect 2494 537 2500 538
rect 2574 542 2580 543
rect 2574 538 2575 542
rect 2579 538 2580 542
rect 2574 537 2580 538
rect 2654 542 2660 543
rect 2654 538 2655 542
rect 2659 538 2660 542
rect 2654 537 2660 538
rect 2750 542 2756 543
rect 2750 538 2751 542
rect 2755 538 2756 542
rect 2750 537 2756 538
rect 2870 542 2876 543
rect 2870 538 2871 542
rect 2875 538 2876 542
rect 2870 537 2876 538
rect 3006 542 3012 543
rect 3006 538 3007 542
rect 3011 538 3012 542
rect 3006 537 3012 538
rect 3166 542 3172 543
rect 3166 538 3167 542
rect 3171 538 3172 542
rect 3166 537 3172 538
rect 3334 542 3340 543
rect 3334 538 3335 542
rect 3339 538 3340 542
rect 3334 537 3340 538
rect 3502 542 3508 543
rect 3502 538 3503 542
rect 3507 538 3508 542
rect 3502 537 3508 538
rect 2176 519 2178 537
rect 2256 519 2258 537
rect 2336 519 2338 537
rect 2416 519 2418 537
rect 2496 519 2498 537
rect 2576 519 2578 537
rect 2656 519 2658 537
rect 2752 519 2754 537
rect 2872 519 2874 537
rect 3008 519 3010 537
rect 3168 519 3170 537
rect 3336 519 3338 537
rect 3504 519 3506 537
rect 3592 519 3594 555
rect 111 518 115 519
rect 111 513 115 514
rect 367 518 371 519
rect 367 513 371 514
rect 463 518 467 519
rect 463 513 467 514
rect 575 518 579 519
rect 575 513 579 514
rect 607 518 611 519
rect 607 513 611 514
rect 695 518 699 519
rect 695 513 699 514
rect 703 518 707 519
rect 703 513 707 514
rect 791 518 795 519
rect 791 513 795 514
rect 839 518 843 519
rect 839 513 843 514
rect 895 518 899 519
rect 895 513 899 514
rect 975 518 979 519
rect 975 513 979 514
rect 999 518 1003 519
rect 999 513 1003 514
rect 1103 518 1107 519
rect 1103 513 1107 514
rect 1111 518 1115 519
rect 1111 513 1115 514
rect 1207 518 1211 519
rect 1207 513 1211 514
rect 1239 518 1243 519
rect 1239 513 1243 514
rect 1311 518 1315 519
rect 1311 513 1315 514
rect 1359 518 1363 519
rect 1359 513 1363 514
rect 1407 518 1411 519
rect 1407 513 1411 514
rect 1471 518 1475 519
rect 1471 513 1475 514
rect 1511 518 1515 519
rect 1511 513 1515 514
rect 1583 518 1587 519
rect 1583 513 1587 514
rect 1615 518 1619 519
rect 1615 513 1619 514
rect 1703 518 1707 519
rect 1703 513 1707 514
rect 1719 518 1723 519
rect 1719 513 1723 514
rect 1831 518 1835 519
rect 1831 513 1835 514
rect 1871 518 1875 519
rect 1871 513 1875 514
rect 2159 518 2163 519
rect 2159 513 2163 514
rect 2175 518 2179 519
rect 2175 513 2179 514
rect 2239 518 2243 519
rect 2239 513 2243 514
rect 2255 518 2259 519
rect 2255 513 2259 514
rect 2319 518 2323 519
rect 2319 513 2323 514
rect 2335 518 2339 519
rect 2335 513 2339 514
rect 2399 518 2403 519
rect 2399 513 2403 514
rect 2415 518 2419 519
rect 2415 513 2419 514
rect 2479 518 2483 519
rect 2479 513 2483 514
rect 2495 518 2499 519
rect 2495 513 2499 514
rect 2559 518 2563 519
rect 2559 513 2563 514
rect 2575 518 2579 519
rect 2575 513 2579 514
rect 2639 518 2643 519
rect 2639 513 2643 514
rect 2655 518 2659 519
rect 2655 513 2659 514
rect 2735 518 2739 519
rect 2735 513 2739 514
rect 2751 518 2755 519
rect 2751 513 2755 514
rect 2855 518 2859 519
rect 2855 513 2859 514
rect 2871 518 2875 519
rect 2871 513 2875 514
rect 2991 518 2995 519
rect 2991 513 2995 514
rect 3007 518 3011 519
rect 3007 513 3011 514
rect 3143 518 3147 519
rect 3143 513 3147 514
rect 3167 518 3171 519
rect 3167 513 3171 514
rect 3311 518 3315 519
rect 3311 513 3315 514
rect 3335 518 3339 519
rect 3335 513 3339 514
rect 3479 518 3483 519
rect 3479 513 3483 514
rect 3503 518 3507 519
rect 3503 513 3507 514
rect 3591 518 3595 519
rect 3591 513 3595 514
rect 112 485 114 513
rect 368 503 370 513
rect 464 503 466 513
rect 576 503 578 513
rect 704 503 706 513
rect 840 503 842 513
rect 976 503 978 513
rect 1112 503 1114 513
rect 1240 503 1242 513
rect 1360 503 1362 513
rect 1472 503 1474 513
rect 1584 503 1586 513
rect 1704 503 1706 513
rect 366 502 372 503
rect 366 498 367 502
rect 371 498 372 502
rect 366 497 372 498
rect 462 502 468 503
rect 462 498 463 502
rect 467 498 468 502
rect 462 497 468 498
rect 574 502 580 503
rect 574 498 575 502
rect 579 498 580 502
rect 574 497 580 498
rect 702 502 708 503
rect 702 498 703 502
rect 707 498 708 502
rect 702 497 708 498
rect 838 502 844 503
rect 838 498 839 502
rect 843 498 844 502
rect 838 497 844 498
rect 974 502 980 503
rect 974 498 975 502
rect 979 498 980 502
rect 974 497 980 498
rect 1110 502 1116 503
rect 1110 498 1111 502
rect 1115 498 1116 502
rect 1110 497 1116 498
rect 1238 502 1244 503
rect 1238 498 1239 502
rect 1243 498 1244 502
rect 1238 497 1244 498
rect 1358 502 1364 503
rect 1358 498 1359 502
rect 1363 498 1364 502
rect 1358 497 1364 498
rect 1470 502 1476 503
rect 1470 498 1471 502
rect 1475 498 1476 502
rect 1470 497 1476 498
rect 1582 502 1588 503
rect 1582 498 1583 502
rect 1587 498 1588 502
rect 1582 497 1588 498
rect 1702 502 1708 503
rect 1702 498 1703 502
rect 1707 498 1708 502
rect 1702 497 1708 498
rect 1832 485 1834 513
rect 1872 485 1874 513
rect 2160 503 2162 513
rect 2240 503 2242 513
rect 2320 503 2322 513
rect 2400 503 2402 513
rect 2480 503 2482 513
rect 2560 503 2562 513
rect 2640 503 2642 513
rect 2736 503 2738 513
rect 2856 503 2858 513
rect 2992 503 2994 513
rect 3144 503 3146 513
rect 3312 503 3314 513
rect 3480 503 3482 513
rect 2158 502 2164 503
rect 2158 498 2159 502
rect 2163 498 2164 502
rect 2158 497 2164 498
rect 2238 502 2244 503
rect 2238 498 2239 502
rect 2243 498 2244 502
rect 2238 497 2244 498
rect 2318 502 2324 503
rect 2318 498 2319 502
rect 2323 498 2324 502
rect 2318 497 2324 498
rect 2398 502 2404 503
rect 2398 498 2399 502
rect 2403 498 2404 502
rect 2398 497 2404 498
rect 2478 502 2484 503
rect 2478 498 2479 502
rect 2483 498 2484 502
rect 2478 497 2484 498
rect 2558 502 2564 503
rect 2558 498 2559 502
rect 2563 498 2564 502
rect 2558 497 2564 498
rect 2638 502 2644 503
rect 2638 498 2639 502
rect 2643 498 2644 502
rect 2638 497 2644 498
rect 2734 502 2740 503
rect 2734 498 2735 502
rect 2739 498 2740 502
rect 2734 497 2740 498
rect 2854 502 2860 503
rect 2854 498 2855 502
rect 2859 498 2860 502
rect 2854 497 2860 498
rect 2990 502 2996 503
rect 2990 498 2991 502
rect 2995 498 2996 502
rect 2990 497 2996 498
rect 3142 502 3148 503
rect 3142 498 3143 502
rect 3147 498 3148 502
rect 3142 497 3148 498
rect 3310 502 3316 503
rect 3310 498 3311 502
rect 3315 498 3316 502
rect 3310 497 3316 498
rect 3478 502 3484 503
rect 3478 498 3479 502
rect 3483 498 3484 502
rect 3478 497 3484 498
rect 3592 485 3594 513
rect 110 484 116 485
rect 110 480 111 484
rect 115 480 116 484
rect 110 479 116 480
rect 1830 484 1836 485
rect 1830 480 1831 484
rect 1835 480 1836 484
rect 1830 479 1836 480
rect 1870 484 1876 485
rect 1870 480 1871 484
rect 1875 480 1876 484
rect 1870 479 1876 480
rect 3590 484 3596 485
rect 3590 480 3591 484
rect 3595 480 3596 484
rect 3590 479 3596 480
rect 110 467 116 468
rect 110 463 111 467
rect 115 463 116 467
rect 1830 467 1836 468
rect 110 462 116 463
rect 358 464 364 465
rect 112 431 114 462
rect 358 460 359 464
rect 363 460 364 464
rect 358 459 364 460
rect 454 464 460 465
rect 454 460 455 464
rect 459 460 460 464
rect 454 459 460 460
rect 566 464 572 465
rect 566 460 567 464
rect 571 460 572 464
rect 566 459 572 460
rect 694 464 700 465
rect 694 460 695 464
rect 699 460 700 464
rect 694 459 700 460
rect 830 464 836 465
rect 830 460 831 464
rect 835 460 836 464
rect 830 459 836 460
rect 966 464 972 465
rect 966 460 967 464
rect 971 460 972 464
rect 966 459 972 460
rect 1102 464 1108 465
rect 1102 460 1103 464
rect 1107 460 1108 464
rect 1102 459 1108 460
rect 1230 464 1236 465
rect 1230 460 1231 464
rect 1235 460 1236 464
rect 1230 459 1236 460
rect 1350 464 1356 465
rect 1350 460 1351 464
rect 1355 460 1356 464
rect 1350 459 1356 460
rect 1462 464 1468 465
rect 1462 460 1463 464
rect 1467 460 1468 464
rect 1462 459 1468 460
rect 1574 464 1580 465
rect 1574 460 1575 464
rect 1579 460 1580 464
rect 1574 459 1580 460
rect 1694 464 1700 465
rect 1694 460 1695 464
rect 1699 460 1700 464
rect 1830 463 1831 467
rect 1835 463 1836 467
rect 1830 462 1836 463
rect 1870 467 1876 468
rect 1870 463 1871 467
rect 1875 463 1876 467
rect 3590 467 3596 468
rect 1870 462 1876 463
rect 2150 464 2156 465
rect 1694 459 1700 460
rect 360 431 362 459
rect 456 431 458 459
rect 568 431 570 459
rect 696 431 698 459
rect 832 431 834 459
rect 968 431 970 459
rect 1104 431 1106 459
rect 1232 431 1234 459
rect 1352 431 1354 459
rect 1464 431 1466 459
rect 1576 431 1578 459
rect 1696 431 1698 459
rect 1832 431 1834 462
rect 1872 431 1874 462
rect 2150 460 2151 464
rect 2155 460 2156 464
rect 2150 459 2156 460
rect 2230 464 2236 465
rect 2230 460 2231 464
rect 2235 460 2236 464
rect 2230 459 2236 460
rect 2310 464 2316 465
rect 2310 460 2311 464
rect 2315 460 2316 464
rect 2310 459 2316 460
rect 2390 464 2396 465
rect 2390 460 2391 464
rect 2395 460 2396 464
rect 2390 459 2396 460
rect 2470 464 2476 465
rect 2470 460 2471 464
rect 2475 460 2476 464
rect 2470 459 2476 460
rect 2550 464 2556 465
rect 2550 460 2551 464
rect 2555 460 2556 464
rect 2550 459 2556 460
rect 2630 464 2636 465
rect 2630 460 2631 464
rect 2635 460 2636 464
rect 2630 459 2636 460
rect 2726 464 2732 465
rect 2726 460 2727 464
rect 2731 460 2732 464
rect 2726 459 2732 460
rect 2846 464 2852 465
rect 2846 460 2847 464
rect 2851 460 2852 464
rect 2846 459 2852 460
rect 2982 464 2988 465
rect 2982 460 2983 464
rect 2987 460 2988 464
rect 2982 459 2988 460
rect 3134 464 3140 465
rect 3134 460 3135 464
rect 3139 460 3140 464
rect 3134 459 3140 460
rect 3302 464 3308 465
rect 3302 460 3303 464
rect 3307 460 3308 464
rect 3302 459 3308 460
rect 3470 464 3476 465
rect 3470 460 3471 464
rect 3475 460 3476 464
rect 3590 463 3591 467
rect 3595 463 3596 467
rect 3590 462 3596 463
rect 3470 459 3476 460
rect 2152 431 2154 459
rect 2232 431 2234 459
rect 2312 431 2314 459
rect 2392 431 2394 459
rect 2472 431 2474 459
rect 2552 431 2554 459
rect 2632 431 2634 459
rect 2728 431 2730 459
rect 2848 431 2850 459
rect 2984 431 2986 459
rect 3136 431 3138 459
rect 3304 431 3306 459
rect 3472 431 3474 459
rect 3592 431 3594 462
rect 111 430 115 431
rect 111 425 115 426
rect 135 430 139 431
rect 135 425 139 426
rect 223 430 227 431
rect 223 425 227 426
rect 359 430 363 431
rect 359 425 363 426
rect 455 430 459 431
rect 455 425 459 426
rect 511 430 515 431
rect 511 425 515 426
rect 567 430 571 431
rect 567 425 571 426
rect 679 430 683 431
rect 679 425 683 426
rect 695 430 699 431
rect 695 425 699 426
rect 831 430 835 431
rect 831 425 835 426
rect 839 430 843 431
rect 839 425 843 426
rect 967 430 971 431
rect 967 425 971 426
rect 999 430 1003 431
rect 999 425 1003 426
rect 1103 430 1107 431
rect 1103 425 1107 426
rect 1143 430 1147 431
rect 1143 425 1147 426
rect 1231 430 1235 431
rect 1231 425 1235 426
rect 1279 430 1283 431
rect 1279 425 1283 426
rect 1351 430 1355 431
rect 1351 425 1355 426
rect 1415 430 1419 431
rect 1415 425 1419 426
rect 1463 430 1467 431
rect 1463 425 1467 426
rect 1551 430 1555 431
rect 1551 425 1555 426
rect 1575 430 1579 431
rect 1575 425 1579 426
rect 1687 430 1691 431
rect 1687 425 1691 426
rect 1695 430 1699 431
rect 1695 425 1699 426
rect 1831 430 1835 431
rect 1831 425 1835 426
rect 1871 430 1875 431
rect 1871 425 1875 426
rect 2151 430 2155 431
rect 2151 425 2155 426
rect 2159 430 2163 431
rect 2159 425 2163 426
rect 2231 430 2235 431
rect 2231 425 2235 426
rect 2239 430 2243 431
rect 2239 425 2243 426
rect 2311 430 2315 431
rect 2311 425 2315 426
rect 2319 430 2323 431
rect 2319 425 2323 426
rect 2391 430 2395 431
rect 2391 425 2395 426
rect 2399 430 2403 431
rect 2399 425 2403 426
rect 2471 430 2475 431
rect 2471 425 2475 426
rect 2479 430 2483 431
rect 2479 425 2483 426
rect 2551 430 2555 431
rect 2551 425 2555 426
rect 2559 430 2563 431
rect 2559 425 2563 426
rect 2631 430 2635 431
rect 2631 425 2635 426
rect 2639 430 2643 431
rect 2639 425 2643 426
rect 2727 430 2731 431
rect 2727 425 2731 426
rect 2735 430 2739 431
rect 2735 425 2739 426
rect 2839 430 2843 431
rect 2839 425 2843 426
rect 2847 430 2851 431
rect 2847 425 2851 426
rect 2959 430 2963 431
rect 2959 425 2963 426
rect 2983 430 2987 431
rect 2983 425 2987 426
rect 3087 430 3091 431
rect 3087 425 3091 426
rect 3135 430 3139 431
rect 3135 425 3139 426
rect 3231 430 3235 431
rect 3231 425 3235 426
rect 3303 430 3307 431
rect 3303 425 3307 426
rect 3375 430 3379 431
rect 3375 425 3379 426
rect 3471 430 3475 431
rect 3471 425 3475 426
rect 3503 430 3507 431
rect 3503 425 3507 426
rect 3591 430 3595 431
rect 3591 425 3595 426
rect 112 406 114 425
rect 136 409 138 425
rect 224 409 226 425
rect 360 409 362 425
rect 512 409 514 425
rect 680 409 682 425
rect 840 409 842 425
rect 1000 409 1002 425
rect 1144 409 1146 425
rect 1280 409 1282 425
rect 1416 409 1418 425
rect 1552 409 1554 425
rect 1688 409 1690 425
rect 134 408 140 409
rect 110 405 116 406
rect 110 401 111 405
rect 115 401 116 405
rect 134 404 135 408
rect 139 404 140 408
rect 134 403 140 404
rect 222 408 228 409
rect 222 404 223 408
rect 227 404 228 408
rect 222 403 228 404
rect 358 408 364 409
rect 358 404 359 408
rect 363 404 364 408
rect 358 403 364 404
rect 510 408 516 409
rect 510 404 511 408
rect 515 404 516 408
rect 510 403 516 404
rect 678 408 684 409
rect 678 404 679 408
rect 683 404 684 408
rect 678 403 684 404
rect 838 408 844 409
rect 838 404 839 408
rect 843 404 844 408
rect 838 403 844 404
rect 998 408 1004 409
rect 998 404 999 408
rect 1003 404 1004 408
rect 998 403 1004 404
rect 1142 408 1148 409
rect 1142 404 1143 408
rect 1147 404 1148 408
rect 1142 403 1148 404
rect 1278 408 1284 409
rect 1278 404 1279 408
rect 1283 404 1284 408
rect 1278 403 1284 404
rect 1414 408 1420 409
rect 1414 404 1415 408
rect 1419 404 1420 408
rect 1414 403 1420 404
rect 1550 408 1556 409
rect 1550 404 1551 408
rect 1555 404 1556 408
rect 1550 403 1556 404
rect 1686 408 1692 409
rect 1686 404 1687 408
rect 1691 404 1692 408
rect 1832 406 1834 425
rect 1872 406 1874 425
rect 2160 409 2162 425
rect 2240 409 2242 425
rect 2320 409 2322 425
rect 2400 409 2402 425
rect 2480 409 2482 425
rect 2560 409 2562 425
rect 2640 409 2642 425
rect 2736 409 2738 425
rect 2840 409 2842 425
rect 2960 409 2962 425
rect 3088 409 3090 425
rect 3232 409 3234 425
rect 3376 409 3378 425
rect 3504 409 3506 425
rect 2158 408 2164 409
rect 1686 403 1692 404
rect 1830 405 1836 406
rect 110 400 116 401
rect 1830 401 1831 405
rect 1835 401 1836 405
rect 1830 400 1836 401
rect 1870 405 1876 406
rect 1870 401 1871 405
rect 1875 401 1876 405
rect 2158 404 2159 408
rect 2163 404 2164 408
rect 2158 403 2164 404
rect 2238 408 2244 409
rect 2238 404 2239 408
rect 2243 404 2244 408
rect 2238 403 2244 404
rect 2318 408 2324 409
rect 2318 404 2319 408
rect 2323 404 2324 408
rect 2318 403 2324 404
rect 2398 408 2404 409
rect 2398 404 2399 408
rect 2403 404 2404 408
rect 2398 403 2404 404
rect 2478 408 2484 409
rect 2478 404 2479 408
rect 2483 404 2484 408
rect 2478 403 2484 404
rect 2558 408 2564 409
rect 2558 404 2559 408
rect 2563 404 2564 408
rect 2558 403 2564 404
rect 2638 408 2644 409
rect 2638 404 2639 408
rect 2643 404 2644 408
rect 2638 403 2644 404
rect 2734 408 2740 409
rect 2734 404 2735 408
rect 2739 404 2740 408
rect 2734 403 2740 404
rect 2838 408 2844 409
rect 2838 404 2839 408
rect 2843 404 2844 408
rect 2838 403 2844 404
rect 2958 408 2964 409
rect 2958 404 2959 408
rect 2963 404 2964 408
rect 2958 403 2964 404
rect 3086 408 3092 409
rect 3086 404 3087 408
rect 3091 404 3092 408
rect 3086 403 3092 404
rect 3230 408 3236 409
rect 3230 404 3231 408
rect 3235 404 3236 408
rect 3230 403 3236 404
rect 3374 408 3380 409
rect 3374 404 3375 408
rect 3379 404 3380 408
rect 3374 403 3380 404
rect 3502 408 3508 409
rect 3502 404 3503 408
rect 3507 404 3508 408
rect 3592 406 3594 425
rect 3502 403 3508 404
rect 3590 405 3596 406
rect 1870 400 1876 401
rect 3590 401 3591 405
rect 3595 401 3596 405
rect 3590 400 3596 401
rect 110 388 116 389
rect 110 384 111 388
rect 115 384 116 388
rect 110 383 116 384
rect 1830 388 1836 389
rect 1830 384 1831 388
rect 1835 384 1836 388
rect 1830 383 1836 384
rect 1870 388 1876 389
rect 1870 384 1871 388
rect 1875 384 1876 388
rect 1870 383 1876 384
rect 3590 388 3596 389
rect 3590 384 3591 388
rect 3595 384 3596 388
rect 3590 383 3596 384
rect 112 347 114 383
rect 142 370 148 371
rect 142 366 143 370
rect 147 366 148 370
rect 142 365 148 366
rect 230 370 236 371
rect 230 366 231 370
rect 235 366 236 370
rect 230 365 236 366
rect 366 370 372 371
rect 366 366 367 370
rect 371 366 372 370
rect 366 365 372 366
rect 518 370 524 371
rect 518 366 519 370
rect 523 366 524 370
rect 518 365 524 366
rect 686 370 692 371
rect 686 366 687 370
rect 691 366 692 370
rect 686 365 692 366
rect 846 370 852 371
rect 846 366 847 370
rect 851 366 852 370
rect 846 365 852 366
rect 1006 370 1012 371
rect 1006 366 1007 370
rect 1011 366 1012 370
rect 1006 365 1012 366
rect 1150 370 1156 371
rect 1150 366 1151 370
rect 1155 366 1156 370
rect 1150 365 1156 366
rect 1286 370 1292 371
rect 1286 366 1287 370
rect 1291 366 1292 370
rect 1286 365 1292 366
rect 1422 370 1428 371
rect 1422 366 1423 370
rect 1427 366 1428 370
rect 1422 365 1428 366
rect 1558 370 1564 371
rect 1558 366 1559 370
rect 1563 366 1564 370
rect 1558 365 1564 366
rect 1694 370 1700 371
rect 1694 366 1695 370
rect 1699 366 1700 370
rect 1694 365 1700 366
rect 144 347 146 365
rect 232 347 234 365
rect 368 347 370 365
rect 520 347 522 365
rect 688 347 690 365
rect 848 347 850 365
rect 1008 347 1010 365
rect 1152 347 1154 365
rect 1288 347 1290 365
rect 1424 347 1426 365
rect 1560 347 1562 365
rect 1696 347 1698 365
rect 1832 347 1834 383
rect 111 346 115 347
rect 111 341 115 342
rect 143 346 147 347
rect 143 341 147 342
rect 231 346 235 347
rect 231 341 235 342
rect 279 346 283 347
rect 279 341 283 342
rect 367 346 371 347
rect 367 341 371 342
rect 455 346 459 347
rect 455 341 459 342
rect 519 346 523 347
rect 519 341 523 342
rect 639 346 643 347
rect 639 341 643 342
rect 687 346 691 347
rect 687 341 691 342
rect 823 346 827 347
rect 823 341 827 342
rect 847 346 851 347
rect 847 341 851 342
rect 999 346 1003 347
rect 999 341 1003 342
rect 1007 346 1011 347
rect 1007 341 1011 342
rect 1151 346 1155 347
rect 1151 341 1155 342
rect 1167 346 1171 347
rect 1167 341 1171 342
rect 1287 346 1291 347
rect 1287 341 1291 342
rect 1327 346 1331 347
rect 1327 341 1331 342
rect 1423 346 1427 347
rect 1423 341 1427 342
rect 1479 346 1483 347
rect 1479 341 1483 342
rect 1559 346 1563 347
rect 1559 341 1563 342
rect 1623 346 1627 347
rect 1623 341 1627 342
rect 1695 346 1699 347
rect 1695 341 1699 342
rect 1751 346 1755 347
rect 1751 341 1755 342
rect 1831 346 1835 347
rect 1872 343 1874 383
rect 2166 370 2172 371
rect 2166 366 2167 370
rect 2171 366 2172 370
rect 2166 365 2172 366
rect 2246 370 2252 371
rect 2246 366 2247 370
rect 2251 366 2252 370
rect 2246 365 2252 366
rect 2326 370 2332 371
rect 2326 366 2327 370
rect 2331 366 2332 370
rect 2326 365 2332 366
rect 2406 370 2412 371
rect 2406 366 2407 370
rect 2411 366 2412 370
rect 2406 365 2412 366
rect 2486 370 2492 371
rect 2486 366 2487 370
rect 2491 366 2492 370
rect 2486 365 2492 366
rect 2566 370 2572 371
rect 2566 366 2567 370
rect 2571 366 2572 370
rect 2566 365 2572 366
rect 2646 370 2652 371
rect 2646 366 2647 370
rect 2651 366 2652 370
rect 2646 365 2652 366
rect 2742 370 2748 371
rect 2742 366 2743 370
rect 2747 366 2748 370
rect 2742 365 2748 366
rect 2846 370 2852 371
rect 2846 366 2847 370
rect 2851 366 2852 370
rect 2846 365 2852 366
rect 2966 370 2972 371
rect 2966 366 2967 370
rect 2971 366 2972 370
rect 2966 365 2972 366
rect 3094 370 3100 371
rect 3094 366 3095 370
rect 3099 366 3100 370
rect 3094 365 3100 366
rect 3238 370 3244 371
rect 3238 366 3239 370
rect 3243 366 3244 370
rect 3238 365 3244 366
rect 3382 370 3388 371
rect 3382 366 3383 370
rect 3387 366 3388 370
rect 3382 365 3388 366
rect 3510 370 3516 371
rect 3510 366 3511 370
rect 3515 366 3516 370
rect 3510 365 3516 366
rect 2168 343 2170 365
rect 2248 343 2250 365
rect 2328 343 2330 365
rect 2408 343 2410 365
rect 2488 343 2490 365
rect 2568 343 2570 365
rect 2648 343 2650 365
rect 2744 343 2746 365
rect 2848 343 2850 365
rect 2968 343 2970 365
rect 3096 343 3098 365
rect 3240 343 3242 365
rect 3384 343 3386 365
rect 3512 343 3514 365
rect 3592 343 3594 383
rect 1831 341 1835 342
rect 1871 342 1875 343
rect 112 313 114 341
rect 144 331 146 341
rect 280 331 282 341
rect 456 331 458 341
rect 640 331 642 341
rect 824 331 826 341
rect 1000 331 1002 341
rect 1168 331 1170 341
rect 1328 331 1330 341
rect 1480 331 1482 341
rect 1624 331 1626 341
rect 1752 331 1754 341
rect 142 330 148 331
rect 142 326 143 330
rect 147 326 148 330
rect 142 325 148 326
rect 278 330 284 331
rect 278 326 279 330
rect 283 326 284 330
rect 278 325 284 326
rect 454 330 460 331
rect 454 326 455 330
rect 459 326 460 330
rect 454 325 460 326
rect 638 330 644 331
rect 638 326 639 330
rect 643 326 644 330
rect 638 325 644 326
rect 822 330 828 331
rect 822 326 823 330
rect 827 326 828 330
rect 822 325 828 326
rect 998 330 1004 331
rect 998 326 999 330
rect 1003 326 1004 330
rect 998 325 1004 326
rect 1166 330 1172 331
rect 1166 326 1167 330
rect 1171 326 1172 330
rect 1166 325 1172 326
rect 1326 330 1332 331
rect 1326 326 1327 330
rect 1331 326 1332 330
rect 1326 325 1332 326
rect 1478 330 1484 331
rect 1478 326 1479 330
rect 1483 326 1484 330
rect 1478 325 1484 326
rect 1622 330 1628 331
rect 1622 326 1623 330
rect 1627 326 1628 330
rect 1622 325 1628 326
rect 1750 330 1756 331
rect 1750 326 1751 330
rect 1755 326 1756 330
rect 1750 325 1756 326
rect 1832 313 1834 341
rect 1871 337 1875 338
rect 2031 342 2035 343
rect 2031 337 2035 338
rect 2119 342 2123 343
rect 2119 337 2123 338
rect 2167 342 2171 343
rect 2167 337 2171 338
rect 2223 342 2227 343
rect 2223 337 2227 338
rect 2247 342 2251 343
rect 2247 337 2251 338
rect 2327 342 2331 343
rect 2327 337 2331 338
rect 2335 342 2339 343
rect 2335 337 2339 338
rect 2407 342 2411 343
rect 2407 337 2411 338
rect 2447 342 2451 343
rect 2447 337 2451 338
rect 2487 342 2491 343
rect 2487 337 2491 338
rect 2567 342 2571 343
rect 2567 337 2571 338
rect 2647 342 2651 343
rect 2647 337 2651 338
rect 2695 342 2699 343
rect 2695 337 2699 338
rect 2743 342 2747 343
rect 2743 337 2747 338
rect 2839 342 2843 343
rect 2839 337 2843 338
rect 2847 342 2851 343
rect 2847 337 2851 338
rect 2967 342 2971 343
rect 2967 337 2971 338
rect 2999 342 3003 343
rect 2999 337 3003 338
rect 3095 342 3099 343
rect 3095 337 3099 338
rect 3167 342 3171 343
rect 3167 337 3171 338
rect 3239 342 3243 343
rect 3239 337 3243 338
rect 3343 342 3347 343
rect 3343 337 3347 338
rect 3383 342 3387 343
rect 3383 337 3387 338
rect 3511 342 3515 343
rect 3511 337 3515 338
rect 3591 342 3595 343
rect 3591 337 3595 338
rect 110 312 116 313
rect 110 308 111 312
rect 115 308 116 312
rect 110 307 116 308
rect 1830 312 1836 313
rect 1830 308 1831 312
rect 1835 308 1836 312
rect 1872 309 1874 337
rect 2032 327 2034 337
rect 2120 327 2122 337
rect 2224 327 2226 337
rect 2336 327 2338 337
rect 2448 327 2450 337
rect 2568 327 2570 337
rect 2696 327 2698 337
rect 2840 327 2842 337
rect 3000 327 3002 337
rect 3168 327 3170 337
rect 3344 327 3346 337
rect 3512 327 3514 337
rect 2030 326 2036 327
rect 2030 322 2031 326
rect 2035 322 2036 326
rect 2030 321 2036 322
rect 2118 326 2124 327
rect 2118 322 2119 326
rect 2123 322 2124 326
rect 2118 321 2124 322
rect 2222 326 2228 327
rect 2222 322 2223 326
rect 2227 322 2228 326
rect 2222 321 2228 322
rect 2334 326 2340 327
rect 2334 322 2335 326
rect 2339 322 2340 326
rect 2334 321 2340 322
rect 2446 326 2452 327
rect 2446 322 2447 326
rect 2451 322 2452 326
rect 2446 321 2452 322
rect 2566 326 2572 327
rect 2566 322 2567 326
rect 2571 322 2572 326
rect 2566 321 2572 322
rect 2694 326 2700 327
rect 2694 322 2695 326
rect 2699 322 2700 326
rect 2694 321 2700 322
rect 2838 326 2844 327
rect 2838 322 2839 326
rect 2843 322 2844 326
rect 2838 321 2844 322
rect 2998 326 3004 327
rect 2998 322 2999 326
rect 3003 322 3004 326
rect 2998 321 3004 322
rect 3166 326 3172 327
rect 3166 322 3167 326
rect 3171 322 3172 326
rect 3166 321 3172 322
rect 3342 326 3348 327
rect 3342 322 3343 326
rect 3347 322 3348 326
rect 3342 321 3348 322
rect 3510 326 3516 327
rect 3510 322 3511 326
rect 3515 322 3516 326
rect 3510 321 3516 322
rect 3592 309 3594 337
rect 1830 307 1836 308
rect 1870 308 1876 309
rect 1870 304 1871 308
rect 1875 304 1876 308
rect 1870 303 1876 304
rect 3590 308 3596 309
rect 3590 304 3591 308
rect 3595 304 3596 308
rect 3590 303 3596 304
rect 110 295 116 296
rect 110 291 111 295
rect 115 291 116 295
rect 1830 295 1836 296
rect 110 290 116 291
rect 134 292 140 293
rect 112 267 114 290
rect 134 288 135 292
rect 139 288 140 292
rect 134 287 140 288
rect 270 292 276 293
rect 270 288 271 292
rect 275 288 276 292
rect 270 287 276 288
rect 446 292 452 293
rect 446 288 447 292
rect 451 288 452 292
rect 446 287 452 288
rect 630 292 636 293
rect 630 288 631 292
rect 635 288 636 292
rect 630 287 636 288
rect 814 292 820 293
rect 814 288 815 292
rect 819 288 820 292
rect 814 287 820 288
rect 990 292 996 293
rect 990 288 991 292
rect 995 288 996 292
rect 990 287 996 288
rect 1158 292 1164 293
rect 1158 288 1159 292
rect 1163 288 1164 292
rect 1158 287 1164 288
rect 1318 292 1324 293
rect 1318 288 1319 292
rect 1323 288 1324 292
rect 1318 287 1324 288
rect 1470 292 1476 293
rect 1470 288 1471 292
rect 1475 288 1476 292
rect 1470 287 1476 288
rect 1614 292 1620 293
rect 1614 288 1615 292
rect 1619 288 1620 292
rect 1614 287 1620 288
rect 1742 292 1748 293
rect 1742 288 1743 292
rect 1747 288 1748 292
rect 1830 291 1831 295
rect 1835 291 1836 295
rect 1830 290 1836 291
rect 1870 291 1876 292
rect 1742 287 1748 288
rect 136 267 138 287
rect 272 267 274 287
rect 448 267 450 287
rect 632 267 634 287
rect 816 267 818 287
rect 992 267 994 287
rect 1160 267 1162 287
rect 1320 267 1322 287
rect 1472 267 1474 287
rect 1616 267 1618 287
rect 1744 267 1746 287
rect 1832 267 1834 290
rect 1870 287 1871 291
rect 1875 287 1876 291
rect 3590 291 3596 292
rect 1870 286 1876 287
rect 2022 288 2028 289
rect 111 266 115 267
rect 111 261 115 262
rect 135 266 139 267
rect 135 261 139 262
rect 271 266 275 267
rect 271 261 275 262
rect 303 266 307 267
rect 303 261 307 262
rect 391 266 395 267
rect 391 261 395 262
rect 447 266 451 267
rect 447 261 451 262
rect 495 266 499 267
rect 495 261 499 262
rect 599 266 603 267
rect 599 261 603 262
rect 631 266 635 267
rect 631 261 635 262
rect 711 266 715 267
rect 711 261 715 262
rect 815 266 819 267
rect 815 261 819 262
rect 823 266 827 267
rect 823 261 827 262
rect 943 266 947 267
rect 943 261 947 262
rect 991 266 995 267
rect 991 261 995 262
rect 1063 266 1067 267
rect 1063 261 1067 262
rect 1159 266 1163 267
rect 1159 261 1163 262
rect 1175 266 1179 267
rect 1175 261 1179 262
rect 1287 266 1291 267
rect 1287 261 1291 262
rect 1319 266 1323 267
rect 1319 261 1323 262
rect 1407 266 1411 267
rect 1407 261 1411 262
rect 1471 266 1475 267
rect 1471 261 1475 262
rect 1527 266 1531 267
rect 1527 261 1531 262
rect 1615 266 1619 267
rect 1615 261 1619 262
rect 1647 266 1651 267
rect 1647 261 1651 262
rect 1743 266 1747 267
rect 1743 261 1747 262
rect 1831 266 1835 267
rect 1872 263 1874 286
rect 2022 284 2023 288
rect 2027 284 2028 288
rect 2022 283 2028 284
rect 2110 288 2116 289
rect 2110 284 2111 288
rect 2115 284 2116 288
rect 2110 283 2116 284
rect 2214 288 2220 289
rect 2214 284 2215 288
rect 2219 284 2220 288
rect 2214 283 2220 284
rect 2326 288 2332 289
rect 2326 284 2327 288
rect 2331 284 2332 288
rect 2326 283 2332 284
rect 2438 288 2444 289
rect 2438 284 2439 288
rect 2443 284 2444 288
rect 2438 283 2444 284
rect 2558 288 2564 289
rect 2558 284 2559 288
rect 2563 284 2564 288
rect 2558 283 2564 284
rect 2686 288 2692 289
rect 2686 284 2687 288
rect 2691 284 2692 288
rect 2686 283 2692 284
rect 2830 288 2836 289
rect 2830 284 2831 288
rect 2835 284 2836 288
rect 2830 283 2836 284
rect 2990 288 2996 289
rect 2990 284 2991 288
rect 2995 284 2996 288
rect 2990 283 2996 284
rect 3158 288 3164 289
rect 3158 284 3159 288
rect 3163 284 3164 288
rect 3158 283 3164 284
rect 3334 288 3340 289
rect 3334 284 3335 288
rect 3339 284 3340 288
rect 3334 283 3340 284
rect 3502 288 3508 289
rect 3502 284 3503 288
rect 3507 284 3508 288
rect 3590 287 3591 291
rect 3595 287 3596 291
rect 3590 286 3596 287
rect 3502 283 3508 284
rect 2024 263 2026 283
rect 2112 263 2114 283
rect 2216 263 2218 283
rect 2328 263 2330 283
rect 2440 263 2442 283
rect 2560 263 2562 283
rect 2688 263 2690 283
rect 2832 263 2834 283
rect 2992 263 2994 283
rect 3160 263 3162 283
rect 3336 263 3338 283
rect 3504 263 3506 283
rect 3592 263 3594 286
rect 1831 261 1835 262
rect 1871 262 1875 263
rect 112 242 114 261
rect 304 245 306 261
rect 392 245 394 261
rect 496 245 498 261
rect 600 245 602 261
rect 712 245 714 261
rect 824 245 826 261
rect 944 245 946 261
rect 1064 245 1066 261
rect 1176 245 1178 261
rect 1288 245 1290 261
rect 1408 245 1410 261
rect 1528 245 1530 261
rect 1648 245 1650 261
rect 1744 245 1746 261
rect 302 244 308 245
rect 110 241 116 242
rect 110 237 111 241
rect 115 237 116 241
rect 302 240 303 244
rect 307 240 308 244
rect 302 239 308 240
rect 390 244 396 245
rect 390 240 391 244
rect 395 240 396 244
rect 390 239 396 240
rect 494 244 500 245
rect 494 240 495 244
rect 499 240 500 244
rect 494 239 500 240
rect 598 244 604 245
rect 598 240 599 244
rect 603 240 604 244
rect 598 239 604 240
rect 710 244 716 245
rect 710 240 711 244
rect 715 240 716 244
rect 710 239 716 240
rect 822 244 828 245
rect 822 240 823 244
rect 827 240 828 244
rect 822 239 828 240
rect 942 244 948 245
rect 942 240 943 244
rect 947 240 948 244
rect 942 239 948 240
rect 1062 244 1068 245
rect 1062 240 1063 244
rect 1067 240 1068 244
rect 1062 239 1068 240
rect 1174 244 1180 245
rect 1174 240 1175 244
rect 1179 240 1180 244
rect 1174 239 1180 240
rect 1286 244 1292 245
rect 1286 240 1287 244
rect 1291 240 1292 244
rect 1286 239 1292 240
rect 1406 244 1412 245
rect 1406 240 1407 244
rect 1411 240 1412 244
rect 1406 239 1412 240
rect 1526 244 1532 245
rect 1526 240 1527 244
rect 1531 240 1532 244
rect 1526 239 1532 240
rect 1646 244 1652 245
rect 1646 240 1647 244
rect 1651 240 1652 244
rect 1646 239 1652 240
rect 1742 244 1748 245
rect 1742 240 1743 244
rect 1747 240 1748 244
rect 1832 242 1834 261
rect 1871 257 1875 258
rect 2023 262 2027 263
rect 2023 257 2027 258
rect 2071 262 2075 263
rect 2071 257 2075 258
rect 2111 262 2115 263
rect 2111 257 2115 258
rect 2215 262 2219 263
rect 2215 257 2219 258
rect 2319 262 2323 263
rect 2319 257 2323 258
rect 2327 262 2331 263
rect 2327 257 2331 258
rect 2439 262 2443 263
rect 2439 257 2443 258
rect 2543 262 2547 263
rect 2543 257 2547 258
rect 2559 262 2563 263
rect 2559 257 2563 258
rect 2687 262 2691 263
rect 2687 257 2691 258
rect 2743 262 2747 263
rect 2743 257 2747 258
rect 2831 262 2835 263
rect 2831 257 2835 258
rect 2927 262 2931 263
rect 2927 257 2931 258
rect 2991 262 2995 263
rect 2991 257 2995 258
rect 3087 262 3091 263
rect 3087 257 3091 258
rect 3159 262 3163 263
rect 3159 257 3163 258
rect 3239 262 3243 263
rect 3239 257 3243 258
rect 3335 262 3339 263
rect 3335 257 3339 258
rect 3383 262 3387 263
rect 3383 257 3387 258
rect 3503 262 3507 263
rect 3503 257 3507 258
rect 3591 262 3595 263
rect 3591 257 3595 258
rect 1742 239 1748 240
rect 1830 241 1836 242
rect 110 236 116 237
rect 1830 237 1831 241
rect 1835 237 1836 241
rect 1872 238 1874 257
rect 2072 241 2074 257
rect 2320 241 2322 257
rect 2544 241 2546 257
rect 2744 241 2746 257
rect 2928 241 2930 257
rect 3088 241 3090 257
rect 3240 241 3242 257
rect 3384 241 3386 257
rect 3504 241 3506 257
rect 2070 240 2076 241
rect 1830 236 1836 237
rect 1870 237 1876 238
rect 1870 233 1871 237
rect 1875 233 1876 237
rect 2070 236 2071 240
rect 2075 236 2076 240
rect 2070 235 2076 236
rect 2318 240 2324 241
rect 2318 236 2319 240
rect 2323 236 2324 240
rect 2318 235 2324 236
rect 2542 240 2548 241
rect 2542 236 2543 240
rect 2547 236 2548 240
rect 2542 235 2548 236
rect 2742 240 2748 241
rect 2742 236 2743 240
rect 2747 236 2748 240
rect 2742 235 2748 236
rect 2926 240 2932 241
rect 2926 236 2927 240
rect 2931 236 2932 240
rect 2926 235 2932 236
rect 3086 240 3092 241
rect 3086 236 3087 240
rect 3091 236 3092 240
rect 3086 235 3092 236
rect 3238 240 3244 241
rect 3238 236 3239 240
rect 3243 236 3244 240
rect 3238 235 3244 236
rect 3382 240 3388 241
rect 3382 236 3383 240
rect 3387 236 3388 240
rect 3382 235 3388 236
rect 3502 240 3508 241
rect 3502 236 3503 240
rect 3507 236 3508 240
rect 3592 238 3594 257
rect 3502 235 3508 236
rect 3590 237 3596 238
rect 1870 232 1876 233
rect 3590 233 3591 237
rect 3595 233 3596 237
rect 3590 232 3596 233
rect 110 224 116 225
rect 110 220 111 224
rect 115 220 116 224
rect 110 219 116 220
rect 1830 224 1836 225
rect 1830 220 1831 224
rect 1835 220 1836 224
rect 1830 219 1836 220
rect 1870 220 1876 221
rect 112 167 114 219
rect 310 206 316 207
rect 310 202 311 206
rect 315 202 316 206
rect 310 201 316 202
rect 398 206 404 207
rect 398 202 399 206
rect 403 202 404 206
rect 398 201 404 202
rect 502 206 508 207
rect 502 202 503 206
rect 507 202 508 206
rect 502 201 508 202
rect 606 206 612 207
rect 606 202 607 206
rect 611 202 612 206
rect 606 201 612 202
rect 718 206 724 207
rect 718 202 719 206
rect 723 202 724 206
rect 718 201 724 202
rect 830 206 836 207
rect 830 202 831 206
rect 835 202 836 206
rect 830 201 836 202
rect 950 206 956 207
rect 950 202 951 206
rect 955 202 956 206
rect 950 201 956 202
rect 1070 206 1076 207
rect 1070 202 1071 206
rect 1075 202 1076 206
rect 1070 201 1076 202
rect 1182 206 1188 207
rect 1182 202 1183 206
rect 1187 202 1188 206
rect 1182 201 1188 202
rect 1294 206 1300 207
rect 1294 202 1295 206
rect 1299 202 1300 206
rect 1294 201 1300 202
rect 1414 206 1420 207
rect 1414 202 1415 206
rect 1419 202 1420 206
rect 1414 201 1420 202
rect 1534 206 1540 207
rect 1534 202 1535 206
rect 1539 202 1540 206
rect 1534 201 1540 202
rect 1654 206 1660 207
rect 1654 202 1655 206
rect 1659 202 1660 206
rect 1654 201 1660 202
rect 1750 206 1756 207
rect 1750 202 1751 206
rect 1755 202 1756 206
rect 1750 201 1756 202
rect 312 167 314 201
rect 400 167 402 201
rect 504 167 506 201
rect 608 167 610 201
rect 720 167 722 201
rect 832 167 834 201
rect 952 167 954 201
rect 1072 167 1074 201
rect 1184 167 1186 201
rect 1296 167 1298 201
rect 1416 167 1418 201
rect 1536 167 1538 201
rect 1656 167 1658 201
rect 1752 167 1754 201
rect 1832 167 1834 219
rect 1870 216 1871 220
rect 1875 216 1876 220
rect 1870 215 1876 216
rect 3590 220 3596 221
rect 3590 216 3591 220
rect 3595 216 3596 220
rect 3590 215 3596 216
rect 111 166 115 167
rect 111 161 115 162
rect 263 166 267 167
rect 263 161 267 162
rect 311 166 315 167
rect 311 161 315 162
rect 343 166 347 167
rect 343 161 347 162
rect 399 166 403 167
rect 399 161 403 162
rect 423 166 427 167
rect 423 161 427 162
rect 503 166 507 167
rect 503 161 507 162
rect 583 166 587 167
rect 583 161 587 162
rect 607 166 611 167
rect 607 161 611 162
rect 663 166 667 167
rect 663 161 667 162
rect 719 166 723 167
rect 719 161 723 162
rect 743 166 747 167
rect 743 161 747 162
rect 823 166 827 167
rect 823 161 827 162
rect 831 166 835 167
rect 831 161 835 162
rect 903 166 907 167
rect 903 161 907 162
rect 951 166 955 167
rect 951 161 955 162
rect 983 166 987 167
rect 983 161 987 162
rect 1063 166 1067 167
rect 1063 161 1067 162
rect 1071 166 1075 167
rect 1071 161 1075 162
rect 1143 166 1147 167
rect 1143 161 1147 162
rect 1183 166 1187 167
rect 1183 161 1187 162
rect 1223 166 1227 167
rect 1223 161 1227 162
rect 1295 166 1299 167
rect 1295 161 1299 162
rect 1303 166 1307 167
rect 1303 161 1307 162
rect 1383 166 1387 167
rect 1383 161 1387 162
rect 1415 166 1419 167
rect 1415 161 1419 162
rect 1463 166 1467 167
rect 1463 161 1467 162
rect 1535 166 1539 167
rect 1535 161 1539 162
rect 1543 166 1547 167
rect 1543 161 1547 162
rect 1655 166 1659 167
rect 1655 161 1659 162
rect 1751 166 1755 167
rect 1751 161 1755 162
rect 1831 166 1835 167
rect 1872 163 1874 215
rect 2078 202 2084 203
rect 2078 198 2079 202
rect 2083 198 2084 202
rect 2078 197 2084 198
rect 2326 202 2332 203
rect 2326 198 2327 202
rect 2331 198 2332 202
rect 2326 197 2332 198
rect 2550 202 2556 203
rect 2550 198 2551 202
rect 2555 198 2556 202
rect 2550 197 2556 198
rect 2750 202 2756 203
rect 2750 198 2751 202
rect 2755 198 2756 202
rect 2750 197 2756 198
rect 2934 202 2940 203
rect 2934 198 2935 202
rect 2939 198 2940 202
rect 2934 197 2940 198
rect 3094 202 3100 203
rect 3094 198 3095 202
rect 3099 198 3100 202
rect 3094 197 3100 198
rect 3246 202 3252 203
rect 3246 198 3247 202
rect 3251 198 3252 202
rect 3246 197 3252 198
rect 3390 202 3396 203
rect 3390 198 3391 202
rect 3395 198 3396 202
rect 3390 197 3396 198
rect 3510 202 3516 203
rect 3510 198 3511 202
rect 3515 198 3516 202
rect 3510 197 3516 198
rect 2080 163 2082 197
rect 2328 163 2330 197
rect 2552 163 2554 197
rect 2752 163 2754 197
rect 2936 163 2938 197
rect 3096 163 3098 197
rect 3248 163 3250 197
rect 3392 163 3394 197
rect 3512 163 3514 197
rect 3592 163 3594 215
rect 1831 161 1835 162
rect 1871 162 1875 163
rect 112 133 114 161
rect 264 151 266 161
rect 344 151 346 161
rect 424 151 426 161
rect 504 151 506 161
rect 584 151 586 161
rect 664 151 666 161
rect 744 151 746 161
rect 824 151 826 161
rect 904 151 906 161
rect 984 151 986 161
rect 1064 151 1066 161
rect 1144 151 1146 161
rect 1224 151 1226 161
rect 1304 151 1306 161
rect 1384 151 1386 161
rect 1464 151 1466 161
rect 1544 151 1546 161
rect 262 150 268 151
rect 262 146 263 150
rect 267 146 268 150
rect 262 145 268 146
rect 342 150 348 151
rect 342 146 343 150
rect 347 146 348 150
rect 342 145 348 146
rect 422 150 428 151
rect 422 146 423 150
rect 427 146 428 150
rect 422 145 428 146
rect 502 150 508 151
rect 502 146 503 150
rect 507 146 508 150
rect 502 145 508 146
rect 582 150 588 151
rect 582 146 583 150
rect 587 146 588 150
rect 582 145 588 146
rect 662 150 668 151
rect 662 146 663 150
rect 667 146 668 150
rect 662 145 668 146
rect 742 150 748 151
rect 742 146 743 150
rect 747 146 748 150
rect 742 145 748 146
rect 822 150 828 151
rect 822 146 823 150
rect 827 146 828 150
rect 822 145 828 146
rect 902 150 908 151
rect 902 146 903 150
rect 907 146 908 150
rect 902 145 908 146
rect 982 150 988 151
rect 982 146 983 150
rect 987 146 988 150
rect 982 145 988 146
rect 1062 150 1068 151
rect 1062 146 1063 150
rect 1067 146 1068 150
rect 1062 145 1068 146
rect 1142 150 1148 151
rect 1142 146 1143 150
rect 1147 146 1148 150
rect 1142 145 1148 146
rect 1222 150 1228 151
rect 1222 146 1223 150
rect 1227 146 1228 150
rect 1222 145 1228 146
rect 1302 150 1308 151
rect 1302 146 1303 150
rect 1307 146 1308 150
rect 1302 145 1308 146
rect 1382 150 1388 151
rect 1382 146 1383 150
rect 1387 146 1388 150
rect 1382 145 1388 146
rect 1462 150 1468 151
rect 1462 146 1463 150
rect 1467 146 1468 150
rect 1462 145 1468 146
rect 1542 150 1548 151
rect 1542 146 1543 150
rect 1547 146 1548 150
rect 1542 145 1548 146
rect 1832 133 1834 161
rect 1871 157 1875 158
rect 1903 162 1907 163
rect 1903 157 1907 158
rect 1983 162 1987 163
rect 1983 157 1987 158
rect 2063 162 2067 163
rect 2063 157 2067 158
rect 2079 162 2083 163
rect 2079 157 2083 158
rect 2143 162 2147 163
rect 2143 157 2147 158
rect 2223 162 2227 163
rect 2223 157 2227 158
rect 2303 162 2307 163
rect 2303 157 2307 158
rect 2327 162 2331 163
rect 2327 157 2331 158
rect 2399 162 2403 163
rect 2399 157 2403 158
rect 2503 162 2507 163
rect 2503 157 2507 158
rect 2551 162 2555 163
rect 2551 157 2555 158
rect 2607 162 2611 163
rect 2607 157 2611 158
rect 2711 162 2715 163
rect 2711 157 2715 158
rect 2751 162 2755 163
rect 2751 157 2755 158
rect 2815 162 2819 163
rect 2815 157 2819 158
rect 2911 162 2915 163
rect 2911 157 2915 158
rect 2935 162 2939 163
rect 2935 157 2939 158
rect 2999 162 3003 163
rect 2999 157 3003 158
rect 3087 162 3091 163
rect 3087 157 3091 158
rect 3095 162 3099 163
rect 3095 157 3099 158
rect 3175 162 3179 163
rect 3175 157 3179 158
rect 3247 162 3251 163
rect 3247 157 3251 158
rect 3263 162 3267 163
rect 3263 157 3267 158
rect 3351 162 3355 163
rect 3351 157 3355 158
rect 3391 162 3395 163
rect 3391 157 3395 158
rect 3431 162 3435 163
rect 3431 157 3435 158
rect 3511 162 3515 163
rect 3511 157 3515 158
rect 3591 162 3595 163
rect 3591 157 3595 158
rect 110 132 116 133
rect 110 128 111 132
rect 115 128 116 132
rect 110 127 116 128
rect 1830 132 1836 133
rect 1830 128 1831 132
rect 1835 128 1836 132
rect 1872 129 1874 157
rect 1904 147 1906 157
rect 1984 147 1986 157
rect 2064 147 2066 157
rect 2144 147 2146 157
rect 2224 147 2226 157
rect 2304 147 2306 157
rect 2400 147 2402 157
rect 2504 147 2506 157
rect 2608 147 2610 157
rect 2712 147 2714 157
rect 2816 147 2818 157
rect 2912 147 2914 157
rect 3000 147 3002 157
rect 3088 147 3090 157
rect 3176 147 3178 157
rect 3264 147 3266 157
rect 3352 147 3354 157
rect 3432 147 3434 157
rect 3512 147 3514 157
rect 1902 146 1908 147
rect 1902 142 1903 146
rect 1907 142 1908 146
rect 1902 141 1908 142
rect 1982 146 1988 147
rect 1982 142 1983 146
rect 1987 142 1988 146
rect 1982 141 1988 142
rect 2062 146 2068 147
rect 2062 142 2063 146
rect 2067 142 2068 146
rect 2062 141 2068 142
rect 2142 146 2148 147
rect 2142 142 2143 146
rect 2147 142 2148 146
rect 2142 141 2148 142
rect 2222 146 2228 147
rect 2222 142 2223 146
rect 2227 142 2228 146
rect 2222 141 2228 142
rect 2302 146 2308 147
rect 2302 142 2303 146
rect 2307 142 2308 146
rect 2302 141 2308 142
rect 2398 146 2404 147
rect 2398 142 2399 146
rect 2403 142 2404 146
rect 2398 141 2404 142
rect 2502 146 2508 147
rect 2502 142 2503 146
rect 2507 142 2508 146
rect 2502 141 2508 142
rect 2606 146 2612 147
rect 2606 142 2607 146
rect 2611 142 2612 146
rect 2606 141 2612 142
rect 2710 146 2716 147
rect 2710 142 2711 146
rect 2715 142 2716 146
rect 2710 141 2716 142
rect 2814 146 2820 147
rect 2814 142 2815 146
rect 2819 142 2820 146
rect 2814 141 2820 142
rect 2910 146 2916 147
rect 2910 142 2911 146
rect 2915 142 2916 146
rect 2910 141 2916 142
rect 2998 146 3004 147
rect 2998 142 2999 146
rect 3003 142 3004 146
rect 2998 141 3004 142
rect 3086 146 3092 147
rect 3086 142 3087 146
rect 3091 142 3092 146
rect 3086 141 3092 142
rect 3174 146 3180 147
rect 3174 142 3175 146
rect 3179 142 3180 146
rect 3174 141 3180 142
rect 3262 146 3268 147
rect 3262 142 3263 146
rect 3267 142 3268 146
rect 3262 141 3268 142
rect 3350 146 3356 147
rect 3350 142 3351 146
rect 3355 142 3356 146
rect 3350 141 3356 142
rect 3430 146 3436 147
rect 3430 142 3431 146
rect 3435 142 3436 146
rect 3430 141 3436 142
rect 3510 146 3516 147
rect 3510 142 3511 146
rect 3515 142 3516 146
rect 3510 141 3516 142
rect 3592 129 3594 157
rect 1830 127 1836 128
rect 1870 128 1876 129
rect 1870 124 1871 128
rect 1875 124 1876 128
rect 1870 123 1876 124
rect 3590 128 3596 129
rect 3590 124 3591 128
rect 3595 124 3596 128
rect 3590 123 3596 124
rect 110 115 116 116
rect 110 111 111 115
rect 115 111 116 115
rect 1830 115 1836 116
rect 110 110 116 111
rect 254 112 260 113
rect 112 91 114 110
rect 254 108 255 112
rect 259 108 260 112
rect 254 107 260 108
rect 334 112 340 113
rect 334 108 335 112
rect 339 108 340 112
rect 334 107 340 108
rect 414 112 420 113
rect 414 108 415 112
rect 419 108 420 112
rect 414 107 420 108
rect 494 112 500 113
rect 494 108 495 112
rect 499 108 500 112
rect 494 107 500 108
rect 574 112 580 113
rect 574 108 575 112
rect 579 108 580 112
rect 574 107 580 108
rect 654 112 660 113
rect 654 108 655 112
rect 659 108 660 112
rect 654 107 660 108
rect 734 112 740 113
rect 734 108 735 112
rect 739 108 740 112
rect 734 107 740 108
rect 814 112 820 113
rect 814 108 815 112
rect 819 108 820 112
rect 814 107 820 108
rect 894 112 900 113
rect 894 108 895 112
rect 899 108 900 112
rect 894 107 900 108
rect 974 112 980 113
rect 974 108 975 112
rect 979 108 980 112
rect 974 107 980 108
rect 1054 112 1060 113
rect 1054 108 1055 112
rect 1059 108 1060 112
rect 1054 107 1060 108
rect 1134 112 1140 113
rect 1134 108 1135 112
rect 1139 108 1140 112
rect 1134 107 1140 108
rect 1214 112 1220 113
rect 1214 108 1215 112
rect 1219 108 1220 112
rect 1214 107 1220 108
rect 1294 112 1300 113
rect 1294 108 1295 112
rect 1299 108 1300 112
rect 1294 107 1300 108
rect 1374 112 1380 113
rect 1374 108 1375 112
rect 1379 108 1380 112
rect 1374 107 1380 108
rect 1454 112 1460 113
rect 1454 108 1455 112
rect 1459 108 1460 112
rect 1454 107 1460 108
rect 1534 112 1540 113
rect 1534 108 1535 112
rect 1539 108 1540 112
rect 1830 111 1831 115
rect 1835 111 1836 115
rect 1830 110 1836 111
rect 1870 111 1876 112
rect 1534 107 1540 108
rect 256 91 258 107
rect 336 91 338 107
rect 416 91 418 107
rect 496 91 498 107
rect 576 91 578 107
rect 656 91 658 107
rect 736 91 738 107
rect 816 91 818 107
rect 896 91 898 107
rect 976 91 978 107
rect 1056 91 1058 107
rect 1136 91 1138 107
rect 1216 91 1218 107
rect 1296 91 1298 107
rect 1376 91 1378 107
rect 1456 91 1458 107
rect 1536 91 1538 107
rect 1832 91 1834 110
rect 1870 107 1871 111
rect 1875 107 1876 111
rect 3590 111 3596 112
rect 1870 106 1876 107
rect 1894 108 1900 109
rect 111 90 115 91
rect 111 85 115 86
rect 255 90 259 91
rect 255 85 259 86
rect 335 90 339 91
rect 335 85 339 86
rect 415 90 419 91
rect 415 85 419 86
rect 495 90 499 91
rect 495 85 499 86
rect 575 90 579 91
rect 575 85 579 86
rect 655 90 659 91
rect 655 85 659 86
rect 735 90 739 91
rect 735 85 739 86
rect 815 90 819 91
rect 815 85 819 86
rect 895 90 899 91
rect 895 85 899 86
rect 975 90 979 91
rect 975 85 979 86
rect 1055 90 1059 91
rect 1055 85 1059 86
rect 1135 90 1139 91
rect 1135 85 1139 86
rect 1215 90 1219 91
rect 1215 85 1219 86
rect 1295 90 1299 91
rect 1295 85 1299 86
rect 1375 90 1379 91
rect 1375 85 1379 86
rect 1455 90 1459 91
rect 1455 85 1459 86
rect 1535 90 1539 91
rect 1535 85 1539 86
rect 1831 90 1835 91
rect 1872 87 1874 106
rect 1894 104 1895 108
rect 1899 104 1900 108
rect 1894 103 1900 104
rect 1974 108 1980 109
rect 1974 104 1975 108
rect 1979 104 1980 108
rect 1974 103 1980 104
rect 2054 108 2060 109
rect 2054 104 2055 108
rect 2059 104 2060 108
rect 2054 103 2060 104
rect 2134 108 2140 109
rect 2134 104 2135 108
rect 2139 104 2140 108
rect 2134 103 2140 104
rect 2214 108 2220 109
rect 2214 104 2215 108
rect 2219 104 2220 108
rect 2214 103 2220 104
rect 2294 108 2300 109
rect 2294 104 2295 108
rect 2299 104 2300 108
rect 2294 103 2300 104
rect 2390 108 2396 109
rect 2390 104 2391 108
rect 2395 104 2396 108
rect 2390 103 2396 104
rect 2494 108 2500 109
rect 2494 104 2495 108
rect 2499 104 2500 108
rect 2494 103 2500 104
rect 2598 108 2604 109
rect 2598 104 2599 108
rect 2603 104 2604 108
rect 2598 103 2604 104
rect 2702 108 2708 109
rect 2702 104 2703 108
rect 2707 104 2708 108
rect 2702 103 2708 104
rect 2806 108 2812 109
rect 2806 104 2807 108
rect 2811 104 2812 108
rect 2806 103 2812 104
rect 2902 108 2908 109
rect 2902 104 2903 108
rect 2907 104 2908 108
rect 2902 103 2908 104
rect 2990 108 2996 109
rect 2990 104 2991 108
rect 2995 104 2996 108
rect 2990 103 2996 104
rect 3078 108 3084 109
rect 3078 104 3079 108
rect 3083 104 3084 108
rect 3078 103 3084 104
rect 3166 108 3172 109
rect 3166 104 3167 108
rect 3171 104 3172 108
rect 3166 103 3172 104
rect 3254 108 3260 109
rect 3254 104 3255 108
rect 3259 104 3260 108
rect 3254 103 3260 104
rect 3342 108 3348 109
rect 3342 104 3343 108
rect 3347 104 3348 108
rect 3342 103 3348 104
rect 3422 108 3428 109
rect 3422 104 3423 108
rect 3427 104 3428 108
rect 3422 103 3428 104
rect 3502 108 3508 109
rect 3502 104 3503 108
rect 3507 104 3508 108
rect 3590 107 3591 111
rect 3595 107 3596 111
rect 3590 106 3596 107
rect 3502 103 3508 104
rect 1896 87 1898 103
rect 1976 87 1978 103
rect 2056 87 2058 103
rect 2136 87 2138 103
rect 2216 87 2218 103
rect 2296 87 2298 103
rect 2392 87 2394 103
rect 2496 87 2498 103
rect 2600 87 2602 103
rect 2704 87 2706 103
rect 2808 87 2810 103
rect 2904 87 2906 103
rect 2992 87 2994 103
rect 3080 87 3082 103
rect 3168 87 3170 103
rect 3256 87 3258 103
rect 3344 87 3346 103
rect 3424 87 3426 103
rect 3504 87 3506 103
rect 3592 87 3594 106
rect 1831 85 1835 86
rect 1871 86 1875 87
rect 1871 81 1875 82
rect 1895 86 1899 87
rect 1895 81 1899 82
rect 1975 86 1979 87
rect 1975 81 1979 82
rect 2055 86 2059 87
rect 2055 81 2059 82
rect 2135 86 2139 87
rect 2135 81 2139 82
rect 2215 86 2219 87
rect 2215 81 2219 82
rect 2295 86 2299 87
rect 2295 81 2299 82
rect 2391 86 2395 87
rect 2391 81 2395 82
rect 2495 86 2499 87
rect 2495 81 2499 82
rect 2599 86 2603 87
rect 2599 81 2603 82
rect 2703 86 2707 87
rect 2703 81 2707 82
rect 2807 86 2811 87
rect 2807 81 2811 82
rect 2903 86 2907 87
rect 2903 81 2907 82
rect 2991 86 2995 87
rect 2991 81 2995 82
rect 3079 86 3083 87
rect 3079 81 3083 82
rect 3167 86 3171 87
rect 3167 81 3171 82
rect 3255 86 3259 87
rect 3255 81 3259 82
rect 3343 86 3347 87
rect 3343 81 3347 82
rect 3423 86 3427 87
rect 3423 81 3427 82
rect 3503 86 3507 87
rect 3503 81 3507 82
rect 3591 86 3595 87
rect 3591 81 3595 82
<< m4c >>
rect 111 3654 115 3658
rect 143 3654 147 3658
rect 223 3654 227 3658
rect 351 3654 355 3658
rect 495 3654 499 3658
rect 647 3654 651 3658
rect 807 3654 811 3658
rect 975 3654 979 3658
rect 1151 3654 1155 3658
rect 1335 3654 1339 3658
rect 1831 3654 1835 3658
rect 1871 3626 1875 3630
rect 1927 3626 1931 3630
rect 2007 3626 2011 3630
rect 2103 3626 2107 3630
rect 2207 3626 2211 3630
rect 2319 3626 2323 3630
rect 2431 3626 2435 3630
rect 2551 3626 2555 3630
rect 2663 3626 2667 3630
rect 2775 3626 2779 3630
rect 2879 3626 2883 3630
rect 2983 3626 2987 3630
rect 3095 3626 3099 3630
rect 3207 3626 3211 3630
rect 3591 3626 3595 3630
rect 111 3578 115 3582
rect 135 3578 139 3582
rect 215 3578 219 3582
rect 239 3578 243 3582
rect 343 3578 347 3582
rect 359 3578 363 3582
rect 479 3578 483 3582
rect 487 3578 491 3582
rect 607 3578 611 3582
rect 639 3578 643 3582
rect 735 3578 739 3582
rect 799 3578 803 3582
rect 863 3578 867 3582
rect 967 3578 971 3582
rect 983 3578 987 3582
rect 1095 3578 1099 3582
rect 1143 3578 1147 3582
rect 1207 3578 1211 3582
rect 1319 3578 1323 3582
rect 1327 3578 1331 3582
rect 1439 3578 1443 3582
rect 1831 3578 1835 3582
rect 1871 3550 1875 3554
rect 1919 3550 1923 3554
rect 1943 3550 1947 3554
rect 1999 3550 2003 3554
rect 2095 3550 2099 3554
rect 2127 3550 2131 3554
rect 2199 3550 2203 3554
rect 2303 3550 2307 3554
rect 2311 3550 2315 3554
rect 2423 3550 2427 3554
rect 2479 3550 2483 3554
rect 2543 3550 2547 3554
rect 2647 3550 2651 3554
rect 2655 3550 2659 3554
rect 2767 3550 2771 3554
rect 2815 3550 2819 3554
rect 2871 3550 2875 3554
rect 2975 3550 2979 3554
rect 3087 3550 3091 3554
rect 3135 3550 3139 3554
rect 3199 3550 3203 3554
rect 3303 3550 3307 3554
rect 3591 3550 3595 3554
rect 111 3502 115 3506
rect 167 3502 171 3506
rect 247 3502 251 3506
rect 287 3502 291 3506
rect 367 3502 371 3506
rect 415 3502 419 3506
rect 487 3502 491 3506
rect 551 3502 555 3506
rect 615 3502 619 3506
rect 687 3502 691 3506
rect 743 3502 747 3506
rect 823 3502 827 3506
rect 871 3502 875 3506
rect 951 3502 955 3506
rect 991 3502 995 3506
rect 1071 3502 1075 3506
rect 1103 3502 1107 3506
rect 1183 3502 1187 3506
rect 1215 3502 1219 3506
rect 1303 3502 1307 3506
rect 1327 3502 1331 3506
rect 1423 3502 1427 3506
rect 1447 3502 1451 3506
rect 1831 3502 1835 3506
rect 1871 3474 1875 3478
rect 1951 3474 1955 3478
rect 1959 3474 1963 3478
rect 2079 3474 2083 3478
rect 2135 3474 2139 3478
rect 2199 3474 2203 3478
rect 2311 3474 2315 3478
rect 2335 3474 2339 3478
rect 2479 3474 2483 3478
rect 2487 3474 2491 3478
rect 2631 3474 2635 3478
rect 2655 3474 2659 3478
rect 2791 3474 2795 3478
rect 2823 3474 2827 3478
rect 2959 3474 2963 3478
rect 2983 3474 2987 3478
rect 3127 3474 3131 3478
rect 3143 3474 3147 3478
rect 3303 3474 3307 3478
rect 3311 3474 3315 3478
rect 3591 3474 3595 3478
rect 111 3418 115 3422
rect 135 3418 139 3422
rect 159 3418 163 3422
rect 247 3418 251 3422
rect 279 3418 283 3422
rect 375 3418 379 3422
rect 407 3418 411 3422
rect 503 3418 507 3422
rect 543 3418 547 3422
rect 639 3418 643 3422
rect 679 3418 683 3422
rect 775 3418 779 3422
rect 815 3418 819 3422
rect 903 3418 907 3422
rect 943 3418 947 3422
rect 1031 3418 1035 3422
rect 1063 3418 1067 3422
rect 1159 3418 1163 3422
rect 1175 3418 1179 3422
rect 1287 3418 1291 3422
rect 1295 3418 1299 3422
rect 1415 3418 1419 3422
rect 1831 3418 1835 3422
rect 1871 3390 1875 3394
rect 1951 3390 1955 3394
rect 1975 3390 1979 3394
rect 2071 3390 2075 3394
rect 2135 3390 2139 3394
rect 2191 3390 2195 3394
rect 2287 3390 2291 3394
rect 2327 3390 2331 3394
rect 2431 3390 2435 3394
rect 2471 3390 2475 3394
rect 2559 3390 2563 3394
rect 2623 3390 2627 3394
rect 2679 3390 2683 3394
rect 2783 3390 2787 3394
rect 2791 3390 2795 3394
rect 2895 3390 2899 3394
rect 2951 3390 2955 3394
rect 2991 3390 2995 3394
rect 3079 3390 3083 3394
rect 3119 3390 3123 3394
rect 3167 3390 3171 3394
rect 3255 3390 3259 3394
rect 3295 3390 3299 3394
rect 3343 3390 3347 3394
rect 3423 3390 3427 3394
rect 3503 3390 3507 3394
rect 3591 3390 3595 3394
rect 111 3338 115 3342
rect 143 3338 147 3342
rect 255 3338 259 3342
rect 271 3338 275 3342
rect 383 3338 387 3342
rect 391 3338 395 3342
rect 511 3338 515 3342
rect 519 3338 523 3342
rect 647 3338 651 3342
rect 655 3338 659 3342
rect 783 3338 787 3342
rect 791 3338 795 3342
rect 911 3338 915 3342
rect 919 3338 923 3342
rect 1039 3338 1043 3342
rect 1055 3338 1059 3342
rect 1167 3338 1171 3342
rect 1191 3338 1195 3342
rect 1295 3338 1299 3342
rect 1327 3338 1331 3342
rect 1423 3338 1427 3342
rect 1463 3338 1467 3342
rect 1831 3338 1835 3342
rect 1871 3310 1875 3314
rect 1935 3310 1939 3314
rect 1983 3310 1987 3314
rect 2071 3310 2075 3314
rect 2143 3310 2147 3314
rect 2207 3310 2211 3314
rect 2295 3310 2299 3314
rect 2367 3310 2371 3314
rect 2439 3310 2443 3314
rect 2551 3310 2555 3314
rect 2567 3310 2571 3314
rect 2687 3310 2691 3314
rect 2767 3310 2771 3314
rect 2799 3310 2803 3314
rect 2903 3310 2907 3314
rect 2999 3310 3003 3314
rect 3007 3310 3011 3314
rect 3087 3310 3091 3314
rect 3175 3310 3179 3314
rect 3255 3310 3259 3314
rect 3263 3310 3267 3314
rect 3351 3310 3355 3314
rect 3431 3310 3435 3314
rect 3511 3310 3515 3314
rect 3591 3310 3595 3314
rect 111 3258 115 3262
rect 263 3258 267 3262
rect 383 3258 387 3262
rect 471 3258 475 3262
rect 511 3258 515 3262
rect 575 3258 579 3262
rect 647 3258 651 3262
rect 687 3258 691 3262
rect 783 3258 787 3262
rect 807 3258 811 3262
rect 911 3258 915 3262
rect 935 3258 939 3262
rect 1047 3258 1051 3262
rect 1063 3258 1067 3262
rect 1183 3258 1187 3262
rect 1191 3258 1195 3262
rect 1319 3258 1323 3262
rect 1447 3258 1451 3262
rect 1455 3258 1459 3262
rect 1575 3258 1579 3262
rect 1831 3258 1835 3262
rect 1871 3230 1875 3234
rect 1895 3230 1899 3234
rect 1927 3230 1931 3234
rect 2007 3230 2011 3234
rect 2063 3230 2067 3234
rect 2143 3230 2147 3234
rect 2199 3230 2203 3234
rect 2279 3230 2283 3234
rect 2359 3230 2363 3234
rect 2415 3230 2419 3234
rect 2543 3230 2547 3234
rect 2567 3230 2571 3234
rect 2727 3230 2731 3234
rect 2759 3230 2763 3234
rect 2911 3230 2915 3234
rect 2999 3230 3003 3234
rect 3103 3230 3107 3234
rect 3247 3230 3251 3234
rect 3311 3230 3315 3234
rect 3503 3230 3507 3234
rect 3591 3230 3595 3234
rect 111 3174 115 3178
rect 383 3174 387 3178
rect 391 3174 395 3178
rect 463 3174 467 3178
rect 479 3174 483 3178
rect 543 3174 547 3178
rect 583 3174 587 3178
rect 623 3174 627 3178
rect 695 3174 699 3178
rect 711 3174 715 3178
rect 815 3174 819 3178
rect 927 3174 931 3178
rect 943 3174 947 3178
rect 1039 3174 1043 3178
rect 1071 3174 1075 3178
rect 1159 3174 1163 3178
rect 1199 3174 1203 3178
rect 1271 3174 1275 3178
rect 1327 3174 1331 3178
rect 1383 3174 1387 3178
rect 1455 3174 1459 3178
rect 1495 3174 1499 3178
rect 1583 3174 1587 3178
rect 1615 3174 1619 3178
rect 1735 3174 1739 3178
rect 1831 3174 1835 3178
rect 1871 3154 1875 3158
rect 1903 3154 1907 3158
rect 2015 3154 2019 3158
rect 2079 3154 2083 3158
rect 2151 3154 2155 3158
rect 2271 3154 2275 3158
rect 2287 3154 2291 3158
rect 2423 3154 2427 3158
rect 2455 3154 2459 3158
rect 2575 3154 2579 3158
rect 2623 3154 2627 3158
rect 2735 3154 2739 3158
rect 2783 3154 2787 3158
rect 2919 3154 2923 3158
rect 2935 3154 2939 3158
rect 3079 3154 3083 3158
rect 3111 3154 3115 3158
rect 3231 3154 3235 3158
rect 3319 3154 3323 3158
rect 3511 3154 3515 3158
rect 3591 3154 3595 3158
rect 111 3098 115 3102
rect 375 3098 379 3102
rect 455 3098 459 3102
rect 535 3098 539 3102
rect 615 3098 619 3102
rect 703 3098 707 3102
rect 807 3098 811 3102
rect 919 3098 923 3102
rect 943 3098 947 3102
rect 1023 3098 1027 3102
rect 1031 3098 1035 3102
rect 1103 3098 1107 3102
rect 1151 3098 1155 3102
rect 1183 3098 1187 3102
rect 1263 3098 1267 3102
rect 1343 3098 1347 3102
rect 1375 3098 1379 3102
rect 1423 3098 1427 3102
rect 1487 3098 1491 3102
rect 1503 3098 1507 3102
rect 1583 3098 1587 3102
rect 1607 3098 1611 3102
rect 1663 3098 1667 3102
rect 1727 3098 1731 3102
rect 1743 3098 1747 3102
rect 1831 3098 1835 3102
rect 1871 3070 1875 3074
rect 1895 3070 1899 3074
rect 1991 3070 1995 3074
rect 2071 3070 2075 3074
rect 2247 3070 2251 3074
rect 2263 3070 2267 3074
rect 2447 3070 2451 3074
rect 2487 3070 2491 3074
rect 2615 3070 2619 3074
rect 2703 3070 2707 3074
rect 2775 3070 2779 3074
rect 2895 3070 2899 3074
rect 2927 3070 2931 3074
rect 3063 3070 3067 3074
rect 3071 3070 3075 3074
rect 3223 3070 3227 3074
rect 3375 3070 3379 3074
rect 3503 3070 3507 3074
rect 3591 3070 3595 3074
rect 111 3006 115 3010
rect 207 3006 211 3010
rect 327 3006 331 3010
rect 471 3006 475 3010
rect 631 3006 635 3010
rect 807 3006 811 3010
rect 951 3006 955 3010
rect 983 3006 987 3010
rect 1031 3006 1035 3010
rect 1111 3006 1115 3010
rect 1151 3006 1155 3010
rect 1191 3006 1195 3010
rect 1271 3006 1275 3010
rect 1311 3006 1315 3010
rect 1351 3006 1355 3010
rect 1431 3006 1435 3010
rect 1463 3006 1467 3010
rect 1511 3006 1515 3010
rect 1591 3006 1595 3010
rect 1615 3006 1619 3010
rect 1671 3006 1675 3010
rect 1751 3006 1755 3010
rect 1831 3006 1835 3010
rect 1871 2990 1875 2994
rect 1903 2990 1907 2994
rect 1999 2990 2003 2994
rect 2143 2990 2147 2994
rect 2255 2990 2259 2994
rect 2391 2990 2395 2994
rect 2495 2990 2499 2994
rect 2607 2990 2611 2994
rect 2711 2990 2715 2994
rect 2799 2990 2803 2994
rect 2903 2990 2907 2994
rect 2967 2990 2971 2994
rect 3071 2990 3075 2994
rect 3119 2990 3123 2994
rect 3231 2990 3235 2994
rect 3263 2990 3267 2994
rect 3383 2990 3387 2994
rect 3399 2990 3403 2994
rect 3511 2990 3515 2994
rect 3591 2990 3595 2994
rect 111 2930 115 2934
rect 199 2930 203 2934
rect 247 2930 251 2934
rect 319 2930 323 2934
rect 351 2930 355 2934
rect 463 2930 467 2934
rect 471 2930 475 2934
rect 607 2930 611 2934
rect 623 2930 627 2934
rect 751 2930 755 2934
rect 799 2930 803 2934
rect 895 2930 899 2934
rect 975 2930 979 2934
rect 1031 2930 1035 2934
rect 1143 2930 1147 2934
rect 1159 2930 1163 2934
rect 1279 2930 1283 2934
rect 1303 2930 1307 2934
rect 1399 2930 1403 2934
rect 1455 2930 1459 2934
rect 1519 2930 1523 2934
rect 1607 2930 1611 2934
rect 1639 2930 1643 2934
rect 1743 2930 1747 2934
rect 1831 2930 1835 2934
rect 1871 2902 1875 2906
rect 1895 2902 1899 2906
rect 2135 2902 2139 2906
rect 2351 2902 2355 2906
rect 2383 2902 2387 2906
rect 2447 2902 2451 2906
rect 2551 2902 2555 2906
rect 2599 2902 2603 2906
rect 2655 2902 2659 2906
rect 2759 2902 2763 2906
rect 2791 2902 2795 2906
rect 2871 2902 2875 2906
rect 2959 2902 2963 2906
rect 2983 2902 2987 2906
rect 3095 2902 3099 2906
rect 3111 2902 3115 2906
rect 3207 2902 3211 2906
rect 3255 2902 3259 2906
rect 3391 2902 3395 2906
rect 3503 2902 3507 2906
rect 3591 2902 3595 2906
rect 111 2854 115 2858
rect 151 2854 155 2858
rect 255 2854 259 2858
rect 279 2854 283 2858
rect 359 2854 363 2858
rect 407 2854 411 2858
rect 479 2854 483 2858
rect 543 2854 547 2858
rect 615 2854 619 2858
rect 671 2854 675 2858
rect 759 2854 763 2858
rect 799 2854 803 2858
rect 903 2854 907 2858
rect 919 2854 923 2858
rect 1039 2854 1043 2858
rect 1151 2854 1155 2858
rect 1167 2854 1171 2858
rect 1271 2854 1275 2858
rect 1287 2854 1291 2858
rect 1391 2854 1395 2858
rect 1407 2854 1411 2858
rect 1527 2854 1531 2858
rect 1647 2854 1651 2858
rect 1831 2854 1835 2858
rect 1871 2826 1875 2830
rect 2239 2826 2243 2830
rect 2319 2826 2323 2830
rect 2359 2826 2363 2830
rect 2399 2826 2403 2830
rect 2455 2826 2459 2830
rect 2479 2826 2483 2830
rect 2559 2826 2563 2830
rect 2567 2826 2571 2830
rect 2663 2826 2667 2830
rect 2671 2826 2675 2830
rect 2767 2826 2771 2830
rect 2807 2826 2811 2830
rect 2879 2826 2883 2830
rect 2967 2826 2971 2830
rect 2991 2826 2995 2830
rect 3103 2826 3107 2830
rect 3143 2826 3147 2830
rect 3215 2826 3219 2830
rect 3335 2826 3339 2830
rect 3511 2826 3515 2830
rect 3591 2826 3595 2830
rect 111 2770 115 2774
rect 143 2770 147 2774
rect 271 2770 275 2774
rect 295 2770 299 2774
rect 399 2770 403 2774
rect 439 2770 443 2774
rect 535 2770 539 2774
rect 567 2770 571 2774
rect 663 2770 667 2774
rect 687 2770 691 2774
rect 791 2770 795 2774
rect 799 2770 803 2774
rect 903 2770 907 2774
rect 911 2770 915 2774
rect 1007 2770 1011 2774
rect 1031 2770 1035 2774
rect 1103 2770 1107 2774
rect 1143 2770 1147 2774
rect 1199 2770 1203 2774
rect 1263 2770 1267 2774
rect 1303 2770 1307 2774
rect 1383 2770 1387 2774
rect 1831 2770 1835 2774
rect 1871 2738 1875 2742
rect 2047 2738 2051 2742
rect 2135 2738 2139 2742
rect 2231 2738 2235 2742
rect 2311 2738 2315 2742
rect 2327 2738 2331 2742
rect 2391 2738 2395 2742
rect 2423 2738 2427 2742
rect 2471 2738 2475 2742
rect 2519 2738 2523 2742
rect 2559 2738 2563 2742
rect 2615 2738 2619 2742
rect 2663 2738 2667 2742
rect 2727 2738 2731 2742
rect 2799 2738 2803 2742
rect 2855 2738 2859 2742
rect 2959 2738 2963 2742
rect 3007 2738 3011 2742
rect 3135 2738 3139 2742
rect 3175 2738 3179 2742
rect 3327 2738 3331 2742
rect 3351 2738 3355 2742
rect 3503 2738 3507 2742
rect 3591 2738 3595 2742
rect 111 2690 115 2694
rect 143 2690 147 2694
rect 151 2690 155 2694
rect 263 2690 267 2694
rect 303 2690 307 2694
rect 407 2690 411 2694
rect 447 2690 451 2694
rect 543 2690 547 2694
rect 575 2690 579 2694
rect 671 2690 675 2694
rect 695 2690 699 2694
rect 791 2690 795 2694
rect 807 2690 811 2694
rect 903 2690 907 2694
rect 911 2690 915 2694
rect 1015 2690 1019 2694
rect 1111 2690 1115 2694
rect 1119 2690 1123 2694
rect 1207 2690 1211 2694
rect 1215 2690 1219 2694
rect 1311 2690 1315 2694
rect 1319 2690 1323 2694
rect 1423 2690 1427 2694
rect 1831 2690 1835 2694
rect 1871 2662 1875 2666
rect 2055 2662 2059 2666
rect 2071 2662 2075 2666
rect 2143 2662 2147 2666
rect 2239 2662 2243 2666
rect 2295 2662 2299 2666
rect 2335 2662 2339 2666
rect 2431 2662 2435 2666
rect 2527 2662 2531 2666
rect 2567 2662 2571 2666
rect 2623 2662 2627 2666
rect 2735 2662 2739 2666
rect 2863 2662 2867 2666
rect 2871 2662 2875 2666
rect 3015 2662 3019 2666
rect 3183 2662 3187 2666
rect 3199 2662 3203 2666
rect 3359 2662 3363 2666
rect 3511 2662 3515 2666
rect 3591 2662 3595 2666
rect 111 2606 115 2610
rect 135 2606 139 2610
rect 143 2606 147 2610
rect 255 2606 259 2610
rect 311 2606 315 2610
rect 399 2606 403 2610
rect 479 2606 483 2610
rect 535 2606 539 2610
rect 639 2606 643 2610
rect 663 2606 667 2610
rect 783 2606 787 2610
rect 791 2606 795 2610
rect 895 2606 899 2610
rect 927 2606 931 2610
rect 1007 2606 1011 2610
rect 1055 2606 1059 2610
rect 1111 2606 1115 2610
rect 1175 2606 1179 2610
rect 1207 2606 1211 2610
rect 1295 2606 1299 2610
rect 1311 2606 1315 2610
rect 1407 2606 1411 2610
rect 1415 2606 1419 2610
rect 1527 2606 1531 2610
rect 1831 2606 1835 2610
rect 1871 2582 1875 2586
rect 2063 2582 2067 2586
rect 2167 2582 2171 2586
rect 2263 2582 2267 2586
rect 2287 2582 2291 2586
rect 2367 2582 2371 2586
rect 2479 2582 2483 2586
rect 2559 2582 2563 2586
rect 2591 2582 2595 2586
rect 2695 2582 2699 2586
rect 2799 2582 2803 2586
rect 2863 2582 2867 2586
rect 2903 2582 2907 2586
rect 3015 2582 3019 2586
rect 3135 2582 3139 2586
rect 3191 2582 3195 2586
rect 3263 2582 3267 2586
rect 3391 2582 3395 2586
rect 3503 2582 3507 2586
rect 3591 2582 3595 2586
rect 111 2522 115 2526
rect 143 2522 147 2526
rect 151 2522 155 2526
rect 295 2522 299 2526
rect 319 2522 323 2526
rect 447 2522 451 2526
rect 487 2522 491 2526
rect 591 2522 595 2526
rect 647 2522 651 2526
rect 735 2522 739 2526
rect 799 2522 803 2526
rect 879 2522 883 2526
rect 935 2522 939 2526
rect 1015 2522 1019 2526
rect 1063 2522 1067 2526
rect 1143 2522 1147 2526
rect 1183 2522 1187 2526
rect 1271 2522 1275 2526
rect 1303 2522 1307 2526
rect 1399 2522 1403 2526
rect 1415 2522 1419 2526
rect 1535 2522 1539 2526
rect 1831 2522 1835 2526
rect 1871 2506 1875 2510
rect 2135 2506 2139 2510
rect 2175 2506 2179 2510
rect 2223 2506 2227 2510
rect 2271 2506 2275 2510
rect 2319 2506 2323 2510
rect 2375 2506 2379 2510
rect 2423 2506 2427 2510
rect 2487 2506 2491 2510
rect 2535 2506 2539 2510
rect 2599 2506 2603 2510
rect 2655 2506 2659 2510
rect 2703 2506 2707 2510
rect 2783 2506 2787 2510
rect 2807 2506 2811 2510
rect 2911 2506 2915 2510
rect 2919 2506 2923 2510
rect 3023 2506 3027 2510
rect 3063 2506 3067 2510
rect 3143 2506 3147 2510
rect 3215 2506 3219 2510
rect 3271 2506 3275 2510
rect 3375 2506 3379 2510
rect 3399 2506 3403 2510
rect 3511 2506 3515 2510
rect 3591 2506 3595 2510
rect 111 2442 115 2446
rect 135 2442 139 2446
rect 199 2442 203 2446
rect 287 2442 291 2446
rect 351 2442 355 2446
rect 439 2442 443 2446
rect 495 2442 499 2446
rect 583 2442 587 2446
rect 639 2442 643 2446
rect 727 2442 731 2446
rect 783 2442 787 2446
rect 871 2442 875 2446
rect 919 2442 923 2446
rect 1007 2442 1011 2446
rect 1047 2442 1051 2446
rect 1135 2442 1139 2446
rect 1175 2442 1179 2446
rect 1263 2442 1267 2446
rect 1311 2442 1315 2446
rect 1391 2442 1395 2446
rect 1447 2442 1451 2446
rect 1527 2442 1531 2446
rect 1831 2442 1835 2446
rect 1871 2422 1875 2426
rect 1975 2422 1979 2426
rect 2087 2422 2091 2426
rect 2127 2422 2131 2426
rect 2207 2422 2211 2426
rect 2215 2422 2219 2426
rect 2311 2422 2315 2426
rect 2335 2422 2339 2426
rect 2415 2422 2419 2426
rect 2479 2422 2483 2426
rect 2527 2422 2531 2426
rect 2631 2422 2635 2426
rect 2647 2422 2651 2426
rect 2775 2422 2779 2426
rect 2791 2422 2795 2426
rect 2911 2422 2915 2426
rect 2967 2422 2971 2426
rect 3055 2422 3059 2426
rect 3151 2422 3155 2426
rect 3207 2422 3211 2426
rect 3335 2422 3339 2426
rect 3367 2422 3371 2426
rect 3503 2422 3507 2426
rect 3591 2422 3595 2426
rect 111 2358 115 2362
rect 207 2358 211 2362
rect 223 2358 227 2362
rect 327 2358 331 2362
rect 359 2358 363 2362
rect 439 2358 443 2362
rect 503 2358 507 2362
rect 559 2358 563 2362
rect 647 2358 651 2362
rect 679 2358 683 2362
rect 791 2358 795 2362
rect 799 2358 803 2362
rect 911 2358 915 2362
rect 927 2358 931 2362
rect 1023 2358 1027 2362
rect 1055 2358 1059 2362
rect 1135 2358 1139 2362
rect 1183 2358 1187 2362
rect 1247 2358 1251 2362
rect 1319 2358 1323 2362
rect 1367 2358 1371 2362
rect 1455 2358 1459 2362
rect 1831 2358 1835 2362
rect 1871 2342 1875 2346
rect 1903 2342 1907 2346
rect 1983 2342 1987 2346
rect 2015 2342 2019 2346
rect 2095 2342 2099 2346
rect 2167 2342 2171 2346
rect 2215 2342 2219 2346
rect 2319 2342 2323 2346
rect 2343 2342 2347 2346
rect 2471 2342 2475 2346
rect 2487 2342 2491 2346
rect 2623 2342 2627 2346
rect 2639 2342 2643 2346
rect 2775 2342 2779 2346
rect 2799 2342 2803 2346
rect 2927 2342 2931 2346
rect 2975 2342 2979 2346
rect 3087 2342 3091 2346
rect 3159 2342 3163 2346
rect 3247 2342 3251 2346
rect 3343 2342 3347 2346
rect 3415 2342 3419 2346
rect 3511 2342 3515 2346
rect 3591 2342 3595 2346
rect 111 2270 115 2274
rect 215 2270 219 2274
rect 311 2270 315 2274
rect 319 2270 323 2274
rect 407 2270 411 2274
rect 431 2270 435 2274
rect 503 2270 507 2274
rect 551 2270 555 2274
rect 607 2270 611 2274
rect 671 2270 675 2274
rect 711 2270 715 2274
rect 791 2270 795 2274
rect 815 2270 819 2274
rect 903 2270 907 2274
rect 911 2270 915 2274
rect 1007 2270 1011 2274
rect 1015 2270 1019 2274
rect 1103 2270 1107 2274
rect 1127 2270 1131 2274
rect 1199 2270 1203 2274
rect 1239 2270 1243 2274
rect 1303 2270 1307 2274
rect 1359 2270 1363 2274
rect 1831 2270 1835 2274
rect 1871 2266 1875 2270
rect 1895 2266 1899 2270
rect 2007 2266 2011 2270
rect 2031 2266 2035 2270
rect 2159 2266 2163 2270
rect 2207 2266 2211 2270
rect 2311 2266 2315 2270
rect 2391 2266 2395 2270
rect 2463 2266 2467 2270
rect 2575 2266 2579 2270
rect 2615 2266 2619 2270
rect 2767 2266 2771 2270
rect 2919 2266 2923 2270
rect 2951 2266 2955 2270
rect 3079 2266 3083 2270
rect 3143 2266 3147 2270
rect 3239 2266 3243 2270
rect 3335 2266 3339 2270
rect 3407 2266 3411 2270
rect 3503 2266 3507 2270
rect 3591 2266 3595 2270
rect 111 2190 115 2194
rect 319 2190 323 2194
rect 415 2190 419 2194
rect 511 2190 515 2194
rect 519 2190 523 2194
rect 615 2190 619 2194
rect 623 2190 627 2194
rect 719 2190 723 2194
rect 727 2190 731 2194
rect 823 2190 827 2194
rect 831 2190 835 2194
rect 919 2190 923 2194
rect 935 2190 939 2194
rect 1015 2190 1019 2194
rect 1039 2190 1043 2194
rect 1111 2190 1115 2194
rect 1151 2190 1155 2194
rect 1207 2190 1211 2194
rect 1263 2190 1267 2194
rect 1311 2190 1315 2194
rect 1831 2190 1835 2194
rect 1871 2182 1875 2186
rect 1903 2182 1907 2186
rect 1967 2182 1971 2186
rect 2039 2182 2043 2186
rect 2079 2182 2083 2186
rect 2215 2182 2219 2186
rect 2367 2182 2371 2186
rect 2399 2182 2403 2186
rect 2527 2182 2531 2186
rect 2583 2182 2587 2186
rect 2687 2182 2691 2186
rect 2775 2182 2779 2186
rect 2847 2182 2851 2186
rect 2959 2182 2963 2186
rect 2991 2182 2995 2186
rect 3127 2182 3131 2186
rect 3151 2182 3155 2186
rect 3263 2182 3267 2186
rect 3343 2182 3347 2186
rect 3399 2182 3403 2186
rect 3511 2182 3515 2186
rect 3591 2182 3595 2186
rect 111 2114 115 2118
rect 279 2114 283 2118
rect 311 2114 315 2118
rect 399 2114 403 2118
rect 407 2114 411 2118
rect 511 2114 515 2118
rect 615 2114 619 2118
rect 623 2114 627 2118
rect 719 2114 723 2118
rect 735 2114 739 2118
rect 823 2114 827 2118
rect 847 2114 851 2118
rect 927 2114 931 2118
rect 951 2114 955 2118
rect 1031 2114 1035 2118
rect 1047 2114 1051 2118
rect 1143 2114 1147 2118
rect 1239 2114 1243 2118
rect 1255 2114 1259 2118
rect 1343 2114 1347 2118
rect 1831 2114 1835 2118
rect 1871 2106 1875 2110
rect 1959 2106 1963 2110
rect 2071 2106 2075 2110
rect 2207 2106 2211 2110
rect 2287 2106 2291 2110
rect 2359 2106 2363 2110
rect 2391 2106 2395 2110
rect 2503 2106 2507 2110
rect 2519 2106 2523 2110
rect 2623 2106 2627 2110
rect 2679 2106 2683 2110
rect 2743 2106 2747 2110
rect 2839 2106 2843 2110
rect 2855 2106 2859 2110
rect 2967 2106 2971 2110
rect 2983 2106 2987 2110
rect 3079 2106 3083 2110
rect 3119 2106 3123 2110
rect 3191 2106 3195 2110
rect 3255 2106 3259 2110
rect 3303 2106 3307 2110
rect 3391 2106 3395 2110
rect 3415 2106 3419 2110
rect 3503 2106 3507 2110
rect 3591 2106 3595 2110
rect 111 2030 115 2034
rect 183 2030 187 2034
rect 287 2030 291 2034
rect 327 2030 331 2034
rect 407 2030 411 2034
rect 471 2030 475 2034
rect 519 2030 523 2034
rect 623 2030 627 2034
rect 631 2030 635 2034
rect 743 2030 747 2034
rect 767 2030 771 2034
rect 855 2030 859 2034
rect 911 2030 915 2034
rect 959 2030 963 2034
rect 1047 2030 1051 2034
rect 1055 2030 1059 2034
rect 1151 2030 1155 2034
rect 1183 2030 1187 2034
rect 1247 2030 1251 2034
rect 1319 2030 1323 2034
rect 1351 2030 1355 2034
rect 1463 2030 1467 2034
rect 1831 2030 1835 2034
rect 1871 2026 1875 2030
rect 2183 2026 2187 2030
rect 2271 2026 2275 2030
rect 2295 2026 2299 2030
rect 2367 2026 2371 2030
rect 2399 2026 2403 2030
rect 2463 2026 2467 2030
rect 2511 2026 2515 2030
rect 2567 2026 2571 2030
rect 2631 2026 2635 2030
rect 2671 2026 2675 2030
rect 2751 2026 2755 2030
rect 2775 2026 2779 2030
rect 2863 2026 2867 2030
rect 2879 2026 2883 2030
rect 2975 2026 2979 2030
rect 2983 2026 2987 2030
rect 3087 2026 3091 2030
rect 3191 2026 3195 2030
rect 3199 2026 3203 2030
rect 3311 2026 3315 2030
rect 3423 2026 3427 2030
rect 3511 2026 3515 2030
rect 3591 2026 3595 2030
rect 111 1954 115 1958
rect 135 1954 139 1958
rect 175 1954 179 1958
rect 295 1954 299 1958
rect 319 1954 323 1958
rect 463 1954 467 1958
rect 615 1954 619 1958
rect 631 1954 635 1958
rect 759 1954 763 1958
rect 799 1954 803 1958
rect 903 1954 907 1958
rect 951 1954 955 1958
rect 1039 1954 1043 1958
rect 1095 1954 1099 1958
rect 1175 1954 1179 1958
rect 1231 1954 1235 1958
rect 1311 1954 1315 1958
rect 1359 1954 1363 1958
rect 1455 1954 1459 1958
rect 1487 1954 1491 1958
rect 1623 1954 1627 1958
rect 1831 1954 1835 1958
rect 1871 1946 1875 1950
rect 1943 1946 1947 1950
rect 2055 1946 2059 1950
rect 2167 1946 2171 1950
rect 2175 1946 2179 1950
rect 2263 1946 2267 1950
rect 2287 1946 2291 1950
rect 2359 1946 2363 1950
rect 2407 1946 2411 1950
rect 2455 1946 2459 1950
rect 2527 1946 2531 1950
rect 2559 1946 2563 1950
rect 2647 1946 2651 1950
rect 2663 1946 2667 1950
rect 2767 1946 2771 1950
rect 2775 1946 2779 1950
rect 2871 1946 2875 1950
rect 2911 1946 2915 1950
rect 2975 1946 2979 1950
rect 3055 1946 3059 1950
rect 3079 1946 3083 1950
rect 3183 1946 3187 1950
rect 3207 1946 3211 1950
rect 3367 1946 3371 1950
rect 3503 1946 3507 1950
rect 3591 1946 3595 1950
rect 111 1870 115 1874
rect 143 1870 147 1874
rect 303 1870 307 1874
rect 319 1870 323 1874
rect 471 1870 475 1874
rect 519 1870 523 1874
rect 639 1870 643 1874
rect 711 1870 715 1874
rect 807 1870 811 1874
rect 887 1870 891 1874
rect 959 1870 963 1874
rect 1055 1870 1059 1874
rect 1103 1870 1107 1874
rect 1207 1870 1211 1874
rect 1239 1870 1243 1874
rect 1343 1870 1347 1874
rect 1367 1870 1371 1874
rect 1471 1870 1475 1874
rect 1495 1870 1499 1874
rect 1599 1870 1603 1874
rect 1631 1870 1635 1874
rect 1727 1870 1731 1874
rect 1831 1870 1835 1874
rect 1871 1866 1875 1870
rect 1903 1866 1907 1870
rect 1951 1866 1955 1870
rect 1983 1866 1987 1870
rect 2063 1866 2067 1870
rect 2095 1866 2099 1870
rect 2175 1866 2179 1870
rect 2207 1866 2211 1870
rect 2295 1866 2299 1870
rect 2327 1866 2331 1870
rect 2415 1866 2419 1870
rect 2463 1866 2467 1870
rect 2535 1866 2539 1870
rect 2631 1866 2635 1870
rect 2655 1866 2659 1870
rect 2783 1866 2787 1870
rect 2831 1866 2835 1870
rect 2919 1866 2923 1870
rect 3055 1866 3059 1870
rect 3063 1866 3067 1870
rect 3215 1866 3219 1870
rect 3295 1866 3299 1870
rect 3375 1866 3379 1870
rect 3511 1866 3515 1870
rect 3591 1866 3595 1870
rect 111 1794 115 1798
rect 135 1794 139 1798
rect 311 1794 315 1798
rect 503 1794 507 1798
rect 511 1794 515 1798
rect 687 1794 691 1798
rect 703 1794 707 1798
rect 847 1794 851 1798
rect 879 1794 883 1798
rect 991 1794 995 1798
rect 1047 1794 1051 1798
rect 1127 1794 1131 1798
rect 1199 1794 1203 1798
rect 1247 1794 1251 1798
rect 1335 1794 1339 1798
rect 1359 1794 1363 1798
rect 1463 1794 1467 1798
rect 1559 1794 1563 1798
rect 1591 1794 1595 1798
rect 1663 1794 1667 1798
rect 1719 1794 1723 1798
rect 1743 1794 1747 1798
rect 1831 1794 1835 1798
rect 1871 1774 1875 1778
rect 1895 1774 1899 1778
rect 1975 1774 1979 1778
rect 2023 1774 2027 1778
rect 2087 1774 2091 1778
rect 2183 1774 2187 1778
rect 2199 1774 2203 1778
rect 2319 1774 2323 1778
rect 2351 1774 2355 1778
rect 2455 1774 2459 1778
rect 2551 1774 2555 1778
rect 2623 1774 2627 1778
rect 2775 1774 2779 1778
rect 2823 1774 2827 1778
rect 3015 1774 3019 1778
rect 3047 1774 3051 1778
rect 3271 1774 3275 1778
rect 3287 1774 3291 1778
rect 3503 1774 3507 1778
rect 3591 1774 3595 1778
rect 111 1710 115 1714
rect 143 1710 147 1714
rect 239 1710 243 1714
rect 319 1710 323 1714
rect 367 1710 371 1714
rect 487 1710 491 1714
rect 511 1710 515 1714
rect 607 1710 611 1714
rect 695 1710 699 1714
rect 719 1710 723 1714
rect 823 1710 827 1714
rect 855 1710 859 1714
rect 927 1710 931 1714
rect 999 1710 1003 1714
rect 1023 1710 1027 1714
rect 1119 1710 1123 1714
rect 1135 1710 1139 1714
rect 1215 1710 1219 1714
rect 1255 1710 1259 1714
rect 1319 1710 1323 1714
rect 1367 1710 1371 1714
rect 1471 1710 1475 1714
rect 1567 1710 1571 1714
rect 1671 1710 1675 1714
rect 1751 1710 1755 1714
rect 1831 1710 1835 1714
rect 1871 1698 1875 1702
rect 1903 1698 1907 1702
rect 1991 1698 1995 1702
rect 2031 1698 2035 1702
rect 2111 1698 2115 1702
rect 2191 1698 2195 1702
rect 2231 1698 2235 1702
rect 2351 1698 2355 1702
rect 2359 1698 2363 1702
rect 2479 1698 2483 1702
rect 2559 1698 2563 1702
rect 2607 1698 2611 1702
rect 2743 1698 2747 1702
rect 2783 1698 2787 1702
rect 2887 1698 2891 1702
rect 3023 1698 3027 1702
rect 3039 1698 3043 1702
rect 3199 1698 3203 1702
rect 3279 1698 3283 1702
rect 3367 1698 3371 1702
rect 3511 1698 3515 1702
rect 3591 1698 3595 1702
rect 111 1626 115 1630
rect 135 1626 139 1630
rect 175 1626 179 1630
rect 231 1626 235 1630
rect 311 1626 315 1630
rect 359 1626 363 1630
rect 439 1626 443 1630
rect 479 1626 483 1630
rect 567 1626 571 1630
rect 599 1626 603 1630
rect 687 1626 691 1630
rect 711 1626 715 1630
rect 799 1626 803 1630
rect 815 1626 819 1630
rect 903 1626 907 1630
rect 919 1626 923 1630
rect 999 1626 1003 1630
rect 1015 1626 1019 1630
rect 1095 1626 1099 1630
rect 1111 1626 1115 1630
rect 1199 1626 1203 1630
rect 1207 1626 1211 1630
rect 1303 1626 1307 1630
rect 1311 1626 1315 1630
rect 1831 1626 1835 1630
rect 1871 1622 1875 1626
rect 1895 1622 1899 1626
rect 1927 1622 1931 1626
rect 1983 1622 1987 1626
rect 2023 1622 2027 1626
rect 2103 1622 2107 1626
rect 2135 1622 2139 1626
rect 2223 1622 2227 1626
rect 2263 1622 2267 1626
rect 2343 1622 2347 1626
rect 2391 1622 2395 1626
rect 2471 1622 2475 1626
rect 2527 1622 2531 1626
rect 2599 1622 2603 1626
rect 2671 1622 2675 1626
rect 2735 1622 2739 1626
rect 2823 1622 2827 1626
rect 2879 1622 2883 1626
rect 2983 1622 2987 1626
rect 3031 1622 3035 1626
rect 3159 1622 3163 1626
rect 3191 1622 3195 1626
rect 3343 1622 3347 1626
rect 3359 1622 3363 1626
rect 3503 1622 3507 1626
rect 3591 1622 3595 1626
rect 111 1542 115 1546
rect 183 1542 187 1546
rect 239 1542 243 1546
rect 319 1542 323 1546
rect 343 1542 347 1546
rect 447 1542 451 1546
rect 463 1542 467 1546
rect 575 1542 579 1546
rect 591 1542 595 1546
rect 695 1542 699 1546
rect 719 1542 723 1546
rect 807 1542 811 1546
rect 855 1542 859 1546
rect 911 1542 915 1546
rect 983 1542 987 1546
rect 1007 1542 1011 1546
rect 1103 1542 1107 1546
rect 1111 1542 1115 1546
rect 1207 1542 1211 1546
rect 1231 1542 1235 1546
rect 1311 1542 1315 1546
rect 1343 1542 1347 1546
rect 1455 1542 1459 1546
rect 1575 1542 1579 1546
rect 1831 1542 1835 1546
rect 1871 1538 1875 1542
rect 1935 1538 1939 1542
rect 2031 1538 2035 1542
rect 2135 1538 2139 1542
rect 2143 1538 2147 1542
rect 2255 1538 2259 1542
rect 2271 1538 2275 1542
rect 2383 1538 2387 1542
rect 2399 1538 2403 1542
rect 2511 1538 2515 1542
rect 2535 1538 2539 1542
rect 2639 1538 2643 1542
rect 2679 1538 2683 1542
rect 2767 1538 2771 1542
rect 2831 1538 2835 1542
rect 2887 1538 2891 1542
rect 2991 1538 2995 1542
rect 3007 1538 3011 1542
rect 3119 1538 3123 1542
rect 3167 1538 3171 1542
rect 3231 1538 3235 1542
rect 3351 1538 3355 1542
rect 3511 1538 3515 1542
rect 3591 1538 3595 1542
rect 111 1454 115 1458
rect 231 1454 235 1458
rect 279 1454 283 1458
rect 335 1454 339 1458
rect 383 1454 387 1458
rect 455 1454 459 1458
rect 511 1454 515 1458
rect 583 1454 587 1458
rect 655 1454 659 1458
rect 711 1454 715 1458
rect 807 1454 811 1458
rect 847 1454 851 1458
rect 959 1454 963 1458
rect 975 1454 979 1458
rect 1103 1454 1107 1458
rect 1111 1454 1115 1458
rect 1223 1454 1227 1458
rect 1247 1454 1251 1458
rect 1335 1454 1339 1458
rect 1383 1454 1387 1458
rect 1447 1454 1451 1458
rect 1511 1454 1515 1458
rect 1567 1454 1571 1458
rect 1639 1454 1643 1458
rect 1743 1454 1747 1458
rect 1831 1454 1835 1458
rect 1871 1454 1875 1458
rect 2127 1454 2131 1458
rect 2247 1454 2251 1458
rect 2343 1454 2347 1458
rect 2375 1454 2379 1458
rect 2455 1454 2459 1458
rect 2503 1454 2507 1458
rect 2575 1454 2579 1458
rect 2631 1454 2635 1458
rect 2703 1454 2707 1458
rect 2759 1454 2763 1458
rect 2831 1454 2835 1458
rect 2879 1454 2883 1458
rect 2951 1454 2955 1458
rect 2999 1454 3003 1458
rect 3071 1454 3075 1458
rect 3111 1454 3115 1458
rect 3183 1454 3187 1458
rect 3223 1454 3227 1458
rect 3295 1454 3299 1458
rect 3343 1454 3347 1458
rect 3407 1454 3411 1458
rect 3503 1454 3507 1458
rect 3591 1454 3595 1458
rect 1871 1370 1875 1374
rect 2255 1370 2259 1374
rect 2351 1370 2355 1374
rect 2399 1370 2403 1374
rect 2463 1370 2467 1374
rect 2503 1370 2507 1374
rect 2583 1370 2587 1374
rect 2615 1370 2619 1374
rect 2711 1370 2715 1374
rect 2735 1370 2739 1374
rect 2839 1370 2843 1374
rect 2847 1370 2851 1374
rect 2959 1370 2963 1374
rect 3071 1370 3075 1374
rect 3079 1370 3083 1374
rect 3183 1370 3187 1374
rect 3191 1370 3195 1374
rect 3295 1370 3299 1374
rect 3303 1370 3307 1374
rect 3415 1370 3419 1374
rect 3511 1370 3515 1374
rect 3591 1370 3595 1374
rect 111 1362 115 1366
rect 223 1362 227 1366
rect 287 1362 291 1366
rect 335 1362 339 1366
rect 391 1362 395 1366
rect 471 1362 475 1366
rect 519 1362 523 1366
rect 623 1362 627 1366
rect 663 1362 667 1366
rect 783 1362 787 1366
rect 815 1362 819 1366
rect 943 1362 947 1366
rect 967 1362 971 1366
rect 1095 1362 1099 1366
rect 1119 1362 1123 1366
rect 1239 1362 1243 1366
rect 1255 1362 1259 1366
rect 1375 1362 1379 1366
rect 1391 1362 1395 1366
rect 1511 1362 1515 1366
rect 1519 1362 1523 1366
rect 1639 1362 1643 1366
rect 1647 1362 1651 1366
rect 1751 1362 1755 1366
rect 1831 1362 1835 1366
rect 111 1286 115 1290
rect 135 1286 139 1290
rect 215 1286 219 1290
rect 327 1286 331 1290
rect 335 1286 339 1290
rect 463 1286 467 1290
rect 607 1286 611 1290
rect 615 1286 619 1290
rect 751 1286 755 1290
rect 775 1286 779 1290
rect 903 1286 907 1290
rect 935 1286 939 1290
rect 1047 1286 1051 1290
rect 1087 1286 1091 1290
rect 1183 1286 1187 1290
rect 1231 1286 1235 1290
rect 1303 1286 1307 1290
rect 1367 1286 1371 1290
rect 1423 1286 1427 1290
rect 1503 1286 1507 1290
rect 1535 1286 1539 1290
rect 1631 1286 1635 1290
rect 1647 1286 1651 1290
rect 1743 1286 1747 1290
rect 1831 1286 1835 1290
rect 1871 1278 1875 1282
rect 1895 1278 1899 1282
rect 2071 1278 2075 1282
rect 2255 1278 2259 1282
rect 2391 1278 2395 1282
rect 2423 1278 2427 1282
rect 2495 1278 2499 1282
rect 2583 1278 2587 1282
rect 2607 1278 2611 1282
rect 2727 1278 2731 1282
rect 2735 1278 2739 1282
rect 2839 1278 2843 1282
rect 2879 1278 2883 1282
rect 2951 1278 2955 1282
rect 3015 1278 3019 1282
rect 3063 1278 3067 1282
rect 3143 1278 3147 1282
rect 3175 1278 3179 1282
rect 3271 1278 3275 1282
rect 3287 1278 3291 1282
rect 3399 1278 3403 1282
rect 3407 1278 3411 1282
rect 3503 1278 3507 1282
rect 3591 1278 3595 1282
rect 111 1198 115 1202
rect 143 1198 147 1202
rect 223 1198 227 1202
rect 255 1198 259 1202
rect 343 1198 347 1202
rect 383 1198 387 1202
rect 471 1198 475 1202
rect 503 1198 507 1202
rect 615 1198 619 1202
rect 719 1198 723 1202
rect 759 1198 763 1202
rect 815 1198 819 1202
rect 911 1198 915 1202
rect 999 1198 1003 1202
rect 1055 1198 1059 1202
rect 1095 1198 1099 1202
rect 1191 1198 1195 1202
rect 1287 1198 1291 1202
rect 1311 1198 1315 1202
rect 1431 1198 1435 1202
rect 1543 1198 1547 1202
rect 1655 1198 1659 1202
rect 1751 1198 1755 1202
rect 1831 1198 1835 1202
rect 1871 1194 1875 1198
rect 1903 1194 1907 1198
rect 1991 1194 1995 1198
rect 2079 1194 2083 1198
rect 2103 1194 2107 1198
rect 2215 1194 2219 1198
rect 2263 1194 2267 1198
rect 2327 1194 2331 1198
rect 2431 1194 2435 1198
rect 2447 1194 2451 1198
rect 2575 1194 2579 1198
rect 2591 1194 2595 1198
rect 2719 1194 2723 1198
rect 2743 1194 2747 1198
rect 2871 1194 2875 1198
rect 2887 1194 2891 1198
rect 3023 1194 3027 1198
rect 3031 1194 3035 1198
rect 3151 1194 3155 1198
rect 3191 1194 3195 1198
rect 3279 1194 3283 1198
rect 3359 1194 3363 1198
rect 3407 1194 3411 1198
rect 3511 1194 3515 1198
rect 3591 1194 3595 1198
rect 111 1110 115 1114
rect 135 1110 139 1114
rect 247 1110 251 1114
rect 255 1110 259 1114
rect 375 1110 379 1114
rect 399 1110 403 1114
rect 495 1110 499 1114
rect 535 1110 539 1114
rect 607 1110 611 1114
rect 663 1110 667 1114
rect 711 1110 715 1114
rect 783 1110 787 1114
rect 807 1110 811 1114
rect 895 1110 899 1114
rect 903 1110 907 1114
rect 991 1110 995 1114
rect 999 1110 1003 1114
rect 1087 1110 1091 1114
rect 1095 1110 1099 1114
rect 1183 1110 1187 1114
rect 1191 1110 1195 1114
rect 1279 1110 1283 1114
rect 1295 1110 1299 1114
rect 1399 1110 1403 1114
rect 1831 1110 1835 1114
rect 1871 1110 1875 1114
rect 1895 1110 1899 1114
rect 1967 1110 1971 1114
rect 1983 1110 1987 1114
rect 2047 1110 2051 1114
rect 2095 1110 2099 1114
rect 2135 1110 2139 1114
rect 2207 1110 2211 1114
rect 2231 1110 2235 1114
rect 2319 1110 2323 1114
rect 2335 1110 2339 1114
rect 2439 1110 2443 1114
rect 2551 1110 2555 1114
rect 2567 1110 2571 1114
rect 2679 1110 2683 1114
rect 2711 1110 2715 1114
rect 2823 1110 2827 1114
rect 2863 1110 2867 1114
rect 2983 1110 2987 1114
rect 3023 1110 3027 1114
rect 3159 1110 3163 1114
rect 3183 1110 3187 1114
rect 3343 1110 3347 1114
rect 3351 1110 3355 1114
rect 3503 1110 3507 1114
rect 3591 1110 3595 1114
rect 111 1026 115 1030
rect 143 1026 147 1030
rect 263 1026 267 1030
rect 271 1026 275 1030
rect 407 1026 411 1030
rect 423 1026 427 1030
rect 543 1026 547 1030
rect 583 1026 587 1030
rect 671 1026 675 1030
rect 735 1026 739 1030
rect 791 1026 795 1030
rect 887 1026 891 1030
rect 903 1026 907 1030
rect 1007 1026 1011 1030
rect 1031 1026 1035 1030
rect 1103 1026 1107 1030
rect 1159 1026 1163 1030
rect 1199 1026 1203 1030
rect 1279 1026 1283 1030
rect 1303 1026 1307 1030
rect 1399 1026 1403 1030
rect 1407 1026 1411 1030
rect 1519 1026 1523 1030
rect 1639 1026 1643 1030
rect 1831 1026 1835 1030
rect 1871 1026 1875 1030
rect 1975 1026 1979 1030
rect 2031 1026 2035 1030
rect 2055 1026 2059 1030
rect 2127 1026 2131 1030
rect 2143 1026 2147 1030
rect 2231 1026 2235 1030
rect 2239 1026 2243 1030
rect 2343 1026 2347 1030
rect 2351 1026 2355 1030
rect 2447 1026 2451 1030
rect 2471 1026 2475 1030
rect 2559 1026 2563 1030
rect 2599 1026 2603 1030
rect 2687 1026 2691 1030
rect 2727 1026 2731 1030
rect 2831 1026 2835 1030
rect 2855 1026 2859 1030
rect 2983 1026 2987 1030
rect 2991 1026 2995 1030
rect 3111 1026 3115 1030
rect 3167 1026 3171 1030
rect 3247 1026 3251 1030
rect 3351 1026 3355 1030
rect 3391 1026 3395 1030
rect 3511 1026 3515 1030
rect 3591 1026 3595 1030
rect 111 942 115 946
rect 135 942 139 946
rect 215 942 219 946
rect 263 942 267 946
rect 335 942 339 946
rect 415 942 419 946
rect 463 942 467 946
rect 575 942 579 946
rect 599 942 603 946
rect 727 942 731 946
rect 735 942 739 946
rect 863 942 867 946
rect 879 942 883 946
rect 991 942 995 946
rect 1023 942 1027 946
rect 1111 942 1115 946
rect 1151 942 1155 946
rect 1223 942 1227 946
rect 1271 942 1275 946
rect 1335 942 1339 946
rect 1391 942 1395 946
rect 1455 942 1459 946
rect 1511 942 1515 946
rect 1631 942 1635 946
rect 1831 942 1835 946
rect 1871 942 1875 946
rect 1895 942 1899 946
rect 1983 942 1987 946
rect 2023 942 2027 946
rect 2111 942 2115 946
rect 2119 942 2123 946
rect 2223 942 2227 946
rect 2263 942 2267 946
rect 2343 942 2347 946
rect 2423 942 2427 946
rect 2463 942 2467 946
rect 2583 942 2587 946
rect 2591 942 2595 946
rect 2719 942 2723 946
rect 2735 942 2739 946
rect 2847 942 2851 946
rect 2879 942 2883 946
rect 2975 942 2979 946
rect 3015 942 3019 946
rect 3103 942 3107 946
rect 3143 942 3147 946
rect 3239 942 3243 946
rect 3271 942 3275 946
rect 3383 942 3387 946
rect 3399 942 3403 946
rect 3503 942 3507 946
rect 3591 942 3595 946
rect 111 854 115 858
rect 143 854 147 858
rect 223 854 227 858
rect 303 854 307 858
rect 343 854 347 858
rect 391 854 395 858
rect 471 854 475 858
rect 495 854 499 858
rect 599 854 603 858
rect 607 854 611 858
rect 711 854 715 858
rect 743 854 747 858
rect 839 854 843 858
rect 871 854 875 858
rect 991 854 995 858
rect 999 854 1003 858
rect 1119 854 1123 858
rect 1167 854 1171 858
rect 1231 854 1235 858
rect 1343 854 1347 858
rect 1359 854 1363 858
rect 1463 854 1467 858
rect 1567 854 1571 858
rect 1751 854 1755 858
rect 1831 854 1835 858
rect 1871 858 1875 862
rect 1903 858 1907 862
rect 1991 858 1995 862
rect 2039 858 2043 862
rect 2119 858 2123 862
rect 2215 858 2219 862
rect 2271 858 2275 862
rect 2391 858 2395 862
rect 2431 858 2435 862
rect 2567 858 2571 862
rect 2591 858 2595 862
rect 2735 858 2739 862
rect 2743 858 2747 862
rect 2887 858 2891 862
rect 3023 858 3027 862
rect 3031 858 3035 862
rect 3151 858 3155 862
rect 3159 858 3163 862
rect 3279 858 3283 862
rect 3287 858 3291 862
rect 3407 858 3411 862
rect 3511 858 3515 862
rect 3591 858 3595 862
rect 111 774 115 778
rect 135 774 139 778
rect 199 774 203 778
rect 215 774 219 778
rect 287 774 291 778
rect 295 774 299 778
rect 383 774 387 778
rect 391 774 395 778
rect 487 774 491 778
rect 503 774 507 778
rect 591 774 595 778
rect 615 774 619 778
rect 703 774 707 778
rect 735 774 739 778
rect 831 774 835 778
rect 855 774 859 778
rect 983 774 987 778
rect 1111 774 1115 778
rect 1159 774 1163 778
rect 1239 774 1243 778
rect 1351 774 1355 778
rect 1367 774 1371 778
rect 1495 774 1499 778
rect 1559 774 1563 778
rect 1631 774 1635 778
rect 1743 774 1747 778
rect 1831 774 1835 778
rect 1871 766 1875 770
rect 1895 766 1899 770
rect 2023 766 2027 770
rect 2031 766 2035 770
rect 2191 766 2195 770
rect 2207 766 2211 770
rect 2359 766 2363 770
rect 2383 766 2387 770
rect 2519 766 2523 770
rect 2559 766 2563 770
rect 2679 766 2683 770
rect 2727 766 2731 770
rect 2831 766 2835 770
rect 2879 766 2883 770
rect 2975 766 2979 770
rect 3023 766 3027 770
rect 3111 766 3115 770
rect 3151 766 3155 770
rect 3247 766 3251 770
rect 3279 766 3283 770
rect 3383 766 3387 770
rect 3399 766 3403 770
rect 3503 766 3507 770
rect 3591 766 3595 770
rect 111 682 115 686
rect 207 682 211 686
rect 295 682 299 686
rect 383 682 387 686
rect 399 682 403 686
rect 479 682 483 686
rect 511 682 515 686
rect 591 682 595 686
rect 623 682 627 686
rect 719 682 723 686
rect 743 682 747 686
rect 855 682 859 686
rect 863 682 867 686
rect 991 682 995 686
rect 1119 682 1123 686
rect 1127 682 1131 686
rect 1247 682 1251 686
rect 1255 682 1259 686
rect 1375 682 1379 686
rect 1383 682 1387 686
rect 1503 682 1507 686
rect 1631 682 1635 686
rect 1639 682 1643 686
rect 1751 682 1755 686
rect 1831 682 1835 686
rect 1871 686 1875 690
rect 2031 686 2035 690
rect 2095 686 2099 690
rect 2175 686 2179 690
rect 2199 686 2203 690
rect 2263 686 2267 690
rect 2359 686 2363 690
rect 2367 686 2371 690
rect 2463 686 2467 690
rect 2527 686 2531 690
rect 2567 686 2571 690
rect 2679 686 2683 690
rect 2687 686 2691 690
rect 2799 686 2803 690
rect 2839 686 2843 690
rect 2927 686 2931 690
rect 2983 686 2987 690
rect 3071 686 3075 690
rect 3119 686 3123 690
rect 3223 686 3227 690
rect 3255 686 3259 690
rect 3375 686 3379 690
rect 3391 686 3395 690
rect 3511 686 3515 690
rect 3591 686 3595 690
rect 111 598 115 602
rect 375 598 379 602
rect 471 598 475 602
rect 583 598 587 602
rect 599 598 603 602
rect 687 598 691 602
rect 711 598 715 602
rect 783 598 787 602
rect 847 598 851 602
rect 887 598 891 602
rect 983 598 987 602
rect 991 598 995 602
rect 1095 598 1099 602
rect 1119 598 1123 602
rect 1199 598 1203 602
rect 1247 598 1251 602
rect 1303 598 1307 602
rect 1375 598 1379 602
rect 1399 598 1403 602
rect 1495 598 1499 602
rect 1503 598 1507 602
rect 1607 598 1611 602
rect 1623 598 1627 602
rect 1711 598 1715 602
rect 1743 598 1747 602
rect 1831 598 1835 602
rect 1871 598 1875 602
rect 2087 598 2091 602
rect 2167 598 2171 602
rect 2247 598 2251 602
rect 2255 598 2259 602
rect 2327 598 2331 602
rect 2351 598 2355 602
rect 2407 598 2411 602
rect 2455 598 2459 602
rect 2487 598 2491 602
rect 2559 598 2563 602
rect 2567 598 2571 602
rect 2647 598 2651 602
rect 2671 598 2675 602
rect 2743 598 2747 602
rect 2791 598 2795 602
rect 2863 598 2867 602
rect 2919 598 2923 602
rect 2999 598 3003 602
rect 3063 598 3067 602
rect 3159 598 3163 602
rect 3215 598 3219 602
rect 3327 598 3331 602
rect 3367 598 3371 602
rect 3495 598 3499 602
rect 3503 598 3507 602
rect 3591 598 3595 602
rect 111 514 115 518
rect 367 514 371 518
rect 463 514 467 518
rect 575 514 579 518
rect 607 514 611 518
rect 695 514 699 518
rect 703 514 707 518
rect 791 514 795 518
rect 839 514 843 518
rect 895 514 899 518
rect 975 514 979 518
rect 999 514 1003 518
rect 1103 514 1107 518
rect 1111 514 1115 518
rect 1207 514 1211 518
rect 1239 514 1243 518
rect 1311 514 1315 518
rect 1359 514 1363 518
rect 1407 514 1411 518
rect 1471 514 1475 518
rect 1511 514 1515 518
rect 1583 514 1587 518
rect 1615 514 1619 518
rect 1703 514 1707 518
rect 1719 514 1723 518
rect 1831 514 1835 518
rect 1871 514 1875 518
rect 2159 514 2163 518
rect 2175 514 2179 518
rect 2239 514 2243 518
rect 2255 514 2259 518
rect 2319 514 2323 518
rect 2335 514 2339 518
rect 2399 514 2403 518
rect 2415 514 2419 518
rect 2479 514 2483 518
rect 2495 514 2499 518
rect 2559 514 2563 518
rect 2575 514 2579 518
rect 2639 514 2643 518
rect 2655 514 2659 518
rect 2735 514 2739 518
rect 2751 514 2755 518
rect 2855 514 2859 518
rect 2871 514 2875 518
rect 2991 514 2995 518
rect 3007 514 3011 518
rect 3143 514 3147 518
rect 3167 514 3171 518
rect 3311 514 3315 518
rect 3335 514 3339 518
rect 3479 514 3483 518
rect 3503 514 3507 518
rect 3591 514 3595 518
rect 111 426 115 430
rect 135 426 139 430
rect 223 426 227 430
rect 359 426 363 430
rect 455 426 459 430
rect 511 426 515 430
rect 567 426 571 430
rect 679 426 683 430
rect 695 426 699 430
rect 831 426 835 430
rect 839 426 843 430
rect 967 426 971 430
rect 999 426 1003 430
rect 1103 426 1107 430
rect 1143 426 1147 430
rect 1231 426 1235 430
rect 1279 426 1283 430
rect 1351 426 1355 430
rect 1415 426 1419 430
rect 1463 426 1467 430
rect 1551 426 1555 430
rect 1575 426 1579 430
rect 1687 426 1691 430
rect 1695 426 1699 430
rect 1831 426 1835 430
rect 1871 426 1875 430
rect 2151 426 2155 430
rect 2159 426 2163 430
rect 2231 426 2235 430
rect 2239 426 2243 430
rect 2311 426 2315 430
rect 2319 426 2323 430
rect 2391 426 2395 430
rect 2399 426 2403 430
rect 2471 426 2475 430
rect 2479 426 2483 430
rect 2551 426 2555 430
rect 2559 426 2563 430
rect 2631 426 2635 430
rect 2639 426 2643 430
rect 2727 426 2731 430
rect 2735 426 2739 430
rect 2839 426 2843 430
rect 2847 426 2851 430
rect 2959 426 2963 430
rect 2983 426 2987 430
rect 3087 426 3091 430
rect 3135 426 3139 430
rect 3231 426 3235 430
rect 3303 426 3307 430
rect 3375 426 3379 430
rect 3471 426 3475 430
rect 3503 426 3507 430
rect 3591 426 3595 430
rect 111 342 115 346
rect 143 342 147 346
rect 231 342 235 346
rect 279 342 283 346
rect 367 342 371 346
rect 455 342 459 346
rect 519 342 523 346
rect 639 342 643 346
rect 687 342 691 346
rect 823 342 827 346
rect 847 342 851 346
rect 999 342 1003 346
rect 1007 342 1011 346
rect 1151 342 1155 346
rect 1167 342 1171 346
rect 1287 342 1291 346
rect 1327 342 1331 346
rect 1423 342 1427 346
rect 1479 342 1483 346
rect 1559 342 1563 346
rect 1623 342 1627 346
rect 1695 342 1699 346
rect 1751 342 1755 346
rect 1831 342 1835 346
rect 1871 338 1875 342
rect 2031 338 2035 342
rect 2119 338 2123 342
rect 2167 338 2171 342
rect 2223 338 2227 342
rect 2247 338 2251 342
rect 2327 338 2331 342
rect 2335 338 2339 342
rect 2407 338 2411 342
rect 2447 338 2451 342
rect 2487 338 2491 342
rect 2567 338 2571 342
rect 2647 338 2651 342
rect 2695 338 2699 342
rect 2743 338 2747 342
rect 2839 338 2843 342
rect 2847 338 2851 342
rect 2967 338 2971 342
rect 2999 338 3003 342
rect 3095 338 3099 342
rect 3167 338 3171 342
rect 3239 338 3243 342
rect 3343 338 3347 342
rect 3383 338 3387 342
rect 3511 338 3515 342
rect 3591 338 3595 342
rect 111 262 115 266
rect 135 262 139 266
rect 271 262 275 266
rect 303 262 307 266
rect 391 262 395 266
rect 447 262 451 266
rect 495 262 499 266
rect 599 262 603 266
rect 631 262 635 266
rect 711 262 715 266
rect 815 262 819 266
rect 823 262 827 266
rect 943 262 947 266
rect 991 262 995 266
rect 1063 262 1067 266
rect 1159 262 1163 266
rect 1175 262 1179 266
rect 1287 262 1291 266
rect 1319 262 1323 266
rect 1407 262 1411 266
rect 1471 262 1475 266
rect 1527 262 1531 266
rect 1615 262 1619 266
rect 1647 262 1651 266
rect 1743 262 1747 266
rect 1831 262 1835 266
rect 1871 258 1875 262
rect 2023 258 2027 262
rect 2071 258 2075 262
rect 2111 258 2115 262
rect 2215 258 2219 262
rect 2319 258 2323 262
rect 2327 258 2331 262
rect 2439 258 2443 262
rect 2543 258 2547 262
rect 2559 258 2563 262
rect 2687 258 2691 262
rect 2743 258 2747 262
rect 2831 258 2835 262
rect 2927 258 2931 262
rect 2991 258 2995 262
rect 3087 258 3091 262
rect 3159 258 3163 262
rect 3239 258 3243 262
rect 3335 258 3339 262
rect 3383 258 3387 262
rect 3503 258 3507 262
rect 3591 258 3595 262
rect 111 162 115 166
rect 263 162 267 166
rect 311 162 315 166
rect 343 162 347 166
rect 399 162 403 166
rect 423 162 427 166
rect 503 162 507 166
rect 583 162 587 166
rect 607 162 611 166
rect 663 162 667 166
rect 719 162 723 166
rect 743 162 747 166
rect 823 162 827 166
rect 831 162 835 166
rect 903 162 907 166
rect 951 162 955 166
rect 983 162 987 166
rect 1063 162 1067 166
rect 1071 162 1075 166
rect 1143 162 1147 166
rect 1183 162 1187 166
rect 1223 162 1227 166
rect 1295 162 1299 166
rect 1303 162 1307 166
rect 1383 162 1387 166
rect 1415 162 1419 166
rect 1463 162 1467 166
rect 1535 162 1539 166
rect 1543 162 1547 166
rect 1655 162 1659 166
rect 1751 162 1755 166
rect 1831 162 1835 166
rect 1871 158 1875 162
rect 1903 158 1907 162
rect 1983 158 1987 162
rect 2063 158 2067 162
rect 2079 158 2083 162
rect 2143 158 2147 162
rect 2223 158 2227 162
rect 2303 158 2307 162
rect 2327 158 2331 162
rect 2399 158 2403 162
rect 2503 158 2507 162
rect 2551 158 2555 162
rect 2607 158 2611 162
rect 2711 158 2715 162
rect 2751 158 2755 162
rect 2815 158 2819 162
rect 2911 158 2915 162
rect 2935 158 2939 162
rect 2999 158 3003 162
rect 3087 158 3091 162
rect 3095 158 3099 162
rect 3175 158 3179 162
rect 3247 158 3251 162
rect 3263 158 3267 162
rect 3351 158 3355 162
rect 3391 158 3395 162
rect 3431 158 3435 162
rect 3511 158 3515 162
rect 3591 158 3595 162
rect 111 86 115 90
rect 255 86 259 90
rect 335 86 339 90
rect 415 86 419 90
rect 495 86 499 90
rect 575 86 579 90
rect 655 86 659 90
rect 735 86 739 90
rect 815 86 819 90
rect 895 86 899 90
rect 975 86 979 90
rect 1055 86 1059 90
rect 1135 86 1139 90
rect 1215 86 1219 90
rect 1295 86 1299 90
rect 1375 86 1379 90
rect 1455 86 1459 90
rect 1535 86 1539 90
rect 1831 86 1835 90
rect 1871 82 1875 86
rect 1895 82 1899 86
rect 1975 82 1979 86
rect 2055 82 2059 86
rect 2135 82 2139 86
rect 2215 82 2219 86
rect 2295 82 2299 86
rect 2391 82 2395 86
rect 2495 82 2499 86
rect 2599 82 2603 86
rect 2703 82 2707 86
rect 2807 82 2811 86
rect 2903 82 2907 86
rect 2991 82 2995 86
rect 3079 82 3083 86
rect 3167 82 3171 86
rect 3255 82 3259 86
rect 3343 82 3347 86
rect 3423 82 3427 86
rect 3503 82 3507 86
rect 3591 82 3595 86
<< m4 >>
rect 96 3653 97 3659
rect 103 3658 1855 3659
rect 103 3654 111 3658
rect 115 3654 143 3658
rect 147 3654 223 3658
rect 227 3654 351 3658
rect 355 3654 495 3658
rect 499 3654 647 3658
rect 651 3654 807 3658
rect 811 3654 975 3658
rect 979 3654 1151 3658
rect 1155 3654 1335 3658
rect 1339 3654 1831 3658
rect 1835 3654 1855 3658
rect 103 3653 1855 3654
rect 1861 3653 1862 3659
rect 1854 3625 1855 3631
rect 1861 3630 3631 3631
rect 1861 3626 1871 3630
rect 1875 3626 1927 3630
rect 1931 3626 2007 3630
rect 2011 3626 2103 3630
rect 2107 3626 2207 3630
rect 2211 3626 2319 3630
rect 2323 3626 2431 3630
rect 2435 3626 2551 3630
rect 2555 3626 2663 3630
rect 2667 3626 2775 3630
rect 2779 3626 2879 3630
rect 2883 3626 2983 3630
rect 2987 3626 3095 3630
rect 3099 3626 3207 3630
rect 3211 3626 3591 3630
rect 3595 3626 3631 3630
rect 1861 3625 3631 3626
rect 3637 3625 3638 3631
rect 84 3577 85 3583
rect 91 3582 1843 3583
rect 91 3578 111 3582
rect 115 3578 135 3582
rect 139 3578 215 3582
rect 219 3578 239 3582
rect 243 3578 343 3582
rect 347 3578 359 3582
rect 363 3578 479 3582
rect 483 3578 487 3582
rect 491 3578 607 3582
rect 611 3578 639 3582
rect 643 3578 735 3582
rect 739 3578 799 3582
rect 803 3578 863 3582
rect 867 3578 967 3582
rect 971 3578 983 3582
rect 987 3578 1095 3582
rect 1099 3578 1143 3582
rect 1147 3578 1207 3582
rect 1211 3578 1319 3582
rect 1323 3578 1327 3582
rect 1331 3578 1439 3582
rect 1443 3578 1831 3582
rect 1835 3578 1843 3582
rect 91 3577 1843 3578
rect 1849 3577 1850 3583
rect 1842 3549 1843 3555
rect 1849 3554 3619 3555
rect 1849 3550 1871 3554
rect 1875 3550 1919 3554
rect 1923 3550 1943 3554
rect 1947 3550 1999 3554
rect 2003 3550 2095 3554
rect 2099 3550 2127 3554
rect 2131 3550 2199 3554
rect 2203 3550 2303 3554
rect 2307 3550 2311 3554
rect 2315 3550 2423 3554
rect 2427 3550 2479 3554
rect 2483 3550 2543 3554
rect 2547 3550 2647 3554
rect 2651 3550 2655 3554
rect 2659 3550 2767 3554
rect 2771 3550 2815 3554
rect 2819 3550 2871 3554
rect 2875 3550 2975 3554
rect 2979 3550 3087 3554
rect 3091 3550 3135 3554
rect 3139 3550 3199 3554
rect 3203 3550 3303 3554
rect 3307 3550 3591 3554
rect 3595 3550 3619 3554
rect 1849 3549 3619 3550
rect 3625 3549 3626 3555
rect 96 3501 97 3507
rect 103 3506 1855 3507
rect 103 3502 111 3506
rect 115 3502 167 3506
rect 171 3502 247 3506
rect 251 3502 287 3506
rect 291 3502 367 3506
rect 371 3502 415 3506
rect 419 3502 487 3506
rect 491 3502 551 3506
rect 555 3502 615 3506
rect 619 3502 687 3506
rect 691 3502 743 3506
rect 747 3502 823 3506
rect 827 3502 871 3506
rect 875 3502 951 3506
rect 955 3502 991 3506
rect 995 3502 1071 3506
rect 1075 3502 1103 3506
rect 1107 3502 1183 3506
rect 1187 3502 1215 3506
rect 1219 3502 1303 3506
rect 1307 3502 1327 3506
rect 1331 3502 1423 3506
rect 1427 3502 1447 3506
rect 1451 3502 1831 3506
rect 1835 3502 1855 3506
rect 103 3501 1855 3502
rect 1861 3501 1862 3507
rect 1854 3473 1855 3479
rect 1861 3478 3631 3479
rect 1861 3474 1871 3478
rect 1875 3474 1951 3478
rect 1955 3474 1959 3478
rect 1963 3474 2079 3478
rect 2083 3474 2135 3478
rect 2139 3474 2199 3478
rect 2203 3474 2311 3478
rect 2315 3474 2335 3478
rect 2339 3474 2479 3478
rect 2483 3474 2487 3478
rect 2491 3474 2631 3478
rect 2635 3474 2655 3478
rect 2659 3474 2791 3478
rect 2795 3474 2823 3478
rect 2827 3474 2959 3478
rect 2963 3474 2983 3478
rect 2987 3474 3127 3478
rect 3131 3474 3143 3478
rect 3147 3474 3303 3478
rect 3307 3474 3311 3478
rect 3315 3474 3591 3478
rect 3595 3474 3631 3478
rect 1861 3473 3631 3474
rect 3637 3473 3638 3479
rect 84 3417 85 3423
rect 91 3422 1843 3423
rect 91 3418 111 3422
rect 115 3418 135 3422
rect 139 3418 159 3422
rect 163 3418 247 3422
rect 251 3418 279 3422
rect 283 3418 375 3422
rect 379 3418 407 3422
rect 411 3418 503 3422
rect 507 3418 543 3422
rect 547 3418 639 3422
rect 643 3418 679 3422
rect 683 3418 775 3422
rect 779 3418 815 3422
rect 819 3418 903 3422
rect 907 3418 943 3422
rect 947 3418 1031 3422
rect 1035 3418 1063 3422
rect 1067 3418 1159 3422
rect 1163 3418 1175 3422
rect 1179 3418 1287 3422
rect 1291 3418 1295 3422
rect 1299 3418 1415 3422
rect 1419 3418 1831 3422
rect 1835 3418 1843 3422
rect 91 3417 1843 3418
rect 1849 3417 1850 3423
rect 1842 3389 1843 3395
rect 1849 3394 3619 3395
rect 1849 3390 1871 3394
rect 1875 3390 1951 3394
rect 1955 3390 1975 3394
rect 1979 3390 2071 3394
rect 2075 3390 2135 3394
rect 2139 3390 2191 3394
rect 2195 3390 2287 3394
rect 2291 3390 2327 3394
rect 2331 3390 2431 3394
rect 2435 3390 2471 3394
rect 2475 3390 2559 3394
rect 2563 3390 2623 3394
rect 2627 3390 2679 3394
rect 2683 3390 2783 3394
rect 2787 3390 2791 3394
rect 2795 3390 2895 3394
rect 2899 3390 2951 3394
rect 2955 3390 2991 3394
rect 2995 3390 3079 3394
rect 3083 3390 3119 3394
rect 3123 3390 3167 3394
rect 3171 3390 3255 3394
rect 3259 3390 3295 3394
rect 3299 3390 3343 3394
rect 3347 3390 3423 3394
rect 3427 3390 3503 3394
rect 3507 3390 3591 3394
rect 3595 3390 3619 3394
rect 1849 3389 3619 3390
rect 3625 3389 3626 3395
rect 96 3337 97 3343
rect 103 3342 1855 3343
rect 103 3338 111 3342
rect 115 3338 143 3342
rect 147 3338 255 3342
rect 259 3338 271 3342
rect 275 3338 383 3342
rect 387 3338 391 3342
rect 395 3338 511 3342
rect 515 3338 519 3342
rect 523 3338 647 3342
rect 651 3338 655 3342
rect 659 3338 783 3342
rect 787 3338 791 3342
rect 795 3338 911 3342
rect 915 3338 919 3342
rect 923 3338 1039 3342
rect 1043 3338 1055 3342
rect 1059 3338 1167 3342
rect 1171 3338 1191 3342
rect 1195 3338 1295 3342
rect 1299 3338 1327 3342
rect 1331 3338 1423 3342
rect 1427 3338 1463 3342
rect 1467 3338 1831 3342
rect 1835 3338 1855 3342
rect 103 3337 1855 3338
rect 1861 3337 1862 3343
rect 1854 3309 1855 3315
rect 1861 3314 3631 3315
rect 1861 3310 1871 3314
rect 1875 3310 1935 3314
rect 1939 3310 1983 3314
rect 1987 3310 2071 3314
rect 2075 3310 2143 3314
rect 2147 3310 2207 3314
rect 2211 3310 2295 3314
rect 2299 3310 2367 3314
rect 2371 3310 2439 3314
rect 2443 3310 2551 3314
rect 2555 3310 2567 3314
rect 2571 3310 2687 3314
rect 2691 3310 2767 3314
rect 2771 3310 2799 3314
rect 2803 3310 2903 3314
rect 2907 3310 2999 3314
rect 3003 3310 3007 3314
rect 3011 3310 3087 3314
rect 3091 3310 3175 3314
rect 3179 3310 3255 3314
rect 3259 3310 3263 3314
rect 3267 3310 3351 3314
rect 3355 3310 3431 3314
rect 3435 3310 3511 3314
rect 3515 3310 3591 3314
rect 3595 3310 3631 3314
rect 1861 3309 3631 3310
rect 3637 3309 3638 3315
rect 84 3257 85 3263
rect 91 3262 1843 3263
rect 91 3258 111 3262
rect 115 3258 263 3262
rect 267 3258 383 3262
rect 387 3258 471 3262
rect 475 3258 511 3262
rect 515 3258 575 3262
rect 579 3258 647 3262
rect 651 3258 687 3262
rect 691 3258 783 3262
rect 787 3258 807 3262
rect 811 3258 911 3262
rect 915 3258 935 3262
rect 939 3258 1047 3262
rect 1051 3258 1063 3262
rect 1067 3258 1183 3262
rect 1187 3258 1191 3262
rect 1195 3258 1319 3262
rect 1323 3258 1447 3262
rect 1451 3258 1455 3262
rect 1459 3258 1575 3262
rect 1579 3258 1831 3262
rect 1835 3258 1843 3262
rect 91 3257 1843 3258
rect 1849 3257 1850 3263
rect 1842 3229 1843 3235
rect 1849 3234 3619 3235
rect 1849 3230 1871 3234
rect 1875 3230 1895 3234
rect 1899 3230 1927 3234
rect 1931 3230 2007 3234
rect 2011 3230 2063 3234
rect 2067 3230 2143 3234
rect 2147 3230 2199 3234
rect 2203 3230 2279 3234
rect 2283 3230 2359 3234
rect 2363 3230 2415 3234
rect 2419 3230 2543 3234
rect 2547 3230 2567 3234
rect 2571 3230 2727 3234
rect 2731 3230 2759 3234
rect 2763 3230 2911 3234
rect 2915 3230 2999 3234
rect 3003 3230 3103 3234
rect 3107 3230 3247 3234
rect 3251 3230 3311 3234
rect 3315 3230 3503 3234
rect 3507 3230 3591 3234
rect 3595 3230 3619 3234
rect 1849 3229 3619 3230
rect 3625 3229 3626 3235
rect 96 3173 97 3179
rect 103 3178 1855 3179
rect 103 3174 111 3178
rect 115 3174 383 3178
rect 387 3174 391 3178
rect 395 3174 463 3178
rect 467 3174 479 3178
rect 483 3174 543 3178
rect 547 3174 583 3178
rect 587 3174 623 3178
rect 627 3174 695 3178
rect 699 3174 711 3178
rect 715 3174 815 3178
rect 819 3174 927 3178
rect 931 3174 943 3178
rect 947 3174 1039 3178
rect 1043 3174 1071 3178
rect 1075 3174 1159 3178
rect 1163 3174 1199 3178
rect 1203 3174 1271 3178
rect 1275 3174 1327 3178
rect 1331 3174 1383 3178
rect 1387 3174 1455 3178
rect 1459 3174 1495 3178
rect 1499 3174 1583 3178
rect 1587 3174 1615 3178
rect 1619 3174 1735 3178
rect 1739 3174 1831 3178
rect 1835 3174 1855 3178
rect 103 3173 1855 3174
rect 1861 3173 1862 3179
rect 1854 3153 1855 3159
rect 1861 3158 3631 3159
rect 1861 3154 1871 3158
rect 1875 3154 1903 3158
rect 1907 3154 2015 3158
rect 2019 3154 2079 3158
rect 2083 3154 2151 3158
rect 2155 3154 2271 3158
rect 2275 3154 2287 3158
rect 2291 3154 2423 3158
rect 2427 3154 2455 3158
rect 2459 3154 2575 3158
rect 2579 3154 2623 3158
rect 2627 3154 2735 3158
rect 2739 3154 2783 3158
rect 2787 3154 2919 3158
rect 2923 3154 2935 3158
rect 2939 3154 3079 3158
rect 3083 3154 3111 3158
rect 3115 3154 3231 3158
rect 3235 3154 3319 3158
rect 3323 3154 3511 3158
rect 3515 3154 3591 3158
rect 3595 3154 3631 3158
rect 1861 3153 3631 3154
rect 3637 3153 3638 3159
rect 84 3097 85 3103
rect 91 3102 1843 3103
rect 91 3098 111 3102
rect 115 3098 375 3102
rect 379 3098 455 3102
rect 459 3098 535 3102
rect 539 3098 615 3102
rect 619 3098 703 3102
rect 707 3098 807 3102
rect 811 3098 919 3102
rect 923 3098 943 3102
rect 947 3098 1023 3102
rect 1027 3098 1031 3102
rect 1035 3098 1103 3102
rect 1107 3098 1151 3102
rect 1155 3098 1183 3102
rect 1187 3098 1263 3102
rect 1267 3098 1343 3102
rect 1347 3098 1375 3102
rect 1379 3098 1423 3102
rect 1427 3098 1487 3102
rect 1491 3098 1503 3102
rect 1507 3098 1583 3102
rect 1587 3098 1607 3102
rect 1611 3098 1663 3102
rect 1667 3098 1727 3102
rect 1731 3098 1743 3102
rect 1747 3098 1831 3102
rect 1835 3098 1843 3102
rect 91 3097 1843 3098
rect 1849 3097 1850 3103
rect 1842 3069 1843 3075
rect 1849 3074 3619 3075
rect 1849 3070 1871 3074
rect 1875 3070 1895 3074
rect 1899 3070 1991 3074
rect 1995 3070 2071 3074
rect 2075 3070 2247 3074
rect 2251 3070 2263 3074
rect 2267 3070 2447 3074
rect 2451 3070 2487 3074
rect 2491 3070 2615 3074
rect 2619 3070 2703 3074
rect 2707 3070 2775 3074
rect 2779 3070 2895 3074
rect 2899 3070 2927 3074
rect 2931 3070 3063 3074
rect 3067 3070 3071 3074
rect 3075 3070 3223 3074
rect 3227 3070 3375 3074
rect 3379 3070 3503 3074
rect 3507 3070 3591 3074
rect 3595 3070 3619 3074
rect 1849 3069 3619 3070
rect 3625 3069 3626 3075
rect 96 3005 97 3011
rect 103 3010 1855 3011
rect 103 3006 111 3010
rect 115 3006 207 3010
rect 211 3006 327 3010
rect 331 3006 471 3010
rect 475 3006 631 3010
rect 635 3006 807 3010
rect 811 3006 951 3010
rect 955 3006 983 3010
rect 987 3006 1031 3010
rect 1035 3006 1111 3010
rect 1115 3006 1151 3010
rect 1155 3006 1191 3010
rect 1195 3006 1271 3010
rect 1275 3006 1311 3010
rect 1315 3006 1351 3010
rect 1355 3006 1431 3010
rect 1435 3006 1463 3010
rect 1467 3006 1511 3010
rect 1515 3006 1591 3010
rect 1595 3006 1615 3010
rect 1619 3006 1671 3010
rect 1675 3006 1751 3010
rect 1755 3006 1831 3010
rect 1835 3006 1855 3010
rect 103 3005 1855 3006
rect 1861 3005 1862 3011
rect 1854 2989 1855 2995
rect 1861 2994 3631 2995
rect 1861 2990 1871 2994
rect 1875 2990 1903 2994
rect 1907 2990 1999 2994
rect 2003 2990 2143 2994
rect 2147 2990 2255 2994
rect 2259 2990 2391 2994
rect 2395 2990 2495 2994
rect 2499 2990 2607 2994
rect 2611 2990 2711 2994
rect 2715 2990 2799 2994
rect 2803 2990 2903 2994
rect 2907 2990 2967 2994
rect 2971 2990 3071 2994
rect 3075 2990 3119 2994
rect 3123 2990 3231 2994
rect 3235 2990 3263 2994
rect 3267 2990 3383 2994
rect 3387 2990 3399 2994
rect 3403 2990 3511 2994
rect 3515 2990 3591 2994
rect 3595 2990 3631 2994
rect 1861 2989 3631 2990
rect 3637 2989 3638 2995
rect 84 2929 85 2935
rect 91 2934 1843 2935
rect 91 2930 111 2934
rect 115 2930 199 2934
rect 203 2930 247 2934
rect 251 2930 319 2934
rect 323 2930 351 2934
rect 355 2930 463 2934
rect 467 2930 471 2934
rect 475 2930 607 2934
rect 611 2930 623 2934
rect 627 2930 751 2934
rect 755 2930 799 2934
rect 803 2930 895 2934
rect 899 2930 975 2934
rect 979 2930 1031 2934
rect 1035 2930 1143 2934
rect 1147 2930 1159 2934
rect 1163 2930 1279 2934
rect 1283 2930 1303 2934
rect 1307 2930 1399 2934
rect 1403 2930 1455 2934
rect 1459 2930 1519 2934
rect 1523 2930 1607 2934
rect 1611 2930 1639 2934
rect 1643 2930 1743 2934
rect 1747 2930 1831 2934
rect 1835 2930 1843 2934
rect 91 2929 1843 2930
rect 1849 2929 1850 2935
rect 1842 2901 1843 2907
rect 1849 2906 3619 2907
rect 1849 2902 1871 2906
rect 1875 2902 1895 2906
rect 1899 2902 2135 2906
rect 2139 2902 2351 2906
rect 2355 2902 2383 2906
rect 2387 2902 2447 2906
rect 2451 2902 2551 2906
rect 2555 2902 2599 2906
rect 2603 2902 2655 2906
rect 2659 2902 2759 2906
rect 2763 2902 2791 2906
rect 2795 2902 2871 2906
rect 2875 2902 2959 2906
rect 2963 2902 2983 2906
rect 2987 2902 3095 2906
rect 3099 2902 3111 2906
rect 3115 2902 3207 2906
rect 3211 2902 3255 2906
rect 3259 2902 3391 2906
rect 3395 2902 3503 2906
rect 3507 2902 3591 2906
rect 3595 2902 3619 2906
rect 1849 2901 3619 2902
rect 3625 2901 3626 2907
rect 96 2853 97 2859
rect 103 2858 1855 2859
rect 103 2854 111 2858
rect 115 2854 151 2858
rect 155 2854 255 2858
rect 259 2854 279 2858
rect 283 2854 359 2858
rect 363 2854 407 2858
rect 411 2854 479 2858
rect 483 2854 543 2858
rect 547 2854 615 2858
rect 619 2854 671 2858
rect 675 2854 759 2858
rect 763 2854 799 2858
rect 803 2854 903 2858
rect 907 2854 919 2858
rect 923 2854 1039 2858
rect 1043 2854 1151 2858
rect 1155 2854 1167 2858
rect 1171 2854 1271 2858
rect 1275 2854 1287 2858
rect 1291 2854 1391 2858
rect 1395 2854 1407 2858
rect 1411 2854 1527 2858
rect 1531 2854 1647 2858
rect 1651 2854 1831 2858
rect 1835 2854 1855 2858
rect 103 2853 1855 2854
rect 1861 2853 1862 2859
rect 1854 2825 1855 2831
rect 1861 2830 3631 2831
rect 1861 2826 1871 2830
rect 1875 2826 2239 2830
rect 2243 2826 2319 2830
rect 2323 2826 2359 2830
rect 2363 2826 2399 2830
rect 2403 2826 2455 2830
rect 2459 2826 2479 2830
rect 2483 2826 2559 2830
rect 2563 2826 2567 2830
rect 2571 2826 2663 2830
rect 2667 2826 2671 2830
rect 2675 2826 2767 2830
rect 2771 2826 2807 2830
rect 2811 2826 2879 2830
rect 2883 2826 2967 2830
rect 2971 2826 2991 2830
rect 2995 2826 3103 2830
rect 3107 2826 3143 2830
rect 3147 2826 3215 2830
rect 3219 2826 3335 2830
rect 3339 2826 3511 2830
rect 3515 2826 3591 2830
rect 3595 2826 3631 2830
rect 1861 2825 3631 2826
rect 3637 2825 3638 2831
rect 84 2769 85 2775
rect 91 2774 1843 2775
rect 91 2770 111 2774
rect 115 2770 143 2774
rect 147 2770 271 2774
rect 275 2770 295 2774
rect 299 2770 399 2774
rect 403 2770 439 2774
rect 443 2770 535 2774
rect 539 2770 567 2774
rect 571 2770 663 2774
rect 667 2770 687 2774
rect 691 2770 791 2774
rect 795 2770 799 2774
rect 803 2770 903 2774
rect 907 2770 911 2774
rect 915 2770 1007 2774
rect 1011 2770 1031 2774
rect 1035 2770 1103 2774
rect 1107 2770 1143 2774
rect 1147 2770 1199 2774
rect 1203 2770 1263 2774
rect 1267 2770 1303 2774
rect 1307 2770 1383 2774
rect 1387 2770 1831 2774
rect 1835 2770 1843 2774
rect 91 2769 1843 2770
rect 1849 2769 1850 2775
rect 1842 2737 1843 2743
rect 1849 2742 3619 2743
rect 1849 2738 1871 2742
rect 1875 2738 2047 2742
rect 2051 2738 2135 2742
rect 2139 2738 2231 2742
rect 2235 2738 2311 2742
rect 2315 2738 2327 2742
rect 2331 2738 2391 2742
rect 2395 2738 2423 2742
rect 2427 2738 2471 2742
rect 2475 2738 2519 2742
rect 2523 2738 2559 2742
rect 2563 2738 2615 2742
rect 2619 2738 2663 2742
rect 2667 2738 2727 2742
rect 2731 2738 2799 2742
rect 2803 2738 2855 2742
rect 2859 2738 2959 2742
rect 2963 2738 3007 2742
rect 3011 2738 3135 2742
rect 3139 2738 3175 2742
rect 3179 2738 3327 2742
rect 3331 2738 3351 2742
rect 3355 2738 3503 2742
rect 3507 2738 3591 2742
rect 3595 2738 3619 2742
rect 1849 2737 3619 2738
rect 3625 2737 3626 2743
rect 96 2689 97 2695
rect 103 2694 1855 2695
rect 103 2690 111 2694
rect 115 2690 143 2694
rect 147 2690 151 2694
rect 155 2690 263 2694
rect 267 2690 303 2694
rect 307 2690 407 2694
rect 411 2690 447 2694
rect 451 2690 543 2694
rect 547 2690 575 2694
rect 579 2690 671 2694
rect 675 2690 695 2694
rect 699 2690 791 2694
rect 795 2690 807 2694
rect 811 2690 903 2694
rect 907 2690 911 2694
rect 915 2690 1015 2694
rect 1019 2690 1111 2694
rect 1115 2690 1119 2694
rect 1123 2690 1207 2694
rect 1211 2690 1215 2694
rect 1219 2690 1311 2694
rect 1315 2690 1319 2694
rect 1323 2690 1423 2694
rect 1427 2690 1831 2694
rect 1835 2690 1855 2694
rect 103 2689 1855 2690
rect 1861 2689 1862 2695
rect 1854 2661 1855 2667
rect 1861 2666 3631 2667
rect 1861 2662 1871 2666
rect 1875 2662 2055 2666
rect 2059 2662 2071 2666
rect 2075 2662 2143 2666
rect 2147 2662 2239 2666
rect 2243 2662 2295 2666
rect 2299 2662 2335 2666
rect 2339 2662 2431 2666
rect 2435 2662 2527 2666
rect 2531 2662 2567 2666
rect 2571 2662 2623 2666
rect 2627 2662 2735 2666
rect 2739 2662 2863 2666
rect 2867 2662 2871 2666
rect 2875 2662 3015 2666
rect 3019 2662 3183 2666
rect 3187 2662 3199 2666
rect 3203 2662 3359 2666
rect 3363 2662 3511 2666
rect 3515 2662 3591 2666
rect 3595 2662 3631 2666
rect 1861 2661 3631 2662
rect 3637 2661 3638 2667
rect 84 2605 85 2611
rect 91 2610 1843 2611
rect 91 2606 111 2610
rect 115 2606 135 2610
rect 139 2606 143 2610
rect 147 2606 255 2610
rect 259 2606 311 2610
rect 315 2606 399 2610
rect 403 2606 479 2610
rect 483 2606 535 2610
rect 539 2606 639 2610
rect 643 2606 663 2610
rect 667 2606 783 2610
rect 787 2606 791 2610
rect 795 2606 895 2610
rect 899 2606 927 2610
rect 931 2606 1007 2610
rect 1011 2606 1055 2610
rect 1059 2606 1111 2610
rect 1115 2606 1175 2610
rect 1179 2606 1207 2610
rect 1211 2606 1295 2610
rect 1299 2606 1311 2610
rect 1315 2606 1407 2610
rect 1411 2606 1415 2610
rect 1419 2606 1527 2610
rect 1531 2606 1831 2610
rect 1835 2606 1843 2610
rect 91 2605 1843 2606
rect 1849 2605 1850 2611
rect 1842 2581 1843 2587
rect 1849 2586 3619 2587
rect 1849 2582 1871 2586
rect 1875 2582 2063 2586
rect 2067 2582 2167 2586
rect 2171 2582 2263 2586
rect 2267 2582 2287 2586
rect 2291 2582 2367 2586
rect 2371 2582 2479 2586
rect 2483 2582 2559 2586
rect 2563 2582 2591 2586
rect 2595 2582 2695 2586
rect 2699 2582 2799 2586
rect 2803 2582 2863 2586
rect 2867 2582 2903 2586
rect 2907 2582 3015 2586
rect 3019 2582 3135 2586
rect 3139 2582 3191 2586
rect 3195 2582 3263 2586
rect 3267 2582 3391 2586
rect 3395 2582 3503 2586
rect 3507 2582 3591 2586
rect 3595 2582 3619 2586
rect 1849 2581 3619 2582
rect 3625 2581 3626 2587
rect 96 2521 97 2527
rect 103 2526 1855 2527
rect 103 2522 111 2526
rect 115 2522 143 2526
rect 147 2522 151 2526
rect 155 2522 295 2526
rect 299 2522 319 2526
rect 323 2522 447 2526
rect 451 2522 487 2526
rect 491 2522 591 2526
rect 595 2522 647 2526
rect 651 2522 735 2526
rect 739 2522 799 2526
rect 803 2522 879 2526
rect 883 2522 935 2526
rect 939 2522 1015 2526
rect 1019 2522 1063 2526
rect 1067 2522 1143 2526
rect 1147 2522 1183 2526
rect 1187 2522 1271 2526
rect 1275 2522 1303 2526
rect 1307 2522 1399 2526
rect 1403 2522 1415 2526
rect 1419 2522 1535 2526
rect 1539 2522 1831 2526
rect 1835 2522 1855 2526
rect 103 2521 1855 2522
rect 1861 2521 1862 2527
rect 1854 2505 1855 2511
rect 1861 2510 3631 2511
rect 1861 2506 1871 2510
rect 1875 2506 2135 2510
rect 2139 2506 2175 2510
rect 2179 2506 2223 2510
rect 2227 2506 2271 2510
rect 2275 2506 2319 2510
rect 2323 2506 2375 2510
rect 2379 2506 2423 2510
rect 2427 2506 2487 2510
rect 2491 2506 2535 2510
rect 2539 2506 2599 2510
rect 2603 2506 2655 2510
rect 2659 2506 2703 2510
rect 2707 2506 2783 2510
rect 2787 2506 2807 2510
rect 2811 2506 2911 2510
rect 2915 2506 2919 2510
rect 2923 2506 3023 2510
rect 3027 2506 3063 2510
rect 3067 2506 3143 2510
rect 3147 2506 3215 2510
rect 3219 2506 3271 2510
rect 3275 2506 3375 2510
rect 3379 2506 3399 2510
rect 3403 2506 3511 2510
rect 3515 2506 3591 2510
rect 3595 2506 3631 2510
rect 1861 2505 3631 2506
rect 3637 2505 3638 2511
rect 84 2441 85 2447
rect 91 2446 1843 2447
rect 91 2442 111 2446
rect 115 2442 135 2446
rect 139 2442 199 2446
rect 203 2442 287 2446
rect 291 2442 351 2446
rect 355 2442 439 2446
rect 443 2442 495 2446
rect 499 2442 583 2446
rect 587 2442 639 2446
rect 643 2442 727 2446
rect 731 2442 783 2446
rect 787 2442 871 2446
rect 875 2442 919 2446
rect 923 2442 1007 2446
rect 1011 2442 1047 2446
rect 1051 2442 1135 2446
rect 1139 2442 1175 2446
rect 1179 2442 1263 2446
rect 1267 2442 1311 2446
rect 1315 2442 1391 2446
rect 1395 2442 1447 2446
rect 1451 2442 1527 2446
rect 1531 2442 1831 2446
rect 1835 2442 1843 2446
rect 91 2441 1843 2442
rect 1849 2441 1850 2447
rect 1842 2421 1843 2427
rect 1849 2426 3619 2427
rect 1849 2422 1871 2426
rect 1875 2422 1975 2426
rect 1979 2422 2087 2426
rect 2091 2422 2127 2426
rect 2131 2422 2207 2426
rect 2211 2422 2215 2426
rect 2219 2422 2311 2426
rect 2315 2422 2335 2426
rect 2339 2422 2415 2426
rect 2419 2422 2479 2426
rect 2483 2422 2527 2426
rect 2531 2422 2631 2426
rect 2635 2422 2647 2426
rect 2651 2422 2775 2426
rect 2779 2422 2791 2426
rect 2795 2422 2911 2426
rect 2915 2422 2967 2426
rect 2971 2422 3055 2426
rect 3059 2422 3151 2426
rect 3155 2422 3207 2426
rect 3211 2422 3335 2426
rect 3339 2422 3367 2426
rect 3371 2422 3503 2426
rect 3507 2422 3591 2426
rect 3595 2422 3619 2426
rect 1849 2421 3619 2422
rect 3625 2421 3626 2427
rect 96 2357 97 2363
rect 103 2362 1855 2363
rect 103 2358 111 2362
rect 115 2358 207 2362
rect 211 2358 223 2362
rect 227 2358 327 2362
rect 331 2358 359 2362
rect 363 2358 439 2362
rect 443 2358 503 2362
rect 507 2358 559 2362
rect 563 2358 647 2362
rect 651 2358 679 2362
rect 683 2358 791 2362
rect 795 2358 799 2362
rect 803 2358 911 2362
rect 915 2358 927 2362
rect 931 2358 1023 2362
rect 1027 2358 1055 2362
rect 1059 2358 1135 2362
rect 1139 2358 1183 2362
rect 1187 2358 1247 2362
rect 1251 2358 1319 2362
rect 1323 2358 1367 2362
rect 1371 2358 1455 2362
rect 1459 2358 1831 2362
rect 1835 2358 1855 2362
rect 103 2357 1855 2358
rect 1861 2357 1862 2363
rect 1854 2341 1855 2347
rect 1861 2346 3631 2347
rect 1861 2342 1871 2346
rect 1875 2342 1903 2346
rect 1907 2342 1983 2346
rect 1987 2342 2015 2346
rect 2019 2342 2095 2346
rect 2099 2342 2167 2346
rect 2171 2342 2215 2346
rect 2219 2342 2319 2346
rect 2323 2342 2343 2346
rect 2347 2342 2471 2346
rect 2475 2342 2487 2346
rect 2491 2342 2623 2346
rect 2627 2342 2639 2346
rect 2643 2342 2775 2346
rect 2779 2342 2799 2346
rect 2803 2342 2927 2346
rect 2931 2342 2975 2346
rect 2979 2342 3087 2346
rect 3091 2342 3159 2346
rect 3163 2342 3247 2346
rect 3251 2342 3343 2346
rect 3347 2342 3415 2346
rect 3419 2342 3511 2346
rect 3515 2342 3591 2346
rect 3595 2342 3631 2346
rect 1861 2341 3631 2342
rect 3637 2341 3638 2347
rect 84 2269 85 2275
rect 91 2274 1843 2275
rect 91 2270 111 2274
rect 115 2270 215 2274
rect 219 2270 311 2274
rect 315 2270 319 2274
rect 323 2270 407 2274
rect 411 2270 431 2274
rect 435 2270 503 2274
rect 507 2270 551 2274
rect 555 2270 607 2274
rect 611 2270 671 2274
rect 675 2270 711 2274
rect 715 2270 791 2274
rect 795 2270 815 2274
rect 819 2270 903 2274
rect 907 2270 911 2274
rect 915 2270 1007 2274
rect 1011 2270 1015 2274
rect 1019 2270 1103 2274
rect 1107 2270 1127 2274
rect 1131 2270 1199 2274
rect 1203 2270 1239 2274
rect 1243 2270 1303 2274
rect 1307 2270 1359 2274
rect 1363 2270 1831 2274
rect 1835 2270 1843 2274
rect 91 2269 1843 2270
rect 1849 2271 1850 2275
rect 1849 2270 3626 2271
rect 1849 2269 1871 2270
rect 1842 2266 1871 2269
rect 1875 2266 1895 2270
rect 1899 2266 2007 2270
rect 2011 2266 2031 2270
rect 2035 2266 2159 2270
rect 2163 2266 2207 2270
rect 2211 2266 2311 2270
rect 2315 2266 2391 2270
rect 2395 2266 2463 2270
rect 2467 2266 2575 2270
rect 2579 2266 2615 2270
rect 2619 2266 2767 2270
rect 2771 2266 2919 2270
rect 2923 2266 2951 2270
rect 2955 2266 3079 2270
rect 3083 2266 3143 2270
rect 3147 2266 3239 2270
rect 3243 2266 3335 2270
rect 3339 2266 3407 2270
rect 3411 2266 3503 2270
rect 3507 2266 3591 2270
rect 3595 2266 3626 2270
rect 1842 2265 3626 2266
rect 96 2189 97 2195
rect 103 2194 1855 2195
rect 103 2190 111 2194
rect 115 2190 319 2194
rect 323 2190 415 2194
rect 419 2190 511 2194
rect 515 2190 519 2194
rect 523 2190 615 2194
rect 619 2190 623 2194
rect 627 2190 719 2194
rect 723 2190 727 2194
rect 731 2190 823 2194
rect 827 2190 831 2194
rect 835 2190 919 2194
rect 923 2190 935 2194
rect 939 2190 1015 2194
rect 1019 2190 1039 2194
rect 1043 2190 1111 2194
rect 1115 2190 1151 2194
rect 1155 2190 1207 2194
rect 1211 2190 1263 2194
rect 1267 2190 1311 2194
rect 1315 2190 1831 2194
rect 1835 2190 1855 2194
rect 103 2189 1855 2190
rect 1861 2189 1862 2195
rect 1854 2187 1862 2189
rect 1854 2181 1855 2187
rect 1861 2186 3631 2187
rect 1861 2182 1871 2186
rect 1875 2182 1903 2186
rect 1907 2182 1967 2186
rect 1971 2182 2039 2186
rect 2043 2182 2079 2186
rect 2083 2182 2215 2186
rect 2219 2182 2367 2186
rect 2371 2182 2399 2186
rect 2403 2182 2527 2186
rect 2531 2182 2583 2186
rect 2587 2182 2687 2186
rect 2691 2182 2775 2186
rect 2779 2182 2847 2186
rect 2851 2182 2959 2186
rect 2963 2182 2991 2186
rect 2995 2182 3127 2186
rect 3131 2182 3151 2186
rect 3155 2182 3263 2186
rect 3267 2182 3343 2186
rect 3347 2182 3399 2186
rect 3403 2182 3511 2186
rect 3515 2182 3591 2186
rect 3595 2182 3631 2186
rect 1861 2181 3631 2182
rect 3637 2181 3638 2187
rect 84 2113 85 2119
rect 91 2118 1843 2119
rect 91 2114 111 2118
rect 115 2114 279 2118
rect 283 2114 311 2118
rect 315 2114 399 2118
rect 403 2114 407 2118
rect 411 2114 511 2118
rect 515 2114 615 2118
rect 619 2114 623 2118
rect 627 2114 719 2118
rect 723 2114 735 2118
rect 739 2114 823 2118
rect 827 2114 847 2118
rect 851 2114 927 2118
rect 931 2114 951 2118
rect 955 2114 1031 2118
rect 1035 2114 1047 2118
rect 1051 2114 1143 2118
rect 1147 2114 1239 2118
rect 1243 2114 1255 2118
rect 1259 2114 1343 2118
rect 1347 2114 1831 2118
rect 1835 2114 1843 2118
rect 91 2113 1843 2114
rect 1849 2113 1850 2119
rect 1842 2111 1850 2113
rect 1842 2105 1843 2111
rect 1849 2110 3619 2111
rect 1849 2106 1871 2110
rect 1875 2106 1959 2110
rect 1963 2106 2071 2110
rect 2075 2106 2207 2110
rect 2211 2106 2287 2110
rect 2291 2106 2359 2110
rect 2363 2106 2391 2110
rect 2395 2106 2503 2110
rect 2507 2106 2519 2110
rect 2523 2106 2623 2110
rect 2627 2106 2679 2110
rect 2683 2106 2743 2110
rect 2747 2106 2839 2110
rect 2843 2106 2855 2110
rect 2859 2106 2967 2110
rect 2971 2106 2983 2110
rect 2987 2106 3079 2110
rect 3083 2106 3119 2110
rect 3123 2106 3191 2110
rect 3195 2106 3255 2110
rect 3259 2106 3303 2110
rect 3307 2106 3391 2110
rect 3395 2106 3415 2110
rect 3419 2106 3503 2110
rect 3507 2106 3591 2110
rect 3595 2106 3619 2110
rect 1849 2105 3619 2106
rect 3625 2105 3626 2111
rect 96 2029 97 2035
rect 103 2034 1855 2035
rect 103 2030 111 2034
rect 115 2030 183 2034
rect 187 2030 287 2034
rect 291 2030 327 2034
rect 331 2030 407 2034
rect 411 2030 471 2034
rect 475 2030 519 2034
rect 523 2030 623 2034
rect 627 2030 631 2034
rect 635 2030 743 2034
rect 747 2030 767 2034
rect 771 2030 855 2034
rect 859 2030 911 2034
rect 915 2030 959 2034
rect 963 2030 1047 2034
rect 1051 2030 1055 2034
rect 1059 2030 1151 2034
rect 1155 2030 1183 2034
rect 1187 2030 1247 2034
rect 1251 2030 1319 2034
rect 1323 2030 1351 2034
rect 1355 2030 1463 2034
rect 1467 2030 1831 2034
rect 1835 2030 1855 2034
rect 103 2029 1855 2030
rect 1861 2031 1862 2035
rect 1861 2030 3638 2031
rect 1861 2029 1871 2030
rect 1854 2026 1871 2029
rect 1875 2026 2183 2030
rect 2187 2026 2271 2030
rect 2275 2026 2295 2030
rect 2299 2026 2367 2030
rect 2371 2026 2399 2030
rect 2403 2026 2463 2030
rect 2467 2026 2511 2030
rect 2515 2026 2567 2030
rect 2571 2026 2631 2030
rect 2635 2026 2671 2030
rect 2675 2026 2751 2030
rect 2755 2026 2775 2030
rect 2779 2026 2863 2030
rect 2867 2026 2879 2030
rect 2883 2026 2975 2030
rect 2979 2026 2983 2030
rect 2987 2026 3087 2030
rect 3091 2026 3191 2030
rect 3195 2026 3199 2030
rect 3203 2026 3311 2030
rect 3315 2026 3423 2030
rect 3427 2026 3511 2030
rect 3515 2026 3591 2030
rect 3595 2026 3638 2030
rect 1854 2025 3638 2026
rect 84 1953 85 1959
rect 91 1958 1843 1959
rect 91 1954 111 1958
rect 115 1954 135 1958
rect 139 1954 175 1958
rect 179 1954 295 1958
rect 299 1954 319 1958
rect 323 1954 463 1958
rect 467 1954 615 1958
rect 619 1954 631 1958
rect 635 1954 759 1958
rect 763 1954 799 1958
rect 803 1954 903 1958
rect 907 1954 951 1958
rect 955 1954 1039 1958
rect 1043 1954 1095 1958
rect 1099 1954 1175 1958
rect 1179 1954 1231 1958
rect 1235 1954 1311 1958
rect 1315 1954 1359 1958
rect 1363 1954 1455 1958
rect 1459 1954 1487 1958
rect 1491 1954 1623 1958
rect 1627 1954 1831 1958
rect 1835 1954 1843 1958
rect 91 1953 1843 1954
rect 1849 1953 1850 1959
rect 1842 1951 1850 1953
rect 1842 1945 1843 1951
rect 1849 1950 3619 1951
rect 1849 1946 1871 1950
rect 1875 1946 1943 1950
rect 1947 1946 2055 1950
rect 2059 1946 2167 1950
rect 2171 1946 2175 1950
rect 2179 1946 2263 1950
rect 2267 1946 2287 1950
rect 2291 1946 2359 1950
rect 2363 1946 2407 1950
rect 2411 1946 2455 1950
rect 2459 1946 2527 1950
rect 2531 1946 2559 1950
rect 2563 1946 2647 1950
rect 2651 1946 2663 1950
rect 2667 1946 2767 1950
rect 2771 1946 2775 1950
rect 2779 1946 2871 1950
rect 2875 1946 2911 1950
rect 2915 1946 2975 1950
rect 2979 1946 3055 1950
rect 3059 1946 3079 1950
rect 3083 1946 3183 1950
rect 3187 1946 3207 1950
rect 3211 1946 3367 1950
rect 3371 1946 3503 1950
rect 3507 1946 3591 1950
rect 3595 1946 3619 1950
rect 1849 1945 3619 1946
rect 3625 1945 3626 1951
rect 96 1869 97 1875
rect 103 1874 1855 1875
rect 103 1870 111 1874
rect 115 1870 143 1874
rect 147 1870 303 1874
rect 307 1870 319 1874
rect 323 1870 471 1874
rect 475 1870 519 1874
rect 523 1870 639 1874
rect 643 1870 711 1874
rect 715 1870 807 1874
rect 811 1870 887 1874
rect 891 1870 959 1874
rect 963 1870 1055 1874
rect 1059 1870 1103 1874
rect 1107 1870 1207 1874
rect 1211 1870 1239 1874
rect 1243 1870 1343 1874
rect 1347 1870 1367 1874
rect 1371 1870 1471 1874
rect 1475 1870 1495 1874
rect 1499 1870 1599 1874
rect 1603 1870 1631 1874
rect 1635 1870 1727 1874
rect 1731 1870 1831 1874
rect 1835 1870 1855 1874
rect 103 1869 1855 1870
rect 1861 1871 1862 1875
rect 1861 1870 3638 1871
rect 1861 1869 1871 1870
rect 1854 1866 1871 1869
rect 1875 1866 1903 1870
rect 1907 1866 1951 1870
rect 1955 1866 1983 1870
rect 1987 1866 2063 1870
rect 2067 1866 2095 1870
rect 2099 1866 2175 1870
rect 2179 1866 2207 1870
rect 2211 1866 2295 1870
rect 2299 1866 2327 1870
rect 2331 1866 2415 1870
rect 2419 1866 2463 1870
rect 2467 1866 2535 1870
rect 2539 1866 2631 1870
rect 2635 1866 2655 1870
rect 2659 1866 2783 1870
rect 2787 1866 2831 1870
rect 2835 1866 2919 1870
rect 2923 1866 3055 1870
rect 3059 1866 3063 1870
rect 3067 1866 3215 1870
rect 3219 1866 3295 1870
rect 3299 1866 3375 1870
rect 3379 1866 3511 1870
rect 3515 1866 3591 1870
rect 3595 1866 3638 1870
rect 1854 1865 3638 1866
rect 84 1793 85 1799
rect 91 1798 1843 1799
rect 91 1794 111 1798
rect 115 1794 135 1798
rect 139 1794 311 1798
rect 315 1794 503 1798
rect 507 1794 511 1798
rect 515 1794 687 1798
rect 691 1794 703 1798
rect 707 1794 847 1798
rect 851 1794 879 1798
rect 883 1794 991 1798
rect 995 1794 1047 1798
rect 1051 1794 1127 1798
rect 1131 1794 1199 1798
rect 1203 1794 1247 1798
rect 1251 1794 1335 1798
rect 1339 1794 1359 1798
rect 1363 1794 1463 1798
rect 1467 1794 1559 1798
rect 1563 1794 1591 1798
rect 1595 1794 1663 1798
rect 1667 1794 1719 1798
rect 1723 1794 1743 1798
rect 1747 1794 1831 1798
rect 1835 1794 1843 1798
rect 91 1793 1843 1794
rect 1849 1793 1850 1799
rect 1842 1773 1843 1779
rect 1849 1778 3619 1779
rect 1849 1774 1871 1778
rect 1875 1774 1895 1778
rect 1899 1774 1975 1778
rect 1979 1774 2023 1778
rect 2027 1774 2087 1778
rect 2091 1774 2183 1778
rect 2187 1774 2199 1778
rect 2203 1774 2319 1778
rect 2323 1774 2351 1778
rect 2355 1774 2455 1778
rect 2459 1774 2551 1778
rect 2555 1774 2623 1778
rect 2627 1774 2775 1778
rect 2779 1774 2823 1778
rect 2827 1774 3015 1778
rect 3019 1774 3047 1778
rect 3051 1774 3271 1778
rect 3275 1774 3287 1778
rect 3291 1774 3503 1778
rect 3507 1774 3591 1778
rect 3595 1774 3619 1778
rect 1849 1773 3619 1774
rect 3625 1773 3626 1779
rect 96 1709 97 1715
rect 103 1714 1855 1715
rect 103 1710 111 1714
rect 115 1710 143 1714
rect 147 1710 239 1714
rect 243 1710 319 1714
rect 323 1710 367 1714
rect 371 1710 487 1714
rect 491 1710 511 1714
rect 515 1710 607 1714
rect 611 1710 695 1714
rect 699 1710 719 1714
rect 723 1710 823 1714
rect 827 1710 855 1714
rect 859 1710 927 1714
rect 931 1710 999 1714
rect 1003 1710 1023 1714
rect 1027 1710 1119 1714
rect 1123 1710 1135 1714
rect 1139 1710 1215 1714
rect 1219 1710 1255 1714
rect 1259 1710 1319 1714
rect 1323 1710 1367 1714
rect 1371 1710 1471 1714
rect 1475 1710 1567 1714
rect 1571 1710 1671 1714
rect 1675 1710 1751 1714
rect 1755 1710 1831 1714
rect 1835 1710 1855 1714
rect 103 1709 1855 1710
rect 1861 1709 1862 1715
rect 1854 1697 1855 1703
rect 1861 1702 3631 1703
rect 1861 1698 1871 1702
rect 1875 1698 1903 1702
rect 1907 1698 1991 1702
rect 1995 1698 2031 1702
rect 2035 1698 2111 1702
rect 2115 1698 2191 1702
rect 2195 1698 2231 1702
rect 2235 1698 2351 1702
rect 2355 1698 2359 1702
rect 2363 1698 2479 1702
rect 2483 1698 2559 1702
rect 2563 1698 2607 1702
rect 2611 1698 2743 1702
rect 2747 1698 2783 1702
rect 2787 1698 2887 1702
rect 2891 1698 3023 1702
rect 3027 1698 3039 1702
rect 3043 1698 3199 1702
rect 3203 1698 3279 1702
rect 3283 1698 3367 1702
rect 3371 1698 3511 1702
rect 3515 1698 3591 1702
rect 3595 1698 3631 1702
rect 1861 1697 3631 1698
rect 3637 1697 3638 1703
rect 84 1625 85 1631
rect 91 1630 1843 1631
rect 91 1626 111 1630
rect 115 1626 135 1630
rect 139 1626 175 1630
rect 179 1626 231 1630
rect 235 1626 311 1630
rect 315 1626 359 1630
rect 363 1626 439 1630
rect 443 1626 479 1630
rect 483 1626 567 1630
rect 571 1626 599 1630
rect 603 1626 687 1630
rect 691 1626 711 1630
rect 715 1626 799 1630
rect 803 1626 815 1630
rect 819 1626 903 1630
rect 907 1626 919 1630
rect 923 1626 999 1630
rect 1003 1626 1015 1630
rect 1019 1626 1095 1630
rect 1099 1626 1111 1630
rect 1115 1626 1199 1630
rect 1203 1626 1207 1630
rect 1211 1626 1303 1630
rect 1307 1626 1311 1630
rect 1315 1626 1831 1630
rect 1835 1626 1843 1630
rect 91 1625 1843 1626
rect 1849 1627 1850 1631
rect 1849 1626 3626 1627
rect 1849 1625 1871 1626
rect 1842 1622 1871 1625
rect 1875 1622 1895 1626
rect 1899 1622 1927 1626
rect 1931 1622 1983 1626
rect 1987 1622 2023 1626
rect 2027 1622 2103 1626
rect 2107 1622 2135 1626
rect 2139 1622 2223 1626
rect 2227 1622 2263 1626
rect 2267 1622 2343 1626
rect 2347 1622 2391 1626
rect 2395 1622 2471 1626
rect 2475 1622 2527 1626
rect 2531 1622 2599 1626
rect 2603 1622 2671 1626
rect 2675 1622 2735 1626
rect 2739 1622 2823 1626
rect 2827 1622 2879 1626
rect 2883 1622 2983 1626
rect 2987 1622 3031 1626
rect 3035 1622 3159 1626
rect 3163 1622 3191 1626
rect 3195 1622 3343 1626
rect 3347 1622 3359 1626
rect 3363 1622 3503 1626
rect 3507 1622 3591 1626
rect 3595 1622 3626 1626
rect 1842 1621 3626 1622
rect 96 1541 97 1547
rect 103 1546 1855 1547
rect 103 1542 111 1546
rect 115 1542 183 1546
rect 187 1542 239 1546
rect 243 1542 319 1546
rect 323 1542 343 1546
rect 347 1542 447 1546
rect 451 1542 463 1546
rect 467 1542 575 1546
rect 579 1542 591 1546
rect 595 1542 695 1546
rect 699 1542 719 1546
rect 723 1542 807 1546
rect 811 1542 855 1546
rect 859 1542 911 1546
rect 915 1542 983 1546
rect 987 1542 1007 1546
rect 1011 1542 1103 1546
rect 1107 1542 1111 1546
rect 1115 1542 1207 1546
rect 1211 1542 1231 1546
rect 1235 1542 1311 1546
rect 1315 1542 1343 1546
rect 1347 1542 1455 1546
rect 1459 1542 1575 1546
rect 1579 1542 1831 1546
rect 1835 1542 1855 1546
rect 103 1541 1855 1542
rect 1861 1543 1862 1547
rect 1861 1542 3638 1543
rect 1861 1541 1871 1542
rect 1854 1538 1871 1541
rect 1875 1538 1935 1542
rect 1939 1538 2031 1542
rect 2035 1538 2135 1542
rect 2139 1538 2143 1542
rect 2147 1538 2255 1542
rect 2259 1538 2271 1542
rect 2275 1538 2383 1542
rect 2387 1538 2399 1542
rect 2403 1538 2511 1542
rect 2515 1538 2535 1542
rect 2539 1538 2639 1542
rect 2643 1538 2679 1542
rect 2683 1538 2767 1542
rect 2771 1538 2831 1542
rect 2835 1538 2887 1542
rect 2891 1538 2991 1542
rect 2995 1538 3007 1542
rect 3011 1538 3119 1542
rect 3123 1538 3167 1542
rect 3171 1538 3231 1542
rect 3235 1538 3351 1542
rect 3355 1538 3511 1542
rect 3515 1538 3591 1542
rect 3595 1538 3638 1542
rect 1854 1537 3638 1538
rect 84 1453 85 1459
rect 91 1458 1843 1459
rect 91 1454 111 1458
rect 115 1454 231 1458
rect 235 1454 279 1458
rect 283 1454 335 1458
rect 339 1454 383 1458
rect 387 1454 455 1458
rect 459 1454 511 1458
rect 515 1454 583 1458
rect 587 1454 655 1458
rect 659 1454 711 1458
rect 715 1454 807 1458
rect 811 1454 847 1458
rect 851 1454 959 1458
rect 963 1454 975 1458
rect 979 1454 1103 1458
rect 1107 1454 1111 1458
rect 1115 1454 1223 1458
rect 1227 1454 1247 1458
rect 1251 1454 1335 1458
rect 1339 1454 1383 1458
rect 1387 1454 1447 1458
rect 1451 1454 1511 1458
rect 1515 1454 1567 1458
rect 1571 1454 1639 1458
rect 1643 1454 1743 1458
rect 1747 1454 1831 1458
rect 1835 1454 1843 1458
rect 91 1453 1843 1454
rect 1849 1458 3626 1459
rect 1849 1454 1871 1458
rect 1875 1454 2127 1458
rect 2131 1454 2247 1458
rect 2251 1454 2343 1458
rect 2347 1454 2375 1458
rect 2379 1454 2455 1458
rect 2459 1454 2503 1458
rect 2507 1454 2575 1458
rect 2579 1454 2631 1458
rect 2635 1454 2703 1458
rect 2707 1454 2759 1458
rect 2763 1454 2831 1458
rect 2835 1454 2879 1458
rect 2883 1454 2951 1458
rect 2955 1454 2999 1458
rect 3003 1454 3071 1458
rect 3075 1454 3111 1458
rect 3115 1454 3183 1458
rect 3187 1454 3223 1458
rect 3227 1454 3295 1458
rect 3299 1454 3343 1458
rect 3347 1454 3407 1458
rect 3411 1454 3503 1458
rect 3507 1454 3591 1458
rect 3595 1454 3626 1458
rect 1849 1453 3626 1454
rect 1854 1369 1855 1375
rect 1861 1374 3631 1375
rect 1861 1370 1871 1374
rect 1875 1370 2255 1374
rect 2259 1370 2351 1374
rect 2355 1370 2399 1374
rect 2403 1370 2463 1374
rect 2467 1370 2503 1374
rect 2507 1370 2583 1374
rect 2587 1370 2615 1374
rect 2619 1370 2711 1374
rect 2715 1370 2735 1374
rect 2739 1370 2839 1374
rect 2843 1370 2847 1374
rect 2851 1370 2959 1374
rect 2963 1370 3071 1374
rect 3075 1370 3079 1374
rect 3083 1370 3183 1374
rect 3187 1370 3191 1374
rect 3195 1370 3295 1374
rect 3299 1370 3303 1374
rect 3307 1370 3415 1374
rect 3419 1370 3511 1374
rect 3515 1370 3591 1374
rect 3595 1370 3631 1374
rect 1861 1369 3631 1370
rect 3637 1369 3638 1375
rect 1854 1367 1862 1369
rect 96 1361 97 1367
rect 103 1366 1855 1367
rect 103 1362 111 1366
rect 115 1362 223 1366
rect 227 1362 287 1366
rect 291 1362 335 1366
rect 339 1362 391 1366
rect 395 1362 471 1366
rect 475 1362 519 1366
rect 523 1362 623 1366
rect 627 1362 663 1366
rect 667 1362 783 1366
rect 787 1362 815 1366
rect 819 1362 943 1366
rect 947 1362 967 1366
rect 971 1362 1095 1366
rect 1099 1362 1119 1366
rect 1123 1362 1239 1366
rect 1243 1362 1255 1366
rect 1259 1362 1375 1366
rect 1379 1362 1391 1366
rect 1395 1362 1511 1366
rect 1515 1362 1519 1366
rect 1523 1362 1639 1366
rect 1643 1362 1647 1366
rect 1651 1362 1751 1366
rect 1755 1362 1831 1366
rect 1835 1362 1855 1366
rect 103 1361 1855 1362
rect 1861 1361 1862 1367
rect 84 1285 85 1291
rect 91 1290 1843 1291
rect 91 1286 111 1290
rect 115 1286 135 1290
rect 139 1286 215 1290
rect 219 1286 327 1290
rect 331 1286 335 1290
rect 339 1286 463 1290
rect 467 1286 607 1290
rect 611 1286 615 1290
rect 619 1286 751 1290
rect 755 1286 775 1290
rect 779 1286 903 1290
rect 907 1286 935 1290
rect 939 1286 1047 1290
rect 1051 1286 1087 1290
rect 1091 1286 1183 1290
rect 1187 1286 1231 1290
rect 1235 1286 1303 1290
rect 1307 1286 1367 1290
rect 1371 1286 1423 1290
rect 1427 1286 1503 1290
rect 1507 1286 1535 1290
rect 1539 1286 1631 1290
rect 1635 1286 1647 1290
rect 1651 1286 1743 1290
rect 1747 1286 1831 1290
rect 1835 1286 1843 1290
rect 91 1285 1843 1286
rect 1849 1285 1850 1291
rect 1842 1283 1850 1285
rect 1842 1277 1843 1283
rect 1849 1282 3619 1283
rect 1849 1278 1871 1282
rect 1875 1278 1895 1282
rect 1899 1278 2071 1282
rect 2075 1278 2255 1282
rect 2259 1278 2391 1282
rect 2395 1278 2423 1282
rect 2427 1278 2495 1282
rect 2499 1278 2583 1282
rect 2587 1278 2607 1282
rect 2611 1278 2727 1282
rect 2731 1278 2735 1282
rect 2739 1278 2839 1282
rect 2843 1278 2879 1282
rect 2883 1278 2951 1282
rect 2955 1278 3015 1282
rect 3019 1278 3063 1282
rect 3067 1278 3143 1282
rect 3147 1278 3175 1282
rect 3179 1278 3271 1282
rect 3275 1278 3287 1282
rect 3291 1278 3399 1282
rect 3403 1278 3407 1282
rect 3411 1278 3503 1282
rect 3507 1278 3591 1282
rect 3595 1278 3619 1282
rect 1849 1277 3619 1278
rect 3625 1277 3626 1283
rect 96 1197 97 1203
rect 103 1202 1855 1203
rect 103 1198 111 1202
rect 115 1198 143 1202
rect 147 1198 223 1202
rect 227 1198 255 1202
rect 259 1198 343 1202
rect 347 1198 383 1202
rect 387 1198 471 1202
rect 475 1198 503 1202
rect 507 1198 615 1202
rect 619 1198 719 1202
rect 723 1198 759 1202
rect 763 1198 815 1202
rect 819 1198 911 1202
rect 915 1198 999 1202
rect 1003 1198 1055 1202
rect 1059 1198 1095 1202
rect 1099 1198 1191 1202
rect 1195 1198 1287 1202
rect 1291 1198 1311 1202
rect 1315 1198 1431 1202
rect 1435 1198 1543 1202
rect 1547 1198 1655 1202
rect 1659 1198 1751 1202
rect 1755 1198 1831 1202
rect 1835 1198 1855 1202
rect 103 1197 1855 1198
rect 1861 1199 1862 1203
rect 1861 1198 3638 1199
rect 1861 1197 1871 1198
rect 1854 1194 1871 1197
rect 1875 1194 1903 1198
rect 1907 1194 1991 1198
rect 1995 1194 2079 1198
rect 2083 1194 2103 1198
rect 2107 1194 2215 1198
rect 2219 1194 2263 1198
rect 2267 1194 2327 1198
rect 2331 1194 2431 1198
rect 2435 1194 2447 1198
rect 2451 1194 2575 1198
rect 2579 1194 2591 1198
rect 2595 1194 2719 1198
rect 2723 1194 2743 1198
rect 2747 1194 2871 1198
rect 2875 1194 2887 1198
rect 2891 1194 3023 1198
rect 3027 1194 3031 1198
rect 3035 1194 3151 1198
rect 3155 1194 3191 1198
rect 3195 1194 3279 1198
rect 3283 1194 3359 1198
rect 3363 1194 3407 1198
rect 3411 1194 3511 1198
rect 3515 1194 3591 1198
rect 3595 1194 3638 1198
rect 1854 1193 3638 1194
rect 84 1109 85 1115
rect 91 1114 1843 1115
rect 91 1110 111 1114
rect 115 1110 135 1114
rect 139 1110 247 1114
rect 251 1110 255 1114
rect 259 1110 375 1114
rect 379 1110 399 1114
rect 403 1110 495 1114
rect 499 1110 535 1114
rect 539 1110 607 1114
rect 611 1110 663 1114
rect 667 1110 711 1114
rect 715 1110 783 1114
rect 787 1110 807 1114
rect 811 1110 895 1114
rect 899 1110 903 1114
rect 907 1110 991 1114
rect 995 1110 999 1114
rect 1003 1110 1087 1114
rect 1091 1110 1095 1114
rect 1099 1110 1183 1114
rect 1187 1110 1191 1114
rect 1195 1110 1279 1114
rect 1283 1110 1295 1114
rect 1299 1110 1399 1114
rect 1403 1110 1831 1114
rect 1835 1110 1843 1114
rect 91 1109 1843 1110
rect 1849 1114 3626 1115
rect 1849 1110 1871 1114
rect 1875 1110 1895 1114
rect 1899 1110 1967 1114
rect 1971 1110 1983 1114
rect 1987 1110 2047 1114
rect 2051 1110 2095 1114
rect 2099 1110 2135 1114
rect 2139 1110 2207 1114
rect 2211 1110 2231 1114
rect 2235 1110 2319 1114
rect 2323 1110 2335 1114
rect 2339 1110 2439 1114
rect 2443 1110 2551 1114
rect 2555 1110 2567 1114
rect 2571 1110 2679 1114
rect 2683 1110 2711 1114
rect 2715 1110 2823 1114
rect 2827 1110 2863 1114
rect 2867 1110 2983 1114
rect 2987 1110 3023 1114
rect 3027 1110 3159 1114
rect 3163 1110 3183 1114
rect 3187 1110 3343 1114
rect 3347 1110 3351 1114
rect 3355 1110 3503 1114
rect 3507 1110 3591 1114
rect 3595 1110 3626 1114
rect 1849 1109 3626 1110
rect 96 1025 97 1031
rect 103 1030 1855 1031
rect 103 1026 111 1030
rect 115 1026 143 1030
rect 147 1026 263 1030
rect 267 1026 271 1030
rect 275 1026 407 1030
rect 411 1026 423 1030
rect 427 1026 543 1030
rect 547 1026 583 1030
rect 587 1026 671 1030
rect 675 1026 735 1030
rect 739 1026 791 1030
rect 795 1026 887 1030
rect 891 1026 903 1030
rect 907 1026 1007 1030
rect 1011 1026 1031 1030
rect 1035 1026 1103 1030
rect 1107 1026 1159 1030
rect 1163 1026 1199 1030
rect 1203 1026 1279 1030
rect 1283 1026 1303 1030
rect 1307 1026 1399 1030
rect 1403 1026 1407 1030
rect 1411 1026 1519 1030
rect 1523 1026 1639 1030
rect 1643 1026 1831 1030
rect 1835 1026 1855 1030
rect 103 1025 1855 1026
rect 1861 1030 3638 1031
rect 1861 1026 1871 1030
rect 1875 1026 1975 1030
rect 1979 1026 2031 1030
rect 2035 1026 2055 1030
rect 2059 1026 2127 1030
rect 2131 1026 2143 1030
rect 2147 1026 2231 1030
rect 2235 1026 2239 1030
rect 2243 1026 2343 1030
rect 2347 1026 2351 1030
rect 2355 1026 2447 1030
rect 2451 1026 2471 1030
rect 2475 1026 2559 1030
rect 2563 1026 2599 1030
rect 2603 1026 2687 1030
rect 2691 1026 2727 1030
rect 2731 1026 2831 1030
rect 2835 1026 2855 1030
rect 2859 1026 2983 1030
rect 2987 1026 2991 1030
rect 2995 1026 3111 1030
rect 3115 1026 3167 1030
rect 3171 1026 3247 1030
rect 3251 1026 3351 1030
rect 3355 1026 3391 1030
rect 3395 1026 3511 1030
rect 3515 1026 3591 1030
rect 3595 1026 3638 1030
rect 1861 1025 3638 1026
rect 84 941 85 947
rect 91 946 1843 947
rect 91 942 111 946
rect 115 942 135 946
rect 139 942 215 946
rect 219 942 263 946
rect 267 942 335 946
rect 339 942 415 946
rect 419 942 463 946
rect 467 942 575 946
rect 579 942 599 946
rect 603 942 727 946
rect 731 942 735 946
rect 739 942 863 946
rect 867 942 879 946
rect 883 942 991 946
rect 995 942 1023 946
rect 1027 942 1111 946
rect 1115 942 1151 946
rect 1155 942 1223 946
rect 1227 942 1271 946
rect 1275 942 1335 946
rect 1339 942 1391 946
rect 1395 942 1455 946
rect 1459 942 1511 946
rect 1515 942 1631 946
rect 1635 942 1831 946
rect 1835 942 1843 946
rect 91 941 1843 942
rect 1849 946 3626 947
rect 1849 942 1871 946
rect 1875 942 1895 946
rect 1899 942 1983 946
rect 1987 942 2023 946
rect 2027 942 2111 946
rect 2115 942 2119 946
rect 2123 942 2223 946
rect 2227 942 2263 946
rect 2267 942 2343 946
rect 2347 942 2423 946
rect 2427 942 2463 946
rect 2467 942 2583 946
rect 2587 942 2591 946
rect 2595 942 2719 946
rect 2723 942 2735 946
rect 2739 942 2847 946
rect 2851 942 2879 946
rect 2883 942 2975 946
rect 2979 942 3015 946
rect 3019 942 3103 946
rect 3107 942 3143 946
rect 3147 942 3239 946
rect 3243 942 3271 946
rect 3275 942 3383 946
rect 3387 942 3399 946
rect 3403 942 3503 946
rect 3507 942 3591 946
rect 3595 942 3626 946
rect 1849 941 3626 942
rect 1854 862 3638 863
rect 1854 859 1871 862
rect 96 853 97 859
rect 103 858 1855 859
rect 103 854 111 858
rect 115 854 143 858
rect 147 854 223 858
rect 227 854 303 858
rect 307 854 343 858
rect 347 854 391 858
rect 395 854 471 858
rect 475 854 495 858
rect 499 854 599 858
rect 603 854 607 858
rect 611 854 711 858
rect 715 854 743 858
rect 747 854 839 858
rect 843 854 871 858
rect 875 854 991 858
rect 995 854 999 858
rect 1003 854 1119 858
rect 1123 854 1167 858
rect 1171 854 1231 858
rect 1235 854 1343 858
rect 1347 854 1359 858
rect 1363 854 1463 858
rect 1467 854 1567 858
rect 1571 854 1751 858
rect 1755 854 1831 858
rect 1835 854 1855 858
rect 103 853 1855 854
rect 1861 858 1871 859
rect 1875 858 1903 862
rect 1907 858 1991 862
rect 1995 858 2039 862
rect 2043 858 2119 862
rect 2123 858 2215 862
rect 2219 858 2271 862
rect 2275 858 2391 862
rect 2395 858 2431 862
rect 2435 858 2567 862
rect 2571 858 2591 862
rect 2595 858 2735 862
rect 2739 858 2743 862
rect 2747 858 2887 862
rect 2891 858 3023 862
rect 3027 858 3031 862
rect 3035 858 3151 862
rect 3155 858 3159 862
rect 3163 858 3279 862
rect 3283 858 3287 862
rect 3291 858 3407 862
rect 3411 858 3511 862
rect 3515 858 3591 862
rect 3595 858 3638 862
rect 1861 857 3638 858
rect 1861 853 1862 857
rect 84 773 85 779
rect 91 778 1843 779
rect 91 774 111 778
rect 115 774 135 778
rect 139 774 199 778
rect 203 774 215 778
rect 219 774 287 778
rect 291 774 295 778
rect 299 774 383 778
rect 387 774 391 778
rect 395 774 487 778
rect 491 774 503 778
rect 507 774 591 778
rect 595 774 615 778
rect 619 774 703 778
rect 707 774 735 778
rect 739 774 831 778
rect 835 774 855 778
rect 859 774 983 778
rect 987 774 1111 778
rect 1115 774 1159 778
rect 1163 774 1239 778
rect 1243 774 1351 778
rect 1355 774 1367 778
rect 1371 774 1495 778
rect 1499 774 1559 778
rect 1563 774 1631 778
rect 1635 774 1743 778
rect 1747 774 1831 778
rect 1835 774 1843 778
rect 91 773 1843 774
rect 1849 773 1850 779
rect 1842 771 1850 773
rect 1842 765 1843 771
rect 1849 770 3619 771
rect 1849 766 1871 770
rect 1875 766 1895 770
rect 1899 766 2023 770
rect 2027 766 2031 770
rect 2035 766 2191 770
rect 2195 766 2207 770
rect 2211 766 2359 770
rect 2363 766 2383 770
rect 2387 766 2519 770
rect 2523 766 2559 770
rect 2563 766 2679 770
rect 2683 766 2727 770
rect 2731 766 2831 770
rect 2835 766 2879 770
rect 2883 766 2975 770
rect 2979 766 3023 770
rect 3027 766 3111 770
rect 3115 766 3151 770
rect 3155 766 3247 770
rect 3251 766 3279 770
rect 3283 766 3383 770
rect 3387 766 3399 770
rect 3403 766 3503 770
rect 3507 766 3591 770
rect 3595 766 3619 770
rect 1849 765 3619 766
rect 3625 765 3626 771
rect 1854 690 3638 691
rect 1854 687 1871 690
rect 96 681 97 687
rect 103 686 1855 687
rect 103 682 111 686
rect 115 682 207 686
rect 211 682 295 686
rect 299 682 383 686
rect 387 682 399 686
rect 403 682 479 686
rect 483 682 511 686
rect 515 682 591 686
rect 595 682 623 686
rect 627 682 719 686
rect 723 682 743 686
rect 747 682 855 686
rect 859 682 863 686
rect 867 682 991 686
rect 995 682 1119 686
rect 1123 682 1127 686
rect 1131 682 1247 686
rect 1251 682 1255 686
rect 1259 682 1375 686
rect 1379 682 1383 686
rect 1387 682 1503 686
rect 1507 682 1631 686
rect 1635 682 1639 686
rect 1643 682 1751 686
rect 1755 682 1831 686
rect 1835 682 1855 686
rect 103 681 1855 682
rect 1861 686 1871 687
rect 1875 686 2031 690
rect 2035 686 2095 690
rect 2099 686 2175 690
rect 2179 686 2199 690
rect 2203 686 2263 690
rect 2267 686 2359 690
rect 2363 686 2367 690
rect 2371 686 2463 690
rect 2467 686 2527 690
rect 2531 686 2567 690
rect 2571 686 2679 690
rect 2683 686 2687 690
rect 2691 686 2799 690
rect 2803 686 2839 690
rect 2843 686 2927 690
rect 2931 686 2983 690
rect 2987 686 3071 690
rect 3075 686 3119 690
rect 3123 686 3223 690
rect 3227 686 3255 690
rect 3259 686 3375 690
rect 3379 686 3391 690
rect 3395 686 3511 690
rect 3515 686 3591 690
rect 3595 686 3638 690
rect 1861 685 3638 686
rect 1861 681 1862 685
rect 84 597 85 603
rect 91 602 1843 603
rect 91 598 111 602
rect 115 598 375 602
rect 379 598 471 602
rect 475 598 583 602
rect 587 598 599 602
rect 603 598 687 602
rect 691 598 711 602
rect 715 598 783 602
rect 787 598 847 602
rect 851 598 887 602
rect 891 598 983 602
rect 987 598 991 602
rect 995 598 1095 602
rect 1099 598 1119 602
rect 1123 598 1199 602
rect 1203 598 1247 602
rect 1251 598 1303 602
rect 1307 598 1375 602
rect 1379 598 1399 602
rect 1403 598 1495 602
rect 1499 598 1503 602
rect 1507 598 1607 602
rect 1611 598 1623 602
rect 1627 598 1711 602
rect 1715 598 1743 602
rect 1747 598 1831 602
rect 1835 598 1843 602
rect 91 597 1843 598
rect 1849 602 3626 603
rect 1849 598 1871 602
rect 1875 598 2087 602
rect 2091 598 2167 602
rect 2171 598 2247 602
rect 2251 598 2255 602
rect 2259 598 2327 602
rect 2331 598 2351 602
rect 2355 598 2407 602
rect 2411 598 2455 602
rect 2459 598 2487 602
rect 2491 598 2559 602
rect 2563 598 2567 602
rect 2571 598 2647 602
rect 2651 598 2671 602
rect 2675 598 2743 602
rect 2747 598 2791 602
rect 2795 598 2863 602
rect 2867 598 2919 602
rect 2923 598 2999 602
rect 3003 598 3063 602
rect 3067 598 3159 602
rect 3163 598 3215 602
rect 3219 598 3327 602
rect 3331 598 3367 602
rect 3371 598 3495 602
rect 3499 598 3503 602
rect 3507 598 3591 602
rect 3595 598 3626 602
rect 1849 597 3626 598
rect 96 513 97 519
rect 103 518 1855 519
rect 103 514 111 518
rect 115 514 367 518
rect 371 514 463 518
rect 467 514 575 518
rect 579 514 607 518
rect 611 514 695 518
rect 699 514 703 518
rect 707 514 791 518
rect 795 514 839 518
rect 843 514 895 518
rect 899 514 975 518
rect 979 514 999 518
rect 1003 514 1103 518
rect 1107 514 1111 518
rect 1115 514 1207 518
rect 1211 514 1239 518
rect 1243 514 1311 518
rect 1315 514 1359 518
rect 1363 514 1407 518
rect 1411 514 1471 518
rect 1475 514 1511 518
rect 1515 514 1583 518
rect 1587 514 1615 518
rect 1619 514 1703 518
rect 1707 514 1719 518
rect 1723 514 1831 518
rect 1835 514 1855 518
rect 103 513 1855 514
rect 1861 518 3638 519
rect 1861 514 1871 518
rect 1875 514 2159 518
rect 2163 514 2175 518
rect 2179 514 2239 518
rect 2243 514 2255 518
rect 2259 514 2319 518
rect 2323 514 2335 518
rect 2339 514 2399 518
rect 2403 514 2415 518
rect 2419 514 2479 518
rect 2483 514 2495 518
rect 2499 514 2559 518
rect 2563 514 2575 518
rect 2579 514 2639 518
rect 2643 514 2655 518
rect 2659 514 2735 518
rect 2739 514 2751 518
rect 2755 514 2855 518
rect 2859 514 2871 518
rect 2875 514 2991 518
rect 2995 514 3007 518
rect 3011 514 3143 518
rect 3147 514 3167 518
rect 3171 514 3311 518
rect 3315 514 3335 518
rect 3339 514 3479 518
rect 3483 514 3503 518
rect 3507 514 3591 518
rect 3595 514 3638 518
rect 1861 513 3638 514
rect 84 425 85 431
rect 91 430 1843 431
rect 91 426 111 430
rect 115 426 135 430
rect 139 426 223 430
rect 227 426 359 430
rect 363 426 455 430
rect 459 426 511 430
rect 515 426 567 430
rect 571 426 679 430
rect 683 426 695 430
rect 699 426 831 430
rect 835 426 839 430
rect 843 426 967 430
rect 971 426 999 430
rect 1003 426 1103 430
rect 1107 426 1143 430
rect 1147 426 1231 430
rect 1235 426 1279 430
rect 1283 426 1351 430
rect 1355 426 1415 430
rect 1419 426 1463 430
rect 1467 426 1551 430
rect 1555 426 1575 430
rect 1579 426 1687 430
rect 1691 426 1695 430
rect 1699 426 1831 430
rect 1835 426 1843 430
rect 91 425 1843 426
rect 1849 430 3626 431
rect 1849 426 1871 430
rect 1875 426 2151 430
rect 2155 426 2159 430
rect 2163 426 2231 430
rect 2235 426 2239 430
rect 2243 426 2311 430
rect 2315 426 2319 430
rect 2323 426 2391 430
rect 2395 426 2399 430
rect 2403 426 2471 430
rect 2475 426 2479 430
rect 2483 426 2551 430
rect 2555 426 2559 430
rect 2563 426 2631 430
rect 2635 426 2639 430
rect 2643 426 2727 430
rect 2731 426 2735 430
rect 2739 426 2839 430
rect 2843 426 2847 430
rect 2851 426 2959 430
rect 2963 426 2983 430
rect 2987 426 3087 430
rect 3091 426 3135 430
rect 3139 426 3231 430
rect 3235 426 3303 430
rect 3307 426 3375 430
rect 3379 426 3471 430
rect 3475 426 3503 430
rect 3507 426 3591 430
rect 3595 426 3626 430
rect 1849 425 3626 426
rect 96 341 97 347
rect 103 346 1855 347
rect 103 342 111 346
rect 115 342 143 346
rect 147 342 231 346
rect 235 342 279 346
rect 283 342 367 346
rect 371 342 455 346
rect 459 342 519 346
rect 523 342 639 346
rect 643 342 687 346
rect 691 342 823 346
rect 827 342 847 346
rect 851 342 999 346
rect 1003 342 1007 346
rect 1011 342 1151 346
rect 1155 342 1167 346
rect 1171 342 1287 346
rect 1291 342 1327 346
rect 1331 342 1423 346
rect 1427 342 1479 346
rect 1483 342 1559 346
rect 1563 342 1623 346
rect 1627 342 1695 346
rect 1699 342 1751 346
rect 1755 342 1831 346
rect 1835 342 1855 346
rect 103 341 1855 342
rect 1861 343 1862 347
rect 1861 342 3638 343
rect 1861 341 1871 342
rect 1854 338 1871 341
rect 1875 338 2031 342
rect 2035 338 2119 342
rect 2123 338 2167 342
rect 2171 338 2223 342
rect 2227 338 2247 342
rect 2251 338 2327 342
rect 2331 338 2335 342
rect 2339 338 2407 342
rect 2411 338 2447 342
rect 2451 338 2487 342
rect 2491 338 2567 342
rect 2571 338 2647 342
rect 2651 338 2695 342
rect 2699 338 2743 342
rect 2747 338 2839 342
rect 2843 338 2847 342
rect 2851 338 2967 342
rect 2971 338 2999 342
rect 3003 338 3095 342
rect 3099 338 3167 342
rect 3171 338 3239 342
rect 3243 338 3343 342
rect 3347 338 3383 342
rect 3387 338 3511 342
rect 3515 338 3591 342
rect 3595 338 3638 342
rect 1854 337 3638 338
rect 84 261 85 267
rect 91 266 1843 267
rect 91 262 111 266
rect 115 262 135 266
rect 139 262 271 266
rect 275 262 303 266
rect 307 262 391 266
rect 395 262 447 266
rect 451 262 495 266
rect 499 262 599 266
rect 603 262 631 266
rect 635 262 711 266
rect 715 262 815 266
rect 819 262 823 266
rect 827 262 943 266
rect 947 262 991 266
rect 995 262 1063 266
rect 1067 262 1159 266
rect 1163 262 1175 266
rect 1179 262 1287 266
rect 1291 262 1319 266
rect 1323 262 1407 266
rect 1411 262 1471 266
rect 1475 262 1527 266
rect 1531 262 1615 266
rect 1619 262 1647 266
rect 1651 262 1743 266
rect 1747 262 1831 266
rect 1835 262 1843 266
rect 91 261 1843 262
rect 1849 263 1850 267
rect 1849 262 3626 263
rect 1849 261 1871 262
rect 1842 258 1871 261
rect 1875 258 2023 262
rect 2027 258 2071 262
rect 2075 258 2111 262
rect 2115 258 2215 262
rect 2219 258 2319 262
rect 2323 258 2327 262
rect 2331 258 2439 262
rect 2443 258 2543 262
rect 2547 258 2559 262
rect 2563 258 2687 262
rect 2691 258 2743 262
rect 2747 258 2831 262
rect 2835 258 2927 262
rect 2931 258 2991 262
rect 2995 258 3087 262
rect 3091 258 3159 262
rect 3163 258 3239 262
rect 3243 258 3335 262
rect 3339 258 3383 262
rect 3387 258 3503 262
rect 3507 258 3591 262
rect 3595 258 3626 262
rect 1842 257 3626 258
rect 96 161 97 167
rect 103 166 1855 167
rect 103 162 111 166
rect 115 162 263 166
rect 267 162 311 166
rect 315 162 343 166
rect 347 162 399 166
rect 403 162 423 166
rect 427 162 503 166
rect 507 162 583 166
rect 587 162 607 166
rect 611 162 663 166
rect 667 162 719 166
rect 723 162 743 166
rect 747 162 823 166
rect 827 162 831 166
rect 835 162 903 166
rect 907 162 951 166
rect 955 162 983 166
rect 987 162 1063 166
rect 1067 162 1071 166
rect 1075 162 1143 166
rect 1147 162 1183 166
rect 1187 162 1223 166
rect 1227 162 1295 166
rect 1299 162 1303 166
rect 1307 162 1383 166
rect 1387 162 1415 166
rect 1419 162 1463 166
rect 1467 162 1535 166
rect 1539 162 1543 166
rect 1547 162 1655 166
rect 1659 162 1751 166
rect 1755 162 1831 166
rect 1835 162 1855 166
rect 103 161 1855 162
rect 1861 163 1862 167
rect 1861 162 3638 163
rect 1861 161 1871 162
rect 1854 158 1871 161
rect 1875 158 1903 162
rect 1907 158 1983 162
rect 1987 158 2063 162
rect 2067 158 2079 162
rect 2083 158 2143 162
rect 2147 158 2223 162
rect 2227 158 2303 162
rect 2307 158 2327 162
rect 2331 158 2399 162
rect 2403 158 2503 162
rect 2507 158 2551 162
rect 2555 158 2607 162
rect 2611 158 2711 162
rect 2715 158 2751 162
rect 2755 158 2815 162
rect 2819 158 2911 162
rect 2915 158 2935 162
rect 2939 158 2999 162
rect 3003 158 3087 162
rect 3091 158 3095 162
rect 3099 158 3175 162
rect 3179 158 3247 162
rect 3251 158 3263 162
rect 3267 158 3351 162
rect 3355 158 3391 162
rect 3395 158 3431 162
rect 3435 158 3511 162
rect 3515 158 3591 162
rect 3595 158 3638 162
rect 1854 157 3638 158
rect 84 85 85 91
rect 91 90 1843 91
rect 91 86 111 90
rect 115 86 255 90
rect 259 86 335 90
rect 339 86 415 90
rect 419 86 495 90
rect 499 86 575 90
rect 579 86 655 90
rect 659 86 735 90
rect 739 86 815 90
rect 819 86 895 90
rect 899 86 975 90
rect 979 86 1055 90
rect 1059 86 1135 90
rect 1139 86 1215 90
rect 1219 86 1295 90
rect 1299 86 1375 90
rect 1379 86 1455 90
rect 1459 86 1535 90
rect 1539 86 1831 90
rect 1835 86 1843 90
rect 91 85 1843 86
rect 1849 87 1850 91
rect 1849 86 3626 87
rect 1849 85 1871 86
rect 1842 82 1871 85
rect 1875 82 1895 86
rect 1899 82 1975 86
rect 1979 82 2055 86
rect 2059 82 2135 86
rect 2139 82 2215 86
rect 2219 82 2295 86
rect 2299 82 2391 86
rect 2395 82 2495 86
rect 2499 82 2599 86
rect 2603 82 2703 86
rect 2707 82 2807 86
rect 2811 82 2903 86
rect 2907 82 2991 86
rect 2995 82 3079 86
rect 3083 82 3167 86
rect 3171 82 3255 86
rect 3259 82 3343 86
rect 3347 82 3423 86
rect 3427 82 3503 86
rect 3507 82 3591 86
rect 3595 82 3626 86
rect 1842 81 3626 82
<< m5c >>
rect 97 3653 103 3659
rect 1855 3653 1861 3659
rect 1855 3625 1861 3631
rect 3631 3625 3637 3631
rect 85 3577 91 3583
rect 1843 3577 1849 3583
rect 1843 3549 1849 3555
rect 3619 3549 3625 3555
rect 97 3501 103 3507
rect 1855 3501 1861 3507
rect 1855 3473 1861 3479
rect 3631 3473 3637 3479
rect 85 3417 91 3423
rect 1843 3417 1849 3423
rect 1843 3389 1849 3395
rect 3619 3389 3625 3395
rect 97 3337 103 3343
rect 1855 3337 1861 3343
rect 1855 3309 1861 3315
rect 3631 3309 3637 3315
rect 85 3257 91 3263
rect 1843 3257 1849 3263
rect 1843 3229 1849 3235
rect 3619 3229 3625 3235
rect 97 3173 103 3179
rect 1855 3173 1861 3179
rect 1855 3153 1861 3159
rect 3631 3153 3637 3159
rect 85 3097 91 3103
rect 1843 3097 1849 3103
rect 1843 3069 1849 3075
rect 3619 3069 3625 3075
rect 97 3005 103 3011
rect 1855 3005 1861 3011
rect 1855 2989 1861 2995
rect 3631 2989 3637 2995
rect 85 2929 91 2935
rect 1843 2929 1849 2935
rect 1843 2901 1849 2907
rect 3619 2901 3625 2907
rect 97 2853 103 2859
rect 1855 2853 1861 2859
rect 1855 2825 1861 2831
rect 3631 2825 3637 2831
rect 85 2769 91 2775
rect 1843 2769 1849 2775
rect 1843 2737 1849 2743
rect 3619 2737 3625 2743
rect 97 2689 103 2695
rect 1855 2689 1861 2695
rect 1855 2661 1861 2667
rect 3631 2661 3637 2667
rect 85 2605 91 2611
rect 1843 2605 1849 2611
rect 1843 2581 1849 2587
rect 3619 2581 3625 2587
rect 97 2521 103 2527
rect 1855 2521 1861 2527
rect 1855 2505 1861 2511
rect 3631 2505 3637 2511
rect 85 2441 91 2447
rect 1843 2441 1849 2447
rect 1843 2421 1849 2427
rect 3619 2421 3625 2427
rect 97 2357 103 2363
rect 1855 2357 1861 2363
rect 1855 2341 1861 2347
rect 3631 2341 3637 2347
rect 85 2269 91 2275
rect 1843 2269 1849 2275
rect 97 2189 103 2195
rect 1855 2189 1861 2195
rect 1855 2181 1861 2187
rect 3631 2181 3637 2187
rect 85 2113 91 2119
rect 1843 2113 1849 2119
rect 1843 2105 1849 2111
rect 3619 2105 3625 2111
rect 97 2029 103 2035
rect 1855 2029 1861 2035
rect 85 1953 91 1959
rect 1843 1953 1849 1959
rect 1843 1945 1849 1951
rect 3619 1945 3625 1951
rect 97 1869 103 1875
rect 1855 1869 1861 1875
rect 85 1793 91 1799
rect 1843 1793 1849 1799
rect 1843 1773 1849 1779
rect 3619 1773 3625 1779
rect 97 1709 103 1715
rect 1855 1709 1861 1715
rect 1855 1697 1861 1703
rect 3631 1697 3637 1703
rect 85 1625 91 1631
rect 1843 1625 1849 1631
rect 97 1541 103 1547
rect 1855 1541 1861 1547
rect 85 1453 91 1459
rect 1843 1453 1849 1459
rect 1855 1369 1861 1375
rect 3631 1369 3637 1375
rect 97 1361 103 1367
rect 1855 1361 1861 1367
rect 85 1285 91 1291
rect 1843 1285 1849 1291
rect 1843 1277 1849 1283
rect 3619 1277 3625 1283
rect 97 1197 103 1203
rect 1855 1197 1861 1203
rect 85 1109 91 1115
rect 1843 1109 1849 1115
rect 97 1025 103 1031
rect 1855 1025 1861 1031
rect 85 941 91 947
rect 1843 941 1849 947
rect 97 853 103 859
rect 1855 853 1861 859
rect 85 773 91 779
rect 1843 773 1849 779
rect 1843 765 1849 771
rect 3619 765 3625 771
rect 97 681 103 687
rect 1855 681 1861 687
rect 85 597 91 603
rect 1843 597 1849 603
rect 97 513 103 519
rect 1855 513 1861 519
rect 85 425 91 431
rect 1843 425 1849 431
rect 97 341 103 347
rect 1855 341 1861 347
rect 85 261 91 267
rect 1843 261 1849 267
rect 97 161 103 167
rect 1855 161 1861 167
rect 85 85 91 91
rect 1843 85 1849 91
<< m5 >>
rect 84 3583 92 3672
rect 84 3577 85 3583
rect 91 3577 92 3583
rect 84 3423 92 3577
rect 84 3417 85 3423
rect 91 3417 92 3423
rect 84 3263 92 3417
rect 84 3257 85 3263
rect 91 3257 92 3263
rect 84 3103 92 3257
rect 84 3097 85 3103
rect 91 3097 92 3103
rect 84 2935 92 3097
rect 84 2929 85 2935
rect 91 2929 92 2935
rect 84 2775 92 2929
rect 84 2769 85 2775
rect 91 2769 92 2775
rect 84 2611 92 2769
rect 84 2605 85 2611
rect 91 2605 92 2611
rect 84 2447 92 2605
rect 84 2441 85 2447
rect 91 2441 92 2447
rect 84 2275 92 2441
rect 84 2269 85 2275
rect 91 2269 92 2275
rect 84 2119 92 2269
rect 84 2113 85 2119
rect 91 2113 92 2119
rect 84 1959 92 2113
rect 84 1953 85 1959
rect 91 1953 92 1959
rect 84 1799 92 1953
rect 84 1793 85 1799
rect 91 1793 92 1799
rect 84 1631 92 1793
rect 84 1625 85 1631
rect 91 1625 92 1631
rect 84 1459 92 1625
rect 84 1453 85 1459
rect 91 1453 92 1459
rect 84 1291 92 1453
rect 84 1285 85 1291
rect 91 1285 92 1291
rect 84 1115 92 1285
rect 84 1109 85 1115
rect 91 1109 92 1115
rect 84 947 92 1109
rect 84 941 85 947
rect 91 941 92 947
rect 84 779 92 941
rect 84 773 85 779
rect 91 773 92 779
rect 84 603 92 773
rect 84 597 85 603
rect 91 597 92 603
rect 84 431 92 597
rect 84 425 85 431
rect 91 425 92 431
rect 84 267 92 425
rect 84 261 85 267
rect 91 261 92 267
rect 84 91 92 261
rect 84 85 85 91
rect 91 85 92 91
rect 84 72 92 85
rect 96 3659 104 3672
rect 96 3653 97 3659
rect 103 3653 104 3659
rect 96 3507 104 3653
rect 96 3501 97 3507
rect 103 3501 104 3507
rect 96 3343 104 3501
rect 96 3337 97 3343
rect 103 3337 104 3343
rect 96 3179 104 3337
rect 96 3173 97 3179
rect 103 3173 104 3179
rect 96 3011 104 3173
rect 96 3005 97 3011
rect 103 3005 104 3011
rect 96 2859 104 3005
rect 96 2853 97 2859
rect 103 2853 104 2859
rect 96 2695 104 2853
rect 96 2689 97 2695
rect 103 2689 104 2695
rect 96 2527 104 2689
rect 96 2521 97 2527
rect 103 2521 104 2527
rect 96 2363 104 2521
rect 96 2357 97 2363
rect 103 2357 104 2363
rect 96 2195 104 2357
rect 96 2189 97 2195
rect 103 2189 104 2195
rect 96 2035 104 2189
rect 96 2029 97 2035
rect 103 2029 104 2035
rect 96 1875 104 2029
rect 96 1869 97 1875
rect 103 1869 104 1875
rect 96 1715 104 1869
rect 96 1709 97 1715
rect 103 1709 104 1715
rect 96 1547 104 1709
rect 96 1541 97 1547
rect 103 1541 104 1547
rect 96 1367 104 1541
rect 96 1361 97 1367
rect 103 1361 104 1367
rect 96 1203 104 1361
rect 96 1197 97 1203
rect 103 1197 104 1203
rect 96 1031 104 1197
rect 96 1025 97 1031
rect 103 1025 104 1031
rect 96 859 104 1025
rect 96 853 97 859
rect 103 853 104 859
rect 96 687 104 853
rect 96 681 97 687
rect 103 681 104 687
rect 96 519 104 681
rect 96 513 97 519
rect 103 513 104 519
rect 96 347 104 513
rect 96 341 97 347
rect 103 341 104 347
rect 96 167 104 341
rect 96 161 97 167
rect 103 161 104 167
rect 96 72 104 161
rect 1842 3583 1850 3672
rect 1842 3577 1843 3583
rect 1849 3577 1850 3583
rect 1842 3555 1850 3577
rect 1842 3549 1843 3555
rect 1849 3549 1850 3555
rect 1842 3423 1850 3549
rect 1842 3417 1843 3423
rect 1849 3417 1850 3423
rect 1842 3395 1850 3417
rect 1842 3389 1843 3395
rect 1849 3389 1850 3395
rect 1842 3263 1850 3389
rect 1842 3257 1843 3263
rect 1849 3257 1850 3263
rect 1842 3235 1850 3257
rect 1842 3229 1843 3235
rect 1849 3229 1850 3235
rect 1842 3103 1850 3229
rect 1842 3097 1843 3103
rect 1849 3097 1850 3103
rect 1842 3075 1850 3097
rect 1842 3069 1843 3075
rect 1849 3069 1850 3075
rect 1842 2935 1850 3069
rect 1842 2929 1843 2935
rect 1849 2929 1850 2935
rect 1842 2907 1850 2929
rect 1842 2901 1843 2907
rect 1849 2901 1850 2907
rect 1842 2775 1850 2901
rect 1842 2769 1843 2775
rect 1849 2769 1850 2775
rect 1842 2743 1850 2769
rect 1842 2737 1843 2743
rect 1849 2737 1850 2743
rect 1842 2611 1850 2737
rect 1842 2605 1843 2611
rect 1849 2605 1850 2611
rect 1842 2587 1850 2605
rect 1842 2581 1843 2587
rect 1849 2581 1850 2587
rect 1842 2447 1850 2581
rect 1842 2441 1843 2447
rect 1849 2441 1850 2447
rect 1842 2427 1850 2441
rect 1842 2421 1843 2427
rect 1849 2421 1850 2427
rect 1842 2275 1850 2421
rect 1842 2269 1843 2275
rect 1849 2269 1850 2275
rect 1842 2119 1850 2269
rect 1842 2113 1843 2119
rect 1849 2113 1850 2119
rect 1842 2111 1850 2113
rect 1842 2105 1843 2111
rect 1849 2105 1850 2111
rect 1842 1959 1850 2105
rect 1842 1953 1843 1959
rect 1849 1953 1850 1959
rect 1842 1951 1850 1953
rect 1842 1945 1843 1951
rect 1849 1945 1850 1951
rect 1842 1799 1850 1945
rect 1842 1793 1843 1799
rect 1849 1793 1850 1799
rect 1842 1779 1850 1793
rect 1842 1773 1843 1779
rect 1849 1773 1850 1779
rect 1842 1631 1850 1773
rect 1842 1625 1843 1631
rect 1849 1625 1850 1631
rect 1842 1459 1850 1625
rect 1842 1453 1843 1459
rect 1849 1453 1850 1459
rect 1842 1291 1850 1453
rect 1842 1285 1843 1291
rect 1849 1285 1850 1291
rect 1842 1283 1850 1285
rect 1842 1277 1843 1283
rect 1849 1277 1850 1283
rect 1842 1115 1850 1277
rect 1842 1109 1843 1115
rect 1849 1109 1850 1115
rect 1842 947 1850 1109
rect 1842 941 1843 947
rect 1849 941 1850 947
rect 1842 779 1850 941
rect 1842 773 1843 779
rect 1849 773 1850 779
rect 1842 771 1850 773
rect 1842 765 1843 771
rect 1849 765 1850 771
rect 1842 603 1850 765
rect 1842 597 1843 603
rect 1849 597 1850 603
rect 1842 431 1850 597
rect 1842 425 1843 431
rect 1849 425 1850 431
rect 1842 267 1850 425
rect 1842 261 1843 267
rect 1849 261 1850 267
rect 1842 91 1850 261
rect 1842 85 1843 91
rect 1849 85 1850 91
rect 1842 72 1850 85
rect 1854 3659 1862 3672
rect 1854 3653 1855 3659
rect 1861 3653 1862 3659
rect 1854 3631 1862 3653
rect 1854 3625 1855 3631
rect 1861 3625 1862 3631
rect 1854 3507 1862 3625
rect 1854 3501 1855 3507
rect 1861 3501 1862 3507
rect 1854 3479 1862 3501
rect 1854 3473 1855 3479
rect 1861 3473 1862 3479
rect 1854 3343 1862 3473
rect 1854 3337 1855 3343
rect 1861 3337 1862 3343
rect 1854 3315 1862 3337
rect 1854 3309 1855 3315
rect 1861 3309 1862 3315
rect 1854 3179 1862 3309
rect 1854 3173 1855 3179
rect 1861 3173 1862 3179
rect 1854 3159 1862 3173
rect 1854 3153 1855 3159
rect 1861 3153 1862 3159
rect 1854 3011 1862 3153
rect 1854 3005 1855 3011
rect 1861 3005 1862 3011
rect 1854 2995 1862 3005
rect 1854 2989 1855 2995
rect 1861 2989 1862 2995
rect 1854 2859 1862 2989
rect 1854 2853 1855 2859
rect 1861 2853 1862 2859
rect 1854 2831 1862 2853
rect 1854 2825 1855 2831
rect 1861 2825 1862 2831
rect 1854 2695 1862 2825
rect 1854 2689 1855 2695
rect 1861 2689 1862 2695
rect 1854 2667 1862 2689
rect 1854 2661 1855 2667
rect 1861 2661 1862 2667
rect 1854 2527 1862 2661
rect 1854 2521 1855 2527
rect 1861 2521 1862 2527
rect 1854 2511 1862 2521
rect 1854 2505 1855 2511
rect 1861 2505 1862 2511
rect 1854 2363 1862 2505
rect 1854 2357 1855 2363
rect 1861 2357 1862 2363
rect 1854 2347 1862 2357
rect 1854 2341 1855 2347
rect 1861 2341 1862 2347
rect 1854 2195 1862 2341
rect 1854 2189 1855 2195
rect 1861 2189 1862 2195
rect 1854 2187 1862 2189
rect 1854 2181 1855 2187
rect 1861 2181 1862 2187
rect 1854 2035 1862 2181
rect 1854 2029 1855 2035
rect 1861 2029 1862 2035
rect 1854 1875 1862 2029
rect 1854 1869 1855 1875
rect 1861 1869 1862 1875
rect 1854 1715 1862 1869
rect 1854 1709 1855 1715
rect 1861 1709 1862 1715
rect 1854 1703 1862 1709
rect 1854 1697 1855 1703
rect 1861 1697 1862 1703
rect 1854 1547 1862 1697
rect 1854 1541 1855 1547
rect 1861 1541 1862 1547
rect 1854 1375 1862 1541
rect 1854 1369 1855 1375
rect 1861 1369 1862 1375
rect 1854 1367 1862 1369
rect 1854 1361 1855 1367
rect 1861 1361 1862 1367
rect 1854 1203 1862 1361
rect 1854 1197 1855 1203
rect 1861 1197 1862 1203
rect 1854 1031 1862 1197
rect 1854 1025 1855 1031
rect 1861 1025 1862 1031
rect 1854 859 1862 1025
rect 1854 853 1855 859
rect 1861 853 1862 859
rect 1854 687 1862 853
rect 1854 681 1855 687
rect 1861 681 1862 687
rect 1854 519 1862 681
rect 1854 513 1855 519
rect 1861 513 1862 519
rect 1854 347 1862 513
rect 1854 341 1855 347
rect 1861 341 1862 347
rect 1854 167 1862 341
rect 1854 161 1855 167
rect 1861 161 1862 167
rect 1854 72 1862 161
rect 3618 3555 3626 3672
rect 3618 3549 3619 3555
rect 3625 3549 3626 3555
rect 3618 3395 3626 3549
rect 3618 3389 3619 3395
rect 3625 3389 3626 3395
rect 3618 3235 3626 3389
rect 3618 3229 3619 3235
rect 3625 3229 3626 3235
rect 3618 3075 3626 3229
rect 3618 3069 3619 3075
rect 3625 3069 3626 3075
rect 3618 2907 3626 3069
rect 3618 2901 3619 2907
rect 3625 2901 3626 2907
rect 3618 2743 3626 2901
rect 3618 2737 3619 2743
rect 3625 2737 3626 2743
rect 3618 2587 3626 2737
rect 3618 2581 3619 2587
rect 3625 2581 3626 2587
rect 3618 2427 3626 2581
rect 3618 2421 3619 2427
rect 3625 2421 3626 2427
rect 3618 2111 3626 2421
rect 3618 2105 3619 2111
rect 3625 2105 3626 2111
rect 3618 1951 3626 2105
rect 3618 1945 3619 1951
rect 3625 1945 3626 1951
rect 3618 1779 3626 1945
rect 3618 1773 3619 1779
rect 3625 1773 3626 1779
rect 3618 1283 3626 1773
rect 3618 1277 3619 1283
rect 3625 1277 3626 1283
rect 3618 771 3626 1277
rect 3618 765 3619 771
rect 3625 765 3626 771
rect 3618 72 3626 765
rect 3630 3631 3638 3672
rect 3630 3625 3631 3631
rect 3637 3625 3638 3631
rect 3630 3479 3638 3625
rect 3630 3473 3631 3479
rect 3637 3473 3638 3479
rect 3630 3315 3638 3473
rect 3630 3309 3631 3315
rect 3637 3309 3638 3315
rect 3630 3159 3638 3309
rect 3630 3153 3631 3159
rect 3637 3153 3638 3159
rect 3630 2995 3638 3153
rect 3630 2989 3631 2995
rect 3637 2989 3638 2995
rect 3630 2831 3638 2989
rect 3630 2825 3631 2831
rect 3637 2825 3638 2831
rect 3630 2667 3638 2825
rect 3630 2661 3631 2667
rect 3637 2661 3638 2667
rect 3630 2511 3638 2661
rect 3630 2505 3631 2511
rect 3637 2505 3638 2511
rect 3630 2347 3638 2505
rect 3630 2341 3631 2347
rect 3637 2341 3638 2347
rect 3630 2187 3638 2341
rect 3630 2181 3631 2187
rect 3637 2181 3638 2187
rect 3630 1703 3638 2181
rect 3630 1697 3631 1703
rect 3637 1697 3638 1703
rect 3630 1375 3638 1697
rect 3630 1369 3631 1375
rect 3637 1369 3638 1375
rect 3630 72 3638 1369
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__171
timestamp 1731220556
transform 1 0 3584 0 1 3572
box 7 3 12 24
use welltap_svt  __well_tap__170
timestamp 1731220556
transform 1 0 1864 0 1 3572
box 7 3 12 24
use welltap_svt  __well_tap__169
timestamp 1731220556
transform 1 0 3584 0 -1 3532
box 7 3 12 24
use welltap_svt  __well_tap__168
timestamp 1731220556
transform 1 0 1864 0 -1 3532
box 7 3 12 24
use welltap_svt  __well_tap__167
timestamp 1731220556
transform 1 0 3584 0 1 3420
box 7 3 12 24
use welltap_svt  __well_tap__166
timestamp 1731220556
transform 1 0 1864 0 1 3420
box 7 3 12 24
use welltap_svt  __well_tap__165
timestamp 1731220556
transform 1 0 3584 0 -1 3372
box 7 3 12 24
use welltap_svt  __well_tap__164
timestamp 1731220556
transform 1 0 1864 0 -1 3372
box 7 3 12 24
use welltap_svt  __well_tap__163
timestamp 1731220556
transform 1 0 3584 0 1 3256
box 7 3 12 24
use welltap_svt  __well_tap__162
timestamp 1731220556
transform 1 0 1864 0 1 3256
box 7 3 12 24
use welltap_svt  __well_tap__161
timestamp 1731220556
transform 1 0 3584 0 -1 3212
box 7 3 12 24
use welltap_svt  __well_tap__160
timestamp 1731220556
transform 1 0 1864 0 -1 3212
box 7 3 12 24
use welltap_svt  __well_tap__159
timestamp 1731220556
transform 1 0 3584 0 1 3100
box 7 3 12 24
use welltap_svt  __well_tap__158
timestamp 1731220556
transform 1 0 1864 0 1 3100
box 7 3 12 24
use welltap_svt  __well_tap__157
timestamp 1731220556
transform 1 0 3584 0 -1 3052
box 7 3 12 24
use welltap_svt  __well_tap__156
timestamp 1731220556
transform 1 0 1864 0 -1 3052
box 7 3 12 24
use welltap_svt  __well_tap__155
timestamp 1731220556
transform 1 0 3584 0 1 2936
box 7 3 12 24
use welltap_svt  __well_tap__154
timestamp 1731220556
transform 1 0 1864 0 1 2936
box 7 3 12 24
use welltap_svt  __well_tap__153
timestamp 1731220556
transform 1 0 3584 0 -1 2884
box 7 3 12 24
use welltap_svt  __well_tap__152
timestamp 1731220556
transform 1 0 1864 0 -1 2884
box 7 3 12 24
use welltap_svt  __well_tap__151
timestamp 1731220556
transform 1 0 3584 0 1 2772
box 7 3 12 24
use welltap_svt  __well_tap__150
timestamp 1731220556
transform 1 0 1864 0 1 2772
box 7 3 12 24
use welltap_svt  __well_tap__149
timestamp 1731220556
transform 1 0 3584 0 -1 2720
box 7 3 12 24
use welltap_svt  __well_tap__148
timestamp 1731220556
transform 1 0 1864 0 -1 2720
box 7 3 12 24
use welltap_svt  __well_tap__147
timestamp 1731220556
transform 1 0 3584 0 1 2608
box 7 3 12 24
use welltap_svt  __well_tap__146
timestamp 1731220556
transform 1 0 1864 0 1 2608
box 7 3 12 24
use welltap_svt  __well_tap__145
timestamp 1731220556
transform 1 0 3584 0 -1 2564
box 7 3 12 24
use welltap_svt  __well_tap__144
timestamp 1731220556
transform 1 0 1864 0 -1 2564
box 7 3 12 24
use welltap_svt  __well_tap__143
timestamp 1731220556
transform 1 0 3584 0 1 2452
box 7 3 12 24
use welltap_svt  __well_tap__142
timestamp 1731220556
transform 1 0 1864 0 1 2452
box 7 3 12 24
use welltap_svt  __well_tap__141
timestamp 1731220556
transform 1 0 3584 0 -1 2404
box 7 3 12 24
use welltap_svt  __well_tap__140
timestamp 1731220556
transform 1 0 1864 0 -1 2404
box 7 3 12 24
use welltap_svt  __well_tap__139
timestamp 1731220556
transform 1 0 3584 0 1 2288
box 7 3 12 24
use welltap_svt  __well_tap__138
timestamp 1731220556
transform 1 0 1864 0 1 2288
box 7 3 12 24
use welltap_svt  __well_tap__137
timestamp 1731220556
transform 1 0 3584 0 -1 2248
box 7 3 12 24
use welltap_svt  __well_tap__136
timestamp 1731220556
transform 1 0 1864 0 -1 2248
box 7 3 12 24
use welltap_svt  __well_tap__135
timestamp 1731220556
transform 1 0 3584 0 1 2128
box 7 3 12 24
use welltap_svt  __well_tap__134
timestamp 1731220556
transform 1 0 1864 0 1 2128
box 7 3 12 24
use welltap_svt  __well_tap__133
timestamp 1731220556
transform 1 0 3584 0 -1 2088
box 7 3 12 24
use welltap_svt  __well_tap__132
timestamp 1731220556
transform 1 0 1864 0 -1 2088
box 7 3 12 24
use welltap_svt  __well_tap__131
timestamp 1731220556
transform 1 0 3584 0 1 1972
box 7 3 12 24
use welltap_svt  __well_tap__130
timestamp 1731220556
transform 1 0 1864 0 1 1972
box 7 3 12 24
use welltap_svt  __well_tap__129
timestamp 1731220556
transform 1 0 3584 0 -1 1928
box 7 3 12 24
use welltap_svt  __well_tap__128
timestamp 1731220556
transform 1 0 1864 0 -1 1928
box 7 3 12 24
use welltap_svt  __well_tap__127
timestamp 1731220556
transform 1 0 3584 0 1 1812
box 7 3 12 24
use welltap_svt  __well_tap__126
timestamp 1731220556
transform 1 0 1864 0 1 1812
box 7 3 12 24
use welltap_svt  __well_tap__125
timestamp 1731220556
transform 1 0 3584 0 -1 1756
box 7 3 12 24
use welltap_svt  __well_tap__124
timestamp 1731220556
transform 1 0 1864 0 -1 1756
box 7 3 12 24
use welltap_svt  __well_tap__123
timestamp 1731220556
transform 1 0 3584 0 1 1644
box 7 3 12 24
use welltap_svt  __well_tap__122
timestamp 1731220556
transform 1 0 1864 0 1 1644
box 7 3 12 24
use welltap_svt  __well_tap__121
timestamp 1731220556
transform 1 0 3584 0 -1 1604
box 7 3 12 24
use welltap_svt  __well_tap__120
timestamp 1731220556
transform 1 0 1864 0 -1 1604
box 7 3 12 24
use welltap_svt  __well_tap__119
timestamp 1731220556
transform 1 0 3584 0 1 1484
box 7 3 12 24
use welltap_svt  __well_tap__118
timestamp 1731220556
transform 1 0 1864 0 1 1484
box 7 3 12 24
use welltap_svt  __well_tap__117
timestamp 1731220556
transform 1 0 3584 0 -1 1436
box 7 3 12 24
use welltap_svt  __well_tap__116
timestamp 1731220556
transform 1 0 1864 0 -1 1436
box 7 3 12 24
use welltap_svt  __well_tap__115
timestamp 1731220556
transform 1 0 3584 0 1 1316
box 7 3 12 24
use welltap_svt  __well_tap__114
timestamp 1731220556
transform 1 0 1864 0 1 1316
box 7 3 12 24
use welltap_svt  __well_tap__113
timestamp 1731220556
transform 1 0 3584 0 -1 1260
box 7 3 12 24
use welltap_svt  __well_tap__112
timestamp 1731220556
transform 1 0 1864 0 -1 1260
box 7 3 12 24
use welltap_svt  __well_tap__111
timestamp 1731220556
transform 1 0 3584 0 1 1140
box 7 3 12 24
use welltap_svt  __well_tap__110
timestamp 1731220556
transform 1 0 1864 0 1 1140
box 7 3 12 24
use welltap_svt  __well_tap__109
timestamp 1731220556
transform 1 0 3584 0 -1 1092
box 7 3 12 24
use welltap_svt  __well_tap__108
timestamp 1731220556
transform 1 0 1864 0 -1 1092
box 7 3 12 24
use welltap_svt  __well_tap__107
timestamp 1731220556
transform 1 0 3584 0 1 972
box 7 3 12 24
use welltap_svt  __well_tap__106
timestamp 1731220556
transform 1 0 1864 0 1 972
box 7 3 12 24
use welltap_svt  __well_tap__105
timestamp 1731220556
transform 1 0 3584 0 -1 924
box 7 3 12 24
use welltap_svt  __well_tap__104
timestamp 1731220556
transform 1 0 1864 0 -1 924
box 7 3 12 24
use welltap_svt  __well_tap__103
timestamp 1731220556
transform 1 0 3584 0 1 804
box 7 3 12 24
use welltap_svt  __well_tap__102
timestamp 1731220556
transform 1 0 1864 0 1 804
box 7 3 12 24
use welltap_svt  __well_tap__101
timestamp 1731220556
transform 1 0 3584 0 -1 748
box 7 3 12 24
use welltap_svt  __well_tap__100
timestamp 1731220556
transform 1 0 1864 0 -1 748
box 7 3 12 24
use welltap_svt  __well_tap__99
timestamp 1731220556
transform 1 0 3584 0 1 632
box 7 3 12 24
use welltap_svt  __well_tap__98
timestamp 1731220556
transform 1 0 1864 0 1 632
box 7 3 12 24
use welltap_svt  __well_tap__97
timestamp 1731220556
transform 1 0 3584 0 -1 580
box 7 3 12 24
use welltap_svt  __well_tap__96
timestamp 1731220556
transform 1 0 1864 0 -1 580
box 7 3 12 24
use welltap_svt  __well_tap__95
timestamp 1731220556
transform 1 0 3584 0 1 460
box 7 3 12 24
use welltap_svt  __well_tap__94
timestamp 1731220556
transform 1 0 1864 0 1 460
box 7 3 12 24
use welltap_svt  __well_tap__93
timestamp 1731220556
transform 1 0 3584 0 -1 408
box 7 3 12 24
use welltap_svt  __well_tap__92
timestamp 1731220556
transform 1 0 1864 0 -1 408
box 7 3 12 24
use welltap_svt  __well_tap__91
timestamp 1731220556
transform 1 0 3584 0 1 284
box 7 3 12 24
use welltap_svt  __well_tap__90
timestamp 1731220556
transform 1 0 1864 0 1 284
box 7 3 12 24
use welltap_svt  __well_tap__89
timestamp 1731220556
transform 1 0 3584 0 -1 240
box 7 3 12 24
use welltap_svt  __well_tap__88
timestamp 1731220556
transform 1 0 1864 0 -1 240
box 7 3 12 24
use welltap_svt  __well_tap__87
timestamp 1731220556
transform 1 0 3584 0 1 104
box 7 3 12 24
use welltap_svt  __well_tap__86
timestamp 1731220556
transform 1 0 1864 0 1 104
box 7 3 12 24
use welltap_svt  __well_tap__85
timestamp 1731220556
transform 1 0 1824 0 1 3600
box 7 3 12 24
use welltap_svt  __well_tap__84
timestamp 1731220556
transform 1 0 104 0 1 3600
box 7 3 12 24
use welltap_svt  __well_tap__83
timestamp 1731220556
transform 1 0 1824 0 -1 3560
box 7 3 12 24
use welltap_svt  __well_tap__82
timestamp 1731220556
transform 1 0 104 0 -1 3560
box 7 3 12 24
use welltap_svt  __well_tap__81
timestamp 1731220556
transform 1 0 1824 0 1 3448
box 7 3 12 24
use welltap_svt  __well_tap__80
timestamp 1731220556
transform 1 0 104 0 1 3448
box 7 3 12 24
use welltap_svt  __well_tap__79
timestamp 1731220556
transform 1 0 1824 0 -1 3400
box 7 3 12 24
use welltap_svt  __well_tap__78
timestamp 1731220556
transform 1 0 104 0 -1 3400
box 7 3 12 24
use welltap_svt  __well_tap__77
timestamp 1731220556
transform 1 0 1824 0 1 3284
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220556
transform 1 0 104 0 1 3284
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220556
transform 1 0 1824 0 -1 3240
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220556
transform 1 0 104 0 -1 3240
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220556
transform 1 0 1824 0 1 3120
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220556
transform 1 0 104 0 1 3120
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220556
transform 1 0 1824 0 -1 3080
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220556
transform 1 0 104 0 -1 3080
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220556
transform 1 0 1824 0 1 2952
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220556
transform 1 0 104 0 1 2952
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220556
transform 1 0 1824 0 -1 2912
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220556
transform 1 0 104 0 -1 2912
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220556
transform 1 0 1824 0 1 2800
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220556
transform 1 0 104 0 1 2800
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220556
transform 1 0 1824 0 -1 2752
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220556
transform 1 0 104 0 -1 2752
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220556
transform 1 0 1824 0 1 2636
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220556
transform 1 0 104 0 1 2636
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220556
transform 1 0 1824 0 -1 2588
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220556
transform 1 0 104 0 -1 2588
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220556
transform 1 0 1824 0 1 2468
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220556
transform 1 0 104 0 1 2468
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220556
transform 1 0 1824 0 -1 2424
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220556
transform 1 0 104 0 -1 2424
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220556
transform 1 0 1824 0 1 2304
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220556
transform 1 0 104 0 1 2304
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220556
transform 1 0 1824 0 -1 2252
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220556
transform 1 0 104 0 -1 2252
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220556
transform 1 0 1824 0 1 2136
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220556
transform 1 0 104 0 1 2136
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220556
transform 1 0 1824 0 -1 2096
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220556
transform 1 0 104 0 -1 2096
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220556
transform 1 0 1824 0 1 1976
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220556
transform 1 0 104 0 1 1976
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220556
transform 1 0 1824 0 -1 1936
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220556
transform 1 0 104 0 -1 1936
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220556
transform 1 0 1824 0 1 1816
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220556
transform 1 0 104 0 1 1816
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220556
transform 1 0 1824 0 -1 1776
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220556
transform 1 0 104 0 -1 1776
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220556
transform 1 0 1824 0 1 1656
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220556
transform 1 0 104 0 1 1656
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220556
transform 1 0 1824 0 -1 1608
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220556
transform 1 0 104 0 -1 1608
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220556
transform 1 0 1824 0 1 1488
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220556
transform 1 0 104 0 1 1488
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220556
transform 1 0 1824 0 -1 1436
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220556
transform 1 0 104 0 -1 1436
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220556
transform 1 0 1824 0 1 1308
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220556
transform 1 0 104 0 1 1308
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220556
transform 1 0 1824 0 -1 1268
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220556
transform 1 0 104 0 -1 1268
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220556
transform 1 0 1824 0 1 1144
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220556
transform 1 0 104 0 1 1144
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220556
transform 1 0 1824 0 -1 1092
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220556
transform 1 0 104 0 -1 1092
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220556
transform 1 0 1824 0 1 972
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220556
transform 1 0 104 0 1 972
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220556
transform 1 0 1824 0 -1 924
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220556
transform 1 0 104 0 -1 924
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220556
transform 1 0 1824 0 1 800
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220556
transform 1 0 104 0 1 800
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220556
transform 1 0 1824 0 -1 756
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220556
transform 1 0 104 0 -1 756
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220556
transform 1 0 1824 0 1 628
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220556
transform 1 0 104 0 1 628
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220556
transform 1 0 1824 0 -1 580
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220556
transform 1 0 104 0 -1 580
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220556
transform 1 0 1824 0 1 460
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220556
transform 1 0 104 0 1 460
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220556
transform 1 0 1824 0 -1 408
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220556
transform 1 0 104 0 -1 408
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220556
transform 1 0 1824 0 1 288
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220556
transform 1 0 104 0 1 288
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220556
transform 1 0 1824 0 -1 244
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220556
transform 1 0 104 0 -1 244
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220556
transform 1 0 1824 0 1 108
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220556
transform 1 0 104 0 1 108
box 7 3 12 24
use _0_0std_0_0cells_0_0LATCHINV  tst_5999_6
timestamp 1731220556
transform 1 0 3416 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5998_6
timestamp 1731220556
transform 1 0 3496 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5997_6
timestamp 1731220556
transform 1 0 3496 0 -1 260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5996_6
timestamp 1731220556
transform 1 0 3496 0 1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5995_6
timestamp 1731220556
transform 1 0 3496 0 -1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5994_6
timestamp 1731220556
transform 1 0 3368 0 -1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5993_6
timestamp 1731220556
transform 1 0 3376 0 -1 260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5992_6
timestamp 1731220556
transform 1 0 3232 0 -1 260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5991_6
timestamp 1731220556
transform 1 0 3336 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5990_6
timestamp 1731220556
transform 1 0 3248 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5989_6
timestamp 1731220556
transform 1 0 3160 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5988_6
timestamp 1731220556
transform 1 0 3072 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5987_6
timestamp 1731220556
transform 1 0 2984 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5986_6
timestamp 1731220556
transform 1 0 2896 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5985_6
timestamp 1731220556
transform 1 0 2800 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5984_6
timestamp 1731220556
transform 1 0 2696 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5983_6
timestamp 1731220556
transform 1 0 3080 0 -1 260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5982_6
timestamp 1731220556
transform 1 0 2920 0 -1 260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5981_6
timestamp 1731220556
transform 1 0 2736 0 -1 260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5980_6
timestamp 1731220556
transform 1 0 2536 0 -1 260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5979_6
timestamp 1731220556
transform 1 0 3328 0 1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5978_6
timestamp 1731220556
transform 1 0 3152 0 1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5977_6
timestamp 1731220556
transform 1 0 2984 0 1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5976_6
timestamp 1731220556
transform 1 0 2824 0 1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5975_6
timestamp 1731220556
transform 1 0 2680 0 1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5974_6
timestamp 1731220556
transform 1 0 3224 0 -1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5973_6
timestamp 1731220556
transform 1 0 3080 0 -1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5972_6
timestamp 1731220556
transform 1 0 2952 0 -1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5971_6
timestamp 1731220556
transform 1 0 2832 0 -1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5970_6
timestamp 1731220556
transform 1 0 2728 0 -1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5969_6
timestamp 1731220556
transform 1 0 2632 0 -1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5968_6
timestamp 1731220556
transform 1 0 3296 0 1 440
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5967_6
timestamp 1731220556
transform 1 0 3128 0 1 440
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5966_6
timestamp 1731220556
transform 1 0 2976 0 1 440
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5965_6
timestamp 1731220556
transform 1 0 2544 0 1 440
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5964_6
timestamp 1731220556
transform 1 0 2464 0 1 440
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5963_6
timestamp 1731220556
transform 1 0 2400 0 -1 600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5962_6
timestamp 1731220556
transform 1 0 2480 0 -1 600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5961_6
timestamp 1731220556
transform 1 0 2560 0 -1 600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5960_6
timestamp 1731220556
transform 1 0 2624 0 1 440
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5959_6
timestamp 1731220556
transform 1 0 2840 0 1 440
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5958_6
timestamp 1731220556
transform 1 0 2720 0 1 440
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5957_6
timestamp 1731220556
transform 1 0 2640 0 -1 600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5956_6
timestamp 1731220556
transform 1 0 2736 0 -1 600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5955_6
timestamp 1731220556
transform 1 0 2856 0 -1 600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5954_6
timestamp 1731220556
transform 1 0 3320 0 -1 600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5953_6
timestamp 1731220556
transform 1 0 3152 0 -1 600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5952_6
timestamp 1731220556
transform 1 0 2992 0 -1 600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5951_6
timestamp 1731220556
transform 1 0 2912 0 1 612
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5950_6
timestamp 1731220556
transform 1 0 2784 0 1 612
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5949_6
timestamp 1731220556
transform 1 0 2664 0 1 612
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5948_6
timestamp 1731220556
transform 1 0 3208 0 1 612
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5947_6
timestamp 1731220556
transform 1 0 3056 0 1 612
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5946_6
timestamp 1731220556
transform 1 0 2968 0 -1 768
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5945_6
timestamp 1731220556
transform 1 0 2824 0 -1 768
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5944_6
timestamp 1731220556
transform 1 0 2672 0 -1 768
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5943_6
timestamp 1731220556
transform 1 0 3104 0 -1 768
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5942_6
timestamp 1731220556
transform 1 0 3016 0 1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5941_6
timestamp 1731220556
transform 1 0 2872 0 1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5940_6
timestamp 1731220556
transform 1 0 2720 0 1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5939_6
timestamp 1731220556
transform 1 0 3144 0 1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5938_6
timestamp 1731220556
transform 1 0 3272 0 1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5937_6
timestamp 1731220556
transform 1 0 3392 0 1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5936_6
timestamp 1731220556
transform 1 0 3376 0 -1 768
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5935_6
timestamp 1731220556
transform 1 0 3240 0 -1 768
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5934_6
timestamp 1731220556
transform 1 0 3360 0 1 612
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5933_6
timestamp 1731220556
transform 1 0 3464 0 1 440
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5932_6
timestamp 1731220556
transform 1 0 3488 0 -1 600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5931_6
timestamp 1731220556
transform 1 0 3496 0 1 612
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5930_6
timestamp 1731220556
transform 1 0 3496 0 -1 768
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5929_6
timestamp 1731220556
transform 1 0 3496 0 1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5928_6
timestamp 1731220556
transform 1 0 3496 0 -1 944
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5927_6
timestamp 1731220556
transform 1 0 3496 0 1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5926_6
timestamp 1731220556
transform 1 0 3496 0 -1 1112
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5925_6
timestamp 1731220556
transform 1 0 3496 0 1 1120
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5924_6
timestamp 1731220556
transform 1 0 3496 0 -1 1280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5923_6
timestamp 1731220556
transform 1 0 3392 0 -1 1280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5922_6
timestamp 1731220556
transform 1 0 3264 0 -1 1280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5921_6
timestamp 1731220556
transform 1 0 3176 0 1 1120
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5920_6
timestamp 1731220556
transform 1 0 3344 0 1 1120
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5919_6
timestamp 1731220556
transform 1 0 3336 0 -1 1112
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5918_6
timestamp 1731220556
transform 1 0 3376 0 1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5917_6
timestamp 1731220556
transform 1 0 3392 0 -1 944
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5916_6
timestamp 1731220556
transform 1 0 3264 0 -1 944
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5915_6
timestamp 1731220556
transform 1 0 3136 0 -1 944
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5914_6
timestamp 1731220556
transform 1 0 3008 0 -1 944
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5913_6
timestamp 1731220556
transform 1 0 2872 0 -1 944
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5912_6
timestamp 1731220556
transform 1 0 2728 0 -1 944
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5911_6
timestamp 1731220556
transform 1 0 3232 0 1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5910_6
timestamp 1731220556
transform 1 0 3096 0 1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5909_6
timestamp 1731220556
transform 1 0 2968 0 1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5908_6
timestamp 1731220556
transform 1 0 2840 0 1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5907_6
timestamp 1731220556
transform 1 0 2712 0 1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5906_6
timestamp 1731220556
transform 1 0 3152 0 -1 1112
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5905_6
timestamp 1731220556
transform 1 0 2976 0 -1 1112
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5904_6
timestamp 1731220556
transform 1 0 2816 0 -1 1112
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5903_6
timestamp 1731220556
transform 1 0 2672 0 -1 1112
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5902_6
timestamp 1731220556
transform 1 0 2544 0 -1 1112
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5901_6
timestamp 1731220556
transform 1 0 2560 0 1 1120
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5900_6
timestamp 1731220556
transform 1 0 2704 0 1 1120
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5899_6
timestamp 1731220556
transform 1 0 2856 0 1 1120
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5898_6
timestamp 1731220556
transform 1 0 3016 0 1 1120
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5897_6
timestamp 1731220556
transform 1 0 2872 0 -1 1280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5896_6
timestamp 1731220556
transform 1 0 2728 0 -1 1280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5895_6
timestamp 1731220556
transform 1 0 2576 0 -1 1280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5894_6
timestamp 1731220556
transform 1 0 3008 0 -1 1280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5893_6
timestamp 1731220556
transform 1 0 3136 0 -1 1280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5892_6
timestamp 1731220556
transform 1 0 3056 0 1 1296
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5891_6
timestamp 1731220556
transform 1 0 2944 0 1 1296
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5890_6
timestamp 1731220556
transform 1 0 3168 0 1 1296
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5889_6
timestamp 1731220556
transform 1 0 3280 0 1 1296
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5888_6
timestamp 1731220556
transform 1 0 3400 0 1 1296
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5887_6
timestamp 1731220556
transform 1 0 3496 0 -1 1456
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5886_6
timestamp 1731220556
transform 1 0 3400 0 -1 1456
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5885_6
timestamp 1731220556
transform 1 0 3288 0 -1 1456
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5884_6
timestamp 1731220556
transform 1 0 3176 0 -1 1456
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5883_6
timestamp 1731220556
transform 1 0 3064 0 -1 1456
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5882_6
timestamp 1731220556
transform 1 0 2944 0 -1 1456
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5881_6
timestamp 1731220556
transform 1 0 3336 0 1 1464
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5880_6
timestamp 1731220556
transform 1 0 3216 0 1 1464
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5879_6
timestamp 1731220556
transform 1 0 3104 0 1 1464
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5878_6
timestamp 1731220556
transform 1 0 2992 0 1 1464
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5877_6
timestamp 1731220556
transform 1 0 2872 0 1 1464
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5876_6
timestamp 1731220556
transform 1 0 2752 0 1 1464
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5875_6
timestamp 1731220556
transform 1 0 3336 0 -1 1624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5874_6
timestamp 1731220556
transform 1 0 3152 0 -1 1624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5873_6
timestamp 1731220556
transform 1 0 2976 0 -1 1624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5872_6
timestamp 1731220556
transform 1 0 2816 0 -1 1624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5871_6
timestamp 1731220556
transform 1 0 2664 0 -1 1624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5870_6
timestamp 1731220556
transform 1 0 3184 0 1 1624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5869_6
timestamp 1731220556
transform 1 0 3024 0 1 1624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5868_6
timestamp 1731220556
transform 1 0 2872 0 1 1624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5867_6
timestamp 1731220556
transform 1 0 2728 0 1 1624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5866_6
timestamp 1731220556
transform 1 0 2592 0 1 1624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5865_6
timestamp 1731220556
transform 1 0 2464 0 1 1624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5864_6
timestamp 1731220556
transform 1 0 3264 0 -1 1776
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5863_6
timestamp 1731220556
transform 1 0 3008 0 -1 1776
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5862_6
timestamp 1731220556
transform 1 0 2768 0 -1 1776
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5861_6
timestamp 1731220556
transform 1 0 2544 0 -1 1776
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5860_6
timestamp 1731220556
transform 1 0 2344 0 -1 1776
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5859_6
timestamp 1731220556
transform 1 0 2448 0 1 1792
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5858_6
timestamp 1731220556
transform 1 0 2616 0 1 1792
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5857_6
timestamp 1731220556
transform 1 0 3280 0 1 1792
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5856_6
timestamp 1731220556
transform 1 0 3040 0 1 1792
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5855_6
timestamp 1731220556
transform 1 0 2816 0 1 1792
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5854_6
timestamp 1731220556
transform 1 0 2768 0 -1 1948
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5853_6
timestamp 1731220556
transform 1 0 2640 0 -1 1948
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5852_6
timestamp 1731220556
transform 1 0 2520 0 -1 1948
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5851_6
timestamp 1731220556
transform 1 0 3200 0 -1 1948
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5850_6
timestamp 1731220556
transform 1 0 3048 0 -1 1948
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5849_6
timestamp 1731220556
transform 1 0 2904 0 -1 1948
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5848_6
timestamp 1731220556
transform 1 0 2864 0 1 1952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5847_6
timestamp 1731220556
transform 1 0 2760 0 1 1952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5846_6
timestamp 1731220556
transform 1 0 3176 0 1 1952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5845_6
timestamp 1731220556
transform 1 0 3072 0 1 1952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5844_6
timestamp 1731220556
transform 1 0 2968 0 1 1952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5843_6
timestamp 1731220556
transform 1 0 2960 0 -1 2108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5842_6
timestamp 1731220556
transform 1 0 2848 0 -1 2108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5841_6
timestamp 1731220556
transform 1 0 3072 0 -1 2108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5840_6
timestamp 1731220556
transform 1 0 3184 0 -1 2108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5839_6
timestamp 1731220556
transform 1 0 3296 0 -1 2108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5838_6
timestamp 1731220556
transform 1 0 3408 0 -1 2108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5837_6
timestamp 1731220556
transform 1 0 3496 0 1 2108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5836_6
timestamp 1731220556
transform 1 0 3248 0 1 2108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5835_6
timestamp 1731220556
transform 1 0 3112 0 1 2108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5834_6
timestamp 1731220556
transform 1 0 2976 0 1 2108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5833_6
timestamp 1731220556
transform 1 0 2832 0 1 2108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5832_6
timestamp 1731220556
transform 1 0 3328 0 -1 2268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5831_6
timestamp 1731220556
transform 1 0 3136 0 -1 2268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5830_6
timestamp 1731220556
transform 1 0 2944 0 -1 2268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5829_6
timestamp 1731220556
transform 1 0 2760 0 -1 2268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5828_6
timestamp 1731220556
transform 1 0 3232 0 1 2268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5827_6
timestamp 1731220556
transform 1 0 3072 0 1 2268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5826_6
timestamp 1731220556
transform 1 0 2912 0 1 2268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5825_6
timestamp 1731220556
transform 1 0 2760 0 1 2268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5824_6
timestamp 1731220556
transform 1 0 2608 0 1 2268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5823_6
timestamp 1731220556
transform 1 0 3144 0 -1 2424
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5822_6
timestamp 1731220556
transform 1 0 2960 0 -1 2424
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5821_6
timestamp 1731220556
transform 1 0 2784 0 -1 2424
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5820_6
timestamp 1731220556
transform 1 0 2624 0 -1 2424
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5819_6
timestamp 1731220556
transform 1 0 2640 0 1 2432
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5818_6
timestamp 1731220556
transform 1 0 3048 0 1 2432
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5817_6
timestamp 1731220556
transform 1 0 2904 0 1 2432
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5816_6
timestamp 1731220556
transform 1 0 2768 0 1 2432
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5815_6
timestamp 1731220556
transform 1 0 2688 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5814_6
timestamp 1731220556
transform 1 0 2792 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5813_6
timestamp 1731220556
transform 1 0 2896 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5812_6
timestamp 1731220556
transform 1 0 3008 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5811_6
timestamp 1731220556
transform 1 0 3128 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5810_6
timestamp 1731220556
transform 1 0 3384 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5809_6
timestamp 1731220556
transform 1 0 3256 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5808_6
timestamp 1731220556
transform 1 0 3200 0 1 2432
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5807_6
timestamp 1731220556
transform 1 0 3360 0 1 2432
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5806_6
timestamp 1731220556
transform 1 0 3328 0 -1 2424
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5805_6
timestamp 1731220556
transform 1 0 3400 0 1 2268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5804_6
timestamp 1731220556
transform 1 0 3384 0 1 2108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5803_6
timestamp 1731220556
transform 1 0 3360 0 -1 1948
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5802_6
timestamp 1731220556
transform 1 0 3352 0 1 1624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5801_6
timestamp 1731220556
transform 1 0 3496 0 -1 1624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5800_6
timestamp 1731220556
transform 1 0 3496 0 1 1624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5799_6
timestamp 1731220556
transform 1 0 3496 0 -1 1776
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5798_6
timestamp 1731220556
transform 1 0 3496 0 1 1792
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5797_6
timestamp 1731220556
transform 1 0 3496 0 -1 1948
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5796_6
timestamp 1731220556
transform 1 0 3496 0 -1 2108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5795_6
timestamp 1731220556
transform 1 0 3496 0 -1 2268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5794_6
timestamp 1731220556
transform 1 0 3496 0 -1 2424
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5793_6
timestamp 1731220556
transform 1 0 3496 0 1 2432
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5792_6
timestamp 1731220556
transform 1 0 3496 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5791_6
timestamp 1731220556
transform 1 0 3496 0 1 2588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5790_6
timestamp 1731220556
transform 1 0 3496 0 -1 2740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5789_6
timestamp 1731220556
transform 1 0 3496 0 1 2752
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5788_6
timestamp 1731220556
transform 1 0 3496 0 1 2916
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5787_6
timestamp 1731220556
transform 1 0 3496 0 -1 3072
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5786_6
timestamp 1731220556
transform 1 0 3496 0 -1 3232
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5785_6
timestamp 1731220556
transform 1 0 3496 0 1 3236
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5784_6
timestamp 1731220556
transform 1 0 3496 0 -1 3392
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5783_6
timestamp 1731220556
transform 1 0 3416 0 -1 3392
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5782_6
timestamp 1731220556
transform 1 0 3336 0 -1 3392
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5781_6
timestamp 1731220556
transform 1 0 3248 0 -1 3392
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5780_6
timestamp 1731220556
transform 1 0 3160 0 -1 3392
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5779_6
timestamp 1731220556
transform 1 0 3072 0 -1 3392
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5778_6
timestamp 1731220556
transform 1 0 2984 0 -1 3392
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5777_6
timestamp 1731220556
transform 1 0 2888 0 -1 3392
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5776_6
timestamp 1731220556
transform 1 0 2784 0 -1 3392
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5775_6
timestamp 1731220556
transform 1 0 3112 0 1 3400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5774_6
timestamp 1731220556
transform 1 0 3288 0 1 3400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5773_6
timestamp 1731220556
transform 1 0 3296 0 -1 3552
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5772_6
timestamp 1731220556
transform 1 0 3128 0 -1 3552
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5771_6
timestamp 1731220556
transform 1 0 2968 0 -1 3552
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5770_6
timestamp 1731220556
transform 1 0 3192 0 1 3552
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5769_6
timestamp 1731220556
transform 1 0 3080 0 1 3552
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5768_6
timestamp 1731220556
transform 1 0 2968 0 1 3552
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5767_6
timestamp 1731220556
transform 1 0 2864 0 1 3552
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5766_6
timestamp 1731220556
transform 1 0 2760 0 1 3552
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5765_6
timestamp 1731220556
transform 1 0 2648 0 1 3552
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5764_6
timestamp 1731220556
transform 1 0 2640 0 -1 3552
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5763_6
timestamp 1731220556
transform 1 0 2808 0 -1 3552
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5762_6
timestamp 1731220556
transform 1 0 2944 0 1 3400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5761_6
timestamp 1731220556
transform 1 0 2776 0 1 3400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5760_6
timestamp 1731220556
transform 1 0 2672 0 -1 3392
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5759_6
timestamp 1731220556
transform 1 0 2552 0 -1 3392
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5758_6
timestamp 1731220556
transform 1 0 2752 0 1 3236
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5757_6
timestamp 1731220556
transform 1 0 2992 0 1 3236
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5756_6
timestamp 1731220556
transform 1 0 3240 0 1 3236
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5755_6
timestamp 1731220556
transform 1 0 3304 0 -1 3232
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5754_6
timestamp 1731220556
transform 1 0 3096 0 -1 3232
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5753_6
timestamp 1731220556
transform 1 0 2904 0 -1 3232
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5752_6
timestamp 1731220556
transform 1 0 2720 0 -1 3232
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5751_6
timestamp 1731220556
transform 1 0 2560 0 -1 3232
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5750_6
timestamp 1731220556
transform 1 0 2608 0 1 3080
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5749_6
timestamp 1731220556
transform 1 0 2768 0 1 3080
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5748_6
timestamp 1731220556
transform 1 0 3216 0 1 3080
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5747_6
timestamp 1731220556
transform 1 0 3064 0 1 3080
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5746_6
timestamp 1731220556
transform 1 0 2920 0 1 3080
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5745_6
timestamp 1731220556
transform 1 0 2888 0 -1 3072
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5744_6
timestamp 1731220556
transform 1 0 2696 0 -1 3072
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5743_6
timestamp 1731220556
transform 1 0 3056 0 -1 3072
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5742_6
timestamp 1731220556
transform 1 0 3216 0 -1 3072
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5741_6
timestamp 1731220556
transform 1 0 3368 0 -1 3072
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5740_6
timestamp 1731220556
transform 1 0 3384 0 1 2916
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5739_6
timestamp 1731220556
transform 1 0 3248 0 1 2916
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5738_6
timestamp 1731220556
transform 1 0 3104 0 1 2916
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5737_6
timestamp 1731220556
transform 1 0 2952 0 1 2916
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5736_6
timestamp 1731220556
transform 1 0 2784 0 1 2916
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5735_6
timestamp 1731220556
transform 1 0 2592 0 1 2916
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5734_6
timestamp 1731220556
transform 1 0 3200 0 -1 2904
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5733_6
timestamp 1731220556
transform 1 0 3088 0 -1 2904
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5732_6
timestamp 1731220556
transform 1 0 2976 0 -1 2904
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5731_6
timestamp 1731220556
transform 1 0 2864 0 -1 2904
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5730_6
timestamp 1731220556
transform 1 0 3128 0 1 2752
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5729_6
timestamp 1731220556
transform 1 0 3320 0 1 2752
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5728_6
timestamp 1731220556
transform 1 0 3344 0 -1 2740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5727_6
timestamp 1731220556
transform 1 0 3168 0 -1 2740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5726_6
timestamp 1731220556
transform 1 0 3000 0 -1 2740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5725_6
timestamp 1731220556
transform 1 0 2848 0 -1 2740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5724_6
timestamp 1731220556
transform 1 0 2720 0 -1 2740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5723_6
timestamp 1731220556
transform 1 0 2608 0 -1 2740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5722_6
timestamp 1731220556
transform 1 0 2512 0 -1 2740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5721_6
timestamp 1731220556
transform 1 0 2952 0 1 2752
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5720_6
timestamp 1731220556
transform 1 0 2792 0 1 2752
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5719_6
timestamp 1731220556
transform 1 0 2656 0 1 2752
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5718_6
timestamp 1731220556
transform 1 0 2552 0 1 2752
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5717_6
timestamp 1731220556
transform 1 0 2752 0 -1 2904
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5716_6
timestamp 1731220556
transform 1 0 2648 0 -1 2904
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5715_6
timestamp 1731220556
transform 1 0 2544 0 -1 2904
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5714_6
timestamp 1731220556
transform 1 0 2440 0 -1 2904
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5713_6
timestamp 1731220556
transform 1 0 2344 0 -1 2904
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5712_6
timestamp 1731220556
transform 1 0 2464 0 1 2752
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5711_6
timestamp 1731220556
transform 1 0 2384 0 1 2752
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5710_6
timestamp 1731220556
transform 1 0 2304 0 1 2752
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5709_6
timestamp 1731220556
transform 1 0 2224 0 1 2752
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5708_6
timestamp 1731220556
transform 1 0 2416 0 -1 2740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5707_6
timestamp 1731220556
transform 1 0 2320 0 -1 2740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5706_6
timestamp 1731220556
transform 1 0 2224 0 -1 2740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5705_6
timestamp 1731220556
transform 1 0 2128 0 -1 2740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5704_6
timestamp 1731220556
transform 1 0 2040 0 -1 2740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5703_6
timestamp 1731220556
transform 1 0 2056 0 1 2588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5702_6
timestamp 1731220556
transform 1 0 2280 0 1 2588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5701_6
timestamp 1731220556
transform 1 0 2552 0 1 2588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5700_6
timestamp 1731220556
transform 1 0 3184 0 1 2588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5699_6
timestamp 1731220556
transform 1 0 2856 0 1 2588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5698_6
timestamp 1731220556
transform 1 0 2584 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5697_6
timestamp 1731220556
transform 1 0 2360 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5696_6
timestamp 1731220556
transform 1 0 2256 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5695_6
timestamp 1731220556
transform 1 0 2160 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5694_6
timestamp 1731220556
transform 1 0 2472 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5693_6
timestamp 1731220556
transform 1 0 2520 0 1 2432
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5692_6
timestamp 1731220556
transform 1 0 2408 0 1 2432
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5691_6
timestamp 1731220556
transform 1 0 2304 0 1 2432
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5690_6
timestamp 1731220556
transform 1 0 2208 0 1 2432
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5689_6
timestamp 1731220556
transform 1 0 2120 0 1 2432
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5688_6
timestamp 1731220556
transform 1 0 2472 0 -1 2424
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5687_6
timestamp 1731220556
transform 1 0 2328 0 -1 2424
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5686_6
timestamp 1731220556
transform 1 0 2200 0 -1 2424
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5685_6
timestamp 1731220556
transform 1 0 2080 0 -1 2424
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5684_6
timestamp 1731220556
transform 1 0 1968 0 -1 2424
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5683_6
timestamp 1731220556
transform 1 0 2456 0 1 2268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5682_6
timestamp 1731220556
transform 1 0 2304 0 1 2268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5681_6
timestamp 1731220556
transform 1 0 2152 0 1 2268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5680_6
timestamp 1731220556
transform 1 0 2000 0 1 2268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5679_6
timestamp 1731220556
transform 1 0 1888 0 1 2268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5678_6
timestamp 1731220556
transform 1 0 1888 0 -1 2268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5677_6
timestamp 1731220556
transform 1 0 2024 0 -1 2268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5676_6
timestamp 1731220556
transform 1 0 2568 0 -1 2268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5675_6
timestamp 1731220556
transform 1 0 2384 0 -1 2268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5674_6
timestamp 1731220556
transform 1 0 2200 0 -1 2268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5673_6
timestamp 1731220556
transform 1 0 2200 0 1 2108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5672_6
timestamp 1731220556
transform 1 0 2064 0 1 2108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5671_6
timestamp 1731220556
transform 1 0 1952 0 1 2108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5670_6
timestamp 1731220556
transform 1 0 2352 0 1 2108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5669_6
timestamp 1731220556
transform 1 0 2512 0 1 2108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5668_6
timestamp 1731220556
transform 1 0 2672 0 1 2108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5667_6
timestamp 1731220556
transform 1 0 2616 0 -1 2108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5666_6
timestamp 1731220556
transform 1 0 2496 0 -1 2108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5665_6
timestamp 1731220556
transform 1 0 2384 0 -1 2108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5664_6
timestamp 1731220556
transform 1 0 2280 0 -1 2108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5663_6
timestamp 1731220556
transform 1 0 2736 0 -1 2108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5662_6
timestamp 1731220556
transform 1 0 2656 0 1 1952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5661_6
timestamp 1731220556
transform 1 0 2552 0 1 1952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5660_6
timestamp 1731220556
transform 1 0 2448 0 1 1952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5659_6
timestamp 1731220556
transform 1 0 2352 0 1 1952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5658_6
timestamp 1731220556
transform 1 0 2256 0 1 1952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5657_6
timestamp 1731220556
transform 1 0 2168 0 1 1952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5656_6
timestamp 1731220556
transform 1 0 2400 0 -1 1948
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5655_6
timestamp 1731220556
transform 1 0 2280 0 -1 1948
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5654_6
timestamp 1731220556
transform 1 0 2160 0 -1 1948
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5653_6
timestamp 1731220556
transform 1 0 2048 0 -1 1948
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5652_6
timestamp 1731220556
transform 1 0 1936 0 -1 1948
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5651_6
timestamp 1731220556
transform 1 0 2312 0 1 1792
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5650_6
timestamp 1731220556
transform 1 0 2192 0 1 1792
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5649_6
timestamp 1731220556
transform 1 0 2080 0 1 1792
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5648_6
timestamp 1731220556
transform 1 0 1968 0 1 1792
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5647_6
timestamp 1731220556
transform 1 0 1888 0 1 1792
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5646_6
timestamp 1731220556
transform 1 0 1736 0 -1 1796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5645_6
timestamp 1731220556
transform 1 0 1656 0 -1 1796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5644_6
timestamp 1731220556
transform 1 0 1552 0 -1 1796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5643_6
timestamp 1731220556
transform 1 0 1888 0 -1 1776
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5642_6
timestamp 1731220556
transform 1 0 2016 0 -1 1776
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5641_6
timestamp 1731220556
transform 1 0 2176 0 -1 1776
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5640_6
timestamp 1731220556
transform 1 0 2336 0 1 1624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5639_6
timestamp 1731220556
transform 1 0 2216 0 1 1624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5638_6
timestamp 1731220556
transform 1 0 2096 0 1 1624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5637_6
timestamp 1731220556
transform 1 0 1976 0 1 1624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5636_6
timestamp 1731220556
transform 1 0 1888 0 1 1624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5635_6
timestamp 1731220556
transform 1 0 1920 0 -1 1624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5634_6
timestamp 1731220556
transform 1 0 2016 0 -1 1624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5633_6
timestamp 1731220556
transform 1 0 2128 0 -1 1624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5632_6
timestamp 1731220556
transform 1 0 2256 0 -1 1624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5631_6
timestamp 1731220556
transform 1 0 2384 0 -1 1624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5630_6
timestamp 1731220556
transform 1 0 2520 0 -1 1624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5629_6
timestamp 1731220556
transform 1 0 2624 0 1 1464
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5628_6
timestamp 1731220556
transform 1 0 2496 0 1 1464
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5627_6
timestamp 1731220556
transform 1 0 2368 0 1 1464
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5626_6
timestamp 1731220556
transform 1 0 2240 0 1 1464
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5625_6
timestamp 1731220556
transform 1 0 2120 0 1 1464
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5624_6
timestamp 1731220556
transform 1 0 2240 0 -1 1456
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5623_6
timestamp 1731220556
transform 1 0 2336 0 -1 1456
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5622_6
timestamp 1731220556
transform 1 0 2448 0 -1 1456
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5621_6
timestamp 1731220556
transform 1 0 2568 0 -1 1456
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5620_6
timestamp 1731220556
transform 1 0 2696 0 -1 1456
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5619_6
timestamp 1731220556
transform 1 0 2824 0 -1 1456
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5618_6
timestamp 1731220556
transform 1 0 2832 0 1 1296
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5617_6
timestamp 1731220556
transform 1 0 2720 0 1 1296
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5616_6
timestamp 1731220556
transform 1 0 2600 0 1 1296
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5615_6
timestamp 1731220556
transform 1 0 2488 0 1 1296
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5614_6
timestamp 1731220556
transform 1 0 2384 0 1 1296
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5613_6
timestamp 1731220556
transform 1 0 2248 0 -1 1280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5612_6
timestamp 1731220556
transform 1 0 2416 0 -1 1280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5611_6
timestamp 1731220556
transform 1 0 2432 0 1 1120
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5610_6
timestamp 1731220556
transform 1 0 2312 0 1 1120
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5609_6
timestamp 1731220556
transform 1 0 2200 0 1 1120
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5608_6
timestamp 1731220556
transform 1 0 2328 0 -1 1112
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5607_6
timestamp 1731220556
transform 1 0 2432 0 -1 1112
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5606_6
timestamp 1731220556
transform 1 0 2584 0 1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5605_6
timestamp 1731220556
transform 1 0 2456 0 1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5604_6
timestamp 1731220556
transform 1 0 2336 0 1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5603_6
timestamp 1731220556
transform 1 0 2216 0 1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5602_6
timestamp 1731220556
transform 1 0 2112 0 1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5601_6
timestamp 1731220556
transform 1 0 2016 0 1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5600_6
timestamp 1731220556
transform 1 0 2224 0 -1 1112
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5599_6
timestamp 1731220556
transform 1 0 2128 0 -1 1112
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5598_6
timestamp 1731220556
transform 1 0 2040 0 -1 1112
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5597_6
timestamp 1731220556
transform 1 0 1960 0 -1 1112
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5596_6
timestamp 1731220556
transform 1 0 1888 0 1 1120
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5595_6
timestamp 1731220556
transform 1 0 1976 0 1 1120
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5594_6
timestamp 1731220556
transform 1 0 2088 0 1 1120
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5593_6
timestamp 1731220556
transform 1 0 2064 0 -1 1280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5592_6
timestamp 1731220556
transform 1 0 1888 0 -1 1280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5591_6
timestamp 1731220556
transform 1 0 1736 0 -1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5590_6
timestamp 1731220556
transform 1 0 1640 0 -1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5589_6
timestamp 1731220556
transform 1 0 1624 0 1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5588_6
timestamp 1731220556
transform 1 0 1528 0 -1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5587_6
timestamp 1731220556
transform 1 0 1416 0 -1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5586_6
timestamp 1731220556
transform 1 0 1296 0 -1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5585_6
timestamp 1731220556
transform 1 0 1176 0 -1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5584_6
timestamp 1731220556
transform 1 0 1496 0 1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5583_6
timestamp 1731220556
transform 1 0 1360 0 1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5582_6
timestamp 1731220556
transform 1 0 1224 0 1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5581_6
timestamp 1731220556
transform 1 0 1080 0 1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5580_6
timestamp 1731220556
transform 1 0 1736 0 1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5579_6
timestamp 1731220556
transform 1 0 1736 0 -1 1456
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5578_6
timestamp 1731220556
transform 1 0 1632 0 -1 1456
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5577_6
timestamp 1731220556
transform 1 0 1504 0 -1 1456
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5576_6
timestamp 1731220556
transform 1 0 1376 0 -1 1456
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5575_6
timestamp 1731220556
transform 1 0 1240 0 -1 1456
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5574_6
timestamp 1731220556
transform 1 0 1104 0 -1 1456
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5573_6
timestamp 1731220556
transform 1 0 1560 0 1 1468
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5572_6
timestamp 1731220556
transform 1 0 1440 0 1 1468
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5571_6
timestamp 1731220556
transform 1 0 1328 0 1 1468
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5570_6
timestamp 1731220556
transform 1 0 1216 0 1 1468
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5569_6
timestamp 1731220556
transform 1 0 1096 0 1 1468
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5568_6
timestamp 1731220556
transform 1 0 968 0 1 1468
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5567_6
timestamp 1731220556
transform 1 0 1296 0 -1 1628
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5566_6
timestamp 1731220556
transform 1 0 1192 0 -1 1628
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5565_6
timestamp 1731220556
transform 1 0 1088 0 -1 1628
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5564_6
timestamp 1731220556
transform 1 0 992 0 -1 1628
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5563_6
timestamp 1731220556
transform 1 0 896 0 -1 1628
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5562_6
timestamp 1731220556
transform 1 0 792 0 -1 1628
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5561_6
timestamp 1731220556
transform 1 0 808 0 1 1636
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5560_6
timestamp 1731220556
transform 1 0 912 0 1 1636
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5559_6
timestamp 1731220556
transform 1 0 1008 0 1 1636
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5558_6
timestamp 1731220556
transform 1 0 1304 0 1 1636
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5557_6
timestamp 1731220556
transform 1 0 1200 0 1 1636
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5556_6
timestamp 1731220556
transform 1 0 1104 0 1 1636
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5555_6
timestamp 1731220556
transform 1 0 984 0 -1 1796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5554_6
timestamp 1731220556
transform 1 0 1120 0 -1 1796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5553_6
timestamp 1731220556
transform 1 0 1456 0 -1 1796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5552_6
timestamp 1731220556
transform 1 0 1352 0 -1 1796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5551_6
timestamp 1731220556
transform 1 0 1240 0 -1 1796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5550_6
timestamp 1731220556
transform 1 0 1192 0 1 1796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5549_6
timestamp 1731220556
transform 1 0 1040 0 1 1796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5548_6
timestamp 1731220556
transform 1 0 1328 0 1 1796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5547_6
timestamp 1731220556
transform 1 0 1456 0 1 1796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5546_6
timestamp 1731220556
transform 1 0 1584 0 1 1796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5545_6
timestamp 1731220556
transform 1 0 1712 0 1 1796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5544_6
timestamp 1731220556
transform 1 0 1616 0 -1 1956
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5543_6
timestamp 1731220556
transform 1 0 1480 0 -1 1956
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5542_6
timestamp 1731220556
transform 1 0 1352 0 -1 1956
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5541_6
timestamp 1731220556
transform 1 0 1224 0 -1 1956
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5540_6
timestamp 1731220556
transform 1 0 1088 0 -1 1956
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5539_6
timestamp 1731220556
transform 1 0 1448 0 1 1956
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5538_6
timestamp 1731220556
transform 1 0 1304 0 1 1956
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5537_6
timestamp 1731220556
transform 1 0 1168 0 1 1956
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5536_6
timestamp 1731220556
transform 1 0 1032 0 1 1956
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5535_6
timestamp 1731220556
transform 1 0 1336 0 -1 2116
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5534_6
timestamp 1731220556
transform 1 0 1232 0 -1 2116
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5533_6
timestamp 1731220556
transform 1 0 1136 0 -1 2116
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5532_6
timestamp 1731220556
transform 1 0 1040 0 -1 2116
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5531_6
timestamp 1731220556
transform 1 0 1248 0 1 2116
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5530_6
timestamp 1731220556
transform 1 0 1136 0 1 2116
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5529_6
timestamp 1731220556
transform 1 0 1024 0 1 2116
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5528_6
timestamp 1731220556
transform 1 0 1000 0 -1 2272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5527_6
timestamp 1731220556
transform 1 0 904 0 -1 2272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5526_6
timestamp 1731220556
transform 1 0 808 0 -1 2272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5525_6
timestamp 1731220556
transform 1 0 784 0 1 2284
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5524_6
timestamp 1731220556
transform 1 0 896 0 1 2284
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5523_6
timestamp 1731220556
transform 1 0 1008 0 1 2284
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5522_6
timestamp 1731220556
transform 1 0 1040 0 -1 2444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5521_6
timestamp 1731220556
transform 1 0 912 0 -1 2444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5520_6
timestamp 1731220556
transform 1 0 776 0 -1 2444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5519_6
timestamp 1731220556
transform 1 0 632 0 -1 2444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5518_6
timestamp 1731220556
transform 1 0 1000 0 1 2448
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5517_6
timestamp 1731220556
transform 1 0 864 0 1 2448
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5516_6
timestamp 1731220556
transform 1 0 720 0 1 2448
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5515_6
timestamp 1731220556
transform 1 0 576 0 1 2448
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5514_6
timestamp 1731220556
transform 1 0 920 0 -1 2608
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5513_6
timestamp 1731220556
transform 1 0 784 0 -1 2608
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5512_6
timestamp 1731220556
transform 1 0 632 0 -1 2608
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5511_6
timestamp 1731220556
transform 1 0 472 0 -1 2608
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5510_6
timestamp 1731220556
transform 1 0 528 0 1 2616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5509_6
timestamp 1731220556
transform 1 0 656 0 1 2616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5508_6
timestamp 1731220556
transform 1 0 776 0 1 2616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5507_6
timestamp 1731220556
transform 1 0 680 0 -1 2772
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5506_6
timestamp 1731220556
transform 1 0 560 0 -1 2772
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5505_6
timestamp 1731220556
transform 1 0 432 0 -1 2772
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5504_6
timestamp 1731220556
transform 1 0 528 0 1 2780
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5503_6
timestamp 1731220556
transform 1 0 656 0 1 2780
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5502_6
timestamp 1731220556
transform 1 0 784 0 1 2780
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5501_6
timestamp 1731220556
transform 1 0 888 0 -1 2932
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5500_6
timestamp 1731220556
transform 1 0 744 0 -1 2932
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5499_6
timestamp 1731220556
transform 1 0 600 0 -1 2932
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5498_6
timestamp 1731220556
transform 1 0 464 0 -1 2932
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5497_6
timestamp 1731220556
transform 1 0 968 0 1 2932
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5496_6
timestamp 1731220556
transform 1 0 792 0 1 2932
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5495_6
timestamp 1731220556
transform 1 0 616 0 1 2932
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5494_6
timestamp 1731220556
transform 1 0 456 0 1 2932
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5493_6
timestamp 1731220556
transform 1 0 312 0 1 2932
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5492_6
timestamp 1731220556
transform 1 0 192 0 1 2932
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5491_6
timestamp 1731220556
transform 1 0 344 0 -1 2932
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5490_6
timestamp 1731220556
transform 1 0 240 0 -1 2932
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5489_6
timestamp 1731220556
transform 1 0 136 0 1 2780
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5488_6
timestamp 1731220556
transform 1 0 264 0 1 2780
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5487_6
timestamp 1731220556
transform 1 0 392 0 1 2780
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5486_6
timestamp 1731220556
transform 1 0 288 0 -1 2772
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5485_6
timestamp 1731220556
transform 1 0 136 0 -1 2772
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5484_6
timestamp 1731220556
transform 1 0 128 0 1 2616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5483_6
timestamp 1731220556
transform 1 0 392 0 1 2616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5482_6
timestamp 1731220556
transform 1 0 248 0 1 2616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5481_6
timestamp 1731220556
transform 1 0 136 0 -1 2608
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5480_6
timestamp 1731220556
transform 1 0 304 0 -1 2608
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5479_6
timestamp 1731220556
transform 1 0 280 0 1 2448
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5478_6
timestamp 1731220556
transform 1 0 128 0 1 2448
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5477_6
timestamp 1731220556
transform 1 0 432 0 1 2448
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5476_6
timestamp 1731220556
transform 1 0 488 0 -1 2444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5475_6
timestamp 1731220556
transform 1 0 344 0 -1 2444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5474_6
timestamp 1731220556
transform 1 0 192 0 -1 2444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5473_6
timestamp 1731220556
transform 1 0 208 0 1 2284
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5472_6
timestamp 1731220556
transform 1 0 312 0 1 2284
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5471_6
timestamp 1731220556
transform 1 0 424 0 1 2284
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5470_6
timestamp 1731220556
transform 1 0 664 0 1 2284
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5469_6
timestamp 1731220556
transform 1 0 544 0 1 2284
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5468_6
timestamp 1731220556
transform 1 0 496 0 -1 2272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5467_6
timestamp 1731220556
transform 1 0 400 0 -1 2272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5466_6
timestamp 1731220556
transform 1 0 304 0 -1 2272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5465_6
timestamp 1731220556
transform 1 0 600 0 -1 2272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5464_6
timestamp 1731220556
transform 1 0 704 0 -1 2272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5463_6
timestamp 1731220556
transform 1 0 712 0 1 2116
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5462_6
timestamp 1731220556
transform 1 0 608 0 1 2116
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5461_6
timestamp 1731220556
transform 1 0 504 0 1 2116
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5460_6
timestamp 1731220556
transform 1 0 400 0 1 2116
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5459_6
timestamp 1731220556
transform 1 0 304 0 1 2116
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5458_6
timestamp 1731220556
transform 1 0 616 0 -1 2116
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5457_6
timestamp 1731220556
transform 1 0 504 0 -1 2116
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5456_6
timestamp 1731220556
transform 1 0 392 0 -1 2116
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5455_6
timestamp 1731220556
transform 1 0 272 0 -1 2116
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5454_6
timestamp 1731220556
transform 1 0 608 0 1 1956
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5453_6
timestamp 1731220556
transform 1 0 456 0 1 1956
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5452_6
timestamp 1731220556
transform 1 0 312 0 1 1956
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5451_6
timestamp 1731220556
transform 1 0 168 0 1 1956
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5450_6
timestamp 1731220556
transform 1 0 456 0 -1 1956
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5449_6
timestamp 1731220556
transform 1 0 288 0 -1 1956
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5448_6
timestamp 1731220556
transform 1 0 128 0 -1 1956
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5447_6
timestamp 1731220556
transform 1 0 128 0 1 1796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5446_6
timestamp 1731220556
transform 1 0 304 0 1 1796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5445_6
timestamp 1731220556
transform 1 0 504 0 1 1796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5444_6
timestamp 1731220556
transform 1 0 304 0 -1 1796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5443_6
timestamp 1731220556
transform 1 0 128 0 -1 1796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5442_6
timestamp 1731220556
transform 1 0 128 0 1 1636
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5441_6
timestamp 1731220556
transform 1 0 224 0 1 1636
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5440_6
timestamp 1731220556
transform 1 0 352 0 1 1636
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5439_6
timestamp 1731220556
transform 1 0 472 0 1 1636
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5438_6
timestamp 1731220556
transform 1 0 432 0 -1 1628
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5437_6
timestamp 1731220556
transform 1 0 304 0 -1 1628
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5436_6
timestamp 1731220556
transform 1 0 168 0 -1 1628
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5435_6
timestamp 1731220556
transform 1 0 224 0 1 1468
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5434_6
timestamp 1731220556
transform 1 0 328 0 1 1468
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5433_6
timestamp 1731220556
transform 1 0 448 0 1 1468
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5432_6
timestamp 1731220556
transform 1 0 576 0 1 1468
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5431_6
timestamp 1731220556
transform 1 0 504 0 -1 1456
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5430_6
timestamp 1731220556
transform 1 0 376 0 -1 1456
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5429_6
timestamp 1731220556
transform 1 0 272 0 -1 1456
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5428_6
timestamp 1731220556
transform 1 0 648 0 -1 1456
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5427_6
timestamp 1731220556
transform 1 0 768 0 1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5426_6
timestamp 1731220556
transform 1 0 608 0 1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5425_6
timestamp 1731220556
transform 1 0 456 0 1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5424_6
timestamp 1731220556
transform 1 0 320 0 1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5423_6
timestamp 1731220556
transform 1 0 328 0 -1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5422_6
timestamp 1731220556
transform 1 0 600 0 -1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5421_6
timestamp 1731220556
transform 1 0 456 0 -1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5420_6
timestamp 1731220556
transform 1 0 368 0 1 1124
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5419_6
timestamp 1731220556
transform 1 0 392 0 -1 1112
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5418_6
timestamp 1731220556
transform 1 0 248 0 -1 1112
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5417_6
timestamp 1731220556
transform 1 0 256 0 1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5416_6
timestamp 1731220556
transform 1 0 408 0 1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5415_6
timestamp 1731220556
transform 1 0 728 0 -1 944
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5414_6
timestamp 1731220556
transform 1 0 872 0 1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5413_6
timestamp 1731220556
transform 1 0 720 0 1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5412_6
timestamp 1731220556
transform 1 0 568 0 1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5411_6
timestamp 1731220556
transform 1 0 528 0 -1 1112
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5410_6
timestamp 1731220556
transform 1 0 776 0 -1 1112
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5409_6
timestamp 1731220556
transform 1 0 656 0 -1 1112
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5408_6
timestamp 1731220556
transform 1 0 600 0 1 1124
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5407_6
timestamp 1731220556
transform 1 0 488 0 1 1124
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5406_6
timestamp 1731220556
transform 1 0 704 0 1 1124
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5405_6
timestamp 1731220556
transform 1 0 744 0 -1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5404_6
timestamp 1731220556
transform 1 0 896 0 -1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5403_6
timestamp 1731220556
transform 1 0 1040 0 -1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5402_6
timestamp 1731220556
transform 1 0 984 0 1 1124
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5401_6
timestamp 1731220556
transform 1 0 896 0 1 1124
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5400_6
timestamp 1731220556
transform 1 0 800 0 1 1124
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5399_6
timestamp 1731220556
transform 1 0 1080 0 1 1124
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5398_6
timestamp 1731220556
transform 1 0 1272 0 1 1124
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5397_6
timestamp 1731220556
transform 1 0 1176 0 1 1124
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5396_6
timestamp 1731220556
transform 1 0 1088 0 -1 1112
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5395_6
timestamp 1731220556
transform 1 0 992 0 -1 1112
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5394_6
timestamp 1731220556
transform 1 0 888 0 -1 1112
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5393_6
timestamp 1731220556
transform 1 0 1184 0 -1 1112
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5392_6
timestamp 1731220556
transform 1 0 1288 0 -1 1112
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5391_6
timestamp 1731220556
transform 1 0 1392 0 -1 1112
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5390_6
timestamp 1731220556
transform 1 0 1624 0 1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5389_6
timestamp 1731220556
transform 1 0 1504 0 1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5388_6
timestamp 1731220556
transform 1 0 1384 0 1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5387_6
timestamp 1731220556
transform 1 0 1264 0 1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5386_6
timestamp 1731220556
transform 1 0 1144 0 1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5385_6
timestamp 1731220556
transform 1 0 1016 0 1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5384_6
timestamp 1731220556
transform 1 0 1448 0 -1 944
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5383_6
timestamp 1731220556
transform 1 0 1328 0 -1 944
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5382_6
timestamp 1731220556
transform 1 0 1216 0 -1 944
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5381_6
timestamp 1731220556
transform 1 0 1104 0 -1 944
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5380_6
timestamp 1731220556
transform 1 0 984 0 -1 944
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5379_6
timestamp 1731220556
transform 1 0 856 0 -1 944
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5378_6
timestamp 1731220556
transform 1 0 1552 0 1 780
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5377_6
timestamp 1731220556
transform 1 0 1344 0 1 780
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5376_6
timestamp 1731220556
transform 1 0 1152 0 1 780
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5375_6
timestamp 1731220556
transform 1 0 976 0 1 780
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5374_6
timestamp 1731220556
transform 1 0 824 0 1 780
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5373_6
timestamp 1731220556
transform 1 0 696 0 1 780
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5372_6
timestamp 1731220556
transform 1 0 848 0 -1 776
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5371_6
timestamp 1731220556
transform 1 0 976 0 -1 776
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5370_6
timestamp 1731220556
transform 1 0 1104 0 -1 776
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5369_6
timestamp 1731220556
transform 1 0 1360 0 -1 776
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5368_6
timestamp 1731220556
transform 1 0 1232 0 -1 776
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5367_6
timestamp 1731220556
transform 1 0 1112 0 1 608
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5366_6
timestamp 1731220556
transform 1 0 1240 0 1 608
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5365_6
timestamp 1731220556
transform 1 0 1368 0 1 608
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5364_6
timestamp 1731220556
transform 1 0 1296 0 -1 600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5363_6
timestamp 1731220556
transform 1 0 1192 0 -1 600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5362_6
timestamp 1731220556
transform 1 0 1392 0 -1 600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5361_6
timestamp 1731220556
transform 1 0 1456 0 1 440
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5360_6
timestamp 1731220556
transform 1 0 1688 0 1 440
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5359_6
timestamp 1731220556
transform 1 0 1704 0 -1 600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5358_6
timestamp 1731220556
transform 1 0 1600 0 -1 600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5357_6
timestamp 1731220556
transform 1 0 1496 0 -1 600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5356_6
timestamp 1731220556
transform 1 0 1488 0 1 608
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5355_6
timestamp 1731220556
transform 1 0 1736 0 1 608
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5354_6
timestamp 1731220556
transform 1 0 1616 0 1 608
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5353_6
timestamp 1731220556
transform 1 0 1488 0 -1 776
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5352_6
timestamp 1731220556
transform 1 0 1624 0 -1 776
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5351_6
timestamp 1731220556
transform 1 0 1736 0 -1 776
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5350_6
timestamp 1731220556
transform 1 0 1736 0 1 780
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5349_6
timestamp 1731220556
transform 1 0 1888 0 1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5348_6
timestamp 1731220556
transform 1 0 1888 0 -1 944
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5347_6
timestamp 1731220556
transform 1 0 1976 0 -1 944
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5346_6
timestamp 1731220556
transform 1 0 2104 0 -1 944
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5345_6
timestamp 1731220556
transform 1 0 2576 0 -1 944
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5344_6
timestamp 1731220556
transform 1 0 2416 0 -1 944
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5343_6
timestamp 1731220556
transform 1 0 2256 0 -1 944
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5342_6
timestamp 1731220556
transform 1 0 2200 0 1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5341_6
timestamp 1731220556
transform 1 0 2024 0 1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5340_6
timestamp 1731220556
transform 1 0 2376 0 1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5339_6
timestamp 1731220556
transform 1 0 2552 0 1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5338_6
timestamp 1731220556
transform 1 0 2512 0 -1 768
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5337_6
timestamp 1731220556
transform 1 0 2352 0 -1 768
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5336_6
timestamp 1731220556
transform 1 0 2184 0 -1 768
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5335_6
timestamp 1731220556
transform 1 0 2016 0 -1 768
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5334_6
timestamp 1731220556
transform 1 0 2080 0 1 612
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5333_6
timestamp 1731220556
transform 1 0 2160 0 1 612
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5332_6
timestamp 1731220556
transform 1 0 2248 0 1 612
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5331_6
timestamp 1731220556
transform 1 0 2552 0 1 612
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5330_6
timestamp 1731220556
transform 1 0 2448 0 1 612
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5329_6
timestamp 1731220556
transform 1 0 2344 0 1 612
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5328_6
timestamp 1731220556
transform 1 0 2320 0 -1 600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5327_6
timestamp 1731220556
transform 1 0 2240 0 -1 600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5326_6
timestamp 1731220556
transform 1 0 2160 0 -1 600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5325_6
timestamp 1731220556
transform 1 0 2384 0 1 440
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5324_6
timestamp 1731220556
transform 1 0 2304 0 1 440
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5323_6
timestamp 1731220556
transform 1 0 2224 0 1 440
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5322_6
timestamp 1731220556
transform 1 0 2144 0 1 440
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5321_6
timestamp 1731220556
transform 1 0 2552 0 -1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5320_6
timestamp 1731220556
transform 1 0 2472 0 -1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5319_6
timestamp 1731220556
transform 1 0 2392 0 -1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5318_6
timestamp 1731220556
transform 1 0 2312 0 -1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5317_6
timestamp 1731220556
transform 1 0 2232 0 -1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5316_6
timestamp 1731220556
transform 1 0 2152 0 -1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5315_6
timestamp 1731220556
transform 1 0 2552 0 1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5314_6
timestamp 1731220556
transform 1 0 2432 0 1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5313_6
timestamp 1731220556
transform 1 0 2320 0 1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5312_6
timestamp 1731220556
transform 1 0 2208 0 1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5311_6
timestamp 1731220556
transform 1 0 2104 0 1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5310_6
timestamp 1731220556
transform 1 0 2016 0 1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5309_6
timestamp 1731220556
transform 1 0 2064 0 -1 260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5308_6
timestamp 1731220556
transform 1 0 2312 0 -1 260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5307_6
timestamp 1731220556
transform 1 0 2592 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5306_6
timestamp 1731220556
transform 1 0 2488 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5305_6
timestamp 1731220556
transform 1 0 2384 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5304_6
timestamp 1731220556
transform 1 0 2288 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5303_6
timestamp 1731220556
transform 1 0 2208 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5302_6
timestamp 1731220556
transform 1 0 2128 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5301_6
timestamp 1731220556
transform 1 0 2048 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5300_6
timestamp 1731220556
transform 1 0 1968 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5299_6
timestamp 1731220556
transform 1 0 1888 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5298_6
timestamp 1731220556
transform 1 0 1736 0 -1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5297_6
timestamp 1731220556
transform 1 0 1640 0 -1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5296_6
timestamp 1731220556
transform 1 0 1520 0 -1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5295_6
timestamp 1731220556
transform 1 0 1736 0 1 268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5294_6
timestamp 1731220556
transform 1 0 1608 0 1 268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5293_6
timestamp 1731220556
transform 1 0 1464 0 1 268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5292_6
timestamp 1731220556
transform 1 0 1312 0 1 268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5291_6
timestamp 1731220556
transform 1 0 1408 0 -1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5290_6
timestamp 1731220556
transform 1 0 1544 0 -1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5289_6
timestamp 1731220556
transform 1 0 1680 0 -1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5288_6
timestamp 1731220556
transform 1 0 1568 0 1 440
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5287_6
timestamp 1731220556
transform 1 0 1344 0 1 440
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5286_6
timestamp 1731220556
transform 1 0 1224 0 1 440
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5285_6
timestamp 1731220556
transform 1 0 1096 0 1 440
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5284_6
timestamp 1731220556
transform 1 0 1272 0 -1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5283_6
timestamp 1731220556
transform 1 0 1136 0 -1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5282_6
timestamp 1731220556
transform 1 0 992 0 -1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5281_6
timestamp 1731220556
transform 1 0 984 0 1 268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5280_6
timestamp 1731220556
transform 1 0 1152 0 1 268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5279_6
timestamp 1731220556
transform 1 0 1400 0 -1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5278_6
timestamp 1731220556
transform 1 0 1280 0 -1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5277_6
timestamp 1731220556
transform 1 0 1168 0 -1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5276_6
timestamp 1731220556
transform 1 0 1056 0 -1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5275_6
timestamp 1731220556
transform 1 0 936 0 -1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5274_6
timestamp 1731220556
transform 1 0 1528 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5273_6
timestamp 1731220556
transform 1 0 1448 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5272_6
timestamp 1731220556
transform 1 0 1368 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5271_6
timestamp 1731220556
transform 1 0 1288 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5270_6
timestamp 1731220556
transform 1 0 1208 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5269_6
timestamp 1731220556
transform 1 0 1128 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5268_6
timestamp 1731220556
transform 1 0 1048 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5267_6
timestamp 1731220556
transform 1 0 968 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5266_6
timestamp 1731220556
transform 1 0 888 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5265_6
timestamp 1731220556
transform 1 0 808 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5264_6
timestamp 1731220556
transform 1 0 728 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5263_6
timestamp 1731220556
transform 1 0 648 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5262_6
timestamp 1731220556
transform 1 0 568 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5261_6
timestamp 1731220556
transform 1 0 488 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5260_6
timestamp 1731220556
transform 1 0 408 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5259_6
timestamp 1731220556
transform 1 0 328 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5258_6
timestamp 1731220556
transform 1 0 248 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5257_6
timestamp 1731220556
transform 1 0 816 0 -1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5256_6
timestamp 1731220556
transform 1 0 704 0 -1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5255_6
timestamp 1731220556
transform 1 0 592 0 -1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5254_6
timestamp 1731220556
transform 1 0 488 0 -1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5253_6
timestamp 1731220556
transform 1 0 384 0 -1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5252_6
timestamp 1731220556
transform 1 0 296 0 -1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5251_6
timestamp 1731220556
transform 1 0 808 0 1 268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5250_6
timestamp 1731220556
transform 1 0 624 0 1 268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5249_6
timestamp 1731220556
transform 1 0 440 0 1 268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5248_6
timestamp 1731220556
transform 1 0 264 0 1 268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5247_6
timestamp 1731220556
transform 1 0 128 0 1 268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5246_6
timestamp 1731220556
transform 1 0 128 0 -1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5245_6
timestamp 1731220556
transform 1 0 216 0 -1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5244_6
timestamp 1731220556
transform 1 0 352 0 -1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5243_6
timestamp 1731220556
transform 1 0 504 0 -1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5242_6
timestamp 1731220556
transform 1 0 832 0 -1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5241_6
timestamp 1731220556
transform 1 0 672 0 -1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5240_6
timestamp 1731220556
transform 1 0 560 0 1 440
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5239_6
timestamp 1731220556
transform 1 0 448 0 1 440
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5238_6
timestamp 1731220556
transform 1 0 352 0 1 440
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5237_6
timestamp 1731220556
transform 1 0 688 0 1 440
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5236_6
timestamp 1731220556
transform 1 0 824 0 1 440
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5235_6
timestamp 1731220556
transform 1 0 960 0 1 440
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5234_6
timestamp 1731220556
transform 1 0 1088 0 -1 600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5233_6
timestamp 1731220556
transform 1 0 984 0 -1 600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5232_6
timestamp 1731220556
transform 1 0 880 0 -1 600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5231_6
timestamp 1731220556
transform 1 0 776 0 -1 600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5230_6
timestamp 1731220556
transform 1 0 680 0 -1 600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5229_6
timestamp 1731220556
transform 1 0 592 0 -1 600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5228_6
timestamp 1731220556
transform 1 0 976 0 1 608
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5227_6
timestamp 1731220556
transform 1 0 840 0 1 608
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5226_6
timestamp 1731220556
transform 1 0 704 0 1 608
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5225_6
timestamp 1731220556
transform 1 0 576 0 1 608
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5224_6
timestamp 1731220556
transform 1 0 464 0 1 608
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5223_6
timestamp 1731220556
transform 1 0 368 0 1 608
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5222_6
timestamp 1731220556
transform 1 0 728 0 -1 776
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5221_6
timestamp 1731220556
transform 1 0 608 0 -1 776
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5220_6
timestamp 1731220556
transform 1 0 496 0 -1 776
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5219_6
timestamp 1731220556
transform 1 0 384 0 -1 776
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5218_6
timestamp 1731220556
transform 1 0 280 0 -1 776
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5217_6
timestamp 1731220556
transform 1 0 192 0 -1 776
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5216_6
timestamp 1731220556
transform 1 0 584 0 1 780
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5215_6
timestamp 1731220556
transform 1 0 480 0 1 780
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5214_6
timestamp 1731220556
transform 1 0 376 0 1 780
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5213_6
timestamp 1731220556
transform 1 0 288 0 1 780
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5212_6
timestamp 1731220556
transform 1 0 208 0 1 780
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5211_6
timestamp 1731220556
transform 1 0 128 0 1 780
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5210_6
timestamp 1731220556
transform 1 0 592 0 -1 944
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5209_6
timestamp 1731220556
transform 1 0 456 0 -1 944
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5208_6
timestamp 1731220556
transform 1 0 328 0 -1 944
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5207_6
timestamp 1731220556
transform 1 0 208 0 -1 944
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5206_6
timestamp 1731220556
transform 1 0 128 0 -1 944
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5205_6
timestamp 1731220556
transform 1 0 128 0 1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5204_6
timestamp 1731220556
transform 1 0 128 0 -1 1112
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5203_6
timestamp 1731220556
transform 1 0 128 0 1 1124
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5202_6
timestamp 1731220556
transform 1 0 240 0 1 1124
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5201_6
timestamp 1731220556
transform 1 0 208 0 -1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5200_6
timestamp 1731220556
transform 1 0 128 0 -1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5199_6
timestamp 1731220556
transform 1 0 208 0 1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5198_6
timestamp 1731220556
transform 1 0 928 0 1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5197_6
timestamp 1731220556
transform 1 0 952 0 -1 1456
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5196_6
timestamp 1731220556
transform 1 0 800 0 -1 1456
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5195_6
timestamp 1731220556
transform 1 0 840 0 1 1468
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5194_6
timestamp 1731220556
transform 1 0 704 0 1 1468
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5193_6
timestamp 1731220556
transform 1 0 680 0 -1 1628
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5192_6
timestamp 1731220556
transform 1 0 560 0 -1 1628
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5191_6
timestamp 1731220556
transform 1 0 592 0 1 1636
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5190_6
timestamp 1731220556
transform 1 0 704 0 1 1636
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5189_6
timestamp 1731220556
transform 1 0 680 0 -1 1796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5188_6
timestamp 1731220556
transform 1 0 496 0 -1 1796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5187_6
timestamp 1731220556
transform 1 0 840 0 -1 1796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5186_6
timestamp 1731220556
transform 1 0 696 0 1 1796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5185_6
timestamp 1731220556
transform 1 0 872 0 1 1796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5184_6
timestamp 1731220556
transform 1 0 944 0 -1 1956
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5183_6
timestamp 1731220556
transform 1 0 792 0 -1 1956
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5182_6
timestamp 1731220556
transform 1 0 624 0 -1 1956
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5181_6
timestamp 1731220556
transform 1 0 752 0 1 1956
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5180_6
timestamp 1731220556
transform 1 0 896 0 1 1956
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5179_6
timestamp 1731220556
transform 1 0 944 0 -1 2116
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5178_6
timestamp 1731220556
transform 1 0 840 0 -1 2116
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5177_6
timestamp 1731220556
transform 1 0 728 0 -1 2116
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5176_6
timestamp 1731220556
transform 1 0 816 0 1 2116
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5175_6
timestamp 1731220556
transform 1 0 920 0 1 2116
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5174_6
timestamp 1731220556
transform 1 0 1096 0 -1 2272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5173_6
timestamp 1731220556
transform 1 0 1296 0 -1 2272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5172_6
timestamp 1731220556
transform 1 0 1192 0 -1 2272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5171_6
timestamp 1731220556
transform 1 0 1120 0 1 2284
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5170_6
timestamp 1731220556
transform 1 0 1232 0 1 2284
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5169_6
timestamp 1731220556
transform 1 0 1352 0 1 2284
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5168_6
timestamp 1731220556
transform 1 0 1440 0 -1 2444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5167_6
timestamp 1731220556
transform 1 0 1304 0 -1 2444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5166_6
timestamp 1731220556
transform 1 0 1168 0 -1 2444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5165_6
timestamp 1731220556
transform 1 0 1128 0 1 2448
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5164_6
timestamp 1731220556
transform 1 0 1256 0 1 2448
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5163_6
timestamp 1731220556
transform 1 0 1384 0 1 2448
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5162_6
timestamp 1731220556
transform 1 0 1520 0 1 2448
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5161_6
timestamp 1731220556
transform 1 0 1520 0 -1 2608
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5160_6
timestamp 1731220556
transform 1 0 1400 0 -1 2608
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5159_6
timestamp 1731220556
transform 1 0 1288 0 -1 2608
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5158_6
timestamp 1731220556
transform 1 0 1168 0 -1 2608
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5157_6
timestamp 1731220556
transform 1 0 1048 0 -1 2608
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5156_6
timestamp 1731220556
transform 1 0 1408 0 1 2616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5155_6
timestamp 1731220556
transform 1 0 1304 0 1 2616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5154_6
timestamp 1731220556
transform 1 0 1200 0 1 2616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5153_6
timestamp 1731220556
transform 1 0 1104 0 1 2616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5152_6
timestamp 1731220556
transform 1 0 1000 0 1 2616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5151_6
timestamp 1731220556
transform 1 0 888 0 1 2616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5150_6
timestamp 1731220556
transform 1 0 1296 0 -1 2772
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5149_6
timestamp 1731220556
transform 1 0 1192 0 -1 2772
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5148_6
timestamp 1731220556
transform 1 0 1096 0 -1 2772
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5147_6
timestamp 1731220556
transform 1 0 1000 0 -1 2772
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5146_6
timestamp 1731220556
transform 1 0 896 0 -1 2772
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5145_6
timestamp 1731220556
transform 1 0 792 0 -1 2772
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5144_6
timestamp 1731220556
transform 1 0 904 0 1 2780
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5143_6
timestamp 1731220556
transform 1 0 1024 0 1 2780
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5142_6
timestamp 1731220556
transform 1 0 1136 0 1 2780
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5141_6
timestamp 1731220556
transform 1 0 1376 0 1 2780
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5140_6
timestamp 1731220556
transform 1 0 1256 0 1 2780
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5139_6
timestamp 1731220556
transform 1 0 1152 0 -1 2932
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5138_6
timestamp 1731220556
transform 1 0 1024 0 -1 2932
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5137_6
timestamp 1731220556
transform 1 0 1272 0 -1 2932
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5136_6
timestamp 1731220556
transform 1 0 1632 0 -1 2932
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5135_6
timestamp 1731220556
transform 1 0 1512 0 -1 2932
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5134_6
timestamp 1731220556
transform 1 0 1392 0 -1 2932
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5133_6
timestamp 1731220556
transform 1 0 1296 0 1 2932
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5132_6
timestamp 1731220556
transform 1 0 1136 0 1 2932
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5131_6
timestamp 1731220556
transform 1 0 1448 0 1 2932
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5130_6
timestamp 1731220556
transform 1 0 1600 0 1 2932
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5129_6
timestamp 1731220556
transform 1 0 1736 0 1 2932
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5128_6
timestamp 1731220556
transform 1 0 1888 0 1 2916
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5127_6
timestamp 1731220556
transform 1 0 2128 0 1 2916
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5126_6
timestamp 1731220556
transform 1 0 2376 0 1 2916
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5125_6
timestamp 1731220556
transform 1 0 2480 0 -1 3072
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5124_6
timestamp 1731220556
transform 1 0 2240 0 -1 3072
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5123_6
timestamp 1731220556
transform 1 0 1984 0 -1 3072
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5122_6
timestamp 1731220556
transform 1 0 2256 0 1 3080
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5121_6
timestamp 1731220556
transform 1 0 2440 0 1 3080
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5120_6
timestamp 1731220556
transform 1 0 2408 0 -1 3232
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5119_6
timestamp 1731220556
transform 1 0 2272 0 -1 3232
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5118_6
timestamp 1731220556
transform 1 0 2192 0 1 3236
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5117_6
timestamp 1731220556
transform 1 0 2536 0 1 3236
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5116_6
timestamp 1731220556
transform 1 0 2352 0 1 3236
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5115_6
timestamp 1731220556
transform 1 0 2280 0 -1 3392
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5114_6
timestamp 1731220556
transform 1 0 2424 0 -1 3392
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5113_6
timestamp 1731220556
transform 1 0 2616 0 1 3400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5112_6
timestamp 1731220556
transform 1 0 2464 0 1 3400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5111_6
timestamp 1731220556
transform 1 0 2320 0 1 3400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5110_6
timestamp 1731220556
transform 1 0 2296 0 -1 3552
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5109_6
timestamp 1731220556
transform 1 0 2472 0 -1 3552
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5108_6
timestamp 1731220556
transform 1 0 2536 0 1 3552
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5107_6
timestamp 1731220556
transform 1 0 2416 0 1 3552
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5106_6
timestamp 1731220556
transform 1 0 2304 0 1 3552
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5105_6
timestamp 1731220556
transform 1 0 2192 0 1 3552
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5104_6
timestamp 1731220556
transform 1 0 2088 0 1 3552
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5103_6
timestamp 1731220556
transform 1 0 1992 0 1 3552
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5102_6
timestamp 1731220556
transform 1 0 1912 0 1 3552
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5101_6
timestamp 1731220556
transform 1 0 1936 0 -1 3552
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5100_6
timestamp 1731220556
transform 1 0 2120 0 -1 3552
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_599_6
timestamp 1731220556
transform 1 0 2184 0 1 3400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_598_6
timestamp 1731220556
transform 1 0 2064 0 1 3400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_597_6
timestamp 1731220556
transform 1 0 1944 0 1 3400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_596_6
timestamp 1731220556
transform 1 0 1968 0 -1 3392
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_595_6
timestamp 1731220556
transform 1 0 2128 0 -1 3392
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_594_6
timestamp 1731220556
transform 1 0 2056 0 1 3236
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_593_6
timestamp 1731220556
transform 1 0 1920 0 1 3236
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_592_6
timestamp 1731220556
transform 1 0 1888 0 -1 3232
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_591_6
timestamp 1731220556
transform 1 0 2000 0 -1 3232
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_590_6
timestamp 1731220556
transform 1 0 2136 0 -1 3232
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_589_6
timestamp 1731220556
transform 1 0 2064 0 1 3080
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_588_6
timestamp 1731220556
transform 1 0 1888 0 1 3080
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_587_6
timestamp 1731220556
transform 1 0 1736 0 -1 3100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_586_6
timestamp 1731220556
transform 1 0 1656 0 -1 3100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_585_6
timestamp 1731220556
transform 1 0 1576 0 -1 3100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_584_6
timestamp 1731220556
transform 1 0 1496 0 -1 3100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_583_6
timestamp 1731220556
transform 1 0 1416 0 -1 3100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_582_6
timestamp 1731220556
transform 1 0 1336 0 -1 3100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_581_6
timestamp 1731220556
transform 1 0 1256 0 -1 3100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_580_6
timestamp 1731220556
transform 1 0 1176 0 -1 3100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_579_6
timestamp 1731220556
transform 1 0 1096 0 -1 3100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_578_6
timestamp 1731220556
transform 1 0 1016 0 -1 3100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_577_6
timestamp 1731220556
transform 1 0 936 0 -1 3100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_576_6
timestamp 1731220556
transform 1 0 1720 0 1 3100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_575_6
timestamp 1731220556
transform 1 0 1600 0 1 3100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_574_6
timestamp 1731220556
transform 1 0 1480 0 1 3100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_573_6
timestamp 1731220556
transform 1 0 1368 0 1 3100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_572_6
timestamp 1731220556
transform 1 0 1256 0 1 3100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_571_6
timestamp 1731220556
transform 1 0 1568 0 -1 3260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_570_6
timestamp 1731220556
transform 1 0 1440 0 -1 3260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_569_6
timestamp 1731220556
transform 1 0 1312 0 -1 3260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_568_6
timestamp 1731220556
transform 1 0 1184 0 -1 3260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_567_6
timestamp 1731220556
transform 1 0 1176 0 1 3264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_566_6
timestamp 1731220556
transform 1 0 1312 0 1 3264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_565_6
timestamp 1731220556
transform 1 0 1448 0 1 3264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_564_6
timestamp 1731220556
transform 1 0 1408 0 -1 3420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_563_6
timestamp 1731220556
transform 1 0 1280 0 -1 3420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_562_6
timestamp 1731220556
transform 1 0 1152 0 -1 3420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_561_6
timestamp 1731220556
transform 1 0 1168 0 1 3428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_560_6
timestamp 1731220556
transform 1 0 1288 0 1 3428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_559_6
timestamp 1731220556
transform 1 0 1408 0 1 3428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_558_6
timestamp 1731220556
transform 1 0 1432 0 -1 3580
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_557_6
timestamp 1731220556
transform 1 0 1312 0 -1 3580
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_556_6
timestamp 1731220556
transform 1 0 1200 0 -1 3580
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_555_6
timestamp 1731220556
transform 1 0 1320 0 1 3580
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_554_6
timestamp 1731220556
transform 1 0 1136 0 1 3580
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_553_6
timestamp 1731220556
transform 1 0 960 0 1 3580
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_552_6
timestamp 1731220556
transform 1 0 856 0 -1 3580
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_551_6
timestamp 1731220556
transform 1 0 976 0 -1 3580
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_550_6
timestamp 1731220556
transform 1 0 1088 0 -1 3580
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_549_6
timestamp 1731220556
transform 1 0 1056 0 1 3428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_548_6
timestamp 1731220556
transform 1 0 936 0 1 3428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_547_6
timestamp 1731220556
transform 1 0 808 0 1 3428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_546_6
timestamp 1731220556
transform 1 0 768 0 -1 3420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_545_6
timestamp 1731220556
transform 1 0 896 0 -1 3420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_544_6
timestamp 1731220556
transform 1 0 1024 0 -1 3420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_543_6
timestamp 1731220556
transform 1 0 1040 0 1 3264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_542_6
timestamp 1731220556
transform 1 0 904 0 1 3264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_541_6
timestamp 1731220556
transform 1 0 776 0 1 3264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_540_6
timestamp 1731220556
transform 1 0 800 0 -1 3260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_539_6
timestamp 1731220556
transform 1 0 928 0 -1 3260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_538_6
timestamp 1731220556
transform 1 0 1056 0 -1 3260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_537_6
timestamp 1731220556
transform 1 0 1144 0 1 3100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_536_6
timestamp 1731220556
transform 1 0 1024 0 1 3100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_535_6
timestamp 1731220556
transform 1 0 912 0 1 3100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_534_6
timestamp 1731220556
transform 1 0 800 0 1 3100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_533_6
timestamp 1731220556
transform 1 0 696 0 1 3100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_532_6
timestamp 1731220556
transform 1 0 608 0 1 3100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_531_6
timestamp 1731220556
transform 1 0 528 0 1 3100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_530_6
timestamp 1731220556
transform 1 0 448 0 1 3100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_529_6
timestamp 1731220556
transform 1 0 368 0 1 3100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_528_6
timestamp 1731220556
transform 1 0 680 0 -1 3260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_527_6
timestamp 1731220556
transform 1 0 568 0 -1 3260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_526_6
timestamp 1731220556
transform 1 0 464 0 -1 3260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_525_6
timestamp 1731220556
transform 1 0 376 0 -1 3260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_524_6
timestamp 1731220556
transform 1 0 640 0 1 3264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_523_6
timestamp 1731220556
transform 1 0 504 0 1 3264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_522_6
timestamp 1731220556
transform 1 0 376 0 1 3264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_521_6
timestamp 1731220556
transform 1 0 256 0 1 3264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_520_6
timestamp 1731220556
transform 1 0 632 0 -1 3420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_519_6
timestamp 1731220556
transform 1 0 496 0 -1 3420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_518_6
timestamp 1731220556
transform 1 0 368 0 -1 3420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_517_6
timestamp 1731220556
transform 1 0 240 0 -1 3420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_516_6
timestamp 1731220556
transform 1 0 128 0 -1 3420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_515_6
timestamp 1731220556
transform 1 0 152 0 1 3428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_514_6
timestamp 1731220556
transform 1 0 272 0 1 3428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_513_6
timestamp 1731220556
transform 1 0 400 0 1 3428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_512_6
timestamp 1731220556
transform 1 0 536 0 1 3428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_511_6
timestamp 1731220556
transform 1 0 672 0 1 3428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_510_6
timestamp 1731220556
transform 1 0 728 0 -1 3580
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_59_6
timestamp 1731220556
transform 1 0 600 0 -1 3580
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_58_6
timestamp 1731220556
transform 1 0 472 0 -1 3580
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_57_6
timestamp 1731220556
transform 1 0 352 0 -1 3580
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_56_6
timestamp 1731220556
transform 1 0 232 0 -1 3580
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_55_6
timestamp 1731220556
transform 1 0 792 0 1 3580
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_54_6
timestamp 1731220556
transform 1 0 632 0 1 3580
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_53_6
timestamp 1731220556
transform 1 0 480 0 1 3580
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_52_6
timestamp 1731220556
transform 1 0 336 0 1 3580
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_51_6
timestamp 1731220556
transform 1 0 208 0 1 3580
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_50_6
timestamp 1731220556
transform 1 0 128 0 1 3580
box 8 4 70 72
<< end >>
