magic
tech sky130l
timestamp 1730592110
<< m1 >>
rect 18 41 23 46
rect 26 41 31 46
rect 42 44 47 45
rect 34 40 38 44
rect 42 41 43 44
rect 46 41 47 44
rect 42 40 47 41
rect 16 32 20 33
rect 16 29 17 32
rect 24 32 28 33
rect 27 29 28 32
rect 16 28 20 29
rect 10 6 13 15
rect 17 12 20 28
rect 16 8 20 12
rect 34 6 37 40
rect 42 24 45 40
<< m2c >>
rect 43 41 46 44
rect 17 29 20 32
rect 24 29 27 32
rect 10 3 13 6
rect 34 3 37 6
<< m2 >>
rect 42 44 47 45
rect 42 41 43 44
rect 46 41 47 44
rect 42 40 47 41
rect 16 32 28 33
rect 16 29 17 32
rect 20 30 24 32
rect 20 29 21 30
rect 16 28 21 29
rect 23 29 24 30
rect 27 29 28 32
rect 23 28 28 29
rect 9 6 14 7
rect 33 6 38 7
rect 9 3 10 6
rect 13 3 34 6
rect 37 3 38 6
rect 9 2 14 3
rect 33 2 38 3
<< labels >>
rlabel m1 s 22 42 23 45 6 A
port 1 nsew signal input
rlabel m1 s 19 42 22 45 6 A
port 1 nsew signal input
rlabel m1 s 18 41 23 42 6 A
port 1 nsew signal input
rlabel m1 s 18 42 19 45 6 A
port 1 nsew signal input
rlabel m1 s 18 45 23 46 6 A
port 1 nsew signal input
rlabel m1 s 30 42 31 45 6 B
port 2 nsew signal input
rlabel m1 s 27 42 30 45 6 B
port 2 nsew signal input
rlabel m1 s 26 42 27 45 6 B
port 2 nsew signal input
rlabel m1 s 26 45 31 46 6 B
port 2 nsew signal input
rlabel m1 s 26 41 31 42 6 B
port 2 nsew signal input
rlabel m2 s 33 6 38 7 6 Y
port 3 nsew signal output
rlabel m2 s 27 29 28 32 6 Y
port 3 nsew signal output
rlabel m2 s 24 29 27 32 6 Y
port 3 nsew signal output
rlabel m2 s 23 29 24 30 6 Y
port 3 nsew signal output
rlabel m2 s 23 28 28 29 6 Y
port 3 nsew signal output
rlabel m2 s 20 29 21 30 6 Y
port 3 nsew signal output
rlabel m2 s 20 30 24 32 6 Y
port 3 nsew signal output
rlabel m2 s 17 29 20 32 6 Y
port 3 nsew signal output
rlabel m2 s 16 28 21 29 6 Y
port 3 nsew signal output
rlabel m2 s 16 29 17 32 6 Y
port 3 nsew signal output
rlabel m2 s 16 32 28 33 6 Y
port 3 nsew signal output
rlabel m2 s 10 3 13 6 6 Y
port 3 nsew signal output
rlabel m2 s 9 2 14 3 6 Y
port 3 nsew signal output
rlabel m2 s 9 3 10 6 6 Y
port 3 nsew signal output
rlabel m2 s 9 6 14 7 6 Y
port 3 nsew signal output
rlabel m2c s 24 29 27 32 6 Y
port 3 nsew signal output
rlabel m2c s 17 29 20 32 6 Y
port 3 nsew signal output
rlabel m2c s 10 3 13 6 6 Y
port 3 nsew signal output
rlabel m1 s 42 24 45 25 6 Y
port 3 nsew signal output
rlabel m1 s 42 25 45 28 6 Y
port 3 nsew signal output
rlabel m1 s 42 28 45 40 6 Y
port 3 nsew signal output
rlabel m1 s 27 29 28 32 6 Y
port 3 nsew signal output
rlabel m1 s 24 29 27 32 6 Y
port 3 nsew signal output
rlabel m1 s 24 32 28 33 6 Y
port 3 nsew signal output
rlabel m1 s 17 12 20 28 6 Y
port 3 nsew signal output
rlabel m1 s 17 29 20 32 6 Y
port 3 nsew signal output
rlabel m1 s 16 8 20 12 6 Y
port 3 nsew signal output
rlabel m1 s 16 28 20 29 6 Y
port 3 nsew signal output
rlabel m1 s 16 29 17 32 6 Y
port 3 nsew signal output
rlabel m1 s 16 32 20 33 6 Y
port 3 nsew signal output
rlabel m1 s 10 3 13 6 6 Y
port 3 nsew signal output
rlabel m1 s 10 6 13 11 6 Y
port 3 nsew signal output
rlabel m1 s 10 11 13 14 6 Y
port 3 nsew signal output
rlabel m1 s 10 14 13 15 6 Y
port 3 nsew signal output
rlabel m2 s 46 41 47 44 6 Vdd
port 4 nsew power input
rlabel m2 s 43 41 46 44 6 Vdd
port 4 nsew power input
rlabel m2 s 42 40 47 41 6 Vdd
port 4 nsew power input
rlabel m2 s 42 41 43 44 6 Vdd
port 4 nsew power input
rlabel m2 s 42 44 47 45 6 Vdd
port 4 nsew power input
rlabel m2c s 43 41 46 44 6 Vdd
port 4 nsew power input
rlabel m1 s 46 41 47 44 6 Vdd
port 4 nsew power input
rlabel m1 s 43 41 46 44 6 Vdd
port 4 nsew power input
rlabel m1 s 42 40 47 41 6 Vdd
port 4 nsew power input
rlabel m1 s 42 41 43 44 6 Vdd
port 4 nsew power input
rlabel m1 s 42 44 47 45 6 Vdd
port 4 nsew power input
rlabel m2 s 33 2 38 3 6 GND
port 5 nsew ground input
rlabel m2 s 37 3 38 6 6 GND
port 5 nsew ground input
rlabel m2 s 34 3 37 6 6 GND
port 5 nsew ground input
rlabel m2 s 13 3 34 6 6 GND
port 5 nsew ground input
rlabel m2c s 34 3 37 6 6 GND
port 5 nsew ground input
rlabel m1 s 34 3 37 6 6 GND
port 5 nsew ground input
rlabel m1 s 34 6 37 12 6 GND
port 5 nsew ground input
rlabel m1 s 34 12 37 15 6 GND
port 5 nsew ground input
rlabel m1 s 34 15 37 40 6 GND
port 5 nsew ground input
rlabel m1 s 34 40 38 44 6 GND
port 5 nsew ground input
<< properties >>
string LEFsite CoreSite
string LEFclass CORE
string FIXED_BBOX 0 0 56 48
string LEFsymmetry X Y
string LEFview TRUE
<< end >>
