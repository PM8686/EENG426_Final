magic
tech TSMC180
timestamp 1734143975
<< ndiffusion >>
rect 3 21 12 22
rect 3 18 6 21
rect 9 18 12 21
rect 3 17 12 18
rect 14 21 20 22
rect 14 18 15 21
rect 18 18 20 21
rect 14 17 20 18
rect 22 21 28 22
rect 22 18 23 21
rect 26 18 28 21
rect 22 17 28 18
rect 30 20 51 22
rect 30 18 36 20
rect 38 18 51 20
rect 30 17 51 18
<< ndcontact >>
rect 6 18 9 21
rect 15 18 18 21
rect 23 18 26 21
rect 36 18 38 20
<< ntransistor >>
rect 12 17 14 22
rect 20 17 22 22
rect 28 17 30 22
<< pdiffusion >>
rect 3 44 12 53
rect 3 41 5 44
rect 8 41 12 44
rect 3 38 12 41
rect 14 38 20 53
rect 22 46 26 53
rect 22 43 28 46
rect 22 41 24 43
rect 26 41 28 43
rect 22 38 28 41
rect 30 43 51 46
rect 30 41 36 43
rect 38 41 51 43
rect 30 38 51 41
<< pdcontact >>
rect 5 41 8 44
rect 24 41 26 43
rect 36 41 38 43
<< ptransistor >>
rect 12 38 14 53
rect 20 38 22 53
rect 28 38 30 46
<< polysilicon >>
rect 19 66 23 67
rect 19 64 20 66
rect 22 64 23 66
rect 19 63 23 64
rect 11 59 15 60
rect 11 57 12 59
rect 14 57 15 59
rect 11 56 15 57
rect 12 53 14 56
rect 20 53 22 63
rect 28 46 30 49
rect 12 22 14 38
rect 20 22 22 38
rect 28 22 30 38
rect 12 14 14 17
rect 20 14 22 17
rect 28 9 30 17
rect 26 8 31 9
rect 26 5 27 8
rect 30 5 31 8
rect 26 4 31 5
<< polycontact >>
rect 20 64 22 66
rect 12 57 14 59
rect 27 5 30 8
<< m1 >>
rect 19 66 23 67
rect 19 64 20 66
rect 22 64 23 66
rect 19 63 23 64
rect 11 59 15 60
rect 11 57 12 59
rect 14 57 15 59
rect 11 56 15 57
rect 4 44 9 45
rect 24 44 27 60
rect 4 41 5 44
rect 8 41 9 44
rect 4 40 9 41
rect 23 43 27 44
rect 23 41 24 43
rect 26 41 27 43
rect 23 40 27 41
rect 35 43 39 44
rect 35 41 36 43
rect 38 41 39 43
rect 35 40 39 41
rect 5 34 8 40
rect 4 33 9 34
rect 4 30 5 33
rect 8 30 9 33
rect 4 29 9 30
rect 14 33 19 34
rect 14 30 15 33
rect 18 30 19 33
rect 14 29 19 30
rect 15 22 18 29
rect 5 21 10 22
rect 5 18 6 21
rect 9 18 10 21
rect 5 17 10 18
rect 14 21 19 22
rect 14 18 15 21
rect 18 18 19 21
rect 14 17 19 18
rect 22 21 27 22
rect 36 21 39 40
rect 22 18 23 21
rect 26 18 27 21
rect 22 17 27 18
rect 35 20 39 21
rect 35 18 36 20
rect 38 18 39 20
rect 35 17 39 18
rect 15 9 18 17
rect 15 8 20 9
rect 15 5 16 8
rect 19 5 20 8
rect 15 4 20 5
rect 26 8 31 9
rect 26 5 27 8
rect 30 5 31 8
rect 26 4 31 5
<< m2c >>
rect 5 30 8 33
rect 15 30 18 33
rect 6 18 9 21
rect 23 18 26 21
rect 16 5 19 8
rect 27 5 30 8
<< m2 >>
rect 4 33 19 34
rect 4 30 5 33
rect 8 30 15 33
rect 18 30 19 33
rect 4 29 19 30
rect 5 21 27 22
rect 5 18 6 21
rect 9 18 23 21
rect 26 18 27 21
rect 5 17 27 18
rect 15 8 31 9
rect 15 5 16 8
rect 19 5 27 8
rect 30 5 31 8
rect 15 4 31 5
<< labels >>
rlabel m1 s 22 64 23 66 6 A
port 1 nsew signal input
rlabel m1 s 20 64 22 66 6 A
port 1 nsew signal input
rlabel m1 s 19 63 23 64 6 A
port 1 nsew signal input
rlabel m1 s 19 64 20 66 6 A
port 1 nsew signal input
rlabel m1 s 19 66 23 67 6 A
port 1 nsew signal input
rlabel m1 s 14 57 15 59 6 B
port 2 nsew signal input
rlabel m1 s 12 57 14 59 6 B
port 2 nsew signal input
rlabel m1 s 11 56 15 57 6 B
port 2 nsew signal input
rlabel m1 s 11 57 12 59 6 B
port 2 nsew signal input
rlabel m1 s 11 59 15 60 6 B
port 2 nsew signal input
rlabel m1 s 38 41 39 43 6 Y
port 3 nsew signal output
rlabel m1 s 38 18 39 20 6 Y
port 3 nsew signal output
rlabel m1 s 36 41 38 43 6 Y
port 3 nsew signal output
rlabel m1 s 36 18 38 20 6 Y
port 3 nsew signal output
rlabel m1 s 35 41 36 43 6 Y
port 3 nsew signal output
rlabel m1 s 35 18 36 20 6 Y
port 3 nsew signal output
rlabel m1 s 35 20 39 21 6 Y
port 3 nsew signal output
rlabel m1 s 35 40 39 41 6 Y
port 3 nsew signal output
rlabel m1 s 35 43 39 44 6 Y
port 3 nsew signal output
rlabel m1 s 36 21 39 40 6 Y
port 3 nsew signal output
rlabel m1 s 35 17 39 18 6 Y
port 3 nsew signal output
rlabel m1 s 26 41 27 43 6 Vdd
port 4 nsew power input
rlabel m1 s 24 41 26 43 6 Vdd
port 4 nsew power input
rlabel m1 s 24 44 27 60 6 Vdd
port 4 nsew power input
rlabel m1 s 23 40 27 41 6 Vdd
port 4 nsew power input
rlabel m1 s 23 41 24 43 6 Vdd
port 4 nsew power input
rlabel m1 s 23 43 27 44 6 Vdd
port 4 nsew power input
rlabel m2 s 26 18 27 21 6 GND
port 5 nsew ground input
rlabel m2 s 23 18 26 21 6 GND
port 5 nsew ground input
rlabel m2 s 9 18 23 21 6 GND
port 5 nsew ground input
rlabel m2 s 6 18 9 21 6 GND
port 5 nsew ground input
rlabel m2 s 5 17 27 18 6 GND
port 5 nsew ground input
rlabel m2 s 5 18 6 21 6 GND
port 5 nsew ground input
rlabel m2 s 5 21 27 22 6 GND
port 5 nsew ground input
rlabel m2c s 23 18 26 21 6 GND
port 5 nsew ground input
rlabel m2c s 6 18 9 21 6 GND
port 5 nsew ground input
rlabel m1 s 26 18 27 21 6 GND
port 5 nsew ground input
rlabel m1 s 23 18 26 21 6 GND
port 5 nsew ground input
rlabel m1 s 22 18 23 21 6 GND
port 5 nsew ground input
rlabel m1 s 22 21 27 22 6 GND
port 5 nsew ground input
rlabel m1 s 22 17 27 18 6 GND
port 5 nsew ground input
rlabel m1 s 9 18 10 21 6 GND
port 5 nsew ground input
rlabel m1 s 6 18 9 21 6 GND
port 5 nsew ground input
rlabel m1 s 5 17 10 18 6 GND
port 5 nsew ground input
rlabel m1 s 5 18 6 21 6 GND
port 5 nsew ground input
rlabel m1 s 5 21 10 22 6 GND
port 5 nsew ground input
rlabel space 0 0 54 70 1 prboundary
rlabel ndiffusion 31 18 31 18 3 Y
rlabel ndiffusion 31 19 31 19 3 Y
rlabel ndiffusion 31 21 31 21 3 Y
rlabel pdiffusion 31 39 31 39 3 Y
rlabel pdiffusion 31 42 31 42 3 Y
rlabel pdiffusion 31 44 31 44 3 Y
rlabel polysilicon 29 47 29 47 3 _Y
rlabel ntransistor 29 18 29 18 3 _Y
rlabel polysilicon 29 23 29 23 3 _Y
rlabel ptransistor 29 39 29 39 3 _Y
rlabel polysilicon 21 54 21 54 3 A
rlabel pdiffusion 23 39 23 39 3 Vdd
rlabel pdiffusion 23 42 23 42 3 Vdd
rlabel pdiffusion 23 44 23 44 3 Vdd
rlabel pdiffusion 23 47 23 47 3 Vdd
rlabel polysilicon 29 10 29 10 3 _Y
rlabel polysilicon 21 15 21 15 3 A
rlabel ntransistor 21 18 21 18 3 A
rlabel polysilicon 21 23 21 23 3 A
rlabel ptransistor 21 39 21 39 3 A
rlabel polysilicon 13 54 13 54 3 B
rlabel polysilicon 13 15 13 15 3 B
rlabel ntransistor 13 18 13 18 3 B
rlabel polysilicon 13 23 13 23 3 B
rlabel ptransistor 13 39 13 39 3 B
rlabel ndiffusion 4 18 4 18 3 GND
rlabel ndiffusion 4 19 4 19 3 GND
rlabel ndiffusion 4 22 4 22 3 GND
rlabel pdiffusion 4 39 4 39 3 _Y
rlabel pdiffusion 4 42 4 42 3 _Y
rlabel pdiffusion 4 45 4 45 3 _Y
rlabel m1 39 42 39 42 3 Y
port 3 e default output
rlabel m1 39 19 39 19 3 Y
port 3 e default output
rlabel pdcontact 37 42 37 42 3 Y
port 3 e default output
rlabel ndcontact 37 19 37 19 3 Y
port 3 e default output
rlabel m1 36 42 36 42 3 Y
port 3 e default output
rlabel m1 36 19 36 19 3 Y
port 3 e default output
rlabel m1 36 21 36 21 3 Y
port 3 e default output
rlabel m1 36 41 36 41 3 Y
port 3 e default output
rlabel m1 27 42 27 42 3 Vdd
rlabel m1 36 44 36 44 3 Y
port 3 e default output
rlabel m1 37 22 37 22 3 Y
port 3 e
rlabel pdcontact 25 42 25 42 3 Vdd
rlabel m1 25 45 25 45 3 Vdd
rlabel m1 24 41 24 41 3 Vdd
rlabel m1 24 42 24 42 3 Vdd
rlabel m1 24 44 24 44 3 Vdd
rlabel m1 23 19 23 19 3 GND
rlabel m1 23 22 23 22 3 GND
rlabel m1 23 65 23 65 3 A
port 1 e default input
rlabel polycontact 21 65 21 65 3 A
port 1 e
rlabel m1 20 64 20 64 3 A
port 1 e
rlabel m1 20 65 20 65 3 A
port 1 e
rlabel m1 20 67 20 67 3 A
port 1 e
rlabel m1 19 19 19 19 3 _Y
rlabel ndcontact 16 19 16 19 3 _Y
rlabel m1 16 23 16 23 3 _Y
rlabel m1 27 6 27 6 3 _Y
rlabel m1 36 18 36 18 3 Y
port 3 e
rlabel m1 15 19 15 19 3 _Y
rlabel m1 15 22 15 22 3 _Y
rlabel m1 15 30 15 30 3 _Y
rlabel m1 15 31 15 31 3 _Y
rlabel m1 15 34 15 34 3 _Y
rlabel m1 27 5 27 5 3 _Y
rlabel m1 27 9 27 9 3 _Y
rlabel m1 23 18 23 18 3 GND
rlabel m1 15 58 15 58 3 B
port 2 e default input
rlabel polycontact 13 58 13 58 3 B
port 2 e
rlabel m1 16 10 16 10 3 _Y
rlabel m1 15 18 15 18 3 _Y
rlabel m1 12 57 12 57 3 B
port 2 e
rlabel m1 12 58 12 58 3 B
port 2 e
rlabel m1 12 60 12 60 3 B
port 2 e
rlabel m1 9 42 9 42 3 _Y
rlabel m1 6 35 6 35 3 _Y
rlabel pdcontact 6 42 6 42 3 _Y
rlabel m1 5 41 5 41 3 _Y
rlabel m1 5 42 5 42 3 _Y
rlabel m1 5 45 5 45 3 _Y
rlabel m2 31 6 31 6 3 _Y
rlabel m2c 28 6 28 6 3 _Y
rlabel m2 20 6 20 6 3 _Y
rlabel m2 27 19 27 19 3 GND
rlabel m2c 17 6 17 6 3 _Y
rlabel m2c 24 19 24 19 3 GND
rlabel m2 19 31 19 31 3 _Y
rlabel m2 16 5 16 5 3 _Y
rlabel m2 16 6 16 6 3 _Y
rlabel m2 16 9 16 9 3 _Y
rlabel m2 10 19 10 19 3 GND
rlabel m2c 16 31 16 31 3 _Y
rlabel m2c 7 19 7 19 3 GND
rlabel m2 9 31 9 31 3 _Y
rlabel m2 6 18 6 18 3 GND
rlabel m2 6 19 6 19 3 GND
rlabel m2 6 22 6 22 3 GND
rlabel m2c 6 31 6 31 3 _Y
rlabel m2 5 30 5 30 3 _Y
rlabel m2 5 31 5 31 3 _Y
rlabel m2 5 34 5 34 3 _Y
<< properties >>
string FIXED_BBOX 0 0 54 70
string LEFclass CORE
string LEFsite CoreSite
string LEFsymmetry X Y
string LEFview TRUE
<< end >>
