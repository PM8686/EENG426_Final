magic
tech sky130l
timestamp 1729295985
<< ndiffusion >>
rect -1 10 13 12
rect -1 7 2 10
rect 5 7 13 10
rect -1 6 13 7
rect 15 6 20 12
rect 22 11 42 12
rect 22 8 26 11
rect 29 8 42 11
rect 22 6 42 8
<< ndc >>
rect 2 7 5 10
rect 26 8 29 11
<< ntransistor >>
rect 13 6 15 12
rect 20 6 22 12
<< pdiffusion >>
rect -1 19 13 34
rect 15 19 20 34
rect 22 24 42 34
rect 22 21 34 24
rect 37 21 42 24
rect 22 19 42 21
<< pdc >>
rect 34 21 37 24
<< ptransistor >>
rect 13 19 15 34
rect 20 19 22 34
<< polysilicon >>
rect 10 41 15 42
rect 10 38 11 41
rect 14 38 15 41
rect 10 37 15 38
rect 18 41 23 42
rect 18 38 19 41
rect 22 38 23 41
rect 18 37 23 38
rect 13 34 15 37
rect 20 34 22 37
rect 13 12 15 19
rect 20 12 22 19
rect 13 4 15 6
rect 20 4 22 6
<< pc >>
rect 11 38 14 41
rect 19 38 22 41
<< m1 >>
rect 10 41 15 42
rect 10 38 11 41
rect 14 38 15 41
rect 10 37 15 38
rect 18 41 23 42
rect 18 38 19 41
rect 22 38 23 41
rect 18 37 23 38
rect 26 36 30 40
rect 34 36 38 40
rect 8 28 12 29
rect 8 25 9 28
rect 16 28 20 29
rect 19 25 20 28
rect 8 24 12 25
rect 2 10 5 11
rect 9 8 12 24
rect 2 2 5 7
rect 8 4 12 8
rect 26 11 29 36
rect 34 24 37 36
rect 34 20 37 21
rect 26 2 29 8
<< m2c >>
rect 9 25 12 28
rect 16 25 19 28
rect 2 -1 5 2
rect 26 -1 29 2
<< m2 >>
rect 8 28 20 29
rect 8 25 9 28
rect 12 26 16 28
rect 12 25 13 26
rect 8 24 13 25
rect 15 25 16 26
rect 19 25 20 28
rect 15 24 20 25
rect 1 2 6 3
rect 25 2 30 3
rect 1 -1 2 2
rect 5 -1 26 2
rect 29 -1 30 2
rect 1 -2 6 -1
rect 25 -2 30 -1
<< labels >>
rlabel ndiffusion 23 7 23 7 3 GND
rlabel pdiffusion 23 20 23 20 3 Y
rlabel polysilicon 21 13 21 13 3 B
rlabel polysilicon 21 18 21 18 3 B
rlabel ndiffusion 16 7 16 7 3 Y
rlabel polysilicon 14 13 14 13 3 A
rlabel polysilicon 14 18 14 18 3 A
rlabel ndiffusion 9 7 9 7 3 GND
rlabel pdiffusion 9 20 9 20 3 Vdd
rlabel m1 9 5 9 5 3 Y
port 4 e
rlabel m1 27 37 28 38 5 GND
rlabel m1 35 37 36 38 6 Vdd
rlabel pc 12 38 13 39 5 A
rlabel pc 19 38 20 39 5 B
rlabel ndc 3 8 4 9 3 Y
<< end >>
