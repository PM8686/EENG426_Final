magic
tech TSMC180
timestamp 1734136781
<< ndiffusion >>
rect 6 11 12 12
rect 6 9 7 11
rect 9 9 12 11
rect 14 11 20 12
rect 14 9 17 11
rect 19 9 20 11
rect 6 8 10 9
rect 16 8 20 9
<< ndcontact >>
rect 7 9 9 11
rect 17 9 19 11
<< ntransistor >>
rect 12 9 14 12
<< pdiffusion >>
rect 6 31 10 32
rect 16 31 20 32
rect 6 29 7 31
rect 9 29 12 31
rect 6 28 12 29
rect 14 29 17 31
rect 19 29 20 31
rect 14 28 20 29
<< pdcontact >>
rect 7 29 9 31
rect 17 29 19 31
<< ptransistor >>
rect 12 28 14 31
<< polysilicon >>
rect 12 31 14 34
rect 12 12 14 28
rect 12 6 14 9
rect 12 5 20 6
rect 12 3 17 5
rect 19 3 20 5
rect 12 2 20 3
<< polycontact >>
rect 17 3 19 5
<< m1 >>
rect 6 32 9 40
rect 6 31 10 32
rect 6 29 7 31
rect 9 29 10 31
rect 6 28 10 29
rect 16 31 20 32
rect 24 31 27 40
rect 16 29 17 31
rect 19 29 27 31
rect 16 28 27 29
rect 6 12 9 13
rect 6 11 10 12
rect 6 9 7 11
rect 9 9 10 11
rect 6 8 10 9
rect 16 11 20 12
rect 16 9 17 11
rect 19 9 20 11
rect 16 5 20 9
rect 16 3 17 5
rect 19 3 20 5
rect 16 2 20 3
<< labels >>
rlabel ndiffusion 15 10 15 10 3 x
rlabel pdiffusion 15 29 15 29 3 Y
rlabel polysilicon 13 13 13 13 3 x
rlabel polysilicon 13 26 13 26 3 x
rlabel ndiffusion 7 10 7 10 3 GND
rlabel pdiffusion 7 29 7 29 3 Vdd
rlabel m1 7 38 7 38 3 Vdd
port 3 e
rlabel m1 7 11 7 11 2 GND
rlabel m1 25 38 25 38 6 Y
<< end >>
